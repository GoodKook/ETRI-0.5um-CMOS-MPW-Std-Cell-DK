magic
tech scmos
magscale 1 2
timestamp 0
<< metal1 >>
<< metal1 >>
rect 178 5 179 6
rect 161 5 162 6
rect 178 6 179 7
rect 177 6 178 7
rect 162 6 163 7
rect 161 6 162 7
rect 178 7 179 8
rect 177 7 178 8
rect 176 7 177 8
rect 175 7 176 8
rect 174 7 175 8
rect 173 7 174 8
rect 172 7 173 8
rect 171 7 172 8
rect 170 7 171 8
rect 169 7 170 8
rect 168 7 169 8
rect 167 7 168 8
rect 166 7 167 8
rect 165 7 166 8
rect 164 7 165 8
rect 163 7 164 8
rect 162 7 163 8
rect 161 7 162 8
rect 178 8 179 9
rect 177 8 178 9
rect 176 8 177 9
rect 175 8 176 9
rect 174 8 175 9
rect 173 8 174 9
rect 172 8 173 9
rect 171 8 172 9
rect 170 8 171 9
rect 169 8 170 9
rect 168 8 169 9
rect 167 8 168 9
rect 166 8 167 9
rect 165 8 166 9
rect 164 8 165 9
rect 163 8 164 9
rect 162 8 163 9
rect 161 8 162 9
rect 178 9 179 10
rect 177 9 178 10
rect 176 9 177 10
rect 175 9 176 10
rect 174 9 175 10
rect 173 9 174 10
rect 172 9 173 10
rect 171 9 172 10
rect 170 9 171 10
rect 169 9 170 10
rect 168 9 169 10
rect 167 9 168 10
rect 166 9 167 10
rect 165 9 166 10
rect 164 9 165 10
rect 163 9 164 10
rect 162 9 163 10
rect 161 9 162 10
rect 178 10 179 11
rect 177 10 178 11
rect 176 10 177 11
rect 175 10 176 11
rect 174 10 175 11
rect 173 10 174 11
rect 172 10 173 11
rect 171 10 172 11
rect 170 10 171 11
rect 169 10 170 11
rect 168 10 169 11
rect 167 10 168 11
rect 166 10 167 11
rect 165 10 166 11
rect 164 10 165 11
rect 163 10 164 11
rect 162 10 163 11
rect 161 10 162 11
rect 178 11 179 12
rect 177 11 178 12
rect 170 11 171 12
rect 169 11 170 12
rect 162 11 163 12
rect 161 11 162 12
rect 178 12 179 13
rect 171 12 172 13
rect 170 12 171 13
rect 169 12 170 13
rect 168 12 169 13
rect 161 12 162 13
rect 173 13 174 14
rect 172 13 173 14
rect 171 13 172 14
rect 170 13 171 14
rect 169 13 170 14
rect 168 13 169 14
rect 167 13 168 14
rect 174 14 175 15
rect 173 14 174 15
rect 172 14 173 15
rect 171 14 172 15
rect 170 14 171 15
rect 169 14 170 15
rect 168 14 169 15
rect 167 14 168 15
rect 166 14 167 15
rect 176 15 177 16
rect 175 15 176 16
rect 174 15 175 16
rect 173 15 174 16
rect 172 15 173 16
rect 171 15 172 16
rect 170 15 171 16
rect 169 15 170 16
rect 166 15 167 16
rect 165 15 166 16
rect 161 15 162 16
rect 177 16 178 17
rect 176 16 177 17
rect 175 16 176 17
rect 174 16 175 17
rect 173 16 174 17
rect 172 16 173 17
rect 171 16 172 17
rect 165 16 166 17
rect 164 16 165 17
rect 163 16 164 17
rect 161 16 162 17
rect 178 17 179 18
rect 177 17 178 18
rect 176 17 177 18
rect 175 17 176 18
rect 174 17 175 18
rect 173 17 174 18
rect 172 17 173 18
rect 164 17 165 18
rect 163 17 164 18
rect 162 17 163 18
rect 161 17 162 18
rect 178 18 179 19
rect 177 18 178 19
rect 176 18 177 19
rect 175 18 176 19
rect 174 18 175 19
rect 163 18 164 19
rect 162 18 163 19
rect 161 18 162 19
rect 178 19 179 20
rect 177 19 178 20
rect 176 19 177 20
rect 175 19 176 20
rect 162 19 163 20
rect 161 19 162 20
rect 178 20 179 21
rect 177 20 178 21
rect 176 20 177 21
rect 162 20 163 21
rect 161 20 162 21
rect 178 21 179 22
rect 177 21 178 22
rect 161 21 162 22
rect 178 22 179 23
rect 161 22 162 23
rect 39 23 40 24
rect 38 23 39 24
rect 41 24 42 25
rect 40 24 41 25
rect 39 24 40 25
rect 38 24 39 25
rect 37 24 38 25
rect 36 24 37 25
rect 161 25 162 26
rect 41 25 42 26
rect 40 25 41 26
rect 39 25 40 26
rect 38 25 39 26
rect 37 25 38 26
rect 36 25 37 26
rect 35 25 36 26
rect 162 26 163 27
rect 161 26 162 27
rect 46 26 47 27
rect 45 26 46 27
rect 41 26 42 27
rect 40 26 41 27
rect 39 26 40 27
rect 38 26 39 27
rect 37 26 38 27
rect 36 26 37 27
rect 35 26 36 27
rect 34 26 35 27
rect 163 27 164 28
rect 162 27 163 28
rect 161 27 162 28
rect 48 27 49 28
rect 47 27 48 28
rect 46 27 47 28
rect 45 27 46 28
rect 44 27 45 28
rect 41 27 42 28
rect 40 27 41 28
rect 39 27 40 28
rect 38 27 39 28
rect 37 27 38 28
rect 36 27 37 28
rect 35 27 36 28
rect 34 27 35 28
rect 165 28 166 29
rect 164 28 165 29
rect 163 28 164 29
rect 162 28 163 29
rect 161 28 162 29
rect 50 28 51 29
rect 49 28 50 29
rect 48 28 49 29
rect 47 28 48 29
rect 46 28 47 29
rect 45 28 46 29
rect 44 28 45 29
rect 43 28 44 29
rect 40 28 41 29
rect 39 28 40 29
rect 38 28 39 29
rect 37 28 38 29
rect 36 28 37 29
rect 35 28 36 29
rect 34 28 35 29
rect 33 28 34 29
rect 178 29 179 30
rect 167 29 168 30
rect 166 29 167 30
rect 165 29 166 30
rect 164 29 165 30
rect 163 29 164 30
rect 162 29 163 30
rect 161 29 162 30
rect 51 29 52 30
rect 50 29 51 30
rect 49 29 50 30
rect 48 29 49 30
rect 47 29 48 30
rect 46 29 47 30
rect 45 29 46 30
rect 44 29 45 30
rect 43 29 44 30
rect 42 29 43 30
rect 40 29 41 30
rect 39 29 40 30
rect 38 29 39 30
rect 37 29 38 30
rect 36 29 37 30
rect 35 29 36 30
rect 34 29 35 30
rect 33 29 34 30
rect 178 30 179 31
rect 169 30 170 31
rect 168 30 169 31
rect 167 30 168 31
rect 166 30 167 31
rect 165 30 166 31
rect 164 30 165 31
rect 163 30 164 31
rect 162 30 163 31
rect 161 30 162 31
rect 52 30 53 31
rect 51 30 52 31
rect 50 30 51 31
rect 49 30 50 31
rect 48 30 49 31
rect 47 30 48 31
rect 46 30 47 31
rect 45 30 46 31
rect 44 30 45 31
rect 43 30 44 31
rect 42 30 43 31
rect 41 30 42 31
rect 39 30 40 31
rect 38 30 39 31
rect 37 30 38 31
rect 36 30 37 31
rect 35 30 36 31
rect 34 30 35 31
rect 33 30 34 31
rect 32 30 33 31
rect 178 31 179 32
rect 177 31 178 32
rect 176 31 177 32
rect 175 31 176 32
rect 174 31 175 32
rect 173 31 174 32
rect 172 31 173 32
rect 171 31 172 32
rect 170 31 171 32
rect 169 31 170 32
rect 168 31 169 32
rect 167 31 168 32
rect 166 31 167 32
rect 165 31 166 32
rect 164 31 165 32
rect 163 31 164 32
rect 162 31 163 32
rect 161 31 162 32
rect 52 31 53 32
rect 51 31 52 32
rect 50 31 51 32
rect 49 31 50 32
rect 48 31 49 32
rect 47 31 48 32
rect 46 31 47 32
rect 45 31 46 32
rect 44 31 45 32
rect 43 31 44 32
rect 42 31 43 32
rect 41 31 42 32
rect 40 31 41 32
rect 39 31 40 32
rect 38 31 39 32
rect 37 31 38 32
rect 36 31 37 32
rect 35 31 36 32
rect 34 31 35 32
rect 33 31 34 32
rect 32 31 33 32
rect 178 32 179 33
rect 177 32 178 33
rect 176 32 177 33
rect 175 32 176 33
rect 174 32 175 33
rect 173 32 174 33
rect 172 32 173 33
rect 171 32 172 33
rect 170 32 171 33
rect 169 32 170 33
rect 168 32 169 33
rect 167 32 168 33
rect 166 32 167 33
rect 165 32 166 33
rect 161 32 162 33
rect 59 32 60 33
rect 58 32 59 33
rect 57 32 58 33
rect 56 32 57 33
rect 53 32 54 33
rect 52 32 53 33
rect 51 32 52 33
rect 50 32 51 33
rect 49 32 50 33
rect 48 32 49 33
rect 47 32 48 33
rect 46 32 47 33
rect 45 32 46 33
rect 44 32 45 33
rect 43 32 44 33
rect 42 32 43 33
rect 41 32 42 33
rect 40 32 41 33
rect 39 32 40 33
rect 38 32 39 33
rect 37 32 38 33
rect 36 32 37 33
rect 35 32 36 33
rect 34 32 35 33
rect 33 32 34 33
rect 32 32 33 33
rect 31 32 32 33
rect 178 33 179 34
rect 177 33 178 34
rect 176 33 177 34
rect 175 33 176 34
rect 174 33 175 34
rect 173 33 174 34
rect 172 33 173 34
rect 171 33 172 34
rect 170 33 171 34
rect 169 33 170 34
rect 168 33 169 34
rect 167 33 168 34
rect 61 33 62 34
rect 60 33 61 34
rect 59 33 60 34
rect 58 33 59 34
rect 57 33 58 34
rect 56 33 57 34
rect 53 33 54 34
rect 52 33 53 34
rect 51 33 52 34
rect 50 33 51 34
rect 49 33 50 34
rect 48 33 49 34
rect 47 33 48 34
rect 46 33 47 34
rect 45 33 46 34
rect 44 33 45 34
rect 43 33 44 34
rect 42 33 43 34
rect 41 33 42 34
rect 40 33 41 34
rect 39 33 40 34
rect 38 33 39 34
rect 37 33 38 34
rect 36 33 37 34
rect 35 33 36 34
rect 34 33 35 34
rect 33 33 34 34
rect 32 33 33 34
rect 31 33 32 34
rect 178 34 179 35
rect 177 34 178 35
rect 176 34 177 35
rect 175 34 176 35
rect 174 34 175 35
rect 173 34 174 35
rect 172 34 173 35
rect 171 34 172 35
rect 170 34 171 35
rect 169 34 170 35
rect 63 34 64 35
rect 62 34 63 35
rect 61 34 62 35
rect 60 34 61 35
rect 59 34 60 35
rect 58 34 59 35
rect 57 34 58 35
rect 56 34 57 35
rect 53 34 54 35
rect 52 34 53 35
rect 51 34 52 35
rect 50 34 51 35
rect 49 34 50 35
rect 48 34 49 35
rect 47 34 48 35
rect 46 34 47 35
rect 45 34 46 35
rect 44 34 45 35
rect 43 34 44 35
rect 42 34 43 35
rect 41 34 42 35
rect 40 34 41 35
rect 39 34 40 35
rect 38 34 39 35
rect 37 34 38 35
rect 36 34 37 35
rect 35 34 36 35
rect 34 34 35 35
rect 33 34 34 35
rect 32 34 33 35
rect 31 34 32 35
rect 30 34 31 35
rect 178 35 179 36
rect 177 35 178 36
rect 176 35 177 36
rect 175 35 176 36
rect 174 35 175 36
rect 173 35 174 36
rect 172 35 173 36
rect 171 35 172 36
rect 170 35 171 36
rect 169 35 170 36
rect 168 35 169 36
rect 167 35 168 36
rect 65 35 66 36
rect 64 35 65 36
rect 63 35 64 36
rect 62 35 63 36
rect 61 35 62 36
rect 60 35 61 36
rect 59 35 60 36
rect 58 35 59 36
rect 57 35 58 36
rect 56 35 57 36
rect 53 35 54 36
rect 52 35 53 36
rect 51 35 52 36
rect 50 35 51 36
rect 49 35 50 36
rect 48 35 49 36
rect 47 35 48 36
rect 46 35 47 36
rect 45 35 46 36
rect 44 35 45 36
rect 43 35 44 36
rect 42 35 43 36
rect 41 35 42 36
rect 40 35 41 36
rect 39 35 40 36
rect 38 35 39 36
rect 37 35 38 36
rect 36 35 37 36
rect 35 35 36 36
rect 34 35 35 36
rect 33 35 34 36
rect 32 35 33 36
rect 31 35 32 36
rect 30 35 31 36
rect 178 36 179 37
rect 168 36 169 37
rect 167 36 168 37
rect 166 36 167 37
rect 165 36 166 37
rect 161 36 162 37
rect 67 36 68 37
rect 66 36 67 37
rect 65 36 66 37
rect 64 36 65 37
rect 63 36 64 37
rect 62 36 63 37
rect 61 36 62 37
rect 60 36 61 37
rect 59 36 60 37
rect 58 36 59 37
rect 57 36 58 37
rect 56 36 57 37
rect 53 36 54 37
rect 52 36 53 37
rect 51 36 52 37
rect 50 36 51 37
rect 49 36 50 37
rect 48 36 49 37
rect 47 36 48 37
rect 46 36 47 37
rect 45 36 46 37
rect 44 36 45 37
rect 43 36 44 37
rect 42 36 43 37
rect 41 36 42 37
rect 40 36 41 37
rect 39 36 40 37
rect 38 36 39 37
rect 37 36 38 37
rect 36 36 37 37
rect 35 36 36 37
rect 34 36 35 37
rect 33 36 34 37
rect 32 36 33 37
rect 31 36 32 37
rect 30 36 31 37
rect 29 36 30 37
rect 193 37 194 38
rect 192 37 193 38
rect 191 37 192 38
rect 190 37 191 38
rect 189 37 190 38
rect 188 37 189 38
rect 187 37 188 38
rect 178 37 179 38
rect 166 37 167 38
rect 165 37 166 38
rect 164 37 165 38
rect 163 37 164 38
rect 162 37 163 38
rect 161 37 162 38
rect 95 37 96 38
rect 94 37 95 38
rect 93 37 94 38
rect 92 37 93 38
rect 91 37 92 38
rect 90 37 91 38
rect 89 37 90 38
rect 88 37 89 38
rect 87 37 88 38
rect 86 37 87 38
rect 85 37 86 38
rect 68 37 69 38
rect 67 37 68 38
rect 66 37 67 38
rect 65 37 66 38
rect 64 37 65 38
rect 63 37 64 38
rect 62 37 63 38
rect 61 37 62 38
rect 60 37 61 38
rect 59 37 60 38
rect 58 37 59 38
rect 57 37 58 38
rect 56 37 57 38
rect 55 37 56 38
rect 52 37 53 38
rect 51 37 52 38
rect 50 37 51 38
rect 49 37 50 38
rect 48 37 49 38
rect 47 37 48 38
rect 46 37 47 38
rect 45 37 46 38
rect 44 37 45 38
rect 43 37 44 38
rect 42 37 43 38
rect 41 37 42 38
rect 40 37 41 38
rect 39 37 40 38
rect 38 37 39 38
rect 37 37 38 38
rect 36 37 37 38
rect 35 37 36 38
rect 34 37 35 38
rect 33 37 34 38
rect 32 37 33 38
rect 31 37 32 38
rect 30 37 31 38
rect 29 37 30 38
rect 28 37 29 38
rect 194 38 195 39
rect 193 38 194 39
rect 192 38 193 39
rect 191 38 192 39
rect 190 38 191 39
rect 189 38 190 39
rect 188 38 189 39
rect 187 38 188 39
rect 164 38 165 39
rect 163 38 164 39
rect 162 38 163 39
rect 161 38 162 39
rect 99 38 100 39
rect 98 38 99 39
rect 97 38 98 39
rect 96 38 97 39
rect 95 38 96 39
rect 94 38 95 39
rect 93 38 94 39
rect 92 38 93 39
rect 91 38 92 39
rect 90 38 91 39
rect 89 38 90 39
rect 88 38 89 39
rect 87 38 88 39
rect 86 38 87 39
rect 85 38 86 39
rect 84 38 85 39
rect 83 38 84 39
rect 82 38 83 39
rect 68 38 69 39
rect 67 38 68 39
rect 66 38 67 39
rect 65 38 66 39
rect 64 38 65 39
rect 63 38 64 39
rect 62 38 63 39
rect 61 38 62 39
rect 60 38 61 39
rect 59 38 60 39
rect 58 38 59 39
rect 57 38 58 39
rect 56 38 57 39
rect 55 38 56 39
rect 52 38 53 39
rect 51 38 52 39
rect 50 38 51 39
rect 49 38 50 39
rect 48 38 49 39
rect 47 38 48 39
rect 46 38 47 39
rect 45 38 46 39
rect 44 38 45 39
rect 43 38 44 39
rect 42 38 43 39
rect 41 38 42 39
rect 40 38 41 39
rect 39 38 40 39
rect 38 38 39 39
rect 37 38 38 39
rect 36 38 37 39
rect 35 38 36 39
rect 34 38 35 39
rect 33 38 34 39
rect 32 38 33 39
rect 31 38 32 39
rect 30 38 31 39
rect 29 38 30 39
rect 28 38 29 39
rect 195 39 196 40
rect 194 39 195 40
rect 193 39 194 40
rect 187 39 188 40
rect 163 39 164 40
rect 162 39 163 40
rect 161 39 162 40
rect 101 39 102 40
rect 100 39 101 40
rect 99 39 100 40
rect 98 39 99 40
rect 97 39 98 40
rect 96 39 97 40
rect 95 39 96 40
rect 94 39 95 40
rect 93 39 94 40
rect 92 39 93 40
rect 91 39 92 40
rect 90 39 91 40
rect 89 39 90 40
rect 88 39 89 40
rect 87 39 88 40
rect 86 39 87 40
rect 85 39 86 40
rect 84 39 85 40
rect 83 39 84 40
rect 82 39 83 40
rect 81 39 82 40
rect 80 39 81 40
rect 68 39 69 40
rect 67 39 68 40
rect 66 39 67 40
rect 65 39 66 40
rect 64 39 65 40
rect 63 39 64 40
rect 62 39 63 40
rect 61 39 62 40
rect 60 39 61 40
rect 59 39 60 40
rect 58 39 59 40
rect 57 39 58 40
rect 56 39 57 40
rect 55 39 56 40
rect 52 39 53 40
rect 51 39 52 40
rect 50 39 51 40
rect 49 39 50 40
rect 48 39 49 40
rect 47 39 48 40
rect 46 39 47 40
rect 45 39 46 40
rect 44 39 45 40
rect 43 39 44 40
rect 42 39 43 40
rect 41 39 42 40
rect 40 39 41 40
rect 39 39 40 40
rect 38 39 39 40
rect 37 39 38 40
rect 36 39 37 40
rect 35 39 36 40
rect 34 39 35 40
rect 33 39 34 40
rect 32 39 33 40
rect 31 39 32 40
rect 30 39 31 40
rect 29 39 30 40
rect 28 39 29 40
rect 27 39 28 40
rect 195 40 196 41
rect 194 40 195 41
rect 162 40 163 41
rect 161 40 162 41
rect 103 40 104 41
rect 102 40 103 41
rect 101 40 102 41
rect 100 40 101 41
rect 99 40 100 41
rect 98 40 99 41
rect 97 40 98 41
rect 96 40 97 41
rect 95 40 96 41
rect 94 40 95 41
rect 93 40 94 41
rect 92 40 93 41
rect 91 40 92 41
rect 90 40 91 41
rect 89 40 90 41
rect 88 40 89 41
rect 87 40 88 41
rect 86 40 87 41
rect 85 40 86 41
rect 84 40 85 41
rect 83 40 84 41
rect 82 40 83 41
rect 81 40 82 41
rect 80 40 81 41
rect 79 40 80 41
rect 78 40 79 41
rect 67 40 68 41
rect 66 40 67 41
rect 65 40 66 41
rect 64 40 65 41
rect 63 40 64 41
rect 62 40 63 41
rect 61 40 62 41
rect 60 40 61 41
rect 59 40 60 41
rect 58 40 59 41
rect 57 40 58 41
rect 56 40 57 41
rect 55 40 56 41
rect 52 40 53 41
rect 51 40 52 41
rect 50 40 51 41
rect 49 40 50 41
rect 48 40 49 41
rect 47 40 48 41
rect 46 40 47 41
rect 45 40 46 41
rect 44 40 45 41
rect 43 40 44 41
rect 42 40 43 41
rect 41 40 42 41
rect 40 40 41 41
rect 39 40 40 41
rect 38 40 39 41
rect 37 40 38 41
rect 36 40 37 41
rect 35 40 36 41
rect 34 40 35 41
rect 33 40 34 41
rect 32 40 33 41
rect 31 40 32 41
rect 30 40 31 41
rect 29 40 30 41
rect 28 40 29 41
rect 27 40 28 41
rect 26 40 27 41
rect 195 41 196 42
rect 161 41 162 42
rect 105 41 106 42
rect 104 41 105 42
rect 103 41 104 42
rect 102 41 103 42
rect 101 41 102 42
rect 100 41 101 42
rect 99 41 100 42
rect 98 41 99 42
rect 97 41 98 42
rect 96 41 97 42
rect 95 41 96 42
rect 94 41 95 42
rect 93 41 94 42
rect 92 41 93 42
rect 91 41 92 42
rect 90 41 91 42
rect 89 41 90 42
rect 88 41 89 42
rect 87 41 88 42
rect 86 41 87 42
rect 85 41 86 42
rect 84 41 85 42
rect 83 41 84 42
rect 82 41 83 42
rect 81 41 82 42
rect 80 41 81 42
rect 79 41 80 42
rect 78 41 79 42
rect 77 41 78 42
rect 67 41 68 42
rect 66 41 67 42
rect 65 41 66 42
rect 64 41 65 42
rect 63 41 64 42
rect 62 41 63 42
rect 61 41 62 42
rect 60 41 61 42
rect 59 41 60 42
rect 58 41 59 42
rect 57 41 58 42
rect 56 41 57 42
rect 55 41 56 42
rect 52 41 53 42
rect 51 41 52 42
rect 50 41 51 42
rect 49 41 50 42
rect 48 41 49 42
rect 47 41 48 42
rect 46 41 47 42
rect 45 41 46 42
rect 44 41 45 42
rect 43 41 44 42
rect 42 41 43 42
rect 41 41 42 42
rect 40 41 41 42
rect 39 41 40 42
rect 38 41 39 42
rect 37 41 38 42
rect 36 41 37 42
rect 35 41 36 42
rect 34 41 35 42
rect 33 41 34 42
rect 32 41 33 42
rect 31 41 32 42
rect 30 41 31 42
rect 29 41 30 42
rect 28 41 29 42
rect 27 41 28 42
rect 26 41 27 42
rect 195 42 196 43
rect 194 42 195 43
rect 107 42 108 43
rect 106 42 107 43
rect 105 42 106 43
rect 104 42 105 43
rect 103 42 104 43
rect 102 42 103 43
rect 101 42 102 43
rect 100 42 101 43
rect 99 42 100 43
rect 98 42 99 43
rect 97 42 98 43
rect 96 42 97 43
rect 95 42 96 43
rect 94 42 95 43
rect 93 42 94 43
rect 92 42 93 43
rect 91 42 92 43
rect 90 42 91 43
rect 89 42 90 43
rect 88 42 89 43
rect 87 42 88 43
rect 86 42 87 43
rect 85 42 86 43
rect 84 42 85 43
rect 83 42 84 43
rect 82 42 83 43
rect 81 42 82 43
rect 80 42 81 43
rect 79 42 80 43
rect 78 42 79 43
rect 77 42 78 43
rect 76 42 77 43
rect 67 42 68 43
rect 66 42 67 43
rect 65 42 66 43
rect 64 42 65 43
rect 63 42 64 43
rect 62 42 63 43
rect 61 42 62 43
rect 60 42 61 43
rect 59 42 60 43
rect 58 42 59 43
rect 57 42 58 43
rect 56 42 57 43
rect 55 42 56 43
rect 51 42 52 43
rect 50 42 51 43
rect 49 42 50 43
rect 48 42 49 43
rect 47 42 48 43
rect 46 42 47 43
rect 45 42 46 43
rect 44 42 45 43
rect 43 42 44 43
rect 42 42 43 43
rect 41 42 42 43
rect 40 42 41 43
rect 39 42 40 43
rect 38 42 39 43
rect 37 42 38 43
rect 36 42 37 43
rect 35 42 36 43
rect 34 42 35 43
rect 33 42 34 43
rect 32 42 33 43
rect 31 42 32 43
rect 30 42 31 43
rect 29 42 30 43
rect 28 42 29 43
rect 27 42 28 43
rect 26 42 27 43
rect 25 42 26 43
rect 194 43 195 44
rect 193 43 194 44
rect 192 43 193 44
rect 191 43 192 44
rect 190 43 191 44
rect 189 43 190 44
rect 188 43 189 44
rect 187 43 188 44
rect 108 43 109 44
rect 107 43 108 44
rect 106 43 107 44
rect 105 43 106 44
rect 104 43 105 44
rect 103 43 104 44
rect 102 43 103 44
rect 101 43 102 44
rect 100 43 101 44
rect 99 43 100 44
rect 98 43 99 44
rect 97 43 98 44
rect 96 43 97 44
rect 95 43 96 44
rect 94 43 95 44
rect 93 43 94 44
rect 92 43 93 44
rect 91 43 92 44
rect 90 43 91 44
rect 89 43 90 44
rect 88 43 89 44
rect 87 43 88 44
rect 86 43 87 44
rect 85 43 86 44
rect 84 43 85 44
rect 83 43 84 44
rect 82 43 83 44
rect 81 43 82 44
rect 80 43 81 44
rect 79 43 80 44
rect 78 43 79 44
rect 77 43 78 44
rect 76 43 77 44
rect 75 43 76 44
rect 66 43 67 44
rect 65 43 66 44
rect 64 43 65 44
rect 63 43 64 44
rect 62 43 63 44
rect 61 43 62 44
rect 60 43 61 44
rect 59 43 60 44
rect 58 43 59 44
rect 57 43 58 44
rect 56 43 57 44
rect 55 43 56 44
rect 54 43 55 44
rect 51 43 52 44
rect 50 43 51 44
rect 49 43 50 44
rect 48 43 49 44
rect 47 43 48 44
rect 46 43 47 44
rect 45 43 46 44
rect 44 43 45 44
rect 43 43 44 44
rect 42 43 43 44
rect 41 43 42 44
rect 40 43 41 44
rect 39 43 40 44
rect 38 43 39 44
rect 37 43 38 44
rect 36 43 37 44
rect 35 43 36 44
rect 34 43 35 44
rect 33 43 34 44
rect 31 43 32 44
rect 30 43 31 44
rect 29 43 30 44
rect 28 43 29 44
rect 27 43 28 44
rect 26 43 27 44
rect 25 43 26 44
rect 24 43 25 44
rect 188 44 189 45
rect 187 44 188 45
rect 161 44 162 45
rect 109 44 110 45
rect 108 44 109 45
rect 107 44 108 45
rect 106 44 107 45
rect 105 44 106 45
rect 104 44 105 45
rect 103 44 104 45
rect 102 44 103 45
rect 101 44 102 45
rect 100 44 101 45
rect 99 44 100 45
rect 98 44 99 45
rect 97 44 98 45
rect 96 44 97 45
rect 95 44 96 45
rect 94 44 95 45
rect 93 44 94 45
rect 92 44 93 45
rect 91 44 92 45
rect 90 44 91 45
rect 89 44 90 45
rect 88 44 89 45
rect 87 44 88 45
rect 86 44 87 45
rect 85 44 86 45
rect 84 44 85 45
rect 83 44 84 45
rect 82 44 83 45
rect 81 44 82 45
rect 80 44 81 45
rect 79 44 80 45
rect 78 44 79 45
rect 77 44 78 45
rect 76 44 77 45
rect 75 44 76 45
rect 74 44 75 45
rect 66 44 67 45
rect 65 44 66 45
rect 64 44 65 45
rect 63 44 64 45
rect 62 44 63 45
rect 61 44 62 45
rect 60 44 61 45
rect 59 44 60 45
rect 58 44 59 45
rect 57 44 58 45
rect 56 44 57 45
rect 55 44 56 45
rect 54 44 55 45
rect 50 44 51 45
rect 49 44 50 45
rect 48 44 49 45
rect 47 44 48 45
rect 46 44 47 45
rect 45 44 46 45
rect 44 44 45 45
rect 43 44 44 45
rect 42 44 43 45
rect 41 44 42 45
rect 40 44 41 45
rect 39 44 40 45
rect 38 44 39 45
rect 37 44 38 45
rect 36 44 37 45
rect 35 44 36 45
rect 34 44 35 45
rect 33 44 34 45
rect 30 44 31 45
rect 29 44 30 45
rect 28 44 29 45
rect 27 44 28 45
rect 26 44 27 45
rect 25 44 26 45
rect 24 44 25 45
rect 23 44 24 45
rect 161 45 162 46
rect 110 45 111 46
rect 109 45 110 46
rect 108 45 109 46
rect 107 45 108 46
rect 106 45 107 46
rect 105 45 106 46
rect 104 45 105 46
rect 103 45 104 46
rect 102 45 103 46
rect 101 45 102 46
rect 100 45 101 46
rect 99 45 100 46
rect 98 45 99 46
rect 97 45 98 46
rect 96 45 97 46
rect 95 45 96 46
rect 94 45 95 46
rect 93 45 94 46
rect 92 45 93 46
rect 91 45 92 46
rect 90 45 91 46
rect 89 45 90 46
rect 88 45 89 46
rect 87 45 88 46
rect 86 45 87 46
rect 85 45 86 46
rect 84 45 85 46
rect 83 45 84 46
rect 82 45 83 46
rect 81 45 82 46
rect 80 45 81 46
rect 79 45 80 46
rect 78 45 79 46
rect 77 45 78 46
rect 76 45 77 46
rect 75 45 76 46
rect 74 45 75 46
rect 66 45 67 46
rect 65 45 66 46
rect 64 45 65 46
rect 63 45 64 46
rect 62 45 63 46
rect 61 45 62 46
rect 60 45 61 46
rect 59 45 60 46
rect 58 45 59 46
rect 57 45 58 46
rect 56 45 57 46
rect 55 45 56 46
rect 54 45 55 46
rect 49 45 50 46
rect 48 45 49 46
rect 47 45 48 46
rect 46 45 47 46
rect 45 45 46 46
rect 44 45 45 46
rect 43 45 44 46
rect 42 45 43 46
rect 41 45 42 46
rect 40 45 41 46
rect 39 45 40 46
rect 38 45 39 46
rect 37 45 38 46
rect 36 45 37 46
rect 35 45 36 46
rect 34 45 35 46
rect 33 45 34 46
rect 30 45 31 46
rect 29 45 30 46
rect 28 45 29 46
rect 27 45 28 46
rect 26 45 27 46
rect 25 45 26 46
rect 24 45 25 46
rect 23 45 24 46
rect 22 45 23 46
rect 171 46 172 47
rect 170 46 171 47
rect 169 46 170 47
rect 168 46 169 47
rect 167 46 168 47
rect 166 46 167 47
rect 165 46 166 47
rect 164 46 165 47
rect 163 46 164 47
rect 162 46 163 47
rect 161 46 162 47
rect 111 46 112 47
rect 110 46 111 47
rect 109 46 110 47
rect 108 46 109 47
rect 107 46 108 47
rect 106 46 107 47
rect 105 46 106 47
rect 104 46 105 47
rect 103 46 104 47
rect 102 46 103 47
rect 101 46 102 47
rect 100 46 101 47
rect 99 46 100 47
rect 98 46 99 47
rect 97 46 98 47
rect 96 46 97 47
rect 95 46 96 47
rect 94 46 95 47
rect 93 46 94 47
rect 92 46 93 47
rect 91 46 92 47
rect 90 46 91 47
rect 89 46 90 47
rect 88 46 89 47
rect 87 46 88 47
rect 86 46 87 47
rect 85 46 86 47
rect 84 46 85 47
rect 83 46 84 47
rect 82 46 83 47
rect 81 46 82 47
rect 80 46 81 47
rect 79 46 80 47
rect 78 46 79 47
rect 77 46 78 47
rect 76 46 77 47
rect 75 46 76 47
rect 74 46 75 47
rect 73 46 74 47
rect 65 46 66 47
rect 64 46 65 47
rect 63 46 64 47
rect 62 46 63 47
rect 61 46 62 47
rect 60 46 61 47
rect 59 46 60 47
rect 58 46 59 47
rect 57 46 58 47
rect 56 46 57 47
rect 55 46 56 47
rect 54 46 55 47
rect 49 46 50 47
rect 48 46 49 47
rect 47 46 48 47
rect 46 46 47 47
rect 45 46 46 47
rect 44 46 45 47
rect 43 46 44 47
rect 42 46 43 47
rect 41 46 42 47
rect 40 46 41 47
rect 39 46 40 47
rect 38 46 39 47
rect 37 46 38 47
rect 36 46 37 47
rect 35 46 36 47
rect 34 46 35 47
rect 29 46 30 47
rect 28 46 29 47
rect 27 46 28 47
rect 26 46 27 47
rect 25 46 26 47
rect 24 46 25 47
rect 23 46 24 47
rect 22 46 23 47
rect 21 46 22 47
rect 20 46 21 47
rect 175 47 176 48
rect 174 47 175 48
rect 173 47 174 48
rect 172 47 173 48
rect 171 47 172 48
rect 170 47 171 48
rect 169 47 170 48
rect 168 47 169 48
rect 167 47 168 48
rect 166 47 167 48
rect 165 47 166 48
rect 164 47 165 48
rect 163 47 164 48
rect 162 47 163 48
rect 161 47 162 48
rect 112 47 113 48
rect 111 47 112 48
rect 110 47 111 48
rect 109 47 110 48
rect 108 47 109 48
rect 107 47 108 48
rect 106 47 107 48
rect 105 47 106 48
rect 104 47 105 48
rect 103 47 104 48
rect 102 47 103 48
rect 101 47 102 48
rect 100 47 101 48
rect 99 47 100 48
rect 98 47 99 48
rect 97 47 98 48
rect 96 47 97 48
rect 95 47 96 48
rect 94 47 95 48
rect 93 47 94 48
rect 92 47 93 48
rect 91 47 92 48
rect 90 47 91 48
rect 89 47 90 48
rect 88 47 89 48
rect 87 47 88 48
rect 86 47 87 48
rect 85 47 86 48
rect 84 47 85 48
rect 83 47 84 48
rect 82 47 83 48
rect 81 47 82 48
rect 80 47 81 48
rect 79 47 80 48
rect 78 47 79 48
rect 77 47 78 48
rect 76 47 77 48
rect 75 47 76 48
rect 74 47 75 48
rect 73 47 74 48
rect 65 47 66 48
rect 64 47 65 48
rect 63 47 64 48
rect 62 47 63 48
rect 61 47 62 48
rect 60 47 61 48
rect 59 47 60 48
rect 58 47 59 48
rect 57 47 58 48
rect 56 47 57 48
rect 55 47 56 48
rect 54 47 55 48
rect 53 47 54 48
rect 50 47 51 48
rect 49 47 50 48
rect 48 47 49 48
rect 47 47 48 48
rect 46 47 47 48
rect 45 47 46 48
rect 44 47 45 48
rect 43 47 44 48
rect 42 47 43 48
rect 41 47 42 48
rect 40 47 41 48
rect 39 47 40 48
rect 38 47 39 48
rect 37 47 38 48
rect 36 47 37 48
rect 29 47 30 48
rect 28 47 29 48
rect 27 47 28 48
rect 26 47 27 48
rect 25 47 26 48
rect 24 47 25 48
rect 23 47 24 48
rect 22 47 23 48
rect 21 47 22 48
rect 20 47 21 48
rect 19 47 20 48
rect 177 48 178 49
rect 176 48 177 49
rect 175 48 176 49
rect 174 48 175 49
rect 173 48 174 49
rect 172 48 173 49
rect 171 48 172 49
rect 170 48 171 49
rect 169 48 170 49
rect 168 48 169 49
rect 167 48 168 49
rect 166 48 167 49
rect 165 48 166 49
rect 164 48 165 49
rect 163 48 164 49
rect 162 48 163 49
rect 161 48 162 49
rect 113 48 114 49
rect 112 48 113 49
rect 111 48 112 49
rect 110 48 111 49
rect 109 48 110 49
rect 108 48 109 49
rect 107 48 108 49
rect 106 48 107 49
rect 105 48 106 49
rect 104 48 105 49
rect 103 48 104 49
rect 102 48 103 49
rect 101 48 102 49
rect 100 48 101 49
rect 99 48 100 49
rect 98 48 99 49
rect 97 48 98 49
rect 96 48 97 49
rect 95 48 96 49
rect 94 48 95 49
rect 93 48 94 49
rect 92 48 93 49
rect 91 48 92 49
rect 90 48 91 49
rect 89 48 90 49
rect 88 48 89 49
rect 87 48 88 49
rect 86 48 87 49
rect 85 48 86 49
rect 84 48 85 49
rect 83 48 84 49
rect 82 48 83 49
rect 81 48 82 49
rect 80 48 81 49
rect 79 48 80 49
rect 78 48 79 49
rect 77 48 78 49
rect 76 48 77 49
rect 75 48 76 49
rect 74 48 75 49
rect 73 48 74 49
rect 72 48 73 49
rect 65 48 66 49
rect 64 48 65 49
rect 63 48 64 49
rect 62 48 63 49
rect 61 48 62 49
rect 60 48 61 49
rect 59 48 60 49
rect 58 48 59 49
rect 57 48 58 49
rect 56 48 57 49
rect 55 48 56 49
rect 54 48 55 49
rect 53 48 54 49
rect 52 48 53 49
rect 51 48 52 49
rect 50 48 51 49
rect 49 48 50 49
rect 48 48 49 49
rect 47 48 48 49
rect 46 48 47 49
rect 45 48 46 49
rect 44 48 45 49
rect 43 48 44 49
rect 42 48 43 49
rect 41 48 42 49
rect 40 48 41 49
rect 39 48 40 49
rect 38 48 39 49
rect 37 48 38 49
rect 36 48 37 49
rect 35 48 36 49
rect 28 48 29 49
rect 27 48 28 49
rect 26 48 27 49
rect 25 48 26 49
rect 24 48 25 49
rect 23 48 24 49
rect 22 48 23 49
rect 21 48 22 49
rect 20 48 21 49
rect 19 48 20 49
rect 18 48 19 49
rect 17 48 18 49
rect 195 49 196 50
rect 194 49 195 50
rect 193 49 194 50
rect 192 49 193 50
rect 191 49 192 50
rect 190 49 191 50
rect 189 49 190 50
rect 188 49 189 50
rect 187 49 188 50
rect 178 49 179 50
rect 177 49 178 50
rect 176 49 177 50
rect 175 49 176 50
rect 174 49 175 50
rect 173 49 174 50
rect 172 49 173 50
rect 171 49 172 50
rect 170 49 171 50
rect 169 49 170 50
rect 168 49 169 50
rect 167 49 168 50
rect 166 49 167 50
rect 165 49 166 50
rect 164 49 165 50
rect 163 49 164 50
rect 162 49 163 50
rect 161 49 162 50
rect 108 49 109 50
rect 107 49 108 50
rect 106 49 107 50
rect 105 49 106 50
rect 104 49 105 50
rect 103 49 104 50
rect 102 49 103 50
rect 101 49 102 50
rect 100 49 101 50
rect 99 49 100 50
rect 98 49 99 50
rect 97 49 98 50
rect 96 49 97 50
rect 95 49 96 50
rect 94 49 95 50
rect 93 49 94 50
rect 92 49 93 50
rect 91 49 92 50
rect 90 49 91 50
rect 89 49 90 50
rect 88 49 89 50
rect 87 49 88 50
rect 86 49 87 50
rect 85 49 86 50
rect 84 49 85 50
rect 83 49 84 50
rect 82 49 83 50
rect 81 49 82 50
rect 80 49 81 50
rect 79 49 80 50
rect 78 49 79 50
rect 77 49 78 50
rect 76 49 77 50
rect 75 49 76 50
rect 74 49 75 50
rect 73 49 74 50
rect 72 49 73 50
rect 64 49 65 50
rect 63 49 64 50
rect 62 49 63 50
rect 61 49 62 50
rect 60 49 61 50
rect 59 49 60 50
rect 58 49 59 50
rect 57 49 58 50
rect 56 49 57 50
rect 55 49 56 50
rect 54 49 55 50
rect 53 49 54 50
rect 52 49 53 50
rect 51 49 52 50
rect 50 49 51 50
rect 49 49 50 50
rect 48 49 49 50
rect 47 49 48 50
rect 46 49 47 50
rect 45 49 46 50
rect 44 49 45 50
rect 43 49 44 50
rect 42 49 43 50
rect 41 49 42 50
rect 40 49 41 50
rect 39 49 40 50
rect 38 49 39 50
rect 37 49 38 50
rect 36 49 37 50
rect 35 49 36 50
rect 34 49 35 50
rect 33 49 34 50
rect 28 49 29 50
rect 27 49 28 50
rect 26 49 27 50
rect 25 49 26 50
rect 24 49 25 50
rect 23 49 24 50
rect 22 49 23 50
rect 21 49 22 50
rect 20 49 21 50
rect 19 49 20 50
rect 18 49 19 50
rect 17 49 18 50
rect 16 49 17 50
rect 195 50 196 51
rect 194 50 195 51
rect 189 50 190 51
rect 188 50 189 51
rect 187 50 188 51
rect 178 50 179 51
rect 177 50 178 51
rect 176 50 177 51
rect 175 50 176 51
rect 174 50 175 51
rect 173 50 174 51
rect 172 50 173 51
rect 171 50 172 51
rect 170 50 171 51
rect 169 50 170 51
rect 168 50 169 51
rect 167 50 168 51
rect 166 50 167 51
rect 165 50 166 51
rect 164 50 165 51
rect 163 50 164 51
rect 162 50 163 51
rect 161 50 162 51
rect 102 50 103 51
rect 101 50 102 51
rect 100 50 101 51
rect 99 50 100 51
rect 98 50 99 51
rect 97 50 98 51
rect 96 50 97 51
rect 95 50 96 51
rect 94 50 95 51
rect 93 50 94 51
rect 92 50 93 51
rect 91 50 92 51
rect 90 50 91 51
rect 89 50 90 51
rect 88 50 89 51
rect 87 50 88 51
rect 86 50 87 51
rect 85 50 86 51
rect 84 50 85 51
rect 83 50 84 51
rect 82 50 83 51
rect 81 50 82 51
rect 80 50 81 51
rect 79 50 80 51
rect 78 50 79 51
rect 77 50 78 51
rect 76 50 77 51
rect 75 50 76 51
rect 74 50 75 51
rect 73 50 74 51
rect 72 50 73 51
rect 71 50 72 51
rect 64 50 65 51
rect 63 50 64 51
rect 62 50 63 51
rect 61 50 62 51
rect 60 50 61 51
rect 59 50 60 51
rect 58 50 59 51
rect 57 50 58 51
rect 56 50 57 51
rect 55 50 56 51
rect 54 50 55 51
rect 53 50 54 51
rect 52 50 53 51
rect 51 50 52 51
rect 50 50 51 51
rect 49 50 50 51
rect 48 50 49 51
rect 47 50 48 51
rect 46 50 47 51
rect 45 50 46 51
rect 44 50 45 51
rect 43 50 44 51
rect 42 50 43 51
rect 41 50 42 51
rect 40 50 41 51
rect 39 50 40 51
rect 38 50 39 51
rect 37 50 38 51
rect 36 50 37 51
rect 35 50 36 51
rect 34 50 35 51
rect 33 50 34 51
rect 32 50 33 51
rect 28 50 29 51
rect 27 50 28 51
rect 26 50 27 51
rect 25 50 26 51
rect 24 50 25 51
rect 23 50 24 51
rect 22 50 23 51
rect 21 50 22 51
rect 20 50 21 51
rect 19 50 20 51
rect 18 50 19 51
rect 17 50 18 51
rect 16 50 17 51
rect 190 51 191 52
rect 189 51 190 52
rect 188 51 189 52
rect 187 51 188 52
rect 178 51 179 52
rect 177 51 178 52
rect 176 51 177 52
rect 175 51 176 52
rect 162 51 163 52
rect 161 51 162 52
rect 100 51 101 52
rect 99 51 100 52
rect 98 51 99 52
rect 97 51 98 52
rect 96 51 97 52
rect 95 51 96 52
rect 94 51 95 52
rect 93 51 94 52
rect 92 51 93 52
rect 91 51 92 52
rect 90 51 91 52
rect 89 51 90 52
rect 88 51 89 52
rect 87 51 88 52
rect 86 51 87 52
rect 85 51 86 52
rect 84 51 85 52
rect 83 51 84 52
rect 82 51 83 52
rect 81 51 82 52
rect 80 51 81 52
rect 79 51 80 52
rect 78 51 79 52
rect 77 51 78 52
rect 76 51 77 52
rect 75 51 76 52
rect 74 51 75 52
rect 73 51 74 52
rect 72 51 73 52
rect 71 51 72 52
rect 64 51 65 52
rect 63 51 64 52
rect 62 51 63 52
rect 61 51 62 52
rect 60 51 61 52
rect 59 51 60 52
rect 58 51 59 52
rect 57 51 58 52
rect 56 51 57 52
rect 55 51 56 52
rect 54 51 55 52
rect 53 51 54 52
rect 52 51 53 52
rect 51 51 52 52
rect 50 51 51 52
rect 49 51 50 52
rect 48 51 49 52
rect 47 51 48 52
rect 46 51 47 52
rect 45 51 46 52
rect 44 51 45 52
rect 43 51 44 52
rect 42 51 43 52
rect 41 51 42 52
rect 40 51 41 52
rect 39 51 40 52
rect 38 51 39 52
rect 37 51 38 52
rect 36 51 37 52
rect 35 51 36 52
rect 34 51 35 52
rect 33 51 34 52
rect 32 51 33 52
rect 31 51 32 52
rect 27 51 28 52
rect 26 51 27 52
rect 25 51 26 52
rect 24 51 25 52
rect 23 51 24 52
rect 22 51 23 52
rect 21 51 22 52
rect 20 51 21 52
rect 19 51 20 52
rect 18 51 19 52
rect 17 51 18 52
rect 16 51 17 52
rect 15 51 16 52
rect 191 52 192 53
rect 190 52 191 53
rect 189 52 190 53
rect 179 52 180 53
rect 178 52 179 53
rect 177 52 178 53
rect 176 52 177 53
rect 161 52 162 53
rect 98 52 99 53
rect 97 52 98 53
rect 96 52 97 53
rect 95 52 96 53
rect 94 52 95 53
rect 93 52 94 53
rect 92 52 93 53
rect 91 52 92 53
rect 90 52 91 53
rect 89 52 90 53
rect 88 52 89 53
rect 87 52 88 53
rect 86 52 87 53
rect 85 52 86 53
rect 84 52 85 53
rect 83 52 84 53
rect 82 52 83 53
rect 81 52 82 53
rect 80 52 81 53
rect 79 52 80 53
rect 78 52 79 53
rect 77 52 78 53
rect 76 52 77 53
rect 75 52 76 53
rect 74 52 75 53
rect 73 52 74 53
rect 72 52 73 53
rect 71 52 72 53
rect 70 52 71 53
rect 63 52 64 53
rect 62 52 63 53
rect 61 52 62 53
rect 60 52 61 53
rect 59 52 60 53
rect 58 52 59 53
rect 57 52 58 53
rect 56 52 57 53
rect 55 52 56 53
rect 54 52 55 53
rect 53 52 54 53
rect 52 52 53 53
rect 51 52 52 53
rect 50 52 51 53
rect 49 52 50 53
rect 48 52 49 53
rect 47 52 48 53
rect 46 52 47 53
rect 45 52 46 53
rect 44 52 45 53
rect 43 52 44 53
rect 42 52 43 53
rect 41 52 42 53
rect 40 52 41 53
rect 39 52 40 53
rect 38 52 39 53
rect 37 52 38 53
rect 36 52 37 53
rect 35 52 36 53
rect 34 52 35 53
rect 33 52 34 53
rect 32 52 33 53
rect 31 52 32 53
rect 30 52 31 53
rect 27 52 28 53
rect 26 52 27 53
rect 25 52 26 53
rect 24 52 25 53
rect 23 52 24 53
rect 22 52 23 53
rect 21 52 22 53
rect 20 52 21 53
rect 19 52 20 53
rect 18 52 19 53
rect 17 52 18 53
rect 16 52 17 53
rect 15 52 16 53
rect 192 53 193 54
rect 191 53 192 54
rect 190 53 191 54
rect 179 53 180 54
rect 178 53 179 54
rect 177 53 178 54
rect 120 53 121 54
rect 119 53 120 54
rect 118 53 119 54
rect 117 53 118 54
rect 116 53 117 54
rect 115 53 116 54
rect 114 53 115 54
rect 113 53 114 54
rect 96 53 97 54
rect 95 53 96 54
rect 94 53 95 54
rect 93 53 94 54
rect 92 53 93 54
rect 91 53 92 54
rect 90 53 91 54
rect 89 53 90 54
rect 88 53 89 54
rect 87 53 88 54
rect 86 53 87 54
rect 85 53 86 54
rect 84 53 85 54
rect 83 53 84 54
rect 82 53 83 54
rect 81 53 82 54
rect 80 53 81 54
rect 79 53 80 54
rect 78 53 79 54
rect 77 53 78 54
rect 76 53 77 54
rect 75 53 76 54
rect 74 53 75 54
rect 73 53 74 54
rect 72 53 73 54
rect 71 53 72 54
rect 70 53 71 54
rect 63 53 64 54
rect 62 53 63 54
rect 61 53 62 54
rect 60 53 61 54
rect 59 53 60 54
rect 58 53 59 54
rect 57 53 58 54
rect 56 53 57 54
rect 55 53 56 54
rect 54 53 55 54
rect 53 53 54 54
rect 52 53 53 54
rect 51 53 52 54
rect 50 53 51 54
rect 49 53 50 54
rect 48 53 49 54
rect 47 53 48 54
rect 46 53 47 54
rect 45 53 46 54
rect 44 53 45 54
rect 43 53 44 54
rect 42 53 43 54
rect 41 53 42 54
rect 40 53 41 54
rect 39 53 40 54
rect 38 53 39 54
rect 37 53 38 54
rect 36 53 37 54
rect 35 53 36 54
rect 34 53 35 54
rect 33 53 34 54
rect 32 53 33 54
rect 31 53 32 54
rect 30 53 31 54
rect 27 53 28 54
rect 26 53 27 54
rect 25 53 26 54
rect 24 53 25 54
rect 23 53 24 54
rect 22 53 23 54
rect 21 53 22 54
rect 20 53 21 54
rect 19 53 20 54
rect 18 53 19 54
rect 17 53 18 54
rect 16 53 17 54
rect 15 53 16 54
rect 193 54 194 55
rect 192 54 193 55
rect 191 54 192 55
rect 179 54 180 55
rect 178 54 179 55
rect 177 54 178 55
rect 122 54 123 55
rect 121 54 122 55
rect 120 54 121 55
rect 119 54 120 55
rect 118 54 119 55
rect 117 54 118 55
rect 116 54 117 55
rect 115 54 116 55
rect 114 54 115 55
rect 113 54 114 55
rect 112 54 113 55
rect 111 54 112 55
rect 110 54 111 55
rect 95 54 96 55
rect 94 54 95 55
rect 93 54 94 55
rect 92 54 93 55
rect 91 54 92 55
rect 90 54 91 55
rect 89 54 90 55
rect 88 54 89 55
rect 87 54 88 55
rect 86 54 87 55
rect 85 54 86 55
rect 84 54 85 55
rect 83 54 84 55
rect 82 54 83 55
rect 81 54 82 55
rect 80 54 81 55
rect 79 54 80 55
rect 78 54 79 55
rect 77 54 78 55
rect 76 54 77 55
rect 75 54 76 55
rect 74 54 75 55
rect 73 54 74 55
rect 72 54 73 55
rect 71 54 72 55
rect 70 54 71 55
rect 62 54 63 55
rect 61 54 62 55
rect 60 54 61 55
rect 59 54 60 55
rect 58 54 59 55
rect 57 54 58 55
rect 56 54 57 55
rect 55 54 56 55
rect 54 54 55 55
rect 53 54 54 55
rect 52 54 53 55
rect 51 54 52 55
rect 50 54 51 55
rect 49 54 50 55
rect 48 54 49 55
rect 47 54 48 55
rect 46 54 47 55
rect 45 54 46 55
rect 44 54 45 55
rect 43 54 44 55
rect 42 54 43 55
rect 41 54 42 55
rect 40 54 41 55
rect 39 54 40 55
rect 38 54 39 55
rect 37 54 38 55
rect 36 54 37 55
rect 35 54 36 55
rect 34 54 35 55
rect 33 54 34 55
rect 32 54 33 55
rect 31 54 32 55
rect 30 54 31 55
rect 29 54 30 55
rect 27 54 28 55
rect 26 54 27 55
rect 25 54 26 55
rect 24 54 25 55
rect 23 54 24 55
rect 22 54 23 55
rect 21 54 22 55
rect 20 54 21 55
rect 19 54 20 55
rect 18 54 19 55
rect 17 54 18 55
rect 16 54 17 55
rect 15 54 16 55
rect 195 55 196 56
rect 194 55 195 56
rect 193 55 194 56
rect 192 55 193 56
rect 191 55 192 56
rect 189 55 190 56
rect 188 55 189 56
rect 187 55 188 56
rect 179 55 180 56
rect 178 55 179 56
rect 177 55 178 56
rect 123 55 124 56
rect 122 55 123 56
rect 121 55 122 56
rect 120 55 121 56
rect 119 55 120 56
rect 118 55 119 56
rect 117 55 118 56
rect 116 55 117 56
rect 115 55 116 56
rect 114 55 115 56
rect 113 55 114 56
rect 112 55 113 56
rect 111 55 112 56
rect 110 55 111 56
rect 109 55 110 56
rect 108 55 109 56
rect 95 55 96 56
rect 94 55 95 56
rect 93 55 94 56
rect 92 55 93 56
rect 91 55 92 56
rect 90 55 91 56
rect 89 55 90 56
rect 88 55 89 56
rect 87 55 88 56
rect 86 55 87 56
rect 85 55 86 56
rect 84 55 85 56
rect 83 55 84 56
rect 82 55 83 56
rect 81 55 82 56
rect 80 55 81 56
rect 79 55 80 56
rect 78 55 79 56
rect 77 55 78 56
rect 76 55 77 56
rect 75 55 76 56
rect 74 55 75 56
rect 73 55 74 56
rect 72 55 73 56
rect 71 55 72 56
rect 70 55 71 56
rect 69 55 70 56
rect 62 55 63 56
rect 61 55 62 56
rect 60 55 61 56
rect 59 55 60 56
rect 58 55 59 56
rect 57 55 58 56
rect 56 55 57 56
rect 55 55 56 56
rect 54 55 55 56
rect 53 55 54 56
rect 52 55 53 56
rect 51 55 52 56
rect 50 55 51 56
rect 49 55 50 56
rect 48 55 49 56
rect 47 55 48 56
rect 46 55 47 56
rect 45 55 46 56
rect 44 55 45 56
rect 43 55 44 56
rect 42 55 43 56
rect 41 55 42 56
rect 40 55 41 56
rect 39 55 40 56
rect 38 55 39 56
rect 37 55 38 56
rect 36 55 37 56
rect 35 55 36 56
rect 34 55 35 56
rect 33 55 34 56
rect 32 55 33 56
rect 31 55 32 56
rect 30 55 31 56
rect 29 55 30 56
rect 26 55 27 56
rect 25 55 26 56
rect 24 55 25 56
rect 23 55 24 56
rect 22 55 23 56
rect 21 55 22 56
rect 20 55 21 56
rect 19 55 20 56
rect 18 55 19 56
rect 17 55 18 56
rect 16 55 17 56
rect 15 55 16 56
rect 195 56 196 57
rect 194 56 195 57
rect 193 56 194 57
rect 192 56 193 57
rect 191 56 192 57
rect 190 56 191 57
rect 189 56 190 57
rect 188 56 189 57
rect 187 56 188 57
rect 179 56 180 57
rect 178 56 179 57
rect 177 56 178 57
rect 161 56 162 57
rect 125 56 126 57
rect 124 56 125 57
rect 123 56 124 57
rect 122 56 123 57
rect 121 56 122 57
rect 120 56 121 57
rect 119 56 120 57
rect 118 56 119 57
rect 117 56 118 57
rect 116 56 117 57
rect 115 56 116 57
rect 114 56 115 57
rect 113 56 114 57
rect 112 56 113 57
rect 111 56 112 57
rect 110 56 111 57
rect 109 56 110 57
rect 108 56 109 57
rect 107 56 108 57
rect 106 56 107 57
rect 94 56 95 57
rect 93 56 94 57
rect 92 56 93 57
rect 91 56 92 57
rect 90 56 91 57
rect 89 56 90 57
rect 88 56 89 57
rect 87 56 88 57
rect 86 56 87 57
rect 85 56 86 57
rect 84 56 85 57
rect 83 56 84 57
rect 82 56 83 57
rect 81 56 82 57
rect 80 56 81 57
rect 79 56 80 57
rect 78 56 79 57
rect 77 56 78 57
rect 76 56 77 57
rect 75 56 76 57
rect 74 56 75 57
rect 73 56 74 57
rect 72 56 73 57
rect 71 56 72 57
rect 70 56 71 57
rect 69 56 70 57
rect 61 56 62 57
rect 60 56 61 57
rect 59 56 60 57
rect 58 56 59 57
rect 57 56 58 57
rect 56 56 57 57
rect 55 56 56 57
rect 54 56 55 57
rect 53 56 54 57
rect 52 56 53 57
rect 51 56 52 57
rect 50 56 51 57
rect 49 56 50 57
rect 48 56 49 57
rect 47 56 48 57
rect 46 56 47 57
rect 45 56 46 57
rect 44 56 45 57
rect 43 56 44 57
rect 42 56 43 57
rect 41 56 42 57
rect 40 56 41 57
rect 39 56 40 57
rect 38 56 39 57
rect 37 56 38 57
rect 36 56 37 57
rect 35 56 36 57
rect 34 56 35 57
rect 33 56 34 57
rect 32 56 33 57
rect 31 56 32 57
rect 30 56 31 57
rect 29 56 30 57
rect 28 56 29 57
rect 26 56 27 57
rect 25 56 26 57
rect 24 56 25 57
rect 23 56 24 57
rect 22 56 23 57
rect 21 56 22 57
rect 20 56 21 57
rect 19 56 20 57
rect 18 56 19 57
rect 17 56 18 57
rect 16 56 17 57
rect 178 57 179 58
rect 177 57 178 58
rect 176 57 177 58
rect 161 57 162 58
rect 126 57 127 58
rect 125 57 126 58
rect 124 57 125 58
rect 123 57 124 58
rect 122 57 123 58
rect 121 57 122 58
rect 120 57 121 58
rect 119 57 120 58
rect 118 57 119 58
rect 117 57 118 58
rect 116 57 117 58
rect 115 57 116 58
rect 114 57 115 58
rect 113 57 114 58
rect 112 57 113 58
rect 111 57 112 58
rect 110 57 111 58
rect 109 57 110 58
rect 108 57 109 58
rect 107 57 108 58
rect 106 57 107 58
rect 105 57 106 58
rect 93 57 94 58
rect 92 57 93 58
rect 91 57 92 58
rect 90 57 91 58
rect 89 57 90 58
rect 88 57 89 58
rect 87 57 88 58
rect 86 57 87 58
rect 85 57 86 58
rect 84 57 85 58
rect 83 57 84 58
rect 82 57 83 58
rect 81 57 82 58
rect 80 57 81 58
rect 79 57 80 58
rect 78 57 79 58
rect 77 57 78 58
rect 76 57 77 58
rect 75 57 76 58
rect 74 57 75 58
rect 73 57 74 58
rect 72 57 73 58
rect 71 57 72 58
rect 70 57 71 58
rect 69 57 70 58
rect 68 57 69 58
rect 61 57 62 58
rect 60 57 61 58
rect 59 57 60 58
rect 58 57 59 58
rect 57 57 58 58
rect 56 57 57 58
rect 55 57 56 58
rect 54 57 55 58
rect 53 57 54 58
rect 52 57 53 58
rect 51 57 52 58
rect 50 57 51 58
rect 49 57 50 58
rect 48 57 49 58
rect 47 57 48 58
rect 46 57 47 58
rect 45 57 46 58
rect 44 57 45 58
rect 43 57 44 58
rect 42 57 43 58
rect 41 57 42 58
rect 40 57 41 58
rect 39 57 40 58
rect 38 57 39 58
rect 37 57 38 58
rect 36 57 37 58
rect 35 57 36 58
rect 34 57 35 58
rect 33 57 34 58
rect 32 57 33 58
rect 31 57 32 58
rect 30 57 31 58
rect 29 57 30 58
rect 28 57 29 58
rect 27 57 28 58
rect 26 57 27 58
rect 25 57 26 58
rect 24 57 25 58
rect 23 57 24 58
rect 22 57 23 58
rect 21 57 22 58
rect 20 57 21 58
rect 19 57 20 58
rect 18 57 19 58
rect 17 57 18 58
rect 16 57 17 58
rect 178 58 179 59
rect 177 58 178 59
rect 176 58 177 59
rect 175 58 176 59
rect 162 58 163 59
rect 161 58 162 59
rect 127 58 128 59
rect 126 58 127 59
rect 125 58 126 59
rect 124 58 125 59
rect 123 58 124 59
rect 122 58 123 59
rect 121 58 122 59
rect 120 58 121 59
rect 119 58 120 59
rect 118 58 119 59
rect 117 58 118 59
rect 116 58 117 59
rect 115 58 116 59
rect 114 58 115 59
rect 113 58 114 59
rect 112 58 113 59
rect 111 58 112 59
rect 110 58 111 59
rect 109 58 110 59
rect 108 58 109 59
rect 107 58 108 59
rect 106 58 107 59
rect 105 58 106 59
rect 104 58 105 59
rect 103 58 104 59
rect 93 58 94 59
rect 92 58 93 59
rect 91 58 92 59
rect 90 58 91 59
rect 89 58 90 59
rect 88 58 89 59
rect 87 58 88 59
rect 86 58 87 59
rect 85 58 86 59
rect 84 58 85 59
rect 83 58 84 59
rect 82 58 83 59
rect 81 58 82 59
rect 80 58 81 59
rect 79 58 80 59
rect 78 58 79 59
rect 77 58 78 59
rect 76 58 77 59
rect 75 58 76 59
rect 74 58 75 59
rect 73 58 74 59
rect 72 58 73 59
rect 71 58 72 59
rect 70 58 71 59
rect 69 58 70 59
rect 68 58 69 59
rect 60 58 61 59
rect 59 58 60 59
rect 58 58 59 59
rect 57 58 58 59
rect 56 58 57 59
rect 55 58 56 59
rect 54 58 55 59
rect 53 58 54 59
rect 52 58 53 59
rect 51 58 52 59
rect 50 58 51 59
rect 49 58 50 59
rect 48 58 49 59
rect 47 58 48 59
rect 46 58 47 59
rect 45 58 46 59
rect 44 58 45 59
rect 43 58 44 59
rect 42 58 43 59
rect 41 58 42 59
rect 40 58 41 59
rect 39 58 40 59
rect 38 58 39 59
rect 37 58 38 59
rect 36 58 37 59
rect 35 58 36 59
rect 34 58 35 59
rect 33 58 34 59
rect 32 58 33 59
rect 31 58 32 59
rect 30 58 31 59
rect 29 58 30 59
rect 28 58 29 59
rect 27 58 28 59
rect 26 58 27 59
rect 25 58 26 59
rect 24 58 25 59
rect 23 58 24 59
rect 22 58 23 59
rect 21 58 22 59
rect 20 58 21 59
rect 19 58 20 59
rect 18 58 19 59
rect 17 58 18 59
rect 177 59 178 60
rect 176 59 177 60
rect 175 59 176 60
rect 174 59 175 60
rect 173 59 174 60
rect 172 59 173 60
rect 171 59 172 60
rect 170 59 171 60
rect 169 59 170 60
rect 168 59 169 60
rect 167 59 168 60
rect 166 59 167 60
rect 165 59 166 60
rect 164 59 165 60
rect 163 59 164 60
rect 162 59 163 60
rect 161 59 162 60
rect 128 59 129 60
rect 127 59 128 60
rect 126 59 127 60
rect 125 59 126 60
rect 124 59 125 60
rect 123 59 124 60
rect 122 59 123 60
rect 121 59 122 60
rect 120 59 121 60
rect 119 59 120 60
rect 118 59 119 60
rect 117 59 118 60
rect 116 59 117 60
rect 115 59 116 60
rect 114 59 115 60
rect 113 59 114 60
rect 112 59 113 60
rect 111 59 112 60
rect 110 59 111 60
rect 109 59 110 60
rect 108 59 109 60
rect 107 59 108 60
rect 106 59 107 60
rect 105 59 106 60
rect 104 59 105 60
rect 103 59 104 60
rect 102 59 103 60
rect 92 59 93 60
rect 91 59 92 60
rect 90 59 91 60
rect 89 59 90 60
rect 88 59 89 60
rect 87 59 88 60
rect 86 59 87 60
rect 85 59 86 60
rect 84 59 85 60
rect 83 59 84 60
rect 82 59 83 60
rect 81 59 82 60
rect 80 59 81 60
rect 79 59 80 60
rect 78 59 79 60
rect 77 59 78 60
rect 76 59 77 60
rect 75 59 76 60
rect 74 59 75 60
rect 73 59 74 60
rect 72 59 73 60
rect 71 59 72 60
rect 70 59 71 60
rect 69 59 70 60
rect 68 59 69 60
rect 67 59 68 60
rect 59 59 60 60
rect 58 59 59 60
rect 57 59 58 60
rect 56 59 57 60
rect 55 59 56 60
rect 54 59 55 60
rect 53 59 54 60
rect 52 59 53 60
rect 51 59 52 60
rect 50 59 51 60
rect 49 59 50 60
rect 48 59 49 60
rect 47 59 48 60
rect 46 59 47 60
rect 45 59 46 60
rect 44 59 45 60
rect 43 59 44 60
rect 42 59 43 60
rect 41 59 42 60
rect 40 59 41 60
rect 39 59 40 60
rect 38 59 39 60
rect 37 59 38 60
rect 36 59 37 60
rect 35 59 36 60
rect 34 59 35 60
rect 33 59 34 60
rect 32 59 33 60
rect 31 59 32 60
rect 30 59 31 60
rect 29 59 30 60
rect 28 59 29 60
rect 27 59 28 60
rect 26 59 27 60
rect 25 59 26 60
rect 24 59 25 60
rect 23 59 24 60
rect 22 59 23 60
rect 21 59 22 60
rect 20 59 21 60
rect 19 59 20 60
rect 18 59 19 60
rect 176 60 177 61
rect 175 60 176 61
rect 174 60 175 61
rect 173 60 174 61
rect 172 60 173 61
rect 171 60 172 61
rect 170 60 171 61
rect 169 60 170 61
rect 168 60 169 61
rect 167 60 168 61
rect 166 60 167 61
rect 165 60 166 61
rect 164 60 165 61
rect 163 60 164 61
rect 162 60 163 61
rect 161 60 162 61
rect 128 60 129 61
rect 127 60 128 61
rect 126 60 127 61
rect 125 60 126 61
rect 124 60 125 61
rect 123 60 124 61
rect 122 60 123 61
rect 121 60 122 61
rect 120 60 121 61
rect 119 60 120 61
rect 118 60 119 61
rect 117 60 118 61
rect 116 60 117 61
rect 115 60 116 61
rect 114 60 115 61
rect 113 60 114 61
rect 112 60 113 61
rect 111 60 112 61
rect 110 60 111 61
rect 109 60 110 61
rect 108 60 109 61
rect 107 60 108 61
rect 106 60 107 61
rect 105 60 106 61
rect 104 60 105 61
rect 103 60 104 61
rect 102 60 103 61
rect 101 60 102 61
rect 92 60 93 61
rect 91 60 92 61
rect 90 60 91 61
rect 89 60 90 61
rect 88 60 89 61
rect 87 60 88 61
rect 86 60 87 61
rect 85 60 86 61
rect 84 60 85 61
rect 83 60 84 61
rect 82 60 83 61
rect 81 60 82 61
rect 80 60 81 61
rect 79 60 80 61
rect 78 60 79 61
rect 77 60 78 61
rect 76 60 77 61
rect 75 60 76 61
rect 74 60 75 61
rect 73 60 74 61
rect 72 60 73 61
rect 71 60 72 61
rect 70 60 71 61
rect 69 60 70 61
rect 68 60 69 61
rect 67 60 68 61
rect 58 60 59 61
rect 57 60 58 61
rect 56 60 57 61
rect 55 60 56 61
rect 54 60 55 61
rect 53 60 54 61
rect 52 60 53 61
rect 51 60 52 61
rect 50 60 51 61
rect 49 60 50 61
rect 48 60 49 61
rect 47 60 48 61
rect 46 60 47 61
rect 45 60 46 61
rect 44 60 45 61
rect 43 60 44 61
rect 42 60 43 61
rect 41 60 42 61
rect 40 60 41 61
rect 39 60 40 61
rect 38 60 39 61
rect 37 60 38 61
rect 36 60 37 61
rect 35 60 36 61
rect 34 60 35 61
rect 33 60 34 61
rect 32 60 33 61
rect 31 60 32 61
rect 30 60 31 61
rect 29 60 30 61
rect 28 60 29 61
rect 27 60 28 61
rect 26 60 27 61
rect 25 60 26 61
rect 24 60 25 61
rect 23 60 24 61
rect 22 60 23 61
rect 21 60 22 61
rect 20 60 21 61
rect 19 60 20 61
rect 12 60 13 61
rect 195 61 196 62
rect 194 61 195 62
rect 187 61 188 62
rect 173 61 174 62
rect 165 61 166 62
rect 164 61 165 62
rect 163 61 164 62
rect 162 61 163 62
rect 161 61 162 62
rect 129 61 130 62
rect 128 61 129 62
rect 127 61 128 62
rect 126 61 127 62
rect 125 61 126 62
rect 124 61 125 62
rect 123 61 124 62
rect 122 61 123 62
rect 121 61 122 62
rect 120 61 121 62
rect 119 61 120 62
rect 118 61 119 62
rect 117 61 118 62
rect 116 61 117 62
rect 115 61 116 62
rect 114 61 115 62
rect 113 61 114 62
rect 112 61 113 62
rect 111 61 112 62
rect 110 61 111 62
rect 109 61 110 62
rect 108 61 109 62
rect 107 61 108 62
rect 106 61 107 62
rect 105 61 106 62
rect 104 61 105 62
rect 103 61 104 62
rect 102 61 103 62
rect 101 61 102 62
rect 100 61 101 62
rect 91 61 92 62
rect 90 61 91 62
rect 89 61 90 62
rect 88 61 89 62
rect 87 61 88 62
rect 86 61 87 62
rect 85 61 86 62
rect 84 61 85 62
rect 83 61 84 62
rect 82 61 83 62
rect 81 61 82 62
rect 80 61 81 62
rect 79 61 80 62
rect 78 61 79 62
rect 77 61 78 62
rect 76 61 77 62
rect 75 61 76 62
rect 74 61 75 62
rect 73 61 74 62
rect 72 61 73 62
rect 71 61 72 62
rect 70 61 71 62
rect 69 61 70 62
rect 68 61 69 62
rect 67 61 68 62
rect 66 61 67 62
rect 57 61 58 62
rect 56 61 57 62
rect 55 61 56 62
rect 54 61 55 62
rect 53 61 54 62
rect 52 61 53 62
rect 51 61 52 62
rect 50 61 51 62
rect 49 61 50 62
rect 48 61 49 62
rect 47 61 48 62
rect 46 61 47 62
rect 45 61 46 62
rect 44 61 45 62
rect 43 61 44 62
rect 42 61 43 62
rect 41 61 42 62
rect 40 61 41 62
rect 39 61 40 62
rect 38 61 39 62
rect 37 61 38 62
rect 36 61 37 62
rect 35 61 36 62
rect 34 61 35 62
rect 33 61 34 62
rect 32 61 33 62
rect 31 61 32 62
rect 30 61 31 62
rect 29 61 30 62
rect 28 61 29 62
rect 27 61 28 62
rect 26 61 27 62
rect 25 61 26 62
rect 24 61 25 62
rect 23 61 24 62
rect 22 61 23 62
rect 21 61 22 62
rect 20 61 21 62
rect 19 61 20 62
rect 14 61 15 62
rect 13 61 14 62
rect 12 61 13 62
rect 11 61 12 62
rect 10 61 11 62
rect 194 62 195 63
rect 193 62 194 63
rect 192 62 193 63
rect 191 62 192 63
rect 190 62 191 63
rect 189 62 190 63
rect 188 62 189 63
rect 187 62 188 63
rect 162 62 163 63
rect 161 62 162 63
rect 130 62 131 63
rect 129 62 130 63
rect 128 62 129 63
rect 127 62 128 63
rect 126 62 127 63
rect 125 62 126 63
rect 124 62 125 63
rect 123 62 124 63
rect 122 62 123 63
rect 121 62 122 63
rect 120 62 121 63
rect 119 62 120 63
rect 118 62 119 63
rect 117 62 118 63
rect 116 62 117 63
rect 115 62 116 63
rect 114 62 115 63
rect 113 62 114 63
rect 112 62 113 63
rect 111 62 112 63
rect 110 62 111 63
rect 109 62 110 63
rect 108 62 109 63
rect 107 62 108 63
rect 106 62 107 63
rect 105 62 106 63
rect 104 62 105 63
rect 103 62 104 63
rect 102 62 103 63
rect 101 62 102 63
rect 100 62 101 63
rect 91 62 92 63
rect 90 62 91 63
rect 89 62 90 63
rect 88 62 89 63
rect 87 62 88 63
rect 86 62 87 63
rect 85 62 86 63
rect 84 62 85 63
rect 83 62 84 63
rect 82 62 83 63
rect 81 62 82 63
rect 80 62 81 63
rect 79 62 80 63
rect 78 62 79 63
rect 77 62 78 63
rect 76 62 77 63
rect 75 62 76 63
rect 74 62 75 63
rect 73 62 74 63
rect 72 62 73 63
rect 71 62 72 63
rect 70 62 71 63
rect 69 62 70 63
rect 68 62 69 63
rect 67 62 68 63
rect 66 62 67 63
rect 56 62 57 63
rect 55 62 56 63
rect 54 62 55 63
rect 53 62 54 63
rect 52 62 53 63
rect 51 62 52 63
rect 50 62 51 63
rect 49 62 50 63
rect 48 62 49 63
rect 47 62 48 63
rect 46 62 47 63
rect 45 62 46 63
rect 44 62 45 63
rect 43 62 44 63
rect 42 62 43 63
rect 41 62 42 63
rect 40 62 41 63
rect 39 62 40 63
rect 38 62 39 63
rect 37 62 38 63
rect 36 62 37 63
rect 35 62 36 63
rect 34 62 35 63
rect 33 62 34 63
rect 32 62 33 63
rect 31 62 32 63
rect 30 62 31 63
rect 29 62 30 63
rect 28 62 29 63
rect 27 62 28 63
rect 26 62 27 63
rect 25 62 26 63
rect 24 62 25 63
rect 23 62 24 63
rect 22 62 23 63
rect 21 62 22 63
rect 20 62 21 63
rect 19 62 20 63
rect 14 62 15 63
rect 13 62 14 63
rect 12 62 13 63
rect 11 62 12 63
rect 10 62 11 63
rect 9 62 10 63
rect 8 62 9 63
rect 194 63 195 64
rect 193 63 194 64
rect 192 63 193 64
rect 191 63 192 64
rect 190 63 191 64
rect 189 63 190 64
rect 188 63 189 64
rect 187 63 188 64
rect 161 63 162 64
rect 130 63 131 64
rect 129 63 130 64
rect 128 63 129 64
rect 127 63 128 64
rect 126 63 127 64
rect 125 63 126 64
rect 124 63 125 64
rect 123 63 124 64
rect 122 63 123 64
rect 121 63 122 64
rect 120 63 121 64
rect 119 63 120 64
rect 118 63 119 64
rect 117 63 118 64
rect 116 63 117 64
rect 115 63 116 64
rect 114 63 115 64
rect 113 63 114 64
rect 112 63 113 64
rect 111 63 112 64
rect 110 63 111 64
rect 109 63 110 64
rect 108 63 109 64
rect 107 63 108 64
rect 106 63 107 64
rect 105 63 106 64
rect 104 63 105 64
rect 103 63 104 64
rect 102 63 103 64
rect 101 63 102 64
rect 100 63 101 64
rect 99 63 100 64
rect 90 63 91 64
rect 89 63 90 64
rect 88 63 89 64
rect 87 63 88 64
rect 86 63 87 64
rect 85 63 86 64
rect 84 63 85 64
rect 83 63 84 64
rect 82 63 83 64
rect 81 63 82 64
rect 80 63 81 64
rect 79 63 80 64
rect 78 63 79 64
rect 77 63 78 64
rect 76 63 77 64
rect 75 63 76 64
rect 74 63 75 64
rect 73 63 74 64
rect 72 63 73 64
rect 71 63 72 64
rect 70 63 71 64
rect 69 63 70 64
rect 68 63 69 64
rect 67 63 68 64
rect 66 63 67 64
rect 65 63 66 64
rect 55 63 56 64
rect 54 63 55 64
rect 53 63 54 64
rect 52 63 53 64
rect 51 63 52 64
rect 50 63 51 64
rect 49 63 50 64
rect 48 63 49 64
rect 47 63 48 64
rect 46 63 47 64
rect 45 63 46 64
rect 44 63 45 64
rect 43 63 44 64
rect 42 63 43 64
rect 41 63 42 64
rect 40 63 41 64
rect 39 63 40 64
rect 38 63 39 64
rect 37 63 38 64
rect 36 63 37 64
rect 35 63 36 64
rect 34 63 35 64
rect 33 63 34 64
rect 32 63 33 64
rect 31 63 32 64
rect 30 63 31 64
rect 29 63 30 64
rect 28 63 29 64
rect 27 63 28 64
rect 26 63 27 64
rect 25 63 26 64
rect 24 63 25 64
rect 23 63 24 64
rect 22 63 23 64
rect 21 63 22 64
rect 20 63 21 64
rect 19 63 20 64
rect 15 63 16 64
rect 14 63 15 64
rect 13 63 14 64
rect 12 63 13 64
rect 11 63 12 64
rect 10 63 11 64
rect 9 63 10 64
rect 8 63 9 64
rect 131 64 132 65
rect 130 64 131 65
rect 129 64 130 65
rect 128 64 129 65
rect 127 64 128 65
rect 126 64 127 65
rect 125 64 126 65
rect 124 64 125 65
rect 123 64 124 65
rect 122 64 123 65
rect 121 64 122 65
rect 120 64 121 65
rect 119 64 120 65
rect 118 64 119 65
rect 117 64 118 65
rect 116 64 117 65
rect 115 64 116 65
rect 114 64 115 65
rect 113 64 114 65
rect 112 64 113 65
rect 111 64 112 65
rect 110 64 111 65
rect 109 64 110 65
rect 108 64 109 65
rect 107 64 108 65
rect 106 64 107 65
rect 105 64 106 65
rect 104 64 105 65
rect 103 64 104 65
rect 102 64 103 65
rect 101 64 102 65
rect 100 64 101 65
rect 99 64 100 65
rect 98 64 99 65
rect 90 64 91 65
rect 89 64 90 65
rect 88 64 89 65
rect 87 64 88 65
rect 86 64 87 65
rect 85 64 86 65
rect 84 64 85 65
rect 83 64 84 65
rect 82 64 83 65
rect 81 64 82 65
rect 80 64 81 65
rect 79 64 80 65
rect 78 64 79 65
rect 77 64 78 65
rect 76 64 77 65
rect 75 64 76 65
rect 74 64 75 65
rect 73 64 74 65
rect 72 64 73 65
rect 71 64 72 65
rect 70 64 71 65
rect 69 64 70 65
rect 68 64 69 65
rect 67 64 68 65
rect 66 64 67 65
rect 65 64 66 65
rect 64 64 65 65
rect 53 64 54 65
rect 52 64 53 65
rect 51 64 52 65
rect 50 64 51 65
rect 49 64 50 65
rect 48 64 49 65
rect 47 64 48 65
rect 46 64 47 65
rect 45 64 46 65
rect 44 64 45 65
rect 43 64 44 65
rect 42 64 43 65
rect 41 64 42 65
rect 40 64 41 65
rect 39 64 40 65
rect 38 64 39 65
rect 37 64 38 65
rect 36 64 37 65
rect 35 64 36 65
rect 34 64 35 65
rect 33 64 34 65
rect 32 64 33 65
rect 31 64 32 65
rect 30 64 31 65
rect 29 64 30 65
rect 28 64 29 65
rect 27 64 28 65
rect 26 64 27 65
rect 25 64 26 65
rect 24 64 25 65
rect 23 64 24 65
rect 22 64 23 65
rect 21 64 22 65
rect 20 64 21 65
rect 19 64 20 65
rect 18 64 19 65
rect 14 64 15 65
rect 13 64 14 65
rect 12 64 13 65
rect 11 64 12 65
rect 10 64 11 65
rect 9 64 10 65
rect 8 64 9 65
rect 7 64 8 65
rect 161 65 162 66
rect 132 65 133 66
rect 131 65 132 66
rect 130 65 131 66
rect 129 65 130 66
rect 128 65 129 66
rect 127 65 128 66
rect 126 65 127 66
rect 125 65 126 66
rect 124 65 125 66
rect 123 65 124 66
rect 122 65 123 66
rect 121 65 122 66
rect 120 65 121 66
rect 119 65 120 66
rect 118 65 119 66
rect 117 65 118 66
rect 116 65 117 66
rect 115 65 116 66
rect 114 65 115 66
rect 113 65 114 66
rect 112 65 113 66
rect 111 65 112 66
rect 110 65 111 66
rect 109 65 110 66
rect 108 65 109 66
rect 107 65 108 66
rect 106 65 107 66
rect 105 65 106 66
rect 104 65 105 66
rect 103 65 104 66
rect 102 65 103 66
rect 101 65 102 66
rect 100 65 101 66
rect 99 65 100 66
rect 98 65 99 66
rect 90 65 91 66
rect 89 65 90 66
rect 88 65 89 66
rect 87 65 88 66
rect 86 65 87 66
rect 85 65 86 66
rect 84 65 85 66
rect 83 65 84 66
rect 82 65 83 66
rect 81 65 82 66
rect 80 65 81 66
rect 79 65 80 66
rect 78 65 79 66
rect 77 65 78 66
rect 76 65 77 66
rect 75 65 76 66
rect 74 65 75 66
rect 73 65 74 66
rect 72 65 73 66
rect 71 65 72 66
rect 70 65 71 66
rect 69 65 70 66
rect 68 65 69 66
rect 67 65 68 66
rect 66 65 67 66
rect 65 65 66 66
rect 64 65 65 66
rect 63 65 64 66
rect 52 65 53 66
rect 51 65 52 66
rect 50 65 51 66
rect 49 65 50 66
rect 48 65 49 66
rect 47 65 48 66
rect 46 65 47 66
rect 45 65 46 66
rect 44 65 45 66
rect 43 65 44 66
rect 42 65 43 66
rect 41 65 42 66
rect 40 65 41 66
rect 39 65 40 66
rect 38 65 39 66
rect 37 65 38 66
rect 36 65 37 66
rect 35 65 36 66
rect 34 65 35 66
rect 33 65 34 66
rect 32 65 33 66
rect 31 65 32 66
rect 30 65 31 66
rect 29 65 30 66
rect 28 65 29 66
rect 27 65 28 66
rect 26 65 27 66
rect 25 65 26 66
rect 24 65 25 66
rect 23 65 24 66
rect 22 65 23 66
rect 21 65 22 66
rect 20 65 21 66
rect 19 65 20 66
rect 18 65 19 66
rect 14 65 15 66
rect 13 65 14 66
rect 12 65 13 66
rect 11 65 12 66
rect 10 65 11 66
rect 9 65 10 66
rect 8 65 9 66
rect 7 65 8 66
rect 6 65 7 66
rect 178 66 179 67
rect 161 66 162 67
rect 133 66 134 67
rect 132 66 133 67
rect 131 66 132 67
rect 130 66 131 67
rect 129 66 130 67
rect 128 66 129 67
rect 127 66 128 67
rect 126 66 127 67
rect 125 66 126 67
rect 124 66 125 67
rect 123 66 124 67
rect 122 66 123 67
rect 121 66 122 67
rect 120 66 121 67
rect 119 66 120 67
rect 118 66 119 67
rect 117 66 118 67
rect 116 66 117 67
rect 115 66 116 67
rect 114 66 115 67
rect 113 66 114 67
rect 112 66 113 67
rect 111 66 112 67
rect 110 66 111 67
rect 109 66 110 67
rect 108 66 109 67
rect 107 66 108 67
rect 106 66 107 67
rect 105 66 106 67
rect 104 66 105 67
rect 103 66 104 67
rect 102 66 103 67
rect 101 66 102 67
rect 100 66 101 67
rect 99 66 100 67
rect 98 66 99 67
rect 97 66 98 67
rect 89 66 90 67
rect 88 66 89 67
rect 87 66 88 67
rect 86 66 87 67
rect 85 66 86 67
rect 84 66 85 67
rect 83 66 84 67
rect 82 66 83 67
rect 81 66 82 67
rect 80 66 81 67
rect 79 66 80 67
rect 78 66 79 67
rect 77 66 78 67
rect 76 66 77 67
rect 75 66 76 67
rect 74 66 75 67
rect 73 66 74 67
rect 72 66 73 67
rect 71 66 72 67
rect 70 66 71 67
rect 69 66 70 67
rect 68 66 69 67
rect 67 66 68 67
rect 66 66 67 67
rect 65 66 66 67
rect 64 66 65 67
rect 63 66 64 67
rect 62 66 63 67
rect 50 66 51 67
rect 49 66 50 67
rect 48 66 49 67
rect 47 66 48 67
rect 46 66 47 67
rect 45 66 46 67
rect 44 66 45 67
rect 43 66 44 67
rect 42 66 43 67
rect 41 66 42 67
rect 40 66 41 67
rect 39 66 40 67
rect 38 66 39 67
rect 37 66 38 67
rect 36 66 37 67
rect 35 66 36 67
rect 34 66 35 67
rect 33 66 34 67
rect 32 66 33 67
rect 31 66 32 67
rect 30 66 31 67
rect 29 66 30 67
rect 28 66 29 67
rect 27 66 28 67
rect 26 66 27 67
rect 25 66 26 67
rect 24 66 25 67
rect 23 66 24 67
rect 22 66 23 67
rect 21 66 22 67
rect 20 66 21 67
rect 19 66 20 67
rect 18 66 19 67
rect 17 66 18 67
rect 14 66 15 67
rect 13 66 14 67
rect 12 66 13 67
rect 11 66 12 67
rect 10 66 11 67
rect 9 66 10 67
rect 8 66 9 67
rect 7 66 8 67
rect 6 66 7 67
rect 178 67 179 68
rect 177 67 178 68
rect 162 67 163 68
rect 161 67 162 68
rect 134 67 135 68
rect 133 67 134 68
rect 132 67 133 68
rect 131 67 132 68
rect 120 67 121 68
rect 119 67 120 68
rect 118 67 119 68
rect 117 67 118 68
rect 116 67 117 68
rect 115 67 116 68
rect 114 67 115 68
rect 113 67 114 68
rect 112 67 113 68
rect 111 67 112 68
rect 110 67 111 68
rect 109 67 110 68
rect 108 67 109 68
rect 107 67 108 68
rect 106 67 107 68
rect 105 67 106 68
rect 104 67 105 68
rect 103 67 104 68
rect 102 67 103 68
rect 101 67 102 68
rect 100 67 101 68
rect 99 67 100 68
rect 98 67 99 68
rect 97 67 98 68
rect 96 67 97 68
rect 89 67 90 68
rect 88 67 89 68
rect 87 67 88 68
rect 86 67 87 68
rect 85 67 86 68
rect 84 67 85 68
rect 83 67 84 68
rect 82 67 83 68
rect 81 67 82 68
rect 80 67 81 68
rect 79 67 80 68
rect 78 67 79 68
rect 77 67 78 68
rect 76 67 77 68
rect 75 67 76 68
rect 74 67 75 68
rect 73 67 74 68
rect 72 67 73 68
rect 71 67 72 68
rect 70 67 71 68
rect 69 67 70 68
rect 68 67 69 68
rect 67 67 68 68
rect 66 67 67 68
rect 65 67 66 68
rect 64 67 65 68
rect 63 67 64 68
rect 62 67 63 68
rect 49 67 50 68
rect 48 67 49 68
rect 47 67 48 68
rect 46 67 47 68
rect 45 67 46 68
rect 44 67 45 68
rect 43 67 44 68
rect 42 67 43 68
rect 41 67 42 68
rect 40 67 41 68
rect 39 67 40 68
rect 38 67 39 68
rect 37 67 38 68
rect 36 67 37 68
rect 35 67 36 68
rect 34 67 35 68
rect 33 67 34 68
rect 32 67 33 68
rect 31 67 32 68
rect 30 67 31 68
rect 29 67 30 68
rect 28 67 29 68
rect 27 67 28 68
rect 26 67 27 68
rect 25 67 26 68
rect 24 67 25 68
rect 23 67 24 68
rect 22 67 23 68
rect 21 67 22 68
rect 20 67 21 68
rect 19 67 20 68
rect 18 67 19 68
rect 17 67 18 68
rect 13 67 14 68
rect 12 67 13 68
rect 11 67 12 68
rect 10 67 11 68
rect 9 67 10 68
rect 8 67 9 68
rect 7 67 8 68
rect 6 67 7 68
rect 187 68 188 69
rect 178 68 179 69
rect 177 68 178 69
rect 176 68 177 69
rect 175 68 176 69
rect 174 68 175 69
rect 173 68 174 69
rect 172 68 173 69
rect 171 68 172 69
rect 170 68 171 69
rect 169 68 170 69
rect 168 68 169 69
rect 167 68 168 69
rect 166 68 167 69
rect 165 68 166 69
rect 164 68 165 69
rect 163 68 164 69
rect 162 68 163 69
rect 161 68 162 69
rect 117 68 118 69
rect 116 68 117 69
rect 115 68 116 69
rect 114 68 115 69
rect 113 68 114 69
rect 112 68 113 69
rect 111 68 112 69
rect 110 68 111 69
rect 109 68 110 69
rect 108 68 109 69
rect 107 68 108 69
rect 106 68 107 69
rect 105 68 106 69
rect 104 68 105 69
rect 103 68 104 69
rect 102 68 103 69
rect 101 68 102 69
rect 100 68 101 69
rect 99 68 100 69
rect 98 68 99 69
rect 97 68 98 69
rect 96 68 97 69
rect 88 68 89 69
rect 87 68 88 69
rect 86 68 87 69
rect 85 68 86 69
rect 84 68 85 69
rect 83 68 84 69
rect 82 68 83 69
rect 81 68 82 69
rect 80 68 81 69
rect 79 68 80 69
rect 78 68 79 69
rect 77 68 78 69
rect 76 68 77 69
rect 75 68 76 69
rect 74 68 75 69
rect 73 68 74 69
rect 72 68 73 69
rect 71 68 72 69
rect 70 68 71 69
rect 69 68 70 69
rect 68 68 69 69
rect 67 68 68 69
rect 66 68 67 69
rect 65 68 66 69
rect 64 68 65 69
rect 63 68 64 69
rect 62 68 63 69
rect 61 68 62 69
rect 47 68 48 69
rect 46 68 47 69
rect 45 68 46 69
rect 44 68 45 69
rect 43 68 44 69
rect 42 68 43 69
rect 41 68 42 69
rect 40 68 41 69
rect 39 68 40 69
rect 38 68 39 69
rect 37 68 38 69
rect 36 68 37 69
rect 35 68 36 69
rect 34 68 35 69
rect 33 68 34 69
rect 32 68 33 69
rect 31 68 32 69
rect 30 68 31 69
rect 29 68 30 69
rect 28 68 29 69
rect 27 68 28 69
rect 26 68 27 69
rect 25 68 26 69
rect 24 68 25 69
rect 23 68 24 69
rect 22 68 23 69
rect 21 68 22 69
rect 20 68 21 69
rect 19 68 20 69
rect 18 68 19 69
rect 17 68 18 69
rect 13 68 14 69
rect 12 68 13 69
rect 11 68 12 69
rect 10 68 11 69
rect 9 68 10 69
rect 8 68 9 69
rect 7 68 8 69
rect 6 68 7 69
rect 189 69 190 70
rect 188 69 189 70
rect 187 69 188 70
rect 178 69 179 70
rect 177 69 178 70
rect 176 69 177 70
rect 175 69 176 70
rect 174 69 175 70
rect 173 69 174 70
rect 172 69 173 70
rect 171 69 172 70
rect 170 69 171 70
rect 169 69 170 70
rect 168 69 169 70
rect 167 69 168 70
rect 166 69 167 70
rect 165 69 166 70
rect 164 69 165 70
rect 163 69 164 70
rect 162 69 163 70
rect 161 69 162 70
rect 115 69 116 70
rect 114 69 115 70
rect 113 69 114 70
rect 112 69 113 70
rect 111 69 112 70
rect 110 69 111 70
rect 109 69 110 70
rect 108 69 109 70
rect 107 69 108 70
rect 106 69 107 70
rect 105 69 106 70
rect 104 69 105 70
rect 103 69 104 70
rect 102 69 103 70
rect 101 69 102 70
rect 100 69 101 70
rect 99 69 100 70
rect 98 69 99 70
rect 97 69 98 70
rect 96 69 97 70
rect 95 69 96 70
rect 88 69 89 70
rect 87 69 88 70
rect 86 69 87 70
rect 85 69 86 70
rect 84 69 85 70
rect 83 69 84 70
rect 82 69 83 70
rect 81 69 82 70
rect 80 69 81 70
rect 79 69 80 70
rect 78 69 79 70
rect 77 69 78 70
rect 76 69 77 70
rect 75 69 76 70
rect 74 69 75 70
rect 73 69 74 70
rect 72 69 73 70
rect 71 69 72 70
rect 70 69 71 70
rect 69 69 70 70
rect 68 69 69 70
rect 67 69 68 70
rect 66 69 67 70
rect 65 69 66 70
rect 64 69 65 70
rect 63 69 64 70
rect 62 69 63 70
rect 61 69 62 70
rect 60 69 61 70
rect 59 69 60 70
rect 46 69 47 70
rect 45 69 46 70
rect 44 69 45 70
rect 43 69 44 70
rect 42 69 43 70
rect 41 69 42 70
rect 40 69 41 70
rect 39 69 40 70
rect 38 69 39 70
rect 37 69 38 70
rect 36 69 37 70
rect 35 69 36 70
rect 34 69 35 70
rect 33 69 34 70
rect 32 69 33 70
rect 30 69 31 70
rect 29 69 30 70
rect 28 69 29 70
rect 27 69 28 70
rect 26 69 27 70
rect 25 69 26 70
rect 24 69 25 70
rect 23 69 24 70
rect 22 69 23 70
rect 21 69 22 70
rect 20 69 21 70
rect 19 69 20 70
rect 18 69 19 70
rect 17 69 18 70
rect 16 69 17 70
rect 12 69 13 70
rect 11 69 12 70
rect 10 69 11 70
rect 9 69 10 70
rect 8 69 9 70
rect 7 69 8 70
rect 6 69 7 70
rect 191 70 192 71
rect 190 70 191 71
rect 189 70 190 71
rect 188 70 189 71
rect 187 70 188 71
rect 178 70 179 71
rect 177 70 178 71
rect 166 70 167 71
rect 165 70 166 71
rect 164 70 165 71
rect 163 70 164 71
rect 162 70 163 71
rect 161 70 162 71
rect 113 70 114 71
rect 112 70 113 71
rect 111 70 112 71
rect 110 70 111 71
rect 109 70 110 71
rect 108 70 109 71
rect 107 70 108 71
rect 106 70 107 71
rect 105 70 106 71
rect 104 70 105 71
rect 103 70 104 71
rect 102 70 103 71
rect 101 70 102 71
rect 100 70 101 71
rect 99 70 100 71
rect 98 70 99 71
rect 97 70 98 71
rect 96 70 97 71
rect 95 70 96 71
rect 87 70 88 71
rect 86 70 87 71
rect 85 70 86 71
rect 84 70 85 71
rect 83 70 84 71
rect 82 70 83 71
rect 81 70 82 71
rect 80 70 81 71
rect 79 70 80 71
rect 78 70 79 71
rect 77 70 78 71
rect 76 70 77 71
rect 75 70 76 71
rect 74 70 75 71
rect 73 70 74 71
rect 72 70 73 71
rect 71 70 72 71
rect 70 70 71 71
rect 69 70 70 71
rect 68 70 69 71
rect 67 70 68 71
rect 66 70 67 71
rect 65 70 66 71
rect 64 70 65 71
rect 63 70 64 71
rect 62 70 63 71
rect 61 70 62 71
rect 60 70 61 71
rect 59 70 60 71
rect 58 70 59 71
rect 43 70 44 71
rect 42 70 43 71
rect 41 70 42 71
rect 40 70 41 71
rect 39 70 40 71
rect 38 70 39 71
rect 37 70 38 71
rect 36 70 37 71
rect 28 70 29 71
rect 27 70 28 71
rect 26 70 27 71
rect 25 70 26 71
rect 24 70 25 71
rect 23 70 24 71
rect 22 70 23 71
rect 21 70 22 71
rect 20 70 21 71
rect 19 70 20 71
rect 18 70 19 71
rect 17 70 18 71
rect 16 70 17 71
rect 12 70 13 71
rect 11 70 12 71
rect 10 70 11 71
rect 9 70 10 71
rect 8 70 9 71
rect 7 70 8 71
rect 194 71 195 72
rect 193 71 194 72
rect 192 71 193 72
rect 191 71 192 72
rect 190 71 191 72
rect 189 71 190 72
rect 187 71 188 72
rect 178 71 179 72
rect 167 71 168 72
rect 166 71 167 72
rect 165 71 166 72
rect 164 71 165 72
rect 163 71 164 72
rect 162 71 163 72
rect 112 71 113 72
rect 111 71 112 72
rect 110 71 111 72
rect 109 71 110 72
rect 108 71 109 72
rect 107 71 108 72
rect 106 71 107 72
rect 105 71 106 72
rect 104 71 105 72
rect 103 71 104 72
rect 102 71 103 72
rect 101 71 102 72
rect 100 71 101 72
rect 99 71 100 72
rect 98 71 99 72
rect 97 71 98 72
rect 96 71 97 72
rect 95 71 96 72
rect 94 71 95 72
rect 87 71 88 72
rect 86 71 87 72
rect 85 71 86 72
rect 84 71 85 72
rect 83 71 84 72
rect 82 71 83 72
rect 81 71 82 72
rect 80 71 81 72
rect 79 71 80 72
rect 78 71 79 72
rect 77 71 78 72
rect 76 71 77 72
rect 75 71 76 72
rect 74 71 75 72
rect 73 71 74 72
rect 72 71 73 72
rect 71 71 72 72
rect 70 71 71 72
rect 69 71 70 72
rect 68 71 69 72
rect 67 71 68 72
rect 66 71 67 72
rect 65 71 66 72
rect 64 71 65 72
rect 63 71 64 72
rect 62 71 63 72
rect 61 71 62 72
rect 60 71 61 72
rect 59 71 60 72
rect 58 71 59 72
rect 57 71 58 72
rect 27 71 28 72
rect 26 71 27 72
rect 25 71 26 72
rect 24 71 25 72
rect 23 71 24 72
rect 22 71 23 72
rect 21 71 22 72
rect 20 71 21 72
rect 19 71 20 72
rect 18 71 19 72
rect 17 71 18 72
rect 16 71 17 72
rect 12 71 13 72
rect 11 71 12 72
rect 10 71 11 72
rect 9 71 10 72
rect 8 71 9 72
rect 7 71 8 72
rect 195 72 196 73
rect 194 72 195 73
rect 193 72 194 73
rect 192 72 193 73
rect 178 72 179 73
rect 168 72 169 73
rect 167 72 168 73
rect 166 72 167 73
rect 165 72 166 73
rect 164 72 165 73
rect 163 72 164 73
rect 111 72 112 73
rect 110 72 111 73
rect 109 72 110 73
rect 108 72 109 73
rect 107 72 108 73
rect 106 72 107 73
rect 105 72 106 73
rect 104 72 105 73
rect 103 72 104 73
rect 102 72 103 73
rect 101 72 102 73
rect 100 72 101 73
rect 99 72 100 73
rect 98 72 99 73
rect 97 72 98 73
rect 96 72 97 73
rect 95 72 96 73
rect 94 72 95 73
rect 86 72 87 73
rect 85 72 86 73
rect 84 72 85 73
rect 83 72 84 73
rect 82 72 83 73
rect 81 72 82 73
rect 80 72 81 73
rect 79 72 80 73
rect 78 72 79 73
rect 77 72 78 73
rect 76 72 77 73
rect 75 72 76 73
rect 74 72 75 73
rect 73 72 74 73
rect 72 72 73 73
rect 71 72 72 73
rect 70 72 71 73
rect 69 72 70 73
rect 68 72 69 73
rect 67 72 68 73
rect 66 72 67 73
rect 65 72 66 73
rect 64 72 65 73
rect 63 72 64 73
rect 62 72 63 73
rect 61 72 62 73
rect 60 72 61 73
rect 59 72 60 73
rect 58 72 59 73
rect 57 72 58 73
rect 56 72 57 73
rect 55 72 56 73
rect 26 72 27 73
rect 25 72 26 73
rect 24 72 25 73
rect 23 72 24 73
rect 22 72 23 73
rect 21 72 22 73
rect 20 72 21 73
rect 19 72 20 73
rect 18 72 19 73
rect 17 72 18 73
rect 12 72 13 73
rect 11 72 12 73
rect 10 72 11 73
rect 9 72 10 73
rect 8 72 9 73
rect 7 72 8 73
rect 193 73 194 74
rect 192 73 193 74
rect 191 73 192 74
rect 169 73 170 74
rect 168 73 169 74
rect 167 73 168 74
rect 166 73 167 74
rect 165 73 166 74
rect 164 73 165 74
rect 110 73 111 74
rect 109 73 110 74
rect 108 73 109 74
rect 107 73 108 74
rect 106 73 107 74
rect 105 73 106 74
rect 104 73 105 74
rect 103 73 104 74
rect 102 73 103 74
rect 101 73 102 74
rect 100 73 101 74
rect 99 73 100 74
rect 98 73 99 74
rect 97 73 98 74
rect 96 73 97 74
rect 95 73 96 74
rect 94 73 95 74
rect 93 73 94 74
rect 85 73 86 74
rect 84 73 85 74
rect 83 73 84 74
rect 82 73 83 74
rect 81 73 82 74
rect 80 73 81 74
rect 79 73 80 74
rect 78 73 79 74
rect 77 73 78 74
rect 76 73 77 74
rect 75 73 76 74
rect 74 73 75 74
rect 73 73 74 74
rect 72 73 73 74
rect 71 73 72 74
rect 70 73 71 74
rect 69 73 70 74
rect 68 73 69 74
rect 67 73 68 74
rect 66 73 67 74
rect 65 73 66 74
rect 64 73 65 74
rect 63 73 64 74
rect 62 73 63 74
rect 61 73 62 74
rect 60 73 61 74
rect 59 73 60 74
rect 58 73 59 74
rect 57 73 58 74
rect 56 73 57 74
rect 55 73 56 74
rect 54 73 55 74
rect 26 73 27 74
rect 25 73 26 74
rect 24 73 25 74
rect 23 73 24 74
rect 22 73 23 74
rect 21 73 22 74
rect 20 73 21 74
rect 19 73 20 74
rect 18 73 19 74
rect 17 73 18 74
rect 12 73 13 74
rect 11 73 12 74
rect 10 73 11 74
rect 9 73 10 74
rect 8 73 9 74
rect 191 74 192 75
rect 190 74 191 75
rect 189 74 190 75
rect 188 74 189 75
rect 187 74 188 75
rect 170 74 171 75
rect 169 74 170 75
rect 168 74 169 75
rect 167 74 168 75
rect 166 74 167 75
rect 165 74 166 75
rect 109 74 110 75
rect 108 74 109 75
rect 107 74 108 75
rect 106 74 107 75
rect 105 74 106 75
rect 104 74 105 75
rect 103 74 104 75
rect 102 74 103 75
rect 101 74 102 75
rect 100 74 101 75
rect 99 74 100 75
rect 98 74 99 75
rect 97 74 98 75
rect 96 74 97 75
rect 95 74 96 75
rect 94 74 95 75
rect 93 74 94 75
rect 85 74 86 75
rect 84 74 85 75
rect 83 74 84 75
rect 82 74 83 75
rect 81 74 82 75
rect 80 74 81 75
rect 79 74 80 75
rect 78 74 79 75
rect 77 74 78 75
rect 76 74 77 75
rect 75 74 76 75
rect 74 74 75 75
rect 73 74 74 75
rect 72 74 73 75
rect 71 74 72 75
rect 70 74 71 75
rect 69 74 70 75
rect 68 74 69 75
rect 67 74 68 75
rect 66 74 67 75
rect 65 74 66 75
rect 64 74 65 75
rect 63 74 64 75
rect 62 74 63 75
rect 61 74 62 75
rect 60 74 61 75
rect 59 74 60 75
rect 58 74 59 75
rect 57 74 58 75
rect 56 74 57 75
rect 55 74 56 75
rect 54 74 55 75
rect 53 74 54 75
rect 52 74 53 75
rect 25 74 26 75
rect 24 74 25 75
rect 23 74 24 75
rect 22 74 23 75
rect 21 74 22 75
rect 20 74 21 75
rect 19 74 20 75
rect 18 74 19 75
rect 12 74 13 75
rect 11 74 12 75
rect 10 74 11 75
rect 9 74 10 75
rect 8 74 9 75
rect 188 75 189 76
rect 187 75 188 76
rect 172 75 173 76
rect 171 75 172 76
rect 170 75 171 76
rect 169 75 170 76
rect 168 75 169 76
rect 167 75 168 76
rect 166 75 167 76
rect 129 75 130 76
rect 128 75 129 76
rect 127 75 128 76
rect 126 75 127 76
rect 125 75 126 76
rect 124 75 125 76
rect 108 75 109 76
rect 107 75 108 76
rect 106 75 107 76
rect 105 75 106 76
rect 104 75 105 76
rect 103 75 104 76
rect 102 75 103 76
rect 101 75 102 76
rect 100 75 101 76
rect 99 75 100 76
rect 98 75 99 76
rect 97 75 98 76
rect 96 75 97 76
rect 95 75 96 76
rect 94 75 95 76
rect 93 75 94 76
rect 92 75 93 76
rect 84 75 85 76
rect 83 75 84 76
rect 82 75 83 76
rect 81 75 82 76
rect 80 75 81 76
rect 79 75 80 76
rect 78 75 79 76
rect 77 75 78 76
rect 76 75 77 76
rect 75 75 76 76
rect 74 75 75 76
rect 73 75 74 76
rect 72 75 73 76
rect 71 75 72 76
rect 70 75 71 76
rect 69 75 70 76
rect 68 75 69 76
rect 67 75 68 76
rect 66 75 67 76
rect 65 75 66 76
rect 64 75 65 76
rect 63 75 64 76
rect 62 75 63 76
rect 61 75 62 76
rect 60 75 61 76
rect 59 75 60 76
rect 58 75 59 76
rect 57 75 58 76
rect 56 75 57 76
rect 55 75 56 76
rect 54 75 55 76
rect 53 75 54 76
rect 52 75 53 76
rect 51 75 52 76
rect 50 75 51 76
rect 49 75 50 76
rect 24 75 25 76
rect 23 75 24 76
rect 22 75 23 76
rect 21 75 22 76
rect 20 75 21 76
rect 19 75 20 76
rect 18 75 19 76
rect 12 75 13 76
rect 11 75 12 76
rect 10 75 11 76
rect 9 75 10 76
rect 8 75 9 76
rect 173 76 174 77
rect 172 76 173 77
rect 171 76 172 77
rect 170 76 171 77
rect 169 76 170 77
rect 168 76 169 77
rect 133 76 134 77
rect 132 76 133 77
rect 131 76 132 77
rect 130 76 131 77
rect 129 76 130 77
rect 128 76 129 77
rect 127 76 128 77
rect 126 76 127 77
rect 125 76 126 77
rect 124 76 125 77
rect 123 76 124 77
rect 122 76 123 77
rect 121 76 122 77
rect 120 76 121 77
rect 107 76 108 77
rect 106 76 107 77
rect 105 76 106 77
rect 104 76 105 77
rect 103 76 104 77
rect 102 76 103 77
rect 101 76 102 77
rect 100 76 101 77
rect 99 76 100 77
rect 98 76 99 77
rect 97 76 98 77
rect 96 76 97 77
rect 95 76 96 77
rect 94 76 95 77
rect 93 76 94 77
rect 92 76 93 77
rect 83 76 84 77
rect 82 76 83 77
rect 81 76 82 77
rect 80 76 81 77
rect 79 76 80 77
rect 78 76 79 77
rect 77 76 78 77
rect 76 76 77 77
rect 75 76 76 77
rect 74 76 75 77
rect 73 76 74 77
rect 72 76 73 77
rect 71 76 72 77
rect 70 76 71 77
rect 69 76 70 77
rect 68 76 69 77
rect 67 76 68 77
rect 66 76 67 77
rect 65 76 66 77
rect 64 76 65 77
rect 63 76 64 77
rect 62 76 63 77
rect 61 76 62 77
rect 60 76 61 77
rect 59 76 60 77
rect 58 76 59 77
rect 57 76 58 77
rect 56 76 57 77
rect 55 76 56 77
rect 54 76 55 77
rect 53 76 54 77
rect 52 76 53 77
rect 51 76 52 77
rect 50 76 51 77
rect 49 76 50 77
rect 48 76 49 77
rect 47 76 48 77
rect 46 76 47 77
rect 33 76 34 77
rect 32 76 33 77
rect 31 76 32 77
rect 22 76 23 77
rect 21 76 22 77
rect 20 76 21 77
rect 12 76 13 77
rect 11 76 12 77
rect 10 76 11 77
rect 9 76 10 77
rect 8 76 9 77
rect 174 77 175 78
rect 173 77 174 78
rect 172 77 173 78
rect 171 77 172 78
rect 170 77 171 78
rect 169 77 170 78
rect 135 77 136 78
rect 134 77 135 78
rect 133 77 134 78
rect 132 77 133 78
rect 131 77 132 78
rect 130 77 131 78
rect 129 77 130 78
rect 128 77 129 78
rect 127 77 128 78
rect 126 77 127 78
rect 125 77 126 78
rect 124 77 125 78
rect 123 77 124 78
rect 122 77 123 78
rect 121 77 122 78
rect 120 77 121 78
rect 119 77 120 78
rect 118 77 119 78
rect 117 77 118 78
rect 107 77 108 78
rect 106 77 107 78
rect 105 77 106 78
rect 104 77 105 78
rect 103 77 104 78
rect 102 77 103 78
rect 101 77 102 78
rect 100 77 101 78
rect 99 77 100 78
rect 98 77 99 78
rect 97 77 98 78
rect 96 77 97 78
rect 95 77 96 78
rect 94 77 95 78
rect 93 77 94 78
rect 92 77 93 78
rect 91 77 92 78
rect 82 77 83 78
rect 81 77 82 78
rect 80 77 81 78
rect 79 77 80 78
rect 78 77 79 78
rect 77 77 78 78
rect 76 77 77 78
rect 75 77 76 78
rect 74 77 75 78
rect 73 77 74 78
rect 72 77 73 78
rect 71 77 72 78
rect 70 77 71 78
rect 69 77 70 78
rect 68 77 69 78
rect 67 77 68 78
rect 66 77 67 78
rect 65 77 66 78
rect 64 77 65 78
rect 63 77 64 78
rect 62 77 63 78
rect 61 77 62 78
rect 60 77 61 78
rect 59 77 60 78
rect 58 77 59 78
rect 57 77 58 78
rect 56 77 57 78
rect 55 77 56 78
rect 54 77 55 78
rect 53 77 54 78
rect 52 77 53 78
rect 51 77 52 78
rect 50 77 51 78
rect 49 77 50 78
rect 48 77 49 78
rect 47 77 48 78
rect 46 77 47 78
rect 45 77 46 78
rect 44 77 45 78
rect 43 77 44 78
rect 42 77 43 78
rect 41 77 42 78
rect 40 77 41 78
rect 39 77 40 78
rect 38 77 39 78
rect 36 77 37 78
rect 35 77 36 78
rect 34 77 35 78
rect 33 77 34 78
rect 32 77 33 78
rect 31 77 32 78
rect 13 77 14 78
rect 12 77 13 78
rect 11 77 12 78
rect 10 77 11 78
rect 9 77 10 78
rect 8 77 9 78
rect 175 78 176 79
rect 174 78 175 79
rect 173 78 174 79
rect 172 78 173 79
rect 171 78 172 79
rect 170 78 171 79
rect 161 78 162 79
rect 136 78 137 79
rect 135 78 136 79
rect 134 78 135 79
rect 133 78 134 79
rect 132 78 133 79
rect 131 78 132 79
rect 130 78 131 79
rect 129 78 130 79
rect 128 78 129 79
rect 127 78 128 79
rect 126 78 127 79
rect 125 78 126 79
rect 124 78 125 79
rect 123 78 124 79
rect 122 78 123 79
rect 121 78 122 79
rect 120 78 121 79
rect 119 78 120 79
rect 118 78 119 79
rect 117 78 118 79
rect 116 78 117 79
rect 115 78 116 79
rect 106 78 107 79
rect 105 78 106 79
rect 104 78 105 79
rect 103 78 104 79
rect 102 78 103 79
rect 101 78 102 79
rect 100 78 101 79
rect 99 78 100 79
rect 98 78 99 79
rect 97 78 98 79
rect 96 78 97 79
rect 95 78 96 79
rect 94 78 95 79
rect 93 78 94 79
rect 92 78 93 79
rect 91 78 92 79
rect 90 78 91 79
rect 81 78 82 79
rect 80 78 81 79
rect 79 78 80 79
rect 78 78 79 79
rect 77 78 78 79
rect 76 78 77 79
rect 75 78 76 79
rect 74 78 75 79
rect 73 78 74 79
rect 72 78 73 79
rect 71 78 72 79
rect 70 78 71 79
rect 69 78 70 79
rect 68 78 69 79
rect 67 78 68 79
rect 66 78 67 79
rect 65 78 66 79
rect 64 78 65 79
rect 63 78 64 79
rect 62 78 63 79
rect 61 78 62 79
rect 60 78 61 79
rect 59 78 60 79
rect 58 78 59 79
rect 57 78 58 79
rect 56 78 57 79
rect 55 78 56 79
rect 54 78 55 79
rect 53 78 54 79
rect 52 78 53 79
rect 51 78 52 79
rect 50 78 51 79
rect 49 78 50 79
rect 48 78 49 79
rect 47 78 48 79
rect 46 78 47 79
rect 45 78 46 79
rect 44 78 45 79
rect 43 78 44 79
rect 42 78 43 79
rect 41 78 42 79
rect 40 78 41 79
rect 39 78 40 79
rect 38 78 39 79
rect 37 78 38 79
rect 36 78 37 79
rect 35 78 36 79
rect 34 78 35 79
rect 33 78 34 79
rect 32 78 33 79
rect 31 78 32 79
rect 13 78 14 79
rect 12 78 13 79
rect 11 78 12 79
rect 10 78 11 79
rect 9 78 10 79
rect 8 78 9 79
rect 177 79 178 80
rect 176 79 177 80
rect 175 79 176 80
rect 174 79 175 80
rect 173 79 174 80
rect 172 79 173 80
rect 171 79 172 80
rect 161 79 162 80
rect 138 79 139 80
rect 137 79 138 80
rect 136 79 137 80
rect 135 79 136 80
rect 134 79 135 80
rect 133 79 134 80
rect 132 79 133 80
rect 131 79 132 80
rect 130 79 131 80
rect 129 79 130 80
rect 128 79 129 80
rect 127 79 128 80
rect 126 79 127 80
rect 125 79 126 80
rect 124 79 125 80
rect 123 79 124 80
rect 122 79 123 80
rect 121 79 122 80
rect 120 79 121 80
rect 119 79 120 80
rect 118 79 119 80
rect 117 79 118 80
rect 116 79 117 80
rect 115 79 116 80
rect 114 79 115 80
rect 113 79 114 80
rect 105 79 106 80
rect 104 79 105 80
rect 103 79 104 80
rect 102 79 103 80
rect 101 79 102 80
rect 100 79 101 80
rect 99 79 100 80
rect 98 79 99 80
rect 97 79 98 80
rect 96 79 97 80
rect 95 79 96 80
rect 94 79 95 80
rect 93 79 94 80
rect 92 79 93 80
rect 91 79 92 80
rect 90 79 91 80
rect 80 79 81 80
rect 79 79 80 80
rect 78 79 79 80
rect 77 79 78 80
rect 76 79 77 80
rect 75 79 76 80
rect 74 79 75 80
rect 73 79 74 80
rect 72 79 73 80
rect 71 79 72 80
rect 70 79 71 80
rect 69 79 70 80
rect 68 79 69 80
rect 67 79 68 80
rect 66 79 67 80
rect 65 79 66 80
rect 64 79 65 80
rect 63 79 64 80
rect 62 79 63 80
rect 61 79 62 80
rect 60 79 61 80
rect 59 79 60 80
rect 58 79 59 80
rect 57 79 58 80
rect 56 79 57 80
rect 55 79 56 80
rect 54 79 55 80
rect 53 79 54 80
rect 52 79 53 80
rect 51 79 52 80
rect 50 79 51 80
rect 49 79 50 80
rect 48 79 49 80
rect 47 79 48 80
rect 46 79 47 80
rect 45 79 46 80
rect 44 79 45 80
rect 43 79 44 80
rect 42 79 43 80
rect 41 79 42 80
rect 40 79 41 80
rect 39 79 40 80
rect 38 79 39 80
rect 37 79 38 80
rect 36 79 37 80
rect 35 79 36 80
rect 34 79 35 80
rect 33 79 34 80
rect 32 79 33 80
rect 31 79 32 80
rect 14 79 15 80
rect 13 79 14 80
rect 12 79 13 80
rect 11 79 12 80
rect 10 79 11 80
rect 9 79 10 80
rect 8 79 9 80
rect 195 80 196 81
rect 194 80 195 81
rect 187 80 188 81
rect 178 80 179 81
rect 177 80 178 81
rect 176 80 177 81
rect 175 80 176 81
rect 174 80 175 81
rect 173 80 174 81
rect 172 80 173 81
rect 162 80 163 81
rect 161 80 162 81
rect 139 80 140 81
rect 138 80 139 81
rect 137 80 138 81
rect 136 80 137 81
rect 135 80 136 81
rect 134 80 135 81
rect 133 80 134 81
rect 132 80 133 81
rect 131 80 132 81
rect 130 80 131 81
rect 129 80 130 81
rect 128 80 129 81
rect 127 80 128 81
rect 126 80 127 81
rect 125 80 126 81
rect 124 80 125 81
rect 123 80 124 81
rect 122 80 123 81
rect 121 80 122 81
rect 120 80 121 81
rect 119 80 120 81
rect 118 80 119 81
rect 117 80 118 81
rect 116 80 117 81
rect 115 80 116 81
rect 114 80 115 81
rect 113 80 114 81
rect 112 80 113 81
rect 105 80 106 81
rect 104 80 105 81
rect 103 80 104 81
rect 102 80 103 81
rect 101 80 102 81
rect 100 80 101 81
rect 99 80 100 81
rect 98 80 99 81
rect 97 80 98 81
rect 96 80 97 81
rect 95 80 96 81
rect 94 80 95 81
rect 93 80 94 81
rect 92 80 93 81
rect 91 80 92 81
rect 90 80 91 81
rect 89 80 90 81
rect 79 80 80 81
rect 78 80 79 81
rect 77 80 78 81
rect 76 80 77 81
rect 75 80 76 81
rect 74 80 75 81
rect 73 80 74 81
rect 72 80 73 81
rect 71 80 72 81
rect 70 80 71 81
rect 69 80 70 81
rect 68 80 69 81
rect 67 80 68 81
rect 66 80 67 81
rect 65 80 66 81
rect 64 80 65 81
rect 63 80 64 81
rect 62 80 63 81
rect 61 80 62 81
rect 60 80 61 81
rect 59 80 60 81
rect 58 80 59 81
rect 57 80 58 81
rect 56 80 57 81
rect 55 80 56 81
rect 54 80 55 81
rect 53 80 54 81
rect 52 80 53 81
rect 51 80 52 81
rect 50 80 51 81
rect 49 80 50 81
rect 48 80 49 81
rect 47 80 48 81
rect 46 80 47 81
rect 45 80 46 81
rect 44 80 45 81
rect 43 80 44 81
rect 42 80 43 81
rect 41 80 42 81
rect 40 80 41 81
rect 39 80 40 81
rect 38 80 39 81
rect 37 80 38 81
rect 36 80 37 81
rect 35 80 36 81
rect 34 80 35 81
rect 33 80 34 81
rect 32 80 33 81
rect 31 80 32 81
rect 14 80 15 81
rect 13 80 14 81
rect 12 80 13 81
rect 11 80 12 81
rect 10 80 11 81
rect 9 80 10 81
rect 8 80 9 81
rect 194 81 195 82
rect 193 81 194 82
rect 192 81 193 82
rect 191 81 192 82
rect 190 81 191 82
rect 189 81 190 82
rect 188 81 189 82
rect 187 81 188 82
rect 179 81 180 82
rect 178 81 179 82
rect 177 81 178 82
rect 176 81 177 82
rect 175 81 176 82
rect 174 81 175 82
rect 173 81 174 82
rect 172 81 173 82
rect 171 81 172 82
rect 170 81 171 82
rect 169 81 170 82
rect 168 81 169 82
rect 167 81 168 82
rect 166 81 167 82
rect 165 81 166 82
rect 164 81 165 82
rect 163 81 164 82
rect 162 81 163 82
rect 161 81 162 82
rect 140 81 141 82
rect 139 81 140 82
rect 138 81 139 82
rect 137 81 138 82
rect 136 81 137 82
rect 135 81 136 82
rect 134 81 135 82
rect 133 81 134 82
rect 132 81 133 82
rect 131 81 132 82
rect 130 81 131 82
rect 129 81 130 82
rect 128 81 129 82
rect 127 81 128 82
rect 126 81 127 82
rect 125 81 126 82
rect 124 81 125 82
rect 123 81 124 82
rect 122 81 123 82
rect 121 81 122 82
rect 120 81 121 82
rect 119 81 120 82
rect 118 81 119 82
rect 117 81 118 82
rect 116 81 117 82
rect 115 81 116 82
rect 114 81 115 82
rect 113 81 114 82
rect 112 81 113 82
rect 111 81 112 82
rect 104 81 105 82
rect 103 81 104 82
rect 102 81 103 82
rect 101 81 102 82
rect 100 81 101 82
rect 99 81 100 82
rect 98 81 99 82
rect 97 81 98 82
rect 96 81 97 82
rect 95 81 96 82
rect 94 81 95 82
rect 93 81 94 82
rect 92 81 93 82
rect 91 81 92 82
rect 90 81 91 82
rect 89 81 90 82
rect 88 81 89 82
rect 78 81 79 82
rect 77 81 78 82
rect 76 81 77 82
rect 75 81 76 82
rect 74 81 75 82
rect 73 81 74 82
rect 72 81 73 82
rect 71 81 72 82
rect 70 81 71 82
rect 69 81 70 82
rect 68 81 69 82
rect 67 81 68 82
rect 66 81 67 82
rect 65 81 66 82
rect 64 81 65 82
rect 63 81 64 82
rect 62 81 63 82
rect 61 81 62 82
rect 60 81 61 82
rect 59 81 60 82
rect 58 81 59 82
rect 57 81 58 82
rect 56 81 57 82
rect 55 81 56 82
rect 54 81 55 82
rect 53 81 54 82
rect 52 81 53 82
rect 51 81 52 82
rect 50 81 51 82
rect 49 81 50 82
rect 48 81 49 82
rect 47 81 48 82
rect 46 81 47 82
rect 45 81 46 82
rect 44 81 45 82
rect 43 81 44 82
rect 42 81 43 82
rect 41 81 42 82
rect 40 81 41 82
rect 39 81 40 82
rect 38 81 39 82
rect 37 81 38 82
rect 36 81 37 82
rect 35 81 36 82
rect 34 81 35 82
rect 33 81 34 82
rect 32 81 33 82
rect 31 81 32 82
rect 23 81 24 82
rect 22 81 23 82
rect 21 81 22 82
rect 15 81 16 82
rect 14 81 15 82
rect 13 81 14 82
rect 12 81 13 82
rect 11 81 12 82
rect 10 81 11 82
rect 9 81 10 82
rect 8 81 9 82
rect 195 82 196 83
rect 194 82 195 83
rect 193 82 194 83
rect 192 82 193 83
rect 191 82 192 83
rect 190 82 191 83
rect 189 82 190 83
rect 188 82 189 83
rect 187 82 188 83
rect 178 82 179 83
rect 177 82 178 83
rect 176 82 177 83
rect 175 82 176 83
rect 174 82 175 83
rect 173 82 174 83
rect 172 82 173 83
rect 171 82 172 83
rect 170 82 171 83
rect 169 82 170 83
rect 168 82 169 83
rect 167 82 168 83
rect 166 82 167 83
rect 165 82 166 83
rect 164 82 165 83
rect 163 82 164 83
rect 162 82 163 83
rect 161 82 162 83
rect 141 82 142 83
rect 140 82 141 83
rect 139 82 140 83
rect 138 82 139 83
rect 137 82 138 83
rect 136 82 137 83
rect 135 82 136 83
rect 134 82 135 83
rect 133 82 134 83
rect 132 82 133 83
rect 131 82 132 83
rect 130 82 131 83
rect 129 82 130 83
rect 128 82 129 83
rect 127 82 128 83
rect 126 82 127 83
rect 125 82 126 83
rect 124 82 125 83
rect 123 82 124 83
rect 122 82 123 83
rect 121 82 122 83
rect 120 82 121 83
rect 119 82 120 83
rect 118 82 119 83
rect 117 82 118 83
rect 116 82 117 83
rect 115 82 116 83
rect 114 82 115 83
rect 113 82 114 83
rect 112 82 113 83
rect 111 82 112 83
rect 110 82 111 83
rect 109 82 110 83
rect 104 82 105 83
rect 103 82 104 83
rect 102 82 103 83
rect 101 82 102 83
rect 100 82 101 83
rect 99 82 100 83
rect 98 82 99 83
rect 97 82 98 83
rect 96 82 97 83
rect 95 82 96 83
rect 94 82 95 83
rect 93 82 94 83
rect 92 82 93 83
rect 91 82 92 83
rect 90 82 91 83
rect 89 82 90 83
rect 88 82 89 83
rect 77 82 78 83
rect 76 82 77 83
rect 75 82 76 83
rect 74 82 75 83
rect 73 82 74 83
rect 72 82 73 83
rect 71 82 72 83
rect 70 82 71 83
rect 69 82 70 83
rect 68 82 69 83
rect 67 82 68 83
rect 66 82 67 83
rect 65 82 66 83
rect 64 82 65 83
rect 63 82 64 83
rect 62 82 63 83
rect 61 82 62 83
rect 60 82 61 83
rect 59 82 60 83
rect 58 82 59 83
rect 57 82 58 83
rect 56 82 57 83
rect 55 82 56 83
rect 54 82 55 83
rect 53 82 54 83
rect 52 82 53 83
rect 51 82 52 83
rect 50 82 51 83
rect 49 82 50 83
rect 48 82 49 83
rect 47 82 48 83
rect 46 82 47 83
rect 45 82 46 83
rect 44 82 45 83
rect 43 82 44 83
rect 42 82 43 83
rect 41 82 42 83
rect 40 82 41 83
rect 39 82 40 83
rect 38 82 39 83
rect 37 82 38 83
rect 36 82 37 83
rect 35 82 36 83
rect 34 82 35 83
rect 33 82 34 83
rect 32 82 33 83
rect 31 82 32 83
rect 24 82 25 83
rect 23 82 24 83
rect 22 82 23 83
rect 21 82 22 83
rect 20 82 21 83
rect 19 82 20 83
rect 18 82 19 83
rect 17 82 18 83
rect 16 82 17 83
rect 15 82 16 83
rect 14 82 15 83
rect 13 82 14 83
rect 12 82 13 83
rect 11 82 12 83
rect 10 82 11 83
rect 9 82 10 83
rect 8 82 9 83
rect 195 83 196 84
rect 191 83 192 84
rect 190 83 191 84
rect 162 83 163 84
rect 161 83 162 84
rect 142 83 143 84
rect 141 83 142 84
rect 140 83 141 84
rect 139 83 140 84
rect 138 83 139 84
rect 137 83 138 84
rect 136 83 137 84
rect 135 83 136 84
rect 134 83 135 84
rect 133 83 134 84
rect 132 83 133 84
rect 131 83 132 84
rect 130 83 131 84
rect 129 83 130 84
rect 128 83 129 84
rect 127 83 128 84
rect 126 83 127 84
rect 125 83 126 84
rect 124 83 125 84
rect 123 83 124 84
rect 122 83 123 84
rect 121 83 122 84
rect 120 83 121 84
rect 119 83 120 84
rect 118 83 119 84
rect 117 83 118 84
rect 116 83 117 84
rect 115 83 116 84
rect 114 83 115 84
rect 113 83 114 84
rect 112 83 113 84
rect 111 83 112 84
rect 110 83 111 84
rect 109 83 110 84
rect 108 83 109 84
rect 103 83 104 84
rect 102 83 103 84
rect 101 83 102 84
rect 100 83 101 84
rect 99 83 100 84
rect 98 83 99 84
rect 97 83 98 84
rect 96 83 97 84
rect 95 83 96 84
rect 94 83 95 84
rect 93 83 94 84
rect 92 83 93 84
rect 91 83 92 84
rect 90 83 91 84
rect 89 83 90 84
rect 88 83 89 84
rect 87 83 88 84
rect 76 83 77 84
rect 75 83 76 84
rect 74 83 75 84
rect 73 83 74 84
rect 72 83 73 84
rect 71 83 72 84
rect 70 83 71 84
rect 69 83 70 84
rect 68 83 69 84
rect 67 83 68 84
rect 66 83 67 84
rect 65 83 66 84
rect 64 83 65 84
rect 63 83 64 84
rect 62 83 63 84
rect 61 83 62 84
rect 60 83 61 84
rect 59 83 60 84
rect 58 83 59 84
rect 57 83 58 84
rect 56 83 57 84
rect 55 83 56 84
rect 54 83 55 84
rect 53 83 54 84
rect 52 83 53 84
rect 51 83 52 84
rect 50 83 51 84
rect 49 83 50 84
rect 48 83 49 84
rect 47 83 48 84
rect 46 83 47 84
rect 45 83 46 84
rect 44 83 45 84
rect 43 83 44 84
rect 42 83 43 84
rect 41 83 42 84
rect 40 83 41 84
rect 39 83 40 84
rect 38 83 39 84
rect 37 83 38 84
rect 36 83 37 84
rect 35 83 36 84
rect 34 83 35 84
rect 33 83 34 84
rect 32 83 33 84
rect 25 83 26 84
rect 24 83 25 84
rect 23 83 24 84
rect 22 83 23 84
rect 21 83 22 84
rect 20 83 21 84
rect 19 83 20 84
rect 18 83 19 84
rect 17 83 18 84
rect 16 83 17 84
rect 15 83 16 84
rect 14 83 15 84
rect 13 83 14 84
rect 12 83 13 84
rect 11 83 12 84
rect 10 83 11 84
rect 9 83 10 84
rect 8 83 9 84
rect 191 84 192 85
rect 190 84 191 85
rect 187 84 188 85
rect 161 84 162 85
rect 143 84 144 85
rect 142 84 143 85
rect 141 84 142 85
rect 140 84 141 85
rect 139 84 140 85
rect 138 84 139 85
rect 137 84 138 85
rect 136 84 137 85
rect 135 84 136 85
rect 134 84 135 85
rect 133 84 134 85
rect 132 84 133 85
rect 131 84 132 85
rect 130 84 131 85
rect 129 84 130 85
rect 128 84 129 85
rect 127 84 128 85
rect 126 84 127 85
rect 125 84 126 85
rect 124 84 125 85
rect 123 84 124 85
rect 122 84 123 85
rect 121 84 122 85
rect 120 84 121 85
rect 119 84 120 85
rect 118 84 119 85
rect 117 84 118 85
rect 116 84 117 85
rect 115 84 116 85
rect 114 84 115 85
rect 113 84 114 85
rect 112 84 113 85
rect 111 84 112 85
rect 110 84 111 85
rect 109 84 110 85
rect 108 84 109 85
rect 107 84 108 85
rect 106 84 107 85
rect 102 84 103 85
rect 101 84 102 85
rect 100 84 101 85
rect 99 84 100 85
rect 98 84 99 85
rect 97 84 98 85
rect 96 84 97 85
rect 95 84 96 85
rect 94 84 95 85
rect 93 84 94 85
rect 92 84 93 85
rect 91 84 92 85
rect 90 84 91 85
rect 89 84 90 85
rect 88 84 89 85
rect 87 84 88 85
rect 86 84 87 85
rect 75 84 76 85
rect 74 84 75 85
rect 73 84 74 85
rect 72 84 73 85
rect 71 84 72 85
rect 70 84 71 85
rect 69 84 70 85
rect 68 84 69 85
rect 67 84 68 85
rect 66 84 67 85
rect 65 84 66 85
rect 64 84 65 85
rect 63 84 64 85
rect 62 84 63 85
rect 61 84 62 85
rect 60 84 61 85
rect 59 84 60 85
rect 58 84 59 85
rect 57 84 58 85
rect 56 84 57 85
rect 55 84 56 85
rect 54 84 55 85
rect 53 84 54 85
rect 52 84 53 85
rect 51 84 52 85
rect 50 84 51 85
rect 49 84 50 85
rect 48 84 49 85
rect 47 84 48 85
rect 46 84 47 85
rect 45 84 46 85
rect 44 84 45 85
rect 43 84 44 85
rect 42 84 43 85
rect 41 84 42 85
rect 40 84 41 85
rect 39 84 40 85
rect 38 84 39 85
rect 37 84 38 85
rect 36 84 37 85
rect 35 84 36 85
rect 34 84 35 85
rect 33 84 34 85
rect 32 84 33 85
rect 25 84 26 85
rect 24 84 25 85
rect 23 84 24 85
rect 22 84 23 85
rect 21 84 22 85
rect 20 84 21 85
rect 19 84 20 85
rect 18 84 19 85
rect 17 84 18 85
rect 16 84 17 85
rect 15 84 16 85
rect 14 84 15 85
rect 13 84 14 85
rect 12 84 13 85
rect 11 84 12 85
rect 10 84 11 85
rect 9 84 10 85
rect 8 84 9 85
rect 195 85 196 86
rect 194 85 195 86
rect 191 85 192 86
rect 190 85 191 86
rect 188 85 189 86
rect 187 85 188 86
rect 144 85 145 86
rect 143 85 144 86
rect 142 85 143 86
rect 141 85 142 86
rect 140 85 141 86
rect 139 85 140 86
rect 138 85 139 86
rect 137 85 138 86
rect 136 85 137 86
rect 135 85 136 86
rect 134 85 135 86
rect 133 85 134 86
rect 132 85 133 86
rect 131 85 132 86
rect 130 85 131 86
rect 129 85 130 86
rect 128 85 129 86
rect 127 85 128 86
rect 126 85 127 86
rect 125 85 126 86
rect 124 85 125 86
rect 123 85 124 86
rect 122 85 123 86
rect 121 85 122 86
rect 120 85 121 86
rect 119 85 120 86
rect 118 85 119 86
rect 117 85 118 86
rect 116 85 117 86
rect 115 85 116 86
rect 114 85 115 86
rect 113 85 114 86
rect 112 85 113 86
rect 111 85 112 86
rect 110 85 111 86
rect 109 85 110 86
rect 108 85 109 86
rect 107 85 108 86
rect 106 85 107 86
rect 105 85 106 86
rect 102 85 103 86
rect 101 85 102 86
rect 100 85 101 86
rect 99 85 100 86
rect 98 85 99 86
rect 97 85 98 86
rect 96 85 97 86
rect 95 85 96 86
rect 94 85 95 86
rect 93 85 94 86
rect 92 85 93 86
rect 91 85 92 86
rect 90 85 91 86
rect 89 85 90 86
rect 88 85 89 86
rect 87 85 88 86
rect 86 85 87 86
rect 85 85 86 86
rect 73 85 74 86
rect 72 85 73 86
rect 71 85 72 86
rect 70 85 71 86
rect 69 85 70 86
rect 68 85 69 86
rect 67 85 68 86
rect 66 85 67 86
rect 65 85 66 86
rect 64 85 65 86
rect 63 85 64 86
rect 62 85 63 86
rect 61 85 62 86
rect 60 85 61 86
rect 59 85 60 86
rect 58 85 59 86
rect 57 85 58 86
rect 56 85 57 86
rect 55 85 56 86
rect 54 85 55 86
rect 53 85 54 86
rect 52 85 53 86
rect 51 85 52 86
rect 50 85 51 86
rect 49 85 50 86
rect 48 85 49 86
rect 47 85 48 86
rect 46 85 47 86
rect 45 85 46 86
rect 44 85 45 86
rect 43 85 44 86
rect 42 85 43 86
rect 41 85 42 86
rect 40 85 41 86
rect 39 85 40 86
rect 38 85 39 86
rect 37 85 38 86
rect 36 85 37 86
rect 35 85 36 86
rect 34 85 35 86
rect 33 85 34 86
rect 26 85 27 86
rect 25 85 26 86
rect 24 85 25 86
rect 23 85 24 86
rect 22 85 23 86
rect 21 85 22 86
rect 20 85 21 86
rect 19 85 20 86
rect 18 85 19 86
rect 17 85 18 86
rect 16 85 17 86
rect 15 85 16 86
rect 14 85 15 86
rect 13 85 14 86
rect 12 85 13 86
rect 11 85 12 86
rect 10 85 11 86
rect 9 85 10 86
rect 8 85 9 86
rect 7 85 8 86
rect 194 86 195 87
rect 193 86 194 87
rect 188 86 189 87
rect 171 86 172 87
rect 170 86 171 87
rect 169 86 170 87
rect 168 86 169 87
rect 144 86 145 87
rect 143 86 144 87
rect 142 86 143 87
rect 141 86 142 87
rect 140 86 141 87
rect 139 86 140 87
rect 138 86 139 87
rect 137 86 138 87
rect 136 86 137 87
rect 135 86 136 87
rect 134 86 135 87
rect 133 86 134 87
rect 132 86 133 87
rect 131 86 132 87
rect 130 86 131 87
rect 129 86 130 87
rect 128 86 129 87
rect 127 86 128 87
rect 126 86 127 87
rect 125 86 126 87
rect 124 86 125 87
rect 123 86 124 87
rect 122 86 123 87
rect 121 86 122 87
rect 120 86 121 87
rect 119 86 120 87
rect 118 86 119 87
rect 117 86 118 87
rect 116 86 117 87
rect 115 86 116 87
rect 114 86 115 87
rect 113 86 114 87
rect 112 86 113 87
rect 111 86 112 87
rect 110 86 111 87
rect 109 86 110 87
rect 108 86 109 87
rect 107 86 108 87
rect 106 86 107 87
rect 105 86 106 87
rect 104 86 105 87
rect 103 86 104 87
rect 102 86 103 87
rect 101 86 102 87
rect 100 86 101 87
rect 99 86 100 87
rect 98 86 99 87
rect 97 86 98 87
rect 96 86 97 87
rect 95 86 96 87
rect 94 86 95 87
rect 93 86 94 87
rect 92 86 93 87
rect 91 86 92 87
rect 90 86 91 87
rect 89 86 90 87
rect 88 86 89 87
rect 87 86 88 87
rect 86 86 87 87
rect 85 86 86 87
rect 84 86 85 87
rect 71 86 72 87
rect 70 86 71 87
rect 69 86 70 87
rect 68 86 69 87
rect 67 86 68 87
rect 66 86 67 87
rect 65 86 66 87
rect 64 86 65 87
rect 63 86 64 87
rect 62 86 63 87
rect 61 86 62 87
rect 60 86 61 87
rect 59 86 60 87
rect 58 86 59 87
rect 57 86 58 87
rect 56 86 57 87
rect 55 86 56 87
rect 54 86 55 87
rect 53 86 54 87
rect 52 86 53 87
rect 51 86 52 87
rect 50 86 51 87
rect 49 86 50 87
rect 48 86 49 87
rect 47 86 48 87
rect 46 86 47 87
rect 45 86 46 87
rect 44 86 45 87
rect 43 86 44 87
rect 42 86 43 87
rect 41 86 42 87
rect 40 86 41 87
rect 39 86 40 87
rect 38 86 39 87
rect 37 86 38 87
rect 36 86 37 87
rect 35 86 36 87
rect 34 86 35 87
rect 27 86 28 87
rect 26 86 27 87
rect 25 86 26 87
rect 24 86 25 87
rect 23 86 24 87
rect 22 86 23 87
rect 21 86 22 87
rect 20 86 21 87
rect 19 86 20 87
rect 18 86 19 87
rect 17 86 18 87
rect 16 86 17 87
rect 15 86 16 87
rect 14 86 15 87
rect 13 86 14 87
rect 12 86 13 87
rect 11 86 12 87
rect 10 86 11 87
rect 9 86 10 87
rect 8 86 9 87
rect 7 86 8 87
rect 174 87 175 88
rect 173 87 174 88
rect 172 87 173 88
rect 171 87 172 88
rect 170 87 171 88
rect 169 87 170 88
rect 168 87 169 88
rect 167 87 168 88
rect 166 87 167 88
rect 165 87 166 88
rect 145 87 146 88
rect 144 87 145 88
rect 143 87 144 88
rect 142 87 143 88
rect 141 87 142 88
rect 140 87 141 88
rect 139 87 140 88
rect 138 87 139 88
rect 137 87 138 88
rect 136 87 137 88
rect 135 87 136 88
rect 134 87 135 88
rect 133 87 134 88
rect 132 87 133 88
rect 131 87 132 88
rect 130 87 131 88
rect 129 87 130 88
rect 128 87 129 88
rect 127 87 128 88
rect 126 87 127 88
rect 125 87 126 88
rect 124 87 125 88
rect 123 87 124 88
rect 122 87 123 88
rect 121 87 122 88
rect 120 87 121 88
rect 119 87 120 88
rect 118 87 119 88
rect 117 87 118 88
rect 116 87 117 88
rect 115 87 116 88
rect 114 87 115 88
rect 113 87 114 88
rect 112 87 113 88
rect 111 87 112 88
rect 110 87 111 88
rect 109 87 110 88
rect 108 87 109 88
rect 107 87 108 88
rect 106 87 107 88
rect 105 87 106 88
rect 104 87 105 88
rect 103 87 104 88
rect 102 87 103 88
rect 101 87 102 88
rect 100 87 101 88
rect 99 87 100 88
rect 98 87 99 88
rect 97 87 98 88
rect 96 87 97 88
rect 95 87 96 88
rect 94 87 95 88
rect 93 87 94 88
rect 92 87 93 88
rect 91 87 92 88
rect 90 87 91 88
rect 89 87 90 88
rect 88 87 89 88
rect 87 87 88 88
rect 86 87 87 88
rect 85 87 86 88
rect 84 87 85 88
rect 83 87 84 88
rect 69 87 70 88
rect 68 87 69 88
rect 67 87 68 88
rect 66 87 67 88
rect 65 87 66 88
rect 64 87 65 88
rect 63 87 64 88
rect 62 87 63 88
rect 61 87 62 88
rect 60 87 61 88
rect 59 87 60 88
rect 58 87 59 88
rect 57 87 58 88
rect 56 87 57 88
rect 55 87 56 88
rect 54 87 55 88
rect 53 87 54 88
rect 52 87 53 88
rect 51 87 52 88
rect 50 87 51 88
rect 49 87 50 88
rect 48 87 49 88
rect 47 87 48 88
rect 46 87 47 88
rect 45 87 46 88
rect 44 87 45 88
rect 43 87 44 88
rect 42 87 43 88
rect 41 87 42 88
rect 40 87 41 88
rect 39 87 40 88
rect 38 87 39 88
rect 37 87 38 88
rect 36 87 37 88
rect 27 87 28 88
rect 26 87 27 88
rect 25 87 26 88
rect 24 87 25 88
rect 23 87 24 88
rect 22 87 23 88
rect 21 87 22 88
rect 20 87 21 88
rect 19 87 20 88
rect 18 87 19 88
rect 17 87 18 88
rect 16 87 17 88
rect 15 87 16 88
rect 14 87 15 88
rect 13 87 14 88
rect 12 87 13 88
rect 11 87 12 88
rect 10 87 11 88
rect 9 87 10 88
rect 8 87 9 88
rect 7 87 8 88
rect 175 88 176 89
rect 174 88 175 89
rect 173 88 174 89
rect 172 88 173 89
rect 171 88 172 89
rect 170 88 171 89
rect 169 88 170 89
rect 168 88 169 89
rect 167 88 168 89
rect 166 88 167 89
rect 165 88 166 89
rect 164 88 165 89
rect 145 88 146 89
rect 144 88 145 89
rect 143 88 144 89
rect 142 88 143 89
rect 141 88 142 89
rect 140 88 141 89
rect 139 88 140 89
rect 138 88 139 89
rect 137 88 138 89
rect 136 88 137 89
rect 135 88 136 89
rect 134 88 135 89
rect 133 88 134 89
rect 132 88 133 89
rect 131 88 132 89
rect 130 88 131 89
rect 129 88 130 89
rect 128 88 129 89
rect 127 88 128 89
rect 126 88 127 89
rect 125 88 126 89
rect 124 88 125 89
rect 123 88 124 89
rect 122 88 123 89
rect 121 88 122 89
rect 120 88 121 89
rect 119 88 120 89
rect 118 88 119 89
rect 117 88 118 89
rect 116 88 117 89
rect 115 88 116 89
rect 114 88 115 89
rect 113 88 114 89
rect 112 88 113 89
rect 111 88 112 89
rect 110 88 111 89
rect 109 88 110 89
rect 108 88 109 89
rect 107 88 108 89
rect 106 88 107 89
rect 105 88 106 89
rect 104 88 105 89
rect 103 88 104 89
rect 102 88 103 89
rect 101 88 102 89
rect 100 88 101 89
rect 99 88 100 89
rect 98 88 99 89
rect 97 88 98 89
rect 96 88 97 89
rect 95 88 96 89
rect 94 88 95 89
rect 93 88 94 89
rect 92 88 93 89
rect 91 88 92 89
rect 90 88 91 89
rect 89 88 90 89
rect 88 88 89 89
rect 87 88 88 89
rect 86 88 87 89
rect 85 88 86 89
rect 84 88 85 89
rect 83 88 84 89
rect 82 88 83 89
rect 81 88 82 89
rect 66 88 67 89
rect 65 88 66 89
rect 64 88 65 89
rect 63 88 64 89
rect 62 88 63 89
rect 61 88 62 89
rect 60 88 61 89
rect 59 88 60 89
rect 58 88 59 89
rect 57 88 58 89
rect 56 88 57 89
rect 55 88 56 89
rect 54 88 55 89
rect 53 88 54 89
rect 52 88 53 89
rect 51 88 52 89
rect 50 88 51 89
rect 49 88 50 89
rect 48 88 49 89
rect 47 88 48 89
rect 46 88 47 89
rect 45 88 46 89
rect 44 88 45 89
rect 43 88 44 89
rect 42 88 43 89
rect 41 88 42 89
rect 40 88 41 89
rect 39 88 40 89
rect 38 88 39 89
rect 37 88 38 89
rect 28 88 29 89
rect 27 88 28 89
rect 26 88 27 89
rect 25 88 26 89
rect 24 88 25 89
rect 23 88 24 89
rect 22 88 23 89
rect 21 88 22 89
rect 20 88 21 89
rect 19 88 20 89
rect 18 88 19 89
rect 17 88 18 89
rect 16 88 17 89
rect 15 88 16 89
rect 14 88 15 89
rect 13 88 14 89
rect 12 88 13 89
rect 11 88 12 89
rect 10 88 11 89
rect 9 88 10 89
rect 8 88 9 89
rect 7 88 8 89
rect 176 89 177 90
rect 175 89 176 90
rect 174 89 175 90
rect 173 89 174 90
rect 172 89 173 90
rect 171 89 172 90
rect 170 89 171 90
rect 169 89 170 90
rect 168 89 169 90
rect 167 89 168 90
rect 166 89 167 90
rect 165 89 166 90
rect 164 89 165 90
rect 163 89 164 90
rect 146 89 147 90
rect 145 89 146 90
rect 144 89 145 90
rect 143 89 144 90
rect 142 89 143 90
rect 141 89 142 90
rect 140 89 141 90
rect 139 89 140 90
rect 138 89 139 90
rect 137 89 138 90
rect 136 89 137 90
rect 135 89 136 90
rect 134 89 135 90
rect 133 89 134 90
rect 132 89 133 90
rect 131 89 132 90
rect 130 89 131 90
rect 129 89 130 90
rect 128 89 129 90
rect 127 89 128 90
rect 126 89 127 90
rect 125 89 126 90
rect 124 89 125 90
rect 123 89 124 90
rect 122 89 123 90
rect 121 89 122 90
rect 120 89 121 90
rect 119 89 120 90
rect 118 89 119 90
rect 117 89 118 90
rect 116 89 117 90
rect 115 89 116 90
rect 114 89 115 90
rect 113 89 114 90
rect 112 89 113 90
rect 111 89 112 90
rect 110 89 111 90
rect 109 89 110 90
rect 108 89 109 90
rect 107 89 108 90
rect 106 89 107 90
rect 105 89 106 90
rect 104 89 105 90
rect 103 89 104 90
rect 102 89 103 90
rect 101 89 102 90
rect 100 89 101 90
rect 99 89 100 90
rect 98 89 99 90
rect 97 89 98 90
rect 96 89 97 90
rect 95 89 96 90
rect 94 89 95 90
rect 93 89 94 90
rect 92 89 93 90
rect 91 89 92 90
rect 90 89 91 90
rect 89 89 90 90
rect 88 89 89 90
rect 87 89 88 90
rect 86 89 87 90
rect 85 89 86 90
rect 84 89 85 90
rect 83 89 84 90
rect 82 89 83 90
rect 81 89 82 90
rect 80 89 81 90
rect 63 89 64 90
rect 62 89 63 90
rect 61 89 62 90
rect 60 89 61 90
rect 59 89 60 90
rect 58 89 59 90
rect 57 89 58 90
rect 56 89 57 90
rect 55 89 56 90
rect 54 89 55 90
rect 53 89 54 90
rect 52 89 53 90
rect 51 89 52 90
rect 50 89 51 90
rect 49 89 50 90
rect 48 89 49 90
rect 47 89 48 90
rect 46 89 47 90
rect 45 89 46 90
rect 44 89 45 90
rect 43 89 44 90
rect 42 89 43 90
rect 41 89 42 90
rect 40 89 41 90
rect 39 89 40 90
rect 29 89 30 90
rect 28 89 29 90
rect 27 89 28 90
rect 26 89 27 90
rect 25 89 26 90
rect 24 89 25 90
rect 23 89 24 90
rect 22 89 23 90
rect 21 89 22 90
rect 20 89 21 90
rect 19 89 20 90
rect 18 89 19 90
rect 17 89 18 90
rect 16 89 17 90
rect 15 89 16 90
rect 14 89 15 90
rect 13 89 14 90
rect 12 89 13 90
rect 11 89 12 90
rect 10 89 11 90
rect 9 89 10 90
rect 8 89 9 90
rect 7 89 8 90
rect 6 89 7 90
rect 187 90 188 91
rect 177 90 178 91
rect 176 90 177 91
rect 175 90 176 91
rect 174 90 175 91
rect 173 90 174 91
rect 172 90 173 91
rect 171 90 172 91
rect 170 90 171 91
rect 169 90 170 91
rect 168 90 169 91
rect 167 90 168 91
rect 166 90 167 91
rect 165 90 166 91
rect 164 90 165 91
rect 163 90 164 91
rect 162 90 163 91
rect 146 90 147 91
rect 145 90 146 91
rect 144 90 145 91
rect 143 90 144 91
rect 142 90 143 91
rect 141 90 142 91
rect 140 90 141 91
rect 139 90 140 91
rect 138 90 139 91
rect 124 90 125 91
rect 123 90 124 91
rect 122 90 123 91
rect 121 90 122 91
rect 120 90 121 91
rect 119 90 120 91
rect 118 90 119 91
rect 117 90 118 91
rect 116 90 117 91
rect 115 90 116 91
rect 114 90 115 91
rect 113 90 114 91
rect 112 90 113 91
rect 111 90 112 91
rect 110 90 111 91
rect 109 90 110 91
rect 108 90 109 91
rect 107 90 108 91
rect 106 90 107 91
rect 105 90 106 91
rect 104 90 105 91
rect 103 90 104 91
rect 102 90 103 91
rect 101 90 102 91
rect 100 90 101 91
rect 99 90 100 91
rect 98 90 99 91
rect 97 90 98 91
rect 96 90 97 91
rect 95 90 96 91
rect 94 90 95 91
rect 93 90 94 91
rect 92 90 93 91
rect 91 90 92 91
rect 90 90 91 91
rect 89 90 90 91
rect 88 90 89 91
rect 87 90 88 91
rect 86 90 87 91
rect 85 90 86 91
rect 84 90 85 91
rect 83 90 84 91
rect 82 90 83 91
rect 81 90 82 91
rect 80 90 81 91
rect 79 90 80 91
rect 78 90 79 91
rect 62 90 63 91
rect 61 90 62 91
rect 60 90 61 91
rect 59 90 60 91
rect 58 90 59 91
rect 57 90 58 91
rect 56 90 57 91
rect 55 90 56 91
rect 54 90 55 91
rect 53 90 54 91
rect 52 90 53 91
rect 51 90 52 91
rect 50 90 51 91
rect 49 90 50 91
rect 48 90 49 91
rect 47 90 48 91
rect 46 90 47 91
rect 45 90 46 91
rect 44 90 45 91
rect 43 90 44 91
rect 42 90 43 91
rect 30 90 31 91
rect 29 90 30 91
rect 28 90 29 91
rect 27 90 28 91
rect 26 90 27 91
rect 25 90 26 91
rect 24 90 25 91
rect 23 90 24 91
rect 22 90 23 91
rect 21 90 22 91
rect 20 90 21 91
rect 19 90 20 91
rect 18 90 19 91
rect 17 90 18 91
rect 16 90 17 91
rect 15 90 16 91
rect 14 90 15 91
rect 13 90 14 91
rect 12 90 13 91
rect 11 90 12 91
rect 10 90 11 91
rect 9 90 10 91
rect 8 90 9 91
rect 7 90 8 91
rect 6 90 7 91
rect 195 91 196 92
rect 194 91 195 92
rect 193 91 194 92
rect 192 91 193 92
rect 191 91 192 92
rect 190 91 191 92
rect 189 91 190 92
rect 188 91 189 92
rect 187 91 188 92
rect 178 91 179 92
rect 177 91 178 92
rect 176 91 177 92
rect 175 91 176 92
rect 174 91 175 92
rect 173 91 174 92
rect 165 91 166 92
rect 164 91 165 92
rect 163 91 164 92
rect 162 91 163 92
rect 147 91 148 92
rect 146 91 147 92
rect 145 91 146 92
rect 144 91 145 92
rect 143 91 144 92
rect 142 91 143 92
rect 121 91 122 92
rect 120 91 121 92
rect 119 91 120 92
rect 118 91 119 92
rect 117 91 118 92
rect 116 91 117 92
rect 115 91 116 92
rect 114 91 115 92
rect 113 91 114 92
rect 112 91 113 92
rect 111 91 112 92
rect 110 91 111 92
rect 109 91 110 92
rect 108 91 109 92
rect 107 91 108 92
rect 106 91 107 92
rect 105 91 106 92
rect 104 91 105 92
rect 103 91 104 92
rect 102 91 103 92
rect 101 91 102 92
rect 100 91 101 92
rect 99 91 100 92
rect 98 91 99 92
rect 97 91 98 92
rect 96 91 97 92
rect 95 91 96 92
rect 94 91 95 92
rect 93 91 94 92
rect 92 91 93 92
rect 91 91 92 92
rect 90 91 91 92
rect 89 91 90 92
rect 88 91 89 92
rect 87 91 88 92
rect 86 91 87 92
rect 85 91 86 92
rect 84 91 85 92
rect 83 91 84 92
rect 82 91 83 92
rect 81 91 82 92
rect 80 91 81 92
rect 79 91 80 92
rect 78 91 79 92
rect 77 91 78 92
rect 76 91 77 92
rect 75 91 76 92
rect 61 91 62 92
rect 60 91 61 92
rect 59 91 60 92
rect 58 91 59 92
rect 57 91 58 92
rect 56 91 57 92
rect 55 91 56 92
rect 54 91 55 92
rect 53 91 54 92
rect 52 91 53 92
rect 51 91 52 92
rect 50 91 51 92
rect 49 91 50 92
rect 48 91 49 92
rect 47 91 48 92
rect 46 91 47 92
rect 45 91 46 92
rect 44 91 45 92
rect 31 91 32 92
rect 30 91 31 92
rect 29 91 30 92
rect 28 91 29 92
rect 27 91 28 92
rect 26 91 27 92
rect 25 91 26 92
rect 24 91 25 92
rect 23 91 24 92
rect 22 91 23 92
rect 21 91 22 92
rect 20 91 21 92
rect 19 91 20 92
rect 18 91 19 92
rect 17 91 18 92
rect 16 91 17 92
rect 15 91 16 92
rect 14 91 15 92
rect 13 91 14 92
rect 12 91 13 92
rect 11 91 12 92
rect 10 91 11 92
rect 9 91 10 92
rect 8 91 9 92
rect 7 91 8 92
rect 6 91 7 92
rect 195 92 196 93
rect 194 92 195 93
rect 193 92 194 93
rect 192 92 193 93
rect 191 92 192 93
rect 190 92 191 93
rect 189 92 190 93
rect 188 92 189 93
rect 187 92 188 93
rect 178 92 179 93
rect 177 92 178 93
rect 176 92 177 93
rect 175 92 176 93
rect 163 92 164 93
rect 162 92 163 93
rect 161 92 162 93
rect 147 92 148 93
rect 146 92 147 93
rect 145 92 146 93
rect 119 92 120 93
rect 118 92 119 93
rect 117 92 118 93
rect 116 92 117 93
rect 115 92 116 93
rect 114 92 115 93
rect 113 92 114 93
rect 112 92 113 93
rect 111 92 112 93
rect 110 92 111 93
rect 109 92 110 93
rect 108 92 109 93
rect 107 92 108 93
rect 106 92 107 93
rect 105 92 106 93
rect 104 92 105 93
rect 103 92 104 93
rect 102 92 103 93
rect 101 92 102 93
rect 100 92 101 93
rect 99 92 100 93
rect 98 92 99 93
rect 97 92 98 93
rect 96 92 97 93
rect 95 92 96 93
rect 94 92 95 93
rect 93 92 94 93
rect 92 92 93 93
rect 91 92 92 93
rect 90 92 91 93
rect 89 92 90 93
rect 88 92 89 93
rect 87 92 88 93
rect 86 92 87 93
rect 85 92 86 93
rect 84 92 85 93
rect 83 92 84 93
rect 82 92 83 93
rect 81 92 82 93
rect 80 92 81 93
rect 79 92 80 93
rect 78 92 79 93
rect 77 92 78 93
rect 76 92 77 93
rect 75 92 76 93
rect 74 92 75 93
rect 73 92 74 93
rect 61 92 62 93
rect 60 92 61 93
rect 59 92 60 93
rect 58 92 59 93
rect 57 92 58 93
rect 56 92 57 93
rect 55 92 56 93
rect 54 92 55 93
rect 53 92 54 93
rect 52 92 53 93
rect 51 92 52 93
rect 50 92 51 93
rect 49 92 50 93
rect 48 92 49 93
rect 47 92 48 93
rect 46 92 47 93
rect 45 92 46 93
rect 32 92 33 93
rect 31 92 32 93
rect 30 92 31 93
rect 29 92 30 93
rect 28 92 29 93
rect 27 92 28 93
rect 26 92 27 93
rect 25 92 26 93
rect 24 92 25 93
rect 23 92 24 93
rect 22 92 23 93
rect 21 92 22 93
rect 20 92 21 93
rect 19 92 20 93
rect 18 92 19 93
rect 17 92 18 93
rect 16 92 17 93
rect 15 92 16 93
rect 14 92 15 93
rect 13 92 14 93
rect 12 92 13 93
rect 11 92 12 93
rect 10 92 11 93
rect 9 92 10 93
rect 8 92 9 93
rect 7 92 8 93
rect 6 92 7 93
rect 195 93 196 94
rect 191 93 192 94
rect 187 93 188 94
rect 178 93 179 94
rect 177 93 178 94
rect 162 93 163 94
rect 161 93 162 94
rect 147 93 148 94
rect 117 93 118 94
rect 116 93 117 94
rect 115 93 116 94
rect 114 93 115 94
rect 113 93 114 94
rect 112 93 113 94
rect 111 93 112 94
rect 110 93 111 94
rect 109 93 110 94
rect 108 93 109 94
rect 107 93 108 94
rect 106 93 107 94
rect 105 93 106 94
rect 104 93 105 94
rect 103 93 104 94
rect 102 93 103 94
rect 101 93 102 94
rect 100 93 101 94
rect 99 93 100 94
rect 98 93 99 94
rect 97 93 98 94
rect 96 93 97 94
rect 95 93 96 94
rect 94 93 95 94
rect 93 93 94 94
rect 92 93 93 94
rect 91 93 92 94
rect 90 93 91 94
rect 89 93 90 94
rect 88 93 89 94
rect 87 93 88 94
rect 86 93 87 94
rect 85 93 86 94
rect 84 93 85 94
rect 83 93 84 94
rect 82 93 83 94
rect 81 93 82 94
rect 80 93 81 94
rect 79 93 80 94
rect 78 93 79 94
rect 77 93 78 94
rect 76 93 77 94
rect 75 93 76 94
rect 74 93 75 94
rect 73 93 74 94
rect 72 93 73 94
rect 71 93 72 94
rect 61 93 62 94
rect 60 93 61 94
rect 59 93 60 94
rect 58 93 59 94
rect 57 93 58 94
rect 56 93 57 94
rect 55 93 56 94
rect 54 93 55 94
rect 53 93 54 94
rect 52 93 53 94
rect 51 93 52 94
rect 50 93 51 94
rect 49 93 50 94
rect 48 93 49 94
rect 47 93 48 94
rect 34 93 35 94
rect 33 93 34 94
rect 32 93 33 94
rect 31 93 32 94
rect 30 93 31 94
rect 29 93 30 94
rect 28 93 29 94
rect 27 93 28 94
rect 26 93 27 94
rect 25 93 26 94
rect 24 93 25 94
rect 23 93 24 94
rect 22 93 23 94
rect 21 93 22 94
rect 20 93 21 94
rect 19 93 20 94
rect 18 93 19 94
rect 17 93 18 94
rect 16 93 17 94
rect 15 93 16 94
rect 14 93 15 94
rect 13 93 14 94
rect 12 93 13 94
rect 11 93 12 94
rect 10 93 11 94
rect 9 93 10 94
rect 8 93 9 94
rect 7 93 8 94
rect 6 93 7 94
rect 193 94 194 95
rect 192 94 193 95
rect 191 94 192 95
rect 190 94 191 95
rect 187 94 188 95
rect 179 94 180 95
rect 178 94 179 95
rect 177 94 178 95
rect 162 94 163 95
rect 161 94 162 95
rect 115 94 116 95
rect 114 94 115 95
rect 113 94 114 95
rect 112 94 113 95
rect 111 94 112 95
rect 110 94 111 95
rect 109 94 110 95
rect 108 94 109 95
rect 107 94 108 95
rect 106 94 107 95
rect 105 94 106 95
rect 104 94 105 95
rect 103 94 104 95
rect 102 94 103 95
rect 101 94 102 95
rect 100 94 101 95
rect 99 94 100 95
rect 98 94 99 95
rect 97 94 98 95
rect 96 94 97 95
rect 95 94 96 95
rect 94 94 95 95
rect 93 94 94 95
rect 92 94 93 95
rect 91 94 92 95
rect 90 94 91 95
rect 89 94 90 95
rect 88 94 89 95
rect 87 94 88 95
rect 86 94 87 95
rect 85 94 86 95
rect 84 94 85 95
rect 83 94 84 95
rect 82 94 83 95
rect 81 94 82 95
rect 80 94 81 95
rect 79 94 80 95
rect 78 94 79 95
rect 77 94 78 95
rect 76 94 77 95
rect 75 94 76 95
rect 74 94 75 95
rect 73 94 74 95
rect 72 94 73 95
rect 71 94 72 95
rect 70 94 71 95
rect 69 94 70 95
rect 61 94 62 95
rect 60 94 61 95
rect 59 94 60 95
rect 58 94 59 95
rect 57 94 58 95
rect 56 94 57 95
rect 55 94 56 95
rect 54 94 55 95
rect 53 94 54 95
rect 52 94 53 95
rect 51 94 52 95
rect 50 94 51 95
rect 49 94 50 95
rect 48 94 49 95
rect 35 94 36 95
rect 34 94 35 95
rect 33 94 34 95
rect 32 94 33 95
rect 31 94 32 95
rect 30 94 31 95
rect 29 94 30 95
rect 28 94 29 95
rect 27 94 28 95
rect 26 94 27 95
rect 25 94 26 95
rect 24 94 25 95
rect 23 94 24 95
rect 22 94 23 95
rect 21 94 22 95
rect 20 94 21 95
rect 19 94 20 95
rect 18 94 19 95
rect 17 94 18 95
rect 16 94 17 95
rect 15 94 16 95
rect 14 94 15 95
rect 13 94 14 95
rect 12 94 13 95
rect 11 94 12 95
rect 10 94 11 95
rect 9 94 10 95
rect 8 94 9 95
rect 7 94 8 95
rect 6 94 7 95
rect 5 94 6 95
rect 194 95 195 96
rect 193 95 194 96
rect 192 95 193 96
rect 191 95 192 96
rect 190 95 191 96
rect 189 95 190 96
rect 188 95 189 96
rect 187 95 188 96
rect 179 95 180 96
rect 178 95 179 96
rect 161 95 162 96
rect 160 95 161 96
rect 114 95 115 96
rect 113 95 114 96
rect 112 95 113 96
rect 111 95 112 96
rect 110 95 111 96
rect 109 95 110 96
rect 108 95 109 96
rect 107 95 108 96
rect 106 95 107 96
rect 105 95 106 96
rect 104 95 105 96
rect 103 95 104 96
rect 102 95 103 96
rect 101 95 102 96
rect 100 95 101 96
rect 99 95 100 96
rect 98 95 99 96
rect 97 95 98 96
rect 96 95 97 96
rect 95 95 96 96
rect 94 95 95 96
rect 93 95 94 96
rect 92 95 93 96
rect 91 95 92 96
rect 90 95 91 96
rect 89 95 90 96
rect 88 95 89 96
rect 87 95 88 96
rect 86 95 87 96
rect 85 95 86 96
rect 84 95 85 96
rect 83 95 84 96
rect 82 95 83 96
rect 81 95 82 96
rect 80 95 81 96
rect 79 95 80 96
rect 78 95 79 96
rect 77 95 78 96
rect 76 95 77 96
rect 75 95 76 96
rect 74 95 75 96
rect 73 95 74 96
rect 72 95 73 96
rect 71 95 72 96
rect 70 95 71 96
rect 69 95 70 96
rect 68 95 69 96
rect 61 95 62 96
rect 60 95 61 96
rect 59 95 60 96
rect 58 95 59 96
rect 57 95 58 96
rect 56 95 57 96
rect 55 95 56 96
rect 54 95 55 96
rect 53 95 54 96
rect 52 95 53 96
rect 51 95 52 96
rect 50 95 51 96
rect 49 95 50 96
rect 48 95 49 96
rect 37 95 38 96
rect 36 95 37 96
rect 35 95 36 96
rect 34 95 35 96
rect 33 95 34 96
rect 32 95 33 96
rect 31 95 32 96
rect 30 95 31 96
rect 29 95 30 96
rect 28 95 29 96
rect 27 95 28 96
rect 26 95 27 96
rect 25 95 26 96
rect 24 95 25 96
rect 23 95 24 96
rect 22 95 23 96
rect 21 95 22 96
rect 20 95 21 96
rect 19 95 20 96
rect 18 95 19 96
rect 17 95 18 96
rect 16 95 17 96
rect 15 95 16 96
rect 14 95 15 96
rect 13 95 14 96
rect 12 95 13 96
rect 11 95 12 96
rect 10 95 11 96
rect 9 95 10 96
rect 8 95 9 96
rect 7 95 8 96
rect 6 95 7 96
rect 5 95 6 96
rect 195 96 196 97
rect 194 96 195 97
rect 193 96 194 97
rect 190 96 191 97
rect 189 96 190 97
rect 188 96 189 97
rect 187 96 188 97
rect 179 96 180 97
rect 178 96 179 97
rect 170 96 171 97
rect 161 96 162 97
rect 160 96 161 97
rect 113 96 114 97
rect 112 96 113 97
rect 111 96 112 97
rect 110 96 111 97
rect 109 96 110 97
rect 108 96 109 97
rect 107 96 108 97
rect 106 96 107 97
rect 105 96 106 97
rect 104 96 105 97
rect 103 96 104 97
rect 102 96 103 97
rect 101 96 102 97
rect 100 96 101 97
rect 99 96 100 97
rect 98 96 99 97
rect 97 96 98 97
rect 96 96 97 97
rect 95 96 96 97
rect 94 96 95 97
rect 93 96 94 97
rect 92 96 93 97
rect 91 96 92 97
rect 90 96 91 97
rect 89 96 90 97
rect 88 96 89 97
rect 87 96 88 97
rect 86 96 87 97
rect 85 96 86 97
rect 84 96 85 97
rect 83 96 84 97
rect 82 96 83 97
rect 81 96 82 97
rect 80 96 81 97
rect 79 96 80 97
rect 78 96 79 97
rect 77 96 78 97
rect 76 96 77 97
rect 75 96 76 97
rect 74 96 75 97
rect 73 96 74 97
rect 72 96 73 97
rect 71 96 72 97
rect 70 96 71 97
rect 69 96 70 97
rect 61 96 62 97
rect 60 96 61 97
rect 59 96 60 97
rect 58 96 59 97
rect 57 96 58 97
rect 56 96 57 97
rect 55 96 56 97
rect 54 96 55 97
rect 53 96 54 97
rect 52 96 53 97
rect 51 96 52 97
rect 50 96 51 97
rect 49 96 50 97
rect 39 96 40 97
rect 38 96 39 97
rect 37 96 38 97
rect 36 96 37 97
rect 35 96 36 97
rect 34 96 35 97
rect 33 96 34 97
rect 32 96 33 97
rect 31 96 32 97
rect 30 96 31 97
rect 29 96 30 97
rect 28 96 29 97
rect 27 96 28 97
rect 26 96 27 97
rect 25 96 26 97
rect 24 96 25 97
rect 23 96 24 97
rect 22 96 23 97
rect 21 96 22 97
rect 20 96 21 97
rect 19 96 20 97
rect 18 96 19 97
rect 17 96 18 97
rect 16 96 17 97
rect 15 96 16 97
rect 14 96 15 97
rect 13 96 14 97
rect 12 96 13 97
rect 11 96 12 97
rect 10 96 11 97
rect 9 96 10 97
rect 8 96 9 97
rect 7 96 8 97
rect 6 96 7 97
rect 5 96 6 97
rect 195 97 196 98
rect 194 97 195 98
rect 179 97 180 98
rect 178 97 179 98
rect 171 97 172 98
rect 170 97 171 98
rect 161 97 162 98
rect 160 97 161 98
rect 112 97 113 98
rect 111 97 112 98
rect 110 97 111 98
rect 109 97 110 98
rect 108 97 109 98
rect 107 97 108 98
rect 106 97 107 98
rect 105 97 106 98
rect 104 97 105 98
rect 103 97 104 98
rect 102 97 103 98
rect 101 97 102 98
rect 100 97 101 98
rect 99 97 100 98
rect 98 97 99 98
rect 97 97 98 98
rect 96 97 97 98
rect 95 97 96 98
rect 94 97 95 98
rect 93 97 94 98
rect 92 97 93 98
rect 91 97 92 98
rect 90 97 91 98
rect 89 97 90 98
rect 88 97 89 98
rect 87 97 88 98
rect 86 97 87 98
rect 85 97 86 98
rect 84 97 85 98
rect 83 97 84 98
rect 82 97 83 98
rect 81 97 82 98
rect 80 97 81 98
rect 79 97 80 98
rect 78 97 79 98
rect 77 97 78 98
rect 76 97 77 98
rect 75 97 76 98
rect 74 97 75 98
rect 73 97 74 98
rect 72 97 73 98
rect 71 97 72 98
rect 70 97 71 98
rect 61 97 62 98
rect 60 97 61 98
rect 59 97 60 98
rect 58 97 59 98
rect 57 97 58 98
rect 56 97 57 98
rect 55 97 56 98
rect 54 97 55 98
rect 53 97 54 98
rect 52 97 53 98
rect 51 97 52 98
rect 50 97 51 98
rect 41 97 42 98
rect 40 97 41 98
rect 39 97 40 98
rect 38 97 39 98
rect 37 97 38 98
rect 36 97 37 98
rect 35 97 36 98
rect 34 97 35 98
rect 33 97 34 98
rect 32 97 33 98
rect 31 97 32 98
rect 30 97 31 98
rect 29 97 30 98
rect 28 97 29 98
rect 27 97 28 98
rect 26 97 27 98
rect 25 97 26 98
rect 24 97 25 98
rect 23 97 24 98
rect 22 97 23 98
rect 21 97 22 98
rect 20 97 21 98
rect 19 97 20 98
rect 18 97 19 98
rect 17 97 18 98
rect 16 97 17 98
rect 15 97 16 98
rect 14 97 15 98
rect 12 97 13 98
rect 11 97 12 98
rect 10 97 11 98
rect 9 97 10 98
rect 8 97 9 98
rect 7 97 8 98
rect 6 97 7 98
rect 5 97 6 98
rect 179 98 180 99
rect 178 98 179 99
rect 171 98 172 99
rect 170 98 171 99
rect 161 98 162 99
rect 160 98 161 99
rect 111 98 112 99
rect 110 98 111 99
rect 109 98 110 99
rect 108 98 109 99
rect 107 98 108 99
rect 106 98 107 99
rect 105 98 106 99
rect 104 98 105 99
rect 103 98 104 99
rect 102 98 103 99
rect 101 98 102 99
rect 100 98 101 99
rect 99 98 100 99
rect 98 98 99 99
rect 97 98 98 99
rect 96 98 97 99
rect 95 98 96 99
rect 94 98 95 99
rect 93 98 94 99
rect 92 98 93 99
rect 91 98 92 99
rect 90 98 91 99
rect 89 98 90 99
rect 88 98 89 99
rect 87 98 88 99
rect 86 98 87 99
rect 85 98 86 99
rect 84 98 85 99
rect 83 98 84 99
rect 82 98 83 99
rect 81 98 82 99
rect 80 98 81 99
rect 79 98 80 99
rect 78 98 79 99
rect 77 98 78 99
rect 76 98 77 99
rect 75 98 76 99
rect 74 98 75 99
rect 73 98 74 99
rect 72 98 73 99
rect 62 98 63 99
rect 61 98 62 99
rect 60 98 61 99
rect 59 98 60 99
rect 58 98 59 99
rect 57 98 58 99
rect 56 98 57 99
rect 55 98 56 99
rect 54 98 55 99
rect 53 98 54 99
rect 52 98 53 99
rect 51 98 52 99
rect 50 98 51 99
rect 42 98 43 99
rect 41 98 42 99
rect 40 98 41 99
rect 39 98 40 99
rect 38 98 39 99
rect 37 98 38 99
rect 36 98 37 99
rect 35 98 36 99
rect 34 98 35 99
rect 33 98 34 99
rect 32 98 33 99
rect 31 98 32 99
rect 30 98 31 99
rect 29 98 30 99
rect 28 98 29 99
rect 27 98 28 99
rect 26 98 27 99
rect 25 98 26 99
rect 24 98 25 99
rect 23 98 24 99
rect 22 98 23 99
rect 21 98 22 99
rect 20 98 21 99
rect 19 98 20 99
rect 18 98 19 99
rect 17 98 18 99
rect 16 98 17 99
rect 15 98 16 99
rect 14 98 15 99
rect 11 98 12 99
rect 10 98 11 99
rect 9 98 10 99
rect 8 98 9 99
rect 7 98 8 99
rect 6 98 7 99
rect 5 98 6 99
rect 179 99 180 100
rect 178 99 179 100
rect 177 99 178 100
rect 176 99 177 100
rect 175 99 176 100
rect 174 99 175 100
rect 173 99 174 100
rect 172 99 173 100
rect 171 99 172 100
rect 170 99 171 100
rect 162 99 163 100
rect 161 99 162 100
rect 160 99 161 100
rect 129 99 130 100
rect 128 99 129 100
rect 127 99 128 100
rect 126 99 127 100
rect 125 99 126 100
rect 124 99 125 100
rect 123 99 124 100
rect 122 99 123 100
rect 121 99 122 100
rect 120 99 121 100
rect 119 99 120 100
rect 118 99 119 100
rect 117 99 118 100
rect 110 99 111 100
rect 109 99 110 100
rect 108 99 109 100
rect 107 99 108 100
rect 106 99 107 100
rect 105 99 106 100
rect 104 99 105 100
rect 103 99 104 100
rect 102 99 103 100
rect 101 99 102 100
rect 100 99 101 100
rect 99 99 100 100
rect 98 99 99 100
rect 97 99 98 100
rect 96 99 97 100
rect 95 99 96 100
rect 94 99 95 100
rect 93 99 94 100
rect 92 99 93 100
rect 91 99 92 100
rect 90 99 91 100
rect 89 99 90 100
rect 88 99 89 100
rect 87 99 88 100
rect 86 99 87 100
rect 85 99 86 100
rect 84 99 85 100
rect 83 99 84 100
rect 82 99 83 100
rect 81 99 82 100
rect 80 99 81 100
rect 79 99 80 100
rect 78 99 79 100
rect 77 99 78 100
rect 76 99 77 100
rect 75 99 76 100
rect 74 99 75 100
rect 62 99 63 100
rect 61 99 62 100
rect 60 99 61 100
rect 59 99 60 100
rect 58 99 59 100
rect 57 99 58 100
rect 56 99 57 100
rect 55 99 56 100
rect 54 99 55 100
rect 53 99 54 100
rect 52 99 53 100
rect 51 99 52 100
rect 50 99 51 100
rect 43 99 44 100
rect 42 99 43 100
rect 41 99 42 100
rect 40 99 41 100
rect 39 99 40 100
rect 38 99 39 100
rect 37 99 38 100
rect 36 99 37 100
rect 35 99 36 100
rect 34 99 35 100
rect 33 99 34 100
rect 32 99 33 100
rect 31 99 32 100
rect 30 99 31 100
rect 29 99 30 100
rect 28 99 29 100
rect 27 99 28 100
rect 26 99 27 100
rect 25 99 26 100
rect 24 99 25 100
rect 23 99 24 100
rect 22 99 23 100
rect 21 99 22 100
rect 20 99 21 100
rect 19 99 20 100
rect 18 99 19 100
rect 17 99 18 100
rect 16 99 17 100
rect 15 99 16 100
rect 14 99 15 100
rect 11 99 12 100
rect 10 99 11 100
rect 9 99 10 100
rect 8 99 9 100
rect 7 99 8 100
rect 6 99 7 100
rect 5 99 6 100
rect 178 100 179 101
rect 177 100 178 101
rect 176 100 177 101
rect 175 100 176 101
rect 174 100 175 101
rect 173 100 174 101
rect 172 100 173 101
rect 171 100 172 101
rect 170 100 171 101
rect 163 100 164 101
rect 162 100 163 101
rect 161 100 162 101
rect 133 100 134 101
rect 132 100 133 101
rect 131 100 132 101
rect 130 100 131 101
rect 129 100 130 101
rect 128 100 129 101
rect 127 100 128 101
rect 126 100 127 101
rect 125 100 126 101
rect 124 100 125 101
rect 123 100 124 101
rect 122 100 123 101
rect 121 100 122 101
rect 120 100 121 101
rect 119 100 120 101
rect 118 100 119 101
rect 117 100 118 101
rect 116 100 117 101
rect 115 100 116 101
rect 114 100 115 101
rect 113 100 114 101
rect 110 100 111 101
rect 109 100 110 101
rect 108 100 109 101
rect 107 100 108 101
rect 106 100 107 101
rect 105 100 106 101
rect 104 100 105 101
rect 103 100 104 101
rect 102 100 103 101
rect 101 100 102 101
rect 100 100 101 101
rect 99 100 100 101
rect 98 100 99 101
rect 97 100 98 101
rect 96 100 97 101
rect 95 100 96 101
rect 94 100 95 101
rect 93 100 94 101
rect 92 100 93 101
rect 91 100 92 101
rect 90 100 91 101
rect 89 100 90 101
rect 88 100 89 101
rect 87 100 88 101
rect 86 100 87 101
rect 85 100 86 101
rect 84 100 85 101
rect 83 100 84 101
rect 82 100 83 101
rect 81 100 82 101
rect 80 100 81 101
rect 79 100 80 101
rect 78 100 79 101
rect 77 100 78 101
rect 76 100 77 101
rect 63 100 64 101
rect 62 100 63 101
rect 61 100 62 101
rect 60 100 61 101
rect 59 100 60 101
rect 58 100 59 101
rect 57 100 58 101
rect 56 100 57 101
rect 55 100 56 101
rect 54 100 55 101
rect 53 100 54 101
rect 52 100 53 101
rect 51 100 52 101
rect 44 100 45 101
rect 43 100 44 101
rect 42 100 43 101
rect 41 100 42 101
rect 40 100 41 101
rect 39 100 40 101
rect 38 100 39 101
rect 37 100 38 101
rect 36 100 37 101
rect 35 100 36 101
rect 34 100 35 101
rect 33 100 34 101
rect 32 100 33 101
rect 31 100 32 101
rect 30 100 31 101
rect 29 100 30 101
rect 28 100 29 101
rect 27 100 28 101
rect 26 100 27 101
rect 25 100 26 101
rect 24 100 25 101
rect 23 100 24 101
rect 22 100 23 101
rect 21 100 22 101
rect 20 100 21 101
rect 19 100 20 101
rect 18 100 19 101
rect 17 100 18 101
rect 16 100 17 101
rect 15 100 16 101
rect 11 100 12 101
rect 10 100 11 101
rect 9 100 10 101
rect 8 100 9 101
rect 7 100 8 101
rect 6 100 7 101
rect 5 100 6 101
rect 4 100 5 101
rect 194 101 195 102
rect 193 101 194 102
rect 189 101 190 102
rect 188 101 189 102
rect 178 101 179 102
rect 177 101 178 102
rect 176 101 177 102
rect 175 101 176 102
rect 174 101 175 102
rect 173 101 174 102
rect 172 101 173 102
rect 171 101 172 102
rect 170 101 171 102
rect 164 101 165 102
rect 163 101 164 102
rect 162 101 163 102
rect 161 101 162 102
rect 133 101 134 102
rect 132 101 133 102
rect 131 101 132 102
rect 130 101 131 102
rect 129 101 130 102
rect 128 101 129 102
rect 127 101 128 102
rect 126 101 127 102
rect 125 101 126 102
rect 124 101 125 102
rect 123 101 124 102
rect 122 101 123 102
rect 121 101 122 102
rect 120 101 121 102
rect 119 101 120 102
rect 118 101 119 102
rect 117 101 118 102
rect 116 101 117 102
rect 115 101 116 102
rect 114 101 115 102
rect 113 101 114 102
rect 112 101 113 102
rect 111 101 112 102
rect 109 101 110 102
rect 108 101 109 102
rect 107 101 108 102
rect 106 101 107 102
rect 105 101 106 102
rect 104 101 105 102
rect 103 101 104 102
rect 102 101 103 102
rect 101 101 102 102
rect 100 101 101 102
rect 99 101 100 102
rect 98 101 99 102
rect 97 101 98 102
rect 96 101 97 102
rect 91 101 92 102
rect 90 101 91 102
rect 89 101 90 102
rect 88 101 89 102
rect 87 101 88 102
rect 86 101 87 102
rect 85 101 86 102
rect 84 101 85 102
rect 83 101 84 102
rect 82 101 83 102
rect 81 101 82 102
rect 80 101 81 102
rect 79 101 80 102
rect 64 101 65 102
rect 63 101 64 102
rect 62 101 63 102
rect 61 101 62 102
rect 60 101 61 102
rect 59 101 60 102
rect 58 101 59 102
rect 57 101 58 102
rect 56 101 57 102
rect 55 101 56 102
rect 54 101 55 102
rect 53 101 54 102
rect 52 101 53 102
rect 51 101 52 102
rect 45 101 46 102
rect 44 101 45 102
rect 43 101 44 102
rect 42 101 43 102
rect 41 101 42 102
rect 40 101 41 102
rect 39 101 40 102
rect 38 101 39 102
rect 37 101 38 102
rect 36 101 37 102
rect 35 101 36 102
rect 34 101 35 102
rect 33 101 34 102
rect 32 101 33 102
rect 31 101 32 102
rect 30 101 31 102
rect 29 101 30 102
rect 28 101 29 102
rect 27 101 28 102
rect 26 101 27 102
rect 25 101 26 102
rect 24 101 25 102
rect 23 101 24 102
rect 22 101 23 102
rect 21 101 22 102
rect 20 101 21 102
rect 19 101 20 102
rect 18 101 19 102
rect 17 101 18 102
rect 16 101 17 102
rect 15 101 16 102
rect 11 101 12 102
rect 10 101 11 102
rect 9 101 10 102
rect 8 101 9 102
rect 7 101 8 102
rect 6 101 7 102
rect 5 101 6 102
rect 195 102 196 103
rect 194 102 195 103
rect 190 102 191 103
rect 189 102 190 103
rect 188 102 189 103
rect 187 102 188 103
rect 178 102 179 103
rect 177 102 178 103
rect 176 102 177 103
rect 175 102 176 103
rect 174 102 175 103
rect 173 102 174 103
rect 172 102 173 103
rect 171 102 172 103
rect 170 102 171 103
rect 165 102 166 103
rect 164 102 165 103
rect 163 102 164 103
rect 162 102 163 103
rect 161 102 162 103
rect 131 102 132 103
rect 130 102 131 103
rect 129 102 130 103
rect 128 102 129 103
rect 127 102 128 103
rect 126 102 127 103
rect 125 102 126 103
rect 124 102 125 103
rect 123 102 124 103
rect 122 102 123 103
rect 121 102 122 103
rect 120 102 121 103
rect 119 102 120 103
rect 118 102 119 103
rect 117 102 118 103
rect 116 102 117 103
rect 115 102 116 103
rect 114 102 115 103
rect 113 102 114 103
rect 112 102 113 103
rect 111 102 112 103
rect 110 102 111 103
rect 109 102 110 103
rect 108 102 109 103
rect 107 102 108 103
rect 106 102 107 103
rect 105 102 106 103
rect 104 102 105 103
rect 103 102 104 103
rect 102 102 103 103
rect 101 102 102 103
rect 100 102 101 103
rect 99 102 100 103
rect 98 102 99 103
rect 97 102 98 103
rect 96 102 97 103
rect 65 102 66 103
rect 64 102 65 103
rect 63 102 64 103
rect 62 102 63 103
rect 61 102 62 103
rect 60 102 61 103
rect 59 102 60 103
rect 58 102 59 103
rect 57 102 58 103
rect 56 102 57 103
rect 55 102 56 103
rect 54 102 55 103
rect 53 102 54 103
rect 52 102 53 103
rect 51 102 52 103
rect 45 102 46 103
rect 44 102 45 103
rect 43 102 44 103
rect 42 102 43 103
rect 41 102 42 103
rect 40 102 41 103
rect 39 102 40 103
rect 38 102 39 103
rect 37 102 38 103
rect 36 102 37 103
rect 35 102 36 103
rect 34 102 35 103
rect 33 102 34 103
rect 32 102 33 103
rect 31 102 32 103
rect 30 102 31 103
rect 29 102 30 103
rect 28 102 29 103
rect 27 102 28 103
rect 26 102 27 103
rect 25 102 26 103
rect 24 102 25 103
rect 23 102 24 103
rect 22 102 23 103
rect 21 102 22 103
rect 20 102 21 103
rect 19 102 20 103
rect 18 102 19 103
rect 17 102 18 103
rect 16 102 17 103
rect 15 102 16 103
rect 11 102 12 103
rect 10 102 11 103
rect 9 102 10 103
rect 8 102 9 103
rect 7 102 8 103
rect 6 102 7 103
rect 5 102 6 103
rect 4 102 5 103
rect 195 103 196 104
rect 191 103 192 104
rect 190 103 191 104
rect 189 103 190 104
rect 187 103 188 104
rect 186 103 187 104
rect 171 103 172 104
rect 170 103 171 104
rect 130 103 131 104
rect 129 103 130 104
rect 128 103 129 104
rect 127 103 128 104
rect 126 103 127 104
rect 125 103 126 104
rect 124 103 125 104
rect 123 103 124 104
rect 122 103 123 104
rect 121 103 122 104
rect 120 103 121 104
rect 119 103 120 104
rect 118 103 119 104
rect 117 103 118 104
rect 116 103 117 104
rect 115 103 116 104
rect 114 103 115 104
rect 113 103 114 104
rect 112 103 113 104
rect 111 103 112 104
rect 110 103 111 104
rect 109 103 110 104
rect 108 103 109 104
rect 107 103 108 104
rect 106 103 107 104
rect 105 103 106 104
rect 104 103 105 104
rect 103 103 104 104
rect 102 103 103 104
rect 101 103 102 104
rect 100 103 101 104
rect 99 103 100 104
rect 98 103 99 104
rect 97 103 98 104
rect 96 103 97 104
rect 95 103 96 104
rect 66 103 67 104
rect 65 103 66 104
rect 64 103 65 104
rect 63 103 64 104
rect 62 103 63 104
rect 61 103 62 104
rect 60 103 61 104
rect 59 103 60 104
rect 58 103 59 104
rect 57 103 58 104
rect 56 103 57 104
rect 55 103 56 104
rect 54 103 55 104
rect 53 103 54 104
rect 52 103 53 104
rect 51 103 52 104
rect 46 103 47 104
rect 45 103 46 104
rect 44 103 45 104
rect 43 103 44 104
rect 42 103 43 104
rect 41 103 42 104
rect 40 103 41 104
rect 39 103 40 104
rect 38 103 39 104
rect 37 103 38 104
rect 36 103 37 104
rect 35 103 36 104
rect 34 103 35 104
rect 33 103 34 104
rect 32 103 33 104
rect 31 103 32 104
rect 30 103 31 104
rect 29 103 30 104
rect 28 103 29 104
rect 27 103 28 104
rect 26 103 27 104
rect 25 103 26 104
rect 24 103 25 104
rect 23 103 24 104
rect 22 103 23 104
rect 21 103 22 104
rect 20 103 21 104
rect 19 103 20 104
rect 18 103 19 104
rect 17 103 18 104
rect 16 103 17 104
rect 11 103 12 104
rect 10 103 11 104
rect 9 103 10 104
rect 8 103 9 104
rect 7 103 8 104
rect 6 103 7 104
rect 5 103 6 104
rect 4 103 5 104
rect 195 104 196 105
rect 192 104 193 105
rect 191 104 192 105
rect 190 104 191 105
rect 187 104 188 105
rect 186 104 187 105
rect 171 104 172 105
rect 170 104 171 105
rect 128 104 129 105
rect 127 104 128 105
rect 126 104 127 105
rect 125 104 126 105
rect 124 104 125 105
rect 123 104 124 105
rect 122 104 123 105
rect 121 104 122 105
rect 120 104 121 105
rect 119 104 120 105
rect 118 104 119 105
rect 117 104 118 105
rect 116 104 117 105
rect 115 104 116 105
rect 114 104 115 105
rect 113 104 114 105
rect 112 104 113 105
rect 111 104 112 105
rect 110 104 111 105
rect 109 104 110 105
rect 108 104 109 105
rect 107 104 108 105
rect 106 104 107 105
rect 105 104 106 105
rect 104 104 105 105
rect 103 104 104 105
rect 102 104 103 105
rect 101 104 102 105
rect 100 104 101 105
rect 99 104 100 105
rect 98 104 99 105
rect 97 104 98 105
rect 96 104 97 105
rect 95 104 96 105
rect 67 104 68 105
rect 66 104 67 105
rect 65 104 66 105
rect 64 104 65 105
rect 63 104 64 105
rect 62 104 63 105
rect 61 104 62 105
rect 60 104 61 105
rect 59 104 60 105
rect 58 104 59 105
rect 57 104 58 105
rect 56 104 57 105
rect 55 104 56 105
rect 54 104 55 105
rect 53 104 54 105
rect 52 104 53 105
rect 46 104 47 105
rect 45 104 46 105
rect 44 104 45 105
rect 43 104 44 105
rect 42 104 43 105
rect 41 104 42 105
rect 40 104 41 105
rect 39 104 40 105
rect 38 104 39 105
rect 37 104 38 105
rect 36 104 37 105
rect 35 104 36 105
rect 34 104 35 105
rect 33 104 34 105
rect 32 104 33 105
rect 31 104 32 105
rect 30 104 31 105
rect 29 104 30 105
rect 28 104 29 105
rect 27 104 28 105
rect 26 104 27 105
rect 25 104 26 105
rect 24 104 25 105
rect 23 104 24 105
rect 22 104 23 105
rect 21 104 22 105
rect 20 104 21 105
rect 19 104 20 105
rect 18 104 19 105
rect 17 104 18 105
rect 16 104 17 105
rect 11 104 12 105
rect 10 104 11 105
rect 9 104 10 105
rect 8 104 9 105
rect 7 104 8 105
rect 6 104 7 105
rect 5 104 6 105
rect 4 104 5 105
rect 194 105 195 106
rect 193 105 194 106
rect 192 105 193 106
rect 191 105 192 106
rect 190 105 191 106
rect 187 105 188 106
rect 186 105 187 106
rect 127 105 128 106
rect 126 105 127 106
rect 125 105 126 106
rect 124 105 125 106
rect 123 105 124 106
rect 122 105 123 106
rect 121 105 122 106
rect 120 105 121 106
rect 119 105 120 106
rect 118 105 119 106
rect 117 105 118 106
rect 116 105 117 106
rect 115 105 116 106
rect 114 105 115 106
rect 113 105 114 106
rect 112 105 113 106
rect 111 105 112 106
rect 110 105 111 106
rect 109 105 110 106
rect 108 105 109 106
rect 107 105 108 106
rect 106 105 107 106
rect 105 105 106 106
rect 104 105 105 106
rect 103 105 104 106
rect 102 105 103 106
rect 101 105 102 106
rect 100 105 101 106
rect 99 105 100 106
rect 98 105 99 106
rect 97 105 98 106
rect 96 105 97 106
rect 95 105 96 106
rect 69 105 70 106
rect 68 105 69 106
rect 67 105 68 106
rect 66 105 67 106
rect 65 105 66 106
rect 64 105 65 106
rect 63 105 64 106
rect 62 105 63 106
rect 61 105 62 106
rect 60 105 61 106
rect 59 105 60 106
rect 58 105 59 106
rect 57 105 58 106
rect 56 105 57 106
rect 55 105 56 106
rect 54 105 55 106
rect 53 105 54 106
rect 52 105 53 106
rect 46 105 47 106
rect 45 105 46 106
rect 44 105 45 106
rect 43 105 44 106
rect 42 105 43 106
rect 41 105 42 106
rect 40 105 41 106
rect 39 105 40 106
rect 38 105 39 106
rect 37 105 38 106
rect 36 105 37 106
rect 35 105 36 106
rect 34 105 35 106
rect 33 105 34 106
rect 32 105 33 106
rect 31 105 32 106
rect 30 105 31 106
rect 29 105 30 106
rect 28 105 29 106
rect 27 105 28 106
rect 25 105 26 106
rect 24 105 25 106
rect 23 105 24 106
rect 22 105 23 106
rect 21 105 22 106
rect 20 105 21 106
rect 19 105 20 106
rect 18 105 19 106
rect 17 105 18 106
rect 16 105 17 106
rect 12 105 13 106
rect 11 105 12 106
rect 10 105 11 106
rect 9 105 10 106
rect 8 105 9 106
rect 7 105 8 106
rect 6 105 7 106
rect 5 105 6 106
rect 4 105 5 106
rect 193 106 194 107
rect 192 106 193 107
rect 191 106 192 107
rect 188 106 189 107
rect 187 106 188 107
rect 126 106 127 107
rect 125 106 126 107
rect 124 106 125 107
rect 123 106 124 107
rect 122 106 123 107
rect 121 106 122 107
rect 120 106 121 107
rect 119 106 120 107
rect 118 106 119 107
rect 117 106 118 107
rect 116 106 117 107
rect 115 106 116 107
rect 114 106 115 107
rect 113 106 114 107
rect 112 106 113 107
rect 111 106 112 107
rect 110 106 111 107
rect 109 106 110 107
rect 108 106 109 107
rect 107 106 108 107
rect 106 106 107 107
rect 105 106 106 107
rect 104 106 105 107
rect 103 106 104 107
rect 102 106 103 107
rect 101 106 102 107
rect 100 106 101 107
rect 99 106 100 107
rect 98 106 99 107
rect 97 106 98 107
rect 96 106 97 107
rect 95 106 96 107
rect 71 106 72 107
rect 70 106 71 107
rect 69 106 70 107
rect 68 106 69 107
rect 67 106 68 107
rect 66 106 67 107
rect 65 106 66 107
rect 64 106 65 107
rect 63 106 64 107
rect 62 106 63 107
rect 61 106 62 107
rect 60 106 61 107
rect 59 106 60 107
rect 58 106 59 107
rect 57 106 58 107
rect 56 106 57 107
rect 55 106 56 107
rect 54 106 55 107
rect 53 106 54 107
rect 52 106 53 107
rect 47 106 48 107
rect 46 106 47 107
rect 45 106 46 107
rect 44 106 45 107
rect 43 106 44 107
rect 42 106 43 107
rect 41 106 42 107
rect 40 106 41 107
rect 39 106 40 107
rect 38 106 39 107
rect 37 106 38 107
rect 36 106 37 107
rect 35 106 36 107
rect 34 106 35 107
rect 33 106 34 107
rect 32 106 33 107
rect 31 106 32 107
rect 30 106 31 107
rect 25 106 26 107
rect 24 106 25 107
rect 23 106 24 107
rect 22 106 23 107
rect 21 106 22 107
rect 20 106 21 107
rect 19 106 20 107
rect 18 106 19 107
rect 17 106 18 107
rect 12 106 13 107
rect 11 106 12 107
rect 10 106 11 107
rect 9 106 10 107
rect 8 106 9 107
rect 7 106 8 107
rect 6 106 7 107
rect 5 106 6 107
rect 4 106 5 107
rect 125 107 126 108
rect 124 107 125 108
rect 123 107 124 108
rect 122 107 123 108
rect 121 107 122 108
rect 120 107 121 108
rect 119 107 120 108
rect 118 107 119 108
rect 117 107 118 108
rect 116 107 117 108
rect 115 107 116 108
rect 114 107 115 108
rect 113 107 114 108
rect 112 107 113 108
rect 111 107 112 108
rect 110 107 111 108
rect 109 107 110 108
rect 108 107 109 108
rect 107 107 108 108
rect 106 107 107 108
rect 105 107 106 108
rect 104 107 105 108
rect 103 107 104 108
rect 102 107 103 108
rect 101 107 102 108
rect 100 107 101 108
rect 99 107 100 108
rect 98 107 99 108
rect 97 107 98 108
rect 96 107 97 108
rect 95 107 96 108
rect 94 107 95 108
rect 75 107 76 108
rect 74 107 75 108
rect 73 107 74 108
rect 72 107 73 108
rect 71 107 72 108
rect 70 107 71 108
rect 69 107 70 108
rect 68 107 69 108
rect 67 107 68 108
rect 66 107 67 108
rect 65 107 66 108
rect 64 107 65 108
rect 63 107 64 108
rect 62 107 63 108
rect 61 107 62 108
rect 60 107 61 108
rect 59 107 60 108
rect 58 107 59 108
rect 57 107 58 108
rect 56 107 57 108
rect 55 107 56 108
rect 54 107 55 108
rect 53 107 54 108
rect 52 107 53 108
rect 47 107 48 108
rect 46 107 47 108
rect 45 107 46 108
rect 44 107 45 108
rect 43 107 44 108
rect 42 107 43 108
rect 41 107 42 108
rect 40 107 41 108
rect 39 107 40 108
rect 38 107 39 108
rect 37 107 38 108
rect 36 107 37 108
rect 35 107 36 108
rect 34 107 35 108
rect 33 107 34 108
rect 32 107 33 108
rect 31 107 32 108
rect 25 107 26 108
rect 24 107 25 108
rect 23 107 24 108
rect 22 107 23 108
rect 21 107 22 108
rect 20 107 21 108
rect 19 107 20 108
rect 18 107 19 108
rect 17 107 18 108
rect 12 107 13 108
rect 11 107 12 108
rect 10 107 11 108
rect 9 107 10 108
rect 8 107 9 108
rect 7 107 8 108
rect 6 107 7 108
rect 5 107 6 108
rect 4 107 5 108
rect 124 108 125 109
rect 123 108 124 109
rect 122 108 123 109
rect 121 108 122 109
rect 120 108 121 109
rect 119 108 120 109
rect 118 108 119 109
rect 117 108 118 109
rect 116 108 117 109
rect 115 108 116 109
rect 114 108 115 109
rect 113 108 114 109
rect 112 108 113 109
rect 111 108 112 109
rect 110 108 111 109
rect 109 108 110 109
rect 108 108 109 109
rect 107 108 108 109
rect 106 108 107 109
rect 105 108 106 109
rect 104 108 105 109
rect 103 108 104 109
rect 102 108 103 109
rect 101 108 102 109
rect 100 108 101 109
rect 99 108 100 109
rect 98 108 99 109
rect 97 108 98 109
rect 96 108 97 109
rect 95 108 96 109
rect 94 108 95 109
rect 85 108 86 109
rect 84 108 85 109
rect 80 108 81 109
rect 79 108 80 109
rect 78 108 79 109
rect 77 108 78 109
rect 76 108 77 109
rect 75 108 76 109
rect 74 108 75 109
rect 73 108 74 109
rect 72 108 73 109
rect 71 108 72 109
rect 70 108 71 109
rect 69 108 70 109
rect 68 108 69 109
rect 67 108 68 109
rect 66 108 67 109
rect 65 108 66 109
rect 64 108 65 109
rect 63 108 64 109
rect 62 108 63 109
rect 61 108 62 109
rect 60 108 61 109
rect 59 108 60 109
rect 58 108 59 109
rect 57 108 58 109
rect 56 108 57 109
rect 55 108 56 109
rect 54 108 55 109
rect 53 108 54 109
rect 52 108 53 109
rect 47 108 48 109
rect 46 108 47 109
rect 45 108 46 109
rect 44 108 45 109
rect 43 108 44 109
rect 42 108 43 109
rect 41 108 42 109
rect 40 108 41 109
rect 39 108 40 109
rect 38 108 39 109
rect 37 108 38 109
rect 36 108 37 109
rect 35 108 36 109
rect 34 108 35 109
rect 33 108 34 109
rect 32 108 33 109
rect 25 108 26 109
rect 24 108 25 109
rect 23 108 24 109
rect 22 108 23 109
rect 21 108 22 109
rect 20 108 21 109
rect 19 108 20 109
rect 18 108 19 109
rect 17 108 18 109
rect 13 108 14 109
rect 12 108 13 109
rect 11 108 12 109
rect 10 108 11 109
rect 9 108 10 109
rect 8 108 9 109
rect 7 108 8 109
rect 6 108 7 109
rect 5 108 6 109
rect 4 108 5 109
rect 123 109 124 110
rect 122 109 123 110
rect 121 109 122 110
rect 120 109 121 110
rect 119 109 120 110
rect 118 109 119 110
rect 117 109 118 110
rect 116 109 117 110
rect 115 109 116 110
rect 114 109 115 110
rect 113 109 114 110
rect 112 109 113 110
rect 111 109 112 110
rect 110 109 111 110
rect 109 109 110 110
rect 108 109 109 110
rect 107 109 108 110
rect 106 109 107 110
rect 105 109 106 110
rect 104 109 105 110
rect 103 109 104 110
rect 102 109 103 110
rect 101 109 102 110
rect 100 109 101 110
rect 99 109 100 110
rect 98 109 99 110
rect 97 109 98 110
rect 96 109 97 110
rect 95 109 96 110
rect 94 109 95 110
rect 85 109 86 110
rect 84 109 85 110
rect 83 109 84 110
rect 82 109 83 110
rect 81 109 82 110
rect 80 109 81 110
rect 79 109 80 110
rect 78 109 79 110
rect 77 109 78 110
rect 76 109 77 110
rect 75 109 76 110
rect 74 109 75 110
rect 73 109 74 110
rect 72 109 73 110
rect 71 109 72 110
rect 70 109 71 110
rect 69 109 70 110
rect 68 109 69 110
rect 67 109 68 110
rect 66 109 67 110
rect 65 109 66 110
rect 64 109 65 110
rect 63 109 64 110
rect 62 109 63 110
rect 61 109 62 110
rect 60 109 61 110
rect 59 109 60 110
rect 58 109 59 110
rect 57 109 58 110
rect 56 109 57 110
rect 55 109 56 110
rect 54 109 55 110
rect 53 109 54 110
rect 47 109 48 110
rect 46 109 47 110
rect 45 109 46 110
rect 44 109 45 110
rect 43 109 44 110
rect 42 109 43 110
rect 41 109 42 110
rect 40 109 41 110
rect 39 109 40 110
rect 38 109 39 110
rect 37 109 38 110
rect 36 109 37 110
rect 35 109 36 110
rect 34 109 35 110
rect 33 109 34 110
rect 32 109 33 110
rect 26 109 27 110
rect 25 109 26 110
rect 24 109 25 110
rect 23 109 24 110
rect 22 109 23 110
rect 21 109 22 110
rect 20 109 21 110
rect 19 109 20 110
rect 18 109 19 110
rect 17 109 18 110
rect 13 109 14 110
rect 12 109 13 110
rect 11 109 12 110
rect 10 109 11 110
rect 9 109 10 110
rect 8 109 9 110
rect 7 109 8 110
rect 6 109 7 110
rect 5 109 6 110
rect 4 109 5 110
rect 187 110 188 111
rect 122 110 123 111
rect 121 110 122 111
rect 120 110 121 111
rect 119 110 120 111
rect 118 110 119 111
rect 117 110 118 111
rect 116 110 117 111
rect 115 110 116 111
rect 114 110 115 111
rect 113 110 114 111
rect 112 110 113 111
rect 111 110 112 111
rect 110 110 111 111
rect 109 110 110 111
rect 108 110 109 111
rect 107 110 108 111
rect 106 110 107 111
rect 105 110 106 111
rect 104 110 105 111
rect 103 110 104 111
rect 102 110 103 111
rect 101 110 102 111
rect 100 110 101 111
rect 99 110 100 111
rect 98 110 99 111
rect 97 110 98 111
rect 96 110 97 111
rect 95 110 96 111
rect 94 110 95 111
rect 93 110 94 111
rect 85 110 86 111
rect 84 110 85 111
rect 83 110 84 111
rect 82 110 83 111
rect 81 110 82 111
rect 80 110 81 111
rect 79 110 80 111
rect 78 110 79 111
rect 77 110 78 111
rect 76 110 77 111
rect 75 110 76 111
rect 74 110 75 111
rect 73 110 74 111
rect 72 110 73 111
rect 71 110 72 111
rect 70 110 71 111
rect 69 110 70 111
rect 68 110 69 111
rect 67 110 68 111
rect 66 110 67 111
rect 65 110 66 111
rect 64 110 65 111
rect 63 110 64 111
rect 62 110 63 111
rect 61 110 62 111
rect 60 110 61 111
rect 59 110 60 111
rect 58 110 59 111
rect 57 110 58 111
rect 56 110 57 111
rect 55 110 56 111
rect 54 110 55 111
rect 53 110 54 111
rect 47 110 48 111
rect 46 110 47 111
rect 45 110 46 111
rect 44 110 45 111
rect 43 110 44 111
rect 42 110 43 111
rect 41 110 42 111
rect 40 110 41 111
rect 39 110 40 111
rect 38 110 39 111
rect 37 110 38 111
rect 36 110 37 111
rect 35 110 36 111
rect 34 110 35 111
rect 33 110 34 111
rect 26 110 27 111
rect 25 110 26 111
rect 24 110 25 111
rect 23 110 24 111
rect 22 110 23 111
rect 21 110 22 111
rect 20 110 21 111
rect 19 110 20 111
rect 18 110 19 111
rect 13 110 14 111
rect 12 110 13 111
rect 11 110 12 111
rect 10 110 11 111
rect 9 110 10 111
rect 8 110 9 111
rect 7 110 8 111
rect 6 110 7 111
rect 5 110 6 111
rect 4 110 5 111
rect 195 111 196 112
rect 194 111 195 112
rect 193 111 194 112
rect 192 111 193 112
rect 191 111 192 112
rect 190 111 191 112
rect 189 111 190 112
rect 188 111 189 112
rect 187 111 188 112
rect 122 111 123 112
rect 121 111 122 112
rect 120 111 121 112
rect 119 111 120 112
rect 118 111 119 112
rect 117 111 118 112
rect 116 111 117 112
rect 115 111 116 112
rect 114 111 115 112
rect 113 111 114 112
rect 112 111 113 112
rect 111 111 112 112
rect 110 111 111 112
rect 109 111 110 112
rect 108 111 109 112
rect 107 111 108 112
rect 106 111 107 112
rect 105 111 106 112
rect 104 111 105 112
rect 103 111 104 112
rect 102 111 103 112
rect 101 111 102 112
rect 100 111 101 112
rect 99 111 100 112
rect 98 111 99 112
rect 97 111 98 112
rect 96 111 97 112
rect 95 111 96 112
rect 94 111 95 112
rect 93 111 94 112
rect 84 111 85 112
rect 83 111 84 112
rect 82 111 83 112
rect 81 111 82 112
rect 80 111 81 112
rect 79 111 80 112
rect 78 111 79 112
rect 77 111 78 112
rect 76 111 77 112
rect 75 111 76 112
rect 74 111 75 112
rect 73 111 74 112
rect 72 111 73 112
rect 71 111 72 112
rect 70 111 71 112
rect 69 111 70 112
rect 68 111 69 112
rect 67 111 68 112
rect 66 111 67 112
rect 65 111 66 112
rect 64 111 65 112
rect 63 111 64 112
rect 62 111 63 112
rect 61 111 62 112
rect 60 111 61 112
rect 59 111 60 112
rect 58 111 59 112
rect 57 111 58 112
rect 56 111 57 112
rect 55 111 56 112
rect 54 111 55 112
rect 53 111 54 112
rect 47 111 48 112
rect 46 111 47 112
rect 45 111 46 112
rect 44 111 45 112
rect 43 111 44 112
rect 42 111 43 112
rect 41 111 42 112
rect 40 111 41 112
rect 39 111 40 112
rect 38 111 39 112
rect 37 111 38 112
rect 36 111 37 112
rect 35 111 36 112
rect 34 111 35 112
rect 27 111 28 112
rect 26 111 27 112
rect 25 111 26 112
rect 24 111 25 112
rect 23 111 24 112
rect 22 111 23 112
rect 21 111 22 112
rect 20 111 21 112
rect 19 111 20 112
rect 18 111 19 112
rect 13 111 14 112
rect 12 111 13 112
rect 11 111 12 112
rect 10 111 11 112
rect 9 111 10 112
rect 8 111 9 112
rect 7 111 8 112
rect 6 111 7 112
rect 5 111 6 112
rect 4 111 5 112
rect 195 112 196 113
rect 194 112 195 113
rect 193 112 194 113
rect 192 112 193 113
rect 191 112 192 113
rect 190 112 191 113
rect 189 112 190 113
rect 188 112 189 113
rect 187 112 188 113
rect 121 112 122 113
rect 120 112 121 113
rect 119 112 120 113
rect 118 112 119 113
rect 117 112 118 113
rect 116 112 117 113
rect 115 112 116 113
rect 114 112 115 113
rect 113 112 114 113
rect 112 112 113 113
rect 111 112 112 113
rect 110 112 111 113
rect 109 112 110 113
rect 108 112 109 113
rect 107 112 108 113
rect 106 112 107 113
rect 105 112 106 113
rect 104 112 105 113
rect 103 112 104 113
rect 102 112 103 113
rect 101 112 102 113
rect 100 112 101 113
rect 99 112 100 113
rect 98 112 99 113
rect 97 112 98 113
rect 96 112 97 113
rect 95 112 96 113
rect 94 112 95 113
rect 93 112 94 113
rect 84 112 85 113
rect 83 112 84 113
rect 82 112 83 113
rect 81 112 82 113
rect 80 112 81 113
rect 79 112 80 113
rect 78 112 79 113
rect 77 112 78 113
rect 76 112 77 113
rect 75 112 76 113
rect 74 112 75 113
rect 73 112 74 113
rect 72 112 73 113
rect 71 112 72 113
rect 70 112 71 113
rect 69 112 70 113
rect 68 112 69 113
rect 67 112 68 113
rect 66 112 67 113
rect 65 112 66 113
rect 64 112 65 113
rect 63 112 64 113
rect 62 112 63 113
rect 61 112 62 113
rect 60 112 61 113
rect 59 112 60 113
rect 58 112 59 113
rect 57 112 58 113
rect 56 112 57 113
rect 55 112 56 113
rect 54 112 55 113
rect 48 112 49 113
rect 47 112 48 113
rect 46 112 47 113
rect 45 112 46 113
rect 44 112 45 113
rect 43 112 44 113
rect 42 112 43 113
rect 41 112 42 113
rect 40 112 41 113
rect 39 112 40 113
rect 38 112 39 113
rect 37 112 38 113
rect 36 112 37 113
rect 35 112 36 113
rect 34 112 35 113
rect 27 112 28 113
rect 26 112 27 113
rect 25 112 26 113
rect 24 112 25 113
rect 23 112 24 113
rect 22 112 23 113
rect 21 112 22 113
rect 20 112 21 113
rect 19 112 20 113
rect 18 112 19 113
rect 13 112 14 113
rect 12 112 13 113
rect 11 112 12 113
rect 10 112 11 113
rect 9 112 10 113
rect 8 112 9 113
rect 7 112 8 113
rect 6 112 7 113
rect 5 112 6 113
rect 4 112 5 113
rect 194 113 195 114
rect 187 113 188 114
rect 178 113 179 114
rect 161 113 162 114
rect 120 113 121 114
rect 119 113 120 114
rect 118 113 119 114
rect 117 113 118 114
rect 116 113 117 114
rect 115 113 116 114
rect 114 113 115 114
rect 113 113 114 114
rect 112 113 113 114
rect 111 113 112 114
rect 110 113 111 114
rect 109 113 110 114
rect 108 113 109 114
rect 107 113 108 114
rect 106 113 107 114
rect 105 113 106 114
rect 104 113 105 114
rect 103 113 104 114
rect 102 113 103 114
rect 101 113 102 114
rect 100 113 101 114
rect 99 113 100 114
rect 98 113 99 114
rect 97 113 98 114
rect 96 113 97 114
rect 95 113 96 114
rect 94 113 95 114
rect 93 113 94 114
rect 92 113 93 114
rect 83 113 84 114
rect 82 113 83 114
rect 81 113 82 114
rect 80 113 81 114
rect 79 113 80 114
rect 78 113 79 114
rect 77 113 78 114
rect 76 113 77 114
rect 75 113 76 114
rect 74 113 75 114
rect 73 113 74 114
rect 72 113 73 114
rect 71 113 72 114
rect 70 113 71 114
rect 69 113 70 114
rect 68 113 69 114
rect 67 113 68 114
rect 66 113 67 114
rect 65 113 66 114
rect 64 113 65 114
rect 63 113 64 114
rect 62 113 63 114
rect 61 113 62 114
rect 60 113 61 114
rect 59 113 60 114
rect 58 113 59 114
rect 57 113 58 114
rect 56 113 57 114
rect 55 113 56 114
rect 54 113 55 114
rect 48 113 49 114
rect 47 113 48 114
rect 46 113 47 114
rect 45 113 46 114
rect 44 113 45 114
rect 43 113 44 114
rect 42 113 43 114
rect 41 113 42 114
rect 40 113 41 114
rect 39 113 40 114
rect 38 113 39 114
rect 37 113 38 114
rect 36 113 37 114
rect 35 113 36 114
rect 28 113 29 114
rect 27 113 28 114
rect 26 113 27 114
rect 25 113 26 114
rect 24 113 25 114
rect 23 113 24 114
rect 22 113 23 114
rect 21 113 22 114
rect 20 113 21 114
rect 19 113 20 114
rect 18 113 19 114
rect 14 113 15 114
rect 13 113 14 114
rect 12 113 13 114
rect 11 113 12 114
rect 10 113 11 114
rect 9 113 10 114
rect 8 113 9 114
rect 7 113 8 114
rect 6 113 7 114
rect 5 113 6 114
rect 4 113 5 114
rect 178 114 179 115
rect 162 114 163 115
rect 161 114 162 115
rect 119 114 120 115
rect 118 114 119 115
rect 117 114 118 115
rect 116 114 117 115
rect 115 114 116 115
rect 114 114 115 115
rect 113 114 114 115
rect 112 114 113 115
rect 111 114 112 115
rect 110 114 111 115
rect 109 114 110 115
rect 108 114 109 115
rect 107 114 108 115
rect 106 114 107 115
rect 105 114 106 115
rect 104 114 105 115
rect 103 114 104 115
rect 102 114 103 115
rect 101 114 102 115
rect 100 114 101 115
rect 99 114 100 115
rect 98 114 99 115
rect 97 114 98 115
rect 96 114 97 115
rect 95 114 96 115
rect 94 114 95 115
rect 93 114 94 115
rect 92 114 93 115
rect 83 114 84 115
rect 82 114 83 115
rect 81 114 82 115
rect 80 114 81 115
rect 79 114 80 115
rect 78 114 79 115
rect 77 114 78 115
rect 76 114 77 115
rect 75 114 76 115
rect 74 114 75 115
rect 73 114 74 115
rect 72 114 73 115
rect 71 114 72 115
rect 70 114 71 115
rect 69 114 70 115
rect 68 114 69 115
rect 67 114 68 115
rect 66 114 67 115
rect 65 114 66 115
rect 64 114 65 115
rect 63 114 64 115
rect 62 114 63 115
rect 61 114 62 115
rect 60 114 61 115
rect 59 114 60 115
rect 58 114 59 115
rect 57 114 58 115
rect 56 114 57 115
rect 55 114 56 115
rect 54 114 55 115
rect 48 114 49 115
rect 47 114 48 115
rect 46 114 47 115
rect 45 114 46 115
rect 44 114 45 115
rect 43 114 44 115
rect 42 114 43 115
rect 41 114 42 115
rect 40 114 41 115
rect 39 114 40 115
rect 38 114 39 115
rect 37 114 38 115
rect 36 114 37 115
rect 35 114 36 115
rect 28 114 29 115
rect 27 114 28 115
rect 26 114 27 115
rect 25 114 26 115
rect 24 114 25 115
rect 23 114 24 115
rect 22 114 23 115
rect 21 114 22 115
rect 20 114 21 115
rect 19 114 20 115
rect 18 114 19 115
rect 14 114 15 115
rect 13 114 14 115
rect 12 114 13 115
rect 11 114 12 115
rect 10 114 11 115
rect 9 114 10 115
rect 8 114 9 115
rect 7 114 8 115
rect 6 114 7 115
rect 5 114 6 115
rect 4 114 5 115
rect 178 115 179 116
rect 177 115 178 116
rect 176 115 177 116
rect 175 115 176 116
rect 174 115 175 116
rect 173 115 174 116
rect 172 115 173 116
rect 171 115 172 116
rect 170 115 171 116
rect 169 115 170 116
rect 168 115 169 116
rect 167 115 168 116
rect 166 115 167 116
rect 165 115 166 116
rect 164 115 165 116
rect 163 115 164 116
rect 162 115 163 116
rect 161 115 162 116
rect 119 115 120 116
rect 118 115 119 116
rect 117 115 118 116
rect 116 115 117 116
rect 115 115 116 116
rect 114 115 115 116
rect 113 115 114 116
rect 112 115 113 116
rect 111 115 112 116
rect 110 115 111 116
rect 109 115 110 116
rect 108 115 109 116
rect 107 115 108 116
rect 106 115 107 116
rect 105 115 106 116
rect 104 115 105 116
rect 103 115 104 116
rect 102 115 103 116
rect 101 115 102 116
rect 100 115 101 116
rect 99 115 100 116
rect 98 115 99 116
rect 97 115 98 116
rect 96 115 97 116
rect 95 115 96 116
rect 94 115 95 116
rect 93 115 94 116
rect 92 115 93 116
rect 91 115 92 116
rect 82 115 83 116
rect 81 115 82 116
rect 80 115 81 116
rect 79 115 80 116
rect 78 115 79 116
rect 77 115 78 116
rect 76 115 77 116
rect 75 115 76 116
rect 74 115 75 116
rect 73 115 74 116
rect 72 115 73 116
rect 71 115 72 116
rect 70 115 71 116
rect 69 115 70 116
rect 68 115 69 116
rect 67 115 68 116
rect 66 115 67 116
rect 65 115 66 116
rect 64 115 65 116
rect 63 115 64 116
rect 62 115 63 116
rect 61 115 62 116
rect 60 115 61 116
rect 59 115 60 116
rect 58 115 59 116
rect 57 115 58 116
rect 56 115 57 116
rect 55 115 56 116
rect 48 115 49 116
rect 47 115 48 116
rect 46 115 47 116
rect 45 115 46 116
rect 44 115 45 116
rect 43 115 44 116
rect 42 115 43 116
rect 41 115 42 116
rect 40 115 41 116
rect 39 115 40 116
rect 38 115 39 116
rect 37 115 38 116
rect 36 115 37 116
rect 35 115 36 116
rect 28 115 29 116
rect 27 115 28 116
rect 26 115 27 116
rect 25 115 26 116
rect 24 115 25 116
rect 23 115 24 116
rect 22 115 23 116
rect 21 115 22 116
rect 20 115 21 116
rect 19 115 20 116
rect 18 115 19 116
rect 14 115 15 116
rect 13 115 14 116
rect 12 115 13 116
rect 11 115 12 116
rect 10 115 11 116
rect 9 115 10 116
rect 8 115 9 116
rect 7 115 8 116
rect 6 115 7 116
rect 5 115 6 116
rect 4 115 5 116
rect 178 116 179 117
rect 177 116 178 117
rect 176 116 177 117
rect 175 116 176 117
rect 174 116 175 117
rect 173 116 174 117
rect 172 116 173 117
rect 171 116 172 117
rect 170 116 171 117
rect 169 116 170 117
rect 168 116 169 117
rect 167 116 168 117
rect 166 116 167 117
rect 165 116 166 117
rect 164 116 165 117
rect 163 116 164 117
rect 162 116 163 117
rect 161 116 162 117
rect 118 116 119 117
rect 117 116 118 117
rect 116 116 117 117
rect 115 116 116 117
rect 114 116 115 117
rect 113 116 114 117
rect 112 116 113 117
rect 111 116 112 117
rect 110 116 111 117
rect 109 116 110 117
rect 108 116 109 117
rect 107 116 108 117
rect 106 116 107 117
rect 105 116 106 117
rect 104 116 105 117
rect 103 116 104 117
rect 102 116 103 117
rect 101 116 102 117
rect 100 116 101 117
rect 99 116 100 117
rect 98 116 99 117
rect 97 116 98 117
rect 96 116 97 117
rect 95 116 96 117
rect 94 116 95 117
rect 93 116 94 117
rect 92 116 93 117
rect 91 116 92 117
rect 82 116 83 117
rect 81 116 82 117
rect 80 116 81 117
rect 79 116 80 117
rect 78 116 79 117
rect 77 116 78 117
rect 76 116 77 117
rect 75 116 76 117
rect 74 116 75 117
rect 73 116 74 117
rect 72 116 73 117
rect 71 116 72 117
rect 70 116 71 117
rect 69 116 70 117
rect 68 116 69 117
rect 67 116 68 117
rect 66 116 67 117
rect 65 116 66 117
rect 64 116 65 117
rect 63 116 64 117
rect 62 116 63 117
rect 61 116 62 117
rect 60 116 61 117
rect 59 116 60 117
rect 58 116 59 117
rect 57 116 58 117
rect 56 116 57 117
rect 55 116 56 117
rect 49 116 50 117
rect 48 116 49 117
rect 47 116 48 117
rect 46 116 47 117
rect 45 116 46 117
rect 44 116 45 117
rect 43 116 44 117
rect 42 116 43 117
rect 41 116 42 117
rect 40 116 41 117
rect 39 116 40 117
rect 38 116 39 117
rect 37 116 38 117
rect 36 116 37 117
rect 35 116 36 117
rect 29 116 30 117
rect 28 116 29 117
rect 27 116 28 117
rect 26 116 27 117
rect 25 116 26 117
rect 24 116 25 117
rect 23 116 24 117
rect 22 116 23 117
rect 21 116 22 117
rect 20 116 21 117
rect 19 116 20 117
rect 18 116 19 117
rect 14 116 15 117
rect 13 116 14 117
rect 12 116 13 117
rect 11 116 12 117
rect 10 116 11 117
rect 9 116 10 117
rect 8 116 9 117
rect 7 116 8 117
rect 6 116 7 117
rect 5 116 6 117
rect 4 116 5 117
rect 188 117 189 118
rect 187 117 188 118
rect 178 117 179 118
rect 177 117 178 118
rect 176 117 177 118
rect 175 117 176 118
rect 174 117 175 118
rect 173 117 174 118
rect 172 117 173 118
rect 171 117 172 118
rect 170 117 171 118
rect 169 117 170 118
rect 168 117 169 118
rect 167 117 168 118
rect 166 117 167 118
rect 165 117 166 118
rect 164 117 165 118
rect 163 117 164 118
rect 162 117 163 118
rect 161 117 162 118
rect 117 117 118 118
rect 116 117 117 118
rect 115 117 116 118
rect 114 117 115 118
rect 113 117 114 118
rect 112 117 113 118
rect 111 117 112 118
rect 110 117 111 118
rect 109 117 110 118
rect 108 117 109 118
rect 107 117 108 118
rect 106 117 107 118
rect 105 117 106 118
rect 104 117 105 118
rect 103 117 104 118
rect 102 117 103 118
rect 101 117 102 118
rect 100 117 101 118
rect 99 117 100 118
rect 98 117 99 118
rect 97 117 98 118
rect 96 117 97 118
rect 95 117 96 118
rect 94 117 95 118
rect 93 117 94 118
rect 92 117 93 118
rect 91 117 92 118
rect 90 117 91 118
rect 81 117 82 118
rect 80 117 81 118
rect 79 117 80 118
rect 78 117 79 118
rect 77 117 78 118
rect 76 117 77 118
rect 75 117 76 118
rect 74 117 75 118
rect 73 117 74 118
rect 72 117 73 118
rect 71 117 72 118
rect 70 117 71 118
rect 69 117 70 118
rect 68 117 69 118
rect 67 117 68 118
rect 66 117 67 118
rect 65 117 66 118
rect 64 117 65 118
rect 63 117 64 118
rect 62 117 63 118
rect 61 117 62 118
rect 60 117 61 118
rect 59 117 60 118
rect 58 117 59 118
rect 57 117 58 118
rect 56 117 57 118
rect 49 117 50 118
rect 48 117 49 118
rect 47 117 48 118
rect 46 117 47 118
rect 45 117 46 118
rect 44 117 45 118
rect 43 117 44 118
rect 42 117 43 118
rect 41 117 42 118
rect 40 117 41 118
rect 39 117 40 118
rect 38 117 39 118
rect 37 117 38 118
rect 36 117 37 118
rect 29 117 30 118
rect 28 117 29 118
rect 27 117 28 118
rect 26 117 27 118
rect 25 117 26 118
rect 24 117 25 118
rect 23 117 24 118
rect 22 117 23 118
rect 21 117 22 118
rect 20 117 21 118
rect 19 117 20 118
rect 18 117 19 118
rect 14 117 15 118
rect 13 117 14 118
rect 12 117 13 118
rect 11 117 12 118
rect 10 117 11 118
rect 9 117 10 118
rect 8 117 9 118
rect 7 117 8 118
rect 6 117 7 118
rect 5 117 6 118
rect 4 117 5 118
rect 187 118 188 119
rect 178 118 179 119
rect 177 118 178 119
rect 176 118 177 119
rect 175 118 176 119
rect 174 118 175 119
rect 173 118 174 119
rect 172 118 173 119
rect 171 118 172 119
rect 170 118 171 119
rect 169 118 170 119
rect 168 118 169 119
rect 167 118 168 119
rect 166 118 167 119
rect 165 118 166 119
rect 164 118 165 119
rect 163 118 164 119
rect 162 118 163 119
rect 161 118 162 119
rect 116 118 117 119
rect 115 118 116 119
rect 114 118 115 119
rect 113 118 114 119
rect 112 118 113 119
rect 111 118 112 119
rect 110 118 111 119
rect 109 118 110 119
rect 108 118 109 119
rect 107 118 108 119
rect 106 118 107 119
rect 105 118 106 119
rect 104 118 105 119
rect 103 118 104 119
rect 102 118 103 119
rect 101 118 102 119
rect 100 118 101 119
rect 99 118 100 119
rect 98 118 99 119
rect 97 118 98 119
rect 96 118 97 119
rect 95 118 96 119
rect 94 118 95 119
rect 93 118 94 119
rect 92 118 93 119
rect 91 118 92 119
rect 90 118 91 119
rect 80 118 81 119
rect 79 118 80 119
rect 78 118 79 119
rect 77 118 78 119
rect 76 118 77 119
rect 75 118 76 119
rect 74 118 75 119
rect 73 118 74 119
rect 72 118 73 119
rect 71 118 72 119
rect 70 118 71 119
rect 69 118 70 119
rect 68 118 69 119
rect 67 118 68 119
rect 66 118 67 119
rect 65 118 66 119
rect 64 118 65 119
rect 63 118 64 119
rect 62 118 63 119
rect 61 118 62 119
rect 60 118 61 119
rect 59 118 60 119
rect 58 118 59 119
rect 57 118 58 119
rect 56 118 57 119
rect 49 118 50 119
rect 48 118 49 119
rect 47 118 48 119
rect 46 118 47 119
rect 45 118 46 119
rect 44 118 45 119
rect 43 118 44 119
rect 42 118 43 119
rect 41 118 42 119
rect 40 118 41 119
rect 39 118 40 119
rect 38 118 39 119
rect 37 118 38 119
rect 36 118 37 119
rect 29 118 30 119
rect 28 118 29 119
rect 27 118 28 119
rect 26 118 27 119
rect 25 118 26 119
rect 24 118 25 119
rect 23 118 24 119
rect 22 118 23 119
rect 21 118 22 119
rect 20 118 21 119
rect 19 118 20 119
rect 18 118 19 119
rect 15 118 16 119
rect 14 118 15 119
rect 13 118 14 119
rect 12 118 13 119
rect 11 118 12 119
rect 10 118 11 119
rect 9 118 10 119
rect 8 118 9 119
rect 7 118 8 119
rect 6 118 7 119
rect 5 118 6 119
rect 4 118 5 119
rect 178 119 179 120
rect 177 119 178 120
rect 170 119 171 120
rect 169 119 170 120
rect 168 119 169 120
rect 163 119 164 120
rect 162 119 163 120
rect 161 119 162 120
rect 115 119 116 120
rect 114 119 115 120
rect 113 119 114 120
rect 112 119 113 120
rect 111 119 112 120
rect 110 119 111 120
rect 109 119 110 120
rect 108 119 109 120
rect 107 119 108 120
rect 106 119 107 120
rect 105 119 106 120
rect 104 119 105 120
rect 103 119 104 120
rect 102 119 103 120
rect 101 119 102 120
rect 100 119 101 120
rect 99 119 100 120
rect 98 119 99 120
rect 97 119 98 120
rect 96 119 97 120
rect 95 119 96 120
rect 94 119 95 120
rect 93 119 94 120
rect 92 119 93 120
rect 91 119 92 120
rect 90 119 91 120
rect 89 119 90 120
rect 80 119 81 120
rect 79 119 80 120
rect 78 119 79 120
rect 77 119 78 120
rect 76 119 77 120
rect 75 119 76 120
rect 74 119 75 120
rect 73 119 74 120
rect 72 119 73 120
rect 71 119 72 120
rect 70 119 71 120
rect 69 119 70 120
rect 68 119 69 120
rect 67 119 68 120
rect 66 119 67 120
rect 65 119 66 120
rect 64 119 65 120
rect 63 119 64 120
rect 62 119 63 120
rect 61 119 62 120
rect 60 119 61 120
rect 59 119 60 120
rect 58 119 59 120
rect 57 119 58 120
rect 50 119 51 120
rect 49 119 50 120
rect 48 119 49 120
rect 47 119 48 120
rect 46 119 47 120
rect 45 119 46 120
rect 44 119 45 120
rect 43 119 44 120
rect 42 119 43 120
rect 41 119 42 120
rect 40 119 41 120
rect 39 119 40 120
rect 38 119 39 120
rect 37 119 38 120
rect 36 119 37 120
rect 30 119 31 120
rect 29 119 30 120
rect 28 119 29 120
rect 27 119 28 120
rect 26 119 27 120
rect 25 119 26 120
rect 24 119 25 120
rect 23 119 24 120
rect 22 119 23 120
rect 21 119 22 120
rect 20 119 21 120
rect 19 119 20 120
rect 18 119 19 120
rect 15 119 16 120
rect 14 119 15 120
rect 13 119 14 120
rect 12 119 13 120
rect 11 119 12 120
rect 10 119 11 120
rect 9 119 10 120
rect 8 119 9 120
rect 7 119 8 120
rect 6 119 7 120
rect 5 119 6 120
rect 4 119 5 120
rect 195 120 196 121
rect 194 120 195 121
rect 193 120 194 121
rect 192 120 193 121
rect 191 120 192 121
rect 190 120 191 121
rect 189 120 190 121
rect 188 120 189 121
rect 187 120 188 121
rect 178 120 179 121
rect 169 120 170 121
rect 168 120 169 121
rect 161 120 162 121
rect 114 120 115 121
rect 113 120 114 121
rect 112 120 113 121
rect 111 120 112 121
rect 110 120 111 121
rect 109 120 110 121
rect 108 120 109 121
rect 107 120 108 121
rect 106 120 107 121
rect 105 120 106 121
rect 104 120 105 121
rect 103 120 104 121
rect 102 120 103 121
rect 101 120 102 121
rect 100 120 101 121
rect 99 120 100 121
rect 98 120 99 121
rect 97 120 98 121
rect 96 120 97 121
rect 95 120 96 121
rect 94 120 95 121
rect 93 120 94 121
rect 92 120 93 121
rect 91 120 92 121
rect 90 120 91 121
rect 89 120 90 121
rect 88 120 89 121
rect 79 120 80 121
rect 78 120 79 121
rect 77 120 78 121
rect 76 120 77 121
rect 75 120 76 121
rect 74 120 75 121
rect 73 120 74 121
rect 72 120 73 121
rect 71 120 72 121
rect 70 120 71 121
rect 69 120 70 121
rect 68 120 69 121
rect 67 120 68 121
rect 66 120 67 121
rect 65 120 66 121
rect 64 120 65 121
rect 63 120 64 121
rect 62 120 63 121
rect 61 120 62 121
rect 60 120 61 121
rect 59 120 60 121
rect 58 120 59 121
rect 57 120 58 121
rect 50 120 51 121
rect 49 120 50 121
rect 48 120 49 121
rect 47 120 48 121
rect 46 120 47 121
rect 45 120 46 121
rect 44 120 45 121
rect 43 120 44 121
rect 42 120 43 121
rect 41 120 42 121
rect 40 120 41 121
rect 39 120 40 121
rect 38 120 39 121
rect 37 120 38 121
rect 36 120 37 121
rect 30 120 31 121
rect 29 120 30 121
rect 28 120 29 121
rect 27 120 28 121
rect 26 120 27 121
rect 25 120 26 121
rect 24 120 25 121
rect 23 120 24 121
rect 22 120 23 121
rect 21 120 22 121
rect 20 120 21 121
rect 19 120 20 121
rect 15 120 16 121
rect 14 120 15 121
rect 13 120 14 121
rect 12 120 13 121
rect 11 120 12 121
rect 10 120 11 121
rect 9 120 10 121
rect 8 120 9 121
rect 7 120 8 121
rect 6 120 7 121
rect 5 120 6 121
rect 4 120 5 121
rect 194 121 195 122
rect 193 121 194 122
rect 192 121 193 122
rect 191 121 192 122
rect 190 121 191 122
rect 189 121 190 122
rect 188 121 189 122
rect 187 121 188 122
rect 178 121 179 122
rect 169 121 170 122
rect 168 121 169 122
rect 161 121 162 122
rect 113 121 114 122
rect 112 121 113 122
rect 111 121 112 122
rect 110 121 111 122
rect 109 121 110 122
rect 108 121 109 122
rect 107 121 108 122
rect 106 121 107 122
rect 105 121 106 122
rect 104 121 105 122
rect 103 121 104 122
rect 102 121 103 122
rect 101 121 102 122
rect 100 121 101 122
rect 99 121 100 122
rect 98 121 99 122
rect 97 121 98 122
rect 96 121 97 122
rect 95 121 96 122
rect 94 121 95 122
rect 93 121 94 122
rect 92 121 93 122
rect 91 121 92 122
rect 90 121 91 122
rect 89 121 90 122
rect 88 121 89 122
rect 78 121 79 122
rect 77 121 78 122
rect 76 121 77 122
rect 75 121 76 122
rect 74 121 75 122
rect 73 121 74 122
rect 72 121 73 122
rect 71 121 72 122
rect 70 121 71 122
rect 69 121 70 122
rect 68 121 69 122
rect 67 121 68 122
rect 66 121 67 122
rect 65 121 66 122
rect 64 121 65 122
rect 63 121 64 122
rect 62 121 63 122
rect 61 121 62 122
rect 60 121 61 122
rect 59 121 60 122
rect 58 121 59 122
rect 51 121 52 122
rect 50 121 51 122
rect 49 121 50 122
rect 48 121 49 122
rect 47 121 48 122
rect 46 121 47 122
rect 45 121 46 122
rect 44 121 45 122
rect 43 121 44 122
rect 42 121 43 122
rect 41 121 42 122
rect 40 121 41 122
rect 39 121 40 122
rect 38 121 39 122
rect 37 121 38 122
rect 30 121 31 122
rect 29 121 30 122
rect 28 121 29 122
rect 27 121 28 122
rect 26 121 27 122
rect 25 121 26 122
rect 24 121 25 122
rect 23 121 24 122
rect 22 121 23 122
rect 21 121 22 122
rect 20 121 21 122
rect 19 121 20 122
rect 15 121 16 122
rect 14 121 15 122
rect 13 121 14 122
rect 12 121 13 122
rect 11 121 12 122
rect 10 121 11 122
rect 9 121 10 122
rect 8 121 9 122
rect 7 121 8 122
rect 6 121 7 122
rect 5 121 6 122
rect 194 122 195 123
rect 192 122 193 123
rect 191 122 192 123
rect 190 122 191 123
rect 189 122 190 123
rect 187 122 188 123
rect 169 122 170 123
rect 168 122 169 123
rect 112 122 113 123
rect 111 122 112 123
rect 110 122 111 123
rect 109 122 110 123
rect 108 122 109 123
rect 107 122 108 123
rect 106 122 107 123
rect 105 122 106 123
rect 104 122 105 123
rect 103 122 104 123
rect 102 122 103 123
rect 101 122 102 123
rect 100 122 101 123
rect 99 122 100 123
rect 98 122 99 123
rect 97 122 98 123
rect 96 122 97 123
rect 95 122 96 123
rect 94 122 95 123
rect 93 122 94 123
rect 92 122 93 123
rect 91 122 92 123
rect 90 122 91 123
rect 89 122 90 123
rect 88 122 89 123
rect 87 122 88 123
rect 77 122 78 123
rect 76 122 77 123
rect 75 122 76 123
rect 74 122 75 123
rect 73 122 74 123
rect 72 122 73 123
rect 71 122 72 123
rect 70 122 71 123
rect 69 122 70 123
rect 68 122 69 123
rect 67 122 68 123
rect 66 122 67 123
rect 65 122 66 123
rect 64 122 65 123
rect 63 122 64 123
rect 62 122 63 123
rect 61 122 62 123
rect 60 122 61 123
rect 59 122 60 123
rect 51 122 52 123
rect 50 122 51 123
rect 49 122 50 123
rect 48 122 49 123
rect 47 122 48 123
rect 46 122 47 123
rect 45 122 46 123
rect 44 122 45 123
rect 43 122 44 123
rect 42 122 43 123
rect 41 122 42 123
rect 40 122 41 123
rect 39 122 40 123
rect 38 122 39 123
rect 37 122 38 123
rect 30 122 31 123
rect 29 122 30 123
rect 28 122 29 123
rect 27 122 28 123
rect 26 122 27 123
rect 25 122 26 123
rect 24 122 25 123
rect 23 122 24 123
rect 22 122 23 123
rect 21 122 22 123
rect 20 122 21 123
rect 19 122 20 123
rect 15 122 16 123
rect 14 122 15 123
rect 13 122 14 123
rect 12 122 13 123
rect 11 122 12 123
rect 10 122 11 123
rect 9 122 10 123
rect 8 122 9 123
rect 7 122 8 123
rect 6 122 7 123
rect 5 122 6 123
rect 187 123 188 124
rect 169 123 170 124
rect 168 123 169 124
rect 111 123 112 124
rect 110 123 111 124
rect 109 123 110 124
rect 108 123 109 124
rect 107 123 108 124
rect 106 123 107 124
rect 105 123 106 124
rect 104 123 105 124
rect 103 123 104 124
rect 102 123 103 124
rect 101 123 102 124
rect 100 123 101 124
rect 99 123 100 124
rect 98 123 99 124
rect 97 123 98 124
rect 96 123 97 124
rect 95 123 96 124
rect 94 123 95 124
rect 93 123 94 124
rect 92 123 93 124
rect 91 123 92 124
rect 90 123 91 124
rect 89 123 90 124
rect 88 123 89 124
rect 87 123 88 124
rect 86 123 87 124
rect 76 123 77 124
rect 75 123 76 124
rect 74 123 75 124
rect 73 123 74 124
rect 72 123 73 124
rect 71 123 72 124
rect 70 123 71 124
rect 69 123 70 124
rect 68 123 69 124
rect 67 123 68 124
rect 66 123 67 124
rect 65 123 66 124
rect 64 123 65 124
rect 63 123 64 124
rect 62 123 63 124
rect 61 123 62 124
rect 60 123 61 124
rect 51 123 52 124
rect 50 123 51 124
rect 49 123 50 124
rect 48 123 49 124
rect 47 123 48 124
rect 46 123 47 124
rect 45 123 46 124
rect 44 123 45 124
rect 43 123 44 124
rect 42 123 43 124
rect 41 123 42 124
rect 40 123 41 124
rect 39 123 40 124
rect 38 123 39 124
rect 37 123 38 124
rect 31 123 32 124
rect 30 123 31 124
rect 29 123 30 124
rect 28 123 29 124
rect 27 123 28 124
rect 26 123 27 124
rect 25 123 26 124
rect 24 123 25 124
rect 23 123 24 124
rect 22 123 23 124
rect 21 123 22 124
rect 20 123 21 124
rect 19 123 20 124
rect 15 123 16 124
rect 14 123 15 124
rect 13 123 14 124
rect 12 123 13 124
rect 11 123 12 124
rect 10 123 11 124
rect 9 123 10 124
rect 8 123 9 124
rect 7 123 8 124
rect 6 123 7 124
rect 5 123 6 124
rect 188 124 189 125
rect 187 124 188 125
rect 186 124 187 125
rect 178 124 179 125
rect 169 124 170 125
rect 168 124 169 125
rect 161 124 162 125
rect 109 124 110 125
rect 108 124 109 125
rect 107 124 108 125
rect 106 124 107 125
rect 105 124 106 125
rect 104 124 105 125
rect 103 124 104 125
rect 102 124 103 125
rect 101 124 102 125
rect 100 124 101 125
rect 99 124 100 125
rect 98 124 99 125
rect 97 124 98 125
rect 96 124 97 125
rect 95 124 96 125
rect 94 124 95 125
rect 93 124 94 125
rect 92 124 93 125
rect 91 124 92 125
rect 90 124 91 125
rect 89 124 90 125
rect 88 124 89 125
rect 87 124 88 125
rect 86 124 87 125
rect 74 124 75 125
rect 73 124 74 125
rect 72 124 73 125
rect 71 124 72 125
rect 70 124 71 125
rect 69 124 70 125
rect 68 124 69 125
rect 67 124 68 125
rect 66 124 67 125
rect 65 124 66 125
rect 64 124 65 125
rect 63 124 64 125
rect 62 124 63 125
rect 52 124 53 125
rect 51 124 52 125
rect 50 124 51 125
rect 49 124 50 125
rect 48 124 49 125
rect 47 124 48 125
rect 46 124 47 125
rect 45 124 46 125
rect 44 124 45 125
rect 43 124 44 125
rect 42 124 43 125
rect 41 124 42 125
rect 40 124 41 125
rect 39 124 40 125
rect 38 124 39 125
rect 37 124 38 125
rect 31 124 32 125
rect 30 124 31 125
rect 29 124 30 125
rect 28 124 29 125
rect 27 124 28 125
rect 26 124 27 125
rect 25 124 26 125
rect 24 124 25 125
rect 23 124 24 125
rect 22 124 23 125
rect 21 124 22 125
rect 20 124 21 125
rect 15 124 16 125
rect 14 124 15 125
rect 13 124 14 125
rect 12 124 13 125
rect 11 124 12 125
rect 10 124 11 125
rect 9 124 10 125
rect 8 124 9 125
rect 7 124 8 125
rect 6 124 7 125
rect 178 125 179 126
rect 169 125 170 126
rect 168 125 169 126
rect 161 125 162 126
rect 108 125 109 126
rect 107 125 108 126
rect 106 125 107 126
rect 105 125 106 126
rect 104 125 105 126
rect 103 125 104 126
rect 102 125 103 126
rect 101 125 102 126
rect 100 125 101 126
rect 99 125 100 126
rect 98 125 99 126
rect 97 125 98 126
rect 96 125 97 126
rect 95 125 96 126
rect 94 125 95 126
rect 93 125 94 126
rect 92 125 93 126
rect 91 125 92 126
rect 90 125 91 126
rect 89 125 90 126
rect 88 125 89 126
rect 87 125 88 126
rect 86 125 87 126
rect 85 125 86 126
rect 73 125 74 126
rect 72 125 73 126
rect 71 125 72 126
rect 70 125 71 126
rect 69 125 70 126
rect 68 125 69 126
rect 67 125 68 126
rect 66 125 67 126
rect 65 125 66 126
rect 64 125 65 126
rect 52 125 53 126
rect 51 125 52 126
rect 50 125 51 126
rect 49 125 50 126
rect 48 125 49 126
rect 47 125 48 126
rect 46 125 47 126
rect 45 125 46 126
rect 44 125 45 126
rect 43 125 44 126
rect 42 125 43 126
rect 41 125 42 126
rect 40 125 41 126
rect 39 125 40 126
rect 38 125 39 126
rect 31 125 32 126
rect 30 125 31 126
rect 29 125 30 126
rect 28 125 29 126
rect 27 125 28 126
rect 26 125 27 126
rect 25 125 26 126
rect 24 125 25 126
rect 23 125 24 126
rect 22 125 23 126
rect 21 125 22 126
rect 20 125 21 126
rect 15 125 16 126
rect 14 125 15 126
rect 13 125 14 126
rect 12 125 13 126
rect 11 125 12 126
rect 10 125 11 126
rect 9 125 10 126
rect 8 125 9 126
rect 7 125 8 126
rect 6 125 7 126
rect 178 126 179 127
rect 177 126 178 127
rect 170 126 171 127
rect 169 126 170 127
rect 168 126 169 127
rect 162 126 163 127
rect 161 126 162 127
rect 107 126 108 127
rect 106 126 107 127
rect 105 126 106 127
rect 104 126 105 127
rect 103 126 104 127
rect 102 126 103 127
rect 101 126 102 127
rect 100 126 101 127
rect 99 126 100 127
rect 98 126 99 127
rect 97 126 98 127
rect 96 126 97 127
rect 95 126 96 127
rect 94 126 95 127
rect 93 126 94 127
rect 92 126 93 127
rect 91 126 92 127
rect 90 126 91 127
rect 89 126 90 127
rect 88 126 89 127
rect 87 126 88 127
rect 86 126 87 127
rect 85 126 86 127
rect 84 126 85 127
rect 70 126 71 127
rect 69 126 70 127
rect 68 126 69 127
rect 67 126 68 127
rect 66 126 67 127
rect 53 126 54 127
rect 52 126 53 127
rect 51 126 52 127
rect 50 126 51 127
rect 49 126 50 127
rect 48 126 49 127
rect 47 126 48 127
rect 46 126 47 127
rect 45 126 46 127
rect 44 126 45 127
rect 43 126 44 127
rect 42 126 43 127
rect 41 126 42 127
rect 40 126 41 127
rect 39 126 40 127
rect 38 126 39 127
rect 32 126 33 127
rect 31 126 32 127
rect 30 126 31 127
rect 29 126 30 127
rect 28 126 29 127
rect 27 126 28 127
rect 26 126 27 127
rect 25 126 26 127
rect 24 126 25 127
rect 23 126 24 127
rect 22 126 23 127
rect 21 126 22 127
rect 20 126 21 127
rect 16 126 17 127
rect 15 126 16 127
rect 14 126 15 127
rect 13 126 14 127
rect 12 126 13 127
rect 11 126 12 127
rect 10 126 11 127
rect 9 126 10 127
rect 8 126 9 127
rect 7 126 8 127
rect 178 127 179 128
rect 177 127 178 128
rect 176 127 177 128
rect 175 127 176 128
rect 174 127 175 128
rect 173 127 174 128
rect 172 127 173 128
rect 171 127 172 128
rect 170 127 171 128
rect 169 127 170 128
rect 168 127 169 128
rect 167 127 168 128
rect 166 127 167 128
rect 165 127 166 128
rect 164 127 165 128
rect 163 127 164 128
rect 162 127 163 128
rect 161 127 162 128
rect 105 127 106 128
rect 104 127 105 128
rect 103 127 104 128
rect 102 127 103 128
rect 101 127 102 128
rect 100 127 101 128
rect 99 127 100 128
rect 98 127 99 128
rect 97 127 98 128
rect 96 127 97 128
rect 95 127 96 128
rect 94 127 95 128
rect 93 127 94 128
rect 92 127 93 128
rect 91 127 92 128
rect 90 127 91 128
rect 89 127 90 128
rect 88 127 89 128
rect 87 127 88 128
rect 86 127 87 128
rect 85 127 86 128
rect 84 127 85 128
rect 83 127 84 128
rect 54 127 55 128
rect 53 127 54 128
rect 52 127 53 128
rect 51 127 52 128
rect 50 127 51 128
rect 49 127 50 128
rect 48 127 49 128
rect 47 127 48 128
rect 46 127 47 128
rect 45 127 46 128
rect 44 127 45 128
rect 43 127 44 128
rect 42 127 43 128
rect 41 127 42 128
rect 40 127 41 128
rect 39 127 40 128
rect 32 127 33 128
rect 31 127 32 128
rect 30 127 31 128
rect 29 127 30 128
rect 28 127 29 128
rect 27 127 28 128
rect 26 127 27 128
rect 25 127 26 128
rect 24 127 25 128
rect 23 127 24 128
rect 22 127 23 128
rect 21 127 22 128
rect 16 127 17 128
rect 15 127 16 128
rect 14 127 15 128
rect 13 127 14 128
rect 12 127 13 128
rect 11 127 12 128
rect 10 127 11 128
rect 9 127 10 128
rect 8 127 9 128
rect 7 127 8 128
rect 178 128 179 129
rect 177 128 178 129
rect 176 128 177 129
rect 175 128 176 129
rect 174 128 175 129
rect 173 128 174 129
rect 172 128 173 129
rect 171 128 172 129
rect 170 128 171 129
rect 169 128 170 129
rect 168 128 169 129
rect 167 128 168 129
rect 166 128 167 129
rect 165 128 166 129
rect 164 128 165 129
rect 163 128 164 129
rect 162 128 163 129
rect 161 128 162 129
rect 103 128 104 129
rect 102 128 103 129
rect 101 128 102 129
rect 100 128 101 129
rect 99 128 100 129
rect 98 128 99 129
rect 97 128 98 129
rect 96 128 97 129
rect 95 128 96 129
rect 94 128 95 129
rect 93 128 94 129
rect 92 128 93 129
rect 91 128 92 129
rect 90 128 91 129
rect 89 128 90 129
rect 88 128 89 129
rect 87 128 88 129
rect 86 128 87 129
rect 85 128 86 129
rect 84 128 85 129
rect 83 128 84 129
rect 82 128 83 129
rect 55 128 56 129
rect 54 128 55 129
rect 53 128 54 129
rect 52 128 53 129
rect 51 128 52 129
rect 50 128 51 129
rect 49 128 50 129
rect 48 128 49 129
rect 47 128 48 129
rect 46 128 47 129
rect 45 128 46 129
rect 44 128 45 129
rect 43 128 44 129
rect 42 128 43 129
rect 41 128 42 129
rect 40 128 41 129
rect 39 128 40 129
rect 32 128 33 129
rect 31 128 32 129
rect 30 128 31 129
rect 29 128 30 129
rect 28 128 29 129
rect 27 128 28 129
rect 26 128 27 129
rect 25 128 26 129
rect 24 128 25 129
rect 23 128 24 129
rect 22 128 23 129
rect 21 128 22 129
rect 16 128 17 129
rect 15 128 16 129
rect 14 128 15 129
rect 13 128 14 129
rect 12 128 13 129
rect 11 128 12 129
rect 10 128 11 129
rect 9 128 10 129
rect 8 128 9 129
rect 187 129 188 130
rect 178 129 179 130
rect 177 129 178 130
rect 176 129 177 130
rect 175 129 176 130
rect 174 129 175 130
rect 173 129 174 130
rect 172 129 173 130
rect 171 129 172 130
rect 170 129 171 130
rect 169 129 170 130
rect 168 129 169 130
rect 167 129 168 130
rect 166 129 167 130
rect 165 129 166 130
rect 164 129 165 130
rect 163 129 164 130
rect 162 129 163 130
rect 161 129 162 130
rect 101 129 102 130
rect 100 129 101 130
rect 99 129 100 130
rect 98 129 99 130
rect 97 129 98 130
rect 96 129 97 130
rect 95 129 96 130
rect 94 129 95 130
rect 93 129 94 130
rect 92 129 93 130
rect 91 129 92 130
rect 90 129 91 130
rect 89 129 90 130
rect 88 129 89 130
rect 87 129 88 130
rect 86 129 87 130
rect 85 129 86 130
rect 84 129 85 130
rect 83 129 84 130
rect 82 129 83 130
rect 81 129 82 130
rect 56 129 57 130
rect 55 129 56 130
rect 54 129 55 130
rect 53 129 54 130
rect 52 129 53 130
rect 51 129 52 130
rect 50 129 51 130
rect 49 129 50 130
rect 48 129 49 130
rect 47 129 48 130
rect 46 129 47 130
rect 45 129 46 130
rect 44 129 45 130
rect 43 129 44 130
rect 42 129 43 130
rect 41 129 42 130
rect 40 129 41 130
rect 33 129 34 130
rect 32 129 33 130
rect 31 129 32 130
rect 30 129 31 130
rect 29 129 30 130
rect 28 129 29 130
rect 27 129 28 130
rect 26 129 27 130
rect 25 129 26 130
rect 24 129 25 130
rect 23 129 24 130
rect 22 129 23 130
rect 21 129 22 130
rect 16 129 17 130
rect 15 129 16 130
rect 14 129 15 130
rect 13 129 14 130
rect 12 129 13 130
rect 11 129 12 130
rect 10 129 11 130
rect 9 129 10 130
rect 8 129 9 130
rect 189 130 190 131
rect 188 130 189 131
rect 187 130 188 131
rect 178 130 179 131
rect 177 130 178 131
rect 176 130 177 131
rect 175 130 176 131
rect 174 130 175 131
rect 173 130 174 131
rect 172 130 173 131
rect 171 130 172 131
rect 170 130 171 131
rect 169 130 170 131
rect 168 130 169 131
rect 167 130 168 131
rect 166 130 167 131
rect 165 130 166 131
rect 164 130 165 131
rect 163 130 164 131
rect 162 130 163 131
rect 161 130 162 131
rect 99 130 100 131
rect 98 130 99 131
rect 97 130 98 131
rect 96 130 97 131
rect 95 130 96 131
rect 94 130 95 131
rect 93 130 94 131
rect 92 130 93 131
rect 91 130 92 131
rect 90 130 91 131
rect 89 130 90 131
rect 88 130 89 131
rect 87 130 88 131
rect 86 130 87 131
rect 85 130 86 131
rect 84 130 85 131
rect 83 130 84 131
rect 82 130 83 131
rect 81 130 82 131
rect 80 130 81 131
rect 57 130 58 131
rect 56 130 57 131
rect 55 130 56 131
rect 54 130 55 131
rect 53 130 54 131
rect 52 130 53 131
rect 51 130 52 131
rect 50 130 51 131
rect 49 130 50 131
rect 48 130 49 131
rect 47 130 48 131
rect 46 130 47 131
rect 45 130 46 131
rect 44 130 45 131
rect 43 130 44 131
rect 42 130 43 131
rect 41 130 42 131
rect 33 130 34 131
rect 32 130 33 131
rect 31 130 32 131
rect 30 130 31 131
rect 29 130 30 131
rect 28 130 29 131
rect 27 130 28 131
rect 26 130 27 131
rect 25 130 26 131
rect 24 130 25 131
rect 23 130 24 131
rect 22 130 23 131
rect 17 130 18 131
rect 16 130 17 131
rect 15 130 16 131
rect 14 130 15 131
rect 13 130 14 131
rect 12 130 13 131
rect 11 130 12 131
rect 10 130 11 131
rect 9 130 10 131
rect 195 131 196 132
rect 194 131 195 132
rect 193 131 194 132
rect 192 131 193 132
rect 191 131 192 132
rect 190 131 191 132
rect 189 131 190 132
rect 188 131 189 132
rect 187 131 188 132
rect 178 131 179 132
rect 177 131 178 132
rect 161 131 162 132
rect 96 131 97 132
rect 95 131 96 132
rect 94 131 95 132
rect 93 131 94 132
rect 92 131 93 132
rect 91 131 92 132
rect 90 131 91 132
rect 89 131 90 132
rect 88 131 89 132
rect 87 131 88 132
rect 86 131 87 132
rect 85 131 86 132
rect 84 131 85 132
rect 83 131 84 132
rect 82 131 83 132
rect 81 131 82 132
rect 80 131 81 132
rect 79 131 80 132
rect 59 131 60 132
rect 58 131 59 132
rect 57 131 58 132
rect 56 131 57 132
rect 55 131 56 132
rect 54 131 55 132
rect 53 131 54 132
rect 52 131 53 132
rect 51 131 52 132
rect 50 131 51 132
rect 49 131 50 132
rect 48 131 49 132
rect 47 131 48 132
rect 46 131 47 132
rect 45 131 46 132
rect 44 131 45 132
rect 43 131 44 132
rect 42 131 43 132
rect 41 131 42 132
rect 34 131 35 132
rect 33 131 34 132
rect 32 131 33 132
rect 31 131 32 132
rect 30 131 31 132
rect 29 131 30 132
rect 28 131 29 132
rect 27 131 28 132
rect 26 131 27 132
rect 25 131 26 132
rect 24 131 25 132
rect 23 131 24 132
rect 22 131 23 132
rect 17 131 18 132
rect 16 131 17 132
rect 15 131 16 132
rect 14 131 15 132
rect 13 131 14 132
rect 12 131 13 132
rect 11 131 12 132
rect 10 131 11 132
rect 194 132 195 133
rect 193 132 194 133
rect 192 132 193 133
rect 191 132 192 133
rect 190 132 191 133
rect 178 132 179 133
rect 161 132 162 133
rect 91 132 92 133
rect 90 132 91 133
rect 89 132 90 133
rect 88 132 89 133
rect 87 132 88 133
rect 86 132 87 133
rect 85 132 86 133
rect 84 132 85 133
rect 83 132 84 133
rect 81 132 82 133
rect 60 132 61 133
rect 59 132 60 133
rect 58 132 59 133
rect 57 132 58 133
rect 56 132 57 133
rect 55 132 56 133
rect 54 132 55 133
rect 53 132 54 133
rect 52 132 53 133
rect 51 132 52 133
rect 50 132 51 133
rect 49 132 50 133
rect 48 132 49 133
rect 47 132 48 133
rect 46 132 47 133
rect 45 132 46 133
rect 44 132 45 133
rect 43 132 44 133
rect 42 132 43 133
rect 34 132 35 133
rect 33 132 34 133
rect 32 132 33 133
rect 31 132 32 133
rect 30 132 31 133
rect 29 132 30 133
rect 28 132 29 133
rect 27 132 28 133
rect 26 132 27 133
rect 25 132 26 133
rect 24 132 25 133
rect 23 132 24 133
rect 22 132 23 133
rect 17 132 18 133
rect 16 132 17 133
rect 15 132 16 133
rect 14 132 15 133
rect 13 132 14 133
rect 12 132 13 133
rect 11 132 12 133
rect 194 133 195 134
rect 193 133 194 134
rect 192 133 193 134
rect 191 133 192 134
rect 190 133 191 134
rect 189 133 190 134
rect 62 133 63 134
rect 61 133 62 134
rect 60 133 61 134
rect 59 133 60 134
rect 58 133 59 134
rect 57 133 58 134
rect 56 133 57 134
rect 55 133 56 134
rect 54 133 55 134
rect 53 133 54 134
rect 52 133 53 134
rect 51 133 52 134
rect 50 133 51 134
rect 49 133 50 134
rect 48 133 49 134
rect 47 133 48 134
rect 46 133 47 134
rect 45 133 46 134
rect 44 133 45 134
rect 43 133 44 134
rect 35 133 36 134
rect 34 133 35 134
rect 33 133 34 134
rect 32 133 33 134
rect 31 133 32 134
rect 30 133 31 134
rect 29 133 30 134
rect 28 133 29 134
rect 27 133 28 134
rect 26 133 27 134
rect 25 133 26 134
rect 24 133 25 134
rect 23 133 24 134
rect 18 133 19 134
rect 17 133 18 134
rect 16 133 17 134
rect 15 133 16 134
rect 14 133 15 134
rect 13 133 14 134
rect 12 133 13 134
rect 11 133 12 134
rect 189 134 190 135
rect 188 134 189 135
rect 187 134 188 135
rect 64 134 65 135
rect 63 134 64 135
rect 62 134 63 135
rect 61 134 62 135
rect 60 134 61 135
rect 59 134 60 135
rect 58 134 59 135
rect 57 134 58 135
rect 56 134 57 135
rect 55 134 56 135
rect 54 134 55 135
rect 53 134 54 135
rect 52 134 53 135
rect 51 134 52 135
rect 50 134 51 135
rect 49 134 50 135
rect 48 134 49 135
rect 47 134 48 135
rect 46 134 47 135
rect 45 134 46 135
rect 44 134 45 135
rect 36 134 37 135
rect 35 134 36 135
rect 34 134 35 135
rect 33 134 34 135
rect 32 134 33 135
rect 31 134 32 135
rect 30 134 31 135
rect 29 134 30 135
rect 28 134 29 135
rect 27 134 28 135
rect 26 134 27 135
rect 25 134 26 135
rect 24 134 25 135
rect 23 134 24 135
rect 18 134 19 135
rect 17 134 18 135
rect 16 134 17 135
rect 15 134 16 135
rect 14 134 15 135
rect 13 134 14 135
rect 12 134 13 135
rect 187 135 188 136
rect 67 135 68 136
rect 66 135 67 136
rect 65 135 66 136
rect 64 135 65 136
rect 63 135 64 136
rect 62 135 63 136
rect 61 135 62 136
rect 60 135 61 136
rect 59 135 60 136
rect 58 135 59 136
rect 57 135 58 136
rect 56 135 57 136
rect 55 135 56 136
rect 54 135 55 136
rect 53 135 54 136
rect 52 135 53 136
rect 51 135 52 136
rect 50 135 51 136
rect 49 135 50 136
rect 48 135 49 136
rect 47 135 48 136
rect 46 135 47 136
rect 45 135 46 136
rect 36 135 37 136
rect 35 135 36 136
rect 34 135 35 136
rect 33 135 34 136
rect 32 135 33 136
rect 31 135 32 136
rect 30 135 31 136
rect 29 135 30 136
rect 28 135 29 136
rect 27 135 28 136
rect 26 135 27 136
rect 25 135 26 136
rect 24 135 25 136
rect 23 135 24 136
rect 18 135 19 136
rect 17 135 18 136
rect 16 135 17 136
rect 15 135 16 136
rect 14 135 15 136
rect 13 135 14 136
rect 178 136 179 137
rect 161 136 162 137
rect 70 136 71 137
rect 69 136 70 137
rect 68 136 69 137
rect 67 136 68 137
rect 66 136 67 137
rect 65 136 66 137
rect 64 136 65 137
rect 63 136 64 137
rect 62 136 63 137
rect 61 136 62 137
rect 60 136 61 137
rect 59 136 60 137
rect 58 136 59 137
rect 57 136 58 137
rect 56 136 57 137
rect 55 136 56 137
rect 54 136 55 137
rect 53 136 54 137
rect 52 136 53 137
rect 51 136 52 137
rect 50 136 51 137
rect 49 136 50 137
rect 48 136 49 137
rect 47 136 48 137
rect 46 136 47 137
rect 45 136 46 137
rect 37 136 38 137
rect 36 136 37 137
rect 35 136 36 137
rect 34 136 35 137
rect 33 136 34 137
rect 32 136 33 137
rect 31 136 32 137
rect 30 136 31 137
rect 29 136 30 137
rect 28 136 29 137
rect 27 136 28 137
rect 26 136 27 137
rect 25 136 26 137
rect 24 136 25 137
rect 19 136 20 137
rect 18 136 19 137
rect 17 136 18 137
rect 16 136 17 137
rect 15 136 16 137
rect 14 136 15 137
rect 178 137 179 138
rect 161 137 162 138
rect 74 137 75 138
rect 73 137 74 138
rect 72 137 73 138
rect 71 137 72 138
rect 70 137 71 138
rect 69 137 70 138
rect 68 137 69 138
rect 67 137 68 138
rect 66 137 67 138
rect 65 137 66 138
rect 64 137 65 138
rect 63 137 64 138
rect 62 137 63 138
rect 61 137 62 138
rect 60 137 61 138
rect 59 137 60 138
rect 58 137 59 138
rect 57 137 58 138
rect 56 137 57 138
rect 55 137 56 138
rect 54 137 55 138
rect 53 137 54 138
rect 52 137 53 138
rect 51 137 52 138
rect 50 137 51 138
rect 49 137 50 138
rect 48 137 49 138
rect 47 137 48 138
rect 46 137 47 138
rect 38 137 39 138
rect 37 137 38 138
rect 36 137 37 138
rect 35 137 36 138
rect 34 137 35 138
rect 33 137 34 138
rect 32 137 33 138
rect 31 137 32 138
rect 30 137 31 138
rect 29 137 30 138
rect 28 137 29 138
rect 27 137 28 138
rect 26 137 27 138
rect 25 137 26 138
rect 24 137 25 138
rect 19 137 20 138
rect 18 137 19 138
rect 17 137 18 138
rect 16 137 17 138
rect 15 137 16 138
rect 178 138 179 139
rect 177 138 178 139
rect 176 138 177 139
rect 175 138 176 139
rect 174 138 175 139
rect 173 138 174 139
rect 172 138 173 139
rect 171 138 172 139
rect 170 138 171 139
rect 169 138 170 139
rect 168 138 169 139
rect 167 138 168 139
rect 166 138 167 139
rect 165 138 166 139
rect 164 138 165 139
rect 163 138 164 139
rect 162 138 163 139
rect 161 138 162 139
rect 73 138 74 139
rect 72 138 73 139
rect 71 138 72 139
rect 70 138 71 139
rect 69 138 70 139
rect 68 138 69 139
rect 67 138 68 139
rect 66 138 67 139
rect 65 138 66 139
rect 64 138 65 139
rect 63 138 64 139
rect 62 138 63 139
rect 61 138 62 139
rect 60 138 61 139
rect 59 138 60 139
rect 58 138 59 139
rect 57 138 58 139
rect 56 138 57 139
rect 55 138 56 139
rect 54 138 55 139
rect 53 138 54 139
rect 52 138 53 139
rect 51 138 52 139
rect 50 138 51 139
rect 49 138 50 139
rect 48 138 49 139
rect 47 138 48 139
rect 39 138 40 139
rect 38 138 39 139
rect 37 138 38 139
rect 36 138 37 139
rect 35 138 36 139
rect 34 138 35 139
rect 33 138 34 139
rect 32 138 33 139
rect 31 138 32 139
rect 30 138 31 139
rect 29 138 30 139
rect 28 138 29 139
rect 27 138 28 139
rect 26 138 27 139
rect 25 138 26 139
rect 20 138 21 139
rect 19 138 20 139
rect 18 138 19 139
rect 17 138 18 139
rect 16 138 17 139
rect 178 139 179 140
rect 177 139 178 140
rect 176 139 177 140
rect 175 139 176 140
rect 174 139 175 140
rect 173 139 174 140
rect 172 139 173 140
rect 171 139 172 140
rect 170 139 171 140
rect 169 139 170 140
rect 168 139 169 140
rect 167 139 168 140
rect 166 139 167 140
rect 165 139 166 140
rect 164 139 165 140
rect 163 139 164 140
rect 162 139 163 140
rect 161 139 162 140
rect 72 139 73 140
rect 71 139 72 140
rect 70 139 71 140
rect 69 139 70 140
rect 68 139 69 140
rect 67 139 68 140
rect 66 139 67 140
rect 65 139 66 140
rect 64 139 65 140
rect 63 139 64 140
rect 62 139 63 140
rect 61 139 62 140
rect 60 139 61 140
rect 59 139 60 140
rect 58 139 59 140
rect 57 139 58 140
rect 56 139 57 140
rect 55 139 56 140
rect 54 139 55 140
rect 53 139 54 140
rect 52 139 53 140
rect 51 139 52 140
rect 50 139 51 140
rect 49 139 50 140
rect 48 139 49 140
rect 39 139 40 140
rect 38 139 39 140
rect 37 139 38 140
rect 36 139 37 140
rect 35 139 36 140
rect 34 139 35 140
rect 33 139 34 140
rect 32 139 33 140
rect 31 139 32 140
rect 30 139 31 140
rect 29 139 30 140
rect 28 139 29 140
rect 27 139 28 140
rect 26 139 27 140
rect 25 139 26 140
rect 20 139 21 140
rect 19 139 20 140
rect 18 139 19 140
rect 17 139 18 140
rect 178 140 179 141
rect 177 140 178 141
rect 176 140 177 141
rect 175 140 176 141
rect 174 140 175 141
rect 173 140 174 141
rect 172 140 173 141
rect 171 140 172 141
rect 170 140 171 141
rect 169 140 170 141
rect 168 140 169 141
rect 167 140 168 141
rect 166 140 167 141
rect 165 140 166 141
rect 164 140 165 141
rect 163 140 164 141
rect 162 140 163 141
rect 161 140 162 141
rect 70 140 71 141
rect 69 140 70 141
rect 68 140 69 141
rect 67 140 68 141
rect 66 140 67 141
rect 65 140 66 141
rect 64 140 65 141
rect 63 140 64 141
rect 62 140 63 141
rect 61 140 62 141
rect 60 140 61 141
rect 59 140 60 141
rect 58 140 59 141
rect 57 140 58 141
rect 56 140 57 141
rect 55 140 56 141
rect 54 140 55 141
rect 53 140 54 141
rect 52 140 53 141
rect 51 140 52 141
rect 50 140 51 141
rect 49 140 50 141
rect 40 140 41 141
rect 39 140 40 141
rect 38 140 39 141
rect 37 140 38 141
rect 36 140 37 141
rect 35 140 36 141
rect 34 140 35 141
rect 33 140 34 141
rect 32 140 33 141
rect 31 140 32 141
rect 30 140 31 141
rect 29 140 30 141
rect 28 140 29 141
rect 27 140 28 141
rect 26 140 27 141
rect 25 140 26 141
rect 21 140 22 141
rect 20 140 21 141
rect 19 140 20 141
rect 18 140 19 141
rect 178 141 179 142
rect 177 141 178 142
rect 176 141 177 142
rect 175 141 176 142
rect 174 141 175 142
rect 173 141 174 142
rect 172 141 173 142
rect 171 141 172 142
rect 170 141 171 142
rect 169 141 170 142
rect 168 141 169 142
rect 167 141 168 142
rect 166 141 167 142
rect 165 141 166 142
rect 164 141 165 142
rect 163 141 164 142
rect 162 141 163 142
rect 161 141 162 142
rect 68 141 69 142
rect 67 141 68 142
rect 66 141 67 142
rect 65 141 66 142
rect 64 141 65 142
rect 63 141 64 142
rect 62 141 63 142
rect 61 141 62 142
rect 60 141 61 142
rect 59 141 60 142
rect 58 141 59 142
rect 57 141 58 142
rect 56 141 57 142
rect 55 141 56 142
rect 54 141 55 142
rect 53 141 54 142
rect 52 141 53 142
rect 51 141 52 142
rect 41 141 42 142
rect 40 141 41 142
rect 39 141 40 142
rect 38 141 39 142
rect 37 141 38 142
rect 36 141 37 142
rect 35 141 36 142
rect 34 141 35 142
rect 33 141 34 142
rect 32 141 33 142
rect 31 141 32 142
rect 30 141 31 142
rect 29 141 30 142
rect 28 141 29 142
rect 27 141 28 142
rect 26 141 27 142
rect 21 141 22 142
rect 178 142 179 143
rect 177 142 178 143
rect 170 142 171 143
rect 169 142 170 143
rect 168 142 169 143
rect 162 142 163 143
rect 161 142 162 143
rect 63 142 64 143
rect 62 142 63 143
rect 61 142 62 143
rect 60 142 61 143
rect 59 142 60 143
rect 58 142 59 143
rect 57 142 58 143
rect 56 142 57 143
rect 55 142 56 143
rect 54 142 55 143
rect 42 142 43 143
rect 41 142 42 143
rect 40 142 41 143
rect 39 142 40 143
rect 38 142 39 143
rect 37 142 38 143
rect 36 142 37 143
rect 35 142 36 143
rect 34 142 35 143
rect 33 142 34 143
rect 32 142 33 143
rect 31 142 32 143
rect 30 142 31 143
rect 29 142 30 143
rect 28 142 29 143
rect 27 142 28 143
rect 26 142 27 143
rect 178 143 179 144
rect 170 143 171 144
rect 169 143 170 144
rect 161 143 162 144
rect 43 143 44 144
rect 42 143 43 144
rect 41 143 42 144
rect 40 143 41 144
rect 39 143 40 144
rect 38 143 39 144
rect 37 143 38 144
rect 36 143 37 144
rect 35 143 36 144
rect 34 143 35 144
rect 33 143 34 144
rect 32 143 33 144
rect 31 143 32 144
rect 30 143 31 144
rect 29 143 30 144
rect 28 143 29 144
rect 27 143 28 144
rect 178 144 179 145
rect 170 144 171 145
rect 169 144 170 145
rect 161 144 162 145
rect 45 144 46 145
rect 44 144 45 145
rect 43 144 44 145
rect 42 144 43 145
rect 41 144 42 145
rect 40 144 41 145
rect 39 144 40 145
rect 38 144 39 145
rect 37 144 38 145
rect 36 144 37 145
rect 35 144 36 145
rect 34 144 35 145
rect 33 144 34 145
rect 32 144 33 145
rect 31 144 32 145
rect 30 144 31 145
rect 29 144 30 145
rect 28 144 29 145
rect 178 145 179 146
rect 170 145 171 146
rect 169 145 170 146
rect 161 145 162 146
rect 46 145 47 146
rect 45 145 46 146
rect 44 145 45 146
rect 43 145 44 146
rect 42 145 43 146
rect 41 145 42 146
rect 40 145 41 146
rect 39 145 40 146
rect 38 145 39 146
rect 37 145 38 146
rect 36 145 37 146
rect 35 145 36 146
rect 34 145 35 146
rect 33 145 34 146
rect 32 145 33 146
rect 31 145 32 146
rect 30 145 31 146
rect 29 145 30 146
rect 178 146 179 147
rect 171 146 172 147
rect 170 146 171 147
rect 169 146 170 147
rect 168 146 169 147
rect 162 146 163 147
rect 161 146 162 147
rect 48 146 49 147
rect 47 146 48 147
rect 46 146 47 147
rect 45 146 46 147
rect 44 146 45 147
rect 43 146 44 147
rect 42 146 43 147
rect 41 146 42 147
rect 40 146 41 147
rect 39 146 40 147
rect 38 146 39 147
rect 37 146 38 147
rect 36 146 37 147
rect 35 146 36 147
rect 34 146 35 147
rect 33 146 34 147
rect 32 146 33 147
rect 31 146 32 147
rect 30 146 31 147
rect 178 147 179 148
rect 177 147 178 148
rect 172 147 173 148
rect 171 147 172 148
rect 170 147 171 148
rect 169 147 170 148
rect 168 147 169 148
rect 167 147 168 148
rect 162 147 163 148
rect 161 147 162 148
rect 49 147 50 148
rect 48 147 49 148
rect 47 147 48 148
rect 46 147 47 148
rect 45 147 46 148
rect 44 147 45 148
rect 43 147 44 148
rect 42 147 43 148
rect 41 147 42 148
rect 40 147 41 148
rect 39 147 40 148
rect 38 147 39 148
rect 37 147 38 148
rect 36 147 37 148
rect 35 147 36 148
rect 34 147 35 148
rect 33 147 34 148
rect 32 147 33 148
rect 178 148 179 149
rect 177 148 178 149
rect 176 148 177 149
rect 165 148 166 149
rect 164 148 165 149
rect 163 148 164 149
rect 162 148 163 149
rect 161 148 162 149
rect 49 148 50 149
rect 48 148 49 149
rect 47 148 48 149
rect 46 148 47 149
rect 45 148 46 149
rect 44 148 45 149
rect 43 148 44 149
rect 42 148 43 149
rect 41 148 42 149
rect 40 148 41 149
rect 39 148 40 149
rect 38 148 39 149
rect 37 148 38 149
rect 36 148 37 149
rect 35 148 36 149
rect 178 149 179 150
rect 177 149 178 150
rect 176 149 177 150
rect 175 149 176 150
rect 174 149 175 150
rect 164 149 165 150
rect 163 149 164 150
rect 162 149 163 150
rect 45 149 46 150
rect 44 149 45 150
rect 43 149 44 150
rect 42 149 43 150
rect 41 149 42 150
rect 40 149 41 150
rect 176 150 177 151
rect 175 150 176 151
rect 174 150 175 151
rect 178 153 179 154
rect 161 153 162 154
rect 178 154 179 155
rect 161 154 162 155
rect 178 155 179 156
rect 177 155 178 156
rect 176 155 177 156
rect 175 155 176 156
rect 174 155 175 156
rect 173 155 174 156
rect 172 155 173 156
rect 171 155 172 156
rect 170 155 171 156
rect 169 155 170 156
rect 168 155 169 156
rect 167 155 168 156
rect 166 155 167 156
rect 165 155 166 156
rect 164 155 165 156
rect 163 155 164 156
rect 162 155 163 156
rect 161 155 162 156
rect 178 156 179 157
rect 177 156 178 157
rect 176 156 177 157
rect 175 156 176 157
rect 174 156 175 157
rect 173 156 174 157
rect 172 156 173 157
rect 171 156 172 157
rect 170 156 171 157
rect 169 156 170 157
rect 168 156 169 157
rect 167 156 168 157
rect 166 156 167 157
rect 165 156 166 157
rect 164 156 165 157
rect 163 156 164 157
rect 162 156 163 157
rect 161 156 162 157
rect 178 157 179 158
rect 177 157 178 158
rect 176 157 177 158
rect 175 157 176 158
rect 174 157 175 158
rect 173 157 174 158
rect 172 157 173 158
rect 171 157 172 158
rect 170 157 171 158
rect 169 157 170 158
rect 168 157 169 158
rect 167 157 168 158
rect 166 157 167 158
rect 165 157 166 158
rect 164 157 165 158
rect 163 157 164 158
rect 162 157 163 158
rect 161 157 162 158
rect 178 158 179 159
rect 177 158 178 159
rect 176 158 177 159
rect 175 158 176 159
rect 174 158 175 159
rect 173 158 174 159
rect 172 158 173 159
rect 171 158 172 159
rect 170 158 171 159
rect 169 158 170 159
rect 168 158 169 159
rect 167 158 168 159
rect 166 158 167 159
rect 165 158 166 159
rect 164 158 165 159
rect 163 158 164 159
rect 162 158 163 159
rect 161 158 162 159
rect 178 159 179 160
rect 177 159 178 160
rect 176 159 177 160
rect 175 159 176 160
rect 174 159 175 160
rect 173 159 174 160
rect 172 159 173 160
rect 171 159 172 160
rect 170 159 171 160
rect 169 159 170 160
rect 168 159 169 160
rect 167 159 168 160
rect 166 159 167 160
rect 165 159 166 160
rect 164 159 165 160
rect 163 159 164 160
rect 162 159 163 160
rect 161 159 162 160
rect 178 160 179 161
rect 177 160 178 161
rect 170 160 171 161
rect 169 160 170 161
rect 161 160 162 161
rect 178 161 179 162
rect 170 161 171 162
rect 169 161 170 162
rect 161 161 162 162
rect 178 162 179 163
rect 170 162 171 163
rect 169 162 170 163
rect 161 162 162 163
rect 178 163 179 164
rect 170 163 171 164
rect 169 163 170 164
rect 168 163 169 164
rect 162 163 163 164
rect 161 163 162 164
rect 178 164 179 165
rect 177 164 178 165
rect 172 164 173 165
rect 171 164 172 165
rect 170 164 171 165
rect 169 164 170 165
rect 168 164 169 165
rect 167 164 168 165
rect 162 164 163 165
rect 161 164 162 165
rect 178 165 179 166
rect 177 165 178 166
rect 176 165 177 166
rect 171 165 172 166
rect 170 165 171 166
rect 169 165 170 166
rect 168 165 169 166
rect 167 165 168 166
rect 164 165 165 166
rect 163 165 164 166
rect 162 165 163 166
rect 161 165 162 166
rect 178 166 179 167
rect 177 166 178 167
rect 176 166 177 167
rect 175 166 176 167
rect 164 166 165 167
rect 163 166 164 167
rect 162 166 163 167
rect 161 166 162 167
rect 177 167 178 168
rect 176 167 177 168
rect 175 167 176 168
rect 174 167 175 168
rect 141 174 142 175
rect 140 174 141 175
rect 139 174 140 175
rect 138 174 139 175
rect 137 174 138 175
rect 136 174 137 175
rect 135 174 136 175
rect 134 174 135 175
rect 133 174 134 175
rect 132 174 133 175
rect 131 174 132 175
rect 130 174 131 175
rect 129 174 130 175
rect 128 174 129 175
rect 127 174 128 175
rect 126 174 127 175
rect 125 174 126 175
rect 124 174 125 175
rect 123 174 124 175
rect 122 174 123 175
rect 121 174 122 175
rect 120 174 121 175
rect 119 174 120 175
rect 118 174 119 175
rect 117 174 118 175
rect 116 174 117 175
rect 115 174 116 175
rect 114 174 115 175
rect 113 174 114 175
rect 112 174 113 175
rect 111 174 112 175
rect 110 174 111 175
rect 109 174 110 175
rect 108 174 109 175
rect 107 174 108 175
rect 106 174 107 175
rect 105 174 106 175
rect 104 174 105 175
rect 103 174 104 175
rect 102 174 103 175
rect 101 174 102 175
rect 100 174 101 175
rect 143 175 144 176
rect 142 175 143 176
rect 141 175 142 176
rect 140 175 141 176
rect 139 175 140 176
rect 138 175 139 176
rect 137 175 138 176
rect 136 175 137 176
rect 135 175 136 176
rect 134 175 135 176
rect 133 175 134 176
rect 132 175 133 176
rect 131 175 132 176
rect 130 175 131 176
rect 129 175 130 176
rect 128 175 129 176
rect 127 175 128 176
rect 126 175 127 176
rect 125 175 126 176
rect 124 175 125 176
rect 123 175 124 176
rect 122 175 123 176
rect 121 175 122 176
rect 120 175 121 176
rect 119 175 120 176
rect 118 175 119 176
rect 117 175 118 176
rect 116 175 117 176
rect 115 175 116 176
rect 114 175 115 176
rect 113 175 114 176
rect 112 175 113 176
rect 111 175 112 176
rect 110 175 111 176
rect 109 175 110 176
rect 108 175 109 176
rect 107 175 108 176
rect 106 175 107 176
rect 105 175 106 176
rect 104 175 105 176
rect 103 175 104 176
rect 102 175 103 176
rect 101 175 102 176
rect 100 175 101 176
rect 194 176 195 177
rect 193 176 194 177
rect 192 176 193 177
rect 191 176 192 177
rect 190 176 191 177
rect 189 176 190 177
rect 188 176 189 177
rect 187 176 188 177
rect 170 176 171 177
rect 165 176 166 177
rect 164 176 165 177
rect 163 176 164 177
rect 144 176 145 177
rect 143 176 144 177
rect 142 176 143 177
rect 141 176 142 177
rect 140 176 141 177
rect 139 176 140 177
rect 138 176 139 177
rect 137 176 138 177
rect 136 176 137 177
rect 135 176 136 177
rect 134 176 135 177
rect 133 176 134 177
rect 132 176 133 177
rect 131 176 132 177
rect 130 176 131 177
rect 129 176 130 177
rect 128 176 129 177
rect 127 176 128 177
rect 126 176 127 177
rect 125 176 126 177
rect 124 176 125 177
rect 123 176 124 177
rect 122 176 123 177
rect 121 176 122 177
rect 120 176 121 177
rect 119 176 120 177
rect 118 176 119 177
rect 117 176 118 177
rect 116 176 117 177
rect 115 176 116 177
rect 114 176 115 177
rect 113 176 114 177
rect 112 176 113 177
rect 111 176 112 177
rect 110 176 111 177
rect 109 176 110 177
rect 108 176 109 177
rect 107 176 108 177
rect 106 176 107 177
rect 105 176 106 177
rect 104 176 105 177
rect 103 176 104 177
rect 102 176 103 177
rect 101 176 102 177
rect 100 176 101 177
rect 195 177 196 178
rect 194 177 195 178
rect 193 177 194 178
rect 192 177 193 178
rect 191 177 192 178
rect 190 177 191 178
rect 189 177 190 178
rect 188 177 189 178
rect 187 177 188 178
rect 172 177 173 178
rect 171 177 172 178
rect 170 177 171 178
rect 169 177 170 178
rect 168 177 169 178
rect 165 177 166 178
rect 164 177 165 178
rect 163 177 164 178
rect 145 177 146 178
rect 144 177 145 178
rect 143 177 144 178
rect 142 177 143 178
rect 141 177 142 178
rect 140 177 141 178
rect 139 177 140 178
rect 138 177 139 178
rect 137 177 138 178
rect 136 177 137 178
rect 135 177 136 178
rect 134 177 135 178
rect 133 177 134 178
rect 132 177 133 178
rect 131 177 132 178
rect 130 177 131 178
rect 129 177 130 178
rect 128 177 129 178
rect 127 177 128 178
rect 126 177 127 178
rect 125 177 126 178
rect 124 177 125 178
rect 123 177 124 178
rect 122 177 123 178
rect 121 177 122 178
rect 120 177 121 178
rect 119 177 120 178
rect 118 177 119 178
rect 117 177 118 178
rect 116 177 117 178
rect 115 177 116 178
rect 114 177 115 178
rect 113 177 114 178
rect 112 177 113 178
rect 111 177 112 178
rect 110 177 111 178
rect 109 177 110 178
rect 108 177 109 178
rect 107 177 108 178
rect 106 177 107 178
rect 105 177 106 178
rect 104 177 105 178
rect 103 177 104 178
rect 102 177 103 178
rect 101 177 102 178
rect 100 177 101 178
rect 194 178 195 179
rect 193 178 194 179
rect 192 178 193 179
rect 191 178 192 179
rect 190 178 191 179
rect 189 178 190 179
rect 188 178 189 179
rect 187 178 188 179
rect 172 178 173 179
rect 171 178 172 179
rect 170 178 171 179
rect 169 178 170 179
rect 168 178 169 179
rect 167 178 168 179
rect 165 178 166 179
rect 164 178 165 179
rect 163 178 164 179
rect 146 178 147 179
rect 145 178 146 179
rect 144 178 145 179
rect 143 178 144 179
rect 142 178 143 179
rect 141 178 142 179
rect 140 178 141 179
rect 139 178 140 179
rect 138 178 139 179
rect 137 178 138 179
rect 136 178 137 179
rect 135 178 136 179
rect 134 178 135 179
rect 133 178 134 179
rect 132 178 133 179
rect 131 178 132 179
rect 130 178 131 179
rect 129 178 130 179
rect 128 178 129 179
rect 127 178 128 179
rect 126 178 127 179
rect 125 178 126 179
rect 124 178 125 179
rect 123 178 124 179
rect 122 178 123 179
rect 121 178 122 179
rect 120 178 121 179
rect 119 178 120 179
rect 118 178 119 179
rect 117 178 118 179
rect 116 178 117 179
rect 115 178 116 179
rect 114 178 115 179
rect 113 178 114 179
rect 112 178 113 179
rect 111 178 112 179
rect 110 178 111 179
rect 109 178 110 179
rect 108 178 109 179
rect 107 178 108 179
rect 106 178 107 179
rect 105 178 106 179
rect 104 178 105 179
rect 103 178 104 179
rect 102 178 103 179
rect 101 178 102 179
rect 100 178 101 179
rect 194 179 195 180
rect 191 179 192 180
rect 190 179 191 180
rect 187 179 188 180
rect 180 179 181 180
rect 179 179 180 180
rect 178 179 179 180
rect 177 179 178 180
rect 176 179 177 180
rect 173 179 174 180
rect 172 179 173 180
rect 171 179 172 180
rect 170 179 171 180
rect 169 179 170 180
rect 168 179 169 180
rect 167 179 168 180
rect 165 179 166 180
rect 164 179 165 180
rect 163 179 164 180
rect 161 179 162 180
rect 160 179 161 180
rect 146 179 147 180
rect 145 179 146 180
rect 144 179 145 180
rect 143 179 144 180
rect 142 179 143 180
rect 141 179 142 180
rect 140 179 141 180
rect 139 179 140 180
rect 138 179 139 180
rect 137 179 138 180
rect 136 179 137 180
rect 135 179 136 180
rect 134 179 135 180
rect 133 179 134 180
rect 132 179 133 180
rect 131 179 132 180
rect 130 179 131 180
rect 129 179 130 180
rect 128 179 129 180
rect 127 179 128 180
rect 126 179 127 180
rect 125 179 126 180
rect 124 179 125 180
rect 123 179 124 180
rect 122 179 123 180
rect 121 179 122 180
rect 120 179 121 180
rect 119 179 120 180
rect 118 179 119 180
rect 117 179 118 180
rect 116 179 117 180
rect 115 179 116 180
rect 114 179 115 180
rect 113 179 114 180
rect 112 179 113 180
rect 111 179 112 180
rect 110 179 111 180
rect 109 179 110 180
rect 108 179 109 180
rect 107 179 108 180
rect 106 179 107 180
rect 105 179 106 180
rect 104 179 105 180
rect 103 179 104 180
rect 102 179 103 180
rect 101 179 102 180
rect 100 179 101 180
rect 194 180 195 181
rect 191 180 192 181
rect 190 180 191 181
rect 187 180 188 181
rect 181 180 182 181
rect 180 180 181 181
rect 179 180 180 181
rect 178 180 179 181
rect 177 180 178 181
rect 176 180 177 181
rect 175 180 176 181
rect 173 180 174 181
rect 172 180 173 181
rect 171 180 172 181
rect 170 180 171 181
rect 169 180 170 181
rect 168 180 169 181
rect 167 180 168 181
rect 165 180 166 181
rect 164 180 165 181
rect 163 180 164 181
rect 161 180 162 181
rect 160 180 161 181
rect 147 180 148 181
rect 146 180 147 181
rect 145 180 146 181
rect 144 180 145 181
rect 143 180 144 181
rect 142 180 143 181
rect 141 180 142 181
rect 140 180 141 181
rect 139 180 140 181
rect 138 180 139 181
rect 137 180 138 181
rect 136 180 137 181
rect 135 180 136 181
rect 134 180 135 181
rect 133 180 134 181
rect 132 180 133 181
rect 131 180 132 181
rect 130 180 131 181
rect 129 180 130 181
rect 128 180 129 181
rect 127 180 128 181
rect 126 180 127 181
rect 125 180 126 181
rect 124 180 125 181
rect 123 180 124 181
rect 122 180 123 181
rect 121 180 122 181
rect 120 180 121 181
rect 119 180 120 181
rect 118 180 119 181
rect 117 180 118 181
rect 116 180 117 181
rect 115 180 116 181
rect 114 180 115 181
rect 113 180 114 181
rect 112 180 113 181
rect 111 180 112 181
rect 110 180 111 181
rect 109 180 110 181
rect 108 180 109 181
rect 107 180 108 181
rect 106 180 107 181
rect 105 180 106 181
rect 104 180 105 181
rect 103 180 104 181
rect 102 180 103 181
rect 101 180 102 181
rect 100 180 101 181
rect 60 180 61 181
rect 59 180 60 181
rect 58 180 59 181
rect 57 180 58 181
rect 195 181 196 182
rect 194 181 195 182
rect 191 181 192 182
rect 190 181 191 182
rect 187 181 188 182
rect 181 181 182 182
rect 180 181 181 182
rect 179 181 180 182
rect 178 181 179 182
rect 177 181 178 182
rect 176 181 177 182
rect 175 181 176 182
rect 173 181 174 182
rect 172 181 173 182
rect 171 181 172 182
rect 169 181 170 182
rect 168 181 169 182
rect 167 181 168 182
rect 166 181 167 182
rect 165 181 166 182
rect 164 181 165 182
rect 163 181 164 182
rect 161 181 162 182
rect 160 181 161 182
rect 147 181 148 182
rect 146 181 147 182
rect 145 181 146 182
rect 144 181 145 182
rect 143 181 144 182
rect 142 181 143 182
rect 141 181 142 182
rect 140 181 141 182
rect 139 181 140 182
rect 138 181 139 182
rect 137 181 138 182
rect 136 181 137 182
rect 135 181 136 182
rect 134 181 135 182
rect 133 181 134 182
rect 132 181 133 182
rect 131 181 132 182
rect 130 181 131 182
rect 129 181 130 182
rect 128 181 129 182
rect 127 181 128 182
rect 126 181 127 182
rect 125 181 126 182
rect 124 181 125 182
rect 123 181 124 182
rect 122 181 123 182
rect 121 181 122 182
rect 120 181 121 182
rect 119 181 120 182
rect 118 181 119 182
rect 117 181 118 182
rect 116 181 117 182
rect 115 181 116 182
rect 114 181 115 182
rect 113 181 114 182
rect 112 181 113 182
rect 111 181 112 182
rect 110 181 111 182
rect 109 181 110 182
rect 108 181 109 182
rect 107 181 108 182
rect 106 181 107 182
rect 105 181 106 182
rect 104 181 105 182
rect 103 181 104 182
rect 102 181 103 182
rect 101 181 102 182
rect 100 181 101 182
rect 60 181 61 182
rect 59 181 60 182
rect 58 181 59 182
rect 57 181 58 182
rect 27 181 28 182
rect 26 181 27 182
rect 181 182 182 183
rect 180 182 181 183
rect 179 182 180 183
rect 178 182 179 183
rect 177 182 178 183
rect 176 182 177 183
rect 175 182 176 183
rect 173 182 174 183
rect 172 182 173 183
rect 168 182 169 183
rect 167 182 168 183
rect 166 182 167 183
rect 165 182 166 183
rect 164 182 165 183
rect 163 182 164 183
rect 161 182 162 183
rect 160 182 161 183
rect 147 182 148 183
rect 146 182 147 183
rect 145 182 146 183
rect 144 182 145 183
rect 143 182 144 183
rect 142 182 143 183
rect 141 182 142 183
rect 140 182 141 183
rect 139 182 140 183
rect 138 182 139 183
rect 137 182 138 183
rect 136 182 137 183
rect 135 182 136 183
rect 134 182 135 183
rect 133 182 134 183
rect 132 182 133 183
rect 131 182 132 183
rect 130 182 131 183
rect 129 182 130 183
rect 128 182 129 183
rect 127 182 128 183
rect 126 182 127 183
rect 125 182 126 183
rect 124 182 125 183
rect 123 182 124 183
rect 122 182 123 183
rect 121 182 122 183
rect 120 182 121 183
rect 119 182 120 183
rect 118 182 119 183
rect 117 182 118 183
rect 116 182 117 183
rect 115 182 116 183
rect 114 182 115 183
rect 113 182 114 183
rect 112 182 113 183
rect 111 182 112 183
rect 110 182 111 183
rect 109 182 110 183
rect 108 182 109 183
rect 107 182 108 183
rect 106 182 107 183
rect 105 182 106 183
rect 104 182 105 183
rect 103 182 104 183
rect 102 182 103 183
rect 101 182 102 183
rect 100 182 101 183
rect 60 182 61 183
rect 59 182 60 183
rect 58 182 59 183
rect 57 182 58 183
rect 27 182 28 183
rect 26 182 27 183
rect 25 182 26 183
rect 24 182 25 183
rect 16 182 17 183
rect 194 183 195 184
rect 193 183 194 184
rect 192 183 193 184
rect 191 183 192 184
rect 190 183 191 184
rect 189 183 190 184
rect 188 183 189 184
rect 187 183 188 184
rect 186 183 187 184
rect 181 183 182 184
rect 180 183 181 184
rect 179 183 180 184
rect 178 183 179 184
rect 177 183 178 184
rect 176 183 177 184
rect 173 183 174 184
rect 172 183 173 184
rect 168 183 169 184
rect 167 183 168 184
rect 166 183 167 184
rect 165 183 166 184
rect 164 183 165 184
rect 163 183 164 184
rect 161 183 162 184
rect 160 183 161 184
rect 147 183 148 184
rect 146 183 147 184
rect 145 183 146 184
rect 144 183 145 184
rect 143 183 144 184
rect 142 183 143 184
rect 141 183 142 184
rect 140 183 141 184
rect 139 183 140 184
rect 138 183 139 184
rect 137 183 138 184
rect 136 183 137 184
rect 135 183 136 184
rect 134 183 135 184
rect 133 183 134 184
rect 132 183 133 184
rect 131 183 132 184
rect 130 183 131 184
rect 129 183 130 184
rect 128 183 129 184
rect 127 183 128 184
rect 126 183 127 184
rect 125 183 126 184
rect 124 183 125 184
rect 123 183 124 184
rect 122 183 123 184
rect 121 183 122 184
rect 120 183 121 184
rect 119 183 120 184
rect 118 183 119 184
rect 117 183 118 184
rect 116 183 117 184
rect 115 183 116 184
rect 114 183 115 184
rect 113 183 114 184
rect 112 183 113 184
rect 111 183 112 184
rect 110 183 111 184
rect 109 183 110 184
rect 108 183 109 184
rect 107 183 108 184
rect 106 183 107 184
rect 105 183 106 184
rect 104 183 105 184
rect 103 183 104 184
rect 102 183 103 184
rect 101 183 102 184
rect 100 183 101 184
rect 76 183 77 184
rect 75 183 76 184
rect 74 183 75 184
rect 73 183 74 184
rect 72 183 73 184
rect 71 183 72 184
rect 70 183 71 184
rect 69 183 70 184
rect 68 183 69 184
rect 67 183 68 184
rect 66 183 67 184
rect 65 183 66 184
rect 64 183 65 184
rect 63 183 64 184
rect 62 183 63 184
rect 61 183 62 184
rect 60 183 61 184
rect 59 183 60 184
rect 58 183 59 184
rect 57 183 58 184
rect 56 183 57 184
rect 55 183 56 184
rect 54 183 55 184
rect 53 183 54 184
rect 52 183 53 184
rect 27 183 28 184
rect 26 183 27 184
rect 25 183 26 184
rect 24 183 25 184
rect 23 183 24 184
rect 17 183 18 184
rect 16 183 17 184
rect 15 183 16 184
rect 194 184 195 185
rect 193 184 194 185
rect 192 184 193 185
rect 191 184 192 185
rect 190 184 191 185
rect 189 184 190 185
rect 188 184 189 185
rect 187 184 188 185
rect 186 184 187 185
rect 181 184 182 185
rect 180 184 181 185
rect 179 184 180 185
rect 178 184 179 185
rect 173 184 174 185
rect 172 184 173 185
rect 168 184 169 185
rect 167 184 168 185
rect 166 184 167 185
rect 165 184 166 185
rect 164 184 165 185
rect 163 184 164 185
rect 161 184 162 185
rect 160 184 161 185
rect 147 184 148 185
rect 146 184 147 185
rect 145 184 146 185
rect 144 184 145 185
rect 143 184 144 185
rect 142 184 143 185
rect 141 184 142 185
rect 140 184 141 185
rect 139 184 140 185
rect 138 184 139 185
rect 137 184 138 185
rect 136 184 137 185
rect 135 184 136 185
rect 134 184 135 185
rect 133 184 134 185
rect 132 184 133 185
rect 131 184 132 185
rect 130 184 131 185
rect 129 184 130 185
rect 128 184 129 185
rect 127 184 128 185
rect 126 184 127 185
rect 125 184 126 185
rect 124 184 125 185
rect 123 184 124 185
rect 122 184 123 185
rect 121 184 122 185
rect 120 184 121 185
rect 119 184 120 185
rect 118 184 119 185
rect 117 184 118 185
rect 116 184 117 185
rect 115 184 116 185
rect 114 184 115 185
rect 113 184 114 185
rect 112 184 113 185
rect 111 184 112 185
rect 110 184 111 185
rect 109 184 110 185
rect 108 184 109 185
rect 107 184 108 185
rect 106 184 107 185
rect 105 184 106 185
rect 104 184 105 185
rect 103 184 104 185
rect 102 184 103 185
rect 101 184 102 185
rect 100 184 101 185
rect 76 184 77 185
rect 75 184 76 185
rect 74 184 75 185
rect 73 184 74 185
rect 72 184 73 185
rect 71 184 72 185
rect 70 184 71 185
rect 69 184 70 185
rect 68 184 69 185
rect 67 184 68 185
rect 66 184 67 185
rect 65 184 66 185
rect 64 184 65 185
rect 63 184 64 185
rect 62 184 63 185
rect 61 184 62 185
rect 60 184 61 185
rect 59 184 60 185
rect 58 184 59 185
rect 57 184 58 185
rect 56 184 57 185
rect 55 184 56 185
rect 54 184 55 185
rect 53 184 54 185
rect 52 184 53 185
rect 51 184 52 185
rect 50 184 51 185
rect 27 184 28 185
rect 26 184 27 185
rect 25 184 26 185
rect 24 184 25 185
rect 23 184 24 185
rect 22 184 23 185
rect 17 184 18 185
rect 16 184 17 185
rect 15 184 16 185
rect 14 184 15 185
rect 181 185 182 186
rect 180 185 181 186
rect 179 185 180 186
rect 178 185 179 186
rect 173 185 174 186
rect 172 185 173 186
rect 171 185 172 186
rect 169 185 170 186
rect 168 185 169 186
rect 167 185 168 186
rect 166 185 167 186
rect 165 185 166 186
rect 164 185 165 186
rect 163 185 164 186
rect 161 185 162 186
rect 160 185 161 186
rect 147 185 148 186
rect 146 185 147 186
rect 145 185 146 186
rect 144 185 145 186
rect 143 185 144 186
rect 142 185 143 186
rect 141 185 142 186
rect 140 185 141 186
rect 139 185 140 186
rect 138 185 139 186
rect 137 185 138 186
rect 136 185 137 186
rect 135 185 136 186
rect 134 185 135 186
rect 133 185 134 186
rect 132 185 133 186
rect 131 185 132 186
rect 130 185 131 186
rect 129 185 130 186
rect 128 185 129 186
rect 127 185 128 186
rect 126 185 127 186
rect 125 185 126 186
rect 124 185 125 186
rect 123 185 124 186
rect 122 185 123 186
rect 121 185 122 186
rect 120 185 121 186
rect 119 185 120 186
rect 118 185 119 186
rect 117 185 118 186
rect 116 185 117 186
rect 115 185 116 186
rect 114 185 115 186
rect 113 185 114 186
rect 112 185 113 186
rect 111 185 112 186
rect 110 185 111 186
rect 109 185 110 186
rect 108 185 109 186
rect 107 185 108 186
rect 106 185 107 186
rect 105 185 106 186
rect 104 185 105 186
rect 103 185 104 186
rect 102 185 103 186
rect 101 185 102 186
rect 100 185 101 186
rect 76 185 77 186
rect 75 185 76 186
rect 74 185 75 186
rect 73 185 74 186
rect 72 185 73 186
rect 71 185 72 186
rect 70 185 71 186
rect 69 185 70 186
rect 68 185 69 186
rect 67 185 68 186
rect 66 185 67 186
rect 65 185 66 186
rect 64 185 65 186
rect 63 185 64 186
rect 62 185 63 186
rect 61 185 62 186
rect 60 185 61 186
rect 59 185 60 186
rect 58 185 59 186
rect 57 185 58 186
rect 56 185 57 186
rect 55 185 56 186
rect 54 185 55 186
rect 53 185 54 186
rect 52 185 53 186
rect 51 185 52 186
rect 50 185 51 186
rect 27 185 28 186
rect 26 185 27 186
rect 25 185 26 186
rect 24 185 25 186
rect 23 185 24 186
rect 22 185 23 186
rect 21 185 22 186
rect 17 185 18 186
rect 16 185 17 186
rect 15 185 16 186
rect 14 185 15 186
rect 13 185 14 186
rect 194 186 195 187
rect 193 186 194 187
rect 192 186 193 187
rect 191 186 192 187
rect 190 186 191 187
rect 181 186 182 187
rect 180 186 181 187
rect 179 186 180 187
rect 178 186 179 187
rect 173 186 174 187
rect 172 186 173 187
rect 171 186 172 187
rect 169 186 170 187
rect 168 186 169 187
rect 167 186 168 187
rect 166 186 167 187
rect 165 186 166 187
rect 164 186 165 187
rect 163 186 164 187
rect 161 186 162 187
rect 160 186 161 187
rect 147 186 148 187
rect 146 186 147 187
rect 145 186 146 187
rect 144 186 145 187
rect 143 186 144 187
rect 142 186 143 187
rect 141 186 142 187
rect 140 186 141 187
rect 139 186 140 187
rect 138 186 139 187
rect 137 186 138 187
rect 136 186 137 187
rect 135 186 136 187
rect 134 186 135 187
rect 133 186 134 187
rect 132 186 133 187
rect 131 186 132 187
rect 130 186 131 187
rect 129 186 130 187
rect 128 186 129 187
rect 127 186 128 187
rect 126 186 127 187
rect 125 186 126 187
rect 124 186 125 187
rect 123 186 124 187
rect 122 186 123 187
rect 121 186 122 187
rect 120 186 121 187
rect 119 186 120 187
rect 118 186 119 187
rect 117 186 118 187
rect 116 186 117 187
rect 115 186 116 187
rect 114 186 115 187
rect 113 186 114 187
rect 112 186 113 187
rect 111 186 112 187
rect 110 186 111 187
rect 109 186 110 187
rect 108 186 109 187
rect 107 186 108 187
rect 106 186 107 187
rect 105 186 106 187
rect 104 186 105 187
rect 103 186 104 187
rect 102 186 103 187
rect 101 186 102 187
rect 100 186 101 187
rect 76 186 77 187
rect 75 186 76 187
rect 74 186 75 187
rect 73 186 74 187
rect 72 186 73 187
rect 71 186 72 187
rect 70 186 71 187
rect 69 186 70 187
rect 68 186 69 187
rect 67 186 68 187
rect 66 186 67 187
rect 65 186 66 187
rect 64 186 65 187
rect 63 186 64 187
rect 62 186 63 187
rect 61 186 62 187
rect 60 186 61 187
rect 59 186 60 187
rect 58 186 59 187
rect 57 186 58 187
rect 56 186 57 187
rect 55 186 56 187
rect 54 186 55 187
rect 53 186 54 187
rect 52 186 53 187
rect 51 186 52 187
rect 50 186 51 187
rect 49 186 50 187
rect 27 186 28 187
rect 26 186 27 187
rect 25 186 26 187
rect 23 186 24 187
rect 22 186 23 187
rect 21 186 22 187
rect 20 186 21 187
rect 15 186 16 187
rect 14 186 15 187
rect 13 186 14 187
rect 194 187 195 188
rect 193 187 194 188
rect 192 187 193 188
rect 191 187 192 188
rect 190 187 191 188
rect 189 187 190 188
rect 181 187 182 188
rect 180 187 181 188
rect 179 187 180 188
rect 178 187 179 188
rect 173 187 174 188
rect 172 187 173 188
rect 171 187 172 188
rect 170 187 171 188
rect 169 187 170 188
rect 168 187 169 188
rect 167 187 168 188
rect 165 187 166 188
rect 164 187 165 188
rect 163 187 164 188
rect 161 187 162 188
rect 160 187 161 188
rect 147 187 148 188
rect 146 187 147 188
rect 145 187 146 188
rect 144 187 145 188
rect 143 187 144 188
rect 142 187 143 188
rect 141 187 142 188
rect 140 187 141 188
rect 139 187 140 188
rect 138 187 139 188
rect 137 187 138 188
rect 136 187 137 188
rect 135 187 136 188
rect 134 187 135 188
rect 133 187 134 188
rect 132 187 133 188
rect 131 187 132 188
rect 130 187 131 188
rect 129 187 130 188
rect 128 187 129 188
rect 127 187 128 188
rect 126 187 127 188
rect 125 187 126 188
rect 124 187 125 188
rect 123 187 124 188
rect 122 187 123 188
rect 121 187 122 188
rect 120 187 121 188
rect 119 187 120 188
rect 118 187 119 188
rect 117 187 118 188
rect 116 187 117 188
rect 115 187 116 188
rect 114 187 115 188
rect 113 187 114 188
rect 112 187 113 188
rect 111 187 112 188
rect 110 187 111 188
rect 109 187 110 188
rect 108 187 109 188
rect 107 187 108 188
rect 106 187 107 188
rect 105 187 106 188
rect 104 187 105 188
rect 103 187 104 188
rect 102 187 103 188
rect 101 187 102 188
rect 100 187 101 188
rect 76 187 77 188
rect 75 187 76 188
rect 74 187 75 188
rect 73 187 74 188
rect 72 187 73 188
rect 71 187 72 188
rect 70 187 71 188
rect 69 187 70 188
rect 68 187 69 188
rect 67 187 68 188
rect 66 187 67 188
rect 65 187 66 188
rect 64 187 65 188
rect 63 187 64 188
rect 62 187 63 188
rect 61 187 62 188
rect 60 187 61 188
rect 59 187 60 188
rect 58 187 59 188
rect 57 187 58 188
rect 56 187 57 188
rect 55 187 56 188
rect 54 187 55 188
rect 53 187 54 188
rect 52 187 53 188
rect 51 187 52 188
rect 50 187 51 188
rect 49 187 50 188
rect 27 187 28 188
rect 26 187 27 188
rect 25 187 26 188
rect 22 187 23 188
rect 21 187 22 188
rect 20 187 21 188
rect 19 187 20 188
rect 15 187 16 188
rect 14 187 15 188
rect 13 187 14 188
rect 195 188 196 189
rect 194 188 195 189
rect 192 188 193 189
rect 190 188 191 189
rect 189 188 190 189
rect 181 188 182 189
rect 180 188 181 189
rect 179 188 180 189
rect 178 188 179 189
rect 173 188 174 189
rect 172 188 173 189
rect 171 188 172 189
rect 170 188 171 189
rect 169 188 170 189
rect 168 188 169 189
rect 167 188 168 189
rect 165 188 166 189
rect 164 188 165 189
rect 163 188 164 189
rect 147 188 148 189
rect 146 188 147 189
rect 145 188 146 189
rect 144 188 145 189
rect 143 188 144 189
rect 142 188 143 189
rect 141 188 142 189
rect 140 188 141 189
rect 139 188 140 189
rect 138 188 139 189
rect 137 188 138 189
rect 136 188 137 189
rect 135 188 136 189
rect 134 188 135 189
rect 133 188 134 189
rect 132 188 133 189
rect 131 188 132 189
rect 130 188 131 189
rect 129 188 130 189
rect 128 188 129 189
rect 127 188 128 189
rect 126 188 127 189
rect 125 188 126 189
rect 124 188 125 189
rect 123 188 124 189
rect 122 188 123 189
rect 121 188 122 189
rect 120 188 121 189
rect 119 188 120 189
rect 118 188 119 189
rect 117 188 118 189
rect 116 188 117 189
rect 115 188 116 189
rect 114 188 115 189
rect 113 188 114 189
rect 112 188 113 189
rect 111 188 112 189
rect 110 188 111 189
rect 109 188 110 189
rect 108 188 109 189
rect 107 188 108 189
rect 106 188 107 189
rect 105 188 106 189
rect 104 188 105 189
rect 103 188 104 189
rect 102 188 103 189
rect 101 188 102 189
rect 100 188 101 189
rect 76 188 77 189
rect 75 188 76 189
rect 74 188 75 189
rect 73 188 74 189
rect 72 188 73 189
rect 71 188 72 189
rect 70 188 71 189
rect 69 188 70 189
rect 68 188 69 189
rect 67 188 68 189
rect 66 188 67 189
rect 65 188 66 189
rect 64 188 65 189
rect 63 188 64 189
rect 62 188 63 189
rect 61 188 62 189
rect 60 188 61 189
rect 59 188 60 189
rect 58 188 59 189
rect 57 188 58 189
rect 56 188 57 189
rect 55 188 56 189
rect 54 188 55 189
rect 53 188 54 189
rect 52 188 53 189
rect 51 188 52 189
rect 50 188 51 189
rect 49 188 50 189
rect 27 188 28 189
rect 26 188 27 189
rect 25 188 26 189
rect 21 188 22 189
rect 20 188 21 189
rect 19 188 20 189
rect 18 188 19 189
rect 15 188 16 189
rect 14 188 15 189
rect 13 188 14 189
rect 195 189 196 190
rect 194 189 195 190
rect 192 189 193 190
rect 191 189 192 190
rect 190 189 191 190
rect 189 189 190 190
rect 181 189 182 190
rect 180 189 181 190
rect 179 189 180 190
rect 178 189 179 190
rect 172 189 173 190
rect 171 189 172 190
rect 170 189 171 190
rect 169 189 170 190
rect 168 189 169 190
rect 165 189 166 190
rect 164 189 165 190
rect 163 189 164 190
rect 147 189 148 190
rect 146 189 147 190
rect 145 189 146 190
rect 144 189 145 190
rect 143 189 144 190
rect 142 189 143 190
rect 141 189 142 190
rect 140 189 141 190
rect 139 189 140 190
rect 138 189 139 190
rect 137 189 138 190
rect 136 189 137 190
rect 135 189 136 190
rect 134 189 135 190
rect 133 189 134 190
rect 132 189 133 190
rect 131 189 132 190
rect 130 189 131 190
rect 129 189 130 190
rect 128 189 129 190
rect 127 189 128 190
rect 126 189 127 190
rect 125 189 126 190
rect 124 189 125 190
rect 123 189 124 190
rect 122 189 123 190
rect 121 189 122 190
rect 120 189 121 190
rect 119 189 120 190
rect 118 189 119 190
rect 117 189 118 190
rect 116 189 117 190
rect 115 189 116 190
rect 114 189 115 190
rect 113 189 114 190
rect 112 189 113 190
rect 111 189 112 190
rect 110 189 111 190
rect 109 189 110 190
rect 108 189 109 190
rect 107 189 108 190
rect 106 189 107 190
rect 105 189 106 190
rect 104 189 105 190
rect 103 189 104 190
rect 102 189 103 190
rect 101 189 102 190
rect 100 189 101 190
rect 60 189 61 190
rect 59 189 60 190
rect 58 189 59 190
rect 57 189 58 190
rect 52 189 53 190
rect 51 189 52 190
rect 50 189 51 190
rect 49 189 50 190
rect 27 189 28 190
rect 26 189 27 190
rect 25 189 26 190
rect 20 189 21 190
rect 19 189 20 190
rect 18 189 19 190
rect 17 189 18 190
rect 16 189 17 190
rect 15 189 16 190
rect 14 189 15 190
rect 13 189 14 190
rect 194 190 195 191
rect 192 190 193 191
rect 191 190 192 191
rect 190 190 191 191
rect 189 190 190 191
rect 181 190 182 191
rect 180 190 181 191
rect 179 190 180 191
rect 178 190 179 191
rect 171 190 172 191
rect 170 190 171 191
rect 169 190 170 191
rect 165 190 166 191
rect 164 190 165 191
rect 163 190 164 191
rect 147 190 148 191
rect 146 190 147 191
rect 145 190 146 191
rect 144 190 145 191
rect 143 190 144 191
rect 142 190 143 191
rect 141 190 142 191
rect 140 190 141 191
rect 139 190 140 191
rect 138 190 139 191
rect 137 190 138 191
rect 136 190 137 191
rect 135 190 136 191
rect 134 190 135 191
rect 133 190 134 191
rect 132 190 133 191
rect 131 190 132 191
rect 130 190 131 191
rect 129 190 130 191
rect 128 190 129 191
rect 127 190 128 191
rect 126 190 127 191
rect 125 190 126 191
rect 124 190 125 191
rect 123 190 124 191
rect 122 190 123 191
rect 121 190 122 191
rect 120 190 121 191
rect 119 190 120 191
rect 118 190 119 191
rect 117 190 118 191
rect 116 190 117 191
rect 115 190 116 191
rect 114 190 115 191
rect 113 190 114 191
rect 112 190 113 191
rect 111 190 112 191
rect 110 190 111 191
rect 109 190 110 191
rect 108 190 109 191
rect 107 190 108 191
rect 106 190 107 191
rect 105 190 106 191
rect 104 190 105 191
rect 103 190 104 191
rect 102 190 103 191
rect 101 190 102 191
rect 100 190 101 191
rect 60 190 61 191
rect 59 190 60 191
rect 58 190 59 191
rect 57 190 58 191
rect 52 190 53 191
rect 51 190 52 191
rect 50 190 51 191
rect 49 190 50 191
rect 26 190 27 191
rect 25 190 26 191
rect 19 190 20 191
rect 18 190 19 191
rect 17 190 18 191
rect 16 190 17 191
rect 15 190 16 191
rect 14 190 15 191
rect 194 191 195 192
rect 192 191 193 192
rect 191 191 192 192
rect 181 191 182 192
rect 180 191 181 192
rect 179 191 180 192
rect 178 191 179 192
rect 164 191 165 192
rect 163 191 164 192
rect 147 191 148 192
rect 146 191 147 192
rect 145 191 146 192
rect 144 191 145 192
rect 143 191 144 192
rect 142 191 143 192
rect 141 191 142 192
rect 140 191 141 192
rect 139 191 140 192
rect 138 191 139 192
rect 137 191 138 192
rect 136 191 137 192
rect 135 191 136 192
rect 134 191 135 192
rect 133 191 134 192
rect 132 191 133 192
rect 131 191 132 192
rect 130 191 131 192
rect 129 191 130 192
rect 128 191 129 192
rect 127 191 128 192
rect 126 191 127 192
rect 125 191 126 192
rect 124 191 125 192
rect 123 191 124 192
rect 122 191 123 192
rect 121 191 122 192
rect 120 191 121 192
rect 119 191 120 192
rect 118 191 119 192
rect 117 191 118 192
rect 116 191 117 192
rect 115 191 116 192
rect 114 191 115 192
rect 113 191 114 192
rect 112 191 113 192
rect 111 191 112 192
rect 110 191 111 192
rect 109 191 110 192
rect 108 191 109 192
rect 107 191 108 192
rect 106 191 107 192
rect 105 191 106 192
rect 104 191 105 192
rect 103 191 104 192
rect 102 191 103 192
rect 101 191 102 192
rect 100 191 101 192
rect 60 191 61 192
rect 59 191 60 192
rect 58 191 59 192
rect 57 191 58 192
rect 52 191 53 192
rect 51 191 52 192
rect 50 191 51 192
rect 49 191 50 192
rect 18 191 19 192
rect 17 191 18 192
rect 16 191 17 192
rect 15 191 16 192
rect 193 192 194 193
rect 192 192 193 193
rect 191 192 192 193
rect 181 192 182 193
rect 180 192 181 193
rect 179 192 180 193
rect 178 192 179 193
rect 147 192 148 193
rect 146 192 147 193
rect 145 192 146 193
rect 144 192 145 193
rect 143 192 144 193
rect 142 192 143 193
rect 141 192 142 193
rect 140 192 141 193
rect 139 192 140 193
rect 138 192 139 193
rect 137 192 138 193
rect 136 192 137 193
rect 135 192 136 193
rect 134 192 135 193
rect 133 192 134 193
rect 132 192 133 193
rect 131 192 132 193
rect 130 192 131 193
rect 129 192 130 193
rect 128 192 129 193
rect 127 192 128 193
rect 126 192 127 193
rect 125 192 126 193
rect 124 192 125 193
rect 123 192 124 193
rect 122 192 123 193
rect 121 192 122 193
rect 120 192 121 193
rect 119 192 120 193
rect 118 192 119 193
rect 117 192 118 193
rect 116 192 117 193
rect 115 192 116 193
rect 114 192 115 193
rect 113 192 114 193
rect 112 192 113 193
rect 111 192 112 193
rect 110 192 111 193
rect 109 192 110 193
rect 108 192 109 193
rect 107 192 108 193
rect 106 192 107 193
rect 105 192 106 193
rect 104 192 105 193
rect 103 192 104 193
rect 102 192 103 193
rect 101 192 102 193
rect 100 192 101 193
rect 60 192 61 193
rect 59 192 60 193
rect 58 192 59 193
rect 57 192 58 193
rect 52 192 53 193
rect 51 192 52 193
rect 50 192 51 193
rect 49 192 50 193
rect 194 193 195 194
rect 193 193 194 194
rect 192 193 193 194
rect 191 193 192 194
rect 190 193 191 194
rect 189 193 190 194
rect 181 193 182 194
rect 180 193 181 194
rect 179 193 180 194
rect 178 193 179 194
rect 147 193 148 194
rect 146 193 147 194
rect 145 193 146 194
rect 144 193 145 194
rect 143 193 144 194
rect 142 193 143 194
rect 141 193 142 194
rect 140 193 141 194
rect 139 193 140 194
rect 138 193 139 194
rect 137 193 138 194
rect 136 193 137 194
rect 135 193 136 194
rect 134 193 135 194
rect 133 193 134 194
rect 132 193 133 194
rect 131 193 132 194
rect 130 193 131 194
rect 129 193 130 194
rect 128 193 129 194
rect 127 193 128 194
rect 126 193 127 194
rect 125 193 126 194
rect 124 193 125 194
rect 123 193 124 194
rect 122 193 123 194
rect 121 193 122 194
rect 120 193 121 194
rect 119 193 120 194
rect 118 193 119 194
rect 117 193 118 194
rect 116 193 117 194
rect 115 193 116 194
rect 114 193 115 194
rect 113 193 114 194
rect 112 193 113 194
rect 111 193 112 194
rect 110 193 111 194
rect 109 193 110 194
rect 108 193 109 194
rect 107 193 108 194
rect 106 193 107 194
rect 105 193 106 194
rect 104 193 105 194
rect 103 193 104 194
rect 102 193 103 194
rect 101 193 102 194
rect 100 193 101 194
rect 51 193 52 194
rect 50 193 51 194
rect 49 193 50 194
rect 25 193 26 194
rect 24 193 25 194
rect 23 193 24 194
rect 22 193 23 194
rect 21 193 22 194
rect 20 193 21 194
rect 19 193 20 194
rect 194 194 195 195
rect 193 194 194 195
rect 190 194 191 195
rect 189 194 190 195
rect 181 194 182 195
rect 180 194 181 195
rect 179 194 180 195
rect 178 194 179 195
rect 175 194 176 195
rect 174 194 175 195
rect 173 194 174 195
rect 172 194 173 195
rect 171 194 172 195
rect 170 194 171 195
rect 169 194 170 195
rect 168 194 169 195
rect 167 194 168 195
rect 166 194 167 195
rect 165 194 166 195
rect 164 194 165 195
rect 163 194 164 195
rect 162 194 163 195
rect 161 194 162 195
rect 160 194 161 195
rect 147 194 148 195
rect 146 194 147 195
rect 145 194 146 195
rect 144 194 145 195
rect 143 194 144 195
rect 142 194 143 195
rect 141 194 142 195
rect 140 194 141 195
rect 139 194 140 195
rect 138 194 139 195
rect 137 194 138 195
rect 136 194 137 195
rect 135 194 136 195
rect 134 194 135 195
rect 133 194 134 195
rect 132 194 133 195
rect 131 194 132 195
rect 130 194 131 195
rect 129 194 130 195
rect 128 194 129 195
rect 127 194 128 195
rect 126 194 127 195
rect 125 194 126 195
rect 124 194 125 195
rect 123 194 124 195
rect 122 194 123 195
rect 121 194 122 195
rect 120 194 121 195
rect 119 194 120 195
rect 118 194 119 195
rect 117 194 118 195
rect 116 194 117 195
rect 115 194 116 195
rect 114 194 115 195
rect 113 194 114 195
rect 112 194 113 195
rect 111 194 112 195
rect 110 194 111 195
rect 109 194 110 195
rect 108 194 109 195
rect 107 194 108 195
rect 106 194 107 195
rect 105 194 106 195
rect 104 194 105 195
rect 103 194 104 195
rect 102 194 103 195
rect 101 194 102 195
rect 100 194 101 195
rect 26 194 27 195
rect 25 194 26 195
rect 24 194 25 195
rect 23 194 24 195
rect 22 194 23 195
rect 21 194 22 195
rect 20 194 21 195
rect 19 194 20 195
rect 18 194 19 195
rect 17 194 18 195
rect 16 194 17 195
rect 195 195 196 196
rect 194 195 195 196
rect 190 195 191 196
rect 189 195 190 196
rect 181 195 182 196
rect 180 195 181 196
rect 179 195 180 196
rect 178 195 179 196
rect 175 195 176 196
rect 174 195 175 196
rect 173 195 174 196
rect 172 195 173 196
rect 171 195 172 196
rect 170 195 171 196
rect 169 195 170 196
rect 168 195 169 196
rect 167 195 168 196
rect 166 195 167 196
rect 165 195 166 196
rect 164 195 165 196
rect 163 195 164 196
rect 162 195 163 196
rect 161 195 162 196
rect 160 195 161 196
rect 147 195 148 196
rect 146 195 147 196
rect 145 195 146 196
rect 144 195 145 196
rect 143 195 144 196
rect 142 195 143 196
rect 141 195 142 196
rect 140 195 141 196
rect 139 195 140 196
rect 138 195 139 196
rect 137 195 138 196
rect 136 195 137 196
rect 135 195 136 196
rect 134 195 135 196
rect 133 195 134 196
rect 132 195 133 196
rect 131 195 132 196
rect 130 195 131 196
rect 129 195 130 196
rect 128 195 129 196
rect 127 195 128 196
rect 126 195 127 196
rect 125 195 126 196
rect 124 195 125 196
rect 123 195 124 196
rect 122 195 123 196
rect 121 195 122 196
rect 120 195 121 196
rect 119 195 120 196
rect 118 195 119 196
rect 117 195 118 196
rect 116 195 117 196
rect 115 195 116 196
rect 114 195 115 196
rect 113 195 114 196
rect 112 195 113 196
rect 111 195 112 196
rect 110 195 111 196
rect 109 195 110 196
rect 108 195 109 196
rect 107 195 108 196
rect 106 195 107 196
rect 105 195 106 196
rect 104 195 105 196
rect 103 195 104 196
rect 102 195 103 196
rect 101 195 102 196
rect 100 195 101 196
rect 76 195 77 196
rect 75 195 76 196
rect 74 195 75 196
rect 73 195 74 196
rect 72 195 73 196
rect 71 195 72 196
rect 70 195 71 196
rect 69 195 70 196
rect 68 195 69 196
rect 67 195 68 196
rect 66 195 67 196
rect 65 195 66 196
rect 64 195 65 196
rect 63 195 64 196
rect 62 195 63 196
rect 61 195 62 196
rect 60 195 61 196
rect 59 195 60 196
rect 58 195 59 196
rect 57 195 58 196
rect 53 195 54 196
rect 52 195 53 196
rect 51 195 52 196
rect 50 195 51 196
rect 49 195 50 196
rect 27 195 28 196
rect 26 195 27 196
rect 25 195 26 196
rect 24 195 25 196
rect 23 195 24 196
rect 22 195 23 196
rect 21 195 22 196
rect 20 195 21 196
rect 19 195 20 196
rect 18 195 19 196
rect 17 195 18 196
rect 16 195 17 196
rect 15 195 16 196
rect 195 196 196 197
rect 194 196 195 197
rect 190 196 191 197
rect 189 196 190 197
rect 181 196 182 197
rect 180 196 181 197
rect 179 196 180 197
rect 178 196 179 197
rect 175 196 176 197
rect 174 196 175 197
rect 173 196 174 197
rect 172 196 173 197
rect 171 196 172 197
rect 170 196 171 197
rect 169 196 170 197
rect 168 196 169 197
rect 167 196 168 197
rect 166 196 167 197
rect 165 196 166 197
rect 164 196 165 197
rect 163 196 164 197
rect 162 196 163 197
rect 161 196 162 197
rect 160 196 161 197
rect 147 196 148 197
rect 146 196 147 197
rect 145 196 146 197
rect 144 196 145 197
rect 143 196 144 197
rect 142 196 143 197
rect 141 196 142 197
rect 140 196 141 197
rect 139 196 140 197
rect 138 196 139 197
rect 137 196 138 197
rect 136 196 137 197
rect 135 196 136 197
rect 134 196 135 197
rect 133 196 134 197
rect 132 196 133 197
rect 131 196 132 197
rect 130 196 131 197
rect 129 196 130 197
rect 128 196 129 197
rect 127 196 128 197
rect 126 196 127 197
rect 125 196 126 197
rect 124 196 125 197
rect 123 196 124 197
rect 122 196 123 197
rect 121 196 122 197
rect 120 196 121 197
rect 119 196 120 197
rect 118 196 119 197
rect 117 196 118 197
rect 116 196 117 197
rect 115 196 116 197
rect 114 196 115 197
rect 113 196 114 197
rect 112 196 113 197
rect 111 196 112 197
rect 110 196 111 197
rect 109 196 110 197
rect 108 196 109 197
rect 107 196 108 197
rect 106 196 107 197
rect 105 196 106 197
rect 104 196 105 197
rect 103 196 104 197
rect 102 196 103 197
rect 101 196 102 197
rect 100 196 101 197
rect 76 196 77 197
rect 75 196 76 197
rect 74 196 75 197
rect 73 196 74 197
rect 72 196 73 197
rect 71 196 72 197
rect 70 196 71 197
rect 69 196 70 197
rect 68 196 69 197
rect 67 196 68 197
rect 66 196 67 197
rect 65 196 66 197
rect 64 196 65 197
rect 63 196 64 197
rect 62 196 63 197
rect 61 196 62 197
rect 60 196 61 197
rect 59 196 60 197
rect 58 196 59 197
rect 57 196 58 197
rect 53 196 54 197
rect 52 196 53 197
rect 51 196 52 197
rect 50 196 51 197
rect 49 196 50 197
rect 27 196 28 197
rect 26 196 27 197
rect 25 196 26 197
rect 19 196 20 197
rect 18 196 19 197
rect 17 196 18 197
rect 16 196 17 197
rect 15 196 16 197
rect 14 196 15 197
rect 189 197 190 198
rect 180 197 181 198
rect 179 197 180 198
rect 168 197 169 198
rect 167 197 168 198
rect 166 197 167 198
rect 147 197 148 198
rect 146 197 147 198
rect 145 197 146 198
rect 144 197 145 198
rect 143 197 144 198
rect 142 197 143 198
rect 141 197 142 198
rect 140 197 141 198
rect 139 197 140 198
rect 138 197 139 198
rect 137 197 138 198
rect 135 197 136 198
rect 134 197 135 198
rect 133 197 134 198
rect 132 197 133 198
rect 131 197 132 198
rect 130 197 131 198
rect 129 197 130 198
rect 128 197 129 198
rect 127 197 128 198
rect 126 197 127 198
rect 125 197 126 198
rect 124 197 125 198
rect 123 197 124 198
rect 122 197 123 198
rect 121 197 122 198
rect 120 197 121 198
rect 119 197 120 198
rect 118 197 119 198
rect 116 197 117 198
rect 115 197 116 198
rect 114 197 115 198
rect 113 197 114 198
rect 112 197 113 198
rect 110 197 111 198
rect 109 197 110 198
rect 108 197 109 198
rect 107 197 108 198
rect 106 197 107 198
rect 105 197 106 198
rect 104 197 105 198
rect 103 197 104 198
rect 102 197 103 198
rect 101 197 102 198
rect 100 197 101 198
rect 76 197 77 198
rect 75 197 76 198
rect 74 197 75 198
rect 73 197 74 198
rect 72 197 73 198
rect 71 197 72 198
rect 70 197 71 198
rect 69 197 70 198
rect 68 197 69 198
rect 67 197 68 198
rect 66 197 67 198
rect 65 197 66 198
rect 64 197 65 198
rect 63 197 64 198
rect 62 197 63 198
rect 61 197 62 198
rect 60 197 61 198
rect 59 197 60 198
rect 58 197 59 198
rect 57 197 58 198
rect 53 197 54 198
rect 52 197 53 198
rect 51 197 52 198
rect 50 197 51 198
rect 49 197 50 198
rect 27 197 28 198
rect 26 197 27 198
rect 25 197 26 198
rect 16 197 17 198
rect 15 197 16 198
rect 14 197 15 198
rect 13 197 14 198
rect 193 198 194 199
rect 192 198 193 199
rect 191 198 192 199
rect 190 198 191 199
rect 189 198 190 199
rect 188 198 189 199
rect 168 198 169 199
rect 167 198 168 199
rect 166 198 167 199
rect 147 198 148 199
rect 146 198 147 199
rect 145 198 146 199
rect 144 198 145 199
rect 143 198 144 199
rect 142 198 143 199
rect 141 198 142 199
rect 140 198 141 199
rect 139 198 140 199
rect 138 198 139 199
rect 129 198 130 199
rect 128 198 129 199
rect 127 198 128 199
rect 126 198 127 199
rect 125 198 126 199
rect 124 198 125 199
rect 123 198 124 199
rect 122 198 123 199
rect 121 198 122 199
rect 120 198 121 199
rect 119 198 120 199
rect 110 198 111 199
rect 109 198 110 199
rect 108 198 109 199
rect 107 198 108 199
rect 106 198 107 199
rect 105 198 106 199
rect 104 198 105 199
rect 103 198 104 199
rect 102 198 103 199
rect 101 198 102 199
rect 100 198 101 199
rect 76 198 77 199
rect 75 198 76 199
rect 74 198 75 199
rect 73 198 74 199
rect 72 198 73 199
rect 71 198 72 199
rect 70 198 71 199
rect 69 198 70 199
rect 68 198 69 199
rect 67 198 68 199
rect 66 198 67 199
rect 65 198 66 199
rect 64 198 65 199
rect 63 198 64 199
rect 62 198 63 199
rect 61 198 62 199
rect 60 198 61 199
rect 59 198 60 199
rect 58 198 59 199
rect 57 198 58 199
rect 53 198 54 199
rect 52 198 53 199
rect 51 198 52 199
rect 50 198 51 199
rect 49 198 50 199
rect 27 198 28 199
rect 26 198 27 199
rect 25 198 26 199
rect 15 198 16 199
rect 14 198 15 199
rect 13 198 14 199
rect 194 199 195 200
rect 193 199 194 200
rect 192 199 193 200
rect 191 199 192 200
rect 190 199 191 200
rect 189 199 190 200
rect 188 199 189 200
rect 187 199 188 200
rect 168 199 169 200
rect 167 199 168 200
rect 166 199 167 200
rect 147 199 148 200
rect 146 199 147 200
rect 145 199 146 200
rect 144 199 145 200
rect 143 199 144 200
rect 142 199 143 200
rect 141 199 142 200
rect 140 199 141 200
rect 139 199 140 200
rect 138 199 139 200
rect 128 199 129 200
rect 127 199 128 200
rect 126 199 127 200
rect 125 199 126 200
rect 124 199 125 200
rect 123 199 124 200
rect 122 199 123 200
rect 121 199 122 200
rect 120 199 121 200
rect 119 199 120 200
rect 110 199 111 200
rect 109 199 110 200
rect 108 199 109 200
rect 107 199 108 200
rect 106 199 107 200
rect 105 199 106 200
rect 104 199 105 200
rect 103 199 104 200
rect 102 199 103 200
rect 101 199 102 200
rect 100 199 101 200
rect 76 199 77 200
rect 75 199 76 200
rect 74 199 75 200
rect 73 199 74 200
rect 72 199 73 200
rect 71 199 72 200
rect 70 199 71 200
rect 69 199 70 200
rect 68 199 69 200
rect 67 199 68 200
rect 66 199 67 200
rect 65 199 66 200
rect 64 199 65 200
rect 63 199 64 200
rect 62 199 63 200
rect 61 199 62 200
rect 60 199 61 200
rect 59 199 60 200
rect 58 199 59 200
rect 57 199 58 200
rect 53 199 54 200
rect 52 199 53 200
rect 51 199 52 200
rect 50 199 51 200
rect 49 199 50 200
rect 26 199 27 200
rect 25 199 26 200
rect 24 199 25 200
rect 23 199 24 200
rect 15 199 16 200
rect 14 199 15 200
rect 13 199 14 200
rect 194 200 195 201
rect 193 200 194 201
rect 192 200 193 201
rect 191 200 192 201
rect 190 200 191 201
rect 189 200 190 201
rect 188 200 189 201
rect 187 200 188 201
rect 147 200 148 201
rect 146 200 147 201
rect 145 200 146 201
rect 144 200 145 201
rect 143 200 144 201
rect 142 200 143 201
rect 141 200 142 201
rect 140 200 141 201
rect 139 200 140 201
rect 138 200 139 201
rect 128 200 129 201
rect 127 200 128 201
rect 126 200 127 201
rect 125 200 126 201
rect 124 200 125 201
rect 123 200 124 201
rect 122 200 123 201
rect 121 200 122 201
rect 120 200 121 201
rect 119 200 120 201
rect 110 200 111 201
rect 109 200 110 201
rect 108 200 109 201
rect 107 200 108 201
rect 106 200 107 201
rect 105 200 106 201
rect 104 200 105 201
rect 103 200 104 201
rect 102 200 103 201
rect 101 200 102 201
rect 100 200 101 201
rect 76 200 77 201
rect 75 200 76 201
rect 74 200 75 201
rect 73 200 74 201
rect 72 200 73 201
rect 71 200 72 201
rect 70 200 71 201
rect 69 200 70 201
rect 68 200 69 201
rect 67 200 68 201
rect 66 200 67 201
rect 65 200 66 201
rect 64 200 65 201
rect 63 200 64 201
rect 62 200 63 201
rect 61 200 62 201
rect 60 200 61 201
rect 59 200 60 201
rect 58 200 59 201
rect 57 200 58 201
rect 53 200 54 201
rect 52 200 53 201
rect 51 200 52 201
rect 50 200 51 201
rect 49 200 50 201
rect 26 200 27 201
rect 25 200 26 201
rect 24 200 25 201
rect 23 200 24 201
rect 22 200 23 201
rect 21 200 22 201
rect 20 200 21 201
rect 19 200 20 201
rect 15 200 16 201
rect 14 200 15 201
rect 13 200 14 201
rect 194 201 195 202
rect 189 201 190 202
rect 147 201 148 202
rect 146 201 147 202
rect 145 201 146 202
rect 144 201 145 202
rect 143 201 144 202
rect 142 201 143 202
rect 141 201 142 202
rect 140 201 141 202
rect 139 201 140 202
rect 138 201 139 202
rect 128 201 129 202
rect 127 201 128 202
rect 126 201 127 202
rect 125 201 126 202
rect 124 201 125 202
rect 123 201 124 202
rect 122 201 123 202
rect 121 201 122 202
rect 120 201 121 202
rect 119 201 120 202
rect 110 201 111 202
rect 109 201 110 202
rect 108 201 109 202
rect 107 201 108 202
rect 106 201 107 202
rect 105 201 106 202
rect 104 201 105 202
rect 103 201 104 202
rect 102 201 103 202
rect 101 201 102 202
rect 100 201 101 202
rect 25 201 26 202
rect 24 201 25 202
rect 23 201 24 202
rect 22 201 23 202
rect 21 201 22 202
rect 20 201 21 202
rect 19 201 20 202
rect 18 201 19 202
rect 17 201 18 202
rect 16 201 17 202
rect 15 201 16 202
rect 14 201 15 202
rect 13 201 14 202
rect 194 202 195 203
rect 193 202 194 203
rect 192 202 193 203
rect 191 202 192 203
rect 190 202 191 203
rect 189 202 190 203
rect 147 202 148 203
rect 146 202 147 203
rect 145 202 146 203
rect 144 202 145 203
rect 143 202 144 203
rect 142 202 143 203
rect 141 202 142 203
rect 140 202 141 203
rect 139 202 140 203
rect 138 202 139 203
rect 128 202 129 203
rect 127 202 128 203
rect 126 202 127 203
rect 125 202 126 203
rect 124 202 125 203
rect 123 202 124 203
rect 122 202 123 203
rect 121 202 122 203
rect 120 202 121 203
rect 119 202 120 203
rect 110 202 111 203
rect 109 202 110 203
rect 108 202 109 203
rect 107 202 108 203
rect 106 202 107 203
rect 105 202 106 203
rect 104 202 105 203
rect 103 202 104 203
rect 102 202 103 203
rect 101 202 102 203
rect 100 202 101 203
rect 23 202 24 203
rect 22 202 23 203
rect 21 202 22 203
rect 20 202 21 203
rect 19 202 20 203
rect 18 202 19 203
rect 17 202 18 203
rect 16 202 17 203
rect 15 202 16 203
rect 14 202 15 203
rect 195 203 196 204
rect 194 203 195 204
rect 193 203 194 204
rect 192 203 193 204
rect 191 203 192 204
rect 190 203 191 204
rect 189 203 190 204
rect 147 203 148 204
rect 146 203 147 204
rect 145 203 146 204
rect 144 203 145 204
rect 143 203 144 204
rect 142 203 143 204
rect 141 203 142 204
rect 140 203 141 204
rect 139 203 140 204
rect 138 203 139 204
rect 128 203 129 204
rect 127 203 128 204
rect 126 203 127 204
rect 125 203 126 204
rect 124 203 125 204
rect 123 203 124 204
rect 122 203 123 204
rect 121 203 122 204
rect 120 203 121 204
rect 119 203 120 204
rect 110 203 111 204
rect 109 203 110 204
rect 108 203 109 204
rect 107 203 108 204
rect 106 203 107 204
rect 105 203 106 204
rect 104 203 105 204
rect 103 203 104 204
rect 102 203 103 204
rect 101 203 102 204
rect 100 203 101 204
rect 20 203 21 204
rect 19 203 20 204
rect 18 203 19 204
rect 17 203 18 204
rect 16 203 17 204
rect 194 204 195 205
rect 193 204 194 205
rect 192 204 193 205
rect 191 204 192 205
rect 190 204 191 205
rect 189 204 190 205
rect 147 204 148 205
rect 146 204 147 205
rect 145 204 146 205
rect 144 204 145 205
rect 143 204 144 205
rect 142 204 143 205
rect 141 204 142 205
rect 140 204 141 205
rect 139 204 140 205
rect 138 204 139 205
rect 128 204 129 205
rect 127 204 128 205
rect 126 204 127 205
rect 125 204 126 205
rect 124 204 125 205
rect 123 204 124 205
rect 122 204 123 205
rect 121 204 122 205
rect 120 204 121 205
rect 119 204 120 205
rect 110 204 111 205
rect 109 204 110 205
rect 108 204 109 205
rect 107 204 108 205
rect 106 204 107 205
rect 105 204 106 205
rect 104 204 105 205
rect 103 204 104 205
rect 102 204 103 205
rect 101 204 102 205
rect 100 204 101 205
rect 190 205 191 206
rect 189 205 190 206
rect 147 205 148 206
rect 146 205 147 206
rect 145 205 146 206
rect 144 205 145 206
rect 143 205 144 206
rect 142 205 143 206
rect 141 205 142 206
rect 140 205 141 206
rect 139 205 140 206
rect 138 205 139 206
rect 128 205 129 206
rect 127 205 128 206
rect 126 205 127 206
rect 125 205 126 206
rect 124 205 125 206
rect 123 205 124 206
rect 122 205 123 206
rect 121 205 122 206
rect 120 205 121 206
rect 119 205 120 206
rect 110 205 111 206
rect 109 205 110 206
rect 108 205 109 206
rect 107 205 108 206
rect 106 205 107 206
rect 105 205 106 206
rect 104 205 105 206
rect 103 205 104 206
rect 102 205 103 206
rect 101 205 102 206
rect 100 205 101 206
rect 27 205 28 206
rect 26 205 27 206
rect 25 205 26 206
rect 193 206 194 207
rect 192 206 193 207
rect 191 206 192 207
rect 190 206 191 207
rect 189 206 190 207
rect 147 206 148 207
rect 146 206 147 207
rect 145 206 146 207
rect 144 206 145 207
rect 143 206 144 207
rect 142 206 143 207
rect 141 206 142 207
rect 140 206 141 207
rect 139 206 140 207
rect 138 206 139 207
rect 128 206 129 207
rect 127 206 128 207
rect 126 206 127 207
rect 125 206 126 207
rect 124 206 125 207
rect 123 206 124 207
rect 122 206 123 207
rect 121 206 122 207
rect 120 206 121 207
rect 119 206 120 207
rect 110 206 111 207
rect 109 206 110 207
rect 108 206 109 207
rect 107 206 108 207
rect 106 206 107 207
rect 105 206 106 207
rect 104 206 105 207
rect 103 206 104 207
rect 102 206 103 207
rect 101 206 102 207
rect 100 206 101 207
rect 76 206 77 207
rect 75 206 76 207
rect 74 206 75 207
rect 73 206 74 207
rect 72 206 73 207
rect 71 206 72 207
rect 70 206 71 207
rect 69 206 70 207
rect 68 206 69 207
rect 67 206 68 207
rect 66 206 67 207
rect 65 206 66 207
rect 64 206 65 207
rect 63 206 64 207
rect 62 206 63 207
rect 61 206 62 207
rect 60 206 61 207
rect 59 206 60 207
rect 58 206 59 207
rect 57 206 58 207
rect 27 206 28 207
rect 26 206 27 207
rect 25 206 26 207
rect 24 206 25 207
rect 17 206 18 207
rect 16 206 17 207
rect 194 207 195 208
rect 193 207 194 208
rect 192 207 193 208
rect 191 207 192 208
rect 190 207 191 208
rect 147 207 148 208
rect 146 207 147 208
rect 145 207 146 208
rect 144 207 145 208
rect 143 207 144 208
rect 142 207 143 208
rect 141 207 142 208
rect 140 207 141 208
rect 139 207 140 208
rect 138 207 139 208
rect 128 207 129 208
rect 127 207 128 208
rect 126 207 127 208
rect 125 207 126 208
rect 124 207 125 208
rect 123 207 124 208
rect 122 207 123 208
rect 121 207 122 208
rect 120 207 121 208
rect 119 207 120 208
rect 110 207 111 208
rect 109 207 110 208
rect 108 207 109 208
rect 107 207 108 208
rect 106 207 107 208
rect 105 207 106 208
rect 104 207 105 208
rect 103 207 104 208
rect 102 207 103 208
rect 101 207 102 208
rect 100 207 101 208
rect 76 207 77 208
rect 75 207 76 208
rect 74 207 75 208
rect 73 207 74 208
rect 72 207 73 208
rect 71 207 72 208
rect 70 207 71 208
rect 69 207 70 208
rect 68 207 69 208
rect 67 207 68 208
rect 66 207 67 208
rect 65 207 66 208
rect 64 207 65 208
rect 63 207 64 208
rect 62 207 63 208
rect 61 207 62 208
rect 60 207 61 208
rect 59 207 60 208
rect 58 207 59 208
rect 57 207 58 208
rect 27 207 28 208
rect 26 207 27 208
rect 25 207 26 208
rect 24 207 25 208
rect 23 207 24 208
rect 17 207 18 208
rect 16 207 17 208
rect 15 207 16 208
rect 14 207 15 208
rect 194 208 195 209
rect 193 208 194 209
rect 192 208 193 209
rect 191 208 192 209
rect 190 208 191 209
rect 189 208 190 209
rect 147 208 148 209
rect 146 208 147 209
rect 145 208 146 209
rect 144 208 145 209
rect 143 208 144 209
rect 142 208 143 209
rect 141 208 142 209
rect 140 208 141 209
rect 139 208 140 209
rect 138 208 139 209
rect 128 208 129 209
rect 127 208 128 209
rect 126 208 127 209
rect 125 208 126 209
rect 124 208 125 209
rect 123 208 124 209
rect 122 208 123 209
rect 121 208 122 209
rect 120 208 121 209
rect 119 208 120 209
rect 110 208 111 209
rect 109 208 110 209
rect 108 208 109 209
rect 107 208 108 209
rect 106 208 107 209
rect 105 208 106 209
rect 104 208 105 209
rect 103 208 104 209
rect 102 208 103 209
rect 101 208 102 209
rect 100 208 101 209
rect 76 208 77 209
rect 75 208 76 209
rect 74 208 75 209
rect 73 208 74 209
rect 72 208 73 209
rect 71 208 72 209
rect 70 208 71 209
rect 69 208 70 209
rect 68 208 69 209
rect 67 208 68 209
rect 66 208 67 209
rect 65 208 66 209
rect 64 208 65 209
rect 63 208 64 209
rect 62 208 63 209
rect 61 208 62 209
rect 60 208 61 209
rect 59 208 60 209
rect 58 208 59 209
rect 57 208 58 209
rect 27 208 28 209
rect 26 208 27 209
rect 25 208 26 209
rect 24 208 25 209
rect 23 208 24 209
rect 22 208 23 209
rect 17 208 18 209
rect 16 208 17 209
rect 15 208 16 209
rect 14 208 15 209
rect 13 208 14 209
rect 195 209 196 210
rect 194 209 195 210
rect 190 209 191 210
rect 189 209 190 210
rect 169 209 170 210
rect 147 209 148 210
rect 146 209 147 210
rect 145 209 146 210
rect 144 209 145 210
rect 143 209 144 210
rect 142 209 143 210
rect 141 209 142 210
rect 140 209 141 210
rect 139 209 140 210
rect 138 209 139 210
rect 128 209 129 210
rect 127 209 128 210
rect 126 209 127 210
rect 125 209 126 210
rect 124 209 125 210
rect 123 209 124 210
rect 122 209 123 210
rect 121 209 122 210
rect 120 209 121 210
rect 119 209 120 210
rect 110 209 111 210
rect 109 209 110 210
rect 108 209 109 210
rect 107 209 108 210
rect 106 209 107 210
rect 105 209 106 210
rect 104 209 105 210
rect 103 209 104 210
rect 102 209 103 210
rect 101 209 102 210
rect 100 209 101 210
rect 76 209 77 210
rect 75 209 76 210
rect 74 209 75 210
rect 73 209 74 210
rect 72 209 73 210
rect 71 209 72 210
rect 70 209 71 210
rect 69 209 70 210
rect 68 209 69 210
rect 67 209 68 210
rect 66 209 67 210
rect 65 209 66 210
rect 64 209 65 210
rect 63 209 64 210
rect 62 209 63 210
rect 61 209 62 210
rect 60 209 61 210
rect 59 209 60 210
rect 58 209 59 210
rect 57 209 58 210
rect 27 209 28 210
rect 26 209 27 210
rect 25 209 26 210
rect 24 209 25 210
rect 23 209 24 210
rect 22 209 23 210
rect 21 209 22 210
rect 16 209 17 210
rect 15 209 16 210
rect 14 209 15 210
rect 13 209 14 210
rect 195 210 196 211
rect 194 210 195 211
rect 190 210 191 211
rect 189 210 190 211
rect 171 210 172 211
rect 170 210 171 211
rect 169 210 170 211
rect 168 210 169 211
rect 147 210 148 211
rect 146 210 147 211
rect 145 210 146 211
rect 144 210 145 211
rect 143 210 144 211
rect 142 210 143 211
rect 141 210 142 211
rect 140 210 141 211
rect 139 210 140 211
rect 138 210 139 211
rect 128 210 129 211
rect 127 210 128 211
rect 126 210 127 211
rect 125 210 126 211
rect 124 210 125 211
rect 123 210 124 211
rect 122 210 123 211
rect 121 210 122 211
rect 120 210 121 211
rect 119 210 120 211
rect 110 210 111 211
rect 109 210 110 211
rect 108 210 109 211
rect 107 210 108 211
rect 106 210 107 211
rect 105 210 106 211
rect 104 210 105 211
rect 103 210 104 211
rect 102 210 103 211
rect 101 210 102 211
rect 100 210 101 211
rect 76 210 77 211
rect 75 210 76 211
rect 74 210 75 211
rect 73 210 74 211
rect 72 210 73 211
rect 71 210 72 211
rect 70 210 71 211
rect 69 210 70 211
rect 68 210 69 211
rect 67 210 68 211
rect 66 210 67 211
rect 65 210 66 211
rect 64 210 65 211
rect 63 210 64 211
rect 62 210 63 211
rect 61 210 62 211
rect 60 210 61 211
rect 59 210 60 211
rect 58 210 59 211
rect 57 210 58 211
rect 27 210 28 211
rect 26 210 27 211
rect 25 210 26 211
rect 23 210 24 211
rect 22 210 23 211
rect 21 210 22 211
rect 20 210 21 211
rect 15 210 16 211
rect 14 210 15 211
rect 13 210 14 211
rect 194 211 195 212
rect 193 211 194 212
rect 192 211 193 212
rect 191 211 192 212
rect 190 211 191 212
rect 189 211 190 212
rect 171 211 172 212
rect 170 211 171 212
rect 169 211 170 212
rect 168 211 169 212
rect 147 211 148 212
rect 146 211 147 212
rect 145 211 146 212
rect 144 211 145 212
rect 143 211 144 212
rect 142 211 143 212
rect 141 211 142 212
rect 140 211 141 212
rect 139 211 140 212
rect 138 211 139 212
rect 128 211 129 212
rect 127 211 128 212
rect 126 211 127 212
rect 125 211 126 212
rect 124 211 125 212
rect 123 211 124 212
rect 122 211 123 212
rect 121 211 122 212
rect 120 211 121 212
rect 119 211 120 212
rect 110 211 111 212
rect 109 211 110 212
rect 108 211 109 212
rect 107 211 108 212
rect 106 211 107 212
rect 105 211 106 212
rect 104 211 105 212
rect 103 211 104 212
rect 102 211 103 212
rect 101 211 102 212
rect 100 211 101 212
rect 64 211 65 212
rect 63 211 64 212
rect 62 211 63 212
rect 61 211 62 212
rect 60 211 61 212
rect 59 211 60 212
rect 58 211 59 212
rect 27 211 28 212
rect 26 211 27 212
rect 25 211 26 212
rect 22 211 23 212
rect 21 211 22 212
rect 20 211 21 212
rect 19 211 20 212
rect 15 211 16 212
rect 14 211 15 212
rect 13 211 14 212
rect 194 212 195 213
rect 193 212 194 213
rect 192 212 193 213
rect 191 212 192 213
rect 190 212 191 213
rect 176 212 177 213
rect 175 212 176 213
rect 171 212 172 213
rect 170 212 171 213
rect 169 212 170 213
rect 168 212 169 213
rect 162 212 163 213
rect 161 212 162 213
rect 147 212 148 213
rect 146 212 147 213
rect 145 212 146 213
rect 144 212 145 213
rect 143 212 144 213
rect 142 212 143 213
rect 141 212 142 213
rect 140 212 141 213
rect 139 212 140 213
rect 138 212 139 213
rect 128 212 129 213
rect 127 212 128 213
rect 126 212 127 213
rect 125 212 126 213
rect 124 212 125 213
rect 123 212 124 213
rect 122 212 123 213
rect 121 212 122 213
rect 120 212 121 213
rect 119 212 120 213
rect 110 212 111 213
rect 109 212 110 213
rect 108 212 109 213
rect 107 212 108 213
rect 106 212 107 213
rect 105 212 106 213
rect 104 212 105 213
rect 103 212 104 213
rect 102 212 103 213
rect 101 212 102 213
rect 100 212 101 213
rect 62 212 63 213
rect 61 212 62 213
rect 60 212 61 213
rect 59 212 60 213
rect 58 212 59 213
rect 57 212 58 213
rect 27 212 28 213
rect 26 212 27 213
rect 25 212 26 213
rect 21 212 22 213
rect 20 212 21 213
rect 19 212 20 213
rect 18 212 19 213
rect 17 212 18 213
rect 16 212 17 213
rect 15 212 16 213
rect 14 212 15 213
rect 13 212 14 213
rect 177 213 178 214
rect 176 213 177 214
rect 175 213 176 214
rect 174 213 175 214
rect 171 213 172 214
rect 170 213 171 214
rect 169 213 170 214
rect 168 213 169 214
rect 163 213 164 214
rect 162 213 163 214
rect 161 213 162 214
rect 160 213 161 214
rect 147 213 148 214
rect 146 213 147 214
rect 145 213 146 214
rect 144 213 145 214
rect 143 213 144 214
rect 142 213 143 214
rect 141 213 142 214
rect 140 213 141 214
rect 139 213 140 214
rect 138 213 139 214
rect 128 213 129 214
rect 127 213 128 214
rect 126 213 127 214
rect 125 213 126 214
rect 124 213 125 214
rect 123 213 124 214
rect 122 213 123 214
rect 121 213 122 214
rect 120 213 121 214
rect 119 213 120 214
rect 110 213 111 214
rect 109 213 110 214
rect 108 213 109 214
rect 107 213 108 214
rect 106 213 107 214
rect 105 213 106 214
rect 104 213 105 214
rect 103 213 104 214
rect 102 213 103 214
rect 101 213 102 214
rect 100 213 101 214
rect 61 213 62 214
rect 60 213 61 214
rect 59 213 60 214
rect 58 213 59 214
rect 57 213 58 214
rect 27 213 28 214
rect 26 213 27 214
rect 25 213 26 214
rect 20 213 21 214
rect 19 213 20 214
rect 18 213 19 214
rect 17 213 18 214
rect 16 213 17 214
rect 15 213 16 214
rect 14 213 15 214
rect 13 213 14 214
rect 194 214 195 215
rect 193 214 194 215
rect 192 214 193 215
rect 191 214 192 215
rect 190 214 191 215
rect 189 214 190 215
rect 177 214 178 215
rect 176 214 177 215
rect 175 214 176 215
rect 174 214 175 215
rect 171 214 172 215
rect 170 214 171 215
rect 169 214 170 215
rect 168 214 169 215
rect 163 214 164 215
rect 162 214 163 215
rect 161 214 162 215
rect 160 214 161 215
rect 147 214 148 215
rect 146 214 147 215
rect 145 214 146 215
rect 144 214 145 215
rect 143 214 144 215
rect 142 214 143 215
rect 141 214 142 215
rect 140 214 141 215
rect 139 214 140 215
rect 138 214 139 215
rect 128 214 129 215
rect 127 214 128 215
rect 126 214 127 215
rect 125 214 126 215
rect 124 214 125 215
rect 123 214 124 215
rect 122 214 123 215
rect 121 214 122 215
rect 120 214 121 215
rect 119 214 120 215
rect 110 214 111 215
rect 109 214 110 215
rect 108 214 109 215
rect 107 214 108 215
rect 106 214 107 215
rect 105 214 106 215
rect 104 214 105 215
rect 103 214 104 215
rect 102 214 103 215
rect 101 214 102 215
rect 100 214 101 215
rect 61 214 62 215
rect 60 214 61 215
rect 59 214 60 215
rect 58 214 59 215
rect 57 214 58 215
rect 56 214 57 215
rect 19 214 20 215
rect 18 214 19 215
rect 17 214 18 215
rect 16 214 17 215
rect 15 214 16 215
rect 14 214 15 215
rect 195 215 196 216
rect 194 215 195 216
rect 193 215 194 216
rect 192 215 193 216
rect 191 215 192 216
rect 190 215 191 216
rect 189 215 190 216
rect 177 215 178 216
rect 176 215 177 216
rect 175 215 176 216
rect 174 215 175 216
rect 171 215 172 216
rect 170 215 171 216
rect 169 215 170 216
rect 168 215 169 216
rect 163 215 164 216
rect 162 215 163 216
rect 161 215 162 216
rect 160 215 161 216
rect 147 215 148 216
rect 146 215 147 216
rect 145 215 146 216
rect 144 215 145 216
rect 143 215 144 216
rect 142 215 143 216
rect 141 215 142 216
rect 140 215 141 216
rect 139 215 140 216
rect 138 215 139 216
rect 128 215 129 216
rect 127 215 128 216
rect 126 215 127 216
rect 125 215 126 216
rect 124 215 125 216
rect 123 215 124 216
rect 122 215 123 216
rect 121 215 122 216
rect 120 215 121 216
rect 119 215 120 216
rect 110 215 111 216
rect 109 215 110 216
rect 108 215 109 216
rect 107 215 108 216
rect 106 215 107 216
rect 105 215 106 216
rect 104 215 105 216
rect 103 215 104 216
rect 102 215 103 216
rect 101 215 102 216
rect 100 215 101 216
rect 61 215 62 216
rect 60 215 61 216
rect 59 215 60 216
rect 58 215 59 216
rect 57 215 58 216
rect 56 215 57 216
rect 17 215 18 216
rect 16 215 17 216
rect 190 216 191 217
rect 189 216 190 217
rect 177 216 178 217
rect 176 216 177 217
rect 175 216 176 217
rect 174 216 175 217
rect 171 216 172 217
rect 170 216 171 217
rect 169 216 170 217
rect 168 216 169 217
rect 163 216 164 217
rect 162 216 163 217
rect 161 216 162 217
rect 160 216 161 217
rect 147 216 148 217
rect 146 216 147 217
rect 145 216 146 217
rect 144 216 145 217
rect 143 216 144 217
rect 142 216 143 217
rect 141 216 142 217
rect 140 216 141 217
rect 139 216 140 217
rect 138 216 139 217
rect 128 216 129 217
rect 127 216 128 217
rect 126 216 127 217
rect 125 216 126 217
rect 124 216 125 217
rect 123 216 124 217
rect 122 216 123 217
rect 121 216 122 217
rect 120 216 121 217
rect 119 216 120 217
rect 110 216 111 217
rect 109 216 110 217
rect 108 216 109 217
rect 107 216 108 217
rect 106 216 107 217
rect 105 216 106 217
rect 104 216 105 217
rect 103 216 104 217
rect 102 216 103 217
rect 101 216 102 217
rect 100 216 101 217
rect 61 216 62 217
rect 60 216 61 217
rect 59 216 60 217
rect 58 216 59 217
rect 57 216 58 217
rect 24 216 25 217
rect 23 216 24 217
rect 22 216 23 217
rect 190 217 191 218
rect 189 217 190 218
rect 177 217 178 218
rect 176 217 177 218
rect 175 217 176 218
rect 174 217 175 218
rect 171 217 172 218
rect 170 217 171 218
rect 169 217 170 218
rect 168 217 169 218
rect 163 217 164 218
rect 162 217 163 218
rect 161 217 162 218
rect 160 217 161 218
rect 147 217 148 218
rect 146 217 147 218
rect 145 217 146 218
rect 144 217 145 218
rect 143 217 144 218
rect 142 217 143 218
rect 141 217 142 218
rect 140 217 141 218
rect 139 217 140 218
rect 138 217 139 218
rect 128 217 129 218
rect 127 217 128 218
rect 126 217 127 218
rect 125 217 126 218
rect 124 217 125 218
rect 123 217 124 218
rect 122 217 123 218
rect 121 217 122 218
rect 120 217 121 218
rect 119 217 120 218
rect 110 217 111 218
rect 109 217 110 218
rect 108 217 109 218
rect 107 217 108 218
rect 106 217 107 218
rect 105 217 106 218
rect 104 217 105 218
rect 103 217 104 218
rect 102 217 103 218
rect 101 217 102 218
rect 100 217 101 218
rect 83 217 84 218
rect 82 217 83 218
rect 81 217 82 218
rect 61 217 62 218
rect 60 217 61 218
rect 59 217 60 218
rect 58 217 59 218
rect 57 217 58 218
rect 24 217 25 218
rect 23 217 24 218
rect 22 217 23 218
rect 21 217 22 218
rect 194 218 195 219
rect 193 218 194 219
rect 192 218 193 219
rect 191 218 192 219
rect 190 218 191 219
rect 189 218 190 219
rect 177 218 178 219
rect 176 218 177 219
rect 175 218 176 219
rect 174 218 175 219
rect 171 218 172 219
rect 170 218 171 219
rect 169 218 170 219
rect 168 218 169 219
rect 163 218 164 219
rect 162 218 163 219
rect 161 218 162 219
rect 160 218 161 219
rect 147 218 148 219
rect 146 218 147 219
rect 145 218 146 219
rect 144 218 145 219
rect 143 218 144 219
rect 142 218 143 219
rect 141 218 142 219
rect 140 218 141 219
rect 139 218 140 219
rect 138 218 139 219
rect 128 218 129 219
rect 127 218 128 219
rect 126 218 127 219
rect 125 218 126 219
rect 124 218 125 219
rect 123 218 124 219
rect 122 218 123 219
rect 121 218 122 219
rect 120 218 121 219
rect 119 218 120 219
rect 110 218 111 219
rect 109 218 110 219
rect 108 218 109 219
rect 107 218 108 219
rect 106 218 107 219
rect 105 218 106 219
rect 104 218 105 219
rect 103 218 104 219
rect 102 218 103 219
rect 101 218 102 219
rect 100 218 101 219
rect 84 218 85 219
rect 83 218 84 219
rect 82 218 83 219
rect 81 218 82 219
rect 58 218 59 219
rect 57 218 58 219
rect 24 218 25 219
rect 23 218 24 219
rect 22 218 23 219
rect 21 218 22 219
rect 20 218 21 219
rect 195 219 196 220
rect 194 219 195 220
rect 193 219 194 220
rect 192 219 193 220
rect 191 219 192 220
rect 190 219 191 220
rect 189 219 190 220
rect 177 219 178 220
rect 176 219 177 220
rect 175 219 176 220
rect 174 219 175 220
rect 171 219 172 220
rect 170 219 171 220
rect 169 219 170 220
rect 168 219 169 220
rect 163 219 164 220
rect 162 219 163 220
rect 161 219 162 220
rect 160 219 161 220
rect 147 219 148 220
rect 146 219 147 220
rect 145 219 146 220
rect 144 219 145 220
rect 143 219 144 220
rect 142 219 143 220
rect 141 219 142 220
rect 140 219 141 220
rect 139 219 140 220
rect 138 219 139 220
rect 128 219 129 220
rect 127 219 128 220
rect 126 219 127 220
rect 125 219 126 220
rect 124 219 125 220
rect 123 219 124 220
rect 122 219 123 220
rect 121 219 122 220
rect 120 219 121 220
rect 119 219 120 220
rect 110 219 111 220
rect 109 219 110 220
rect 108 219 109 220
rect 107 219 108 220
rect 106 219 107 220
rect 105 219 106 220
rect 104 219 105 220
rect 103 219 104 220
rect 102 219 103 220
rect 101 219 102 220
rect 100 219 101 220
rect 84 219 85 220
rect 83 219 84 220
rect 82 219 83 220
rect 81 219 82 220
rect 24 219 25 220
rect 23 219 24 220
rect 22 219 23 220
rect 21 219 22 220
rect 20 219 21 220
rect 19 219 20 220
rect 177 220 178 221
rect 176 220 177 221
rect 175 220 176 221
rect 174 220 175 221
rect 173 220 174 221
rect 172 220 173 221
rect 171 220 172 221
rect 170 220 171 221
rect 169 220 170 221
rect 168 220 169 221
rect 163 220 164 221
rect 162 220 163 221
rect 161 220 162 221
rect 160 220 161 221
rect 147 220 148 221
rect 146 220 147 221
rect 145 220 146 221
rect 144 220 145 221
rect 143 220 144 221
rect 142 220 143 221
rect 141 220 142 221
rect 140 220 141 221
rect 139 220 140 221
rect 138 220 139 221
rect 128 220 129 221
rect 127 220 128 221
rect 126 220 127 221
rect 125 220 126 221
rect 124 220 125 221
rect 123 220 124 221
rect 122 220 123 221
rect 121 220 122 221
rect 120 220 121 221
rect 119 220 120 221
rect 110 220 111 221
rect 109 220 110 221
rect 108 220 109 221
rect 107 220 108 221
rect 106 220 107 221
rect 105 220 106 221
rect 104 220 105 221
rect 103 220 104 221
rect 102 220 103 221
rect 101 220 102 221
rect 100 220 101 221
rect 84 220 85 221
rect 83 220 84 221
rect 82 220 83 221
rect 81 220 82 221
rect 24 220 25 221
rect 23 220 24 221
rect 22 220 23 221
rect 20 220 21 221
rect 19 220 20 221
rect 18 220 19 221
rect 194 221 195 222
rect 193 221 194 222
rect 192 221 193 222
rect 191 221 192 222
rect 190 221 191 222
rect 189 221 190 222
rect 187 221 188 222
rect 186 221 187 222
rect 177 221 178 222
rect 176 221 177 222
rect 175 221 176 222
rect 174 221 175 222
rect 173 221 174 222
rect 172 221 173 222
rect 171 221 172 222
rect 170 221 171 222
rect 169 221 170 222
rect 168 221 169 222
rect 163 221 164 222
rect 162 221 163 222
rect 161 221 162 222
rect 160 221 161 222
rect 147 221 148 222
rect 146 221 147 222
rect 145 221 146 222
rect 144 221 145 222
rect 143 221 144 222
rect 142 221 143 222
rect 141 221 142 222
rect 140 221 141 222
rect 139 221 140 222
rect 138 221 139 222
rect 128 221 129 222
rect 127 221 128 222
rect 126 221 127 222
rect 125 221 126 222
rect 124 221 125 222
rect 123 221 124 222
rect 122 221 123 222
rect 121 221 122 222
rect 120 221 121 222
rect 119 221 120 222
rect 110 221 111 222
rect 109 221 110 222
rect 108 221 109 222
rect 107 221 108 222
rect 106 221 107 222
rect 105 221 106 222
rect 104 221 105 222
rect 103 221 104 222
rect 102 221 103 222
rect 101 221 102 222
rect 100 221 101 222
rect 84 221 85 222
rect 83 221 84 222
rect 82 221 83 222
rect 81 221 82 222
rect 27 221 28 222
rect 26 221 27 222
rect 24 221 25 222
rect 23 221 24 222
rect 22 221 23 222
rect 19 221 20 222
rect 18 221 19 222
rect 17 221 18 222
rect 16 221 17 222
rect 194 222 195 223
rect 193 222 194 223
rect 192 222 193 223
rect 191 222 192 223
rect 190 222 191 223
rect 189 222 190 223
rect 187 222 188 223
rect 186 222 187 223
rect 177 222 178 223
rect 176 222 177 223
rect 175 222 176 223
rect 174 222 175 223
rect 173 222 174 223
rect 172 222 173 223
rect 171 222 172 223
rect 170 222 171 223
rect 169 222 170 223
rect 168 222 169 223
rect 163 222 164 223
rect 162 222 163 223
rect 161 222 162 223
rect 160 222 161 223
rect 147 222 148 223
rect 146 222 147 223
rect 145 222 146 223
rect 144 222 145 223
rect 143 222 144 223
rect 142 222 143 223
rect 141 222 142 223
rect 140 222 141 223
rect 139 222 140 223
rect 138 222 139 223
rect 128 222 129 223
rect 127 222 128 223
rect 126 222 127 223
rect 125 222 126 223
rect 124 222 125 223
rect 123 222 124 223
rect 122 222 123 223
rect 121 222 122 223
rect 120 222 121 223
rect 119 222 120 223
rect 110 222 111 223
rect 109 222 110 223
rect 108 222 109 223
rect 107 222 108 223
rect 106 222 107 223
rect 105 222 106 223
rect 104 222 105 223
rect 103 222 104 223
rect 102 222 103 223
rect 101 222 102 223
rect 100 222 101 223
rect 84 222 85 223
rect 83 222 84 223
rect 82 222 83 223
rect 81 222 82 223
rect 27 222 28 223
rect 26 222 27 223
rect 25 222 26 223
rect 24 222 25 223
rect 23 222 24 223
rect 22 222 23 223
rect 21 222 22 223
rect 18 222 19 223
rect 17 222 18 223
rect 16 222 17 223
rect 15 222 16 223
rect 177 223 178 224
rect 176 223 177 224
rect 175 223 176 224
rect 174 223 175 224
rect 171 223 172 224
rect 170 223 171 224
rect 169 223 170 224
rect 168 223 169 224
rect 163 223 164 224
rect 162 223 163 224
rect 161 223 162 224
rect 160 223 161 224
rect 147 223 148 224
rect 146 223 147 224
rect 145 223 146 224
rect 144 223 145 224
rect 143 223 144 224
rect 142 223 143 224
rect 141 223 142 224
rect 140 223 141 224
rect 139 223 140 224
rect 138 223 139 224
rect 128 223 129 224
rect 127 223 128 224
rect 126 223 127 224
rect 125 223 126 224
rect 124 223 125 224
rect 123 223 124 224
rect 122 223 123 224
rect 121 223 122 224
rect 120 223 121 224
rect 119 223 120 224
rect 110 223 111 224
rect 109 223 110 224
rect 108 223 109 224
rect 107 223 108 224
rect 106 223 107 224
rect 105 223 106 224
rect 104 223 105 224
rect 103 223 104 224
rect 102 223 103 224
rect 101 223 102 224
rect 100 223 101 224
rect 84 223 85 224
rect 83 223 84 224
rect 82 223 83 224
rect 81 223 82 224
rect 27 223 28 224
rect 26 223 27 224
rect 25 223 26 224
rect 24 223 25 224
rect 23 223 24 224
rect 22 223 23 224
rect 21 223 22 224
rect 20 223 21 224
rect 19 223 20 224
rect 18 223 19 224
rect 17 223 18 224
rect 16 223 17 224
rect 15 223 16 224
rect 14 223 15 224
rect 193 224 194 225
rect 192 224 193 225
rect 191 224 192 225
rect 190 224 191 225
rect 177 224 178 225
rect 176 224 177 225
rect 175 224 176 225
rect 174 224 175 225
rect 171 224 172 225
rect 170 224 171 225
rect 169 224 170 225
rect 168 224 169 225
rect 163 224 164 225
rect 162 224 163 225
rect 161 224 162 225
rect 160 224 161 225
rect 147 224 148 225
rect 146 224 147 225
rect 145 224 146 225
rect 144 224 145 225
rect 143 224 144 225
rect 142 224 143 225
rect 141 224 142 225
rect 140 224 141 225
rect 139 224 140 225
rect 138 224 139 225
rect 128 224 129 225
rect 127 224 128 225
rect 126 224 127 225
rect 125 224 126 225
rect 124 224 125 225
rect 123 224 124 225
rect 122 224 123 225
rect 121 224 122 225
rect 120 224 121 225
rect 119 224 120 225
rect 110 224 111 225
rect 109 224 110 225
rect 108 224 109 225
rect 107 224 108 225
rect 106 224 107 225
rect 105 224 106 225
rect 104 224 105 225
rect 103 224 104 225
rect 102 224 103 225
rect 101 224 102 225
rect 100 224 101 225
rect 84 224 85 225
rect 83 224 84 225
rect 82 224 83 225
rect 81 224 82 225
rect 25 224 26 225
rect 24 224 25 225
rect 23 224 24 225
rect 22 224 23 225
rect 21 224 22 225
rect 20 224 21 225
rect 19 224 20 225
rect 18 224 19 225
rect 17 224 18 225
rect 16 224 17 225
rect 15 224 16 225
rect 14 224 15 225
rect 13 224 14 225
rect 194 225 195 226
rect 193 225 194 226
rect 192 225 193 226
rect 191 225 192 226
rect 190 225 191 226
rect 189 225 190 226
rect 177 225 178 226
rect 176 225 177 226
rect 175 225 176 226
rect 174 225 175 226
rect 171 225 172 226
rect 170 225 171 226
rect 169 225 170 226
rect 168 225 169 226
rect 163 225 164 226
rect 162 225 163 226
rect 161 225 162 226
rect 160 225 161 226
rect 147 225 148 226
rect 146 225 147 226
rect 145 225 146 226
rect 144 225 145 226
rect 143 225 144 226
rect 142 225 143 226
rect 141 225 142 226
rect 140 225 141 226
rect 139 225 140 226
rect 138 225 139 226
rect 128 225 129 226
rect 127 225 128 226
rect 126 225 127 226
rect 125 225 126 226
rect 124 225 125 226
rect 123 225 124 226
rect 122 225 123 226
rect 121 225 122 226
rect 120 225 121 226
rect 119 225 120 226
rect 110 225 111 226
rect 109 225 110 226
rect 108 225 109 226
rect 107 225 108 226
rect 106 225 107 226
rect 105 225 106 226
rect 104 225 105 226
rect 103 225 104 226
rect 102 225 103 226
rect 101 225 102 226
rect 100 225 101 226
rect 84 225 85 226
rect 83 225 84 226
rect 82 225 83 226
rect 81 225 82 226
rect 24 225 25 226
rect 23 225 24 226
rect 22 225 23 226
rect 20 225 21 226
rect 19 225 20 226
rect 18 225 19 226
rect 17 225 18 226
rect 16 225 17 226
rect 15 225 16 226
rect 14 225 15 226
rect 13 225 14 226
rect 194 226 195 227
rect 193 226 194 227
rect 190 226 191 227
rect 189 226 190 227
rect 177 226 178 227
rect 176 226 177 227
rect 175 226 176 227
rect 174 226 175 227
rect 171 226 172 227
rect 170 226 171 227
rect 169 226 170 227
rect 168 226 169 227
rect 163 226 164 227
rect 162 226 163 227
rect 161 226 162 227
rect 160 226 161 227
rect 147 226 148 227
rect 146 226 147 227
rect 145 226 146 227
rect 144 226 145 227
rect 143 226 144 227
rect 142 226 143 227
rect 141 226 142 227
rect 140 226 141 227
rect 139 226 140 227
rect 138 226 139 227
rect 128 226 129 227
rect 127 226 128 227
rect 126 226 127 227
rect 125 226 126 227
rect 124 226 125 227
rect 123 226 124 227
rect 122 226 123 227
rect 121 226 122 227
rect 120 226 121 227
rect 119 226 120 227
rect 110 226 111 227
rect 109 226 110 227
rect 108 226 109 227
rect 107 226 108 227
rect 106 226 107 227
rect 105 226 106 227
rect 104 226 105 227
rect 103 226 104 227
rect 102 226 103 227
rect 101 226 102 227
rect 100 226 101 227
rect 84 226 85 227
rect 83 226 84 227
rect 82 226 83 227
rect 81 226 82 227
rect 23 226 24 227
rect 22 226 23 227
rect 16 226 17 227
rect 15 226 16 227
rect 14 226 15 227
rect 13 226 14 227
rect 195 227 196 228
rect 194 227 195 228
rect 190 227 191 228
rect 189 227 190 228
rect 181 227 182 228
rect 180 227 181 228
rect 179 227 180 228
rect 178 227 179 228
rect 177 227 178 228
rect 176 227 177 228
rect 175 227 176 228
rect 174 227 175 228
rect 171 227 172 228
rect 170 227 171 228
rect 169 227 170 228
rect 168 227 169 228
rect 167 227 168 228
rect 166 227 167 228
rect 165 227 166 228
rect 164 227 165 228
rect 163 227 164 228
rect 162 227 163 228
rect 161 227 162 228
rect 160 227 161 228
rect 147 227 148 228
rect 146 227 147 228
rect 145 227 146 228
rect 144 227 145 228
rect 143 227 144 228
rect 142 227 143 228
rect 141 227 142 228
rect 140 227 141 228
rect 139 227 140 228
rect 138 227 139 228
rect 128 227 129 228
rect 127 227 128 228
rect 126 227 127 228
rect 125 227 126 228
rect 124 227 125 228
rect 123 227 124 228
rect 122 227 123 228
rect 121 227 122 228
rect 120 227 121 228
rect 119 227 120 228
rect 110 227 111 228
rect 109 227 110 228
rect 108 227 109 228
rect 107 227 108 228
rect 106 227 107 228
rect 105 227 106 228
rect 104 227 105 228
rect 103 227 104 228
rect 102 227 103 228
rect 101 227 102 228
rect 100 227 101 228
rect 84 227 85 228
rect 83 227 84 228
rect 82 227 83 228
rect 81 227 82 228
rect 194 228 195 229
rect 189 228 190 229
rect 181 228 182 229
rect 180 228 181 229
rect 179 228 180 229
rect 178 228 179 229
rect 177 228 178 229
rect 176 228 177 229
rect 175 228 176 229
rect 174 228 175 229
rect 171 228 172 229
rect 170 228 171 229
rect 169 228 170 229
rect 168 228 169 229
rect 167 228 168 229
rect 166 228 167 229
rect 165 228 166 229
rect 164 228 165 229
rect 163 228 164 229
rect 162 228 163 229
rect 161 228 162 229
rect 160 228 161 229
rect 147 228 148 229
rect 146 228 147 229
rect 145 228 146 229
rect 144 228 145 229
rect 143 228 144 229
rect 142 228 143 229
rect 141 228 142 229
rect 140 228 141 229
rect 139 228 140 229
rect 138 228 139 229
rect 128 228 129 229
rect 127 228 128 229
rect 126 228 127 229
rect 125 228 126 229
rect 124 228 125 229
rect 123 228 124 229
rect 122 228 123 229
rect 121 228 122 229
rect 120 228 121 229
rect 119 228 120 229
rect 110 228 111 229
rect 109 228 110 229
rect 108 228 109 229
rect 107 228 108 229
rect 106 228 107 229
rect 105 228 106 229
rect 104 228 105 229
rect 103 228 104 229
rect 102 228 103 229
rect 101 228 102 229
rect 100 228 101 229
rect 84 228 85 229
rect 83 228 84 229
rect 82 228 83 229
rect 81 228 82 229
rect 23 228 24 229
rect 22 228 23 229
rect 21 228 22 229
rect 194 229 195 230
rect 191 229 192 230
rect 190 229 191 230
rect 181 229 182 230
rect 180 229 181 230
rect 179 229 180 230
rect 178 229 179 230
rect 177 229 178 230
rect 176 229 177 230
rect 175 229 176 230
rect 174 229 175 230
rect 171 229 172 230
rect 170 229 171 230
rect 169 229 170 230
rect 168 229 169 230
rect 167 229 168 230
rect 166 229 167 230
rect 165 229 166 230
rect 164 229 165 230
rect 163 229 164 230
rect 162 229 163 230
rect 161 229 162 230
rect 160 229 161 230
rect 147 229 148 230
rect 146 229 147 230
rect 145 229 146 230
rect 144 229 145 230
rect 143 229 144 230
rect 142 229 143 230
rect 141 229 142 230
rect 140 229 141 230
rect 139 229 140 230
rect 138 229 139 230
rect 128 229 129 230
rect 127 229 128 230
rect 126 229 127 230
rect 125 229 126 230
rect 124 229 125 230
rect 123 229 124 230
rect 122 229 123 230
rect 121 229 122 230
rect 120 229 121 230
rect 119 229 120 230
rect 110 229 111 230
rect 109 229 110 230
rect 108 229 109 230
rect 107 229 108 230
rect 106 229 107 230
rect 105 229 106 230
rect 104 229 105 230
rect 103 229 104 230
rect 102 229 103 230
rect 101 229 102 230
rect 100 229 101 230
rect 84 229 85 230
rect 83 229 84 230
rect 82 229 83 230
rect 81 229 82 230
rect 23 229 24 230
rect 22 229 23 230
rect 21 229 22 230
rect 195 230 196 231
rect 194 230 195 231
rect 192 230 193 231
rect 191 230 192 231
rect 190 230 191 231
rect 189 230 190 231
rect 181 230 182 231
rect 180 230 181 231
rect 179 230 180 231
rect 178 230 179 231
rect 177 230 178 231
rect 176 230 177 231
rect 175 230 176 231
rect 174 230 175 231
rect 171 230 172 231
rect 170 230 171 231
rect 169 230 170 231
rect 168 230 169 231
rect 167 230 168 231
rect 166 230 167 231
rect 165 230 166 231
rect 164 230 165 231
rect 163 230 164 231
rect 162 230 163 231
rect 161 230 162 231
rect 160 230 161 231
rect 147 230 148 231
rect 146 230 147 231
rect 145 230 146 231
rect 144 230 145 231
rect 143 230 144 231
rect 142 230 143 231
rect 141 230 142 231
rect 140 230 141 231
rect 139 230 140 231
rect 138 230 139 231
rect 128 230 129 231
rect 127 230 128 231
rect 126 230 127 231
rect 125 230 126 231
rect 124 230 125 231
rect 123 230 124 231
rect 122 230 123 231
rect 121 230 122 231
rect 120 230 121 231
rect 119 230 120 231
rect 110 230 111 231
rect 109 230 110 231
rect 108 230 109 231
rect 107 230 108 231
rect 106 230 107 231
rect 105 230 106 231
rect 104 230 105 231
rect 103 230 104 231
rect 102 230 103 231
rect 101 230 102 231
rect 100 230 101 231
rect 84 230 85 231
rect 83 230 84 231
rect 82 230 83 231
rect 81 230 82 231
rect 23 230 24 231
rect 22 230 23 231
rect 21 230 22 231
rect 195 231 196 232
rect 194 231 195 232
rect 192 231 193 232
rect 191 231 192 232
rect 190 231 191 232
rect 189 231 190 232
rect 171 231 172 232
rect 170 231 171 232
rect 169 231 170 232
rect 168 231 169 232
rect 162 231 163 232
rect 161 231 162 232
rect 147 231 148 232
rect 146 231 147 232
rect 145 231 146 232
rect 144 231 145 232
rect 143 231 144 232
rect 142 231 143 232
rect 141 231 142 232
rect 140 231 141 232
rect 139 231 140 232
rect 138 231 139 232
rect 128 231 129 232
rect 127 231 128 232
rect 126 231 127 232
rect 125 231 126 232
rect 124 231 125 232
rect 123 231 124 232
rect 122 231 123 232
rect 121 231 122 232
rect 120 231 121 232
rect 119 231 120 232
rect 110 231 111 232
rect 109 231 110 232
rect 108 231 109 232
rect 107 231 108 232
rect 106 231 107 232
rect 105 231 106 232
rect 104 231 105 232
rect 103 231 104 232
rect 102 231 103 232
rect 101 231 102 232
rect 100 231 101 232
rect 84 231 85 232
rect 83 231 84 232
rect 82 231 83 232
rect 81 231 82 232
rect 23 231 24 232
rect 22 231 23 232
rect 21 231 22 232
rect 195 232 196 233
rect 194 232 195 233
rect 193 232 194 233
rect 192 232 193 233
rect 190 232 191 233
rect 189 232 190 233
rect 171 232 172 233
rect 170 232 171 233
rect 169 232 170 233
rect 168 232 169 233
rect 147 232 148 233
rect 146 232 147 233
rect 145 232 146 233
rect 144 232 145 233
rect 143 232 144 233
rect 142 232 143 233
rect 141 232 142 233
rect 140 232 141 233
rect 139 232 140 233
rect 138 232 139 233
rect 128 232 129 233
rect 127 232 128 233
rect 126 232 127 233
rect 125 232 126 233
rect 124 232 125 233
rect 123 232 124 233
rect 122 232 123 233
rect 121 232 122 233
rect 120 232 121 233
rect 119 232 120 233
rect 110 232 111 233
rect 109 232 110 233
rect 108 232 109 233
rect 107 232 108 233
rect 106 232 107 233
rect 105 232 106 233
rect 104 232 105 233
rect 103 232 104 233
rect 102 232 103 233
rect 101 232 102 233
rect 100 232 101 233
rect 84 232 85 233
rect 83 232 84 233
rect 82 232 83 233
rect 81 232 82 233
rect 23 232 24 233
rect 22 232 23 233
rect 21 232 22 233
rect 194 233 195 234
rect 193 233 194 234
rect 192 233 193 234
rect 190 233 191 234
rect 189 233 190 234
rect 171 233 172 234
rect 170 233 171 234
rect 169 233 170 234
rect 168 233 169 234
rect 147 233 148 234
rect 146 233 147 234
rect 145 233 146 234
rect 144 233 145 234
rect 143 233 144 234
rect 142 233 143 234
rect 141 233 142 234
rect 140 233 141 234
rect 139 233 140 234
rect 138 233 139 234
rect 128 233 129 234
rect 127 233 128 234
rect 126 233 127 234
rect 125 233 126 234
rect 124 233 125 234
rect 123 233 124 234
rect 122 233 123 234
rect 121 233 122 234
rect 120 233 121 234
rect 119 233 120 234
rect 110 233 111 234
rect 109 233 110 234
rect 108 233 109 234
rect 107 233 108 234
rect 106 233 107 234
rect 105 233 106 234
rect 104 233 105 234
rect 103 233 104 234
rect 102 233 103 234
rect 101 233 102 234
rect 100 233 101 234
rect 84 233 85 234
rect 83 233 84 234
rect 82 233 83 234
rect 81 233 82 234
rect 23 233 24 234
rect 22 233 23 234
rect 21 233 22 234
rect 170 234 171 235
rect 169 234 170 235
rect 147 234 148 235
rect 146 234 147 235
rect 145 234 146 235
rect 144 234 145 235
rect 143 234 144 235
rect 142 234 143 235
rect 141 234 142 235
rect 140 234 141 235
rect 139 234 140 235
rect 138 234 139 235
rect 128 234 129 235
rect 127 234 128 235
rect 126 234 127 235
rect 125 234 126 235
rect 124 234 125 235
rect 123 234 124 235
rect 122 234 123 235
rect 121 234 122 235
rect 120 234 121 235
rect 119 234 120 235
rect 110 234 111 235
rect 109 234 110 235
rect 108 234 109 235
rect 107 234 108 235
rect 106 234 107 235
rect 105 234 106 235
rect 104 234 105 235
rect 103 234 104 235
rect 102 234 103 235
rect 101 234 102 235
rect 100 234 101 235
rect 84 234 85 235
rect 83 234 84 235
rect 82 234 83 235
rect 81 234 82 235
rect 147 235 148 236
rect 146 235 147 236
rect 145 235 146 236
rect 144 235 145 236
rect 143 235 144 236
rect 142 235 143 236
rect 141 235 142 236
rect 140 235 141 236
rect 139 235 140 236
rect 138 235 139 236
rect 128 235 129 236
rect 127 235 128 236
rect 126 235 127 236
rect 125 235 126 236
rect 124 235 125 236
rect 123 235 124 236
rect 122 235 123 236
rect 121 235 122 236
rect 120 235 121 236
rect 119 235 120 236
rect 110 235 111 236
rect 109 235 110 236
rect 108 235 109 236
rect 107 235 108 236
rect 106 235 107 236
rect 105 235 106 236
rect 104 235 105 236
rect 103 235 104 236
rect 102 235 103 236
rect 101 235 102 236
rect 100 235 101 236
rect 84 235 85 236
rect 83 235 84 236
rect 82 235 83 236
rect 81 235 82 236
rect 24 235 25 236
rect 23 235 24 236
rect 147 236 148 237
rect 146 236 147 237
rect 145 236 146 237
rect 144 236 145 237
rect 143 236 144 237
rect 142 236 143 237
rect 141 236 142 237
rect 140 236 141 237
rect 139 236 140 237
rect 138 236 139 237
rect 128 236 129 237
rect 127 236 128 237
rect 126 236 127 237
rect 125 236 126 237
rect 124 236 125 237
rect 123 236 124 237
rect 122 236 123 237
rect 121 236 122 237
rect 120 236 121 237
rect 119 236 120 237
rect 110 236 111 237
rect 109 236 110 237
rect 108 236 109 237
rect 107 236 108 237
rect 106 236 107 237
rect 105 236 106 237
rect 104 236 105 237
rect 103 236 104 237
rect 102 236 103 237
rect 101 236 102 237
rect 100 236 101 237
rect 84 236 85 237
rect 83 236 84 237
rect 82 236 83 237
rect 81 236 82 237
rect 26 236 27 237
rect 25 236 26 237
rect 24 236 25 237
rect 23 236 24 237
rect 147 237 148 238
rect 146 237 147 238
rect 145 237 146 238
rect 144 237 145 238
rect 143 237 144 238
rect 142 237 143 238
rect 141 237 142 238
rect 140 237 141 238
rect 139 237 140 238
rect 138 237 139 238
rect 128 237 129 238
rect 127 237 128 238
rect 126 237 127 238
rect 125 237 126 238
rect 124 237 125 238
rect 123 237 124 238
rect 122 237 123 238
rect 121 237 122 238
rect 120 237 121 238
rect 119 237 120 238
rect 110 237 111 238
rect 109 237 110 238
rect 108 237 109 238
rect 107 237 108 238
rect 106 237 107 238
rect 105 237 106 238
rect 104 237 105 238
rect 103 237 104 238
rect 102 237 103 238
rect 101 237 102 238
rect 100 237 101 238
rect 84 237 85 238
rect 83 237 84 238
rect 82 237 83 238
rect 81 237 82 238
rect 26 237 27 238
rect 25 237 26 238
rect 24 237 25 238
rect 23 237 24 238
rect 17 237 18 238
rect 16 237 17 238
rect 15 237 16 238
rect 194 238 195 239
rect 193 238 194 239
rect 192 238 193 239
rect 190 238 191 239
rect 189 238 190 239
rect 147 238 148 239
rect 146 238 147 239
rect 145 238 146 239
rect 144 238 145 239
rect 143 238 144 239
rect 142 238 143 239
rect 141 238 142 239
rect 140 238 141 239
rect 139 238 140 239
rect 138 238 139 239
rect 128 238 129 239
rect 127 238 128 239
rect 126 238 127 239
rect 125 238 126 239
rect 124 238 125 239
rect 123 238 124 239
rect 122 238 123 239
rect 121 238 122 239
rect 120 238 121 239
rect 119 238 120 239
rect 110 238 111 239
rect 109 238 110 239
rect 108 238 109 239
rect 107 238 108 239
rect 106 238 107 239
rect 105 238 106 239
rect 104 238 105 239
rect 103 238 104 239
rect 102 238 103 239
rect 101 238 102 239
rect 100 238 101 239
rect 84 238 85 239
rect 83 238 84 239
rect 82 238 83 239
rect 81 238 82 239
rect 27 238 28 239
rect 26 238 27 239
rect 25 238 26 239
rect 24 238 25 239
rect 17 238 18 239
rect 16 238 17 239
rect 15 238 16 239
rect 14 238 15 239
rect 194 239 195 240
rect 193 239 194 240
rect 192 239 193 240
rect 191 239 192 240
rect 190 239 191 240
rect 189 239 190 240
rect 147 239 148 240
rect 146 239 147 240
rect 145 239 146 240
rect 144 239 145 240
rect 143 239 144 240
rect 142 239 143 240
rect 141 239 142 240
rect 140 239 141 240
rect 139 239 140 240
rect 138 239 139 240
rect 128 239 129 240
rect 127 239 128 240
rect 126 239 127 240
rect 125 239 126 240
rect 124 239 125 240
rect 123 239 124 240
rect 122 239 123 240
rect 121 239 122 240
rect 120 239 121 240
rect 119 239 120 240
rect 110 239 111 240
rect 109 239 110 240
rect 108 239 109 240
rect 107 239 108 240
rect 106 239 107 240
rect 105 239 106 240
rect 104 239 105 240
rect 103 239 104 240
rect 102 239 103 240
rect 101 239 102 240
rect 100 239 101 240
rect 83 239 84 240
rect 82 239 83 240
rect 81 239 82 240
rect 27 239 28 240
rect 26 239 27 240
rect 25 239 26 240
rect 17 239 18 240
rect 16 239 17 240
rect 15 239 16 240
rect 14 239 15 240
rect 13 239 14 240
rect 195 240 196 241
rect 194 240 195 241
rect 192 240 193 241
rect 191 240 192 241
rect 190 240 191 241
rect 189 240 190 241
rect 147 240 148 241
rect 146 240 147 241
rect 145 240 146 241
rect 144 240 145 241
rect 143 240 144 241
rect 142 240 143 241
rect 141 240 142 241
rect 140 240 141 241
rect 139 240 140 241
rect 138 240 139 241
rect 128 240 129 241
rect 127 240 128 241
rect 126 240 127 241
rect 125 240 126 241
rect 124 240 125 241
rect 123 240 124 241
rect 122 240 123 241
rect 121 240 122 241
rect 120 240 121 241
rect 119 240 120 241
rect 110 240 111 241
rect 109 240 110 241
rect 108 240 109 241
rect 107 240 108 241
rect 106 240 107 241
rect 105 240 106 241
rect 104 240 105 241
rect 103 240 104 241
rect 102 240 103 241
rect 101 240 102 241
rect 100 240 101 241
rect 27 240 28 241
rect 26 240 27 241
rect 25 240 26 241
rect 20 240 21 241
rect 19 240 20 241
rect 15 240 16 241
rect 14 240 15 241
rect 13 240 14 241
rect 194 241 195 242
rect 193 241 194 242
rect 192 241 193 242
rect 191 241 192 242
rect 190 241 191 242
rect 189 241 190 242
rect 147 241 148 242
rect 146 241 147 242
rect 145 241 146 242
rect 144 241 145 242
rect 143 241 144 242
rect 142 241 143 242
rect 141 241 142 242
rect 140 241 141 242
rect 139 241 140 242
rect 138 241 139 242
rect 128 241 129 242
rect 127 241 128 242
rect 126 241 127 242
rect 125 241 126 242
rect 124 241 125 242
rect 123 241 124 242
rect 122 241 123 242
rect 121 241 122 242
rect 120 241 121 242
rect 119 241 120 242
rect 110 241 111 242
rect 109 241 110 242
rect 108 241 109 242
rect 107 241 108 242
rect 106 241 107 242
rect 105 241 106 242
rect 104 241 105 242
rect 103 241 104 242
rect 102 241 103 242
rect 101 241 102 242
rect 100 241 101 242
rect 27 241 28 242
rect 26 241 27 242
rect 25 241 26 242
rect 21 241 22 242
rect 20 241 21 242
rect 19 241 20 242
rect 18 241 19 242
rect 15 241 16 242
rect 14 241 15 242
rect 13 241 14 242
rect 195 242 196 243
rect 194 242 195 243
rect 193 242 194 243
rect 192 242 193 243
rect 191 242 192 243
rect 190 242 191 243
rect 189 242 190 243
rect 147 242 148 243
rect 146 242 147 243
rect 145 242 146 243
rect 144 242 145 243
rect 143 242 144 243
rect 142 242 143 243
rect 141 242 142 243
rect 140 242 141 243
rect 139 242 140 243
rect 138 242 139 243
rect 128 242 129 243
rect 127 242 128 243
rect 126 242 127 243
rect 125 242 126 243
rect 124 242 125 243
rect 123 242 124 243
rect 122 242 123 243
rect 121 242 122 243
rect 120 242 121 243
rect 119 242 120 243
rect 110 242 111 243
rect 109 242 110 243
rect 108 242 109 243
rect 107 242 108 243
rect 106 242 107 243
rect 105 242 106 243
rect 104 242 105 243
rect 103 242 104 243
rect 102 242 103 243
rect 101 242 102 243
rect 100 242 101 243
rect 84 242 85 243
rect 83 242 84 243
rect 82 242 83 243
rect 81 242 82 243
rect 80 242 81 243
rect 79 242 80 243
rect 78 242 79 243
rect 77 242 78 243
rect 76 242 77 243
rect 75 242 76 243
rect 74 242 75 243
rect 73 242 74 243
rect 72 242 73 243
rect 71 242 72 243
rect 70 242 71 243
rect 69 242 70 243
rect 68 242 69 243
rect 67 242 68 243
rect 66 242 67 243
rect 65 242 66 243
rect 64 242 65 243
rect 63 242 64 243
rect 62 242 63 243
rect 61 242 62 243
rect 60 242 61 243
rect 59 242 60 243
rect 58 242 59 243
rect 57 242 58 243
rect 26 242 27 243
rect 25 242 26 243
rect 24 242 25 243
rect 23 242 24 243
rect 22 242 23 243
rect 21 242 22 243
rect 20 242 21 243
rect 19 242 20 243
rect 18 242 19 243
rect 15 242 16 243
rect 14 242 15 243
rect 13 242 14 243
rect 194 243 195 244
rect 193 243 194 244
rect 192 243 193 244
rect 191 243 192 244
rect 190 243 191 244
rect 147 243 148 244
rect 146 243 147 244
rect 145 243 146 244
rect 144 243 145 244
rect 143 243 144 244
rect 142 243 143 244
rect 141 243 142 244
rect 140 243 141 244
rect 139 243 140 244
rect 138 243 139 244
rect 128 243 129 244
rect 127 243 128 244
rect 126 243 127 244
rect 125 243 126 244
rect 124 243 125 244
rect 123 243 124 244
rect 122 243 123 244
rect 121 243 122 244
rect 120 243 121 244
rect 119 243 120 244
rect 110 243 111 244
rect 109 243 110 244
rect 108 243 109 244
rect 107 243 108 244
rect 106 243 107 244
rect 105 243 106 244
rect 104 243 105 244
rect 103 243 104 244
rect 102 243 103 244
rect 101 243 102 244
rect 100 243 101 244
rect 84 243 85 244
rect 83 243 84 244
rect 82 243 83 244
rect 81 243 82 244
rect 80 243 81 244
rect 79 243 80 244
rect 78 243 79 244
rect 77 243 78 244
rect 76 243 77 244
rect 75 243 76 244
rect 74 243 75 244
rect 73 243 74 244
rect 72 243 73 244
rect 71 243 72 244
rect 70 243 71 244
rect 69 243 70 244
rect 68 243 69 244
rect 67 243 68 244
rect 66 243 67 244
rect 65 243 66 244
rect 64 243 65 244
rect 63 243 64 244
rect 62 243 63 244
rect 61 243 62 244
rect 60 243 61 244
rect 59 243 60 244
rect 58 243 59 244
rect 57 243 58 244
rect 26 243 27 244
rect 25 243 26 244
rect 24 243 25 244
rect 23 243 24 244
rect 22 243 23 244
rect 21 243 22 244
rect 20 243 21 244
rect 19 243 20 244
rect 18 243 19 244
rect 17 243 18 244
rect 16 243 17 244
rect 15 243 16 244
rect 14 243 15 244
rect 13 243 14 244
rect 147 244 148 245
rect 146 244 147 245
rect 145 244 146 245
rect 144 244 145 245
rect 143 244 144 245
rect 142 244 143 245
rect 141 244 142 245
rect 140 244 141 245
rect 139 244 140 245
rect 138 244 139 245
rect 128 244 129 245
rect 127 244 128 245
rect 126 244 127 245
rect 125 244 126 245
rect 124 244 125 245
rect 123 244 124 245
rect 122 244 123 245
rect 121 244 122 245
rect 120 244 121 245
rect 119 244 120 245
rect 110 244 111 245
rect 109 244 110 245
rect 108 244 109 245
rect 107 244 108 245
rect 106 244 107 245
rect 105 244 106 245
rect 104 244 105 245
rect 103 244 104 245
rect 102 244 103 245
rect 101 244 102 245
rect 100 244 101 245
rect 84 244 85 245
rect 83 244 84 245
rect 82 244 83 245
rect 81 244 82 245
rect 80 244 81 245
rect 79 244 80 245
rect 78 244 79 245
rect 77 244 78 245
rect 76 244 77 245
rect 75 244 76 245
rect 74 244 75 245
rect 73 244 74 245
rect 72 244 73 245
rect 71 244 72 245
rect 70 244 71 245
rect 69 244 70 245
rect 68 244 69 245
rect 67 244 68 245
rect 66 244 67 245
rect 65 244 66 245
rect 64 244 65 245
rect 63 244 64 245
rect 62 244 63 245
rect 61 244 62 245
rect 60 244 61 245
rect 59 244 60 245
rect 58 244 59 245
rect 57 244 58 245
rect 25 244 26 245
rect 24 244 25 245
rect 23 244 24 245
rect 22 244 23 245
rect 21 244 22 245
rect 19 244 20 245
rect 18 244 19 245
rect 17 244 18 245
rect 16 244 17 245
rect 15 244 16 245
rect 14 244 15 245
rect 195 245 196 246
rect 194 245 195 246
rect 193 245 194 246
rect 192 245 193 246
rect 191 245 192 246
rect 190 245 191 246
rect 189 245 190 246
rect 171 245 172 246
rect 170 245 171 246
rect 147 245 148 246
rect 146 245 147 246
rect 145 245 146 246
rect 144 245 145 246
rect 143 245 144 246
rect 142 245 143 246
rect 141 245 142 246
rect 140 245 141 246
rect 139 245 140 246
rect 138 245 139 246
rect 128 245 129 246
rect 127 245 128 246
rect 126 245 127 246
rect 125 245 126 246
rect 124 245 125 246
rect 123 245 124 246
rect 122 245 123 246
rect 121 245 122 246
rect 120 245 121 246
rect 119 245 120 246
rect 110 245 111 246
rect 109 245 110 246
rect 108 245 109 246
rect 107 245 108 246
rect 106 245 107 246
rect 105 245 106 246
rect 104 245 105 246
rect 103 245 104 246
rect 102 245 103 246
rect 101 245 102 246
rect 100 245 101 246
rect 84 245 85 246
rect 83 245 84 246
rect 82 245 83 246
rect 81 245 82 246
rect 80 245 81 246
rect 79 245 80 246
rect 78 245 79 246
rect 77 245 78 246
rect 76 245 77 246
rect 75 245 76 246
rect 74 245 75 246
rect 73 245 74 246
rect 72 245 73 246
rect 71 245 72 246
rect 70 245 71 246
rect 69 245 70 246
rect 68 245 69 246
rect 67 245 68 246
rect 66 245 67 246
rect 65 245 66 246
rect 64 245 65 246
rect 63 245 64 246
rect 62 245 63 246
rect 61 245 62 246
rect 60 245 61 246
rect 59 245 60 246
rect 58 245 59 246
rect 57 245 58 246
rect 23 245 24 246
rect 22 245 23 246
rect 18 245 19 246
rect 17 245 18 246
rect 16 245 17 246
rect 15 245 16 246
rect 194 246 195 247
rect 193 246 194 247
rect 192 246 193 247
rect 191 246 192 247
rect 190 246 191 247
rect 189 246 190 247
rect 172 246 173 247
rect 171 246 172 247
rect 170 246 171 247
rect 163 246 164 247
rect 162 246 163 247
rect 161 246 162 247
rect 147 246 148 247
rect 146 246 147 247
rect 145 246 146 247
rect 144 246 145 247
rect 143 246 144 247
rect 142 246 143 247
rect 141 246 142 247
rect 140 246 141 247
rect 139 246 140 247
rect 138 246 139 247
rect 128 246 129 247
rect 127 246 128 247
rect 126 246 127 247
rect 125 246 126 247
rect 124 246 125 247
rect 123 246 124 247
rect 122 246 123 247
rect 121 246 122 247
rect 120 246 121 247
rect 119 246 120 247
rect 110 246 111 247
rect 109 246 110 247
rect 108 246 109 247
rect 107 246 108 247
rect 106 246 107 247
rect 105 246 106 247
rect 104 246 105 247
rect 103 246 104 247
rect 102 246 103 247
rect 101 246 102 247
rect 100 246 101 247
rect 84 246 85 247
rect 83 246 84 247
rect 82 246 83 247
rect 81 246 82 247
rect 80 246 81 247
rect 79 246 80 247
rect 78 246 79 247
rect 77 246 78 247
rect 76 246 77 247
rect 75 246 76 247
rect 74 246 75 247
rect 73 246 74 247
rect 72 246 73 247
rect 71 246 72 247
rect 70 246 71 247
rect 69 246 70 247
rect 68 246 69 247
rect 67 246 68 247
rect 66 246 67 247
rect 65 246 66 247
rect 64 246 65 247
rect 63 246 64 247
rect 62 246 63 247
rect 61 246 62 247
rect 60 246 61 247
rect 59 246 60 247
rect 58 246 59 247
rect 57 246 58 247
rect 190 247 191 248
rect 189 247 190 248
rect 172 247 173 248
rect 171 247 172 248
rect 170 247 171 248
rect 169 247 170 248
rect 163 247 164 248
rect 162 247 163 248
rect 161 247 162 248
rect 147 247 148 248
rect 146 247 147 248
rect 145 247 146 248
rect 144 247 145 248
rect 143 247 144 248
rect 142 247 143 248
rect 141 247 142 248
rect 140 247 141 248
rect 139 247 140 248
rect 138 247 139 248
rect 128 247 129 248
rect 127 247 128 248
rect 126 247 127 248
rect 125 247 126 248
rect 124 247 125 248
rect 123 247 124 248
rect 122 247 123 248
rect 121 247 122 248
rect 120 247 121 248
rect 119 247 120 248
rect 110 247 111 248
rect 109 247 110 248
rect 108 247 109 248
rect 107 247 108 248
rect 106 247 107 248
rect 105 247 106 248
rect 104 247 105 248
rect 103 247 104 248
rect 102 247 103 248
rect 101 247 102 248
rect 100 247 101 248
rect 74 247 75 248
rect 73 247 74 248
rect 72 247 73 248
rect 71 247 72 248
rect 70 247 71 248
rect 69 247 70 248
rect 68 247 69 248
rect 64 247 65 248
rect 63 247 64 248
rect 62 247 63 248
rect 61 247 62 248
rect 60 247 61 248
rect 59 247 60 248
rect 194 248 195 249
rect 193 248 194 249
rect 192 248 193 249
rect 191 248 192 249
rect 190 248 191 249
rect 189 248 190 249
rect 172 248 173 249
rect 171 248 172 249
rect 170 248 171 249
rect 169 248 170 249
rect 168 248 169 249
rect 163 248 164 249
rect 162 248 163 249
rect 161 248 162 249
rect 147 248 148 249
rect 146 248 147 249
rect 145 248 146 249
rect 144 248 145 249
rect 143 248 144 249
rect 142 248 143 249
rect 141 248 142 249
rect 140 248 141 249
rect 139 248 140 249
rect 138 248 139 249
rect 128 248 129 249
rect 127 248 128 249
rect 126 248 127 249
rect 125 248 126 249
rect 124 248 125 249
rect 123 248 124 249
rect 122 248 123 249
rect 121 248 122 249
rect 120 248 121 249
rect 119 248 120 249
rect 110 248 111 249
rect 109 248 110 249
rect 108 248 109 249
rect 107 248 108 249
rect 106 248 107 249
rect 105 248 106 249
rect 104 248 105 249
rect 103 248 104 249
rect 102 248 103 249
rect 101 248 102 249
rect 100 248 101 249
rect 75 248 76 249
rect 74 248 75 249
rect 73 248 74 249
rect 72 248 73 249
rect 71 248 72 249
rect 61 248 62 249
rect 60 248 61 249
rect 59 248 60 249
rect 58 248 59 249
rect 195 249 196 250
rect 194 249 195 250
rect 193 249 194 250
rect 192 249 193 250
rect 191 249 192 250
rect 190 249 191 250
rect 189 249 190 250
rect 180 249 181 250
rect 179 249 180 250
rect 178 249 179 250
rect 177 249 178 250
rect 176 249 177 250
rect 175 249 176 250
rect 174 249 175 250
rect 171 249 172 250
rect 170 249 171 250
rect 169 249 170 250
rect 168 249 169 250
rect 167 249 168 250
rect 163 249 164 250
rect 162 249 163 250
rect 161 249 162 250
rect 147 249 148 250
rect 146 249 147 250
rect 145 249 146 250
rect 144 249 145 250
rect 143 249 144 250
rect 142 249 143 250
rect 141 249 142 250
rect 140 249 141 250
rect 139 249 140 250
rect 138 249 139 250
rect 128 249 129 250
rect 127 249 128 250
rect 126 249 127 250
rect 125 249 126 250
rect 124 249 125 250
rect 123 249 124 250
rect 122 249 123 250
rect 121 249 122 250
rect 120 249 121 250
rect 119 249 120 250
rect 110 249 111 250
rect 109 249 110 250
rect 108 249 109 250
rect 107 249 108 250
rect 106 249 107 250
rect 105 249 106 250
rect 104 249 105 250
rect 103 249 104 250
rect 102 249 103 250
rect 101 249 102 250
rect 100 249 101 250
rect 75 249 76 250
rect 74 249 75 250
rect 73 249 74 250
rect 72 249 73 250
rect 60 249 61 250
rect 59 249 60 250
rect 58 249 59 250
rect 57 249 58 250
rect 194 250 195 251
rect 193 250 194 251
rect 192 250 193 251
rect 191 250 192 251
rect 190 250 191 251
rect 181 250 182 251
rect 180 250 181 251
rect 179 250 180 251
rect 178 250 179 251
rect 177 250 178 251
rect 176 250 177 251
rect 175 250 176 251
rect 174 250 175 251
rect 171 250 172 251
rect 170 250 171 251
rect 169 250 170 251
rect 168 250 169 251
rect 167 250 168 251
rect 166 250 167 251
rect 163 250 164 251
rect 162 250 163 251
rect 161 250 162 251
rect 76 250 77 251
rect 75 250 76 251
rect 74 250 75 251
rect 73 250 74 251
rect 60 250 61 251
rect 59 250 60 251
rect 58 250 59 251
rect 57 250 58 251
rect 193 251 194 252
rect 192 251 193 252
rect 191 251 192 252
rect 181 251 182 252
rect 180 251 181 252
rect 179 251 180 252
rect 178 251 179 252
rect 177 251 178 252
rect 176 251 177 252
rect 175 251 176 252
rect 174 251 175 252
rect 170 251 171 252
rect 169 251 170 252
rect 168 251 169 252
rect 167 251 168 252
rect 166 251 167 252
rect 165 251 166 252
rect 164 251 165 252
rect 163 251 164 252
rect 162 251 163 252
rect 161 251 162 252
rect 76 251 77 252
rect 75 251 76 252
rect 74 251 75 252
rect 73 251 74 252
rect 60 251 61 252
rect 59 251 60 252
rect 58 251 59 252
rect 57 251 58 252
rect 194 252 195 253
rect 193 252 194 253
rect 192 252 193 253
rect 191 252 192 253
rect 190 252 191 253
rect 189 252 190 253
rect 181 252 182 253
rect 180 252 181 253
rect 179 252 180 253
rect 178 252 179 253
rect 177 252 178 253
rect 176 252 177 253
rect 175 252 176 253
rect 174 252 175 253
rect 169 252 170 253
rect 168 252 169 253
rect 167 252 168 253
rect 166 252 167 253
rect 165 252 166 253
rect 164 252 165 253
rect 163 252 164 253
rect 162 252 163 253
rect 161 252 162 253
rect 76 252 77 253
rect 75 252 76 253
rect 74 252 75 253
rect 73 252 74 253
rect 60 252 61 253
rect 59 252 60 253
rect 58 252 59 253
rect 57 252 58 253
rect 56 252 57 253
rect 194 253 195 254
rect 193 253 194 254
rect 192 253 193 254
rect 191 253 192 254
rect 190 253 191 254
rect 189 253 190 254
rect 181 253 182 254
rect 180 253 181 254
rect 179 253 180 254
rect 178 253 179 254
rect 169 253 170 254
rect 168 253 169 254
rect 167 253 168 254
rect 166 253 167 254
rect 165 253 166 254
rect 164 253 165 254
rect 163 253 164 254
rect 162 253 163 254
rect 161 253 162 254
rect 76 253 77 254
rect 75 253 76 254
rect 74 253 75 254
rect 73 253 74 254
rect 60 253 61 254
rect 59 253 60 254
rect 58 253 59 254
rect 57 253 58 254
rect 56 253 57 254
rect 27 253 28 254
rect 26 253 27 254
rect 25 253 26 254
rect 24 253 25 254
rect 195 254 196 255
rect 194 254 195 255
rect 190 254 191 255
rect 189 254 190 255
rect 181 254 182 255
rect 180 254 181 255
rect 179 254 180 255
rect 178 254 179 255
rect 170 254 171 255
rect 169 254 170 255
rect 168 254 169 255
rect 167 254 168 255
rect 166 254 167 255
rect 165 254 166 255
rect 164 254 165 255
rect 163 254 164 255
rect 162 254 163 255
rect 161 254 162 255
rect 76 254 77 255
rect 75 254 76 255
rect 74 254 75 255
rect 73 254 74 255
rect 72 254 73 255
rect 61 254 62 255
rect 60 254 61 255
rect 59 254 60 255
rect 58 254 59 255
rect 57 254 58 255
rect 56 254 57 255
rect 27 254 28 255
rect 26 254 27 255
rect 25 254 26 255
rect 24 254 25 255
rect 23 254 24 255
rect 22 254 23 255
rect 21 254 22 255
rect 20 254 21 255
rect 19 254 20 255
rect 195 255 196 256
rect 194 255 195 256
rect 193 255 194 256
rect 192 255 193 256
rect 191 255 192 256
rect 190 255 191 256
rect 189 255 190 256
rect 188 255 189 256
rect 187 255 188 256
rect 186 255 187 256
rect 181 255 182 256
rect 180 255 181 256
rect 179 255 180 256
rect 178 255 179 256
rect 170 255 171 256
rect 169 255 170 256
rect 168 255 169 256
rect 167 255 168 256
rect 166 255 167 256
rect 163 255 164 256
rect 162 255 163 256
rect 161 255 162 256
rect 76 255 77 256
rect 75 255 76 256
rect 74 255 75 256
rect 73 255 74 256
rect 72 255 73 256
rect 71 255 72 256
rect 70 255 71 256
rect 63 255 64 256
rect 62 255 63 256
rect 61 255 62 256
rect 60 255 61 256
rect 59 255 60 256
rect 58 255 59 256
rect 57 255 58 256
rect 27 255 28 256
rect 26 255 27 256
rect 25 255 26 256
rect 24 255 25 256
rect 23 255 24 256
rect 22 255 23 256
rect 21 255 22 256
rect 20 255 21 256
rect 19 255 20 256
rect 18 255 19 256
rect 17 255 18 256
rect 16 255 17 256
rect 15 255 16 256
rect 14 255 15 256
rect 195 256 196 257
rect 194 256 195 257
rect 193 256 194 257
rect 192 256 193 257
rect 191 256 192 257
rect 190 256 191 257
rect 189 256 190 257
rect 188 256 189 257
rect 187 256 188 257
rect 186 256 187 257
rect 181 256 182 257
rect 180 256 181 257
rect 179 256 180 257
rect 178 256 179 257
rect 171 256 172 257
rect 170 256 171 257
rect 169 256 170 257
rect 168 256 169 257
rect 163 256 164 257
rect 162 256 163 257
rect 161 256 162 257
rect 76 256 77 257
rect 75 256 76 257
rect 74 256 75 257
rect 73 256 74 257
rect 72 256 73 257
rect 71 256 72 257
rect 70 256 71 257
rect 69 256 70 257
rect 68 256 69 257
rect 67 256 68 257
rect 66 256 67 257
rect 65 256 66 257
rect 64 256 65 257
rect 63 256 64 257
rect 62 256 63 257
rect 61 256 62 257
rect 60 256 61 257
rect 59 256 60 257
rect 58 256 59 257
rect 57 256 58 257
rect 24 256 25 257
rect 23 256 24 257
rect 22 256 23 257
rect 21 256 22 257
rect 20 256 21 257
rect 19 256 20 257
rect 18 256 19 257
rect 17 256 18 257
rect 16 256 17 257
rect 15 256 16 257
rect 14 256 15 257
rect 13 256 14 257
rect 12 256 13 257
rect 194 257 195 258
rect 193 257 194 258
rect 192 257 193 258
rect 191 257 192 258
rect 190 257 191 258
rect 189 257 190 258
rect 188 257 189 258
rect 187 257 188 258
rect 186 257 187 258
rect 181 257 182 258
rect 180 257 181 258
rect 179 257 180 258
rect 178 257 179 258
rect 171 257 172 258
rect 170 257 171 258
rect 169 257 170 258
rect 168 257 169 258
rect 163 257 164 258
rect 162 257 163 258
rect 161 257 162 258
rect 75 257 76 258
rect 74 257 75 258
rect 73 257 74 258
rect 72 257 73 258
rect 71 257 72 258
rect 70 257 71 258
rect 69 257 70 258
rect 68 257 69 258
rect 67 257 68 258
rect 66 257 67 258
rect 65 257 66 258
rect 64 257 65 258
rect 63 257 64 258
rect 62 257 63 258
rect 61 257 62 258
rect 60 257 61 258
rect 59 257 60 258
rect 58 257 59 258
rect 18 257 19 258
rect 17 257 18 258
rect 16 257 17 258
rect 15 257 16 258
rect 14 257 15 258
rect 13 257 14 258
rect 12 257 13 258
rect 181 258 182 259
rect 180 258 181 259
rect 179 258 180 259
rect 178 258 179 259
rect 172 258 173 259
rect 171 258 172 259
rect 170 258 171 259
rect 169 258 170 259
rect 163 258 164 259
rect 162 258 163 259
rect 161 258 162 259
rect 74 258 75 259
rect 73 258 74 259
rect 72 258 73 259
rect 71 258 72 259
rect 70 258 71 259
rect 69 258 70 259
rect 68 258 69 259
rect 67 258 68 259
rect 66 258 67 259
rect 65 258 66 259
rect 64 258 65 259
rect 63 258 64 259
rect 62 258 63 259
rect 61 258 62 259
rect 60 258 61 259
rect 59 258 60 259
rect 27 258 28 259
rect 26 258 27 259
rect 25 258 26 259
rect 24 258 25 259
rect 23 258 24 259
rect 22 258 23 259
rect 21 258 22 259
rect 20 258 21 259
rect 19 258 20 259
rect 18 258 19 259
rect 17 258 18 259
rect 16 258 17 259
rect 15 258 16 259
rect 14 258 15 259
rect 13 258 14 259
rect 12 258 13 259
rect 181 259 182 260
rect 180 259 181 260
rect 179 259 180 260
rect 178 259 179 260
rect 171 259 172 260
rect 170 259 171 260
rect 167 259 168 260
rect 166 259 167 260
rect 165 259 166 260
rect 164 259 165 260
rect 163 259 164 260
rect 162 259 163 260
rect 161 259 162 260
rect 73 259 74 260
rect 72 259 73 260
rect 71 259 72 260
rect 70 259 71 260
rect 69 259 70 260
rect 68 259 69 260
rect 67 259 68 260
rect 66 259 67 260
rect 65 259 66 260
rect 64 259 65 260
rect 63 259 64 260
rect 62 259 63 260
rect 61 259 62 260
rect 60 259 61 260
rect 27 259 28 260
rect 26 259 27 260
rect 25 259 26 260
rect 24 259 25 260
rect 23 259 24 260
rect 22 259 23 260
rect 21 259 22 260
rect 20 259 21 260
rect 19 259 20 260
rect 18 259 19 260
rect 17 259 18 260
rect 16 259 17 260
rect 15 259 16 260
rect 14 259 15 260
rect 13 259 14 260
rect 12 259 13 260
rect 181 260 182 261
rect 180 260 181 261
rect 179 260 180 261
rect 178 260 179 261
rect 170 260 171 261
rect 167 260 168 261
rect 166 260 167 261
rect 165 260 166 261
rect 164 260 165 261
rect 71 260 72 261
rect 70 260 71 261
rect 69 260 70 261
rect 68 260 69 261
rect 67 260 68 261
rect 66 260 67 261
rect 65 260 66 261
rect 64 260 65 261
rect 63 260 64 261
rect 62 260 63 261
rect 61 260 62 261
rect 27 260 28 261
rect 26 260 27 261
rect 25 260 26 261
rect 24 260 25 261
rect 23 260 24 261
rect 22 260 23 261
rect 21 260 22 261
rect 20 260 21 261
rect 19 260 20 261
rect 18 260 19 261
rect 17 260 18 261
rect 16 260 17 261
rect 15 260 16 261
rect 14 260 15 261
rect 13 260 14 261
rect 187 261 188 262
rect 181 261 182 262
rect 180 261 181 262
rect 179 261 180 262
rect 178 261 179 262
rect 167 261 168 262
rect 166 261 167 262
rect 165 261 166 262
rect 164 261 165 262
rect 67 261 68 262
rect 66 261 67 262
rect 65 261 66 262
rect 27 261 28 262
rect 26 261 27 262
rect 25 261 26 262
rect 24 261 25 262
rect 23 261 24 262
rect 22 261 23 262
rect 21 261 22 262
rect 187 262 188 263
rect 181 262 182 263
rect 180 262 181 263
rect 179 262 180 263
rect 178 262 179 263
rect 167 262 168 263
rect 166 262 167 263
rect 165 262 166 263
rect 164 262 165 263
rect 25 262 26 263
rect 24 262 25 263
rect 23 262 24 263
rect 22 262 23 263
rect 21 262 22 263
rect 20 262 21 263
rect 19 262 20 263
rect 188 263 189 264
rect 187 263 188 264
rect 181 263 182 264
rect 180 263 181 264
rect 179 263 180 264
rect 178 263 179 264
rect 175 263 176 264
rect 174 263 175 264
rect 173 263 174 264
rect 172 263 173 264
rect 171 263 172 264
rect 170 263 171 264
rect 169 263 170 264
rect 168 263 169 264
rect 167 263 168 264
rect 166 263 167 264
rect 165 263 166 264
rect 164 263 165 264
rect 163 263 164 264
rect 162 263 163 264
rect 161 263 162 264
rect 160 263 161 264
rect 110 263 111 264
rect 109 263 110 264
rect 108 263 109 264
rect 107 263 108 264
rect 106 263 107 264
rect 105 263 106 264
rect 104 263 105 264
rect 103 263 104 264
rect 102 263 103 264
rect 101 263 102 264
rect 100 263 101 264
rect 23 263 24 264
rect 22 263 23 264
rect 21 263 22 264
rect 20 263 21 264
rect 19 263 20 264
rect 18 263 19 264
rect 17 263 18 264
rect 195 264 196 265
rect 194 264 195 265
rect 193 264 194 265
rect 192 264 193 265
rect 191 264 192 265
rect 190 264 191 265
rect 189 264 190 265
rect 188 264 189 265
rect 187 264 188 265
rect 181 264 182 265
rect 180 264 181 265
rect 179 264 180 265
rect 178 264 179 265
rect 175 264 176 265
rect 174 264 175 265
rect 173 264 174 265
rect 172 264 173 265
rect 171 264 172 265
rect 170 264 171 265
rect 169 264 170 265
rect 168 264 169 265
rect 167 264 168 265
rect 166 264 167 265
rect 165 264 166 265
rect 164 264 165 265
rect 163 264 164 265
rect 162 264 163 265
rect 161 264 162 265
rect 160 264 161 265
rect 110 264 111 265
rect 109 264 110 265
rect 108 264 109 265
rect 107 264 108 265
rect 106 264 107 265
rect 105 264 106 265
rect 104 264 105 265
rect 103 264 104 265
rect 102 264 103 265
rect 101 264 102 265
rect 100 264 101 265
rect 71 264 72 265
rect 70 264 71 265
rect 69 264 70 265
rect 68 264 69 265
rect 67 264 68 265
rect 66 264 67 265
rect 65 264 66 265
rect 64 264 65 265
rect 63 264 64 265
rect 62 264 63 265
rect 27 264 28 265
rect 20 264 21 265
rect 19 264 20 265
rect 18 264 19 265
rect 17 264 18 265
rect 16 264 17 265
rect 15 264 16 265
rect 194 265 195 266
rect 193 265 194 266
rect 192 265 193 266
rect 191 265 192 266
rect 190 265 191 266
rect 189 265 190 266
rect 188 265 189 266
rect 187 265 188 266
rect 181 265 182 266
rect 180 265 181 266
rect 179 265 180 266
rect 178 265 179 266
rect 175 265 176 266
rect 174 265 175 266
rect 173 265 174 266
rect 172 265 173 266
rect 171 265 172 266
rect 170 265 171 266
rect 169 265 170 266
rect 168 265 169 266
rect 167 265 168 266
rect 166 265 167 266
rect 165 265 166 266
rect 164 265 165 266
rect 163 265 164 266
rect 162 265 163 266
rect 161 265 162 266
rect 160 265 161 266
rect 110 265 111 266
rect 109 265 110 266
rect 108 265 109 266
rect 107 265 108 266
rect 106 265 107 266
rect 105 265 106 266
rect 104 265 105 266
rect 103 265 104 266
rect 102 265 103 266
rect 101 265 102 266
rect 100 265 101 266
rect 73 265 74 266
rect 72 265 73 266
rect 71 265 72 266
rect 70 265 71 266
rect 69 265 70 266
rect 68 265 69 266
rect 67 265 68 266
rect 66 265 67 266
rect 65 265 66 266
rect 64 265 65 266
rect 63 265 64 266
rect 62 265 63 266
rect 61 265 62 266
rect 60 265 61 266
rect 27 265 28 266
rect 26 265 27 266
rect 25 265 26 266
rect 24 265 25 266
rect 23 265 24 266
rect 22 265 23 266
rect 18 265 19 266
rect 17 265 18 266
rect 16 265 17 266
rect 15 265 16 266
rect 14 265 15 266
rect 13 265 14 266
rect 187 266 188 267
rect 181 266 182 267
rect 180 266 181 267
rect 179 266 180 267
rect 178 266 179 267
rect 175 266 176 267
rect 174 266 175 267
rect 173 266 174 267
rect 172 266 173 267
rect 171 266 172 267
rect 170 266 171 267
rect 169 266 170 267
rect 168 266 169 267
rect 167 266 168 267
rect 166 266 167 267
rect 165 266 166 267
rect 164 266 165 267
rect 163 266 164 267
rect 162 266 163 267
rect 161 266 162 267
rect 160 266 161 267
rect 110 266 111 267
rect 109 266 110 267
rect 108 266 109 267
rect 107 266 108 267
rect 106 266 107 267
rect 105 266 106 267
rect 104 266 105 267
rect 103 266 104 267
rect 102 266 103 267
rect 101 266 102 267
rect 100 266 101 267
rect 74 266 75 267
rect 73 266 74 267
rect 72 266 73 267
rect 71 266 72 267
rect 70 266 71 267
rect 69 266 70 267
rect 68 266 69 267
rect 67 266 68 267
rect 66 266 67 267
rect 65 266 66 267
rect 64 266 65 267
rect 63 266 64 267
rect 62 266 63 267
rect 61 266 62 267
rect 60 266 61 267
rect 59 266 60 267
rect 27 266 28 267
rect 26 266 27 267
rect 25 266 26 267
rect 24 266 25 267
rect 23 266 24 267
rect 22 266 23 267
rect 21 266 22 267
rect 20 266 21 267
rect 19 266 20 267
rect 18 266 19 267
rect 17 266 18 267
rect 16 266 17 267
rect 15 266 16 267
rect 14 266 15 267
rect 13 266 14 267
rect 12 266 13 267
rect 193 267 194 268
rect 192 267 193 268
rect 191 267 192 268
rect 190 267 191 268
rect 187 267 188 268
rect 180 267 181 268
rect 179 267 180 268
rect 110 267 111 268
rect 109 267 110 268
rect 108 267 109 268
rect 107 267 108 268
rect 106 267 107 268
rect 105 267 106 268
rect 104 267 105 268
rect 103 267 104 268
rect 102 267 103 268
rect 101 267 102 268
rect 100 267 101 268
rect 75 267 76 268
rect 74 267 75 268
rect 73 267 74 268
rect 72 267 73 268
rect 71 267 72 268
rect 70 267 71 268
rect 69 267 70 268
rect 68 267 69 268
rect 67 267 68 268
rect 66 267 67 268
rect 65 267 66 268
rect 64 267 65 268
rect 63 267 64 268
rect 62 267 63 268
rect 61 267 62 268
rect 60 267 61 268
rect 59 267 60 268
rect 58 267 59 268
rect 26 267 27 268
rect 25 267 26 268
rect 24 267 25 268
rect 23 267 24 268
rect 22 267 23 268
rect 21 267 22 268
rect 20 267 21 268
rect 19 267 20 268
rect 18 267 19 268
rect 17 267 18 268
rect 16 267 17 268
rect 15 267 16 268
rect 14 267 15 268
rect 13 267 14 268
rect 12 267 13 268
rect 194 268 195 269
rect 193 268 194 269
rect 192 268 193 269
rect 191 268 192 269
rect 190 268 191 269
rect 189 268 190 269
rect 110 268 111 269
rect 109 268 110 269
rect 108 268 109 269
rect 107 268 108 269
rect 106 268 107 269
rect 105 268 106 269
rect 104 268 105 269
rect 103 268 104 269
rect 102 268 103 269
rect 101 268 102 269
rect 100 268 101 269
rect 75 268 76 269
rect 74 268 75 269
rect 73 268 74 269
rect 72 268 73 269
rect 71 268 72 269
rect 70 268 71 269
rect 69 268 70 269
rect 68 268 69 269
rect 67 268 68 269
rect 66 268 67 269
rect 65 268 66 269
rect 64 268 65 269
rect 63 268 64 269
rect 62 268 63 269
rect 61 268 62 269
rect 60 268 61 269
rect 59 268 60 269
rect 58 268 59 269
rect 21 268 22 269
rect 20 268 21 269
rect 19 268 20 269
rect 18 268 19 269
rect 17 268 18 269
rect 16 268 17 269
rect 15 268 16 269
rect 14 268 15 269
rect 13 268 14 269
rect 12 268 13 269
rect 195 269 196 270
rect 194 269 195 270
rect 193 269 194 270
rect 192 269 193 270
rect 191 269 192 270
rect 190 269 191 270
rect 189 269 190 270
rect 110 269 111 270
rect 109 269 110 270
rect 108 269 109 270
rect 107 269 108 270
rect 106 269 107 270
rect 105 269 106 270
rect 104 269 105 270
rect 103 269 104 270
rect 102 269 103 270
rect 101 269 102 270
rect 100 269 101 270
rect 76 269 77 270
rect 75 269 76 270
rect 74 269 75 270
rect 73 269 74 270
rect 72 269 73 270
rect 71 269 72 270
rect 70 269 71 270
rect 69 269 70 270
rect 68 269 69 270
rect 67 269 68 270
rect 66 269 67 270
rect 65 269 66 270
rect 64 269 65 270
rect 63 269 64 270
rect 62 269 63 270
rect 61 269 62 270
rect 60 269 61 270
rect 59 269 60 270
rect 58 269 59 270
rect 57 269 58 270
rect 16 269 17 270
rect 15 269 16 270
rect 14 269 15 270
rect 13 269 14 270
rect 12 269 13 270
rect 195 270 196 271
rect 194 270 195 271
rect 192 270 193 271
rect 190 270 191 271
rect 189 270 190 271
rect 110 270 111 271
rect 109 270 110 271
rect 108 270 109 271
rect 107 270 108 271
rect 106 270 107 271
rect 105 270 106 271
rect 104 270 105 271
rect 103 270 104 271
rect 102 270 103 271
rect 101 270 102 271
rect 100 270 101 271
rect 76 270 77 271
rect 75 270 76 271
rect 74 270 75 271
rect 73 270 74 271
rect 72 270 73 271
rect 68 270 69 271
rect 67 270 68 271
rect 66 270 67 271
rect 65 270 66 271
rect 61 270 62 271
rect 60 270 61 271
rect 59 270 60 271
rect 58 270 59 271
rect 57 270 58 271
rect 31 270 32 271
rect 30 270 31 271
rect 195 271 196 272
rect 194 271 195 272
rect 192 271 193 272
rect 191 271 192 272
rect 190 271 191 272
rect 189 271 190 272
rect 110 271 111 272
rect 109 271 110 272
rect 108 271 109 272
rect 107 271 108 272
rect 106 271 107 272
rect 105 271 106 272
rect 104 271 105 272
rect 103 271 104 272
rect 102 271 103 272
rect 101 271 102 272
rect 100 271 101 272
rect 76 271 77 272
rect 75 271 76 272
rect 74 271 75 272
rect 73 271 74 272
rect 72 271 73 272
rect 68 271 69 272
rect 67 271 68 272
rect 66 271 67 272
rect 65 271 66 272
rect 60 271 61 272
rect 59 271 60 272
rect 58 271 59 272
rect 57 271 58 272
rect 56 271 57 272
rect 31 271 32 272
rect 30 271 31 272
rect 17 271 18 272
rect 194 272 195 273
rect 192 272 193 273
rect 191 272 192 273
rect 190 272 191 273
rect 110 272 111 273
rect 109 272 110 273
rect 108 272 109 273
rect 107 272 108 273
rect 106 272 107 273
rect 105 272 106 273
rect 104 272 105 273
rect 103 272 104 273
rect 102 272 103 273
rect 101 272 102 273
rect 100 272 101 273
rect 76 272 77 273
rect 75 272 76 273
rect 74 272 75 273
rect 73 272 74 273
rect 68 272 69 273
rect 67 272 68 273
rect 66 272 67 273
rect 65 272 66 273
rect 60 272 61 273
rect 59 272 60 273
rect 58 272 59 273
rect 57 272 58 273
rect 56 272 57 273
rect 31 272 32 273
rect 30 272 31 273
rect 29 272 30 273
rect 23 272 24 273
rect 22 272 23 273
rect 21 272 22 273
rect 20 272 21 273
rect 19 272 20 273
rect 18 272 19 273
rect 17 272 18 273
rect 16 272 17 273
rect 110 273 111 274
rect 109 273 110 274
rect 108 273 109 274
rect 107 273 108 274
rect 106 273 107 274
rect 105 273 106 274
rect 104 273 105 274
rect 103 273 104 274
rect 102 273 103 274
rect 101 273 102 274
rect 100 273 101 274
rect 76 273 77 274
rect 75 273 76 274
rect 74 273 75 274
rect 73 273 74 274
rect 68 273 69 274
rect 67 273 68 274
rect 66 273 67 274
rect 65 273 66 274
rect 60 273 61 274
rect 59 273 60 274
rect 58 273 59 274
rect 57 273 58 274
rect 56 273 57 274
rect 31 273 32 274
rect 30 273 31 274
rect 29 273 30 274
rect 28 273 29 274
rect 27 273 28 274
rect 26 273 27 274
rect 25 273 26 274
rect 24 273 25 274
rect 23 273 24 274
rect 22 273 23 274
rect 21 273 22 274
rect 20 273 21 274
rect 19 273 20 274
rect 18 273 19 274
rect 17 273 18 274
rect 16 273 17 274
rect 194 274 195 275
rect 193 274 194 275
rect 192 274 193 275
rect 191 274 192 275
rect 190 274 191 275
rect 189 274 190 275
rect 188 274 189 275
rect 187 274 188 275
rect 186 274 187 275
rect 110 274 111 275
rect 109 274 110 275
rect 108 274 109 275
rect 107 274 108 275
rect 106 274 107 275
rect 105 274 106 275
rect 104 274 105 275
rect 103 274 104 275
rect 102 274 103 275
rect 101 274 102 275
rect 100 274 101 275
rect 76 274 77 275
rect 75 274 76 275
rect 74 274 75 275
rect 73 274 74 275
rect 68 274 69 275
rect 67 274 68 275
rect 66 274 67 275
rect 65 274 66 275
rect 60 274 61 275
rect 59 274 60 275
rect 58 274 59 275
rect 57 274 58 275
rect 56 274 57 275
rect 30 274 31 275
rect 29 274 30 275
rect 28 274 29 275
rect 27 274 28 275
rect 26 274 27 275
rect 25 274 26 275
rect 24 274 25 275
rect 23 274 24 275
rect 22 274 23 275
rect 21 274 22 275
rect 20 274 21 275
rect 19 274 20 275
rect 18 274 19 275
rect 17 274 18 275
rect 194 275 195 276
rect 193 275 194 276
rect 192 275 193 276
rect 191 275 192 276
rect 190 275 191 276
rect 189 275 190 276
rect 188 275 189 276
rect 187 275 188 276
rect 186 275 187 276
rect 110 275 111 276
rect 109 275 110 276
rect 108 275 109 276
rect 107 275 108 276
rect 106 275 107 276
rect 105 275 106 276
rect 104 275 105 276
rect 103 275 104 276
rect 102 275 103 276
rect 101 275 102 276
rect 100 275 101 276
rect 76 275 77 276
rect 75 275 76 276
rect 74 275 75 276
rect 73 275 74 276
rect 68 275 69 276
rect 67 275 68 276
rect 66 275 67 276
rect 65 275 66 276
rect 60 275 61 276
rect 59 275 60 276
rect 58 275 59 276
rect 57 275 58 276
rect 29 275 30 276
rect 28 275 29 276
rect 27 275 28 276
rect 26 275 27 276
rect 25 275 26 276
rect 24 275 25 276
rect 23 275 24 276
rect 110 276 111 277
rect 109 276 110 277
rect 108 276 109 277
rect 107 276 108 277
rect 106 276 107 277
rect 105 276 106 277
rect 104 276 105 277
rect 103 276 104 277
rect 102 276 103 277
rect 101 276 102 277
rect 100 276 101 277
rect 76 276 77 277
rect 75 276 76 277
rect 74 276 75 277
rect 73 276 74 277
rect 72 276 73 277
rect 71 276 72 277
rect 68 276 69 277
rect 67 276 68 277
rect 66 276 67 277
rect 65 276 66 277
rect 62 276 63 277
rect 61 276 62 277
rect 60 276 61 277
rect 59 276 60 277
rect 58 276 59 277
rect 57 276 58 277
rect 27 276 28 277
rect 26 276 27 277
rect 25 276 26 277
rect 24 276 25 277
rect 23 276 24 277
rect 22 276 23 277
rect 194 277 195 278
rect 193 277 194 278
rect 192 277 193 278
rect 191 277 192 278
rect 190 277 191 278
rect 110 277 111 278
rect 109 277 110 278
rect 108 277 109 278
rect 107 277 108 278
rect 106 277 107 278
rect 105 277 106 278
rect 104 277 105 278
rect 103 277 104 278
rect 102 277 103 278
rect 101 277 102 278
rect 100 277 101 278
rect 76 277 77 278
rect 75 277 76 278
rect 74 277 75 278
rect 73 277 74 278
rect 72 277 73 278
rect 71 277 72 278
rect 70 277 71 278
rect 68 277 69 278
rect 67 277 68 278
rect 66 277 67 278
rect 65 277 66 278
rect 64 277 65 278
rect 63 277 64 278
rect 62 277 63 278
rect 61 277 62 278
rect 60 277 61 278
rect 59 277 60 278
rect 58 277 59 278
rect 57 277 58 278
rect 26 277 27 278
rect 25 277 26 278
rect 24 277 25 278
rect 23 277 24 278
rect 22 277 23 278
rect 21 277 22 278
rect 20 277 21 278
rect 194 278 195 279
rect 193 278 194 279
rect 192 278 193 279
rect 191 278 192 279
rect 190 278 191 279
rect 189 278 190 279
rect 176 278 177 279
rect 110 278 111 279
rect 109 278 110 279
rect 108 278 109 279
rect 107 278 108 279
rect 106 278 107 279
rect 105 278 106 279
rect 104 278 105 279
rect 103 278 104 279
rect 102 278 103 279
rect 101 278 102 279
rect 100 278 101 279
rect 75 278 76 279
rect 74 278 75 279
rect 73 278 74 279
rect 72 278 73 279
rect 71 278 72 279
rect 68 278 69 279
rect 67 278 68 279
rect 66 278 67 279
rect 65 278 66 279
rect 64 278 65 279
rect 63 278 64 279
rect 62 278 63 279
rect 61 278 62 279
rect 60 278 61 279
rect 59 278 60 279
rect 58 278 59 279
rect 24 278 25 279
rect 23 278 24 279
rect 22 278 23 279
rect 21 278 22 279
rect 20 278 21 279
rect 19 278 20 279
rect 18 278 19 279
rect 195 279 196 280
rect 194 279 195 280
rect 192 279 193 280
rect 191 279 192 280
rect 190 279 191 280
rect 189 279 190 280
rect 177 279 178 280
rect 176 279 177 280
rect 175 279 176 280
rect 164 279 165 280
rect 110 279 111 280
rect 109 279 110 280
rect 108 279 109 280
rect 107 279 108 280
rect 106 279 107 280
rect 105 279 106 280
rect 104 279 105 280
rect 103 279 104 280
rect 102 279 103 280
rect 101 279 102 280
rect 100 279 101 280
rect 75 279 76 280
rect 74 279 75 280
rect 73 279 74 280
rect 72 279 73 280
rect 71 279 72 280
rect 68 279 69 280
rect 67 279 68 280
rect 66 279 67 280
rect 65 279 66 280
rect 64 279 65 280
rect 63 279 64 280
rect 62 279 63 280
rect 61 279 62 280
rect 60 279 61 280
rect 59 279 60 280
rect 22 279 23 280
rect 21 279 22 280
rect 20 279 21 280
rect 19 279 20 280
rect 18 279 19 280
rect 17 279 18 280
rect 195 280 196 281
rect 194 280 195 281
rect 192 280 193 281
rect 190 280 191 281
rect 189 280 190 281
rect 177 280 178 281
rect 176 280 177 281
rect 175 280 176 281
rect 174 280 175 281
rect 164 280 165 281
rect 163 280 164 281
rect 162 280 163 281
rect 110 280 111 281
rect 109 280 110 281
rect 108 280 109 281
rect 107 280 108 281
rect 106 280 107 281
rect 105 280 106 281
rect 104 280 105 281
rect 103 280 104 281
rect 102 280 103 281
rect 101 280 102 281
rect 100 280 101 281
rect 74 280 75 281
rect 73 280 74 281
rect 72 280 73 281
rect 71 280 72 281
rect 68 280 69 281
rect 67 280 68 281
rect 66 280 67 281
rect 65 280 66 281
rect 64 280 65 281
rect 63 280 64 281
rect 62 280 63 281
rect 61 280 62 281
rect 60 280 61 281
rect 20 280 21 281
rect 19 280 20 281
rect 18 280 19 281
rect 17 280 18 281
rect 16 280 17 281
rect 194 281 195 282
rect 192 281 193 282
rect 191 281 192 282
rect 190 281 191 282
rect 189 281 190 282
rect 177 281 178 282
rect 176 281 177 282
rect 175 281 176 282
rect 174 281 175 282
rect 173 281 174 282
rect 164 281 165 282
rect 163 281 164 282
rect 162 281 163 282
rect 110 281 111 282
rect 109 281 110 282
rect 108 281 109 282
rect 107 281 108 282
rect 106 281 107 282
rect 105 281 106 282
rect 104 281 105 282
rect 103 281 104 282
rect 102 281 103 282
rect 101 281 102 282
rect 100 281 101 282
rect 72 281 73 282
rect 71 281 72 282
rect 68 281 69 282
rect 67 281 68 282
rect 66 281 67 282
rect 65 281 66 282
rect 64 281 65 282
rect 63 281 64 282
rect 62 281 63 282
rect 61 281 62 282
rect 18 281 19 282
rect 17 281 18 282
rect 16 281 17 282
rect 194 282 195 283
rect 192 282 193 283
rect 191 282 192 283
rect 190 282 191 283
rect 177 282 178 283
rect 176 282 177 283
rect 175 282 176 283
rect 174 282 175 283
rect 173 282 174 283
rect 172 282 173 283
rect 164 282 165 283
rect 163 282 164 283
rect 162 282 163 283
rect 110 282 111 283
rect 109 282 110 283
rect 108 282 109 283
rect 107 282 108 283
rect 106 282 107 283
rect 105 282 106 283
rect 104 282 105 283
rect 103 282 104 283
rect 102 282 103 283
rect 101 282 102 283
rect 100 282 101 283
rect 67 282 68 283
rect 66 282 67 283
rect 65 282 66 283
rect 193 283 194 284
rect 192 283 193 284
rect 191 283 192 284
rect 176 283 177 284
rect 175 283 176 284
rect 174 283 175 284
rect 173 283 174 284
rect 172 283 173 284
rect 171 283 172 284
rect 164 283 165 284
rect 163 283 164 284
rect 162 283 163 284
rect 110 283 111 284
rect 109 283 110 284
rect 108 283 109 284
rect 107 283 108 284
rect 106 283 107 284
rect 105 283 106 284
rect 104 283 105 284
rect 103 283 104 284
rect 102 283 103 284
rect 101 283 102 284
rect 100 283 101 284
rect 194 284 195 285
rect 193 284 194 285
rect 192 284 193 285
rect 191 284 192 285
rect 190 284 191 285
rect 189 284 190 285
rect 175 284 176 285
rect 174 284 175 285
rect 173 284 174 285
rect 172 284 173 285
rect 171 284 172 285
rect 170 284 171 285
rect 169 284 170 285
rect 168 284 169 285
rect 167 284 168 285
rect 164 284 165 285
rect 163 284 164 285
rect 162 284 163 285
rect 110 284 111 285
rect 109 284 110 285
rect 108 284 109 285
rect 107 284 108 285
rect 106 284 107 285
rect 105 284 106 285
rect 104 284 105 285
rect 103 284 104 285
rect 102 284 103 285
rect 101 284 102 285
rect 100 284 101 285
rect 194 285 195 286
rect 193 285 194 286
rect 192 285 193 286
rect 191 285 192 286
rect 190 285 191 286
rect 189 285 190 286
rect 174 285 175 286
rect 173 285 174 286
rect 172 285 173 286
rect 171 285 172 286
rect 170 285 171 286
rect 169 285 170 286
rect 168 285 169 286
rect 167 285 168 286
rect 166 285 167 286
rect 165 285 166 286
rect 164 285 165 286
rect 163 285 164 286
rect 162 285 163 286
rect 110 285 111 286
rect 109 285 110 286
rect 108 285 109 286
rect 107 285 108 286
rect 106 285 107 286
rect 105 285 106 286
rect 104 285 105 286
rect 103 285 104 286
rect 102 285 103 286
rect 101 285 102 286
rect 100 285 101 286
rect 195 286 196 287
rect 194 286 195 287
rect 190 286 191 287
rect 189 286 190 287
rect 172 286 173 287
rect 171 286 172 287
rect 170 286 171 287
rect 169 286 170 287
rect 168 286 169 287
rect 167 286 168 287
rect 166 286 167 287
rect 165 286 166 287
rect 164 286 165 287
rect 163 286 164 287
rect 162 286 163 287
rect 110 286 111 287
rect 109 286 110 287
rect 108 286 109 287
rect 107 286 108 287
rect 106 286 107 287
rect 105 286 106 287
rect 104 286 105 287
rect 103 286 104 287
rect 102 286 103 287
rect 101 286 102 287
rect 100 286 101 287
rect 195 287 196 288
rect 194 287 195 288
rect 190 287 191 288
rect 189 287 190 288
rect 172 287 173 288
rect 171 287 172 288
rect 170 287 171 288
rect 169 287 170 288
rect 168 287 169 288
rect 167 287 168 288
rect 166 287 167 288
rect 165 287 166 288
rect 164 287 165 288
rect 163 287 164 288
rect 162 287 163 288
rect 110 287 111 288
rect 109 287 110 288
rect 108 287 109 288
rect 107 287 108 288
rect 106 287 107 288
rect 105 287 106 288
rect 104 287 105 288
rect 103 287 104 288
rect 102 287 103 288
rect 101 287 102 288
rect 100 287 101 288
rect 194 288 195 289
rect 193 288 194 289
rect 191 288 192 289
rect 174 288 175 289
rect 173 288 174 289
rect 172 288 173 289
rect 171 288 172 289
rect 170 288 171 289
rect 169 288 170 289
rect 168 288 169 289
rect 167 288 168 289
rect 166 288 167 289
rect 165 288 166 289
rect 164 288 165 289
rect 163 288 164 289
rect 162 288 163 289
rect 110 288 111 289
rect 109 288 110 289
rect 108 288 109 289
rect 107 288 108 289
rect 106 288 107 289
rect 105 288 106 289
rect 104 288 105 289
rect 103 288 104 289
rect 102 288 103 289
rect 101 288 102 289
rect 100 288 101 289
rect 194 289 195 290
rect 193 289 194 290
rect 192 289 193 290
rect 191 289 192 290
rect 190 289 191 290
rect 175 289 176 290
rect 174 289 175 290
rect 173 289 174 290
rect 172 289 173 290
rect 171 289 172 290
rect 170 289 171 290
rect 169 289 170 290
rect 164 289 165 290
rect 163 289 164 290
rect 162 289 163 290
rect 110 289 111 290
rect 109 289 110 290
rect 108 289 109 290
rect 107 289 108 290
rect 106 289 107 290
rect 105 289 106 290
rect 104 289 105 290
rect 103 289 104 290
rect 102 289 103 290
rect 101 289 102 290
rect 100 289 101 290
rect 23 289 24 290
rect 22 289 23 290
rect 21 289 22 290
rect 20 289 21 290
rect 19 289 20 290
rect 194 290 195 291
rect 193 290 194 291
rect 192 290 193 291
rect 191 290 192 291
rect 190 290 191 291
rect 189 290 190 291
rect 175 290 176 291
rect 174 290 175 291
rect 173 290 174 291
rect 172 290 173 291
rect 171 290 172 291
rect 164 290 165 291
rect 163 290 164 291
rect 162 290 163 291
rect 147 290 148 291
rect 146 290 147 291
rect 145 290 146 291
rect 144 290 145 291
rect 143 290 144 291
rect 142 290 143 291
rect 141 290 142 291
rect 140 290 141 291
rect 139 290 140 291
rect 138 290 139 291
rect 137 290 138 291
rect 136 290 137 291
rect 135 290 136 291
rect 134 290 135 291
rect 133 290 134 291
rect 132 290 133 291
rect 131 290 132 291
rect 130 290 131 291
rect 129 290 130 291
rect 128 290 129 291
rect 127 290 128 291
rect 126 290 127 291
rect 125 290 126 291
rect 124 290 125 291
rect 123 290 124 291
rect 122 290 123 291
rect 121 290 122 291
rect 120 290 121 291
rect 119 290 120 291
rect 118 290 119 291
rect 117 290 118 291
rect 116 290 117 291
rect 115 290 116 291
rect 114 290 115 291
rect 113 290 114 291
rect 112 290 113 291
rect 111 290 112 291
rect 110 290 111 291
rect 109 290 110 291
rect 108 290 109 291
rect 107 290 108 291
rect 106 290 107 291
rect 105 290 106 291
rect 104 290 105 291
rect 103 290 104 291
rect 102 290 103 291
rect 101 290 102 291
rect 100 290 101 291
rect 25 290 26 291
rect 24 290 25 291
rect 23 290 24 291
rect 22 290 23 291
rect 21 290 22 291
rect 20 290 21 291
rect 19 290 20 291
rect 18 290 19 291
rect 17 290 18 291
rect 16 290 17 291
rect 195 291 196 292
rect 194 291 195 292
rect 190 291 191 292
rect 189 291 190 292
rect 176 291 177 292
rect 175 291 176 292
rect 174 291 175 292
rect 173 291 174 292
rect 164 291 165 292
rect 163 291 164 292
rect 162 291 163 292
rect 147 291 148 292
rect 146 291 147 292
rect 145 291 146 292
rect 144 291 145 292
rect 143 291 144 292
rect 142 291 143 292
rect 141 291 142 292
rect 140 291 141 292
rect 139 291 140 292
rect 138 291 139 292
rect 137 291 138 292
rect 136 291 137 292
rect 135 291 136 292
rect 134 291 135 292
rect 133 291 134 292
rect 132 291 133 292
rect 131 291 132 292
rect 130 291 131 292
rect 129 291 130 292
rect 128 291 129 292
rect 127 291 128 292
rect 126 291 127 292
rect 125 291 126 292
rect 124 291 125 292
rect 123 291 124 292
rect 122 291 123 292
rect 121 291 122 292
rect 120 291 121 292
rect 119 291 120 292
rect 118 291 119 292
rect 117 291 118 292
rect 116 291 117 292
rect 115 291 116 292
rect 114 291 115 292
rect 113 291 114 292
rect 112 291 113 292
rect 111 291 112 292
rect 110 291 111 292
rect 109 291 110 292
rect 108 291 109 292
rect 107 291 108 292
rect 106 291 107 292
rect 105 291 106 292
rect 104 291 105 292
rect 103 291 104 292
rect 102 291 103 292
rect 101 291 102 292
rect 100 291 101 292
rect 26 291 27 292
rect 25 291 26 292
rect 24 291 25 292
rect 23 291 24 292
rect 22 291 23 292
rect 21 291 22 292
rect 20 291 21 292
rect 19 291 20 292
rect 18 291 19 292
rect 17 291 18 292
rect 16 291 17 292
rect 15 291 16 292
rect 195 292 196 293
rect 194 292 195 293
rect 190 292 191 293
rect 189 292 190 293
rect 177 292 178 293
rect 176 292 177 293
rect 175 292 176 293
rect 174 292 175 293
rect 173 292 174 293
rect 164 292 165 293
rect 163 292 164 293
rect 162 292 163 293
rect 147 292 148 293
rect 146 292 147 293
rect 145 292 146 293
rect 144 292 145 293
rect 143 292 144 293
rect 142 292 143 293
rect 141 292 142 293
rect 140 292 141 293
rect 139 292 140 293
rect 138 292 139 293
rect 137 292 138 293
rect 136 292 137 293
rect 135 292 136 293
rect 134 292 135 293
rect 133 292 134 293
rect 132 292 133 293
rect 131 292 132 293
rect 130 292 131 293
rect 129 292 130 293
rect 128 292 129 293
rect 127 292 128 293
rect 126 292 127 293
rect 125 292 126 293
rect 124 292 125 293
rect 123 292 124 293
rect 122 292 123 293
rect 121 292 122 293
rect 120 292 121 293
rect 119 292 120 293
rect 118 292 119 293
rect 117 292 118 293
rect 116 292 117 293
rect 115 292 116 293
rect 114 292 115 293
rect 113 292 114 293
rect 112 292 113 293
rect 111 292 112 293
rect 110 292 111 293
rect 109 292 110 293
rect 108 292 109 293
rect 107 292 108 293
rect 106 292 107 293
rect 105 292 106 293
rect 104 292 105 293
rect 103 292 104 293
rect 102 292 103 293
rect 101 292 102 293
rect 100 292 101 293
rect 27 292 28 293
rect 26 292 27 293
rect 25 292 26 293
rect 24 292 25 293
rect 23 292 24 293
rect 22 292 23 293
rect 21 292 22 293
rect 20 292 21 293
rect 19 292 20 293
rect 18 292 19 293
rect 17 292 18 293
rect 16 292 17 293
rect 15 292 16 293
rect 14 292 15 293
rect 194 293 195 294
rect 193 293 194 294
rect 192 293 193 294
rect 191 293 192 294
rect 190 293 191 294
rect 189 293 190 294
rect 176 293 177 294
rect 175 293 176 294
rect 174 293 175 294
rect 164 293 165 294
rect 163 293 164 294
rect 162 293 163 294
rect 147 293 148 294
rect 146 293 147 294
rect 145 293 146 294
rect 144 293 145 294
rect 143 293 144 294
rect 142 293 143 294
rect 141 293 142 294
rect 140 293 141 294
rect 139 293 140 294
rect 138 293 139 294
rect 137 293 138 294
rect 136 293 137 294
rect 135 293 136 294
rect 134 293 135 294
rect 133 293 134 294
rect 132 293 133 294
rect 131 293 132 294
rect 130 293 131 294
rect 129 293 130 294
rect 128 293 129 294
rect 127 293 128 294
rect 126 293 127 294
rect 125 293 126 294
rect 124 293 125 294
rect 123 293 124 294
rect 122 293 123 294
rect 121 293 122 294
rect 120 293 121 294
rect 119 293 120 294
rect 118 293 119 294
rect 117 293 118 294
rect 116 293 117 294
rect 115 293 116 294
rect 114 293 115 294
rect 113 293 114 294
rect 112 293 113 294
rect 111 293 112 294
rect 110 293 111 294
rect 109 293 110 294
rect 108 293 109 294
rect 107 293 108 294
rect 106 293 107 294
rect 105 293 106 294
rect 104 293 105 294
rect 103 293 104 294
rect 102 293 103 294
rect 101 293 102 294
rect 100 293 101 294
rect 27 293 28 294
rect 26 293 27 294
rect 25 293 26 294
rect 24 293 25 294
rect 17 293 18 294
rect 16 293 17 294
rect 15 293 16 294
rect 14 293 15 294
rect 13 293 14 294
rect 194 294 195 295
rect 193 294 194 295
rect 192 294 193 295
rect 191 294 192 295
rect 190 294 191 295
rect 175 294 176 295
rect 147 294 148 295
rect 146 294 147 295
rect 145 294 146 295
rect 144 294 145 295
rect 143 294 144 295
rect 142 294 143 295
rect 141 294 142 295
rect 140 294 141 295
rect 139 294 140 295
rect 138 294 139 295
rect 137 294 138 295
rect 136 294 137 295
rect 135 294 136 295
rect 134 294 135 295
rect 133 294 134 295
rect 132 294 133 295
rect 131 294 132 295
rect 130 294 131 295
rect 129 294 130 295
rect 128 294 129 295
rect 127 294 128 295
rect 126 294 127 295
rect 125 294 126 295
rect 124 294 125 295
rect 123 294 124 295
rect 122 294 123 295
rect 121 294 122 295
rect 120 294 121 295
rect 119 294 120 295
rect 118 294 119 295
rect 117 294 118 295
rect 116 294 117 295
rect 115 294 116 295
rect 114 294 115 295
rect 113 294 114 295
rect 112 294 113 295
rect 111 294 112 295
rect 110 294 111 295
rect 109 294 110 295
rect 108 294 109 295
rect 107 294 108 295
rect 106 294 107 295
rect 105 294 106 295
rect 104 294 105 295
rect 103 294 104 295
rect 102 294 103 295
rect 101 294 102 295
rect 100 294 101 295
rect 27 294 28 295
rect 26 294 27 295
rect 25 294 26 295
rect 15 294 16 295
rect 14 294 15 295
rect 13 294 14 295
rect 192 295 193 296
rect 147 295 148 296
rect 146 295 147 296
rect 145 295 146 296
rect 144 295 145 296
rect 143 295 144 296
rect 142 295 143 296
rect 141 295 142 296
rect 140 295 141 296
rect 139 295 140 296
rect 138 295 139 296
rect 137 295 138 296
rect 136 295 137 296
rect 135 295 136 296
rect 134 295 135 296
rect 133 295 134 296
rect 132 295 133 296
rect 131 295 132 296
rect 130 295 131 296
rect 129 295 130 296
rect 128 295 129 296
rect 127 295 128 296
rect 126 295 127 296
rect 125 295 126 296
rect 124 295 125 296
rect 123 295 124 296
rect 122 295 123 296
rect 121 295 122 296
rect 120 295 121 296
rect 119 295 120 296
rect 118 295 119 296
rect 117 295 118 296
rect 116 295 117 296
rect 115 295 116 296
rect 114 295 115 296
rect 113 295 114 296
rect 112 295 113 296
rect 111 295 112 296
rect 110 295 111 296
rect 109 295 110 296
rect 108 295 109 296
rect 107 295 108 296
rect 106 295 107 296
rect 105 295 106 296
rect 104 295 105 296
rect 103 295 104 296
rect 102 295 103 296
rect 101 295 102 296
rect 100 295 101 296
rect 27 295 28 296
rect 26 295 27 296
rect 25 295 26 296
rect 15 295 16 296
rect 14 295 15 296
rect 13 295 14 296
rect 12 295 13 296
rect 194 296 195 297
rect 193 296 194 297
rect 192 296 193 297
rect 191 296 192 297
rect 190 296 191 297
rect 189 296 190 297
rect 180 296 181 297
rect 179 296 180 297
rect 178 296 179 297
rect 177 296 178 297
rect 176 296 177 297
rect 175 296 176 297
rect 174 296 175 297
rect 173 296 174 297
rect 172 296 173 297
rect 171 296 172 297
rect 170 296 171 297
rect 169 296 170 297
rect 168 296 169 297
rect 167 296 168 297
rect 166 296 167 297
rect 165 296 166 297
rect 164 296 165 297
rect 163 296 164 297
rect 162 296 163 297
rect 161 296 162 297
rect 147 296 148 297
rect 146 296 147 297
rect 145 296 146 297
rect 144 296 145 297
rect 143 296 144 297
rect 142 296 143 297
rect 141 296 142 297
rect 140 296 141 297
rect 139 296 140 297
rect 138 296 139 297
rect 137 296 138 297
rect 136 296 137 297
rect 135 296 136 297
rect 134 296 135 297
rect 133 296 134 297
rect 132 296 133 297
rect 131 296 132 297
rect 130 296 131 297
rect 129 296 130 297
rect 128 296 129 297
rect 127 296 128 297
rect 126 296 127 297
rect 125 296 126 297
rect 124 296 125 297
rect 123 296 124 297
rect 122 296 123 297
rect 121 296 122 297
rect 120 296 121 297
rect 119 296 120 297
rect 118 296 119 297
rect 117 296 118 297
rect 116 296 117 297
rect 115 296 116 297
rect 114 296 115 297
rect 113 296 114 297
rect 112 296 113 297
rect 111 296 112 297
rect 110 296 111 297
rect 109 296 110 297
rect 108 296 109 297
rect 107 296 108 297
rect 106 296 107 297
rect 105 296 106 297
rect 104 296 105 297
rect 103 296 104 297
rect 102 296 103 297
rect 101 296 102 297
rect 100 296 101 297
rect 67 296 68 297
rect 66 296 67 297
rect 65 296 66 297
rect 27 296 28 297
rect 26 296 27 297
rect 25 296 26 297
rect 14 296 15 297
rect 13 296 14 297
rect 12 296 13 297
rect 195 297 196 298
rect 194 297 195 298
rect 193 297 194 298
rect 192 297 193 298
rect 191 297 192 298
rect 190 297 191 298
rect 189 297 190 298
rect 181 297 182 298
rect 180 297 181 298
rect 179 297 180 298
rect 178 297 179 298
rect 177 297 178 298
rect 176 297 177 298
rect 175 297 176 298
rect 174 297 175 298
rect 173 297 174 298
rect 172 297 173 298
rect 171 297 172 298
rect 170 297 171 298
rect 169 297 170 298
rect 168 297 169 298
rect 167 297 168 298
rect 166 297 167 298
rect 165 297 166 298
rect 164 297 165 298
rect 163 297 164 298
rect 162 297 163 298
rect 161 297 162 298
rect 160 297 161 298
rect 147 297 148 298
rect 146 297 147 298
rect 145 297 146 298
rect 144 297 145 298
rect 143 297 144 298
rect 142 297 143 298
rect 141 297 142 298
rect 140 297 141 298
rect 139 297 140 298
rect 138 297 139 298
rect 137 297 138 298
rect 136 297 137 298
rect 135 297 136 298
rect 134 297 135 298
rect 133 297 134 298
rect 132 297 133 298
rect 131 297 132 298
rect 130 297 131 298
rect 129 297 130 298
rect 128 297 129 298
rect 127 297 128 298
rect 126 297 127 298
rect 125 297 126 298
rect 124 297 125 298
rect 123 297 124 298
rect 122 297 123 298
rect 121 297 122 298
rect 120 297 121 298
rect 119 297 120 298
rect 118 297 119 298
rect 117 297 118 298
rect 116 297 117 298
rect 115 297 116 298
rect 114 297 115 298
rect 113 297 114 298
rect 112 297 113 298
rect 111 297 112 298
rect 110 297 111 298
rect 109 297 110 298
rect 108 297 109 298
rect 107 297 108 298
rect 106 297 107 298
rect 105 297 106 298
rect 104 297 105 298
rect 103 297 104 298
rect 102 297 103 298
rect 101 297 102 298
rect 100 297 101 298
rect 73 297 74 298
rect 72 297 73 298
rect 71 297 72 298
rect 70 297 71 298
rect 69 297 70 298
rect 68 297 69 298
rect 67 297 68 298
rect 66 297 67 298
rect 65 297 66 298
rect 64 297 65 298
rect 63 297 64 298
rect 62 297 63 298
rect 61 297 62 298
rect 60 297 61 298
rect 59 297 60 298
rect 27 297 28 298
rect 26 297 27 298
rect 25 297 26 298
rect 14 297 15 298
rect 13 297 14 298
rect 12 297 13 298
rect 190 298 191 299
rect 189 298 190 299
rect 181 298 182 299
rect 180 298 181 299
rect 179 298 180 299
rect 178 298 179 299
rect 177 298 178 299
rect 176 298 177 299
rect 175 298 176 299
rect 174 298 175 299
rect 173 298 174 299
rect 172 298 173 299
rect 171 298 172 299
rect 170 298 171 299
rect 169 298 170 299
rect 168 298 169 299
rect 167 298 168 299
rect 166 298 167 299
rect 165 298 166 299
rect 164 298 165 299
rect 163 298 164 299
rect 162 298 163 299
rect 161 298 162 299
rect 160 298 161 299
rect 147 298 148 299
rect 146 298 147 299
rect 145 298 146 299
rect 144 298 145 299
rect 143 298 144 299
rect 142 298 143 299
rect 141 298 142 299
rect 140 298 141 299
rect 139 298 140 299
rect 138 298 139 299
rect 137 298 138 299
rect 136 298 137 299
rect 135 298 136 299
rect 134 298 135 299
rect 133 298 134 299
rect 132 298 133 299
rect 131 298 132 299
rect 130 298 131 299
rect 129 298 130 299
rect 128 298 129 299
rect 127 298 128 299
rect 126 298 127 299
rect 125 298 126 299
rect 124 298 125 299
rect 123 298 124 299
rect 122 298 123 299
rect 121 298 122 299
rect 120 298 121 299
rect 119 298 120 299
rect 118 298 119 299
rect 117 298 118 299
rect 116 298 117 299
rect 115 298 116 299
rect 114 298 115 299
rect 113 298 114 299
rect 112 298 113 299
rect 111 298 112 299
rect 110 298 111 299
rect 109 298 110 299
rect 108 298 109 299
rect 107 298 108 299
rect 106 298 107 299
rect 105 298 106 299
rect 104 298 105 299
rect 103 298 104 299
rect 102 298 103 299
rect 101 298 102 299
rect 100 298 101 299
rect 76 298 77 299
rect 75 298 76 299
rect 74 298 75 299
rect 73 298 74 299
rect 72 298 73 299
rect 71 298 72 299
rect 70 298 71 299
rect 69 298 70 299
rect 68 298 69 299
rect 67 298 68 299
rect 66 298 67 299
rect 65 298 66 299
rect 64 298 65 299
rect 63 298 64 299
rect 62 298 63 299
rect 61 298 62 299
rect 60 298 61 299
rect 59 298 60 299
rect 58 298 59 299
rect 57 298 58 299
rect 56 298 57 299
rect 27 298 28 299
rect 26 298 27 299
rect 25 298 26 299
rect 24 298 25 299
rect 14 298 15 299
rect 13 298 14 299
rect 12 298 13 299
rect 190 299 191 300
rect 189 299 190 300
rect 181 299 182 300
rect 180 299 181 300
rect 179 299 180 300
rect 178 299 179 300
rect 177 299 178 300
rect 176 299 177 300
rect 175 299 176 300
rect 174 299 175 300
rect 173 299 174 300
rect 172 299 173 300
rect 171 299 172 300
rect 170 299 171 300
rect 169 299 170 300
rect 168 299 169 300
rect 167 299 168 300
rect 166 299 167 300
rect 165 299 166 300
rect 164 299 165 300
rect 163 299 164 300
rect 162 299 163 300
rect 161 299 162 300
rect 160 299 161 300
rect 147 299 148 300
rect 146 299 147 300
rect 145 299 146 300
rect 144 299 145 300
rect 143 299 144 300
rect 142 299 143 300
rect 141 299 142 300
rect 140 299 141 300
rect 139 299 140 300
rect 138 299 139 300
rect 137 299 138 300
rect 136 299 137 300
rect 135 299 136 300
rect 134 299 135 300
rect 133 299 134 300
rect 132 299 133 300
rect 131 299 132 300
rect 130 299 131 300
rect 129 299 130 300
rect 128 299 129 300
rect 127 299 128 300
rect 126 299 127 300
rect 125 299 126 300
rect 124 299 125 300
rect 123 299 124 300
rect 122 299 123 300
rect 121 299 122 300
rect 120 299 121 300
rect 119 299 120 300
rect 118 299 119 300
rect 117 299 118 300
rect 116 299 117 300
rect 115 299 116 300
rect 114 299 115 300
rect 113 299 114 300
rect 112 299 113 300
rect 111 299 112 300
rect 110 299 111 300
rect 109 299 110 300
rect 108 299 109 300
rect 107 299 108 300
rect 106 299 107 300
rect 105 299 106 300
rect 104 299 105 300
rect 103 299 104 300
rect 102 299 103 300
rect 101 299 102 300
rect 100 299 101 300
rect 79 299 80 300
rect 78 299 79 300
rect 77 299 78 300
rect 76 299 77 300
rect 75 299 76 300
rect 74 299 75 300
rect 73 299 74 300
rect 72 299 73 300
rect 71 299 72 300
rect 70 299 71 300
rect 69 299 70 300
rect 68 299 69 300
rect 67 299 68 300
rect 66 299 67 300
rect 65 299 66 300
rect 64 299 65 300
rect 63 299 64 300
rect 62 299 63 300
rect 61 299 62 300
rect 60 299 61 300
rect 59 299 60 300
rect 58 299 59 300
rect 57 299 58 300
rect 56 299 57 300
rect 55 299 56 300
rect 54 299 55 300
rect 26 299 27 300
rect 25 299 26 300
rect 24 299 25 300
rect 23 299 24 300
rect 15 299 16 300
rect 14 299 15 300
rect 13 299 14 300
rect 12 299 13 300
rect 195 300 196 301
rect 194 300 195 301
rect 193 300 194 301
rect 192 300 193 301
rect 191 300 192 301
rect 190 300 191 301
rect 189 300 190 301
rect 171 300 172 301
rect 170 300 171 301
rect 169 300 170 301
rect 168 300 169 301
rect 147 300 148 301
rect 146 300 147 301
rect 145 300 146 301
rect 144 300 145 301
rect 143 300 144 301
rect 142 300 143 301
rect 141 300 142 301
rect 140 300 141 301
rect 139 300 140 301
rect 138 300 139 301
rect 137 300 138 301
rect 136 300 137 301
rect 135 300 136 301
rect 134 300 135 301
rect 133 300 134 301
rect 132 300 133 301
rect 131 300 132 301
rect 130 300 131 301
rect 129 300 130 301
rect 128 300 129 301
rect 127 300 128 301
rect 126 300 127 301
rect 125 300 126 301
rect 124 300 125 301
rect 123 300 124 301
rect 122 300 123 301
rect 121 300 122 301
rect 120 300 121 301
rect 119 300 120 301
rect 118 300 119 301
rect 117 300 118 301
rect 116 300 117 301
rect 115 300 116 301
rect 114 300 115 301
rect 113 300 114 301
rect 112 300 113 301
rect 111 300 112 301
rect 110 300 111 301
rect 109 300 110 301
rect 108 300 109 301
rect 107 300 108 301
rect 106 300 107 301
rect 105 300 106 301
rect 104 300 105 301
rect 103 300 104 301
rect 102 300 103 301
rect 101 300 102 301
rect 100 300 101 301
rect 80 300 81 301
rect 79 300 80 301
rect 78 300 79 301
rect 77 300 78 301
rect 76 300 77 301
rect 75 300 76 301
rect 74 300 75 301
rect 73 300 74 301
rect 72 300 73 301
rect 71 300 72 301
rect 70 300 71 301
rect 69 300 70 301
rect 68 300 69 301
rect 67 300 68 301
rect 66 300 67 301
rect 65 300 66 301
rect 64 300 65 301
rect 63 300 64 301
rect 62 300 63 301
rect 61 300 62 301
rect 60 300 61 301
rect 59 300 60 301
rect 58 300 59 301
rect 57 300 58 301
rect 56 300 57 301
rect 55 300 56 301
rect 54 300 55 301
rect 53 300 54 301
rect 52 300 53 301
rect 25 300 26 301
rect 24 300 25 301
rect 23 300 24 301
rect 17 300 18 301
rect 16 300 17 301
rect 15 300 16 301
rect 14 300 15 301
rect 13 300 14 301
rect 194 301 195 302
rect 193 301 194 302
rect 192 301 193 302
rect 191 301 192 302
rect 190 301 191 302
rect 189 301 190 302
rect 171 301 172 302
rect 170 301 171 302
rect 169 301 170 302
rect 168 301 169 302
rect 147 301 148 302
rect 146 301 147 302
rect 145 301 146 302
rect 144 301 145 302
rect 143 301 144 302
rect 142 301 143 302
rect 141 301 142 302
rect 140 301 141 302
rect 139 301 140 302
rect 138 301 139 302
rect 137 301 138 302
rect 136 301 137 302
rect 135 301 136 302
rect 134 301 135 302
rect 133 301 134 302
rect 132 301 133 302
rect 131 301 132 302
rect 130 301 131 302
rect 129 301 130 302
rect 128 301 129 302
rect 127 301 128 302
rect 126 301 127 302
rect 125 301 126 302
rect 124 301 125 302
rect 123 301 124 302
rect 122 301 123 302
rect 121 301 122 302
rect 120 301 121 302
rect 119 301 120 302
rect 118 301 119 302
rect 117 301 118 302
rect 116 301 117 302
rect 115 301 116 302
rect 114 301 115 302
rect 113 301 114 302
rect 112 301 113 302
rect 111 301 112 302
rect 110 301 111 302
rect 109 301 110 302
rect 108 301 109 302
rect 107 301 108 302
rect 106 301 107 302
rect 105 301 106 302
rect 104 301 105 302
rect 103 301 104 302
rect 102 301 103 302
rect 101 301 102 302
rect 100 301 101 302
rect 82 301 83 302
rect 81 301 82 302
rect 80 301 81 302
rect 79 301 80 302
rect 78 301 79 302
rect 77 301 78 302
rect 76 301 77 302
rect 75 301 76 302
rect 74 301 75 302
rect 73 301 74 302
rect 72 301 73 302
rect 71 301 72 302
rect 70 301 71 302
rect 69 301 70 302
rect 68 301 69 302
rect 67 301 68 302
rect 66 301 67 302
rect 65 301 66 302
rect 64 301 65 302
rect 63 301 64 302
rect 62 301 63 302
rect 61 301 62 302
rect 60 301 61 302
rect 59 301 60 302
rect 58 301 59 302
rect 57 301 58 302
rect 56 301 57 302
rect 55 301 56 302
rect 54 301 55 302
rect 53 301 54 302
rect 52 301 53 302
rect 51 301 52 302
rect 24 301 25 302
rect 23 301 24 302
rect 17 301 18 302
rect 16 301 17 302
rect 15 301 16 302
rect 14 301 15 302
rect 190 302 191 303
rect 189 302 190 303
rect 171 302 172 303
rect 170 302 171 303
rect 169 302 170 303
rect 168 302 169 303
rect 147 302 148 303
rect 146 302 147 303
rect 145 302 146 303
rect 144 302 145 303
rect 143 302 144 303
rect 142 302 143 303
rect 141 302 142 303
rect 140 302 141 303
rect 139 302 140 303
rect 138 302 139 303
rect 137 302 138 303
rect 136 302 137 303
rect 135 302 136 303
rect 134 302 135 303
rect 133 302 134 303
rect 132 302 133 303
rect 131 302 132 303
rect 130 302 131 303
rect 129 302 130 303
rect 128 302 129 303
rect 127 302 128 303
rect 126 302 127 303
rect 125 302 126 303
rect 124 302 125 303
rect 123 302 124 303
rect 122 302 123 303
rect 121 302 122 303
rect 120 302 121 303
rect 119 302 120 303
rect 118 302 119 303
rect 117 302 118 303
rect 116 302 117 303
rect 115 302 116 303
rect 114 302 115 303
rect 113 302 114 303
rect 112 302 113 303
rect 111 302 112 303
rect 110 302 111 303
rect 109 302 110 303
rect 108 302 109 303
rect 107 302 108 303
rect 106 302 107 303
rect 105 302 106 303
rect 104 302 105 303
rect 103 302 104 303
rect 102 302 103 303
rect 101 302 102 303
rect 100 302 101 303
rect 83 302 84 303
rect 82 302 83 303
rect 81 302 82 303
rect 80 302 81 303
rect 79 302 80 303
rect 78 302 79 303
rect 77 302 78 303
rect 76 302 77 303
rect 75 302 76 303
rect 74 302 75 303
rect 73 302 74 303
rect 59 302 60 303
rect 58 302 59 303
rect 57 302 58 303
rect 56 302 57 303
rect 55 302 56 303
rect 54 302 55 303
rect 53 302 54 303
rect 52 302 53 303
rect 51 302 52 303
rect 50 302 51 303
rect 49 302 50 303
rect 16 302 17 303
rect 15 302 16 303
rect 194 303 195 304
rect 193 303 194 304
rect 192 303 193 304
rect 191 303 192 304
rect 190 303 191 304
rect 189 303 190 304
rect 170 303 171 304
rect 169 303 170 304
rect 147 303 148 304
rect 146 303 147 304
rect 145 303 146 304
rect 144 303 145 304
rect 143 303 144 304
rect 142 303 143 304
rect 141 303 142 304
rect 140 303 141 304
rect 139 303 140 304
rect 138 303 139 304
rect 137 303 138 304
rect 136 303 137 304
rect 135 303 136 304
rect 134 303 135 304
rect 133 303 134 304
rect 132 303 133 304
rect 131 303 132 304
rect 130 303 131 304
rect 129 303 130 304
rect 128 303 129 304
rect 127 303 128 304
rect 126 303 127 304
rect 125 303 126 304
rect 124 303 125 304
rect 123 303 124 304
rect 122 303 123 304
rect 121 303 122 304
rect 120 303 121 304
rect 119 303 120 304
rect 118 303 119 304
rect 117 303 118 304
rect 116 303 117 304
rect 115 303 116 304
rect 114 303 115 304
rect 113 303 114 304
rect 112 303 113 304
rect 111 303 112 304
rect 110 303 111 304
rect 109 303 110 304
rect 108 303 109 304
rect 107 303 108 304
rect 106 303 107 304
rect 105 303 106 304
rect 104 303 105 304
rect 103 303 104 304
rect 102 303 103 304
rect 101 303 102 304
rect 100 303 101 304
rect 84 303 85 304
rect 83 303 84 304
rect 82 303 83 304
rect 81 303 82 304
rect 80 303 81 304
rect 79 303 80 304
rect 78 303 79 304
rect 55 303 56 304
rect 54 303 55 304
rect 53 303 54 304
rect 52 303 53 304
rect 51 303 52 304
rect 50 303 51 304
rect 49 303 50 304
rect 195 304 196 305
rect 194 304 195 305
rect 193 304 194 305
rect 192 304 193 305
rect 191 304 192 305
rect 190 304 191 305
rect 189 304 190 305
rect 147 304 148 305
rect 146 304 147 305
rect 145 304 146 305
rect 144 304 145 305
rect 143 304 144 305
rect 142 304 143 305
rect 141 304 142 305
rect 140 304 141 305
rect 139 304 140 305
rect 138 304 139 305
rect 137 304 138 305
rect 136 304 137 305
rect 135 304 136 305
rect 134 304 135 305
rect 133 304 134 305
rect 132 304 133 305
rect 131 304 132 305
rect 130 304 131 305
rect 129 304 130 305
rect 128 304 129 305
rect 127 304 128 305
rect 126 304 127 305
rect 125 304 126 305
rect 124 304 125 305
rect 123 304 124 305
rect 122 304 123 305
rect 121 304 122 305
rect 120 304 121 305
rect 119 304 120 305
rect 118 304 119 305
rect 117 304 118 305
rect 116 304 117 305
rect 115 304 116 305
rect 114 304 115 305
rect 113 304 114 305
rect 112 304 113 305
rect 111 304 112 305
rect 110 304 111 305
rect 109 304 110 305
rect 108 304 109 305
rect 107 304 108 305
rect 106 304 107 305
rect 105 304 106 305
rect 104 304 105 305
rect 103 304 104 305
rect 102 304 103 305
rect 101 304 102 305
rect 100 304 101 305
rect 84 304 85 305
rect 83 304 84 305
rect 82 304 83 305
rect 81 304 82 305
rect 80 304 81 305
rect 53 304 54 305
rect 52 304 53 305
rect 51 304 52 305
rect 50 304 51 305
rect 49 304 50 305
rect 27 304 28 305
rect 26 304 27 305
rect 25 304 26 305
rect 24 304 25 305
rect 23 304 24 305
rect 194 305 195 306
rect 193 305 194 306
rect 192 305 193 306
rect 191 305 192 306
rect 190 305 191 306
rect 147 305 148 306
rect 146 305 147 306
rect 145 305 146 306
rect 144 305 145 306
rect 143 305 144 306
rect 142 305 143 306
rect 141 305 142 306
rect 140 305 141 306
rect 139 305 140 306
rect 138 305 139 306
rect 137 305 138 306
rect 136 305 137 306
rect 135 305 136 306
rect 134 305 135 306
rect 133 305 134 306
rect 132 305 133 306
rect 131 305 132 306
rect 130 305 131 306
rect 129 305 130 306
rect 128 305 129 306
rect 127 305 128 306
rect 126 305 127 306
rect 125 305 126 306
rect 124 305 125 306
rect 123 305 124 306
rect 122 305 123 306
rect 121 305 122 306
rect 120 305 121 306
rect 119 305 120 306
rect 118 305 119 306
rect 117 305 118 306
rect 116 305 117 306
rect 115 305 116 306
rect 114 305 115 306
rect 113 305 114 306
rect 112 305 113 306
rect 111 305 112 306
rect 110 305 111 306
rect 109 305 110 306
rect 108 305 109 306
rect 107 305 108 306
rect 106 305 107 306
rect 105 305 106 306
rect 104 305 105 306
rect 103 305 104 306
rect 102 305 103 306
rect 101 305 102 306
rect 100 305 101 306
rect 84 305 85 306
rect 83 305 84 306
rect 50 305 51 306
rect 49 305 50 306
rect 27 305 28 306
rect 26 305 27 306
rect 25 305 26 306
rect 24 305 25 306
rect 23 305 24 306
rect 22 305 23 306
rect 21 305 22 306
rect 20 305 21 306
rect 19 305 20 306
rect 18 305 19 306
rect 194 306 195 307
rect 190 306 191 307
rect 147 306 148 307
rect 146 306 147 307
rect 145 306 146 307
rect 144 306 145 307
rect 143 306 144 307
rect 142 306 143 307
rect 141 306 142 307
rect 140 306 141 307
rect 139 306 140 307
rect 138 306 139 307
rect 137 306 138 307
rect 136 306 137 307
rect 135 306 136 307
rect 134 306 135 307
rect 133 306 134 307
rect 132 306 133 307
rect 131 306 132 307
rect 130 306 131 307
rect 129 306 130 307
rect 128 306 129 307
rect 127 306 128 307
rect 126 306 127 307
rect 125 306 126 307
rect 124 306 125 307
rect 123 306 124 307
rect 122 306 123 307
rect 121 306 122 307
rect 120 306 121 307
rect 119 306 120 307
rect 118 306 119 307
rect 117 306 118 307
rect 116 306 117 307
rect 115 306 116 307
rect 114 306 115 307
rect 113 306 114 307
rect 112 306 113 307
rect 111 306 112 307
rect 110 306 111 307
rect 109 306 110 307
rect 108 306 109 307
rect 107 306 108 307
rect 106 306 107 307
rect 105 306 106 307
rect 104 306 105 307
rect 103 306 104 307
rect 102 306 103 307
rect 101 306 102 307
rect 100 306 101 307
rect 27 306 28 307
rect 26 306 27 307
rect 25 306 26 307
rect 24 306 25 307
rect 23 306 24 307
rect 22 306 23 307
rect 21 306 22 307
rect 20 306 21 307
rect 19 306 20 307
rect 18 306 19 307
rect 17 306 18 307
rect 16 306 17 307
rect 15 306 16 307
rect 14 306 15 307
rect 13 306 14 307
rect 195 307 196 308
rect 194 307 195 308
rect 193 307 194 308
rect 192 307 193 308
rect 191 307 192 308
rect 190 307 191 308
rect 189 307 190 308
rect 147 307 148 308
rect 146 307 147 308
rect 145 307 146 308
rect 144 307 145 308
rect 143 307 144 308
rect 142 307 143 308
rect 141 307 142 308
rect 140 307 141 308
rect 139 307 140 308
rect 138 307 139 308
rect 137 307 138 308
rect 136 307 137 308
rect 135 307 136 308
rect 134 307 135 308
rect 133 307 134 308
rect 132 307 133 308
rect 131 307 132 308
rect 130 307 131 308
rect 129 307 130 308
rect 128 307 129 308
rect 127 307 128 308
rect 126 307 127 308
rect 125 307 126 308
rect 124 307 125 308
rect 123 307 124 308
rect 122 307 123 308
rect 121 307 122 308
rect 120 307 121 308
rect 119 307 120 308
rect 118 307 119 308
rect 117 307 118 308
rect 116 307 117 308
rect 115 307 116 308
rect 114 307 115 308
rect 113 307 114 308
rect 112 307 113 308
rect 111 307 112 308
rect 110 307 111 308
rect 109 307 110 308
rect 108 307 109 308
rect 107 307 108 308
rect 106 307 107 308
rect 105 307 106 308
rect 104 307 105 308
rect 103 307 104 308
rect 102 307 103 308
rect 101 307 102 308
rect 100 307 101 308
rect 23 307 24 308
rect 22 307 23 308
rect 21 307 22 308
rect 20 307 21 308
rect 19 307 20 308
rect 18 307 19 308
rect 17 307 18 308
rect 16 307 17 308
rect 15 307 16 308
rect 14 307 15 308
rect 13 307 14 308
rect 12 307 13 308
rect 194 308 195 309
rect 193 308 194 309
rect 192 308 193 309
rect 191 308 192 309
rect 190 308 191 309
rect 189 308 190 309
rect 147 308 148 309
rect 146 308 147 309
rect 145 308 146 309
rect 144 308 145 309
rect 143 308 144 309
rect 142 308 143 309
rect 141 308 142 309
rect 140 308 141 309
rect 139 308 140 309
rect 138 308 139 309
rect 137 308 138 309
rect 136 308 137 309
rect 135 308 136 309
rect 134 308 135 309
rect 133 308 134 309
rect 132 308 133 309
rect 131 308 132 309
rect 130 308 131 309
rect 129 308 130 309
rect 128 308 129 309
rect 127 308 128 309
rect 126 308 127 309
rect 125 308 126 309
rect 124 308 125 309
rect 123 308 124 309
rect 122 308 123 309
rect 121 308 122 309
rect 120 308 121 309
rect 119 308 120 309
rect 118 308 119 309
rect 117 308 118 309
rect 116 308 117 309
rect 115 308 116 309
rect 114 308 115 309
rect 113 308 114 309
rect 112 308 113 309
rect 111 308 112 309
rect 110 308 111 309
rect 109 308 110 309
rect 108 308 109 309
rect 107 308 108 309
rect 106 308 107 309
rect 105 308 106 309
rect 104 308 105 309
rect 103 308 104 309
rect 102 308 103 309
rect 101 308 102 309
rect 100 308 101 309
rect 19 308 20 309
rect 18 308 19 309
rect 17 308 18 309
rect 16 308 17 309
rect 15 308 16 309
rect 14 308 15 309
rect 13 308 14 309
rect 12 308 13 309
rect 190 309 191 310
rect 189 309 190 310
rect 147 309 148 310
rect 146 309 147 310
rect 145 309 146 310
rect 144 309 145 310
rect 143 309 144 310
rect 142 309 143 310
rect 141 309 142 310
rect 140 309 141 310
rect 139 309 140 310
rect 138 309 139 310
rect 137 309 138 310
rect 136 309 137 310
rect 135 309 136 310
rect 134 309 135 310
rect 133 309 134 310
rect 132 309 133 310
rect 131 309 132 310
rect 130 309 131 310
rect 129 309 130 310
rect 128 309 129 310
rect 127 309 128 310
rect 126 309 127 310
rect 125 309 126 310
rect 124 309 125 310
rect 123 309 124 310
rect 122 309 123 310
rect 121 309 122 310
rect 120 309 121 310
rect 119 309 120 310
rect 118 309 119 310
rect 117 309 118 310
rect 116 309 117 310
rect 115 309 116 310
rect 114 309 115 310
rect 113 309 114 310
rect 112 309 113 310
rect 111 309 112 310
rect 110 309 111 310
rect 109 309 110 310
rect 108 309 109 310
rect 107 309 108 310
rect 106 309 107 310
rect 105 309 106 310
rect 104 309 105 310
rect 103 309 104 310
rect 102 309 103 310
rect 101 309 102 310
rect 100 309 101 310
rect 18 309 19 310
rect 17 309 18 310
rect 14 309 15 310
rect 13 309 14 310
rect 194 310 195 311
rect 193 310 194 311
rect 192 310 193 311
rect 191 310 192 311
rect 190 310 191 311
rect 189 310 190 311
rect 147 310 148 311
rect 146 310 147 311
rect 145 310 146 311
rect 144 310 145 311
rect 143 310 144 311
rect 142 310 143 311
rect 141 310 142 311
rect 140 310 141 311
rect 139 310 140 311
rect 138 310 139 311
rect 137 310 138 311
rect 136 310 137 311
rect 135 310 136 311
rect 134 310 135 311
rect 133 310 134 311
rect 132 310 133 311
rect 131 310 132 311
rect 130 310 131 311
rect 129 310 130 311
rect 128 310 129 311
rect 127 310 128 311
rect 126 310 127 311
rect 125 310 126 311
rect 124 310 125 311
rect 123 310 124 311
rect 122 310 123 311
rect 121 310 122 311
rect 120 310 121 311
rect 119 310 120 311
rect 118 310 119 311
rect 117 310 118 311
rect 116 310 117 311
rect 115 310 116 311
rect 114 310 115 311
rect 113 310 114 311
rect 112 310 113 311
rect 111 310 112 311
rect 110 310 111 311
rect 109 310 110 311
rect 108 310 109 311
rect 107 310 108 311
rect 106 310 107 311
rect 105 310 106 311
rect 104 310 105 311
rect 103 310 104 311
rect 102 310 103 311
rect 101 310 102 311
rect 100 310 101 311
rect 76 310 77 311
rect 75 310 76 311
rect 74 310 75 311
rect 73 310 74 311
rect 72 310 73 311
rect 71 310 72 311
rect 70 310 71 311
rect 69 310 70 311
rect 68 310 69 311
rect 67 310 68 311
rect 66 310 67 311
rect 65 310 66 311
rect 64 310 65 311
rect 63 310 64 311
rect 62 310 63 311
rect 61 310 62 311
rect 60 310 61 311
rect 59 310 60 311
rect 58 310 59 311
rect 57 310 58 311
rect 56 310 57 311
rect 55 310 56 311
rect 54 310 55 311
rect 53 310 54 311
rect 52 310 53 311
rect 51 310 52 311
rect 50 310 51 311
rect 49 310 50 311
rect 18 310 19 311
rect 17 310 18 311
rect 195 311 196 312
rect 194 311 195 312
rect 193 311 194 312
rect 192 311 193 312
rect 191 311 192 312
rect 190 311 191 312
rect 189 311 190 312
rect 147 311 148 312
rect 146 311 147 312
rect 145 311 146 312
rect 144 311 145 312
rect 143 311 144 312
rect 142 311 143 312
rect 141 311 142 312
rect 140 311 141 312
rect 139 311 140 312
rect 138 311 139 312
rect 137 311 138 312
rect 136 311 137 312
rect 135 311 136 312
rect 134 311 135 312
rect 133 311 134 312
rect 132 311 133 312
rect 131 311 132 312
rect 130 311 131 312
rect 129 311 130 312
rect 128 311 129 312
rect 127 311 128 312
rect 126 311 127 312
rect 125 311 126 312
rect 124 311 125 312
rect 123 311 124 312
rect 122 311 123 312
rect 121 311 122 312
rect 120 311 121 312
rect 119 311 120 312
rect 118 311 119 312
rect 117 311 118 312
rect 116 311 117 312
rect 115 311 116 312
rect 114 311 115 312
rect 113 311 114 312
rect 112 311 113 312
rect 111 311 112 312
rect 110 311 111 312
rect 109 311 110 312
rect 108 311 109 312
rect 107 311 108 312
rect 106 311 107 312
rect 105 311 106 312
rect 104 311 105 312
rect 103 311 104 312
rect 102 311 103 312
rect 101 311 102 312
rect 100 311 101 312
rect 76 311 77 312
rect 75 311 76 312
rect 74 311 75 312
rect 73 311 74 312
rect 72 311 73 312
rect 71 311 72 312
rect 70 311 71 312
rect 69 311 70 312
rect 68 311 69 312
rect 67 311 68 312
rect 66 311 67 312
rect 65 311 66 312
rect 64 311 65 312
rect 63 311 64 312
rect 62 311 63 312
rect 61 311 62 312
rect 60 311 61 312
rect 59 311 60 312
rect 58 311 59 312
rect 57 311 58 312
rect 56 311 57 312
rect 55 311 56 312
rect 54 311 55 312
rect 53 311 54 312
rect 52 311 53 312
rect 51 311 52 312
rect 50 311 51 312
rect 49 311 50 312
rect 27 311 28 312
rect 26 311 27 312
rect 25 311 26 312
rect 24 311 25 312
rect 23 311 24 312
rect 18 311 19 312
rect 17 311 18 312
rect 16 311 17 312
rect 190 312 191 313
rect 189 312 190 313
rect 172 312 173 313
rect 147 312 148 313
rect 146 312 147 313
rect 145 312 146 313
rect 144 312 145 313
rect 143 312 144 313
rect 142 312 143 313
rect 141 312 142 313
rect 140 312 141 313
rect 139 312 140 313
rect 138 312 139 313
rect 137 312 138 313
rect 136 312 137 313
rect 135 312 136 313
rect 134 312 135 313
rect 133 312 134 313
rect 132 312 133 313
rect 131 312 132 313
rect 130 312 131 313
rect 129 312 130 313
rect 128 312 129 313
rect 127 312 128 313
rect 126 312 127 313
rect 125 312 126 313
rect 124 312 125 313
rect 123 312 124 313
rect 122 312 123 313
rect 121 312 122 313
rect 120 312 121 313
rect 119 312 120 313
rect 118 312 119 313
rect 117 312 118 313
rect 116 312 117 313
rect 115 312 116 313
rect 114 312 115 313
rect 113 312 114 313
rect 112 312 113 313
rect 111 312 112 313
rect 110 312 111 313
rect 109 312 110 313
rect 108 312 109 313
rect 107 312 108 313
rect 106 312 107 313
rect 105 312 106 313
rect 104 312 105 313
rect 103 312 104 313
rect 102 312 103 313
rect 101 312 102 313
rect 100 312 101 313
rect 76 312 77 313
rect 75 312 76 313
rect 74 312 75 313
rect 73 312 74 313
rect 72 312 73 313
rect 71 312 72 313
rect 70 312 71 313
rect 69 312 70 313
rect 68 312 69 313
rect 67 312 68 313
rect 66 312 67 313
rect 65 312 66 313
rect 64 312 65 313
rect 63 312 64 313
rect 62 312 63 313
rect 61 312 62 313
rect 60 312 61 313
rect 59 312 60 313
rect 58 312 59 313
rect 57 312 58 313
rect 56 312 57 313
rect 55 312 56 313
rect 54 312 55 313
rect 53 312 54 313
rect 52 312 53 313
rect 51 312 52 313
rect 50 312 51 313
rect 49 312 50 313
rect 27 312 28 313
rect 26 312 27 313
rect 25 312 26 313
rect 24 312 25 313
rect 23 312 24 313
rect 22 312 23 313
rect 21 312 22 313
rect 20 312 21 313
rect 19 312 20 313
rect 18 312 19 313
rect 17 312 18 313
rect 16 312 17 313
rect 190 313 191 314
rect 189 313 190 314
rect 173 313 174 314
rect 172 313 173 314
rect 171 313 172 314
rect 147 313 148 314
rect 146 313 147 314
rect 145 313 146 314
rect 144 313 145 314
rect 143 313 144 314
rect 142 313 143 314
rect 141 313 142 314
rect 140 313 141 314
rect 139 313 140 314
rect 138 313 139 314
rect 137 313 138 314
rect 136 313 137 314
rect 135 313 136 314
rect 134 313 135 314
rect 133 313 134 314
rect 132 313 133 314
rect 131 313 132 314
rect 130 313 131 314
rect 129 313 130 314
rect 128 313 129 314
rect 127 313 128 314
rect 126 313 127 314
rect 125 313 126 314
rect 124 313 125 314
rect 123 313 124 314
rect 122 313 123 314
rect 121 313 122 314
rect 120 313 121 314
rect 119 313 120 314
rect 118 313 119 314
rect 117 313 118 314
rect 116 313 117 314
rect 115 313 116 314
rect 114 313 115 314
rect 113 313 114 314
rect 112 313 113 314
rect 111 313 112 314
rect 110 313 111 314
rect 109 313 110 314
rect 108 313 109 314
rect 107 313 108 314
rect 106 313 107 314
rect 105 313 106 314
rect 104 313 105 314
rect 103 313 104 314
rect 102 313 103 314
rect 101 313 102 314
rect 100 313 101 314
rect 76 313 77 314
rect 75 313 76 314
rect 74 313 75 314
rect 73 313 74 314
rect 72 313 73 314
rect 71 313 72 314
rect 70 313 71 314
rect 69 313 70 314
rect 68 313 69 314
rect 67 313 68 314
rect 66 313 67 314
rect 65 313 66 314
rect 64 313 65 314
rect 63 313 64 314
rect 62 313 63 314
rect 61 313 62 314
rect 60 313 61 314
rect 59 313 60 314
rect 58 313 59 314
rect 57 313 58 314
rect 56 313 57 314
rect 55 313 56 314
rect 54 313 55 314
rect 53 313 54 314
rect 52 313 53 314
rect 51 313 52 314
rect 50 313 51 314
rect 49 313 50 314
rect 27 313 28 314
rect 26 313 27 314
rect 25 313 26 314
rect 24 313 25 314
rect 23 313 24 314
rect 22 313 23 314
rect 21 313 22 314
rect 20 313 21 314
rect 19 313 20 314
rect 18 313 19 314
rect 17 313 18 314
rect 16 313 17 314
rect 194 314 195 315
rect 193 314 194 315
rect 192 314 193 315
rect 191 314 192 315
rect 190 314 191 315
rect 189 314 190 315
rect 173 314 174 315
rect 172 314 173 315
rect 171 314 172 315
rect 110 314 111 315
rect 109 314 110 315
rect 108 314 109 315
rect 107 314 108 315
rect 106 314 107 315
rect 105 314 106 315
rect 104 314 105 315
rect 103 314 104 315
rect 102 314 103 315
rect 101 314 102 315
rect 100 314 101 315
rect 76 314 77 315
rect 75 314 76 315
rect 74 314 75 315
rect 73 314 74 315
rect 72 314 73 315
rect 71 314 72 315
rect 70 314 71 315
rect 69 314 70 315
rect 68 314 69 315
rect 67 314 68 315
rect 66 314 67 315
rect 65 314 66 315
rect 64 314 65 315
rect 63 314 64 315
rect 62 314 63 315
rect 61 314 62 315
rect 60 314 61 315
rect 59 314 60 315
rect 58 314 59 315
rect 57 314 58 315
rect 56 314 57 315
rect 55 314 56 315
rect 54 314 55 315
rect 53 314 54 315
rect 52 314 53 315
rect 51 314 52 315
rect 50 314 51 315
rect 49 314 50 315
rect 24 314 25 315
rect 23 314 24 315
rect 22 314 23 315
rect 21 314 22 315
rect 20 314 21 315
rect 19 314 20 315
rect 18 314 19 315
rect 17 314 18 315
rect 194 315 195 316
rect 193 315 194 316
rect 192 315 193 316
rect 191 315 192 316
rect 190 315 191 316
rect 179 315 180 316
rect 178 315 179 316
rect 177 315 178 316
rect 173 315 174 316
rect 172 315 173 316
rect 171 315 172 316
rect 110 315 111 316
rect 109 315 110 316
rect 108 315 109 316
rect 107 315 108 316
rect 106 315 107 316
rect 105 315 106 316
rect 104 315 105 316
rect 103 315 104 316
rect 102 315 103 316
rect 101 315 102 316
rect 100 315 101 316
rect 76 315 77 316
rect 75 315 76 316
rect 74 315 75 316
rect 73 315 74 316
rect 72 315 73 316
rect 71 315 72 316
rect 70 315 71 316
rect 69 315 70 316
rect 68 315 69 316
rect 67 315 68 316
rect 66 315 67 316
rect 65 315 66 316
rect 64 315 65 316
rect 63 315 64 316
rect 62 315 63 316
rect 61 315 62 316
rect 60 315 61 316
rect 59 315 60 316
rect 58 315 59 316
rect 57 315 58 316
rect 56 315 57 316
rect 55 315 56 316
rect 54 315 55 316
rect 53 315 54 316
rect 52 315 53 316
rect 51 315 52 316
rect 50 315 51 316
rect 49 315 50 316
rect 19 315 20 316
rect 180 316 181 317
rect 179 316 180 317
rect 178 316 179 317
rect 177 316 178 317
rect 176 316 177 317
rect 173 316 174 317
rect 172 316 173 317
rect 171 316 172 317
rect 169 316 170 317
rect 168 316 169 317
rect 167 316 168 317
rect 166 316 167 317
rect 165 316 166 317
rect 164 316 165 317
rect 163 316 164 317
rect 162 316 163 317
rect 161 316 162 317
rect 160 316 161 317
rect 110 316 111 317
rect 109 316 110 317
rect 108 316 109 317
rect 107 316 108 317
rect 106 316 107 317
rect 105 316 106 317
rect 104 316 105 317
rect 103 316 104 317
rect 102 316 103 317
rect 101 316 102 317
rect 100 316 101 317
rect 64 316 65 317
rect 63 316 64 317
rect 62 316 63 317
rect 61 316 62 317
rect 60 316 61 317
rect 53 316 54 317
rect 52 316 53 317
rect 51 316 52 317
rect 50 316 51 317
rect 49 316 50 317
rect 194 317 195 318
rect 193 317 194 318
rect 192 317 193 318
rect 191 317 192 318
rect 190 317 191 318
rect 189 317 190 318
rect 180 317 181 318
rect 179 317 180 318
rect 178 317 179 318
rect 177 317 178 318
rect 176 317 177 318
rect 175 317 176 318
rect 173 317 174 318
rect 172 317 173 318
rect 171 317 172 318
rect 169 317 170 318
rect 168 317 169 318
rect 167 317 168 318
rect 166 317 167 318
rect 165 317 166 318
rect 164 317 165 318
rect 163 317 164 318
rect 162 317 163 318
rect 161 317 162 318
rect 160 317 161 318
rect 110 317 111 318
rect 109 317 110 318
rect 108 317 109 318
rect 107 317 108 318
rect 106 317 107 318
rect 105 317 106 318
rect 104 317 105 318
rect 103 317 104 318
rect 102 317 103 318
rect 101 317 102 318
rect 100 317 101 318
rect 64 317 65 318
rect 63 317 64 318
rect 62 317 63 318
rect 61 317 62 318
rect 60 317 61 318
rect 53 317 54 318
rect 52 317 53 318
rect 51 317 52 318
rect 50 317 51 318
rect 49 317 50 318
rect 27 317 28 318
rect 26 317 27 318
rect 25 317 26 318
rect 24 317 25 318
rect 23 317 24 318
rect 195 318 196 319
rect 194 318 195 319
rect 193 318 194 319
rect 192 318 193 319
rect 191 318 192 319
rect 190 318 191 319
rect 189 318 190 319
rect 181 318 182 319
rect 180 318 181 319
rect 179 318 180 319
rect 178 318 179 319
rect 177 318 178 319
rect 176 318 177 319
rect 175 318 176 319
rect 173 318 174 319
rect 172 318 173 319
rect 171 318 172 319
rect 169 318 170 319
rect 168 318 169 319
rect 167 318 168 319
rect 166 318 167 319
rect 165 318 166 319
rect 164 318 165 319
rect 163 318 164 319
rect 162 318 163 319
rect 161 318 162 319
rect 160 318 161 319
rect 110 318 111 319
rect 109 318 110 319
rect 108 318 109 319
rect 107 318 108 319
rect 106 318 107 319
rect 105 318 106 319
rect 104 318 105 319
rect 103 318 104 319
rect 102 318 103 319
rect 101 318 102 319
rect 100 318 101 319
rect 64 318 65 319
rect 63 318 64 319
rect 62 318 63 319
rect 61 318 62 319
rect 60 318 61 319
rect 53 318 54 319
rect 52 318 53 319
rect 51 318 52 319
rect 50 318 51 319
rect 49 318 50 319
rect 27 318 28 319
rect 26 318 27 319
rect 25 318 26 319
rect 24 318 25 319
rect 23 318 24 319
rect 22 318 23 319
rect 21 318 22 319
rect 20 318 21 319
rect 19 318 20 319
rect 18 318 19 319
rect 194 319 195 320
rect 181 319 182 320
rect 180 319 181 320
rect 179 319 180 320
rect 178 319 179 320
rect 177 319 178 320
rect 176 319 177 320
rect 175 319 176 320
rect 173 319 174 320
rect 172 319 173 320
rect 171 319 172 320
rect 169 319 170 320
rect 168 319 169 320
rect 167 319 168 320
rect 166 319 167 320
rect 165 319 166 320
rect 164 319 165 320
rect 163 319 164 320
rect 162 319 163 320
rect 161 319 162 320
rect 160 319 161 320
rect 110 319 111 320
rect 109 319 110 320
rect 108 319 109 320
rect 107 319 108 320
rect 106 319 107 320
rect 105 319 106 320
rect 104 319 105 320
rect 103 319 104 320
rect 102 319 103 320
rect 101 319 102 320
rect 100 319 101 320
rect 64 319 65 320
rect 63 319 64 320
rect 62 319 63 320
rect 61 319 62 320
rect 60 319 61 320
rect 53 319 54 320
rect 52 319 53 320
rect 51 319 52 320
rect 50 319 51 320
rect 49 319 50 320
rect 27 319 28 320
rect 26 319 27 320
rect 25 319 26 320
rect 24 319 25 320
rect 23 319 24 320
rect 22 319 23 320
rect 21 319 22 320
rect 20 319 21 320
rect 19 319 20 320
rect 18 319 19 320
rect 17 319 18 320
rect 14 319 15 320
rect 13 319 14 320
rect 194 320 195 321
rect 181 320 182 321
rect 180 320 181 321
rect 179 320 180 321
rect 177 320 178 321
rect 176 320 177 321
rect 175 320 176 321
rect 173 320 174 321
rect 172 320 173 321
rect 171 320 172 321
rect 169 320 170 321
rect 168 320 169 321
rect 167 320 168 321
rect 165 320 166 321
rect 164 320 165 321
rect 162 320 163 321
rect 161 320 162 321
rect 160 320 161 321
rect 110 320 111 321
rect 109 320 110 321
rect 108 320 109 321
rect 107 320 108 321
rect 106 320 107 321
rect 105 320 106 321
rect 104 320 105 321
rect 103 320 104 321
rect 102 320 103 321
rect 101 320 102 321
rect 100 320 101 321
rect 64 320 65 321
rect 63 320 64 321
rect 62 320 63 321
rect 61 320 62 321
rect 60 320 61 321
rect 53 320 54 321
rect 52 320 53 321
rect 51 320 52 321
rect 50 320 51 321
rect 49 320 50 321
rect 23 320 24 321
rect 22 320 23 321
rect 21 320 22 321
rect 20 320 21 321
rect 19 320 20 321
rect 18 320 19 321
rect 17 320 18 321
rect 16 320 17 321
rect 14 320 15 321
rect 13 320 14 321
rect 12 320 13 321
rect 195 321 196 322
rect 194 321 195 322
rect 193 321 194 322
rect 192 321 193 322
rect 191 321 192 322
rect 190 321 191 322
rect 189 321 190 322
rect 181 321 182 322
rect 180 321 181 322
rect 176 321 177 322
rect 175 321 176 322
rect 173 321 174 322
rect 172 321 173 322
rect 171 321 172 322
rect 169 321 170 322
rect 168 321 169 322
rect 167 321 168 322
rect 165 321 166 322
rect 164 321 165 322
rect 162 321 163 322
rect 161 321 162 322
rect 160 321 161 322
rect 110 321 111 322
rect 109 321 110 322
rect 108 321 109 322
rect 107 321 108 322
rect 106 321 107 322
rect 105 321 106 322
rect 104 321 105 322
rect 103 321 104 322
rect 102 321 103 322
rect 101 321 102 322
rect 100 321 101 322
rect 64 321 65 322
rect 63 321 64 322
rect 62 321 63 322
rect 61 321 62 322
rect 60 321 61 322
rect 53 321 54 322
rect 52 321 53 322
rect 51 321 52 322
rect 50 321 51 322
rect 49 321 50 322
rect 19 321 20 322
rect 18 321 19 322
rect 17 321 18 322
rect 14 321 15 322
rect 13 321 14 322
rect 12 321 13 322
rect 194 322 195 323
rect 193 322 194 323
rect 192 322 193 323
rect 191 322 192 323
rect 190 322 191 323
rect 189 322 190 323
rect 182 322 183 323
rect 181 322 182 323
rect 180 322 181 323
rect 176 322 177 323
rect 175 322 176 323
rect 174 322 175 323
rect 173 322 174 323
rect 172 322 173 323
rect 171 322 172 323
rect 169 322 170 323
rect 168 322 169 323
rect 167 322 168 323
rect 165 322 166 323
rect 164 322 165 323
rect 162 322 163 323
rect 161 322 162 323
rect 160 322 161 323
rect 110 322 111 323
rect 109 322 110 323
rect 108 322 109 323
rect 107 322 108 323
rect 106 322 107 323
rect 105 322 106 323
rect 104 322 105 323
rect 103 322 104 323
rect 102 322 103 323
rect 101 322 102 323
rect 100 322 101 323
rect 64 322 65 323
rect 63 322 64 323
rect 62 322 63 323
rect 61 322 62 323
rect 60 322 61 323
rect 53 322 54 323
rect 52 322 53 323
rect 51 322 52 323
rect 50 322 51 323
rect 49 322 50 323
rect 31 322 32 323
rect 30 322 31 323
rect 29 322 30 323
rect 28 322 29 323
rect 27 322 28 323
rect 26 322 27 323
rect 14 322 15 323
rect 13 322 14 323
rect 182 323 183 324
rect 181 323 182 324
rect 180 323 181 324
rect 176 323 177 324
rect 175 323 176 324
rect 174 323 175 324
rect 173 323 174 324
rect 172 323 173 324
rect 171 323 172 324
rect 170 323 171 324
rect 169 323 170 324
rect 168 323 169 324
rect 167 323 168 324
rect 165 323 166 324
rect 164 323 165 324
rect 162 323 163 324
rect 161 323 162 324
rect 160 323 161 324
rect 110 323 111 324
rect 109 323 110 324
rect 108 323 109 324
rect 107 323 108 324
rect 106 323 107 324
rect 105 323 106 324
rect 104 323 105 324
rect 103 323 104 324
rect 102 323 103 324
rect 101 323 102 324
rect 100 323 101 324
rect 64 323 65 324
rect 63 323 64 324
rect 62 323 63 324
rect 61 323 62 324
rect 60 323 61 324
rect 53 323 54 324
rect 52 323 53 324
rect 51 323 52 324
rect 50 323 51 324
rect 49 323 50 324
rect 31 323 32 324
rect 30 323 31 324
rect 29 323 30 324
rect 28 323 29 324
rect 27 323 28 324
rect 26 323 27 324
rect 25 323 26 324
rect 24 323 25 324
rect 23 323 24 324
rect 22 323 23 324
rect 194 324 195 325
rect 193 324 194 325
rect 192 324 193 325
rect 191 324 192 325
rect 190 324 191 325
rect 189 324 190 325
rect 182 324 183 325
rect 181 324 182 325
rect 180 324 181 325
rect 176 324 177 325
rect 175 324 176 325
rect 174 324 175 325
rect 173 324 174 325
rect 172 324 173 325
rect 171 324 172 325
rect 170 324 171 325
rect 169 324 170 325
rect 168 324 169 325
rect 167 324 168 325
rect 165 324 166 325
rect 164 324 165 325
rect 162 324 163 325
rect 161 324 162 325
rect 160 324 161 325
rect 110 324 111 325
rect 109 324 110 325
rect 108 324 109 325
rect 107 324 108 325
rect 106 324 107 325
rect 105 324 106 325
rect 104 324 105 325
rect 103 324 104 325
rect 102 324 103 325
rect 101 324 102 325
rect 100 324 101 325
rect 64 324 65 325
rect 63 324 64 325
rect 62 324 63 325
rect 61 324 62 325
rect 60 324 61 325
rect 53 324 54 325
rect 52 324 53 325
rect 51 324 52 325
rect 50 324 51 325
rect 49 324 50 325
rect 31 324 32 325
rect 30 324 31 325
rect 29 324 30 325
rect 28 324 29 325
rect 27 324 28 325
rect 26 324 27 325
rect 25 324 26 325
rect 24 324 25 325
rect 23 324 24 325
rect 22 324 23 325
rect 21 324 22 325
rect 20 324 21 325
rect 19 324 20 325
rect 18 324 19 325
rect 17 324 18 325
rect 195 325 196 326
rect 194 325 195 326
rect 193 325 194 326
rect 192 325 193 326
rect 191 325 192 326
rect 190 325 191 326
rect 189 325 190 326
rect 182 325 183 326
rect 181 325 182 326
rect 180 325 181 326
rect 176 325 177 326
rect 175 325 176 326
rect 174 325 175 326
rect 173 325 174 326
rect 172 325 173 326
rect 171 325 172 326
rect 170 325 171 326
rect 169 325 170 326
rect 168 325 169 326
rect 167 325 168 326
rect 165 325 166 326
rect 164 325 165 326
rect 162 325 163 326
rect 161 325 162 326
rect 160 325 161 326
rect 110 325 111 326
rect 109 325 110 326
rect 108 325 109 326
rect 107 325 108 326
rect 106 325 107 326
rect 105 325 106 326
rect 104 325 105 326
rect 103 325 104 326
rect 102 325 103 326
rect 101 325 102 326
rect 100 325 101 326
rect 64 325 65 326
rect 63 325 64 326
rect 62 325 63 326
rect 61 325 62 326
rect 60 325 61 326
rect 53 325 54 326
rect 52 325 53 326
rect 51 325 52 326
rect 50 325 51 326
rect 49 325 50 326
rect 27 325 28 326
rect 26 325 27 326
rect 25 325 26 326
rect 24 325 25 326
rect 23 325 24 326
rect 22 325 23 326
rect 21 325 22 326
rect 20 325 21 326
rect 19 325 20 326
rect 18 325 19 326
rect 17 325 18 326
rect 16 325 17 326
rect 194 326 195 327
rect 191 326 192 327
rect 190 326 191 327
rect 189 326 190 327
rect 182 326 183 327
rect 181 326 182 327
rect 180 326 181 327
rect 176 326 177 327
rect 175 326 176 327
rect 174 326 175 327
rect 173 326 174 327
rect 172 326 173 327
rect 171 326 172 327
rect 170 326 171 327
rect 169 326 170 327
rect 168 326 169 327
rect 167 326 168 327
rect 165 326 166 327
rect 164 326 165 327
rect 162 326 163 327
rect 161 326 162 327
rect 160 326 161 327
rect 110 326 111 327
rect 109 326 110 327
rect 108 326 109 327
rect 107 326 108 327
rect 106 326 107 327
rect 105 326 106 327
rect 104 326 105 327
rect 103 326 104 327
rect 102 326 103 327
rect 101 326 102 327
rect 100 326 101 327
rect 64 326 65 327
rect 63 326 64 327
rect 62 326 63 327
rect 61 326 62 327
rect 60 326 61 327
rect 53 326 54 327
rect 52 326 53 327
rect 51 326 52 327
rect 50 326 51 327
rect 49 326 50 327
rect 26 326 27 327
rect 25 326 26 327
rect 24 326 25 327
rect 23 326 24 327
rect 22 326 23 327
rect 21 326 22 327
rect 20 326 21 327
rect 19 326 20 327
rect 18 326 19 327
rect 17 326 18 327
rect 16 326 17 327
rect 190 327 191 328
rect 189 327 190 328
rect 182 327 183 328
rect 181 327 182 328
rect 180 327 181 328
rect 176 327 177 328
rect 175 327 176 328
rect 174 327 175 328
rect 173 327 174 328
rect 172 327 173 328
rect 171 327 172 328
rect 169 327 170 328
rect 168 327 169 328
rect 167 327 168 328
rect 165 327 166 328
rect 164 327 165 328
rect 162 327 163 328
rect 161 327 162 328
rect 160 327 161 328
rect 110 327 111 328
rect 109 327 110 328
rect 108 327 109 328
rect 107 327 108 328
rect 106 327 107 328
rect 105 327 106 328
rect 104 327 105 328
rect 103 327 104 328
rect 102 327 103 328
rect 101 327 102 328
rect 100 327 101 328
rect 53 327 54 328
rect 52 327 53 328
rect 51 327 52 328
rect 50 327 51 328
rect 49 327 50 328
rect 27 327 28 328
rect 26 327 27 328
rect 25 327 26 328
rect 19 327 20 328
rect 18 327 19 328
rect 17 327 18 328
rect 194 328 195 329
rect 193 328 194 329
rect 192 328 193 329
rect 191 328 192 329
rect 190 328 191 329
rect 189 328 190 329
rect 182 328 183 329
rect 181 328 182 329
rect 180 328 181 329
rect 177 328 178 329
rect 176 328 177 329
rect 175 328 176 329
rect 173 328 174 329
rect 172 328 173 329
rect 171 328 172 329
rect 169 328 170 329
rect 168 328 169 329
rect 167 328 168 329
rect 165 328 166 329
rect 164 328 165 329
rect 162 328 163 329
rect 161 328 162 329
rect 160 328 161 329
rect 110 328 111 329
rect 109 328 110 329
rect 108 328 109 329
rect 107 328 108 329
rect 106 328 107 329
rect 105 328 106 329
rect 104 328 105 329
rect 103 328 104 329
rect 102 328 103 329
rect 101 328 102 329
rect 100 328 101 329
rect 53 328 54 329
rect 52 328 53 329
rect 51 328 52 329
rect 50 328 51 329
rect 49 328 50 329
rect 27 328 28 329
rect 26 328 27 329
rect 18 328 19 329
rect 17 328 18 329
rect 195 329 196 330
rect 194 329 195 330
rect 193 329 194 330
rect 192 329 193 330
rect 191 329 192 330
rect 190 329 191 330
rect 189 329 190 330
rect 181 329 182 330
rect 180 329 181 330
rect 179 329 180 330
rect 177 329 178 330
rect 176 329 177 330
rect 175 329 176 330
rect 173 329 174 330
rect 172 329 173 330
rect 171 329 172 330
rect 169 329 170 330
rect 168 329 169 330
rect 167 329 168 330
rect 165 329 166 330
rect 164 329 165 330
rect 162 329 163 330
rect 161 329 162 330
rect 160 329 161 330
rect 110 329 111 330
rect 109 329 110 330
rect 108 329 109 330
rect 107 329 108 330
rect 106 329 107 330
rect 105 329 106 330
rect 104 329 105 330
rect 103 329 104 330
rect 102 329 103 330
rect 101 329 102 330
rect 100 329 101 330
rect 27 329 28 330
rect 26 329 27 330
rect 25 329 26 330
rect 17 329 18 330
rect 16 329 17 330
rect 181 330 182 331
rect 180 330 181 331
rect 179 330 180 331
rect 177 330 178 331
rect 176 330 177 331
rect 175 330 176 331
rect 173 330 174 331
rect 172 330 173 331
rect 171 330 172 331
rect 169 330 170 331
rect 168 330 169 331
rect 167 330 168 331
rect 165 330 166 331
rect 164 330 165 331
rect 162 330 163 331
rect 161 330 162 331
rect 160 330 161 331
rect 110 330 111 331
rect 109 330 110 331
rect 108 330 109 331
rect 107 330 108 331
rect 106 330 107 331
rect 105 330 106 331
rect 104 330 105 331
rect 103 330 104 331
rect 102 330 103 331
rect 101 330 102 331
rect 100 330 101 331
rect 27 330 28 331
rect 26 330 27 331
rect 25 330 26 331
rect 24 330 25 331
rect 18 330 19 331
rect 17 330 18 331
rect 16 330 17 331
rect 194 331 195 332
rect 193 331 194 332
rect 192 331 193 332
rect 191 331 192 332
rect 190 331 191 332
rect 189 331 190 332
rect 187 331 188 332
rect 186 331 187 332
rect 181 331 182 332
rect 180 331 181 332
rect 179 331 180 332
rect 178 331 179 332
rect 177 331 178 332
rect 176 331 177 332
rect 175 331 176 332
rect 173 331 174 332
rect 172 331 173 332
rect 171 331 172 332
rect 169 331 170 332
rect 168 331 169 332
rect 167 331 168 332
rect 165 331 166 332
rect 164 331 165 332
rect 162 331 163 332
rect 161 331 162 332
rect 160 331 161 332
rect 110 331 111 332
rect 109 331 110 332
rect 108 331 109 332
rect 107 331 108 332
rect 106 331 107 332
rect 105 331 106 332
rect 104 331 105 332
rect 103 331 104 332
rect 102 331 103 332
rect 101 331 102 332
rect 100 331 101 332
rect 26 331 27 332
rect 25 331 26 332
rect 24 331 25 332
rect 23 331 24 332
rect 22 331 23 332
rect 21 331 22 332
rect 20 331 21 332
rect 19 331 20 332
rect 18 331 19 332
rect 17 331 18 332
rect 16 331 17 332
rect 195 332 196 333
rect 194 332 195 333
rect 193 332 194 333
rect 192 332 193 333
rect 191 332 192 333
rect 190 332 191 333
rect 189 332 190 333
rect 187 332 188 333
rect 186 332 187 333
rect 181 332 182 333
rect 180 332 181 333
rect 179 332 180 333
rect 178 332 179 333
rect 177 332 178 333
rect 176 332 177 333
rect 173 332 174 333
rect 172 332 173 333
rect 171 332 172 333
rect 169 332 170 333
rect 168 332 169 333
rect 167 332 168 333
rect 165 332 166 333
rect 164 332 165 333
rect 162 332 163 333
rect 161 332 162 333
rect 160 332 161 333
rect 110 332 111 333
rect 109 332 110 333
rect 108 332 109 333
rect 107 332 108 333
rect 106 332 107 333
rect 105 332 106 333
rect 104 332 105 333
rect 103 332 104 333
rect 102 332 103 333
rect 101 332 102 333
rect 100 332 101 333
rect 25 332 26 333
rect 24 332 25 333
rect 23 332 24 333
rect 22 332 23 333
rect 21 332 22 333
rect 20 332 21 333
rect 19 332 20 333
rect 18 332 19 333
rect 17 332 18 333
rect 194 333 195 334
rect 192 333 193 334
rect 187 333 188 334
rect 180 333 181 334
rect 179 333 180 334
rect 178 333 179 334
rect 177 333 178 334
rect 176 333 177 334
rect 173 333 174 334
rect 172 333 173 334
rect 171 333 172 334
rect 169 333 170 334
rect 168 333 169 334
rect 167 333 168 334
rect 165 333 166 334
rect 164 333 165 334
rect 162 333 163 334
rect 161 333 162 334
rect 160 333 161 334
rect 110 333 111 334
rect 109 333 110 334
rect 108 333 109 334
rect 107 333 108 334
rect 106 333 107 334
rect 105 333 106 334
rect 104 333 105 334
rect 103 333 104 334
rect 102 333 103 334
rect 101 333 102 334
rect 100 333 101 334
rect 76 333 77 334
rect 75 333 76 334
rect 74 333 75 334
rect 73 333 74 334
rect 72 333 73 334
rect 71 333 72 334
rect 70 333 71 334
rect 69 333 70 334
rect 68 333 69 334
rect 67 333 68 334
rect 66 333 67 334
rect 65 333 66 334
rect 64 333 65 334
rect 63 333 64 334
rect 62 333 63 334
rect 61 333 62 334
rect 60 333 61 334
rect 59 333 60 334
rect 58 333 59 334
rect 57 333 58 334
rect 56 333 57 334
rect 55 333 56 334
rect 54 333 55 334
rect 53 333 54 334
rect 52 333 53 334
rect 51 333 52 334
rect 50 333 51 334
rect 49 333 50 334
rect 24 333 25 334
rect 23 333 24 334
rect 22 333 23 334
rect 21 333 22 334
rect 20 333 21 334
rect 19 333 20 334
rect 18 333 19 334
rect 17 333 18 334
rect 193 334 194 335
rect 192 334 193 335
rect 191 334 192 335
rect 190 334 191 335
rect 179 334 180 335
rect 178 334 179 335
rect 177 334 178 335
rect 173 334 174 335
rect 172 334 173 335
rect 171 334 172 335
rect 168 334 169 335
rect 167 334 168 335
rect 110 334 111 335
rect 109 334 110 335
rect 108 334 109 335
rect 107 334 108 335
rect 106 334 107 335
rect 105 334 106 335
rect 104 334 105 335
rect 103 334 104 335
rect 102 334 103 335
rect 101 334 102 335
rect 100 334 101 335
rect 76 334 77 335
rect 75 334 76 335
rect 74 334 75 335
rect 73 334 74 335
rect 72 334 73 335
rect 71 334 72 335
rect 70 334 71 335
rect 69 334 70 335
rect 68 334 69 335
rect 67 334 68 335
rect 66 334 67 335
rect 65 334 66 335
rect 64 334 65 335
rect 63 334 64 335
rect 62 334 63 335
rect 61 334 62 335
rect 60 334 61 335
rect 59 334 60 335
rect 58 334 59 335
rect 57 334 58 335
rect 56 334 57 335
rect 55 334 56 335
rect 54 334 55 335
rect 53 334 54 335
rect 52 334 53 335
rect 51 334 52 335
rect 50 334 51 335
rect 49 334 50 335
rect 22 334 23 335
rect 21 334 22 335
rect 20 334 21 335
rect 19 334 20 335
rect 194 335 195 336
rect 193 335 194 336
rect 192 335 193 336
rect 191 335 192 336
rect 190 335 191 336
rect 189 335 190 336
rect 173 335 174 336
rect 172 335 173 336
rect 171 335 172 336
rect 110 335 111 336
rect 109 335 110 336
rect 108 335 109 336
rect 107 335 108 336
rect 106 335 107 336
rect 105 335 106 336
rect 104 335 105 336
rect 103 335 104 336
rect 102 335 103 336
rect 101 335 102 336
rect 100 335 101 336
rect 76 335 77 336
rect 75 335 76 336
rect 74 335 75 336
rect 73 335 74 336
rect 72 335 73 336
rect 71 335 72 336
rect 70 335 71 336
rect 69 335 70 336
rect 68 335 69 336
rect 67 335 68 336
rect 66 335 67 336
rect 65 335 66 336
rect 64 335 65 336
rect 63 335 64 336
rect 62 335 63 336
rect 61 335 62 336
rect 60 335 61 336
rect 59 335 60 336
rect 58 335 59 336
rect 57 335 58 336
rect 56 335 57 336
rect 55 335 56 336
rect 54 335 55 336
rect 53 335 54 336
rect 52 335 53 336
rect 51 335 52 336
rect 50 335 51 336
rect 49 335 50 336
rect 194 336 195 337
rect 193 336 194 337
rect 190 336 191 337
rect 189 336 190 337
rect 173 336 174 337
rect 172 336 173 337
rect 171 336 172 337
rect 110 336 111 337
rect 109 336 110 337
rect 108 336 109 337
rect 107 336 108 337
rect 106 336 107 337
rect 105 336 106 337
rect 104 336 105 337
rect 103 336 104 337
rect 102 336 103 337
rect 101 336 102 337
rect 100 336 101 337
rect 76 336 77 337
rect 75 336 76 337
rect 74 336 75 337
rect 73 336 74 337
rect 72 336 73 337
rect 71 336 72 337
rect 70 336 71 337
rect 69 336 70 337
rect 68 336 69 337
rect 67 336 68 337
rect 66 336 67 337
rect 65 336 66 337
rect 64 336 65 337
rect 63 336 64 337
rect 62 336 63 337
rect 61 336 62 337
rect 60 336 61 337
rect 59 336 60 337
rect 58 336 59 337
rect 57 336 58 337
rect 56 336 57 337
rect 55 336 56 337
rect 54 336 55 337
rect 53 336 54 337
rect 52 336 53 337
rect 51 336 52 337
rect 50 336 51 337
rect 49 336 50 337
rect 195 337 196 338
rect 194 337 195 338
rect 190 337 191 338
rect 189 337 190 338
rect 172 337 173 338
rect 110 337 111 338
rect 109 337 110 338
rect 108 337 109 338
rect 107 337 108 338
rect 106 337 107 338
rect 105 337 106 338
rect 104 337 105 338
rect 103 337 104 338
rect 102 337 103 338
rect 101 337 102 338
rect 100 337 101 338
rect 76 337 77 338
rect 75 337 76 338
rect 74 337 75 338
rect 73 337 74 338
rect 72 337 73 338
rect 71 337 72 338
rect 70 337 71 338
rect 69 337 70 338
rect 68 337 69 338
rect 67 337 68 338
rect 66 337 67 338
rect 65 337 66 338
rect 64 337 65 338
rect 63 337 64 338
rect 62 337 63 338
rect 61 337 62 338
rect 60 337 61 338
rect 59 337 60 338
rect 58 337 59 338
rect 57 337 58 338
rect 56 337 57 338
rect 55 337 56 338
rect 54 337 55 338
rect 53 337 54 338
rect 52 337 53 338
rect 51 337 52 338
rect 50 337 51 338
rect 49 337 50 338
rect 194 338 195 339
rect 190 338 191 339
rect 189 338 190 339
rect 110 338 111 339
rect 109 338 110 339
rect 108 338 109 339
rect 107 338 108 339
rect 106 338 107 339
rect 105 338 106 339
rect 104 338 105 339
rect 103 338 104 339
rect 102 338 103 339
rect 101 338 102 339
rect 100 338 101 339
rect 76 338 77 339
rect 75 338 76 339
rect 74 338 75 339
rect 73 338 74 339
rect 72 338 73 339
rect 71 338 72 339
rect 70 338 71 339
rect 69 338 70 339
rect 68 338 69 339
rect 67 338 68 339
rect 66 338 67 339
rect 65 338 66 339
rect 64 338 65 339
rect 63 338 64 339
rect 62 338 63 339
rect 61 338 62 339
rect 60 338 61 339
rect 59 338 60 339
rect 58 338 59 339
rect 57 338 58 339
rect 56 338 57 339
rect 55 338 56 339
rect 54 338 55 339
rect 53 338 54 339
rect 52 338 53 339
rect 51 338 52 339
rect 50 338 51 339
rect 49 338 50 339
rect 193 339 194 340
rect 110 339 111 340
rect 109 339 110 340
rect 108 339 109 340
rect 107 339 108 340
rect 106 339 107 340
rect 105 339 106 340
rect 104 339 105 340
rect 103 339 104 340
rect 102 339 103 340
rect 101 339 102 340
rect 100 339 101 340
rect 194 340 195 341
rect 193 340 194 341
rect 192 340 193 341
rect 190 340 191 341
rect 189 340 190 341
rect 110 340 111 341
rect 109 340 110 341
rect 108 340 109 341
rect 107 340 108 341
rect 106 340 107 341
rect 105 340 106 341
rect 104 340 105 341
rect 103 340 104 341
rect 102 340 103 341
rect 101 340 102 341
rect 100 340 101 341
rect 195 341 196 342
rect 194 341 195 342
rect 193 341 194 342
rect 192 341 193 342
rect 191 341 192 342
rect 190 341 191 342
rect 189 341 190 342
rect 27 341 28 342
rect 26 341 27 342
rect 195 342 196 343
rect 194 342 195 343
rect 192 342 193 343
rect 191 342 192 343
rect 190 342 191 343
rect 189 342 190 343
rect 27 342 28 343
rect 26 342 27 343
rect 25 342 26 343
rect 24 342 25 343
rect 23 342 24 343
rect 22 342 23 343
rect 194 343 195 344
rect 193 343 194 344
rect 192 343 193 344
rect 191 343 192 344
rect 190 343 191 344
rect 189 343 190 344
rect 27 343 28 344
rect 26 343 27 344
rect 25 343 26 344
rect 24 343 25 344
rect 23 343 24 344
rect 22 343 23 344
rect 21 343 22 344
rect 20 343 21 344
rect 19 343 20 344
rect 18 343 19 344
rect 17 343 18 344
rect 195 344 196 345
rect 194 344 195 345
rect 193 344 194 345
rect 192 344 193 345
rect 191 344 192 345
rect 190 344 191 345
rect 189 344 190 345
rect 76 344 77 345
rect 75 344 76 345
rect 74 344 75 345
rect 73 344 74 345
rect 72 344 73 345
rect 71 344 72 345
rect 70 344 71 345
rect 69 344 70 345
rect 68 344 69 345
rect 67 344 68 345
rect 66 344 67 345
rect 65 344 66 345
rect 64 344 65 345
rect 63 344 64 345
rect 62 344 63 345
rect 61 344 62 345
rect 60 344 61 345
rect 59 344 60 345
rect 58 344 59 345
rect 57 344 58 345
rect 56 344 57 345
rect 55 344 56 345
rect 54 344 55 345
rect 53 344 54 345
rect 52 344 53 345
rect 51 344 52 345
rect 50 344 51 345
rect 49 344 50 345
rect 26 344 27 345
rect 25 344 26 345
rect 24 344 25 345
rect 23 344 24 345
rect 22 344 23 345
rect 21 344 22 345
rect 20 344 21 345
rect 19 344 20 345
rect 18 344 19 345
rect 17 344 18 345
rect 16 344 17 345
rect 15 344 16 345
rect 14 344 15 345
rect 13 344 14 345
rect 194 345 195 346
rect 76 345 77 346
rect 75 345 76 346
rect 74 345 75 346
rect 73 345 74 346
rect 72 345 73 346
rect 71 345 72 346
rect 70 345 71 346
rect 69 345 70 346
rect 68 345 69 346
rect 67 345 68 346
rect 66 345 67 346
rect 65 345 66 346
rect 64 345 65 346
rect 63 345 64 346
rect 62 345 63 346
rect 61 345 62 346
rect 60 345 61 346
rect 59 345 60 346
rect 58 345 59 346
rect 57 345 58 346
rect 56 345 57 346
rect 55 345 56 346
rect 54 345 55 346
rect 53 345 54 346
rect 52 345 53 346
rect 51 345 52 346
rect 50 345 51 346
rect 49 345 50 346
rect 21 345 22 346
rect 20 345 21 346
rect 19 345 20 346
rect 18 345 19 346
rect 17 345 18 346
rect 16 345 17 346
rect 15 345 16 346
rect 14 345 15 346
rect 13 345 14 346
rect 12 345 13 346
rect 190 346 191 347
rect 189 346 190 347
rect 76 346 77 347
rect 75 346 76 347
rect 74 346 75 347
rect 73 346 74 347
rect 72 346 73 347
rect 71 346 72 347
rect 70 346 71 347
rect 69 346 70 347
rect 68 346 69 347
rect 67 346 68 347
rect 66 346 67 347
rect 65 346 66 347
rect 64 346 65 347
rect 63 346 64 347
rect 62 346 63 347
rect 61 346 62 347
rect 60 346 61 347
rect 59 346 60 347
rect 58 346 59 347
rect 57 346 58 347
rect 56 346 57 347
rect 55 346 56 347
rect 54 346 55 347
rect 53 346 54 347
rect 52 346 53 347
rect 51 346 52 347
rect 50 346 51 347
rect 49 346 50 347
rect 18 346 19 347
rect 17 346 18 347
rect 16 346 17 347
rect 15 346 16 347
rect 14 346 15 347
rect 13 346 14 347
rect 12 346 13 347
rect 194 347 195 348
rect 193 347 194 348
rect 192 347 193 348
rect 191 347 192 348
rect 190 347 191 348
rect 189 347 190 348
rect 188 347 189 348
rect 187 347 188 348
rect 171 347 172 348
rect 76 347 77 348
rect 75 347 76 348
rect 74 347 75 348
rect 73 347 74 348
rect 72 347 73 348
rect 71 347 72 348
rect 70 347 71 348
rect 69 347 70 348
rect 68 347 69 348
rect 67 347 68 348
rect 66 347 67 348
rect 65 347 66 348
rect 64 347 65 348
rect 63 347 64 348
rect 62 347 63 348
rect 61 347 62 348
rect 60 347 61 348
rect 59 347 60 348
rect 58 347 59 348
rect 57 347 58 348
rect 56 347 57 348
rect 55 347 56 348
rect 54 347 55 348
rect 53 347 54 348
rect 52 347 53 348
rect 51 347 52 348
rect 50 347 51 348
rect 49 347 50 348
rect 27 347 28 348
rect 26 347 27 348
rect 25 347 26 348
rect 24 347 25 348
rect 23 347 24 348
rect 22 347 23 348
rect 21 347 22 348
rect 20 347 21 348
rect 19 347 20 348
rect 18 347 19 348
rect 17 347 18 348
rect 16 347 17 348
rect 15 347 16 348
rect 14 347 15 348
rect 13 347 14 348
rect 12 347 13 348
rect 194 348 195 349
rect 193 348 194 349
rect 192 348 193 349
rect 191 348 192 349
rect 190 348 191 349
rect 189 348 190 349
rect 188 348 189 349
rect 187 348 188 349
rect 172 348 173 349
rect 171 348 172 349
rect 170 348 171 349
rect 76 348 77 349
rect 75 348 76 349
rect 74 348 75 349
rect 73 348 74 349
rect 72 348 73 349
rect 71 348 72 349
rect 70 348 71 349
rect 69 348 70 349
rect 68 348 69 349
rect 67 348 68 349
rect 66 348 67 349
rect 65 348 66 349
rect 64 348 65 349
rect 63 348 64 349
rect 62 348 63 349
rect 61 348 62 349
rect 60 348 61 349
rect 59 348 60 349
rect 58 348 59 349
rect 57 348 58 349
rect 56 348 57 349
rect 55 348 56 349
rect 54 348 55 349
rect 53 348 54 349
rect 52 348 53 349
rect 51 348 52 349
rect 50 348 51 349
rect 49 348 50 349
rect 27 348 28 349
rect 26 348 27 349
rect 25 348 26 349
rect 24 348 25 349
rect 23 348 24 349
rect 22 348 23 349
rect 21 348 22 349
rect 20 348 21 349
rect 19 348 20 349
rect 18 348 19 349
rect 17 348 18 349
rect 16 348 17 349
rect 15 348 16 349
rect 14 348 15 349
rect 13 348 14 349
rect 195 349 196 350
rect 194 349 195 350
rect 190 349 191 350
rect 189 349 190 350
rect 172 349 173 350
rect 171 349 172 350
rect 170 349 171 350
rect 76 349 77 350
rect 75 349 76 350
rect 74 349 75 350
rect 73 349 74 350
rect 72 349 73 350
rect 71 349 72 350
rect 70 349 71 350
rect 69 349 70 350
rect 68 349 69 350
rect 67 349 68 350
rect 66 349 67 350
rect 65 349 66 350
rect 64 349 65 350
rect 63 349 64 350
rect 62 349 63 350
rect 61 349 62 350
rect 60 349 61 350
rect 59 349 60 350
rect 58 349 59 350
rect 57 349 58 350
rect 56 349 57 350
rect 55 349 56 350
rect 54 349 55 350
rect 53 349 54 350
rect 52 349 53 350
rect 51 349 52 350
rect 50 349 51 350
rect 49 349 50 350
rect 27 349 28 350
rect 26 349 27 350
rect 25 349 26 350
rect 24 349 25 350
rect 23 349 24 350
rect 22 349 23 350
rect 194 350 195 351
rect 189 350 190 351
rect 172 350 173 351
rect 171 350 172 351
rect 170 350 171 351
rect 169 350 170 351
rect 65 350 66 351
rect 64 350 65 351
rect 63 350 64 351
rect 62 350 63 351
rect 61 350 62 351
rect 60 350 61 351
rect 53 350 54 351
rect 52 350 53 351
rect 51 350 52 351
rect 50 350 51 351
rect 49 350 50 351
rect 26 350 27 351
rect 25 350 26 351
rect 24 350 25 351
rect 23 350 24 351
rect 22 350 23 351
rect 21 350 22 351
rect 20 350 21 351
rect 194 351 195 352
rect 193 351 194 352
rect 192 351 193 352
rect 191 351 192 352
rect 190 351 191 352
rect 189 351 190 352
rect 187 351 188 352
rect 186 351 187 352
rect 171 351 172 352
rect 170 351 171 352
rect 169 351 170 352
rect 168 351 169 352
rect 64 351 65 352
rect 63 351 64 352
rect 62 351 63 352
rect 61 351 62 352
rect 60 351 61 352
rect 53 351 54 352
rect 52 351 53 352
rect 51 351 52 352
rect 50 351 51 352
rect 49 351 50 352
rect 24 351 25 352
rect 23 351 24 352
rect 22 351 23 352
rect 21 351 22 352
rect 20 351 21 352
rect 19 351 20 352
rect 18 351 19 352
rect 194 352 195 353
rect 193 352 194 353
rect 192 352 193 353
rect 191 352 192 353
rect 190 352 191 353
rect 189 352 190 353
rect 187 352 188 353
rect 186 352 187 353
rect 180 352 181 353
rect 179 352 180 353
rect 178 352 179 353
rect 177 352 178 353
rect 176 352 177 353
rect 175 352 176 353
rect 174 352 175 353
rect 171 352 172 353
rect 170 352 171 353
rect 169 352 170 353
rect 168 352 169 353
rect 167 352 168 353
rect 147 352 148 353
rect 146 352 147 353
rect 145 352 146 353
rect 144 352 145 353
rect 143 352 144 353
rect 142 352 143 353
rect 141 352 142 353
rect 140 352 141 353
rect 139 352 140 353
rect 138 352 139 353
rect 137 352 138 353
rect 136 352 137 353
rect 135 352 136 353
rect 134 352 135 353
rect 133 352 134 353
rect 132 352 133 353
rect 131 352 132 353
rect 130 352 131 353
rect 129 352 130 353
rect 128 352 129 353
rect 127 352 128 353
rect 126 352 127 353
rect 125 352 126 353
rect 124 352 125 353
rect 123 352 124 353
rect 122 352 123 353
rect 121 352 122 353
rect 120 352 121 353
rect 119 352 120 353
rect 118 352 119 353
rect 117 352 118 353
rect 116 352 117 353
rect 115 352 116 353
rect 114 352 115 353
rect 113 352 114 353
rect 112 352 113 353
rect 111 352 112 353
rect 110 352 111 353
rect 109 352 110 353
rect 108 352 109 353
rect 107 352 108 353
rect 106 352 107 353
rect 105 352 106 353
rect 104 352 105 353
rect 103 352 104 353
rect 102 352 103 353
rect 101 352 102 353
rect 100 352 101 353
rect 65 352 66 353
rect 64 352 65 353
rect 63 352 64 353
rect 62 352 63 353
rect 61 352 62 353
rect 60 352 61 353
rect 53 352 54 353
rect 52 352 53 353
rect 51 352 52 353
rect 50 352 51 353
rect 49 352 50 353
rect 22 352 23 353
rect 21 352 22 353
rect 20 352 21 353
rect 19 352 20 353
rect 18 352 19 353
rect 17 352 18 353
rect 16 352 17 353
rect 181 353 182 354
rect 180 353 181 354
rect 179 353 180 354
rect 178 353 179 354
rect 177 353 178 354
rect 176 353 177 354
rect 175 353 176 354
rect 174 353 175 354
rect 170 353 171 354
rect 169 353 170 354
rect 168 353 169 354
rect 167 353 168 354
rect 166 353 167 354
rect 165 353 166 354
rect 164 353 165 354
rect 147 353 148 354
rect 146 353 147 354
rect 145 353 146 354
rect 144 353 145 354
rect 143 353 144 354
rect 142 353 143 354
rect 141 353 142 354
rect 140 353 141 354
rect 139 353 140 354
rect 138 353 139 354
rect 137 353 138 354
rect 136 353 137 354
rect 135 353 136 354
rect 134 353 135 354
rect 133 353 134 354
rect 132 353 133 354
rect 131 353 132 354
rect 130 353 131 354
rect 129 353 130 354
rect 128 353 129 354
rect 127 353 128 354
rect 126 353 127 354
rect 125 353 126 354
rect 124 353 125 354
rect 123 353 124 354
rect 122 353 123 354
rect 121 353 122 354
rect 120 353 121 354
rect 119 353 120 354
rect 118 353 119 354
rect 117 353 118 354
rect 116 353 117 354
rect 115 353 116 354
rect 114 353 115 354
rect 113 353 114 354
rect 112 353 113 354
rect 111 353 112 354
rect 110 353 111 354
rect 109 353 110 354
rect 108 353 109 354
rect 107 353 108 354
rect 106 353 107 354
rect 105 353 106 354
rect 104 353 105 354
rect 103 353 104 354
rect 102 353 103 354
rect 101 353 102 354
rect 100 353 101 354
rect 65 353 66 354
rect 64 353 65 354
rect 63 353 64 354
rect 62 353 63 354
rect 61 353 62 354
rect 60 353 61 354
rect 53 353 54 354
rect 52 353 53 354
rect 51 353 52 354
rect 50 353 51 354
rect 49 353 50 354
rect 27 353 28 354
rect 26 353 27 354
rect 25 353 26 354
rect 19 353 20 354
rect 18 353 19 354
rect 17 353 18 354
rect 16 353 17 354
rect 15 353 16 354
rect 14 353 15 354
rect 194 354 195 355
rect 193 354 194 355
rect 192 354 193 355
rect 191 354 192 355
rect 190 354 191 355
rect 181 354 182 355
rect 180 354 181 355
rect 179 354 180 355
rect 178 354 179 355
rect 177 354 178 355
rect 176 354 177 355
rect 175 354 176 355
rect 174 354 175 355
rect 169 354 170 355
rect 168 354 169 355
rect 167 354 168 355
rect 166 354 167 355
rect 165 354 166 355
rect 164 354 165 355
rect 163 354 164 355
rect 162 354 163 355
rect 161 354 162 355
rect 160 354 161 355
rect 147 354 148 355
rect 146 354 147 355
rect 145 354 146 355
rect 144 354 145 355
rect 143 354 144 355
rect 142 354 143 355
rect 141 354 142 355
rect 140 354 141 355
rect 139 354 140 355
rect 138 354 139 355
rect 137 354 138 355
rect 136 354 137 355
rect 135 354 136 355
rect 134 354 135 355
rect 133 354 134 355
rect 132 354 133 355
rect 131 354 132 355
rect 130 354 131 355
rect 129 354 130 355
rect 128 354 129 355
rect 127 354 128 355
rect 126 354 127 355
rect 125 354 126 355
rect 124 354 125 355
rect 123 354 124 355
rect 122 354 123 355
rect 121 354 122 355
rect 120 354 121 355
rect 119 354 120 355
rect 118 354 119 355
rect 117 354 118 355
rect 116 354 117 355
rect 115 354 116 355
rect 114 354 115 355
rect 113 354 114 355
rect 112 354 113 355
rect 111 354 112 355
rect 110 354 111 355
rect 109 354 110 355
rect 108 354 109 355
rect 107 354 108 355
rect 106 354 107 355
rect 105 354 106 355
rect 104 354 105 355
rect 103 354 104 355
rect 102 354 103 355
rect 101 354 102 355
rect 100 354 101 355
rect 65 354 66 355
rect 64 354 65 355
rect 63 354 64 355
rect 62 354 63 355
rect 61 354 62 355
rect 60 354 61 355
rect 53 354 54 355
rect 52 354 53 355
rect 51 354 52 355
rect 50 354 51 355
rect 49 354 50 355
rect 27 354 28 355
rect 26 354 27 355
rect 25 354 26 355
rect 24 354 25 355
rect 23 354 24 355
rect 22 354 23 355
rect 21 354 22 355
rect 20 354 21 355
rect 18 354 19 355
rect 17 354 18 355
rect 16 354 17 355
rect 15 354 16 355
rect 14 354 15 355
rect 13 354 14 355
rect 194 355 195 356
rect 193 355 194 356
rect 192 355 193 356
rect 191 355 192 356
rect 190 355 191 356
rect 189 355 190 356
rect 181 355 182 356
rect 180 355 181 356
rect 179 355 180 356
rect 178 355 179 356
rect 168 355 169 356
rect 167 355 168 356
rect 166 355 167 356
rect 165 355 166 356
rect 164 355 165 356
rect 163 355 164 356
rect 162 355 163 356
rect 161 355 162 356
rect 160 355 161 356
rect 147 355 148 356
rect 146 355 147 356
rect 145 355 146 356
rect 144 355 145 356
rect 143 355 144 356
rect 142 355 143 356
rect 141 355 142 356
rect 140 355 141 356
rect 139 355 140 356
rect 138 355 139 356
rect 137 355 138 356
rect 136 355 137 356
rect 135 355 136 356
rect 134 355 135 356
rect 133 355 134 356
rect 132 355 133 356
rect 131 355 132 356
rect 130 355 131 356
rect 129 355 130 356
rect 128 355 129 356
rect 127 355 128 356
rect 126 355 127 356
rect 125 355 126 356
rect 124 355 125 356
rect 123 355 124 356
rect 122 355 123 356
rect 121 355 122 356
rect 120 355 121 356
rect 119 355 120 356
rect 118 355 119 356
rect 117 355 118 356
rect 116 355 117 356
rect 115 355 116 356
rect 114 355 115 356
rect 113 355 114 356
rect 112 355 113 356
rect 111 355 112 356
rect 110 355 111 356
rect 109 355 110 356
rect 108 355 109 356
rect 107 355 108 356
rect 106 355 107 356
rect 105 355 106 356
rect 104 355 105 356
rect 103 355 104 356
rect 102 355 103 356
rect 101 355 102 356
rect 100 355 101 356
rect 66 355 67 356
rect 65 355 66 356
rect 64 355 65 356
rect 63 355 64 356
rect 62 355 63 356
rect 61 355 62 356
rect 60 355 61 356
rect 53 355 54 356
rect 52 355 53 356
rect 51 355 52 356
rect 50 355 51 356
rect 49 355 50 356
rect 27 355 28 356
rect 26 355 27 356
rect 25 355 26 356
rect 24 355 25 356
rect 23 355 24 356
rect 22 355 23 356
rect 21 355 22 356
rect 20 355 21 356
rect 19 355 20 356
rect 18 355 19 356
rect 17 355 18 356
rect 16 355 17 356
rect 15 355 16 356
rect 14 355 15 356
rect 13 355 14 356
rect 12 355 13 356
rect 194 356 195 357
rect 190 356 191 357
rect 189 356 190 357
rect 181 356 182 357
rect 180 356 181 357
rect 179 356 180 357
rect 178 356 179 357
rect 169 356 170 357
rect 168 356 169 357
rect 167 356 168 357
rect 166 356 167 357
rect 165 356 166 357
rect 164 356 165 357
rect 163 356 164 357
rect 162 356 163 357
rect 161 356 162 357
rect 160 356 161 357
rect 147 356 148 357
rect 146 356 147 357
rect 145 356 146 357
rect 144 356 145 357
rect 143 356 144 357
rect 142 356 143 357
rect 141 356 142 357
rect 140 356 141 357
rect 139 356 140 357
rect 138 356 139 357
rect 137 356 138 357
rect 136 356 137 357
rect 135 356 136 357
rect 134 356 135 357
rect 133 356 134 357
rect 132 356 133 357
rect 131 356 132 357
rect 130 356 131 357
rect 129 356 130 357
rect 128 356 129 357
rect 127 356 128 357
rect 126 356 127 357
rect 125 356 126 357
rect 124 356 125 357
rect 123 356 124 357
rect 122 356 123 357
rect 121 356 122 357
rect 120 356 121 357
rect 119 356 120 357
rect 118 356 119 357
rect 117 356 118 357
rect 116 356 117 357
rect 115 356 116 357
rect 114 356 115 357
rect 113 356 114 357
rect 112 356 113 357
rect 111 356 112 357
rect 110 356 111 357
rect 109 356 110 357
rect 108 356 109 357
rect 107 356 108 357
rect 106 356 107 357
rect 105 356 106 357
rect 104 356 105 357
rect 103 356 104 357
rect 102 356 103 357
rect 101 356 102 357
rect 100 356 101 357
rect 68 356 69 357
rect 67 356 68 357
rect 66 356 67 357
rect 65 356 66 357
rect 64 356 65 357
rect 63 356 64 357
rect 62 356 63 357
rect 61 356 62 357
rect 60 356 61 357
rect 53 356 54 357
rect 52 356 53 357
rect 51 356 52 357
rect 50 356 51 357
rect 49 356 50 357
rect 24 356 25 357
rect 23 356 24 357
rect 22 356 23 357
rect 21 356 22 357
rect 20 356 21 357
rect 19 356 20 357
rect 18 356 19 357
rect 17 356 18 357
rect 16 356 17 357
rect 15 356 16 357
rect 14 356 15 357
rect 13 356 14 357
rect 12 356 13 357
rect 195 357 196 358
rect 194 357 195 358
rect 190 357 191 358
rect 189 357 190 358
rect 181 357 182 358
rect 180 357 181 358
rect 179 357 180 358
rect 178 357 179 358
rect 169 357 170 358
rect 168 357 169 358
rect 167 357 168 358
rect 166 357 167 358
rect 165 357 166 358
rect 164 357 165 358
rect 163 357 164 358
rect 162 357 163 358
rect 161 357 162 358
rect 160 357 161 358
rect 147 357 148 358
rect 146 357 147 358
rect 145 357 146 358
rect 144 357 145 358
rect 143 357 144 358
rect 142 357 143 358
rect 141 357 142 358
rect 140 357 141 358
rect 139 357 140 358
rect 138 357 139 358
rect 137 357 138 358
rect 136 357 137 358
rect 135 357 136 358
rect 134 357 135 358
rect 133 357 134 358
rect 132 357 133 358
rect 131 357 132 358
rect 130 357 131 358
rect 129 357 130 358
rect 128 357 129 358
rect 127 357 128 358
rect 126 357 127 358
rect 125 357 126 358
rect 124 357 125 358
rect 123 357 124 358
rect 122 357 123 358
rect 121 357 122 358
rect 120 357 121 358
rect 119 357 120 358
rect 118 357 119 358
rect 117 357 118 358
rect 116 357 117 358
rect 115 357 116 358
rect 114 357 115 358
rect 113 357 114 358
rect 112 357 113 358
rect 111 357 112 358
rect 110 357 111 358
rect 109 357 110 358
rect 108 357 109 358
rect 107 357 108 358
rect 106 357 107 358
rect 105 357 106 358
rect 104 357 105 358
rect 103 357 104 358
rect 102 357 103 358
rect 101 357 102 358
rect 100 357 101 358
rect 69 357 70 358
rect 68 357 69 358
rect 67 357 68 358
rect 66 357 67 358
rect 65 357 66 358
rect 64 357 65 358
rect 63 357 64 358
rect 62 357 63 358
rect 61 357 62 358
rect 60 357 61 358
rect 53 357 54 358
rect 52 357 53 358
rect 51 357 52 358
rect 50 357 51 358
rect 49 357 50 358
rect 19 357 20 358
rect 18 357 19 358
rect 17 357 18 358
rect 16 357 17 358
rect 15 357 16 358
rect 14 357 15 358
rect 13 357 14 358
rect 12 357 13 358
rect 194 358 195 359
rect 193 358 194 359
rect 192 358 193 359
rect 191 358 192 359
rect 190 358 191 359
rect 189 358 190 359
rect 181 358 182 359
rect 180 358 181 359
rect 179 358 180 359
rect 178 358 179 359
rect 170 358 171 359
rect 169 358 170 359
rect 168 358 169 359
rect 167 358 168 359
rect 166 358 167 359
rect 147 358 148 359
rect 146 358 147 359
rect 145 358 146 359
rect 144 358 145 359
rect 143 358 144 359
rect 142 358 143 359
rect 141 358 142 359
rect 140 358 141 359
rect 139 358 140 359
rect 138 358 139 359
rect 137 358 138 359
rect 136 358 137 359
rect 135 358 136 359
rect 134 358 135 359
rect 133 358 134 359
rect 132 358 133 359
rect 131 358 132 359
rect 130 358 131 359
rect 129 358 130 359
rect 128 358 129 359
rect 127 358 128 359
rect 126 358 127 359
rect 125 358 126 359
rect 124 358 125 359
rect 123 358 124 359
rect 122 358 123 359
rect 121 358 122 359
rect 120 358 121 359
rect 119 358 120 359
rect 118 358 119 359
rect 117 358 118 359
rect 116 358 117 359
rect 115 358 116 359
rect 114 358 115 359
rect 113 358 114 359
rect 112 358 113 359
rect 111 358 112 359
rect 110 358 111 359
rect 109 358 110 359
rect 108 358 109 359
rect 107 358 108 359
rect 106 358 107 359
rect 105 358 106 359
rect 104 358 105 359
rect 103 358 104 359
rect 102 358 103 359
rect 101 358 102 359
rect 100 358 101 359
rect 71 358 72 359
rect 70 358 71 359
rect 69 358 70 359
rect 68 358 69 359
rect 67 358 68 359
rect 66 358 67 359
rect 65 358 66 359
rect 64 358 65 359
rect 63 358 64 359
rect 62 358 63 359
rect 61 358 62 359
rect 60 358 61 359
rect 54 358 55 359
rect 53 358 54 359
rect 52 358 53 359
rect 51 358 52 359
rect 50 358 51 359
rect 49 358 50 359
rect 13 358 14 359
rect 194 359 195 360
rect 193 359 194 360
rect 192 359 193 360
rect 191 359 192 360
rect 190 359 191 360
rect 189 359 190 360
rect 181 359 182 360
rect 180 359 181 360
rect 179 359 180 360
rect 178 359 179 360
rect 171 359 172 360
rect 170 359 171 360
rect 169 359 170 360
rect 168 359 169 360
rect 167 359 168 360
rect 147 359 148 360
rect 146 359 147 360
rect 145 359 146 360
rect 144 359 145 360
rect 143 359 144 360
rect 142 359 143 360
rect 141 359 142 360
rect 140 359 141 360
rect 139 359 140 360
rect 138 359 139 360
rect 137 359 138 360
rect 136 359 137 360
rect 135 359 136 360
rect 134 359 135 360
rect 133 359 134 360
rect 132 359 133 360
rect 131 359 132 360
rect 130 359 131 360
rect 129 359 130 360
rect 128 359 129 360
rect 127 359 128 360
rect 126 359 127 360
rect 125 359 126 360
rect 124 359 125 360
rect 123 359 124 360
rect 122 359 123 360
rect 121 359 122 360
rect 120 359 121 360
rect 119 359 120 360
rect 118 359 119 360
rect 117 359 118 360
rect 116 359 117 360
rect 115 359 116 360
rect 114 359 115 360
rect 113 359 114 360
rect 112 359 113 360
rect 111 359 112 360
rect 110 359 111 360
rect 109 359 110 360
rect 108 359 109 360
rect 107 359 108 360
rect 106 359 107 360
rect 105 359 106 360
rect 104 359 105 360
rect 103 359 104 360
rect 102 359 103 360
rect 101 359 102 360
rect 100 359 101 360
rect 72 359 73 360
rect 71 359 72 360
rect 70 359 71 360
rect 69 359 70 360
rect 68 359 69 360
rect 67 359 68 360
rect 66 359 67 360
rect 65 359 66 360
rect 64 359 65 360
rect 63 359 64 360
rect 62 359 63 360
rect 61 359 62 360
rect 60 359 61 360
rect 54 359 55 360
rect 53 359 54 360
rect 52 359 53 360
rect 51 359 52 360
rect 50 359 51 360
rect 49 359 50 360
rect 27 359 28 360
rect 26 359 27 360
rect 25 359 26 360
rect 192 360 193 361
rect 181 360 182 361
rect 180 360 181 361
rect 179 360 180 361
rect 178 360 179 361
rect 171 360 172 361
rect 170 360 171 361
rect 169 360 170 361
rect 168 360 169 361
rect 147 360 148 361
rect 146 360 147 361
rect 145 360 146 361
rect 144 360 145 361
rect 143 360 144 361
rect 142 360 143 361
rect 141 360 142 361
rect 140 360 141 361
rect 139 360 140 361
rect 138 360 139 361
rect 137 360 138 361
rect 136 360 137 361
rect 135 360 136 361
rect 134 360 135 361
rect 133 360 134 361
rect 132 360 133 361
rect 131 360 132 361
rect 130 360 131 361
rect 129 360 130 361
rect 128 360 129 361
rect 127 360 128 361
rect 126 360 127 361
rect 125 360 126 361
rect 124 360 125 361
rect 123 360 124 361
rect 122 360 123 361
rect 121 360 122 361
rect 120 360 121 361
rect 119 360 120 361
rect 118 360 119 361
rect 117 360 118 361
rect 116 360 117 361
rect 115 360 116 361
rect 114 360 115 361
rect 113 360 114 361
rect 112 360 113 361
rect 111 360 112 361
rect 110 360 111 361
rect 109 360 110 361
rect 108 360 109 361
rect 107 360 108 361
rect 106 360 107 361
rect 105 360 106 361
rect 104 360 105 361
rect 103 360 104 361
rect 102 360 103 361
rect 101 360 102 361
rect 100 360 101 361
rect 73 360 74 361
rect 72 360 73 361
rect 71 360 72 361
rect 70 360 71 361
rect 69 360 70 361
rect 68 360 69 361
rect 67 360 68 361
rect 66 360 67 361
rect 65 360 66 361
rect 64 360 65 361
rect 63 360 64 361
rect 62 360 63 361
rect 61 360 62 361
rect 60 360 61 361
rect 59 360 60 361
rect 55 360 56 361
rect 54 360 55 361
rect 53 360 54 361
rect 52 360 53 361
rect 51 360 52 361
rect 50 360 51 361
rect 49 360 50 361
rect 27 360 28 361
rect 26 360 27 361
rect 25 360 26 361
rect 24 360 25 361
rect 23 360 24 361
rect 22 360 23 361
rect 21 360 22 361
rect 194 361 195 362
rect 193 361 194 362
rect 191 361 192 362
rect 190 361 191 362
rect 189 361 190 362
rect 181 361 182 362
rect 180 361 181 362
rect 179 361 180 362
rect 178 361 179 362
rect 172 361 173 362
rect 171 361 172 362
rect 170 361 171 362
rect 169 361 170 362
rect 147 361 148 362
rect 146 361 147 362
rect 145 361 146 362
rect 144 361 145 362
rect 143 361 144 362
rect 142 361 143 362
rect 141 361 142 362
rect 140 361 141 362
rect 139 361 140 362
rect 138 361 139 362
rect 137 361 138 362
rect 136 361 137 362
rect 135 361 136 362
rect 134 361 135 362
rect 133 361 134 362
rect 132 361 133 362
rect 131 361 132 362
rect 130 361 131 362
rect 129 361 130 362
rect 128 361 129 362
rect 127 361 128 362
rect 126 361 127 362
rect 125 361 126 362
rect 124 361 125 362
rect 123 361 124 362
rect 122 361 123 362
rect 121 361 122 362
rect 120 361 121 362
rect 119 361 120 362
rect 118 361 119 362
rect 117 361 118 362
rect 116 361 117 362
rect 115 361 116 362
rect 114 361 115 362
rect 113 361 114 362
rect 112 361 113 362
rect 111 361 112 362
rect 110 361 111 362
rect 109 361 110 362
rect 108 361 109 362
rect 107 361 108 362
rect 106 361 107 362
rect 105 361 106 362
rect 104 361 105 362
rect 103 361 104 362
rect 102 361 103 362
rect 101 361 102 362
rect 100 361 101 362
rect 75 361 76 362
rect 74 361 75 362
rect 73 361 74 362
rect 72 361 73 362
rect 71 361 72 362
rect 70 361 71 362
rect 69 361 70 362
rect 68 361 69 362
rect 67 361 68 362
rect 66 361 67 362
rect 63 361 64 362
rect 62 361 63 362
rect 61 361 62 362
rect 60 361 61 362
rect 59 361 60 362
rect 58 361 59 362
rect 57 361 58 362
rect 56 361 57 362
rect 55 361 56 362
rect 54 361 55 362
rect 53 361 54 362
rect 52 361 53 362
rect 51 361 52 362
rect 50 361 51 362
rect 27 361 28 362
rect 26 361 27 362
rect 25 361 26 362
rect 24 361 25 362
rect 23 361 24 362
rect 22 361 23 362
rect 21 361 22 362
rect 20 361 21 362
rect 19 361 20 362
rect 18 361 19 362
rect 17 361 18 362
rect 16 361 17 362
rect 195 362 196 363
rect 194 362 195 363
rect 193 362 194 363
rect 192 362 193 363
rect 191 362 192 363
rect 190 362 191 363
rect 189 362 190 363
rect 181 362 182 363
rect 180 362 181 363
rect 179 362 180 363
rect 178 362 179 363
rect 172 362 173 363
rect 171 362 172 363
rect 170 362 171 363
rect 169 362 170 363
rect 147 362 148 363
rect 146 362 147 363
rect 145 362 146 363
rect 144 362 145 363
rect 143 362 144 363
rect 142 362 143 363
rect 141 362 142 363
rect 140 362 141 363
rect 139 362 140 363
rect 138 362 139 363
rect 137 362 138 363
rect 136 362 137 363
rect 135 362 136 363
rect 134 362 135 363
rect 133 362 134 363
rect 132 362 133 363
rect 131 362 132 363
rect 130 362 131 363
rect 129 362 130 363
rect 128 362 129 363
rect 127 362 128 363
rect 126 362 127 363
rect 125 362 126 363
rect 124 362 125 363
rect 123 362 124 363
rect 122 362 123 363
rect 121 362 122 363
rect 120 362 121 363
rect 119 362 120 363
rect 118 362 119 363
rect 117 362 118 363
rect 116 362 117 363
rect 115 362 116 363
rect 114 362 115 363
rect 113 362 114 363
rect 112 362 113 363
rect 111 362 112 363
rect 110 362 111 363
rect 109 362 110 363
rect 108 362 109 363
rect 107 362 108 363
rect 106 362 107 363
rect 105 362 106 363
rect 104 362 105 363
rect 103 362 104 363
rect 102 362 103 363
rect 101 362 102 363
rect 100 362 101 363
rect 76 362 77 363
rect 75 362 76 363
rect 74 362 75 363
rect 73 362 74 363
rect 72 362 73 363
rect 71 362 72 363
rect 70 362 71 363
rect 69 362 70 363
rect 68 362 69 363
rect 67 362 68 363
rect 63 362 64 363
rect 62 362 63 363
rect 61 362 62 363
rect 60 362 61 363
rect 59 362 60 363
rect 58 362 59 363
rect 57 362 58 363
rect 56 362 57 363
rect 55 362 56 363
rect 54 362 55 363
rect 53 362 54 363
rect 52 362 53 363
rect 51 362 52 363
rect 50 362 51 363
rect 26 362 27 363
rect 25 362 26 363
rect 24 362 25 363
rect 23 362 24 363
rect 22 362 23 363
rect 21 362 22 363
rect 20 362 21 363
rect 19 362 20 363
rect 18 362 19 363
rect 17 362 18 363
rect 16 362 17 363
rect 15 362 16 363
rect 14 362 15 363
rect 13 362 14 363
rect 194 363 195 364
rect 191 363 192 364
rect 190 363 191 364
rect 189 363 190 364
rect 181 363 182 364
rect 180 363 181 364
rect 179 363 180 364
rect 178 363 179 364
rect 170 363 171 364
rect 147 363 148 364
rect 146 363 147 364
rect 145 363 146 364
rect 144 363 145 364
rect 143 363 144 364
rect 142 363 143 364
rect 141 363 142 364
rect 140 363 141 364
rect 139 363 140 364
rect 138 363 139 364
rect 137 363 138 364
rect 136 363 137 364
rect 135 363 136 364
rect 134 363 135 364
rect 133 363 134 364
rect 132 363 133 364
rect 131 363 132 364
rect 130 363 131 364
rect 129 363 130 364
rect 128 363 129 364
rect 127 363 128 364
rect 126 363 127 364
rect 125 363 126 364
rect 124 363 125 364
rect 123 363 124 364
rect 122 363 123 364
rect 121 363 122 364
rect 120 363 121 364
rect 119 363 120 364
rect 118 363 119 364
rect 117 363 118 364
rect 116 363 117 364
rect 115 363 116 364
rect 114 363 115 364
rect 113 363 114 364
rect 112 363 113 364
rect 111 363 112 364
rect 110 363 111 364
rect 109 363 110 364
rect 108 363 109 364
rect 107 363 108 364
rect 106 363 107 364
rect 105 363 106 364
rect 104 363 105 364
rect 103 363 104 364
rect 102 363 103 364
rect 101 363 102 364
rect 100 363 101 364
rect 76 363 77 364
rect 75 363 76 364
rect 74 363 75 364
rect 73 363 74 364
rect 72 363 73 364
rect 71 363 72 364
rect 70 363 71 364
rect 69 363 70 364
rect 68 363 69 364
rect 62 363 63 364
rect 61 363 62 364
rect 60 363 61 364
rect 59 363 60 364
rect 58 363 59 364
rect 57 363 58 364
rect 56 363 57 364
rect 55 363 56 364
rect 54 363 55 364
rect 53 363 54 364
rect 52 363 53 364
rect 51 363 52 364
rect 22 363 23 364
rect 21 363 22 364
rect 20 363 21 364
rect 19 363 20 364
rect 18 363 19 364
rect 17 363 18 364
rect 16 363 17 364
rect 15 363 16 364
rect 14 363 15 364
rect 13 363 14 364
rect 12 363 13 364
rect 190 364 191 365
rect 189 364 190 365
rect 181 364 182 365
rect 180 364 181 365
rect 179 364 180 365
rect 178 364 179 365
rect 147 364 148 365
rect 146 364 147 365
rect 145 364 146 365
rect 144 364 145 365
rect 143 364 144 365
rect 142 364 143 365
rect 141 364 142 365
rect 140 364 141 365
rect 139 364 140 365
rect 138 364 139 365
rect 137 364 138 365
rect 136 364 137 365
rect 135 364 136 365
rect 134 364 135 365
rect 133 364 134 365
rect 132 364 133 365
rect 131 364 132 365
rect 130 364 131 365
rect 129 364 130 365
rect 128 364 129 365
rect 127 364 128 365
rect 126 364 127 365
rect 125 364 126 365
rect 124 364 125 365
rect 123 364 124 365
rect 122 364 123 365
rect 121 364 122 365
rect 120 364 121 365
rect 119 364 120 365
rect 118 364 119 365
rect 117 364 118 365
rect 116 364 117 365
rect 115 364 116 365
rect 114 364 115 365
rect 113 364 114 365
rect 112 364 113 365
rect 111 364 112 365
rect 110 364 111 365
rect 109 364 110 365
rect 108 364 109 365
rect 107 364 108 365
rect 106 364 107 365
rect 105 364 106 365
rect 104 364 105 365
rect 103 364 104 365
rect 102 364 103 365
rect 101 364 102 365
rect 100 364 101 365
rect 76 364 77 365
rect 75 364 76 365
rect 74 364 75 365
rect 73 364 74 365
rect 72 364 73 365
rect 71 364 72 365
rect 70 364 71 365
rect 69 364 70 365
rect 62 364 63 365
rect 61 364 62 365
rect 60 364 61 365
rect 59 364 60 365
rect 58 364 59 365
rect 57 364 58 365
rect 56 364 57 365
rect 55 364 56 365
rect 54 364 55 365
rect 53 364 54 365
rect 52 364 53 365
rect 51 364 52 365
rect 21 364 22 365
rect 20 364 21 365
rect 19 364 20 365
rect 17 364 18 365
rect 16 364 17 365
rect 15 364 16 365
rect 14 364 15 365
rect 13 364 14 365
rect 12 364 13 365
rect 194 365 195 366
rect 193 365 194 366
rect 192 365 193 366
rect 191 365 192 366
rect 190 365 191 366
rect 189 365 190 366
rect 181 365 182 366
rect 180 365 181 366
rect 179 365 180 366
rect 178 365 179 366
rect 147 365 148 366
rect 146 365 147 366
rect 145 365 146 366
rect 144 365 145 366
rect 143 365 144 366
rect 142 365 143 366
rect 141 365 142 366
rect 140 365 141 366
rect 139 365 140 366
rect 138 365 139 366
rect 137 365 138 366
rect 136 365 137 366
rect 135 365 136 366
rect 134 365 135 366
rect 133 365 134 366
rect 132 365 133 366
rect 131 365 132 366
rect 130 365 131 366
rect 129 365 130 366
rect 128 365 129 366
rect 127 365 128 366
rect 126 365 127 366
rect 125 365 126 366
rect 124 365 125 366
rect 123 365 124 366
rect 122 365 123 366
rect 121 365 122 366
rect 120 365 121 366
rect 119 365 120 366
rect 118 365 119 366
rect 117 365 118 366
rect 116 365 117 366
rect 115 365 116 366
rect 114 365 115 366
rect 113 365 114 366
rect 112 365 113 366
rect 111 365 112 366
rect 110 365 111 366
rect 109 365 110 366
rect 108 365 109 366
rect 107 365 108 366
rect 106 365 107 366
rect 105 365 106 366
rect 104 365 105 366
rect 103 365 104 366
rect 102 365 103 366
rect 101 365 102 366
rect 100 365 101 366
rect 76 365 77 366
rect 75 365 76 366
rect 74 365 75 366
rect 73 365 74 366
rect 72 365 73 366
rect 71 365 72 366
rect 61 365 62 366
rect 60 365 61 366
rect 59 365 60 366
rect 58 365 59 366
rect 57 365 58 366
rect 56 365 57 366
rect 55 365 56 366
rect 54 365 55 366
rect 53 365 54 366
rect 52 365 53 366
rect 21 365 22 366
rect 20 365 21 366
rect 19 365 20 366
rect 14 365 15 366
rect 13 365 14 366
rect 12 365 13 366
rect 195 366 196 367
rect 194 366 195 367
rect 193 366 194 367
rect 192 366 193 367
rect 191 366 192 367
rect 190 366 191 367
rect 189 366 190 367
rect 181 366 182 367
rect 180 366 181 367
rect 179 366 180 367
rect 178 366 179 367
rect 175 366 176 367
rect 174 366 175 367
rect 173 366 174 367
rect 172 366 173 367
rect 171 366 172 367
rect 170 366 171 367
rect 169 366 170 367
rect 168 366 169 367
rect 167 366 168 367
rect 166 366 167 367
rect 165 366 166 367
rect 164 366 165 367
rect 163 366 164 367
rect 162 366 163 367
rect 161 366 162 367
rect 160 366 161 367
rect 147 366 148 367
rect 146 366 147 367
rect 145 366 146 367
rect 144 366 145 367
rect 143 366 144 367
rect 142 366 143 367
rect 141 366 142 367
rect 140 366 141 367
rect 139 366 140 367
rect 138 366 139 367
rect 137 366 138 367
rect 136 366 137 367
rect 135 366 136 367
rect 134 366 135 367
rect 133 366 134 367
rect 132 366 133 367
rect 131 366 132 367
rect 130 366 131 367
rect 129 366 130 367
rect 128 366 129 367
rect 127 366 128 367
rect 126 366 127 367
rect 125 366 126 367
rect 124 366 125 367
rect 123 366 124 367
rect 122 366 123 367
rect 121 366 122 367
rect 120 366 121 367
rect 119 366 120 367
rect 118 366 119 367
rect 117 366 118 367
rect 116 366 117 367
rect 115 366 116 367
rect 114 366 115 367
rect 113 366 114 367
rect 112 366 113 367
rect 111 366 112 367
rect 110 366 111 367
rect 109 366 110 367
rect 108 366 109 367
rect 107 366 108 367
rect 106 366 107 367
rect 105 366 106 367
rect 104 366 105 367
rect 103 366 104 367
rect 102 366 103 367
rect 101 366 102 367
rect 100 366 101 367
rect 76 366 77 367
rect 75 366 76 367
rect 74 366 75 367
rect 73 366 74 367
rect 59 366 60 367
rect 58 366 59 367
rect 57 366 58 367
rect 56 366 57 367
rect 55 366 56 367
rect 54 366 55 367
rect 21 366 22 367
rect 20 366 21 367
rect 19 366 20 367
rect 14 366 15 367
rect 13 366 14 367
rect 12 366 13 367
rect 181 367 182 368
rect 180 367 181 368
rect 179 367 180 368
rect 178 367 179 368
rect 175 367 176 368
rect 174 367 175 368
rect 173 367 174 368
rect 172 367 173 368
rect 171 367 172 368
rect 170 367 171 368
rect 169 367 170 368
rect 168 367 169 368
rect 167 367 168 368
rect 166 367 167 368
rect 165 367 166 368
rect 164 367 165 368
rect 163 367 164 368
rect 162 367 163 368
rect 161 367 162 368
rect 160 367 161 368
rect 147 367 148 368
rect 146 367 147 368
rect 145 367 146 368
rect 144 367 145 368
rect 143 367 144 368
rect 142 367 143 368
rect 141 367 142 368
rect 140 367 141 368
rect 139 367 140 368
rect 138 367 139 368
rect 137 367 138 368
rect 136 367 137 368
rect 135 367 136 368
rect 134 367 135 368
rect 133 367 134 368
rect 132 367 133 368
rect 131 367 132 368
rect 130 367 131 368
rect 129 367 130 368
rect 128 367 129 368
rect 127 367 128 368
rect 126 367 127 368
rect 125 367 126 368
rect 124 367 125 368
rect 123 367 124 368
rect 122 367 123 368
rect 121 367 122 368
rect 120 367 121 368
rect 119 367 120 368
rect 118 367 119 368
rect 117 367 118 368
rect 116 367 117 368
rect 115 367 116 368
rect 114 367 115 368
rect 113 367 114 368
rect 112 367 113 368
rect 111 367 112 368
rect 110 367 111 368
rect 109 367 110 368
rect 108 367 109 368
rect 107 367 108 368
rect 106 367 107 368
rect 105 367 106 368
rect 104 367 105 368
rect 103 367 104 368
rect 102 367 103 368
rect 101 367 102 368
rect 100 367 101 368
rect 76 367 77 368
rect 75 367 76 368
rect 74 367 75 368
rect 21 367 22 368
rect 20 367 21 368
rect 19 367 20 368
rect 14 367 15 368
rect 13 367 14 368
rect 12 367 13 368
rect 194 368 195 369
rect 191 368 192 369
rect 190 368 191 369
rect 181 368 182 369
rect 180 368 181 369
rect 179 368 180 369
rect 178 368 179 369
rect 175 368 176 369
rect 174 368 175 369
rect 173 368 174 369
rect 172 368 173 369
rect 171 368 172 369
rect 170 368 171 369
rect 169 368 170 369
rect 168 368 169 369
rect 167 368 168 369
rect 166 368 167 369
rect 165 368 166 369
rect 164 368 165 369
rect 163 368 164 369
rect 162 368 163 369
rect 161 368 162 369
rect 160 368 161 369
rect 147 368 148 369
rect 146 368 147 369
rect 145 368 146 369
rect 144 368 145 369
rect 143 368 144 369
rect 142 368 143 369
rect 141 368 142 369
rect 140 368 141 369
rect 139 368 140 369
rect 138 368 139 369
rect 137 368 138 369
rect 136 368 137 369
rect 135 368 136 369
rect 134 368 135 369
rect 133 368 134 369
rect 132 368 133 369
rect 131 368 132 369
rect 130 368 131 369
rect 129 368 130 369
rect 128 368 129 369
rect 127 368 128 369
rect 126 368 127 369
rect 125 368 126 369
rect 124 368 125 369
rect 123 368 124 369
rect 122 368 123 369
rect 121 368 122 369
rect 120 368 121 369
rect 119 368 120 369
rect 118 368 119 369
rect 117 368 118 369
rect 116 368 117 369
rect 115 368 116 369
rect 114 368 115 369
rect 113 368 114 369
rect 112 368 113 369
rect 111 368 112 369
rect 110 368 111 369
rect 109 368 110 369
rect 108 368 109 369
rect 107 368 108 369
rect 106 368 107 369
rect 105 368 106 369
rect 104 368 105 369
rect 103 368 104 369
rect 102 368 103 369
rect 101 368 102 369
rect 100 368 101 369
rect 76 368 77 369
rect 21 368 22 369
rect 20 368 21 369
rect 19 368 20 369
rect 14 368 15 369
rect 13 368 14 369
rect 12 368 13 369
rect 195 369 196 370
rect 194 369 195 370
rect 192 369 193 370
rect 191 369 192 370
rect 190 369 191 370
rect 189 369 190 370
rect 181 369 182 370
rect 180 369 181 370
rect 179 369 180 370
rect 178 369 179 370
rect 175 369 176 370
rect 174 369 175 370
rect 173 369 174 370
rect 172 369 173 370
rect 171 369 172 370
rect 170 369 171 370
rect 169 369 170 370
rect 168 369 169 370
rect 167 369 168 370
rect 166 369 167 370
rect 165 369 166 370
rect 164 369 165 370
rect 163 369 164 370
rect 162 369 163 370
rect 161 369 162 370
rect 160 369 161 370
rect 147 369 148 370
rect 146 369 147 370
rect 145 369 146 370
rect 144 369 145 370
rect 143 369 144 370
rect 142 369 143 370
rect 141 369 142 370
rect 140 369 141 370
rect 139 369 140 370
rect 138 369 139 370
rect 137 369 138 370
rect 136 369 137 370
rect 135 369 136 370
rect 134 369 135 370
rect 133 369 134 370
rect 132 369 133 370
rect 131 369 132 370
rect 130 369 131 370
rect 129 369 130 370
rect 128 369 129 370
rect 127 369 128 370
rect 126 369 127 370
rect 125 369 126 370
rect 124 369 125 370
rect 123 369 124 370
rect 122 369 123 370
rect 121 369 122 370
rect 120 369 121 370
rect 119 369 120 370
rect 118 369 119 370
rect 117 369 118 370
rect 116 369 117 370
rect 115 369 116 370
rect 114 369 115 370
rect 113 369 114 370
rect 112 369 113 370
rect 111 369 112 370
rect 110 369 111 370
rect 109 369 110 370
rect 108 369 109 370
rect 107 369 108 370
rect 106 369 107 370
rect 105 369 106 370
rect 104 369 105 370
rect 103 369 104 370
rect 102 369 103 370
rect 101 369 102 370
rect 100 369 101 370
rect 21 369 22 370
rect 20 369 21 370
rect 19 369 20 370
rect 18 369 19 370
rect 15 369 16 370
rect 14 369 15 370
rect 13 369 14 370
rect 195 370 196 371
rect 194 370 195 371
rect 193 370 194 371
rect 192 370 193 371
rect 191 370 192 371
rect 190 370 191 371
rect 189 370 190 371
rect 180 370 181 371
rect 179 370 180 371
rect 147 370 148 371
rect 146 370 147 371
rect 145 370 146 371
rect 144 370 145 371
rect 143 370 144 371
rect 142 370 143 371
rect 141 370 142 371
rect 140 370 141 371
rect 139 370 140 371
rect 138 370 139 371
rect 137 370 138 371
rect 136 370 137 371
rect 135 370 136 371
rect 134 370 135 371
rect 133 370 134 371
rect 132 370 133 371
rect 131 370 132 371
rect 130 370 131 371
rect 129 370 130 371
rect 128 370 129 371
rect 127 370 128 371
rect 126 370 127 371
rect 125 370 126 371
rect 124 370 125 371
rect 123 370 124 371
rect 122 370 123 371
rect 121 370 122 371
rect 120 370 121 371
rect 119 370 120 371
rect 118 370 119 371
rect 117 370 118 371
rect 116 370 117 371
rect 115 370 116 371
rect 114 370 115 371
rect 113 370 114 371
rect 112 370 113 371
rect 111 370 112 371
rect 110 370 111 371
rect 109 370 110 371
rect 108 370 109 371
rect 107 370 108 371
rect 106 370 107 371
rect 105 370 106 371
rect 104 370 105 371
rect 103 370 104 371
rect 102 370 103 371
rect 101 370 102 371
rect 100 370 101 371
rect 20 370 21 371
rect 19 370 20 371
rect 18 370 19 371
rect 17 370 18 371
rect 16 370 17 371
rect 15 370 16 371
rect 14 370 15 371
rect 13 370 14 371
rect 194 371 195 372
rect 193 371 194 372
rect 192 371 193 372
rect 190 371 191 372
rect 189 371 190 372
rect 147 371 148 372
rect 146 371 147 372
rect 145 371 146 372
rect 144 371 145 372
rect 143 371 144 372
rect 142 371 143 372
rect 141 371 142 372
rect 140 371 141 372
rect 139 371 140 372
rect 138 371 139 372
rect 137 371 138 372
rect 136 371 137 372
rect 135 371 136 372
rect 134 371 135 372
rect 133 371 134 372
rect 132 371 133 372
rect 131 371 132 372
rect 130 371 131 372
rect 129 371 130 372
rect 128 371 129 372
rect 127 371 128 372
rect 126 371 127 372
rect 125 371 126 372
rect 124 371 125 372
rect 123 371 124 372
rect 122 371 123 372
rect 121 371 122 372
rect 120 371 121 372
rect 119 371 120 372
rect 118 371 119 372
rect 117 371 118 372
rect 116 371 117 372
rect 115 371 116 372
rect 114 371 115 372
rect 113 371 114 372
rect 112 371 113 372
rect 111 371 112 372
rect 110 371 111 372
rect 109 371 110 372
rect 108 371 109 372
rect 107 371 108 372
rect 106 371 107 372
rect 105 371 106 372
rect 104 371 105 372
rect 103 371 104 372
rect 102 371 103 372
rect 101 371 102 372
rect 100 371 101 372
rect 72 371 73 372
rect 71 371 72 372
rect 70 371 71 372
rect 69 371 70 372
rect 68 371 69 372
rect 67 371 68 372
rect 66 371 67 372
rect 65 371 66 372
rect 57 371 58 372
rect 56 371 57 372
rect 55 371 56 372
rect 54 371 55 372
rect 20 371 21 372
rect 19 371 20 372
rect 18 371 19 372
rect 17 371 18 372
rect 16 371 17 372
rect 15 371 16 372
rect 14 371 15 372
rect 13 371 14 372
rect 194 372 195 373
rect 193 372 194 373
rect 192 372 193 373
rect 189 372 190 373
rect 147 372 148 373
rect 146 372 147 373
rect 145 372 146 373
rect 144 372 145 373
rect 143 372 144 373
rect 142 372 143 373
rect 141 372 142 373
rect 140 372 141 373
rect 139 372 140 373
rect 138 372 139 373
rect 137 372 138 373
rect 136 372 137 373
rect 135 372 136 373
rect 134 372 135 373
rect 133 372 134 373
rect 132 372 133 373
rect 131 372 132 373
rect 130 372 131 373
rect 129 372 130 373
rect 128 372 129 373
rect 127 372 128 373
rect 126 372 127 373
rect 125 372 126 373
rect 124 372 125 373
rect 123 372 124 373
rect 122 372 123 373
rect 121 372 122 373
rect 120 372 121 373
rect 119 372 120 373
rect 118 372 119 373
rect 117 372 118 373
rect 116 372 117 373
rect 115 372 116 373
rect 114 372 115 373
rect 113 372 114 373
rect 112 372 113 373
rect 111 372 112 373
rect 110 372 111 373
rect 109 372 110 373
rect 108 372 109 373
rect 107 372 108 373
rect 106 372 107 373
rect 105 372 106 373
rect 104 372 105 373
rect 103 372 104 373
rect 102 372 103 373
rect 101 372 102 373
rect 100 372 101 373
rect 73 372 74 373
rect 72 372 73 373
rect 71 372 72 373
rect 70 372 71 373
rect 69 372 70 373
rect 68 372 69 373
rect 67 372 68 373
rect 66 372 67 373
rect 65 372 66 373
rect 64 372 65 373
rect 59 372 60 373
rect 58 372 59 373
rect 57 372 58 373
rect 56 372 57 373
rect 55 372 56 373
rect 54 372 55 373
rect 53 372 54 373
rect 52 372 53 373
rect 18 372 19 373
rect 17 372 18 373
rect 16 372 17 373
rect 15 372 16 373
rect 14 372 15 373
rect 147 373 148 374
rect 146 373 147 374
rect 145 373 146 374
rect 144 373 145 374
rect 143 373 144 374
rect 142 373 143 374
rect 141 373 142 374
rect 140 373 141 374
rect 139 373 140 374
rect 138 373 139 374
rect 137 373 138 374
rect 136 373 137 374
rect 135 373 136 374
rect 134 373 135 374
rect 133 373 134 374
rect 132 373 133 374
rect 131 373 132 374
rect 130 373 131 374
rect 129 373 130 374
rect 128 373 129 374
rect 127 373 128 374
rect 126 373 127 374
rect 125 373 126 374
rect 124 373 125 374
rect 123 373 124 374
rect 122 373 123 374
rect 121 373 122 374
rect 120 373 121 374
rect 119 373 120 374
rect 118 373 119 374
rect 117 373 118 374
rect 116 373 117 374
rect 115 373 116 374
rect 114 373 115 374
rect 113 373 114 374
rect 112 373 113 374
rect 111 373 112 374
rect 110 373 111 374
rect 109 373 110 374
rect 108 373 109 374
rect 107 373 108 374
rect 106 373 107 374
rect 105 373 106 374
rect 104 373 105 374
rect 103 373 104 374
rect 102 373 103 374
rect 101 373 102 374
rect 100 373 101 374
rect 74 373 75 374
rect 73 373 74 374
rect 72 373 73 374
rect 71 373 72 374
rect 70 373 71 374
rect 69 373 70 374
rect 68 373 69 374
rect 67 373 68 374
rect 66 373 67 374
rect 65 373 66 374
rect 64 373 65 374
rect 63 373 64 374
rect 60 373 61 374
rect 59 373 60 374
rect 58 373 59 374
rect 57 373 58 374
rect 56 373 57 374
rect 55 373 56 374
rect 54 373 55 374
rect 53 373 54 374
rect 52 373 53 374
rect 51 373 52 374
rect 147 374 148 375
rect 146 374 147 375
rect 145 374 146 375
rect 144 374 145 375
rect 143 374 144 375
rect 142 374 143 375
rect 141 374 142 375
rect 140 374 141 375
rect 139 374 140 375
rect 138 374 139 375
rect 137 374 138 375
rect 136 374 137 375
rect 135 374 136 375
rect 134 374 135 375
rect 133 374 134 375
rect 132 374 133 375
rect 131 374 132 375
rect 130 374 131 375
rect 129 374 130 375
rect 128 374 129 375
rect 127 374 128 375
rect 126 374 127 375
rect 125 374 126 375
rect 124 374 125 375
rect 123 374 124 375
rect 122 374 123 375
rect 121 374 122 375
rect 120 374 121 375
rect 119 374 120 375
rect 118 374 119 375
rect 117 374 118 375
rect 116 374 117 375
rect 115 374 116 375
rect 114 374 115 375
rect 113 374 114 375
rect 112 374 113 375
rect 111 374 112 375
rect 110 374 111 375
rect 109 374 110 375
rect 108 374 109 375
rect 107 374 108 375
rect 106 374 107 375
rect 105 374 106 375
rect 104 374 105 375
rect 103 374 104 375
rect 102 374 103 375
rect 101 374 102 375
rect 100 374 101 375
rect 75 374 76 375
rect 74 374 75 375
rect 73 374 74 375
rect 72 374 73 375
rect 71 374 72 375
rect 70 374 71 375
rect 69 374 70 375
rect 68 374 69 375
rect 67 374 68 375
rect 66 374 67 375
rect 65 374 66 375
rect 64 374 65 375
rect 63 374 64 375
rect 62 374 63 375
rect 61 374 62 375
rect 60 374 61 375
rect 59 374 60 375
rect 58 374 59 375
rect 57 374 58 375
rect 56 374 57 375
rect 55 374 56 375
rect 54 374 55 375
rect 53 374 54 375
rect 52 374 53 375
rect 51 374 52 375
rect 50 374 51 375
rect 147 375 148 376
rect 146 375 147 376
rect 145 375 146 376
rect 144 375 145 376
rect 143 375 144 376
rect 142 375 143 376
rect 141 375 142 376
rect 140 375 141 376
rect 139 375 140 376
rect 138 375 139 376
rect 137 375 138 376
rect 136 375 137 376
rect 135 375 136 376
rect 134 375 135 376
rect 133 375 134 376
rect 132 375 133 376
rect 131 375 132 376
rect 130 375 131 376
rect 129 375 130 376
rect 128 375 129 376
rect 127 375 128 376
rect 126 375 127 376
rect 125 375 126 376
rect 124 375 125 376
rect 123 375 124 376
rect 122 375 123 376
rect 121 375 122 376
rect 120 375 121 376
rect 119 375 120 376
rect 118 375 119 376
rect 117 375 118 376
rect 116 375 117 376
rect 115 375 116 376
rect 114 375 115 376
rect 113 375 114 376
rect 112 375 113 376
rect 111 375 112 376
rect 110 375 111 376
rect 109 375 110 376
rect 108 375 109 376
rect 107 375 108 376
rect 106 375 107 376
rect 105 375 106 376
rect 104 375 105 376
rect 103 375 104 376
rect 102 375 103 376
rect 101 375 102 376
rect 100 375 101 376
rect 76 375 77 376
rect 75 375 76 376
rect 74 375 75 376
rect 73 375 74 376
rect 72 375 73 376
rect 71 375 72 376
rect 70 375 71 376
rect 69 375 70 376
rect 68 375 69 376
rect 67 375 68 376
rect 66 375 67 376
rect 65 375 66 376
rect 64 375 65 376
rect 63 375 64 376
rect 62 375 63 376
rect 61 375 62 376
rect 60 375 61 376
rect 59 375 60 376
rect 58 375 59 376
rect 57 375 58 376
rect 56 375 57 376
rect 55 375 56 376
rect 54 375 55 376
rect 53 375 54 376
rect 52 375 53 376
rect 51 375 52 376
rect 50 375 51 376
rect 27 375 28 376
rect 26 375 27 376
rect 25 375 26 376
rect 24 375 25 376
rect 23 375 24 376
rect 22 375 23 376
rect 21 375 22 376
rect 20 375 21 376
rect 19 375 20 376
rect 18 375 19 376
rect 17 375 18 376
rect 16 375 17 376
rect 15 375 16 376
rect 14 375 15 376
rect 13 375 14 376
rect 12 375 13 376
rect 110 376 111 377
rect 109 376 110 377
rect 108 376 109 377
rect 107 376 108 377
rect 106 376 107 377
rect 105 376 106 377
rect 104 376 105 377
rect 103 376 104 377
rect 102 376 103 377
rect 101 376 102 377
rect 100 376 101 377
rect 76 376 77 377
rect 75 376 76 377
rect 74 376 75 377
rect 73 376 74 377
rect 72 376 73 377
rect 71 376 72 377
rect 65 376 66 377
rect 64 376 65 377
rect 63 376 64 377
rect 62 376 63 377
rect 61 376 62 377
rect 60 376 61 377
rect 59 376 60 377
rect 58 376 59 377
rect 57 376 58 377
rect 56 376 57 377
rect 55 376 56 377
rect 54 376 55 377
rect 53 376 54 377
rect 52 376 53 377
rect 51 376 52 377
rect 50 376 51 377
rect 27 376 28 377
rect 26 376 27 377
rect 25 376 26 377
rect 24 376 25 377
rect 23 376 24 377
rect 22 376 23 377
rect 21 376 22 377
rect 20 376 21 377
rect 19 376 20 377
rect 18 376 19 377
rect 17 376 18 377
rect 16 376 17 377
rect 15 376 16 377
rect 14 376 15 377
rect 13 376 14 377
rect 12 376 13 377
rect 195 377 196 378
rect 194 377 195 378
rect 193 377 194 378
rect 192 377 193 378
rect 191 377 192 378
rect 190 377 191 378
rect 189 377 190 378
rect 188 377 189 378
rect 187 377 188 378
rect 110 377 111 378
rect 109 377 110 378
rect 108 377 109 378
rect 107 377 108 378
rect 106 377 107 378
rect 105 377 106 378
rect 104 377 105 378
rect 103 377 104 378
rect 102 377 103 378
rect 101 377 102 378
rect 100 377 101 378
rect 76 377 77 378
rect 75 377 76 378
rect 74 377 75 378
rect 73 377 74 378
rect 72 377 73 378
rect 64 377 65 378
rect 63 377 64 378
rect 62 377 63 378
rect 61 377 62 378
rect 60 377 61 378
rect 59 377 60 378
rect 53 377 54 378
rect 52 377 53 378
rect 51 377 52 378
rect 50 377 51 378
rect 49 377 50 378
rect 27 377 28 378
rect 26 377 27 378
rect 25 377 26 378
rect 24 377 25 378
rect 23 377 24 378
rect 22 377 23 378
rect 21 377 22 378
rect 20 377 21 378
rect 19 377 20 378
rect 18 377 19 378
rect 17 377 18 378
rect 16 377 17 378
rect 15 377 16 378
rect 14 377 15 378
rect 13 377 14 378
rect 194 378 195 379
rect 193 378 194 379
rect 192 378 193 379
rect 191 378 192 379
rect 190 378 191 379
rect 189 378 190 379
rect 188 378 189 379
rect 187 378 188 379
rect 110 378 111 379
rect 109 378 110 379
rect 108 378 109 379
rect 107 378 108 379
rect 106 378 107 379
rect 105 378 106 379
rect 104 378 105 379
rect 103 378 104 379
rect 102 378 103 379
rect 101 378 102 379
rect 100 378 101 379
rect 76 378 77 379
rect 75 378 76 379
rect 74 378 75 379
rect 73 378 74 379
rect 63 378 64 379
rect 62 378 63 379
rect 61 378 62 379
rect 60 378 61 379
rect 53 378 54 379
rect 52 378 53 379
rect 51 378 52 379
rect 50 378 51 379
rect 49 378 50 379
rect 27 378 28 379
rect 26 378 27 379
rect 25 378 26 379
rect 24 378 25 379
rect 23 378 24 379
rect 22 378 23 379
rect 191 379 192 380
rect 190 379 191 380
rect 187 379 188 380
rect 110 379 111 380
rect 109 379 110 380
rect 108 379 109 380
rect 107 379 108 380
rect 106 379 107 380
rect 105 379 106 380
rect 104 379 105 380
rect 103 379 104 380
rect 102 379 103 380
rect 101 379 102 380
rect 100 379 101 380
rect 76 379 77 380
rect 75 379 76 380
rect 74 379 75 380
rect 73 379 74 380
rect 63 379 64 380
rect 62 379 63 380
rect 61 379 62 380
rect 60 379 61 380
rect 53 379 54 380
rect 52 379 53 380
rect 51 379 52 380
rect 50 379 51 380
rect 49 379 50 380
rect 26 379 27 380
rect 25 379 26 380
rect 24 379 25 380
rect 23 379 24 380
rect 22 379 23 380
rect 21 379 22 380
rect 20 379 21 380
rect 192 380 193 381
rect 191 380 192 381
rect 190 380 191 381
rect 188 380 189 381
rect 187 380 188 381
rect 110 380 111 381
rect 109 380 110 381
rect 108 380 109 381
rect 107 380 108 381
rect 106 380 107 381
rect 105 380 106 381
rect 104 380 105 381
rect 103 380 104 381
rect 102 380 103 381
rect 101 380 102 381
rect 100 380 101 381
rect 76 380 77 381
rect 75 380 76 381
rect 74 380 75 381
rect 73 380 74 381
rect 63 380 64 381
rect 62 380 63 381
rect 61 380 62 381
rect 60 380 61 381
rect 53 380 54 381
rect 52 380 53 381
rect 51 380 52 381
rect 50 380 51 381
rect 49 380 50 381
rect 24 380 25 381
rect 23 380 24 381
rect 22 380 23 381
rect 21 380 22 381
rect 20 380 21 381
rect 19 380 20 381
rect 18 380 19 381
rect 194 381 195 382
rect 193 381 194 382
rect 192 381 193 382
rect 191 381 192 382
rect 190 381 191 382
rect 189 381 190 382
rect 188 381 189 382
rect 187 381 188 382
rect 110 381 111 382
rect 109 381 110 382
rect 108 381 109 382
rect 107 381 108 382
rect 106 381 107 382
rect 105 381 106 382
rect 104 381 105 382
rect 103 381 104 382
rect 102 381 103 382
rect 101 381 102 382
rect 100 381 101 382
rect 76 381 77 382
rect 75 381 76 382
rect 74 381 75 382
rect 73 381 74 382
rect 64 381 65 382
rect 63 381 64 382
rect 62 381 63 382
rect 61 381 62 382
rect 60 381 61 382
rect 59 381 60 382
rect 53 381 54 382
rect 52 381 53 382
rect 51 381 52 382
rect 50 381 51 382
rect 49 381 50 382
rect 22 381 23 382
rect 21 381 22 382
rect 20 381 21 382
rect 19 381 20 382
rect 18 381 19 382
rect 17 381 18 382
rect 16 381 17 382
rect 194 382 195 383
rect 193 382 194 383
rect 192 382 193 383
rect 190 382 191 383
rect 189 382 190 383
rect 188 382 189 383
rect 187 382 188 383
rect 110 382 111 383
rect 109 382 110 383
rect 108 382 109 383
rect 107 382 108 383
rect 106 382 107 383
rect 105 382 106 383
rect 104 382 105 383
rect 103 382 104 383
rect 102 382 103 383
rect 101 382 102 383
rect 100 382 101 383
rect 76 382 77 383
rect 75 382 76 383
rect 74 382 75 383
rect 73 382 74 383
rect 72 382 73 383
rect 65 382 66 383
rect 64 382 65 383
rect 63 382 64 383
rect 62 382 63 383
rect 61 382 62 383
rect 60 382 61 383
rect 59 382 60 383
rect 58 382 59 383
rect 54 382 55 383
rect 53 382 54 383
rect 52 382 53 383
rect 51 382 52 383
rect 50 382 51 383
rect 49 382 50 383
rect 20 382 21 383
rect 19 382 20 383
rect 18 382 19 383
rect 17 382 18 383
rect 16 382 17 383
rect 15 382 16 383
rect 14 382 15 383
rect 194 383 195 384
rect 192 383 193 384
rect 168 383 169 384
rect 167 383 168 384
rect 166 383 167 384
rect 165 383 166 384
rect 164 383 165 384
rect 163 383 164 384
rect 110 383 111 384
rect 109 383 110 384
rect 108 383 109 384
rect 107 383 108 384
rect 106 383 107 384
rect 105 383 106 384
rect 104 383 105 384
rect 103 383 104 384
rect 102 383 103 384
rect 101 383 102 384
rect 100 383 101 384
rect 76 383 77 384
rect 75 383 76 384
rect 74 383 75 384
rect 73 383 74 384
rect 72 383 73 384
rect 71 383 72 384
rect 70 383 71 384
rect 69 383 70 384
rect 68 383 69 384
rect 67 383 68 384
rect 66 383 67 384
rect 65 383 66 384
rect 64 383 65 384
rect 63 383 64 384
rect 62 383 63 384
rect 61 383 62 384
rect 60 383 61 384
rect 59 383 60 384
rect 58 383 59 384
rect 57 383 58 384
rect 56 383 57 384
rect 55 383 56 384
rect 54 383 55 384
rect 53 383 54 384
rect 52 383 53 384
rect 51 383 52 384
rect 50 383 51 384
rect 17 383 18 384
rect 16 383 17 384
rect 15 383 16 384
rect 14 383 15 384
rect 13 383 14 384
rect 194 384 195 385
rect 193 384 194 385
rect 192 384 193 385
rect 191 384 192 385
rect 190 384 191 385
rect 169 384 170 385
rect 168 384 169 385
rect 167 384 168 385
rect 166 384 167 385
rect 165 384 166 385
rect 164 384 165 385
rect 163 384 164 385
rect 162 384 163 385
rect 126 384 127 385
rect 110 384 111 385
rect 109 384 110 385
rect 108 384 109 385
rect 107 384 108 385
rect 106 384 107 385
rect 105 384 106 385
rect 104 384 105 385
rect 103 384 104 385
rect 102 384 103 385
rect 101 384 102 385
rect 100 384 101 385
rect 75 384 76 385
rect 74 384 75 385
rect 73 384 74 385
rect 72 384 73 385
rect 71 384 72 385
rect 70 384 71 385
rect 69 384 70 385
rect 68 384 69 385
rect 67 384 68 385
rect 66 384 67 385
rect 65 384 66 385
rect 64 384 65 385
rect 63 384 64 385
rect 62 384 63 385
rect 61 384 62 385
rect 60 384 61 385
rect 59 384 60 385
rect 58 384 59 385
rect 57 384 58 385
rect 56 384 57 385
rect 55 384 56 385
rect 54 384 55 385
rect 53 384 54 385
rect 52 384 53 385
rect 51 384 52 385
rect 50 384 51 385
rect 27 384 28 385
rect 26 384 27 385
rect 25 384 26 385
rect 24 384 25 385
rect 23 384 24 385
rect 22 384 23 385
rect 21 384 22 385
rect 20 384 21 385
rect 19 384 20 385
rect 18 384 19 385
rect 17 384 18 385
rect 16 384 17 385
rect 15 384 16 385
rect 14 384 15 385
rect 13 384 14 385
rect 12 384 13 385
rect 194 385 195 386
rect 193 385 194 386
rect 192 385 193 386
rect 191 385 192 386
rect 190 385 191 386
rect 189 385 190 386
rect 170 385 171 386
rect 169 385 170 386
rect 168 385 169 386
rect 167 385 168 386
rect 166 385 167 386
rect 165 385 166 386
rect 164 385 165 386
rect 163 385 164 386
rect 162 385 163 386
rect 161 385 162 386
rect 127 385 128 386
rect 126 385 127 386
rect 125 385 126 386
rect 110 385 111 386
rect 109 385 110 386
rect 108 385 109 386
rect 107 385 108 386
rect 106 385 107 386
rect 105 385 106 386
rect 104 385 105 386
rect 103 385 104 386
rect 102 385 103 386
rect 101 385 102 386
rect 100 385 101 386
rect 75 385 76 386
rect 74 385 75 386
rect 73 385 74 386
rect 72 385 73 386
rect 71 385 72 386
rect 70 385 71 386
rect 69 385 70 386
rect 68 385 69 386
rect 67 385 68 386
rect 66 385 67 386
rect 65 385 66 386
rect 64 385 65 386
rect 63 385 64 386
rect 60 385 61 386
rect 59 385 60 386
rect 58 385 59 386
rect 57 385 58 386
rect 56 385 57 386
rect 55 385 56 386
rect 54 385 55 386
rect 53 385 54 386
rect 52 385 53 386
rect 51 385 52 386
rect 27 385 28 386
rect 26 385 27 386
rect 25 385 26 386
rect 24 385 25 386
rect 23 385 24 386
rect 22 385 23 386
rect 21 385 22 386
rect 20 385 21 386
rect 19 385 20 386
rect 18 385 19 386
rect 17 385 18 386
rect 16 385 17 386
rect 15 385 16 386
rect 14 385 15 386
rect 13 385 14 386
rect 12 385 13 386
rect 195 386 196 387
rect 194 386 195 387
rect 192 386 193 387
rect 190 386 191 387
rect 189 386 190 387
rect 181 386 182 387
rect 180 386 181 387
rect 179 386 180 387
rect 178 386 179 387
rect 177 386 178 387
rect 176 386 177 387
rect 175 386 176 387
rect 174 386 175 387
rect 171 386 172 387
rect 170 386 171 387
rect 169 386 170 387
rect 168 386 169 387
rect 167 386 168 387
rect 164 386 165 387
rect 163 386 164 387
rect 162 386 163 387
rect 161 386 162 387
rect 128 386 129 387
rect 127 386 128 387
rect 126 386 127 387
rect 125 386 126 387
rect 110 386 111 387
rect 109 386 110 387
rect 108 386 109 387
rect 107 386 108 387
rect 106 386 107 387
rect 105 386 106 387
rect 104 386 105 387
rect 103 386 104 387
rect 102 386 103 387
rect 101 386 102 387
rect 100 386 101 387
rect 74 386 75 387
rect 73 386 74 387
rect 72 386 73 387
rect 71 386 72 387
rect 70 386 71 387
rect 69 386 70 387
rect 68 386 69 387
rect 67 386 68 387
rect 66 386 67 387
rect 65 386 66 387
rect 64 386 65 387
rect 63 386 64 387
rect 59 386 60 387
rect 58 386 59 387
rect 57 386 58 387
rect 56 386 57 387
rect 55 386 56 387
rect 54 386 55 387
rect 53 386 54 387
rect 52 386 53 387
rect 27 386 28 387
rect 26 386 27 387
rect 25 386 26 387
rect 24 386 25 387
rect 23 386 24 387
rect 22 386 23 387
rect 21 386 22 387
rect 20 386 21 387
rect 19 386 20 387
rect 18 386 19 387
rect 17 386 18 387
rect 16 386 17 387
rect 15 386 16 387
rect 14 386 15 387
rect 13 386 14 387
rect 195 387 196 388
rect 194 387 195 388
rect 192 387 193 388
rect 190 387 191 388
rect 189 387 190 388
rect 181 387 182 388
rect 180 387 181 388
rect 179 387 180 388
rect 178 387 179 388
rect 177 387 178 388
rect 176 387 177 388
rect 175 387 176 388
rect 174 387 175 388
rect 171 387 172 388
rect 170 387 171 388
rect 169 387 170 388
rect 168 387 169 388
rect 163 387 164 388
rect 162 387 163 388
rect 161 387 162 388
rect 129 387 130 388
rect 128 387 129 388
rect 127 387 128 388
rect 126 387 127 388
rect 125 387 126 388
rect 110 387 111 388
rect 109 387 110 388
rect 108 387 109 388
rect 107 387 108 388
rect 106 387 107 388
rect 105 387 106 388
rect 104 387 105 388
rect 103 387 104 388
rect 102 387 103 388
rect 101 387 102 388
rect 100 387 101 388
rect 73 387 74 388
rect 72 387 73 388
rect 71 387 72 388
rect 70 387 71 388
rect 69 387 70 388
rect 68 387 69 388
rect 67 387 68 388
rect 66 387 67 388
rect 65 387 66 388
rect 64 387 65 388
rect 58 387 59 388
rect 57 387 58 388
rect 56 387 57 388
rect 55 387 56 388
rect 54 387 55 388
rect 27 387 28 388
rect 26 387 27 388
rect 25 387 26 388
rect 24 387 25 388
rect 23 387 24 388
rect 22 387 23 388
rect 195 388 196 389
rect 194 388 195 389
rect 192 388 193 389
rect 191 388 192 389
rect 190 388 191 389
rect 189 388 190 389
rect 181 388 182 389
rect 180 388 181 389
rect 179 388 180 389
rect 178 388 179 389
rect 177 388 178 389
rect 176 388 177 389
rect 175 388 176 389
rect 174 388 175 389
rect 171 388 172 389
rect 170 388 171 389
rect 169 388 170 389
rect 163 388 164 389
rect 162 388 163 389
rect 161 388 162 389
rect 160 388 161 389
rect 129 388 130 389
rect 128 388 129 389
rect 127 388 128 389
rect 126 388 127 389
rect 125 388 126 389
rect 110 388 111 389
rect 109 388 110 389
rect 108 388 109 389
rect 107 388 108 389
rect 106 388 107 389
rect 105 388 106 389
rect 104 388 105 389
rect 103 388 104 389
rect 102 388 103 389
rect 101 388 102 389
rect 100 388 101 389
rect 71 388 72 389
rect 70 388 71 389
rect 69 388 70 389
rect 68 388 69 389
rect 67 388 68 389
rect 66 388 67 389
rect 25 388 26 389
rect 24 388 25 389
rect 23 388 24 389
rect 22 388 23 389
rect 21 388 22 389
rect 20 388 21 389
rect 194 389 195 390
rect 192 389 193 390
rect 191 389 192 390
rect 190 389 191 390
rect 181 389 182 390
rect 180 389 181 390
rect 179 389 180 390
rect 178 389 179 390
rect 177 389 178 390
rect 176 389 177 390
rect 175 389 176 390
rect 174 389 175 390
rect 171 389 172 390
rect 170 389 171 390
rect 169 389 170 390
rect 162 389 163 390
rect 161 389 162 390
rect 160 389 161 390
rect 130 389 131 390
rect 129 389 130 390
rect 128 389 129 390
rect 127 389 128 390
rect 126 389 127 390
rect 125 389 126 390
rect 110 389 111 390
rect 109 389 110 390
rect 108 389 109 390
rect 107 389 108 390
rect 106 389 107 390
rect 105 389 106 390
rect 104 389 105 390
rect 103 389 104 390
rect 102 389 103 390
rect 101 389 102 390
rect 100 389 101 390
rect 23 389 24 390
rect 22 389 23 390
rect 21 389 22 390
rect 20 389 21 390
rect 19 389 20 390
rect 18 389 19 390
rect 194 390 195 391
rect 191 390 192 391
rect 181 390 182 391
rect 180 390 181 391
rect 179 390 180 391
rect 178 390 179 391
rect 171 390 172 391
rect 170 390 171 391
rect 169 390 170 391
rect 163 390 164 391
rect 162 390 163 391
rect 161 390 162 391
rect 160 390 161 391
rect 131 390 132 391
rect 130 390 131 391
rect 129 390 130 391
rect 128 390 129 391
rect 127 390 128 391
rect 126 390 127 391
rect 125 390 126 391
rect 110 390 111 391
rect 109 390 110 391
rect 108 390 109 391
rect 107 390 108 391
rect 106 390 107 391
rect 105 390 106 391
rect 104 390 105 391
rect 103 390 104 391
rect 102 390 103 391
rect 101 390 102 391
rect 100 390 101 391
rect 21 390 22 391
rect 20 390 21 391
rect 19 390 20 391
rect 18 390 19 391
rect 17 390 18 391
rect 16 390 17 391
rect 15 390 16 391
rect 195 391 196 392
rect 194 391 195 392
rect 192 391 193 392
rect 191 391 192 392
rect 190 391 191 392
rect 189 391 190 392
rect 181 391 182 392
rect 180 391 181 392
rect 179 391 180 392
rect 178 391 179 392
rect 171 391 172 392
rect 170 391 171 392
rect 169 391 170 392
rect 168 391 169 392
rect 163 391 164 392
rect 162 391 163 392
rect 161 391 162 392
rect 132 391 133 392
rect 131 391 132 392
rect 130 391 131 392
rect 129 391 130 392
rect 128 391 129 392
rect 127 391 128 392
rect 126 391 127 392
rect 125 391 126 392
rect 110 391 111 392
rect 109 391 110 392
rect 108 391 109 392
rect 107 391 108 392
rect 106 391 107 392
rect 105 391 106 392
rect 104 391 105 392
rect 103 391 104 392
rect 102 391 103 392
rect 101 391 102 392
rect 100 391 101 392
rect 19 391 20 392
rect 18 391 19 392
rect 17 391 18 392
rect 16 391 17 392
rect 15 391 16 392
rect 14 391 15 392
rect 13 391 14 392
rect 195 392 196 393
rect 194 392 195 393
rect 192 392 193 393
rect 191 392 192 393
rect 190 392 191 393
rect 189 392 190 393
rect 181 392 182 393
rect 180 392 181 393
rect 179 392 180 393
rect 178 392 179 393
rect 171 392 172 393
rect 170 392 171 393
rect 169 392 170 393
rect 168 392 169 393
rect 167 392 168 393
rect 164 392 165 393
rect 163 392 164 393
rect 162 392 163 393
rect 161 392 162 393
rect 133 392 134 393
rect 132 392 133 393
rect 131 392 132 393
rect 130 392 131 393
rect 129 392 130 393
rect 128 392 129 393
rect 127 392 128 393
rect 126 392 127 393
rect 125 392 126 393
rect 110 392 111 393
rect 109 392 110 393
rect 108 392 109 393
rect 107 392 108 393
rect 106 392 107 393
rect 105 392 106 393
rect 104 392 105 393
rect 103 392 104 393
rect 102 392 103 393
rect 101 392 102 393
rect 100 392 101 393
rect 84 392 85 393
rect 83 392 84 393
rect 82 392 83 393
rect 51 392 52 393
rect 50 392 51 393
rect 49 392 50 393
rect 17 392 18 393
rect 16 392 17 393
rect 15 392 16 393
rect 14 392 15 393
rect 13 392 14 393
rect 12 392 13 393
rect 195 393 196 394
rect 194 393 195 394
rect 193 393 194 394
rect 192 393 193 394
rect 190 393 191 394
rect 189 393 190 394
rect 181 393 182 394
rect 180 393 181 394
rect 179 393 180 394
rect 178 393 179 394
rect 170 393 171 394
rect 169 393 170 394
rect 168 393 169 394
rect 167 393 168 394
rect 166 393 167 394
rect 165 393 166 394
rect 164 393 165 394
rect 163 393 164 394
rect 162 393 163 394
rect 161 393 162 394
rect 134 393 135 394
rect 133 393 134 394
rect 132 393 133 394
rect 131 393 132 394
rect 130 393 131 394
rect 129 393 130 394
rect 128 393 129 394
rect 127 393 128 394
rect 126 393 127 394
rect 125 393 126 394
rect 110 393 111 394
rect 109 393 110 394
rect 108 393 109 394
rect 107 393 108 394
rect 106 393 107 394
rect 105 393 106 394
rect 104 393 105 394
rect 103 393 104 394
rect 102 393 103 394
rect 101 393 102 394
rect 100 393 101 394
rect 84 393 85 394
rect 83 393 84 394
rect 82 393 83 394
rect 81 393 82 394
rect 80 393 81 394
rect 53 393 54 394
rect 52 393 53 394
rect 51 393 52 394
rect 50 393 51 394
rect 49 393 50 394
rect 15 393 16 394
rect 14 393 15 394
rect 13 393 14 394
rect 12 393 13 394
rect 194 394 195 395
rect 193 394 194 395
rect 192 394 193 395
rect 189 394 190 395
rect 181 394 182 395
rect 180 394 181 395
rect 179 394 180 395
rect 178 394 179 395
rect 170 394 171 395
rect 169 394 170 395
rect 168 394 169 395
rect 167 394 168 395
rect 166 394 167 395
rect 165 394 166 395
rect 164 394 165 395
rect 163 394 164 395
rect 162 394 163 395
rect 134 394 135 395
rect 133 394 134 395
rect 132 394 133 395
rect 131 394 132 395
rect 130 394 131 395
rect 129 394 130 395
rect 128 394 129 395
rect 127 394 128 395
rect 126 394 127 395
rect 125 394 126 395
rect 110 394 111 395
rect 109 394 110 395
rect 108 394 109 395
rect 107 394 108 395
rect 106 394 107 395
rect 105 394 106 395
rect 104 394 105 395
rect 103 394 104 395
rect 102 394 103 395
rect 101 394 102 395
rect 100 394 101 395
rect 84 394 85 395
rect 83 394 84 395
rect 82 394 83 395
rect 81 394 82 395
rect 80 394 81 395
rect 79 394 80 395
rect 78 394 79 395
rect 77 394 78 395
rect 56 394 57 395
rect 55 394 56 395
rect 54 394 55 395
rect 53 394 54 395
rect 52 394 53 395
rect 51 394 52 395
rect 50 394 51 395
rect 49 394 50 395
rect 13 394 14 395
rect 193 395 194 396
rect 192 395 193 396
rect 191 395 192 396
rect 181 395 182 396
rect 180 395 181 396
rect 179 395 180 396
rect 178 395 179 396
rect 169 395 170 396
rect 168 395 169 396
rect 167 395 168 396
rect 166 395 167 396
rect 165 395 166 396
rect 164 395 165 396
rect 163 395 164 396
rect 162 395 163 396
rect 135 395 136 396
rect 134 395 135 396
rect 133 395 134 396
rect 132 395 133 396
rect 131 395 132 396
rect 130 395 131 396
rect 129 395 130 396
rect 128 395 129 396
rect 127 395 128 396
rect 126 395 127 396
rect 125 395 126 396
rect 110 395 111 396
rect 109 395 110 396
rect 108 395 109 396
rect 107 395 108 396
rect 106 395 107 396
rect 105 395 106 396
rect 104 395 105 396
rect 103 395 104 396
rect 102 395 103 396
rect 101 395 102 396
rect 100 395 101 396
rect 83 395 84 396
rect 82 395 83 396
rect 81 395 82 396
rect 80 395 81 396
rect 79 395 80 396
rect 78 395 79 396
rect 77 395 78 396
rect 76 395 77 396
rect 75 395 76 396
rect 74 395 75 396
rect 73 395 74 396
rect 72 395 73 396
rect 61 395 62 396
rect 60 395 61 396
rect 59 395 60 396
rect 58 395 59 396
rect 57 395 58 396
rect 56 395 57 396
rect 55 395 56 396
rect 54 395 55 396
rect 53 395 54 396
rect 52 395 53 396
rect 51 395 52 396
rect 50 395 51 396
rect 194 396 195 397
rect 193 396 194 397
rect 192 396 193 397
rect 191 396 192 397
rect 190 396 191 397
rect 189 396 190 397
rect 181 396 182 397
rect 180 396 181 397
rect 179 396 180 397
rect 178 396 179 397
rect 169 396 170 397
rect 168 396 169 397
rect 167 396 168 397
rect 166 396 167 397
rect 165 396 166 397
rect 164 396 165 397
rect 163 396 164 397
rect 162 396 163 397
rect 136 396 137 397
rect 135 396 136 397
rect 134 396 135 397
rect 133 396 134 397
rect 132 396 133 397
rect 131 396 132 397
rect 130 396 131 397
rect 129 396 130 397
rect 128 396 129 397
rect 127 396 128 397
rect 126 396 127 397
rect 125 396 126 397
rect 110 396 111 397
rect 109 396 110 397
rect 108 396 109 397
rect 107 396 108 397
rect 106 396 107 397
rect 105 396 106 397
rect 104 396 105 397
rect 103 396 104 397
rect 102 396 103 397
rect 101 396 102 397
rect 100 396 101 397
rect 82 396 83 397
rect 81 396 82 397
rect 80 396 81 397
rect 79 396 80 397
rect 78 396 79 397
rect 77 396 78 397
rect 76 396 77 397
rect 75 396 76 397
rect 74 396 75 397
rect 73 396 74 397
rect 72 396 73 397
rect 71 396 72 397
rect 70 396 71 397
rect 69 396 70 397
rect 68 396 69 397
rect 67 396 68 397
rect 66 396 67 397
rect 65 396 66 397
rect 64 396 65 397
rect 63 396 64 397
rect 62 396 63 397
rect 61 396 62 397
rect 60 396 61 397
rect 59 396 60 397
rect 58 396 59 397
rect 57 396 58 397
rect 56 396 57 397
rect 55 396 56 397
rect 54 396 55 397
rect 53 396 54 397
rect 52 396 53 397
rect 51 396 52 397
rect 195 397 196 398
rect 194 397 195 398
rect 193 397 194 398
rect 192 397 193 398
rect 191 397 192 398
rect 190 397 191 398
rect 189 397 190 398
rect 181 397 182 398
rect 180 397 181 398
rect 179 397 180 398
rect 178 397 179 398
rect 169 397 170 398
rect 168 397 169 398
rect 167 397 168 398
rect 165 397 166 398
rect 164 397 165 398
rect 163 397 164 398
rect 162 397 163 398
rect 137 397 138 398
rect 136 397 137 398
rect 135 397 136 398
rect 134 397 135 398
rect 133 397 134 398
rect 132 397 133 398
rect 131 397 132 398
rect 130 397 131 398
rect 129 397 130 398
rect 128 397 129 398
rect 127 397 128 398
rect 126 397 127 398
rect 125 397 126 398
rect 110 397 111 398
rect 109 397 110 398
rect 108 397 109 398
rect 107 397 108 398
rect 106 397 107 398
rect 105 397 106 398
rect 104 397 105 398
rect 103 397 104 398
rect 102 397 103 398
rect 101 397 102 398
rect 100 397 101 398
rect 80 397 81 398
rect 79 397 80 398
rect 78 397 79 398
rect 77 397 78 398
rect 76 397 77 398
rect 75 397 76 398
rect 74 397 75 398
rect 73 397 74 398
rect 72 397 73 398
rect 71 397 72 398
rect 70 397 71 398
rect 69 397 70 398
rect 68 397 69 398
rect 67 397 68 398
rect 66 397 67 398
rect 65 397 66 398
rect 64 397 65 398
rect 63 397 64 398
rect 62 397 63 398
rect 61 397 62 398
rect 60 397 61 398
rect 59 397 60 398
rect 58 397 59 398
rect 57 397 58 398
rect 56 397 57 398
rect 55 397 56 398
rect 54 397 55 398
rect 53 397 54 398
rect 195 398 196 399
rect 194 398 195 399
rect 192 398 193 399
rect 190 398 191 399
rect 189 398 190 399
rect 181 398 182 399
rect 180 398 181 399
rect 179 398 180 399
rect 178 398 179 399
rect 169 398 170 399
rect 168 398 169 399
rect 167 398 168 399
rect 165 398 166 399
rect 164 398 165 399
rect 163 398 164 399
rect 162 398 163 399
rect 138 398 139 399
rect 137 398 138 399
rect 136 398 137 399
rect 135 398 136 399
rect 134 398 135 399
rect 133 398 134 399
rect 132 398 133 399
rect 131 398 132 399
rect 130 398 131 399
rect 129 398 130 399
rect 128 398 129 399
rect 127 398 128 399
rect 126 398 127 399
rect 125 398 126 399
rect 110 398 111 399
rect 109 398 110 399
rect 108 398 109 399
rect 107 398 108 399
rect 106 398 107 399
rect 105 398 106 399
rect 104 398 105 399
rect 103 398 104 399
rect 102 398 103 399
rect 101 398 102 399
rect 100 398 101 399
rect 78 398 79 399
rect 77 398 78 399
rect 76 398 77 399
rect 75 398 76 399
rect 74 398 75 399
rect 73 398 74 399
rect 72 398 73 399
rect 71 398 72 399
rect 70 398 71 399
rect 69 398 70 399
rect 68 398 69 399
rect 67 398 68 399
rect 66 398 67 399
rect 65 398 66 399
rect 64 398 65 399
rect 63 398 64 399
rect 62 398 63 399
rect 61 398 62 399
rect 60 398 61 399
rect 59 398 60 399
rect 58 398 59 399
rect 57 398 58 399
rect 56 398 57 399
rect 55 398 56 399
rect 195 399 196 400
rect 194 399 195 400
rect 192 399 193 400
rect 191 399 192 400
rect 190 399 191 400
rect 189 399 190 400
rect 181 399 182 400
rect 180 399 181 400
rect 179 399 180 400
rect 178 399 179 400
rect 169 399 170 400
rect 168 399 169 400
rect 167 399 168 400
rect 165 399 166 400
rect 164 399 165 400
rect 163 399 164 400
rect 162 399 163 400
rect 138 399 139 400
rect 137 399 138 400
rect 136 399 137 400
rect 135 399 136 400
rect 134 399 135 400
rect 133 399 134 400
rect 132 399 133 400
rect 131 399 132 400
rect 130 399 131 400
rect 129 399 130 400
rect 128 399 129 400
rect 127 399 128 400
rect 126 399 127 400
rect 125 399 126 400
rect 110 399 111 400
rect 109 399 110 400
rect 108 399 109 400
rect 107 399 108 400
rect 106 399 107 400
rect 105 399 106 400
rect 104 399 105 400
rect 103 399 104 400
rect 102 399 103 400
rect 101 399 102 400
rect 100 399 101 400
rect 76 399 77 400
rect 75 399 76 400
rect 74 399 75 400
rect 73 399 74 400
rect 72 399 73 400
rect 71 399 72 400
rect 70 399 71 400
rect 69 399 70 400
rect 68 399 69 400
rect 67 399 68 400
rect 66 399 67 400
rect 65 399 66 400
rect 64 399 65 400
rect 63 399 64 400
rect 62 399 63 400
rect 61 399 62 400
rect 60 399 61 400
rect 59 399 60 400
rect 58 399 59 400
rect 57 399 58 400
rect 194 400 195 401
rect 192 400 193 401
rect 191 400 192 401
rect 190 400 191 401
rect 189 400 190 401
rect 181 400 182 401
rect 180 400 181 401
rect 179 400 180 401
rect 178 400 179 401
rect 175 400 176 401
rect 174 400 175 401
rect 173 400 174 401
rect 172 400 173 401
rect 171 400 172 401
rect 170 400 171 401
rect 169 400 170 401
rect 168 400 169 401
rect 167 400 168 401
rect 166 400 167 401
rect 165 400 166 401
rect 164 400 165 401
rect 163 400 164 401
rect 162 400 163 401
rect 161 400 162 401
rect 160 400 161 401
rect 139 400 140 401
rect 138 400 139 401
rect 137 400 138 401
rect 136 400 137 401
rect 135 400 136 401
rect 134 400 135 401
rect 133 400 134 401
rect 132 400 133 401
rect 131 400 132 401
rect 130 400 131 401
rect 129 400 130 401
rect 128 400 129 401
rect 127 400 128 401
rect 126 400 127 401
rect 125 400 126 401
rect 110 400 111 401
rect 109 400 110 401
rect 108 400 109 401
rect 107 400 108 401
rect 106 400 107 401
rect 105 400 106 401
rect 104 400 105 401
rect 103 400 104 401
rect 102 400 103 401
rect 101 400 102 401
rect 100 400 101 401
rect 72 400 73 401
rect 71 400 72 401
rect 70 400 71 401
rect 69 400 70 401
rect 68 400 69 401
rect 67 400 68 401
rect 66 400 67 401
rect 65 400 66 401
rect 64 400 65 401
rect 63 400 64 401
rect 62 400 63 401
rect 61 400 62 401
rect 60 400 61 401
rect 192 401 193 402
rect 191 401 192 402
rect 181 401 182 402
rect 180 401 181 402
rect 179 401 180 402
rect 178 401 179 402
rect 175 401 176 402
rect 174 401 175 402
rect 173 401 174 402
rect 172 401 173 402
rect 171 401 172 402
rect 170 401 171 402
rect 169 401 170 402
rect 168 401 169 402
rect 167 401 168 402
rect 166 401 167 402
rect 165 401 166 402
rect 164 401 165 402
rect 163 401 164 402
rect 162 401 163 402
rect 161 401 162 402
rect 160 401 161 402
rect 140 401 141 402
rect 139 401 140 402
rect 138 401 139 402
rect 137 401 138 402
rect 136 401 137 402
rect 135 401 136 402
rect 134 401 135 402
rect 133 401 134 402
rect 132 401 133 402
rect 131 401 132 402
rect 130 401 131 402
rect 129 401 130 402
rect 128 401 129 402
rect 127 401 128 402
rect 126 401 127 402
rect 125 401 126 402
rect 110 401 111 402
rect 109 401 110 402
rect 108 401 109 402
rect 107 401 108 402
rect 106 401 107 402
rect 105 401 106 402
rect 104 401 105 402
rect 103 401 104 402
rect 102 401 103 402
rect 101 401 102 402
rect 100 401 101 402
rect 194 402 195 403
rect 193 402 194 403
rect 192 402 193 403
rect 181 402 182 403
rect 180 402 181 403
rect 179 402 180 403
rect 178 402 179 403
rect 175 402 176 403
rect 174 402 175 403
rect 173 402 174 403
rect 172 402 173 403
rect 171 402 172 403
rect 170 402 171 403
rect 169 402 170 403
rect 168 402 169 403
rect 167 402 168 403
rect 166 402 167 403
rect 165 402 166 403
rect 164 402 165 403
rect 163 402 164 403
rect 162 402 163 403
rect 161 402 162 403
rect 160 402 161 403
rect 141 402 142 403
rect 140 402 141 403
rect 139 402 140 403
rect 138 402 139 403
rect 137 402 138 403
rect 136 402 137 403
rect 135 402 136 403
rect 134 402 135 403
rect 133 402 134 403
rect 132 402 133 403
rect 131 402 132 403
rect 130 402 131 403
rect 129 402 130 403
rect 128 402 129 403
rect 127 402 128 403
rect 126 402 127 403
rect 125 402 126 403
rect 110 402 111 403
rect 109 402 110 403
rect 108 402 109 403
rect 107 402 108 403
rect 106 402 107 403
rect 105 402 106 403
rect 104 402 105 403
rect 103 402 104 403
rect 102 402 103 403
rect 101 402 102 403
rect 100 402 101 403
rect 195 403 196 404
rect 194 403 195 404
rect 193 403 194 404
rect 192 403 193 404
rect 190 403 191 404
rect 189 403 190 404
rect 181 403 182 404
rect 180 403 181 404
rect 179 403 180 404
rect 178 403 179 404
rect 175 403 176 404
rect 174 403 175 404
rect 173 403 174 404
rect 172 403 173 404
rect 171 403 172 404
rect 170 403 171 404
rect 169 403 170 404
rect 168 403 169 404
rect 167 403 168 404
rect 166 403 167 404
rect 165 403 166 404
rect 164 403 165 404
rect 163 403 164 404
rect 162 403 163 404
rect 161 403 162 404
rect 160 403 161 404
rect 142 403 143 404
rect 141 403 142 404
rect 140 403 141 404
rect 139 403 140 404
rect 138 403 139 404
rect 137 403 138 404
rect 136 403 137 404
rect 135 403 136 404
rect 134 403 135 404
rect 133 403 134 404
rect 132 403 133 404
rect 131 403 132 404
rect 130 403 131 404
rect 129 403 130 404
rect 128 403 129 404
rect 127 403 128 404
rect 126 403 127 404
rect 125 403 126 404
rect 110 403 111 404
rect 109 403 110 404
rect 108 403 109 404
rect 107 403 108 404
rect 106 403 107 404
rect 105 403 106 404
rect 104 403 105 404
rect 103 403 104 404
rect 102 403 103 404
rect 101 403 102 404
rect 100 403 101 404
rect 195 404 196 405
rect 194 404 195 405
rect 192 404 193 405
rect 191 404 192 405
rect 190 404 191 405
rect 189 404 190 405
rect 180 404 181 405
rect 179 404 180 405
rect 178 404 179 405
rect 174 404 175 405
rect 173 404 174 405
rect 172 404 173 405
rect 171 404 172 405
rect 170 404 171 405
rect 169 404 170 405
rect 168 404 169 405
rect 167 404 168 405
rect 166 404 167 405
rect 165 404 166 405
rect 164 404 165 405
rect 163 404 164 405
rect 162 404 163 405
rect 161 404 162 405
rect 142 404 143 405
rect 141 404 142 405
rect 140 404 141 405
rect 139 404 140 405
rect 138 404 139 405
rect 137 404 138 405
rect 136 404 137 405
rect 135 404 136 405
rect 134 404 135 405
rect 133 404 134 405
rect 132 404 133 405
rect 131 404 132 405
rect 130 404 131 405
rect 129 404 130 405
rect 128 404 129 405
rect 127 404 128 405
rect 126 404 127 405
rect 125 404 126 405
rect 110 404 111 405
rect 109 404 110 405
rect 108 404 109 405
rect 107 404 108 405
rect 106 404 107 405
rect 105 404 106 405
rect 104 404 105 405
rect 103 404 104 405
rect 102 404 103 405
rect 101 404 102 405
rect 100 404 101 405
rect 194 405 195 406
rect 192 405 193 406
rect 191 405 192 406
rect 190 405 191 406
rect 189 405 190 406
rect 143 405 144 406
rect 142 405 143 406
rect 141 405 142 406
rect 140 405 141 406
rect 139 405 140 406
rect 138 405 139 406
rect 137 405 138 406
rect 136 405 137 406
rect 135 405 136 406
rect 134 405 135 406
rect 133 405 134 406
rect 132 405 133 406
rect 131 405 132 406
rect 130 405 131 406
rect 129 405 130 406
rect 128 405 129 406
rect 127 405 128 406
rect 126 405 127 406
rect 125 405 126 406
rect 110 405 111 406
rect 109 405 110 406
rect 108 405 109 406
rect 107 405 108 406
rect 106 405 107 406
rect 105 405 106 406
rect 104 405 105 406
rect 103 405 104 406
rect 102 405 103 406
rect 101 405 102 406
rect 100 405 101 406
rect 195 406 196 407
rect 194 406 195 407
rect 193 406 194 407
rect 192 406 193 407
rect 191 406 192 407
rect 190 406 191 407
rect 189 406 190 407
rect 144 406 145 407
rect 143 406 144 407
rect 142 406 143 407
rect 141 406 142 407
rect 140 406 141 407
rect 139 406 140 407
rect 138 406 139 407
rect 137 406 138 407
rect 136 406 137 407
rect 135 406 136 407
rect 134 406 135 407
rect 133 406 134 407
rect 132 406 133 407
rect 131 406 132 407
rect 130 406 131 407
rect 129 406 130 407
rect 128 406 129 407
rect 127 406 128 407
rect 126 406 127 407
rect 125 406 126 407
rect 110 406 111 407
rect 109 406 110 407
rect 108 406 109 407
rect 107 406 108 407
rect 106 406 107 407
rect 105 406 106 407
rect 104 406 105 407
rect 103 406 104 407
rect 102 406 103 407
rect 101 406 102 407
rect 100 406 101 407
rect 194 407 195 408
rect 193 407 194 408
rect 192 407 193 408
rect 191 407 192 408
rect 190 407 191 408
rect 189 407 190 408
rect 145 407 146 408
rect 144 407 145 408
rect 143 407 144 408
rect 142 407 143 408
rect 141 407 142 408
rect 140 407 141 408
rect 139 407 140 408
rect 138 407 139 408
rect 137 407 138 408
rect 136 407 137 408
rect 135 407 136 408
rect 134 407 135 408
rect 133 407 134 408
rect 132 407 133 408
rect 131 407 132 408
rect 130 407 131 408
rect 129 407 130 408
rect 128 407 129 408
rect 127 407 128 408
rect 126 407 127 408
rect 125 407 126 408
rect 110 407 111 408
rect 109 407 110 408
rect 108 407 109 408
rect 107 407 108 408
rect 106 407 107 408
rect 105 407 106 408
rect 104 407 105 408
rect 103 407 104 408
rect 102 407 103 408
rect 101 407 102 408
rect 100 407 101 408
rect 146 408 147 409
rect 145 408 146 409
rect 144 408 145 409
rect 143 408 144 409
rect 142 408 143 409
rect 141 408 142 409
rect 140 408 141 409
rect 139 408 140 409
rect 138 408 139 409
rect 137 408 138 409
rect 136 408 137 409
rect 135 408 136 409
rect 134 408 135 409
rect 133 408 134 409
rect 132 408 133 409
rect 131 408 132 409
rect 130 408 131 409
rect 129 408 130 409
rect 128 408 129 409
rect 127 408 128 409
rect 126 408 127 409
rect 125 408 126 409
rect 110 408 111 409
rect 109 408 110 409
rect 108 408 109 409
rect 107 408 108 409
rect 106 408 107 409
rect 105 408 106 409
rect 104 408 105 409
rect 103 408 104 409
rect 102 408 103 409
rect 101 408 102 409
rect 100 408 101 409
rect 194 409 195 410
rect 193 409 194 410
rect 192 409 193 410
rect 191 409 192 410
rect 190 409 191 410
rect 189 409 190 410
rect 147 409 148 410
rect 146 409 147 410
rect 145 409 146 410
rect 144 409 145 410
rect 143 409 144 410
rect 142 409 143 410
rect 141 409 142 410
rect 140 409 141 410
rect 139 409 140 410
rect 138 409 139 410
rect 137 409 138 410
rect 136 409 137 410
rect 135 409 136 410
rect 134 409 135 410
rect 133 409 134 410
rect 132 409 133 410
rect 131 409 132 410
rect 130 409 131 410
rect 129 409 130 410
rect 128 409 129 410
rect 127 409 128 410
rect 126 409 127 410
rect 125 409 126 410
rect 110 409 111 410
rect 109 409 110 410
rect 108 409 109 410
rect 107 409 108 410
rect 106 409 107 410
rect 105 409 106 410
rect 104 409 105 410
rect 103 409 104 410
rect 102 409 103 410
rect 101 409 102 410
rect 100 409 101 410
rect 195 410 196 411
rect 194 410 195 411
rect 193 410 194 411
rect 192 410 193 411
rect 191 410 192 411
rect 190 410 191 411
rect 189 410 190 411
rect 147 410 148 411
rect 146 410 147 411
rect 145 410 146 411
rect 144 410 145 411
rect 143 410 144 411
rect 142 410 143 411
rect 141 410 142 411
rect 140 410 141 411
rect 139 410 140 411
rect 138 410 139 411
rect 137 410 138 411
rect 136 410 137 411
rect 135 410 136 411
rect 134 410 135 411
rect 133 410 134 411
rect 132 410 133 411
rect 131 410 132 411
rect 130 410 131 411
rect 129 410 130 411
rect 128 410 129 411
rect 127 410 128 411
rect 126 410 127 411
rect 125 410 126 411
rect 124 410 125 411
rect 123 410 124 411
rect 122 410 123 411
rect 121 410 122 411
rect 120 410 121 411
rect 119 410 120 411
rect 118 410 119 411
rect 117 410 118 411
rect 116 410 117 411
rect 115 410 116 411
rect 114 410 115 411
rect 113 410 114 411
rect 112 410 113 411
rect 111 410 112 411
rect 110 410 111 411
rect 109 410 110 411
rect 108 410 109 411
rect 107 410 108 411
rect 106 410 107 411
rect 105 410 106 411
rect 104 410 105 411
rect 103 410 104 411
rect 102 410 103 411
rect 101 410 102 411
rect 100 410 101 411
rect 190 411 191 412
rect 189 411 190 412
rect 148 411 149 412
rect 147 411 148 412
rect 146 411 147 412
rect 145 411 146 412
rect 144 411 145 412
rect 143 411 144 412
rect 142 411 143 412
rect 141 411 142 412
rect 140 411 141 412
rect 139 411 140 412
rect 138 411 139 412
rect 137 411 138 412
rect 136 411 137 412
rect 135 411 136 412
rect 134 411 135 412
rect 133 411 134 412
rect 132 411 133 412
rect 131 411 132 412
rect 130 411 131 412
rect 129 411 130 412
rect 128 411 129 412
rect 127 411 128 412
rect 126 411 127 412
rect 125 411 126 412
rect 124 411 125 412
rect 123 411 124 412
rect 122 411 123 412
rect 121 411 122 412
rect 120 411 121 412
rect 119 411 120 412
rect 118 411 119 412
rect 117 411 118 412
rect 116 411 117 412
rect 115 411 116 412
rect 114 411 115 412
rect 113 411 114 412
rect 112 411 113 412
rect 111 411 112 412
rect 110 411 111 412
rect 109 411 110 412
rect 108 411 109 412
rect 107 411 108 412
rect 106 411 107 412
rect 105 411 106 412
rect 104 411 105 412
rect 103 411 104 412
rect 102 411 103 412
rect 101 411 102 412
rect 100 411 101 412
rect 190 412 191 413
rect 189 412 190 413
rect 149 412 150 413
rect 148 412 149 413
rect 147 412 148 413
rect 146 412 147 413
rect 145 412 146 413
rect 144 412 145 413
rect 143 412 144 413
rect 142 412 143 413
rect 141 412 142 413
rect 140 412 141 413
rect 139 412 140 413
rect 138 412 139 413
rect 137 412 138 413
rect 136 412 137 413
rect 135 412 136 413
rect 134 412 135 413
rect 133 412 134 413
rect 132 412 133 413
rect 131 412 132 413
rect 130 412 131 413
rect 129 412 130 413
rect 128 412 129 413
rect 127 412 128 413
rect 125 412 126 413
rect 124 412 125 413
rect 123 412 124 413
rect 122 412 123 413
rect 121 412 122 413
rect 120 412 121 413
rect 119 412 120 413
rect 118 412 119 413
rect 117 412 118 413
rect 116 412 117 413
rect 115 412 116 413
rect 114 412 115 413
rect 113 412 114 413
rect 112 412 113 413
rect 111 412 112 413
rect 110 412 111 413
rect 109 412 110 413
rect 108 412 109 413
rect 107 412 108 413
rect 106 412 107 413
rect 105 412 106 413
rect 104 412 105 413
rect 103 412 104 413
rect 102 412 103 413
rect 101 412 102 413
rect 100 412 101 413
rect 194 413 195 414
rect 193 413 194 414
rect 192 413 193 414
rect 191 413 192 414
rect 190 413 191 414
rect 150 413 151 414
rect 149 413 150 414
rect 148 413 149 414
rect 147 413 148 414
rect 146 413 147 414
rect 145 413 146 414
rect 144 413 145 414
rect 143 413 144 414
rect 142 413 143 414
rect 141 413 142 414
rect 140 413 141 414
rect 139 413 140 414
rect 138 413 139 414
rect 137 413 138 414
rect 136 413 137 414
rect 135 413 136 414
rect 134 413 135 414
rect 133 413 134 414
rect 132 413 133 414
rect 131 413 132 414
rect 130 413 131 414
rect 129 413 130 414
rect 128 413 129 414
rect 125 413 126 414
rect 124 413 125 414
rect 123 413 124 414
rect 122 413 123 414
rect 121 413 122 414
rect 120 413 121 414
rect 119 413 120 414
rect 118 413 119 414
rect 117 413 118 414
rect 116 413 117 414
rect 115 413 116 414
rect 114 413 115 414
rect 113 413 114 414
rect 112 413 113 414
rect 111 413 112 414
rect 110 413 111 414
rect 109 413 110 414
rect 108 413 109 414
rect 107 413 108 414
rect 106 413 107 414
rect 105 413 106 414
rect 104 413 105 414
rect 103 413 104 414
rect 102 413 103 414
rect 101 413 102 414
rect 100 413 101 414
rect 194 414 195 415
rect 193 414 194 415
rect 192 414 193 415
rect 191 414 192 415
rect 190 414 191 415
rect 189 414 190 415
rect 151 414 152 415
rect 150 414 151 415
rect 149 414 150 415
rect 148 414 149 415
rect 147 414 148 415
rect 146 414 147 415
rect 145 414 146 415
rect 144 414 145 415
rect 143 414 144 415
rect 142 414 143 415
rect 141 414 142 415
rect 140 414 141 415
rect 139 414 140 415
rect 138 414 139 415
rect 137 414 138 415
rect 136 414 137 415
rect 135 414 136 415
rect 134 414 135 415
rect 133 414 134 415
rect 132 414 133 415
rect 131 414 132 415
rect 130 414 131 415
rect 129 414 130 415
rect 125 414 126 415
rect 124 414 125 415
rect 123 414 124 415
rect 122 414 123 415
rect 121 414 122 415
rect 120 414 121 415
rect 119 414 120 415
rect 118 414 119 415
rect 117 414 118 415
rect 116 414 117 415
rect 115 414 116 415
rect 114 414 115 415
rect 113 414 114 415
rect 112 414 113 415
rect 111 414 112 415
rect 110 414 111 415
rect 109 414 110 415
rect 108 414 109 415
rect 107 414 108 415
rect 106 414 107 415
rect 105 414 106 415
rect 104 414 105 415
rect 103 414 104 415
rect 102 414 103 415
rect 101 414 102 415
rect 100 414 101 415
rect 194 415 195 416
rect 193 415 194 416
rect 190 415 191 416
rect 189 415 190 416
rect 151 415 152 416
rect 150 415 151 416
rect 149 415 150 416
rect 148 415 149 416
rect 147 415 148 416
rect 146 415 147 416
rect 145 415 146 416
rect 144 415 145 416
rect 143 415 144 416
rect 142 415 143 416
rect 141 415 142 416
rect 140 415 141 416
rect 139 415 140 416
rect 138 415 139 416
rect 137 415 138 416
rect 136 415 137 416
rect 135 415 136 416
rect 134 415 135 416
rect 133 415 134 416
rect 132 415 133 416
rect 131 415 132 416
rect 130 415 131 416
rect 129 415 130 416
rect 125 415 126 416
rect 124 415 125 416
rect 123 415 124 416
rect 122 415 123 416
rect 121 415 122 416
rect 120 415 121 416
rect 119 415 120 416
rect 118 415 119 416
rect 117 415 118 416
rect 116 415 117 416
rect 115 415 116 416
rect 114 415 115 416
rect 113 415 114 416
rect 112 415 113 416
rect 111 415 112 416
rect 110 415 111 416
rect 109 415 110 416
rect 108 415 109 416
rect 107 415 108 416
rect 106 415 107 416
rect 105 415 106 416
rect 104 415 105 416
rect 103 415 104 416
rect 102 415 103 416
rect 101 415 102 416
rect 100 415 101 416
rect 195 416 196 417
rect 194 416 195 417
rect 190 416 191 417
rect 189 416 190 417
rect 172 416 173 417
rect 171 416 172 417
rect 170 416 171 417
rect 151 416 152 417
rect 150 416 151 417
rect 149 416 150 417
rect 148 416 149 417
rect 147 416 148 417
rect 146 416 147 417
rect 145 416 146 417
rect 144 416 145 417
rect 143 416 144 417
rect 142 416 143 417
rect 141 416 142 417
rect 140 416 141 417
rect 139 416 140 417
rect 138 416 139 417
rect 137 416 138 417
rect 136 416 137 417
rect 135 416 136 417
rect 134 416 135 417
rect 133 416 134 417
rect 132 416 133 417
rect 131 416 132 417
rect 130 416 131 417
rect 125 416 126 417
rect 124 416 125 417
rect 123 416 124 417
rect 122 416 123 417
rect 121 416 122 417
rect 120 416 121 417
rect 119 416 120 417
rect 118 416 119 417
rect 117 416 118 417
rect 116 416 117 417
rect 115 416 116 417
rect 114 416 115 417
rect 113 416 114 417
rect 112 416 113 417
rect 111 416 112 417
rect 110 416 111 417
rect 109 416 110 417
rect 108 416 109 417
rect 107 416 108 417
rect 106 416 107 417
rect 105 416 106 417
rect 104 416 105 417
rect 103 416 104 417
rect 102 416 103 417
rect 101 416 102 417
rect 100 416 101 417
rect 194 417 195 418
rect 189 417 190 418
rect 172 417 173 418
rect 171 417 172 418
rect 170 417 171 418
rect 151 417 152 418
rect 150 417 151 418
rect 149 417 150 418
rect 148 417 149 418
rect 147 417 148 418
rect 146 417 147 418
rect 145 417 146 418
rect 144 417 145 418
rect 143 417 144 418
rect 142 417 143 418
rect 141 417 142 418
rect 140 417 141 418
rect 139 417 140 418
rect 138 417 139 418
rect 137 417 138 418
rect 136 417 137 418
rect 135 417 136 418
rect 134 417 135 418
rect 133 417 134 418
rect 132 417 133 418
rect 131 417 132 418
rect 125 417 126 418
rect 124 417 125 418
rect 123 417 124 418
rect 122 417 123 418
rect 121 417 122 418
rect 120 417 121 418
rect 119 417 120 418
rect 118 417 119 418
rect 117 417 118 418
rect 116 417 117 418
rect 115 417 116 418
rect 114 417 115 418
rect 113 417 114 418
rect 112 417 113 418
rect 111 417 112 418
rect 110 417 111 418
rect 109 417 110 418
rect 108 417 109 418
rect 107 417 108 418
rect 106 417 107 418
rect 105 417 106 418
rect 104 417 105 418
rect 103 417 104 418
rect 102 417 103 418
rect 101 417 102 418
rect 100 417 101 418
rect 172 418 173 419
rect 171 418 172 419
rect 170 418 171 419
rect 162 418 163 419
rect 151 418 152 419
rect 150 418 151 419
rect 149 418 150 419
rect 148 418 149 419
rect 147 418 148 419
rect 146 418 147 419
rect 145 418 146 419
rect 144 418 145 419
rect 143 418 144 419
rect 142 418 143 419
rect 141 418 142 419
rect 140 418 141 419
rect 139 418 140 419
rect 138 418 139 419
rect 137 418 138 419
rect 136 418 137 419
rect 135 418 136 419
rect 134 418 135 419
rect 133 418 134 419
rect 132 418 133 419
rect 125 418 126 419
rect 124 418 125 419
rect 123 418 124 419
rect 122 418 123 419
rect 121 418 122 419
rect 120 418 121 419
rect 119 418 120 419
rect 118 418 119 419
rect 117 418 118 419
rect 116 418 117 419
rect 115 418 116 419
rect 114 418 115 419
rect 113 418 114 419
rect 112 418 113 419
rect 111 418 112 419
rect 110 418 111 419
rect 109 418 110 419
rect 108 418 109 419
rect 107 418 108 419
rect 106 418 107 419
rect 105 418 106 419
rect 104 418 105 419
rect 103 418 104 419
rect 102 418 103 419
rect 101 418 102 419
rect 100 418 101 419
rect 195 419 196 420
rect 194 419 195 420
rect 193 419 194 420
rect 192 419 193 420
rect 191 419 192 420
rect 190 419 191 420
rect 189 419 190 420
rect 188 419 189 420
rect 187 419 188 420
rect 186 419 187 420
rect 172 419 173 420
rect 171 419 172 420
rect 170 419 171 420
rect 163 419 164 420
rect 162 419 163 420
rect 161 419 162 420
rect 151 419 152 420
rect 150 419 151 420
rect 149 419 150 420
rect 148 419 149 420
rect 147 419 148 420
rect 146 419 147 420
rect 145 419 146 420
rect 144 419 145 420
rect 143 419 144 420
rect 142 419 143 420
rect 141 419 142 420
rect 140 419 141 420
rect 139 419 140 420
rect 138 419 139 420
rect 137 419 138 420
rect 136 419 137 420
rect 135 419 136 420
rect 134 419 135 420
rect 133 419 134 420
rect 125 419 126 420
rect 124 419 125 420
rect 123 419 124 420
rect 122 419 123 420
rect 121 419 122 420
rect 120 419 121 420
rect 119 419 120 420
rect 118 419 119 420
rect 117 419 118 420
rect 116 419 117 420
rect 115 419 116 420
rect 114 419 115 420
rect 113 419 114 420
rect 112 419 113 420
rect 111 419 112 420
rect 110 419 111 420
rect 109 419 110 420
rect 108 419 109 420
rect 107 419 108 420
rect 106 419 107 420
rect 105 419 106 420
rect 104 419 105 420
rect 103 419 104 420
rect 102 419 103 420
rect 101 419 102 420
rect 100 419 101 420
rect 194 420 195 421
rect 193 420 194 421
rect 192 420 193 421
rect 191 420 192 421
rect 190 420 191 421
rect 189 420 190 421
rect 188 420 189 421
rect 187 420 188 421
rect 186 420 187 421
rect 172 420 173 421
rect 171 420 172 421
rect 170 420 171 421
rect 163 420 164 421
rect 162 420 163 421
rect 161 420 162 421
rect 151 420 152 421
rect 150 420 151 421
rect 149 420 150 421
rect 148 420 149 421
rect 147 420 148 421
rect 146 420 147 421
rect 145 420 146 421
rect 144 420 145 421
rect 143 420 144 421
rect 142 420 143 421
rect 141 420 142 421
rect 140 420 141 421
rect 139 420 140 421
rect 138 420 139 421
rect 137 420 138 421
rect 136 420 137 421
rect 135 420 136 421
rect 134 420 135 421
rect 125 420 126 421
rect 124 420 125 421
rect 123 420 124 421
rect 122 420 123 421
rect 121 420 122 421
rect 120 420 121 421
rect 119 420 120 421
rect 118 420 119 421
rect 117 420 118 421
rect 116 420 117 421
rect 115 420 116 421
rect 114 420 115 421
rect 113 420 114 421
rect 112 420 113 421
rect 111 420 112 421
rect 110 420 111 421
rect 109 420 110 421
rect 108 420 109 421
rect 107 420 108 421
rect 106 420 107 421
rect 105 420 106 421
rect 104 420 105 421
rect 103 420 104 421
rect 102 420 103 421
rect 101 420 102 421
rect 100 420 101 421
rect 190 421 191 422
rect 189 421 190 422
rect 172 421 173 422
rect 171 421 172 422
rect 170 421 171 422
rect 163 421 164 422
rect 162 421 163 422
rect 161 421 162 422
rect 151 421 152 422
rect 150 421 151 422
rect 149 421 150 422
rect 148 421 149 422
rect 147 421 148 422
rect 146 421 147 422
rect 145 421 146 422
rect 144 421 145 422
rect 143 421 144 422
rect 142 421 143 422
rect 141 421 142 422
rect 140 421 141 422
rect 139 421 140 422
rect 138 421 139 422
rect 137 421 138 422
rect 136 421 137 422
rect 135 421 136 422
rect 134 421 135 422
rect 125 421 126 422
rect 124 421 125 422
rect 123 421 124 422
rect 122 421 123 422
rect 121 421 122 422
rect 120 421 121 422
rect 119 421 120 422
rect 118 421 119 422
rect 117 421 118 422
rect 116 421 117 422
rect 115 421 116 422
rect 114 421 115 422
rect 113 421 114 422
rect 112 421 113 422
rect 111 421 112 422
rect 110 421 111 422
rect 109 421 110 422
rect 108 421 109 422
rect 107 421 108 422
rect 106 421 107 422
rect 105 421 106 422
rect 104 421 105 422
rect 103 421 104 422
rect 102 421 103 422
rect 101 421 102 422
rect 100 421 101 422
rect 194 422 195 423
rect 193 422 194 423
rect 192 422 193 423
rect 190 422 191 423
rect 189 422 190 423
rect 172 422 173 423
rect 171 422 172 423
rect 170 422 171 423
rect 163 422 164 423
rect 162 422 163 423
rect 161 422 162 423
rect 151 422 152 423
rect 150 422 151 423
rect 149 422 150 423
rect 148 422 149 423
rect 147 422 148 423
rect 146 422 147 423
rect 145 422 146 423
rect 144 422 145 423
rect 143 422 144 423
rect 142 422 143 423
rect 141 422 142 423
rect 140 422 141 423
rect 139 422 140 423
rect 138 422 139 423
rect 137 422 138 423
rect 136 422 137 423
rect 135 422 136 423
rect 125 422 126 423
rect 124 422 125 423
rect 123 422 124 423
rect 122 422 123 423
rect 121 422 122 423
rect 120 422 121 423
rect 119 422 120 423
rect 118 422 119 423
rect 117 422 118 423
rect 116 422 117 423
rect 115 422 116 423
rect 114 422 115 423
rect 113 422 114 423
rect 112 422 113 423
rect 111 422 112 423
rect 110 422 111 423
rect 109 422 110 423
rect 108 422 109 423
rect 107 422 108 423
rect 106 422 107 423
rect 105 422 106 423
rect 104 422 105 423
rect 103 422 104 423
rect 102 422 103 423
rect 101 422 102 423
rect 100 422 101 423
rect 195 423 196 424
rect 194 423 195 424
rect 193 423 194 424
rect 192 423 193 424
rect 191 423 192 424
rect 190 423 191 424
rect 189 423 190 424
rect 172 423 173 424
rect 171 423 172 424
rect 170 423 171 424
rect 163 423 164 424
rect 162 423 163 424
rect 161 423 162 424
rect 151 423 152 424
rect 150 423 151 424
rect 149 423 150 424
rect 148 423 149 424
rect 147 423 148 424
rect 146 423 147 424
rect 145 423 146 424
rect 144 423 145 424
rect 143 423 144 424
rect 142 423 143 424
rect 141 423 142 424
rect 140 423 141 424
rect 139 423 140 424
rect 138 423 139 424
rect 137 423 138 424
rect 136 423 137 424
rect 125 423 126 424
rect 124 423 125 424
rect 123 423 124 424
rect 122 423 123 424
rect 121 423 122 424
rect 120 423 121 424
rect 119 423 120 424
rect 118 423 119 424
rect 117 423 118 424
rect 116 423 117 424
rect 115 423 116 424
rect 114 423 115 424
rect 113 423 114 424
rect 112 423 113 424
rect 111 423 112 424
rect 110 423 111 424
rect 109 423 110 424
rect 108 423 109 424
rect 107 423 108 424
rect 106 423 107 424
rect 105 423 106 424
rect 104 423 105 424
rect 103 423 104 424
rect 102 423 103 424
rect 101 423 102 424
rect 100 423 101 424
rect 172 424 173 425
rect 171 424 172 425
rect 170 424 171 425
rect 163 424 164 425
rect 162 424 163 425
rect 161 424 162 425
rect 151 424 152 425
rect 150 424 151 425
rect 149 424 150 425
rect 148 424 149 425
rect 147 424 148 425
rect 146 424 147 425
rect 145 424 146 425
rect 144 424 145 425
rect 143 424 144 425
rect 142 424 143 425
rect 141 424 142 425
rect 140 424 141 425
rect 139 424 140 425
rect 138 424 139 425
rect 137 424 138 425
rect 125 424 126 425
rect 124 424 125 425
rect 123 424 124 425
rect 122 424 123 425
rect 121 424 122 425
rect 120 424 121 425
rect 119 424 120 425
rect 118 424 119 425
rect 117 424 118 425
rect 116 424 117 425
rect 115 424 116 425
rect 114 424 115 425
rect 113 424 114 425
rect 112 424 113 425
rect 111 424 112 425
rect 110 424 111 425
rect 109 424 110 425
rect 108 424 109 425
rect 107 424 108 425
rect 106 424 107 425
rect 105 424 106 425
rect 104 424 105 425
rect 103 424 104 425
rect 102 424 103 425
rect 101 424 102 425
rect 100 424 101 425
rect 172 425 173 426
rect 171 425 172 426
rect 170 425 171 426
rect 163 425 164 426
rect 162 425 163 426
rect 161 425 162 426
rect 151 425 152 426
rect 150 425 151 426
rect 149 425 150 426
rect 148 425 149 426
rect 147 425 148 426
rect 146 425 147 426
rect 145 425 146 426
rect 144 425 145 426
rect 143 425 144 426
rect 142 425 143 426
rect 141 425 142 426
rect 140 425 141 426
rect 139 425 140 426
rect 138 425 139 426
rect 125 425 126 426
rect 124 425 125 426
rect 123 425 124 426
rect 122 425 123 426
rect 121 425 122 426
rect 120 425 121 426
rect 119 425 120 426
rect 118 425 119 426
rect 117 425 118 426
rect 116 425 117 426
rect 115 425 116 426
rect 114 425 115 426
rect 113 425 114 426
rect 112 425 113 426
rect 111 425 112 426
rect 110 425 111 426
rect 109 425 110 426
rect 108 425 109 426
rect 107 425 108 426
rect 106 425 107 426
rect 105 425 106 426
rect 104 425 105 426
rect 103 425 104 426
rect 102 425 103 426
rect 101 425 102 426
rect 100 425 101 426
rect 181 426 182 427
rect 180 426 181 427
rect 179 426 180 427
rect 178 426 179 427
rect 177 426 178 427
rect 176 426 177 427
rect 175 426 176 427
rect 174 426 175 427
rect 173 426 174 427
rect 172 426 173 427
rect 171 426 172 427
rect 170 426 171 427
rect 163 426 164 427
rect 162 426 163 427
rect 161 426 162 427
rect 151 426 152 427
rect 150 426 151 427
rect 149 426 150 427
rect 148 426 149 427
rect 147 426 148 427
rect 146 426 147 427
rect 145 426 146 427
rect 144 426 145 427
rect 143 426 144 427
rect 142 426 143 427
rect 141 426 142 427
rect 140 426 141 427
rect 139 426 140 427
rect 138 426 139 427
rect 125 426 126 427
rect 124 426 125 427
rect 123 426 124 427
rect 122 426 123 427
rect 121 426 122 427
rect 120 426 121 427
rect 119 426 120 427
rect 118 426 119 427
rect 117 426 118 427
rect 116 426 117 427
rect 115 426 116 427
rect 114 426 115 427
rect 113 426 114 427
rect 112 426 113 427
rect 111 426 112 427
rect 110 426 111 427
rect 109 426 110 427
rect 108 426 109 427
rect 107 426 108 427
rect 106 426 107 427
rect 105 426 106 427
rect 104 426 105 427
rect 103 426 104 427
rect 102 426 103 427
rect 101 426 102 427
rect 181 427 182 428
rect 180 427 181 428
rect 179 427 180 428
rect 178 427 179 428
rect 177 427 178 428
rect 176 427 177 428
rect 175 427 176 428
rect 174 427 175 428
rect 173 427 174 428
rect 172 427 173 428
rect 171 427 172 428
rect 170 427 171 428
rect 163 427 164 428
rect 162 427 163 428
rect 161 427 162 428
rect 151 427 152 428
rect 150 427 151 428
rect 149 427 150 428
rect 148 427 149 428
rect 147 427 148 428
rect 146 427 147 428
rect 145 427 146 428
rect 144 427 145 428
rect 143 427 144 428
rect 142 427 143 428
rect 141 427 142 428
rect 140 427 141 428
rect 139 427 140 428
rect 125 427 126 428
rect 124 427 125 428
rect 123 427 124 428
rect 122 427 123 428
rect 121 427 122 428
rect 120 427 121 428
rect 119 427 120 428
rect 118 427 119 428
rect 117 427 118 428
rect 116 427 117 428
rect 115 427 116 428
rect 114 427 115 428
rect 113 427 114 428
rect 112 427 113 428
rect 111 427 112 428
rect 110 427 111 428
rect 109 427 110 428
rect 108 427 109 428
rect 107 427 108 428
rect 106 427 107 428
rect 105 427 106 428
rect 104 427 105 428
rect 103 427 104 428
rect 102 427 103 428
rect 101 427 102 428
rect 194 428 195 429
rect 193 428 194 429
rect 192 428 193 429
rect 191 428 192 429
rect 190 428 191 429
rect 189 428 190 429
rect 188 428 189 429
rect 187 428 188 429
rect 181 428 182 429
rect 180 428 181 429
rect 179 428 180 429
rect 178 428 179 429
rect 177 428 178 429
rect 176 428 177 429
rect 175 428 176 429
rect 174 428 175 429
rect 173 428 174 429
rect 172 428 173 429
rect 171 428 172 429
rect 170 428 171 429
rect 163 428 164 429
rect 162 428 163 429
rect 161 428 162 429
rect 151 428 152 429
rect 150 428 151 429
rect 149 428 150 429
rect 148 428 149 429
rect 147 428 148 429
rect 146 428 147 429
rect 145 428 146 429
rect 144 428 145 429
rect 143 428 144 429
rect 142 428 143 429
rect 141 428 142 429
rect 140 428 141 429
rect 125 428 126 429
rect 124 428 125 429
rect 123 428 124 429
rect 122 428 123 429
rect 121 428 122 429
rect 120 428 121 429
rect 119 428 120 429
rect 118 428 119 429
rect 117 428 118 429
rect 116 428 117 429
rect 115 428 116 429
rect 114 428 115 429
rect 113 428 114 429
rect 112 428 113 429
rect 111 428 112 429
rect 110 428 111 429
rect 109 428 110 429
rect 108 428 109 429
rect 107 428 108 429
rect 106 428 107 429
rect 105 428 106 429
rect 104 428 105 429
rect 103 428 104 429
rect 102 428 103 429
rect 101 428 102 429
rect 195 429 196 430
rect 194 429 195 430
rect 193 429 194 430
rect 192 429 193 430
rect 191 429 192 430
rect 190 429 191 430
rect 189 429 190 430
rect 188 429 189 430
rect 187 429 188 430
rect 181 429 182 430
rect 180 429 181 430
rect 179 429 180 430
rect 178 429 179 430
rect 177 429 178 430
rect 176 429 177 430
rect 175 429 176 430
rect 174 429 175 430
rect 173 429 174 430
rect 172 429 173 430
rect 171 429 172 430
rect 170 429 171 430
rect 163 429 164 430
rect 162 429 163 430
rect 161 429 162 430
rect 151 429 152 430
rect 150 429 151 430
rect 149 429 150 430
rect 148 429 149 430
rect 147 429 148 430
rect 146 429 147 430
rect 145 429 146 430
rect 144 429 145 430
rect 143 429 144 430
rect 142 429 143 430
rect 141 429 142 430
rect 125 429 126 430
rect 124 429 125 430
rect 123 429 124 430
rect 122 429 123 430
rect 121 429 122 430
rect 120 429 121 430
rect 119 429 120 430
rect 118 429 119 430
rect 117 429 118 430
rect 116 429 117 430
rect 115 429 116 430
rect 114 429 115 430
rect 113 429 114 430
rect 112 429 113 430
rect 111 429 112 430
rect 110 429 111 430
rect 109 429 110 430
rect 108 429 109 430
rect 107 429 108 430
rect 106 429 107 430
rect 105 429 106 430
rect 104 429 105 430
rect 103 429 104 430
rect 102 429 103 430
rect 194 430 195 431
rect 193 430 194 431
rect 192 430 193 431
rect 191 430 192 431
rect 190 430 191 431
rect 189 430 190 431
rect 188 430 189 431
rect 187 430 188 431
rect 172 430 173 431
rect 171 430 172 431
rect 170 430 171 431
rect 163 430 164 431
rect 162 430 163 431
rect 161 430 162 431
rect 151 430 152 431
rect 150 430 151 431
rect 149 430 150 431
rect 148 430 149 431
rect 147 430 148 431
rect 146 430 147 431
rect 145 430 146 431
rect 144 430 145 431
rect 143 430 144 431
rect 142 430 143 431
rect 125 430 126 431
rect 124 430 125 431
rect 123 430 124 431
rect 122 430 123 431
rect 121 430 122 431
rect 120 430 121 431
rect 119 430 120 431
rect 118 430 119 431
rect 117 430 118 431
rect 116 430 117 431
rect 115 430 116 431
rect 114 430 115 431
rect 113 430 114 431
rect 112 430 113 431
rect 111 430 112 431
rect 110 430 111 431
rect 109 430 110 431
rect 108 430 109 431
rect 107 430 108 431
rect 106 430 107 431
rect 105 430 106 431
rect 104 430 105 431
rect 103 430 104 431
rect 172 431 173 432
rect 171 431 172 432
rect 170 431 171 432
rect 163 431 164 432
rect 162 431 163 432
rect 161 431 162 432
rect 151 431 152 432
rect 150 431 151 432
rect 149 431 150 432
rect 148 431 149 432
rect 147 431 148 432
rect 146 431 147 432
rect 145 431 146 432
rect 144 431 145 432
rect 143 431 144 432
rect 142 431 143 432
rect 125 431 126 432
rect 124 431 125 432
rect 123 431 124 432
rect 122 431 123 432
rect 121 431 122 432
rect 120 431 121 432
rect 119 431 120 432
rect 118 431 119 432
rect 117 431 118 432
rect 116 431 117 432
rect 115 431 116 432
rect 114 431 115 432
rect 113 431 114 432
rect 112 431 113 432
rect 111 431 112 432
rect 110 431 111 432
rect 109 431 110 432
rect 108 431 109 432
rect 107 431 108 432
rect 106 431 107 432
rect 105 431 106 432
rect 104 431 105 432
rect 194 432 195 433
rect 193 432 194 433
rect 192 432 193 433
rect 191 432 192 433
rect 190 432 191 433
rect 189 432 190 433
rect 172 432 173 433
rect 171 432 172 433
rect 170 432 171 433
rect 163 432 164 433
rect 162 432 163 433
rect 161 432 162 433
rect 151 432 152 433
rect 150 432 151 433
rect 149 432 150 433
rect 148 432 149 433
rect 147 432 148 433
rect 146 432 147 433
rect 145 432 146 433
rect 144 432 145 433
rect 143 432 144 433
rect 125 432 126 433
rect 124 432 125 433
rect 123 432 124 433
rect 122 432 123 433
rect 121 432 122 433
rect 120 432 121 433
rect 119 432 120 433
rect 118 432 119 433
rect 117 432 118 433
rect 116 432 117 433
rect 115 432 116 433
rect 114 432 115 433
rect 113 432 114 433
rect 112 432 113 433
rect 111 432 112 433
rect 110 432 111 433
rect 109 432 110 433
rect 108 432 109 433
rect 107 432 108 433
rect 106 432 107 433
rect 105 432 106 433
rect 195 433 196 434
rect 194 433 195 434
rect 193 433 194 434
rect 192 433 193 434
rect 191 433 192 434
rect 190 433 191 434
rect 189 433 190 434
rect 172 433 173 434
rect 171 433 172 434
rect 170 433 171 434
rect 169 433 170 434
rect 168 433 169 434
rect 167 433 168 434
rect 166 433 167 434
rect 165 433 166 434
rect 164 433 165 434
rect 163 433 164 434
rect 162 433 163 434
rect 161 433 162 434
rect 151 433 152 434
rect 150 433 151 434
rect 149 433 150 434
rect 148 433 149 434
rect 147 433 148 434
rect 146 433 147 434
rect 145 433 146 434
rect 144 433 145 434
rect 125 433 126 434
rect 124 433 125 434
rect 123 433 124 434
rect 122 433 123 434
rect 121 433 122 434
rect 120 433 121 434
rect 119 433 120 434
rect 118 433 119 434
rect 117 433 118 434
rect 116 433 117 434
rect 115 433 116 434
rect 114 433 115 434
rect 113 433 114 434
rect 112 433 113 434
rect 111 433 112 434
rect 110 433 111 434
rect 109 433 110 434
rect 108 433 109 434
rect 107 433 108 434
rect 106 433 107 434
rect 190 434 191 435
rect 189 434 190 435
rect 172 434 173 435
rect 171 434 172 435
rect 170 434 171 435
rect 169 434 170 435
rect 168 434 169 435
rect 167 434 168 435
rect 166 434 167 435
rect 165 434 166 435
rect 164 434 165 435
rect 163 434 164 435
rect 162 434 163 435
rect 161 434 162 435
rect 151 434 152 435
rect 150 434 151 435
rect 149 434 150 435
rect 148 434 149 435
rect 147 434 148 435
rect 146 434 147 435
rect 145 434 146 435
rect 190 435 191 436
rect 189 435 190 436
rect 172 435 173 436
rect 171 435 172 436
rect 170 435 171 436
rect 169 435 170 436
rect 168 435 169 436
rect 167 435 168 436
rect 166 435 167 436
rect 165 435 166 436
rect 164 435 165 436
rect 163 435 164 436
rect 162 435 163 436
rect 161 435 162 436
rect 151 435 152 436
rect 150 435 151 436
rect 149 435 150 436
rect 148 435 149 436
rect 147 435 148 436
rect 146 435 147 436
rect 194 436 195 437
rect 193 436 194 437
rect 192 436 193 437
rect 191 436 192 437
rect 190 436 191 437
rect 189 436 190 437
rect 172 436 173 437
rect 171 436 172 437
rect 170 436 171 437
rect 168 436 169 437
rect 167 436 168 437
rect 166 436 167 437
rect 165 436 166 437
rect 164 436 165 437
rect 163 436 164 437
rect 162 436 163 437
rect 161 436 162 437
rect 151 436 152 437
rect 150 436 151 437
rect 149 436 150 437
rect 148 436 149 437
rect 147 436 148 437
rect 195 437 196 438
rect 194 437 195 438
rect 193 437 194 438
rect 192 437 193 438
rect 191 437 192 438
rect 190 437 191 438
rect 189 437 190 438
rect 172 437 173 438
rect 171 437 172 438
rect 170 437 171 438
rect 165 437 166 438
rect 164 437 165 438
rect 163 437 164 438
rect 162 437 163 438
rect 161 437 162 438
rect 151 437 152 438
rect 150 437 151 438
rect 149 437 150 438
rect 148 437 149 438
rect 147 437 148 438
rect 190 438 191 439
rect 172 438 173 439
rect 171 438 172 439
rect 170 438 171 439
rect 151 438 152 439
rect 150 438 151 439
rect 149 438 150 439
rect 148 438 149 439
rect 194 439 195 440
rect 191 439 192 440
rect 190 439 191 440
rect 172 439 173 440
rect 171 439 172 440
rect 170 439 171 440
rect 151 439 152 440
rect 150 439 151 440
rect 149 439 150 440
rect 195 440 196 441
rect 194 440 195 441
rect 192 440 193 441
rect 191 440 192 441
rect 190 440 191 441
rect 189 440 190 441
rect 172 440 173 441
rect 171 440 172 441
rect 170 440 171 441
rect 151 440 152 441
rect 150 440 151 441
rect 195 441 196 442
rect 194 441 195 442
rect 193 441 194 442
rect 192 441 193 442
rect 191 441 192 442
rect 190 441 191 442
rect 189 441 190 442
rect 151 441 152 442
rect 150 441 151 442
rect 194 442 195 443
rect 193 442 194 443
rect 192 442 193 443
rect 190 442 191 443
rect 189 442 190 443
rect 194 443 195 444
rect 193 443 194 444
rect 192 443 193 444
rect 190 444 191 445
rect 189 444 190 445
rect 194 445 195 446
rect 193 445 194 446
rect 192 445 193 446
rect 191 445 192 446
rect 190 445 191 446
rect 189 445 190 446
rect 188 445 189 446
rect 195 446 196 447
rect 194 446 195 447
rect 193 446 194 447
rect 192 446 193 447
rect 191 446 192 447
rect 190 446 191 447
rect 189 446 190 447
rect 188 446 189 447
rect 187 446 188 447
rect 195 447 196 448
rect 194 447 195 448
rect 190 447 191 448
rect 189 447 190 448
rect 194 448 195 449
rect 194 449 195 450
rect 193 449 194 450
rect 192 449 193 450
rect 191 449 192 450
rect 190 449 191 450
rect 189 449 190 450
rect 187 449 188 450
rect 186 449 187 450
rect 195 450 196 451
rect 194 450 195 451
rect 193 450 194 451
rect 192 450 193 451
rect 191 450 192 451
rect 190 450 191 451
rect 189 450 190 451
rect 187 450 188 451
rect 186 450 187 451
rect 171 451 172 452
rect 170 451 171 452
rect 169 451 170 452
rect 147 451 148 452
rect 146 451 147 452
rect 145 451 146 452
rect 144 451 145 452
rect 143 451 144 452
rect 142 451 143 452
rect 141 451 142 452
rect 140 451 141 452
rect 139 451 140 452
rect 138 451 139 452
rect 137 451 138 452
rect 136 451 137 452
rect 135 451 136 452
rect 134 451 135 452
rect 133 451 134 452
rect 132 451 133 452
rect 131 451 132 452
rect 130 451 131 452
rect 129 451 130 452
rect 128 451 129 452
rect 127 451 128 452
rect 126 451 127 452
rect 125 451 126 452
rect 124 451 125 452
rect 123 451 124 452
rect 122 451 123 452
rect 121 451 122 452
rect 120 451 121 452
rect 119 451 120 452
rect 118 451 119 452
rect 117 451 118 452
rect 116 451 117 452
rect 115 451 116 452
rect 114 451 115 452
rect 113 451 114 452
rect 112 451 113 452
rect 111 451 112 452
rect 110 451 111 452
rect 109 451 110 452
rect 108 451 109 452
rect 107 451 108 452
rect 106 451 107 452
rect 105 451 106 452
rect 104 451 105 452
rect 103 451 104 452
rect 102 451 103 452
rect 101 451 102 452
rect 100 451 101 452
rect 190 452 191 453
rect 189 452 190 453
rect 171 452 172 453
rect 170 452 171 453
rect 169 452 170 453
rect 168 452 169 453
rect 147 452 148 453
rect 146 452 147 453
rect 145 452 146 453
rect 144 452 145 453
rect 143 452 144 453
rect 142 452 143 453
rect 141 452 142 453
rect 140 452 141 453
rect 139 452 140 453
rect 138 452 139 453
rect 137 452 138 453
rect 136 452 137 453
rect 135 452 136 453
rect 134 452 135 453
rect 133 452 134 453
rect 132 452 133 453
rect 131 452 132 453
rect 130 452 131 453
rect 129 452 130 453
rect 128 452 129 453
rect 127 452 128 453
rect 126 452 127 453
rect 125 452 126 453
rect 124 452 125 453
rect 123 452 124 453
rect 122 452 123 453
rect 121 452 122 453
rect 120 452 121 453
rect 119 452 120 453
rect 118 452 119 453
rect 117 452 118 453
rect 116 452 117 453
rect 115 452 116 453
rect 114 452 115 453
rect 113 452 114 453
rect 112 452 113 453
rect 111 452 112 453
rect 110 452 111 453
rect 109 452 110 453
rect 108 452 109 453
rect 107 452 108 453
rect 106 452 107 453
rect 105 452 106 453
rect 104 452 105 453
rect 103 452 104 453
rect 102 452 103 453
rect 101 452 102 453
rect 100 452 101 453
rect 194 453 195 454
rect 193 453 194 454
rect 192 453 193 454
rect 191 453 192 454
rect 190 453 191 454
rect 189 453 190 454
rect 188 453 189 454
rect 187 453 188 454
rect 171 453 172 454
rect 170 453 171 454
rect 169 453 170 454
rect 168 453 169 454
rect 165 453 166 454
rect 164 453 165 454
rect 163 453 164 454
rect 162 453 163 454
rect 147 453 148 454
rect 146 453 147 454
rect 145 453 146 454
rect 144 453 145 454
rect 143 453 144 454
rect 142 453 143 454
rect 141 453 142 454
rect 140 453 141 454
rect 139 453 140 454
rect 138 453 139 454
rect 137 453 138 454
rect 136 453 137 454
rect 135 453 136 454
rect 134 453 135 454
rect 133 453 134 454
rect 132 453 133 454
rect 131 453 132 454
rect 130 453 131 454
rect 129 453 130 454
rect 128 453 129 454
rect 127 453 128 454
rect 126 453 127 454
rect 125 453 126 454
rect 124 453 125 454
rect 123 453 124 454
rect 122 453 123 454
rect 121 453 122 454
rect 120 453 121 454
rect 119 453 120 454
rect 118 453 119 454
rect 117 453 118 454
rect 116 453 117 454
rect 115 453 116 454
rect 114 453 115 454
rect 113 453 114 454
rect 112 453 113 454
rect 111 453 112 454
rect 110 453 111 454
rect 109 453 110 454
rect 108 453 109 454
rect 107 453 108 454
rect 106 453 107 454
rect 105 453 106 454
rect 104 453 105 454
rect 103 453 104 454
rect 102 453 103 454
rect 101 453 102 454
rect 100 453 101 454
rect 195 454 196 455
rect 194 454 195 455
rect 193 454 194 455
rect 192 454 193 455
rect 191 454 192 455
rect 190 454 191 455
rect 189 454 190 455
rect 188 454 189 455
rect 187 454 188 455
rect 171 454 172 455
rect 170 454 171 455
rect 169 454 170 455
rect 168 454 169 455
rect 166 454 167 455
rect 165 454 166 455
rect 164 454 165 455
rect 163 454 164 455
rect 162 454 163 455
rect 161 454 162 455
rect 147 454 148 455
rect 146 454 147 455
rect 145 454 146 455
rect 144 454 145 455
rect 143 454 144 455
rect 142 454 143 455
rect 141 454 142 455
rect 140 454 141 455
rect 139 454 140 455
rect 138 454 139 455
rect 137 454 138 455
rect 136 454 137 455
rect 135 454 136 455
rect 134 454 135 455
rect 133 454 134 455
rect 132 454 133 455
rect 131 454 132 455
rect 130 454 131 455
rect 129 454 130 455
rect 128 454 129 455
rect 127 454 128 455
rect 126 454 127 455
rect 125 454 126 455
rect 124 454 125 455
rect 123 454 124 455
rect 122 454 123 455
rect 121 454 122 455
rect 120 454 121 455
rect 119 454 120 455
rect 118 454 119 455
rect 117 454 118 455
rect 116 454 117 455
rect 115 454 116 455
rect 114 454 115 455
rect 113 454 114 455
rect 112 454 113 455
rect 111 454 112 455
rect 110 454 111 455
rect 109 454 110 455
rect 108 454 109 455
rect 107 454 108 455
rect 106 454 107 455
rect 105 454 106 455
rect 104 454 105 455
rect 103 454 104 455
rect 102 454 103 455
rect 101 454 102 455
rect 100 454 101 455
rect 195 455 196 456
rect 194 455 195 456
rect 190 455 191 456
rect 189 455 190 456
rect 181 455 182 456
rect 180 455 181 456
rect 179 455 180 456
rect 178 455 179 456
rect 177 455 178 456
rect 176 455 177 456
rect 171 455 172 456
rect 170 455 171 456
rect 169 455 170 456
rect 168 455 169 456
rect 166 455 167 456
rect 165 455 166 456
rect 164 455 165 456
rect 163 455 164 456
rect 162 455 163 456
rect 161 455 162 456
rect 160 455 161 456
rect 147 455 148 456
rect 146 455 147 456
rect 145 455 146 456
rect 144 455 145 456
rect 143 455 144 456
rect 142 455 143 456
rect 141 455 142 456
rect 140 455 141 456
rect 139 455 140 456
rect 138 455 139 456
rect 137 455 138 456
rect 136 455 137 456
rect 135 455 136 456
rect 134 455 135 456
rect 133 455 134 456
rect 132 455 133 456
rect 131 455 132 456
rect 130 455 131 456
rect 129 455 130 456
rect 128 455 129 456
rect 127 455 128 456
rect 126 455 127 456
rect 125 455 126 456
rect 124 455 125 456
rect 123 455 124 456
rect 122 455 123 456
rect 121 455 122 456
rect 120 455 121 456
rect 119 455 120 456
rect 118 455 119 456
rect 117 455 118 456
rect 116 455 117 456
rect 115 455 116 456
rect 114 455 115 456
rect 113 455 114 456
rect 112 455 113 456
rect 111 455 112 456
rect 110 455 111 456
rect 109 455 110 456
rect 108 455 109 456
rect 107 455 108 456
rect 106 455 107 456
rect 105 455 106 456
rect 104 455 105 456
rect 103 455 104 456
rect 102 455 103 456
rect 101 455 102 456
rect 100 455 101 456
rect 194 456 195 457
rect 181 456 182 457
rect 180 456 181 457
rect 179 456 180 457
rect 178 456 179 457
rect 177 456 178 457
rect 176 456 177 457
rect 171 456 172 457
rect 170 456 171 457
rect 169 456 170 457
rect 168 456 169 457
rect 167 456 168 457
rect 166 456 167 457
rect 165 456 166 457
rect 164 456 165 457
rect 163 456 164 457
rect 162 456 163 457
rect 161 456 162 457
rect 160 456 161 457
rect 147 456 148 457
rect 146 456 147 457
rect 145 456 146 457
rect 144 456 145 457
rect 143 456 144 457
rect 142 456 143 457
rect 141 456 142 457
rect 140 456 141 457
rect 139 456 140 457
rect 138 456 139 457
rect 137 456 138 457
rect 136 456 137 457
rect 135 456 136 457
rect 134 456 135 457
rect 133 456 134 457
rect 132 456 133 457
rect 131 456 132 457
rect 130 456 131 457
rect 129 456 130 457
rect 128 456 129 457
rect 127 456 128 457
rect 126 456 127 457
rect 125 456 126 457
rect 124 456 125 457
rect 123 456 124 457
rect 122 456 123 457
rect 121 456 122 457
rect 120 456 121 457
rect 119 456 120 457
rect 118 456 119 457
rect 117 456 118 457
rect 116 456 117 457
rect 115 456 116 457
rect 114 456 115 457
rect 113 456 114 457
rect 112 456 113 457
rect 111 456 112 457
rect 110 456 111 457
rect 109 456 110 457
rect 108 456 109 457
rect 107 456 108 457
rect 106 456 107 457
rect 105 456 106 457
rect 104 456 105 457
rect 103 456 104 457
rect 102 456 103 457
rect 101 456 102 457
rect 100 456 101 457
rect 194 457 195 458
rect 193 457 194 458
rect 192 457 193 458
rect 191 457 192 458
rect 190 457 191 458
rect 189 457 190 458
rect 181 457 182 458
rect 180 457 181 458
rect 179 457 180 458
rect 178 457 179 458
rect 177 457 178 458
rect 176 457 177 458
rect 175 457 176 458
rect 174 457 175 458
rect 173 457 174 458
rect 172 457 173 458
rect 171 457 172 458
rect 170 457 171 458
rect 169 457 170 458
rect 168 457 169 458
rect 167 457 168 458
rect 166 457 167 458
rect 165 457 166 458
rect 164 457 165 458
rect 162 457 163 458
rect 161 457 162 458
rect 160 457 161 458
rect 159 457 160 458
rect 147 457 148 458
rect 146 457 147 458
rect 145 457 146 458
rect 144 457 145 458
rect 143 457 144 458
rect 142 457 143 458
rect 141 457 142 458
rect 140 457 141 458
rect 139 457 140 458
rect 138 457 139 458
rect 137 457 138 458
rect 136 457 137 458
rect 135 457 136 458
rect 134 457 135 458
rect 133 457 134 458
rect 132 457 133 458
rect 131 457 132 458
rect 130 457 131 458
rect 129 457 130 458
rect 128 457 129 458
rect 127 457 128 458
rect 126 457 127 458
rect 125 457 126 458
rect 124 457 125 458
rect 123 457 124 458
rect 122 457 123 458
rect 121 457 122 458
rect 120 457 121 458
rect 119 457 120 458
rect 118 457 119 458
rect 117 457 118 458
rect 116 457 117 458
rect 115 457 116 458
rect 114 457 115 458
rect 113 457 114 458
rect 112 457 113 458
rect 111 457 112 458
rect 110 457 111 458
rect 109 457 110 458
rect 108 457 109 458
rect 107 457 108 458
rect 106 457 107 458
rect 105 457 106 458
rect 104 457 105 458
rect 103 457 104 458
rect 102 457 103 458
rect 101 457 102 458
rect 100 457 101 458
rect 195 458 196 459
rect 194 458 195 459
rect 193 458 194 459
rect 192 458 193 459
rect 191 458 192 459
rect 190 458 191 459
rect 189 458 190 459
rect 181 458 182 459
rect 180 458 181 459
rect 179 458 180 459
rect 178 458 179 459
rect 177 458 178 459
rect 176 458 177 459
rect 175 458 176 459
rect 174 458 175 459
rect 173 458 174 459
rect 172 458 173 459
rect 171 458 172 459
rect 170 458 171 459
rect 169 458 170 459
rect 168 458 169 459
rect 167 458 168 459
rect 166 458 167 459
rect 165 458 166 459
rect 161 458 162 459
rect 160 458 161 459
rect 159 458 160 459
rect 147 458 148 459
rect 146 458 147 459
rect 145 458 146 459
rect 144 458 145 459
rect 143 458 144 459
rect 142 458 143 459
rect 141 458 142 459
rect 140 458 141 459
rect 139 458 140 459
rect 138 458 139 459
rect 137 458 138 459
rect 136 458 137 459
rect 135 458 136 459
rect 134 458 135 459
rect 133 458 134 459
rect 132 458 133 459
rect 131 458 132 459
rect 130 458 131 459
rect 129 458 130 459
rect 128 458 129 459
rect 127 458 128 459
rect 126 458 127 459
rect 125 458 126 459
rect 124 458 125 459
rect 123 458 124 459
rect 122 458 123 459
rect 121 458 122 459
rect 120 458 121 459
rect 119 458 120 459
rect 118 458 119 459
rect 117 458 118 459
rect 116 458 117 459
rect 115 458 116 459
rect 114 458 115 459
rect 113 458 114 459
rect 112 458 113 459
rect 111 458 112 459
rect 110 458 111 459
rect 109 458 110 459
rect 108 458 109 459
rect 107 458 108 459
rect 106 458 107 459
rect 105 458 106 459
rect 104 458 105 459
rect 103 458 104 459
rect 102 458 103 459
rect 101 458 102 459
rect 100 458 101 459
rect 195 459 196 460
rect 194 459 195 460
rect 181 459 182 460
rect 180 459 181 460
rect 179 459 180 460
rect 178 459 179 460
rect 174 459 175 460
rect 173 459 174 460
rect 172 459 173 460
rect 171 459 172 460
rect 170 459 171 460
rect 169 459 170 460
rect 168 459 169 460
rect 167 459 168 460
rect 166 459 167 460
rect 165 459 166 460
rect 161 459 162 460
rect 160 459 161 460
rect 159 459 160 460
rect 147 459 148 460
rect 146 459 147 460
rect 145 459 146 460
rect 144 459 145 460
rect 143 459 144 460
rect 142 459 143 460
rect 141 459 142 460
rect 140 459 141 460
rect 139 459 140 460
rect 138 459 139 460
rect 137 459 138 460
rect 136 459 137 460
rect 135 459 136 460
rect 134 459 135 460
rect 133 459 134 460
rect 132 459 133 460
rect 131 459 132 460
rect 130 459 131 460
rect 129 459 130 460
rect 128 459 129 460
rect 127 459 128 460
rect 126 459 127 460
rect 125 459 126 460
rect 124 459 125 460
rect 123 459 124 460
rect 122 459 123 460
rect 121 459 122 460
rect 120 459 121 460
rect 119 459 120 460
rect 118 459 119 460
rect 117 459 118 460
rect 116 459 117 460
rect 115 459 116 460
rect 114 459 115 460
rect 113 459 114 460
rect 112 459 113 460
rect 111 459 112 460
rect 110 459 111 460
rect 109 459 110 460
rect 108 459 109 460
rect 107 459 108 460
rect 106 459 107 460
rect 105 459 106 460
rect 104 459 105 460
rect 103 459 104 460
rect 102 459 103 460
rect 101 459 102 460
rect 100 459 101 460
rect 194 460 195 461
rect 181 460 182 461
rect 180 460 181 461
rect 179 460 180 461
rect 178 460 179 461
rect 171 460 172 461
rect 170 460 171 461
rect 169 460 170 461
rect 168 460 169 461
rect 167 460 168 461
rect 166 460 167 461
rect 165 460 166 461
rect 161 460 162 461
rect 160 460 161 461
rect 159 460 160 461
rect 147 460 148 461
rect 146 460 147 461
rect 145 460 146 461
rect 144 460 145 461
rect 143 460 144 461
rect 142 460 143 461
rect 141 460 142 461
rect 140 460 141 461
rect 139 460 140 461
rect 138 460 139 461
rect 137 460 138 461
rect 136 460 137 461
rect 135 460 136 461
rect 134 460 135 461
rect 133 460 134 461
rect 132 460 133 461
rect 131 460 132 461
rect 130 460 131 461
rect 129 460 130 461
rect 128 460 129 461
rect 127 460 128 461
rect 126 460 127 461
rect 125 460 126 461
rect 124 460 125 461
rect 123 460 124 461
rect 122 460 123 461
rect 121 460 122 461
rect 120 460 121 461
rect 119 460 120 461
rect 118 460 119 461
rect 117 460 118 461
rect 116 460 117 461
rect 115 460 116 461
rect 114 460 115 461
rect 113 460 114 461
rect 112 460 113 461
rect 111 460 112 461
rect 110 460 111 461
rect 109 460 110 461
rect 108 460 109 461
rect 107 460 108 461
rect 106 460 107 461
rect 105 460 106 461
rect 104 460 105 461
rect 103 460 104 461
rect 102 460 103 461
rect 101 460 102 461
rect 100 460 101 461
rect 195 461 196 462
rect 194 461 195 462
rect 193 461 194 462
rect 192 461 193 462
rect 191 461 192 462
rect 190 461 191 462
rect 189 461 190 462
rect 181 461 182 462
rect 180 461 181 462
rect 179 461 180 462
rect 178 461 179 462
rect 171 461 172 462
rect 170 461 171 462
rect 169 461 170 462
rect 168 461 169 462
rect 167 461 168 462
rect 166 461 167 462
rect 165 461 166 462
rect 161 461 162 462
rect 160 461 161 462
rect 159 461 160 462
rect 147 461 148 462
rect 146 461 147 462
rect 145 461 146 462
rect 144 461 145 462
rect 143 461 144 462
rect 142 461 143 462
rect 141 461 142 462
rect 140 461 141 462
rect 139 461 140 462
rect 138 461 139 462
rect 137 461 138 462
rect 136 461 137 462
rect 135 461 136 462
rect 134 461 135 462
rect 133 461 134 462
rect 132 461 133 462
rect 131 461 132 462
rect 130 461 131 462
rect 129 461 130 462
rect 128 461 129 462
rect 127 461 128 462
rect 126 461 127 462
rect 125 461 126 462
rect 124 461 125 462
rect 123 461 124 462
rect 122 461 123 462
rect 121 461 122 462
rect 120 461 121 462
rect 119 461 120 462
rect 118 461 119 462
rect 117 461 118 462
rect 116 461 117 462
rect 115 461 116 462
rect 114 461 115 462
rect 113 461 114 462
rect 112 461 113 462
rect 111 461 112 462
rect 110 461 111 462
rect 109 461 110 462
rect 108 461 109 462
rect 107 461 108 462
rect 106 461 107 462
rect 105 461 106 462
rect 104 461 105 462
rect 103 461 104 462
rect 102 461 103 462
rect 101 461 102 462
rect 100 461 101 462
rect 194 462 195 463
rect 193 462 194 463
rect 192 462 193 463
rect 191 462 192 463
rect 190 462 191 463
rect 189 462 190 463
rect 181 462 182 463
rect 180 462 181 463
rect 179 462 180 463
rect 178 462 179 463
rect 171 462 172 463
rect 170 462 171 463
rect 169 462 170 463
rect 168 462 169 463
rect 167 462 168 463
rect 166 462 167 463
rect 165 462 166 463
rect 164 462 165 463
rect 162 462 163 463
rect 161 462 162 463
rect 160 462 161 463
rect 147 462 148 463
rect 146 462 147 463
rect 145 462 146 463
rect 144 462 145 463
rect 143 462 144 463
rect 142 462 143 463
rect 141 462 142 463
rect 140 462 141 463
rect 139 462 140 463
rect 138 462 139 463
rect 137 462 138 463
rect 136 462 137 463
rect 135 462 136 463
rect 134 462 135 463
rect 133 462 134 463
rect 132 462 133 463
rect 131 462 132 463
rect 130 462 131 463
rect 129 462 130 463
rect 128 462 129 463
rect 127 462 128 463
rect 126 462 127 463
rect 125 462 126 463
rect 124 462 125 463
rect 123 462 124 463
rect 122 462 123 463
rect 121 462 122 463
rect 120 462 121 463
rect 119 462 120 463
rect 118 462 119 463
rect 117 462 118 463
rect 116 462 117 463
rect 115 462 116 463
rect 114 462 115 463
rect 113 462 114 463
rect 112 462 113 463
rect 111 462 112 463
rect 110 462 111 463
rect 109 462 110 463
rect 108 462 109 463
rect 107 462 108 463
rect 106 462 107 463
rect 105 462 106 463
rect 104 462 105 463
rect 103 462 104 463
rect 102 462 103 463
rect 101 462 102 463
rect 100 462 101 463
rect 181 463 182 464
rect 180 463 181 464
rect 179 463 180 464
rect 178 463 179 464
rect 171 463 172 464
rect 170 463 171 464
rect 169 463 170 464
rect 168 463 169 464
rect 166 463 167 464
rect 165 463 166 464
rect 164 463 165 464
rect 163 463 164 464
rect 162 463 163 464
rect 161 463 162 464
rect 160 463 161 464
rect 147 463 148 464
rect 146 463 147 464
rect 145 463 146 464
rect 144 463 145 464
rect 143 463 144 464
rect 142 463 143 464
rect 141 463 142 464
rect 140 463 141 464
rect 139 463 140 464
rect 138 463 139 464
rect 137 463 138 464
rect 136 463 137 464
rect 135 463 136 464
rect 134 463 135 464
rect 133 463 134 464
rect 132 463 133 464
rect 131 463 132 464
rect 130 463 131 464
rect 129 463 130 464
rect 128 463 129 464
rect 127 463 128 464
rect 126 463 127 464
rect 125 463 126 464
rect 124 463 125 464
rect 123 463 124 464
rect 122 463 123 464
rect 121 463 122 464
rect 120 463 121 464
rect 119 463 120 464
rect 118 463 119 464
rect 117 463 118 464
rect 116 463 117 464
rect 115 463 116 464
rect 114 463 115 464
rect 113 463 114 464
rect 112 463 113 464
rect 111 463 112 464
rect 110 463 111 464
rect 109 463 110 464
rect 108 463 109 464
rect 107 463 108 464
rect 106 463 107 464
rect 105 463 106 464
rect 104 463 105 464
rect 103 463 104 464
rect 102 463 103 464
rect 101 463 102 464
rect 100 463 101 464
rect 193 464 194 465
rect 192 464 193 465
rect 191 464 192 465
rect 190 464 191 465
rect 189 464 190 465
rect 188 464 189 465
rect 181 464 182 465
rect 180 464 181 465
rect 179 464 180 465
rect 178 464 179 465
rect 174 464 175 465
rect 173 464 174 465
rect 172 464 173 465
rect 171 464 172 465
rect 170 464 171 465
rect 169 464 170 465
rect 168 464 169 465
rect 166 464 167 465
rect 165 464 166 465
rect 164 464 165 465
rect 163 464 164 465
rect 162 464 163 465
rect 161 464 162 465
rect 147 464 148 465
rect 146 464 147 465
rect 145 464 146 465
rect 144 464 145 465
rect 143 464 144 465
rect 142 464 143 465
rect 141 464 142 465
rect 140 464 141 465
rect 139 464 140 465
rect 138 464 139 465
rect 137 464 138 465
rect 136 464 137 465
rect 135 464 136 465
rect 134 464 135 465
rect 133 464 134 465
rect 132 464 133 465
rect 131 464 132 465
rect 130 464 131 465
rect 129 464 130 465
rect 128 464 129 465
rect 127 464 128 465
rect 126 464 127 465
rect 125 464 126 465
rect 124 464 125 465
rect 123 464 124 465
rect 122 464 123 465
rect 121 464 122 465
rect 120 464 121 465
rect 119 464 120 465
rect 118 464 119 465
rect 117 464 118 465
rect 116 464 117 465
rect 115 464 116 465
rect 114 464 115 465
rect 113 464 114 465
rect 112 464 113 465
rect 111 464 112 465
rect 110 464 111 465
rect 109 464 110 465
rect 108 464 109 465
rect 107 464 108 465
rect 106 464 107 465
rect 105 464 106 465
rect 104 464 105 465
rect 103 464 104 465
rect 102 464 103 465
rect 101 464 102 465
rect 100 464 101 465
rect 194 465 195 466
rect 193 465 194 466
rect 192 465 193 466
rect 191 465 192 466
rect 190 465 191 466
rect 189 465 190 466
rect 188 465 189 466
rect 187 465 188 466
rect 181 465 182 466
rect 180 465 181 466
rect 179 465 180 466
rect 178 465 179 466
rect 174 465 175 466
rect 173 465 174 466
rect 172 465 173 466
rect 171 465 172 466
rect 170 465 171 466
rect 169 465 170 466
rect 168 465 169 466
rect 165 465 166 466
rect 164 465 165 466
rect 163 465 164 466
rect 162 465 163 466
rect 161 465 162 466
rect 147 465 148 466
rect 146 465 147 466
rect 145 465 146 466
rect 144 465 145 466
rect 143 465 144 466
rect 142 465 143 466
rect 141 465 142 466
rect 140 465 141 466
rect 139 465 140 466
rect 138 465 139 466
rect 137 465 138 466
rect 136 465 137 466
rect 135 465 136 466
rect 134 465 135 466
rect 133 465 134 466
rect 132 465 133 466
rect 131 465 132 466
rect 130 465 131 466
rect 129 465 130 466
rect 128 465 129 466
rect 127 465 128 466
rect 126 465 127 466
rect 125 465 126 466
rect 124 465 125 466
rect 123 465 124 466
rect 122 465 123 466
rect 121 465 122 466
rect 120 465 121 466
rect 119 465 120 466
rect 118 465 119 466
rect 117 465 118 466
rect 116 465 117 466
rect 115 465 116 466
rect 114 465 115 466
rect 113 465 114 466
rect 112 465 113 466
rect 111 465 112 466
rect 110 465 111 466
rect 109 465 110 466
rect 108 465 109 466
rect 107 465 108 466
rect 106 465 107 466
rect 105 465 106 466
rect 104 465 105 466
rect 103 465 104 466
rect 102 465 103 466
rect 101 465 102 466
rect 100 465 101 466
rect 194 466 195 467
rect 193 466 194 467
rect 192 466 193 467
rect 191 466 192 467
rect 190 466 191 467
rect 189 466 190 467
rect 188 466 189 467
rect 187 466 188 467
rect 181 466 182 467
rect 180 466 181 467
rect 179 466 180 467
rect 178 466 179 467
rect 174 466 175 467
rect 173 466 174 467
rect 172 466 173 467
rect 171 466 172 467
rect 170 466 171 467
rect 169 466 170 467
rect 168 466 169 467
rect 164 466 165 467
rect 163 466 164 467
rect 162 466 163 467
rect 147 466 148 467
rect 146 466 147 467
rect 145 466 146 467
rect 144 466 145 467
rect 143 466 144 467
rect 142 466 143 467
rect 141 466 142 467
rect 140 466 141 467
rect 139 466 140 467
rect 138 466 139 467
rect 137 466 138 467
rect 136 466 137 467
rect 135 466 136 467
rect 134 466 135 467
rect 133 466 134 467
rect 132 466 133 467
rect 131 466 132 467
rect 130 466 131 467
rect 129 466 130 467
rect 128 466 129 467
rect 127 466 128 467
rect 126 466 127 467
rect 125 466 126 467
rect 124 466 125 467
rect 123 466 124 467
rect 122 466 123 467
rect 121 466 122 467
rect 120 466 121 467
rect 119 466 120 467
rect 118 466 119 467
rect 117 466 118 467
rect 116 466 117 467
rect 115 466 116 467
rect 114 466 115 467
rect 113 466 114 467
rect 112 466 113 467
rect 111 466 112 467
rect 110 466 111 467
rect 109 466 110 467
rect 108 466 109 467
rect 107 466 108 467
rect 106 466 107 467
rect 105 466 106 467
rect 104 466 105 467
rect 103 466 104 467
rect 102 466 103 467
rect 101 466 102 467
rect 100 466 101 467
rect 195 467 196 468
rect 194 467 195 468
rect 190 467 191 468
rect 189 467 190 468
rect 181 467 182 468
rect 180 467 181 468
rect 179 467 180 468
rect 178 467 179 468
rect 174 467 175 468
rect 173 467 174 468
rect 172 467 173 468
rect 170 467 171 468
rect 169 467 170 468
rect 168 467 169 468
rect 147 467 148 468
rect 146 467 147 468
rect 145 467 146 468
rect 144 467 145 468
rect 143 467 144 468
rect 142 467 143 468
rect 141 467 142 468
rect 140 467 141 468
rect 139 467 140 468
rect 138 467 139 468
rect 137 467 138 468
rect 136 467 137 468
rect 135 467 136 468
rect 134 467 135 468
rect 133 467 134 468
rect 132 467 133 468
rect 131 467 132 468
rect 130 467 131 468
rect 129 467 130 468
rect 128 467 129 468
rect 127 467 128 468
rect 126 467 127 468
rect 125 467 126 468
rect 124 467 125 468
rect 123 467 124 468
rect 122 467 123 468
rect 121 467 122 468
rect 120 467 121 468
rect 119 467 120 468
rect 118 467 119 468
rect 117 467 118 468
rect 116 467 117 468
rect 115 467 116 468
rect 114 467 115 468
rect 113 467 114 468
rect 112 467 113 468
rect 111 467 112 468
rect 110 467 111 468
rect 109 467 110 468
rect 108 467 109 468
rect 107 467 108 468
rect 106 467 107 468
rect 105 467 106 468
rect 104 467 105 468
rect 103 467 104 468
rect 102 467 103 468
rect 101 467 102 468
rect 100 467 101 468
rect 193 468 194 469
rect 192 468 193 469
rect 191 468 192 469
rect 181 468 182 469
rect 180 468 181 469
rect 179 468 180 469
rect 178 468 179 469
rect 174 468 175 469
rect 173 468 174 469
rect 172 468 173 469
rect 170 468 171 469
rect 169 468 170 469
rect 168 468 169 469
rect 147 468 148 469
rect 146 468 147 469
rect 145 468 146 469
rect 144 468 145 469
rect 143 468 144 469
rect 142 468 143 469
rect 141 468 142 469
rect 140 468 141 469
rect 139 468 140 469
rect 138 468 139 469
rect 137 468 138 469
rect 136 468 137 469
rect 135 468 136 469
rect 134 468 135 469
rect 133 468 134 469
rect 132 468 133 469
rect 131 468 132 469
rect 130 468 131 469
rect 129 468 130 469
rect 128 468 129 469
rect 127 468 128 469
rect 126 468 127 469
rect 125 468 126 469
rect 124 468 125 469
rect 123 468 124 469
rect 122 468 123 469
rect 121 468 122 469
rect 120 468 121 469
rect 119 468 120 469
rect 118 468 119 469
rect 117 468 118 469
rect 116 468 117 469
rect 115 468 116 469
rect 114 468 115 469
rect 113 468 114 469
rect 112 468 113 469
rect 111 468 112 469
rect 110 468 111 469
rect 109 468 110 469
rect 108 468 109 469
rect 107 468 108 469
rect 106 468 107 469
rect 105 468 106 469
rect 104 468 105 469
rect 103 468 104 469
rect 102 468 103 469
rect 101 468 102 469
rect 100 468 101 469
rect 194 469 195 470
rect 193 469 194 470
rect 192 469 193 470
rect 191 469 192 470
rect 190 469 191 470
rect 189 469 190 470
rect 181 469 182 470
rect 180 469 181 470
rect 179 469 180 470
rect 178 469 179 470
rect 174 469 175 470
rect 173 469 174 470
rect 172 469 173 470
rect 171 469 172 470
rect 147 469 148 470
rect 146 469 147 470
rect 145 469 146 470
rect 144 469 145 470
rect 143 469 144 470
rect 142 469 143 470
rect 141 469 142 470
rect 140 469 141 470
rect 139 469 140 470
rect 138 469 139 470
rect 137 469 138 470
rect 136 469 137 470
rect 135 469 136 470
rect 134 469 135 470
rect 133 469 134 470
rect 132 469 133 470
rect 131 469 132 470
rect 130 469 131 470
rect 129 469 130 470
rect 128 469 129 470
rect 127 469 128 470
rect 126 469 127 470
rect 125 469 126 470
rect 124 469 125 470
rect 123 469 124 470
rect 122 469 123 470
rect 121 469 122 470
rect 120 469 121 470
rect 119 469 120 470
rect 118 469 119 470
rect 117 469 118 470
rect 116 469 117 470
rect 115 469 116 470
rect 114 469 115 470
rect 113 469 114 470
rect 112 469 113 470
rect 111 469 112 470
rect 110 469 111 470
rect 109 469 110 470
rect 108 469 109 470
rect 107 469 108 470
rect 106 469 107 470
rect 105 469 106 470
rect 104 469 105 470
rect 103 469 104 470
rect 102 469 103 470
rect 101 469 102 470
rect 100 469 101 470
rect 194 470 195 471
rect 193 470 194 471
rect 192 470 193 471
rect 191 470 192 471
rect 190 470 191 471
rect 189 470 190 471
rect 181 470 182 471
rect 180 470 181 471
rect 179 470 180 471
rect 178 470 179 471
rect 176 470 177 471
rect 175 470 176 471
rect 174 470 175 471
rect 173 470 174 471
rect 172 470 173 471
rect 171 470 172 471
rect 170 470 171 471
rect 169 470 170 471
rect 168 470 169 471
rect 167 470 168 471
rect 166 470 167 471
rect 165 470 166 471
rect 164 470 165 471
rect 163 470 164 471
rect 162 470 163 471
rect 161 470 162 471
rect 160 470 161 471
rect 147 470 148 471
rect 146 470 147 471
rect 145 470 146 471
rect 144 470 145 471
rect 143 470 144 471
rect 142 470 143 471
rect 141 470 142 471
rect 140 470 141 471
rect 139 470 140 471
rect 138 470 139 471
rect 137 470 138 471
rect 136 470 137 471
rect 135 470 136 471
rect 134 470 135 471
rect 133 470 134 471
rect 132 470 133 471
rect 131 470 132 471
rect 130 470 131 471
rect 129 470 130 471
rect 128 470 129 471
rect 127 470 128 471
rect 126 470 127 471
rect 125 470 126 471
rect 124 470 125 471
rect 123 470 124 471
rect 122 470 123 471
rect 121 470 122 471
rect 120 470 121 471
rect 119 470 120 471
rect 118 470 119 471
rect 117 470 118 471
rect 116 470 117 471
rect 115 470 116 471
rect 114 470 115 471
rect 113 470 114 471
rect 112 470 113 471
rect 111 470 112 471
rect 110 470 111 471
rect 109 470 110 471
rect 108 470 109 471
rect 107 470 108 471
rect 106 470 107 471
rect 105 470 106 471
rect 104 470 105 471
rect 103 470 104 471
rect 102 470 103 471
rect 101 470 102 471
rect 100 470 101 471
rect 195 471 196 472
rect 194 471 195 472
rect 192 471 193 472
rect 190 471 191 472
rect 189 471 190 472
rect 181 471 182 472
rect 180 471 181 472
rect 179 471 180 472
rect 178 471 179 472
rect 176 471 177 472
rect 175 471 176 472
rect 174 471 175 472
rect 173 471 174 472
rect 172 471 173 472
rect 171 471 172 472
rect 170 471 171 472
rect 169 471 170 472
rect 168 471 169 472
rect 167 471 168 472
rect 166 471 167 472
rect 165 471 166 472
rect 164 471 165 472
rect 163 471 164 472
rect 162 471 163 472
rect 161 471 162 472
rect 160 471 161 472
rect 147 471 148 472
rect 146 471 147 472
rect 145 471 146 472
rect 144 471 145 472
rect 143 471 144 472
rect 142 471 143 472
rect 141 471 142 472
rect 140 471 141 472
rect 139 471 140 472
rect 138 471 139 472
rect 137 471 138 472
rect 136 471 137 472
rect 135 471 136 472
rect 134 471 135 472
rect 133 471 134 472
rect 132 471 133 472
rect 131 471 132 472
rect 130 471 131 472
rect 129 471 130 472
rect 128 471 129 472
rect 127 471 128 472
rect 126 471 127 472
rect 125 471 126 472
rect 124 471 125 472
rect 123 471 124 472
rect 122 471 123 472
rect 121 471 122 472
rect 120 471 121 472
rect 119 471 120 472
rect 118 471 119 472
rect 117 471 118 472
rect 116 471 117 472
rect 115 471 116 472
rect 114 471 115 472
rect 113 471 114 472
rect 112 471 113 472
rect 111 471 112 472
rect 110 471 111 472
rect 109 471 110 472
rect 108 471 109 472
rect 107 471 108 472
rect 106 471 107 472
rect 105 471 106 472
rect 104 471 105 472
rect 103 471 104 472
rect 102 471 103 472
rect 101 471 102 472
rect 100 471 101 472
rect 195 472 196 473
rect 194 472 195 473
rect 192 472 193 473
rect 191 472 192 473
rect 190 472 191 473
rect 189 472 190 473
rect 181 472 182 473
rect 180 472 181 473
rect 179 472 180 473
rect 178 472 179 473
rect 176 472 177 473
rect 175 472 176 473
rect 174 472 175 473
rect 173 472 174 473
rect 172 472 173 473
rect 171 472 172 473
rect 170 472 171 473
rect 169 472 170 473
rect 168 472 169 473
rect 167 472 168 473
rect 166 472 167 473
rect 165 472 166 473
rect 164 472 165 473
rect 163 472 164 473
rect 162 472 163 473
rect 161 472 162 473
rect 160 472 161 473
rect 147 472 148 473
rect 146 472 147 473
rect 145 472 146 473
rect 144 472 145 473
rect 143 472 144 473
rect 142 472 143 473
rect 141 472 142 473
rect 140 472 141 473
rect 139 472 140 473
rect 138 472 139 473
rect 137 472 138 473
rect 136 472 137 473
rect 135 472 136 473
rect 134 472 135 473
rect 133 472 134 473
rect 132 472 133 473
rect 131 472 132 473
rect 130 472 131 473
rect 129 472 130 473
rect 128 472 129 473
rect 127 472 128 473
rect 126 472 127 473
rect 125 472 126 473
rect 124 472 125 473
rect 123 472 124 473
rect 122 472 123 473
rect 121 472 122 473
rect 120 472 121 473
rect 119 472 120 473
rect 118 472 119 473
rect 117 472 118 473
rect 116 472 117 473
rect 115 472 116 473
rect 114 472 115 473
rect 113 472 114 473
rect 112 472 113 473
rect 111 472 112 473
rect 110 472 111 473
rect 109 472 110 473
rect 108 472 109 473
rect 107 472 108 473
rect 106 472 107 473
rect 105 472 106 473
rect 104 472 105 473
rect 103 472 104 473
rect 102 472 103 473
rect 101 472 102 473
rect 100 472 101 473
rect 194 473 195 474
rect 192 473 193 474
rect 191 473 192 474
rect 190 473 191 474
rect 189 473 190 474
rect 180 473 181 474
rect 179 473 180 474
rect 178 473 179 474
rect 175 473 176 474
rect 174 473 175 474
rect 173 473 174 474
rect 172 473 173 474
rect 171 473 172 474
rect 170 473 171 474
rect 169 473 170 474
rect 168 473 169 474
rect 167 473 168 474
rect 166 473 167 474
rect 165 473 166 474
rect 164 473 165 474
rect 163 473 164 474
rect 162 473 163 474
rect 161 473 162 474
rect 160 473 161 474
rect 147 473 148 474
rect 146 473 147 474
rect 145 473 146 474
rect 144 473 145 474
rect 143 473 144 474
rect 142 473 143 474
rect 141 473 142 474
rect 140 473 141 474
rect 139 473 140 474
rect 138 473 139 474
rect 137 473 138 474
rect 136 473 137 474
rect 135 473 136 474
rect 134 473 135 474
rect 133 473 134 474
rect 132 473 133 474
rect 131 473 132 474
rect 130 473 131 474
rect 129 473 130 474
rect 128 473 129 474
rect 127 473 128 474
rect 126 473 127 474
rect 125 473 126 474
rect 124 473 125 474
rect 123 473 124 474
rect 122 473 123 474
rect 121 473 122 474
rect 120 473 121 474
rect 119 473 120 474
rect 118 473 119 474
rect 117 473 118 474
rect 116 473 117 474
rect 115 473 116 474
rect 114 473 115 474
rect 113 473 114 474
rect 112 473 113 474
rect 111 473 112 474
rect 110 473 111 474
rect 109 473 110 474
rect 108 473 109 474
rect 107 473 108 474
rect 106 473 107 474
rect 105 473 106 474
rect 104 473 105 474
rect 103 473 104 474
rect 102 473 103 474
rect 101 473 102 474
rect 100 473 101 474
rect 192 474 193 475
rect 147 474 148 475
rect 146 474 147 475
rect 145 474 146 475
rect 144 474 145 475
rect 143 474 144 475
rect 142 474 143 475
rect 141 474 142 475
rect 140 474 141 475
rect 139 474 140 475
rect 138 474 139 475
rect 137 474 138 475
rect 136 474 137 475
rect 135 474 136 475
rect 134 474 135 475
rect 133 474 134 475
rect 132 474 133 475
rect 131 474 132 475
rect 130 474 131 475
rect 129 474 130 475
rect 128 474 129 475
rect 127 474 128 475
rect 126 474 127 475
rect 125 474 126 475
rect 124 474 125 475
rect 123 474 124 475
rect 122 474 123 475
rect 121 474 122 475
rect 120 474 121 475
rect 119 474 120 475
rect 118 474 119 475
rect 117 474 118 475
rect 116 474 117 475
rect 115 474 116 475
rect 114 474 115 475
rect 113 474 114 475
rect 112 474 113 475
rect 111 474 112 475
rect 110 474 111 475
rect 109 474 110 475
rect 108 474 109 475
rect 107 474 108 475
rect 106 474 107 475
rect 105 474 106 475
rect 104 474 105 475
rect 103 474 104 475
rect 102 474 103 475
rect 101 474 102 475
rect 100 474 101 475
<< metal2 >>
rect 180 7 181 8
rect 163 7 164 8
rect 180 8 181 9
rect 179 8 180 9
rect 164 8 165 9
rect 163 8 164 9
rect 180 9 181 10
rect 179 9 180 10
rect 178 9 179 10
rect 177 9 178 10
rect 176 9 177 10
rect 175 9 176 10
rect 174 9 175 10
rect 173 9 174 10
rect 172 9 173 10
rect 171 9 172 10
rect 170 9 171 10
rect 169 9 170 10
rect 168 9 169 10
rect 167 9 168 10
rect 166 9 167 10
rect 165 9 166 10
rect 164 9 165 10
rect 163 9 164 10
rect 180 10 181 11
rect 179 10 180 11
rect 178 10 179 11
rect 177 10 178 11
rect 176 10 177 11
rect 175 10 176 11
rect 174 10 175 11
rect 173 10 174 11
rect 172 10 173 11
rect 171 10 172 11
rect 170 10 171 11
rect 169 10 170 11
rect 168 10 169 11
rect 167 10 168 11
rect 166 10 167 11
rect 165 10 166 11
rect 164 10 165 11
rect 163 10 164 11
rect 180 11 181 12
rect 179 11 180 12
rect 178 11 179 12
rect 177 11 178 12
rect 176 11 177 12
rect 175 11 176 12
rect 174 11 175 12
rect 173 11 174 12
rect 172 11 173 12
rect 171 11 172 12
rect 170 11 171 12
rect 169 11 170 12
rect 168 11 169 12
rect 167 11 168 12
rect 166 11 167 12
rect 165 11 166 12
rect 164 11 165 12
rect 163 11 164 12
rect 180 12 181 13
rect 179 12 180 13
rect 178 12 179 13
rect 177 12 178 13
rect 176 12 177 13
rect 175 12 176 13
rect 174 12 175 13
rect 173 12 174 13
rect 172 12 173 13
rect 171 12 172 13
rect 170 12 171 13
rect 169 12 170 13
rect 168 12 169 13
rect 167 12 168 13
rect 166 12 167 13
rect 165 12 166 13
rect 164 12 165 13
rect 163 12 164 13
rect 180 13 181 14
rect 179 13 180 14
rect 172 13 173 14
rect 171 13 172 14
rect 164 13 165 14
rect 163 13 164 14
rect 180 14 181 15
rect 173 14 174 15
rect 172 14 173 15
rect 171 14 172 15
rect 170 14 171 15
rect 163 14 164 15
rect 175 15 176 16
rect 174 15 175 16
rect 173 15 174 16
rect 172 15 173 16
rect 171 15 172 16
rect 170 15 171 16
rect 169 15 170 16
rect 176 16 177 17
rect 175 16 176 17
rect 174 16 175 17
rect 173 16 174 17
rect 172 16 173 17
rect 171 16 172 17
rect 170 16 171 17
rect 169 16 170 17
rect 168 16 169 17
rect 178 17 179 18
rect 177 17 178 18
rect 176 17 177 18
rect 175 17 176 18
rect 174 17 175 18
rect 173 17 174 18
rect 172 17 173 18
rect 171 17 172 18
rect 168 17 169 18
rect 167 17 168 18
rect 163 17 164 18
rect 179 18 180 19
rect 178 18 179 19
rect 177 18 178 19
rect 176 18 177 19
rect 175 18 176 19
rect 174 18 175 19
rect 173 18 174 19
rect 167 18 168 19
rect 166 18 167 19
rect 165 18 166 19
rect 163 18 164 19
rect 180 19 181 20
rect 179 19 180 20
rect 178 19 179 20
rect 177 19 178 20
rect 176 19 177 20
rect 175 19 176 20
rect 174 19 175 20
rect 166 19 167 20
rect 165 19 166 20
rect 164 19 165 20
rect 163 19 164 20
rect 180 20 181 21
rect 179 20 180 21
rect 178 20 179 21
rect 177 20 178 21
rect 176 20 177 21
rect 165 20 166 21
rect 164 20 165 21
rect 163 20 164 21
rect 180 21 181 22
rect 179 21 180 22
rect 178 21 179 22
rect 177 21 178 22
rect 164 21 165 22
rect 163 21 164 22
rect 180 22 181 23
rect 179 22 180 23
rect 178 22 179 23
rect 164 22 165 23
rect 163 22 164 23
rect 180 23 181 24
rect 179 23 180 24
rect 163 23 164 24
rect 180 24 181 25
rect 163 24 164 25
rect 41 25 42 26
rect 40 25 41 26
rect 43 26 44 27
rect 42 26 43 27
rect 41 26 42 27
rect 40 26 41 27
rect 39 26 40 27
rect 38 26 39 27
rect 163 27 164 28
rect 43 27 44 28
rect 42 27 43 28
rect 41 27 42 28
rect 40 27 41 28
rect 39 27 40 28
rect 38 27 39 28
rect 37 27 38 28
rect 164 28 165 29
rect 163 28 164 29
rect 48 28 49 29
rect 47 28 48 29
rect 43 28 44 29
rect 42 28 43 29
rect 41 28 42 29
rect 40 28 41 29
rect 39 28 40 29
rect 38 28 39 29
rect 37 28 38 29
rect 36 28 37 29
rect 165 29 166 30
rect 164 29 165 30
rect 163 29 164 30
rect 50 29 51 30
rect 49 29 50 30
rect 48 29 49 30
rect 47 29 48 30
rect 46 29 47 30
rect 43 29 44 30
rect 42 29 43 30
rect 41 29 42 30
rect 40 29 41 30
rect 39 29 40 30
rect 38 29 39 30
rect 37 29 38 30
rect 36 29 37 30
rect 167 30 168 31
rect 166 30 167 31
rect 165 30 166 31
rect 164 30 165 31
rect 163 30 164 31
rect 52 30 53 31
rect 51 30 52 31
rect 50 30 51 31
rect 49 30 50 31
rect 48 30 49 31
rect 47 30 48 31
rect 46 30 47 31
rect 45 30 46 31
rect 42 30 43 31
rect 41 30 42 31
rect 40 30 41 31
rect 39 30 40 31
rect 38 30 39 31
rect 37 30 38 31
rect 36 30 37 31
rect 35 30 36 31
rect 180 31 181 32
rect 169 31 170 32
rect 168 31 169 32
rect 167 31 168 32
rect 166 31 167 32
rect 165 31 166 32
rect 164 31 165 32
rect 163 31 164 32
rect 53 31 54 32
rect 52 31 53 32
rect 51 31 52 32
rect 50 31 51 32
rect 49 31 50 32
rect 48 31 49 32
rect 47 31 48 32
rect 46 31 47 32
rect 45 31 46 32
rect 44 31 45 32
rect 42 31 43 32
rect 41 31 42 32
rect 40 31 41 32
rect 39 31 40 32
rect 38 31 39 32
rect 37 31 38 32
rect 36 31 37 32
rect 35 31 36 32
rect 180 32 181 33
rect 171 32 172 33
rect 170 32 171 33
rect 169 32 170 33
rect 168 32 169 33
rect 167 32 168 33
rect 166 32 167 33
rect 165 32 166 33
rect 164 32 165 33
rect 163 32 164 33
rect 54 32 55 33
rect 53 32 54 33
rect 52 32 53 33
rect 51 32 52 33
rect 50 32 51 33
rect 49 32 50 33
rect 48 32 49 33
rect 47 32 48 33
rect 46 32 47 33
rect 45 32 46 33
rect 44 32 45 33
rect 43 32 44 33
rect 41 32 42 33
rect 40 32 41 33
rect 39 32 40 33
rect 38 32 39 33
rect 37 32 38 33
rect 36 32 37 33
rect 35 32 36 33
rect 34 32 35 33
rect 180 33 181 34
rect 179 33 180 34
rect 178 33 179 34
rect 177 33 178 34
rect 176 33 177 34
rect 175 33 176 34
rect 174 33 175 34
rect 173 33 174 34
rect 172 33 173 34
rect 171 33 172 34
rect 170 33 171 34
rect 169 33 170 34
rect 168 33 169 34
rect 167 33 168 34
rect 166 33 167 34
rect 165 33 166 34
rect 164 33 165 34
rect 163 33 164 34
rect 54 33 55 34
rect 53 33 54 34
rect 52 33 53 34
rect 51 33 52 34
rect 50 33 51 34
rect 49 33 50 34
rect 48 33 49 34
rect 47 33 48 34
rect 46 33 47 34
rect 45 33 46 34
rect 44 33 45 34
rect 43 33 44 34
rect 42 33 43 34
rect 41 33 42 34
rect 40 33 41 34
rect 39 33 40 34
rect 38 33 39 34
rect 37 33 38 34
rect 36 33 37 34
rect 35 33 36 34
rect 34 33 35 34
rect 180 34 181 35
rect 179 34 180 35
rect 178 34 179 35
rect 177 34 178 35
rect 176 34 177 35
rect 175 34 176 35
rect 174 34 175 35
rect 173 34 174 35
rect 172 34 173 35
rect 171 34 172 35
rect 170 34 171 35
rect 169 34 170 35
rect 168 34 169 35
rect 167 34 168 35
rect 163 34 164 35
rect 61 34 62 35
rect 60 34 61 35
rect 59 34 60 35
rect 58 34 59 35
rect 55 34 56 35
rect 54 34 55 35
rect 53 34 54 35
rect 52 34 53 35
rect 51 34 52 35
rect 50 34 51 35
rect 49 34 50 35
rect 48 34 49 35
rect 47 34 48 35
rect 46 34 47 35
rect 45 34 46 35
rect 44 34 45 35
rect 43 34 44 35
rect 42 34 43 35
rect 41 34 42 35
rect 40 34 41 35
rect 39 34 40 35
rect 38 34 39 35
rect 37 34 38 35
rect 36 34 37 35
rect 35 34 36 35
rect 34 34 35 35
rect 33 34 34 35
rect 180 35 181 36
rect 179 35 180 36
rect 178 35 179 36
rect 177 35 178 36
rect 176 35 177 36
rect 175 35 176 36
rect 174 35 175 36
rect 173 35 174 36
rect 172 35 173 36
rect 171 35 172 36
rect 170 35 171 36
rect 169 35 170 36
rect 63 35 64 36
rect 62 35 63 36
rect 61 35 62 36
rect 60 35 61 36
rect 59 35 60 36
rect 58 35 59 36
rect 55 35 56 36
rect 54 35 55 36
rect 53 35 54 36
rect 52 35 53 36
rect 51 35 52 36
rect 50 35 51 36
rect 49 35 50 36
rect 48 35 49 36
rect 47 35 48 36
rect 46 35 47 36
rect 45 35 46 36
rect 44 35 45 36
rect 43 35 44 36
rect 42 35 43 36
rect 41 35 42 36
rect 40 35 41 36
rect 39 35 40 36
rect 38 35 39 36
rect 37 35 38 36
rect 36 35 37 36
rect 35 35 36 36
rect 34 35 35 36
rect 33 35 34 36
rect 180 36 181 37
rect 179 36 180 37
rect 178 36 179 37
rect 177 36 178 37
rect 176 36 177 37
rect 175 36 176 37
rect 174 36 175 37
rect 173 36 174 37
rect 172 36 173 37
rect 171 36 172 37
rect 65 36 66 37
rect 64 36 65 37
rect 63 36 64 37
rect 62 36 63 37
rect 61 36 62 37
rect 60 36 61 37
rect 59 36 60 37
rect 58 36 59 37
rect 55 36 56 37
rect 54 36 55 37
rect 53 36 54 37
rect 52 36 53 37
rect 51 36 52 37
rect 50 36 51 37
rect 49 36 50 37
rect 48 36 49 37
rect 47 36 48 37
rect 46 36 47 37
rect 45 36 46 37
rect 44 36 45 37
rect 43 36 44 37
rect 42 36 43 37
rect 41 36 42 37
rect 40 36 41 37
rect 39 36 40 37
rect 38 36 39 37
rect 37 36 38 37
rect 36 36 37 37
rect 35 36 36 37
rect 34 36 35 37
rect 33 36 34 37
rect 32 36 33 37
rect 180 37 181 38
rect 179 37 180 38
rect 178 37 179 38
rect 177 37 178 38
rect 176 37 177 38
rect 175 37 176 38
rect 174 37 175 38
rect 173 37 174 38
rect 172 37 173 38
rect 171 37 172 38
rect 170 37 171 38
rect 169 37 170 38
rect 67 37 68 38
rect 66 37 67 38
rect 65 37 66 38
rect 64 37 65 38
rect 63 37 64 38
rect 62 37 63 38
rect 61 37 62 38
rect 60 37 61 38
rect 59 37 60 38
rect 58 37 59 38
rect 55 37 56 38
rect 54 37 55 38
rect 53 37 54 38
rect 52 37 53 38
rect 51 37 52 38
rect 50 37 51 38
rect 49 37 50 38
rect 48 37 49 38
rect 47 37 48 38
rect 46 37 47 38
rect 45 37 46 38
rect 44 37 45 38
rect 43 37 44 38
rect 42 37 43 38
rect 41 37 42 38
rect 40 37 41 38
rect 39 37 40 38
rect 38 37 39 38
rect 37 37 38 38
rect 36 37 37 38
rect 35 37 36 38
rect 34 37 35 38
rect 33 37 34 38
rect 32 37 33 38
rect 180 38 181 39
rect 170 38 171 39
rect 169 38 170 39
rect 168 38 169 39
rect 167 38 168 39
rect 163 38 164 39
rect 69 38 70 39
rect 68 38 69 39
rect 67 38 68 39
rect 66 38 67 39
rect 65 38 66 39
rect 64 38 65 39
rect 63 38 64 39
rect 62 38 63 39
rect 61 38 62 39
rect 60 38 61 39
rect 59 38 60 39
rect 58 38 59 39
rect 55 38 56 39
rect 54 38 55 39
rect 53 38 54 39
rect 52 38 53 39
rect 51 38 52 39
rect 50 38 51 39
rect 49 38 50 39
rect 48 38 49 39
rect 47 38 48 39
rect 46 38 47 39
rect 45 38 46 39
rect 44 38 45 39
rect 43 38 44 39
rect 42 38 43 39
rect 41 38 42 39
rect 40 38 41 39
rect 39 38 40 39
rect 38 38 39 39
rect 37 38 38 39
rect 36 38 37 39
rect 35 38 36 39
rect 34 38 35 39
rect 33 38 34 39
rect 32 38 33 39
rect 31 38 32 39
rect 195 39 196 40
rect 194 39 195 40
rect 193 39 194 40
rect 192 39 193 40
rect 191 39 192 40
rect 190 39 191 40
rect 189 39 190 40
rect 180 39 181 40
rect 168 39 169 40
rect 167 39 168 40
rect 166 39 167 40
rect 165 39 166 40
rect 164 39 165 40
rect 163 39 164 40
rect 97 39 98 40
rect 96 39 97 40
rect 95 39 96 40
rect 94 39 95 40
rect 93 39 94 40
rect 92 39 93 40
rect 91 39 92 40
rect 90 39 91 40
rect 89 39 90 40
rect 88 39 89 40
rect 87 39 88 40
rect 70 39 71 40
rect 69 39 70 40
rect 68 39 69 40
rect 67 39 68 40
rect 66 39 67 40
rect 65 39 66 40
rect 64 39 65 40
rect 63 39 64 40
rect 62 39 63 40
rect 61 39 62 40
rect 60 39 61 40
rect 59 39 60 40
rect 58 39 59 40
rect 57 39 58 40
rect 54 39 55 40
rect 53 39 54 40
rect 52 39 53 40
rect 51 39 52 40
rect 50 39 51 40
rect 49 39 50 40
rect 48 39 49 40
rect 47 39 48 40
rect 46 39 47 40
rect 45 39 46 40
rect 44 39 45 40
rect 43 39 44 40
rect 42 39 43 40
rect 41 39 42 40
rect 40 39 41 40
rect 39 39 40 40
rect 38 39 39 40
rect 37 39 38 40
rect 36 39 37 40
rect 35 39 36 40
rect 34 39 35 40
rect 33 39 34 40
rect 32 39 33 40
rect 31 39 32 40
rect 30 39 31 40
rect 196 40 197 41
rect 195 40 196 41
rect 194 40 195 41
rect 193 40 194 41
rect 192 40 193 41
rect 191 40 192 41
rect 190 40 191 41
rect 189 40 190 41
rect 166 40 167 41
rect 165 40 166 41
rect 164 40 165 41
rect 163 40 164 41
rect 101 40 102 41
rect 100 40 101 41
rect 99 40 100 41
rect 98 40 99 41
rect 97 40 98 41
rect 96 40 97 41
rect 95 40 96 41
rect 94 40 95 41
rect 93 40 94 41
rect 92 40 93 41
rect 91 40 92 41
rect 90 40 91 41
rect 89 40 90 41
rect 88 40 89 41
rect 87 40 88 41
rect 86 40 87 41
rect 85 40 86 41
rect 84 40 85 41
rect 70 40 71 41
rect 69 40 70 41
rect 68 40 69 41
rect 67 40 68 41
rect 66 40 67 41
rect 65 40 66 41
rect 64 40 65 41
rect 63 40 64 41
rect 62 40 63 41
rect 61 40 62 41
rect 60 40 61 41
rect 59 40 60 41
rect 58 40 59 41
rect 57 40 58 41
rect 54 40 55 41
rect 53 40 54 41
rect 52 40 53 41
rect 51 40 52 41
rect 50 40 51 41
rect 49 40 50 41
rect 48 40 49 41
rect 47 40 48 41
rect 46 40 47 41
rect 45 40 46 41
rect 44 40 45 41
rect 43 40 44 41
rect 42 40 43 41
rect 41 40 42 41
rect 40 40 41 41
rect 39 40 40 41
rect 38 40 39 41
rect 37 40 38 41
rect 36 40 37 41
rect 35 40 36 41
rect 34 40 35 41
rect 33 40 34 41
rect 32 40 33 41
rect 31 40 32 41
rect 30 40 31 41
rect 197 41 198 42
rect 196 41 197 42
rect 195 41 196 42
rect 189 41 190 42
rect 165 41 166 42
rect 164 41 165 42
rect 163 41 164 42
rect 103 41 104 42
rect 102 41 103 42
rect 101 41 102 42
rect 100 41 101 42
rect 99 41 100 42
rect 98 41 99 42
rect 97 41 98 42
rect 96 41 97 42
rect 95 41 96 42
rect 94 41 95 42
rect 93 41 94 42
rect 92 41 93 42
rect 91 41 92 42
rect 90 41 91 42
rect 89 41 90 42
rect 88 41 89 42
rect 87 41 88 42
rect 86 41 87 42
rect 85 41 86 42
rect 84 41 85 42
rect 83 41 84 42
rect 82 41 83 42
rect 70 41 71 42
rect 69 41 70 42
rect 68 41 69 42
rect 67 41 68 42
rect 66 41 67 42
rect 65 41 66 42
rect 64 41 65 42
rect 63 41 64 42
rect 62 41 63 42
rect 61 41 62 42
rect 60 41 61 42
rect 59 41 60 42
rect 58 41 59 42
rect 57 41 58 42
rect 54 41 55 42
rect 53 41 54 42
rect 52 41 53 42
rect 51 41 52 42
rect 50 41 51 42
rect 49 41 50 42
rect 48 41 49 42
rect 47 41 48 42
rect 46 41 47 42
rect 45 41 46 42
rect 44 41 45 42
rect 43 41 44 42
rect 42 41 43 42
rect 41 41 42 42
rect 40 41 41 42
rect 39 41 40 42
rect 38 41 39 42
rect 37 41 38 42
rect 36 41 37 42
rect 35 41 36 42
rect 34 41 35 42
rect 33 41 34 42
rect 32 41 33 42
rect 31 41 32 42
rect 30 41 31 42
rect 29 41 30 42
rect 197 42 198 43
rect 196 42 197 43
rect 164 42 165 43
rect 163 42 164 43
rect 105 42 106 43
rect 104 42 105 43
rect 103 42 104 43
rect 102 42 103 43
rect 101 42 102 43
rect 100 42 101 43
rect 99 42 100 43
rect 98 42 99 43
rect 97 42 98 43
rect 96 42 97 43
rect 95 42 96 43
rect 94 42 95 43
rect 93 42 94 43
rect 92 42 93 43
rect 91 42 92 43
rect 90 42 91 43
rect 89 42 90 43
rect 88 42 89 43
rect 87 42 88 43
rect 86 42 87 43
rect 85 42 86 43
rect 84 42 85 43
rect 83 42 84 43
rect 82 42 83 43
rect 81 42 82 43
rect 80 42 81 43
rect 69 42 70 43
rect 68 42 69 43
rect 67 42 68 43
rect 66 42 67 43
rect 65 42 66 43
rect 64 42 65 43
rect 63 42 64 43
rect 62 42 63 43
rect 61 42 62 43
rect 60 42 61 43
rect 59 42 60 43
rect 58 42 59 43
rect 57 42 58 43
rect 54 42 55 43
rect 53 42 54 43
rect 52 42 53 43
rect 51 42 52 43
rect 50 42 51 43
rect 49 42 50 43
rect 48 42 49 43
rect 47 42 48 43
rect 46 42 47 43
rect 45 42 46 43
rect 44 42 45 43
rect 43 42 44 43
rect 42 42 43 43
rect 41 42 42 43
rect 40 42 41 43
rect 39 42 40 43
rect 38 42 39 43
rect 37 42 38 43
rect 36 42 37 43
rect 35 42 36 43
rect 34 42 35 43
rect 33 42 34 43
rect 32 42 33 43
rect 31 42 32 43
rect 30 42 31 43
rect 29 42 30 43
rect 28 42 29 43
rect 197 43 198 44
rect 163 43 164 44
rect 107 43 108 44
rect 106 43 107 44
rect 105 43 106 44
rect 104 43 105 44
rect 103 43 104 44
rect 102 43 103 44
rect 101 43 102 44
rect 100 43 101 44
rect 99 43 100 44
rect 98 43 99 44
rect 97 43 98 44
rect 96 43 97 44
rect 95 43 96 44
rect 94 43 95 44
rect 93 43 94 44
rect 92 43 93 44
rect 91 43 92 44
rect 90 43 91 44
rect 89 43 90 44
rect 88 43 89 44
rect 87 43 88 44
rect 86 43 87 44
rect 85 43 86 44
rect 84 43 85 44
rect 83 43 84 44
rect 82 43 83 44
rect 81 43 82 44
rect 80 43 81 44
rect 79 43 80 44
rect 69 43 70 44
rect 68 43 69 44
rect 67 43 68 44
rect 66 43 67 44
rect 65 43 66 44
rect 64 43 65 44
rect 63 43 64 44
rect 62 43 63 44
rect 61 43 62 44
rect 60 43 61 44
rect 59 43 60 44
rect 58 43 59 44
rect 57 43 58 44
rect 54 43 55 44
rect 53 43 54 44
rect 52 43 53 44
rect 51 43 52 44
rect 50 43 51 44
rect 49 43 50 44
rect 48 43 49 44
rect 47 43 48 44
rect 46 43 47 44
rect 45 43 46 44
rect 44 43 45 44
rect 43 43 44 44
rect 42 43 43 44
rect 41 43 42 44
rect 40 43 41 44
rect 39 43 40 44
rect 38 43 39 44
rect 37 43 38 44
rect 36 43 37 44
rect 35 43 36 44
rect 34 43 35 44
rect 33 43 34 44
rect 32 43 33 44
rect 31 43 32 44
rect 30 43 31 44
rect 29 43 30 44
rect 28 43 29 44
rect 197 44 198 45
rect 196 44 197 45
rect 109 44 110 45
rect 108 44 109 45
rect 107 44 108 45
rect 106 44 107 45
rect 105 44 106 45
rect 104 44 105 45
rect 103 44 104 45
rect 102 44 103 45
rect 101 44 102 45
rect 100 44 101 45
rect 99 44 100 45
rect 98 44 99 45
rect 97 44 98 45
rect 96 44 97 45
rect 95 44 96 45
rect 94 44 95 45
rect 93 44 94 45
rect 92 44 93 45
rect 91 44 92 45
rect 90 44 91 45
rect 89 44 90 45
rect 88 44 89 45
rect 87 44 88 45
rect 86 44 87 45
rect 85 44 86 45
rect 84 44 85 45
rect 83 44 84 45
rect 82 44 83 45
rect 81 44 82 45
rect 80 44 81 45
rect 79 44 80 45
rect 78 44 79 45
rect 69 44 70 45
rect 68 44 69 45
rect 67 44 68 45
rect 66 44 67 45
rect 65 44 66 45
rect 64 44 65 45
rect 63 44 64 45
rect 62 44 63 45
rect 61 44 62 45
rect 60 44 61 45
rect 59 44 60 45
rect 58 44 59 45
rect 57 44 58 45
rect 53 44 54 45
rect 52 44 53 45
rect 51 44 52 45
rect 50 44 51 45
rect 49 44 50 45
rect 48 44 49 45
rect 47 44 48 45
rect 46 44 47 45
rect 45 44 46 45
rect 44 44 45 45
rect 43 44 44 45
rect 42 44 43 45
rect 41 44 42 45
rect 40 44 41 45
rect 39 44 40 45
rect 38 44 39 45
rect 37 44 38 45
rect 36 44 37 45
rect 35 44 36 45
rect 34 44 35 45
rect 33 44 34 45
rect 32 44 33 45
rect 31 44 32 45
rect 30 44 31 45
rect 29 44 30 45
rect 28 44 29 45
rect 27 44 28 45
rect 196 45 197 46
rect 195 45 196 46
rect 194 45 195 46
rect 193 45 194 46
rect 192 45 193 46
rect 191 45 192 46
rect 190 45 191 46
rect 189 45 190 46
rect 110 45 111 46
rect 109 45 110 46
rect 108 45 109 46
rect 107 45 108 46
rect 106 45 107 46
rect 105 45 106 46
rect 104 45 105 46
rect 103 45 104 46
rect 102 45 103 46
rect 101 45 102 46
rect 100 45 101 46
rect 99 45 100 46
rect 98 45 99 46
rect 97 45 98 46
rect 96 45 97 46
rect 95 45 96 46
rect 94 45 95 46
rect 93 45 94 46
rect 92 45 93 46
rect 91 45 92 46
rect 90 45 91 46
rect 89 45 90 46
rect 88 45 89 46
rect 87 45 88 46
rect 86 45 87 46
rect 85 45 86 46
rect 84 45 85 46
rect 83 45 84 46
rect 82 45 83 46
rect 81 45 82 46
rect 80 45 81 46
rect 79 45 80 46
rect 78 45 79 46
rect 77 45 78 46
rect 68 45 69 46
rect 67 45 68 46
rect 66 45 67 46
rect 65 45 66 46
rect 64 45 65 46
rect 63 45 64 46
rect 62 45 63 46
rect 61 45 62 46
rect 60 45 61 46
rect 59 45 60 46
rect 58 45 59 46
rect 57 45 58 46
rect 56 45 57 46
rect 53 45 54 46
rect 52 45 53 46
rect 51 45 52 46
rect 50 45 51 46
rect 49 45 50 46
rect 48 45 49 46
rect 47 45 48 46
rect 46 45 47 46
rect 45 45 46 46
rect 44 45 45 46
rect 43 45 44 46
rect 42 45 43 46
rect 41 45 42 46
rect 40 45 41 46
rect 39 45 40 46
rect 38 45 39 46
rect 37 45 38 46
rect 36 45 37 46
rect 35 45 36 46
rect 33 45 34 46
rect 32 45 33 46
rect 31 45 32 46
rect 30 45 31 46
rect 29 45 30 46
rect 28 45 29 46
rect 27 45 28 46
rect 26 45 27 46
rect 190 46 191 47
rect 189 46 190 47
rect 163 46 164 47
rect 111 46 112 47
rect 110 46 111 47
rect 109 46 110 47
rect 108 46 109 47
rect 107 46 108 47
rect 106 46 107 47
rect 105 46 106 47
rect 104 46 105 47
rect 103 46 104 47
rect 102 46 103 47
rect 101 46 102 47
rect 100 46 101 47
rect 99 46 100 47
rect 98 46 99 47
rect 97 46 98 47
rect 96 46 97 47
rect 95 46 96 47
rect 94 46 95 47
rect 93 46 94 47
rect 92 46 93 47
rect 91 46 92 47
rect 90 46 91 47
rect 89 46 90 47
rect 88 46 89 47
rect 87 46 88 47
rect 86 46 87 47
rect 85 46 86 47
rect 84 46 85 47
rect 83 46 84 47
rect 82 46 83 47
rect 81 46 82 47
rect 80 46 81 47
rect 79 46 80 47
rect 78 46 79 47
rect 77 46 78 47
rect 76 46 77 47
rect 68 46 69 47
rect 67 46 68 47
rect 66 46 67 47
rect 65 46 66 47
rect 64 46 65 47
rect 63 46 64 47
rect 62 46 63 47
rect 61 46 62 47
rect 60 46 61 47
rect 59 46 60 47
rect 58 46 59 47
rect 57 46 58 47
rect 56 46 57 47
rect 52 46 53 47
rect 51 46 52 47
rect 50 46 51 47
rect 49 46 50 47
rect 48 46 49 47
rect 47 46 48 47
rect 46 46 47 47
rect 45 46 46 47
rect 44 46 45 47
rect 43 46 44 47
rect 42 46 43 47
rect 41 46 42 47
rect 40 46 41 47
rect 39 46 40 47
rect 38 46 39 47
rect 37 46 38 47
rect 36 46 37 47
rect 35 46 36 47
rect 32 46 33 47
rect 31 46 32 47
rect 30 46 31 47
rect 29 46 30 47
rect 28 46 29 47
rect 27 46 28 47
rect 26 46 27 47
rect 25 46 26 47
rect 163 47 164 48
rect 112 47 113 48
rect 111 47 112 48
rect 110 47 111 48
rect 109 47 110 48
rect 108 47 109 48
rect 107 47 108 48
rect 106 47 107 48
rect 105 47 106 48
rect 104 47 105 48
rect 103 47 104 48
rect 102 47 103 48
rect 101 47 102 48
rect 100 47 101 48
rect 99 47 100 48
rect 98 47 99 48
rect 97 47 98 48
rect 96 47 97 48
rect 95 47 96 48
rect 94 47 95 48
rect 93 47 94 48
rect 92 47 93 48
rect 91 47 92 48
rect 90 47 91 48
rect 89 47 90 48
rect 88 47 89 48
rect 87 47 88 48
rect 86 47 87 48
rect 85 47 86 48
rect 84 47 85 48
rect 83 47 84 48
rect 82 47 83 48
rect 81 47 82 48
rect 80 47 81 48
rect 79 47 80 48
rect 78 47 79 48
rect 77 47 78 48
rect 76 47 77 48
rect 68 47 69 48
rect 67 47 68 48
rect 66 47 67 48
rect 65 47 66 48
rect 64 47 65 48
rect 63 47 64 48
rect 62 47 63 48
rect 61 47 62 48
rect 60 47 61 48
rect 59 47 60 48
rect 58 47 59 48
rect 57 47 58 48
rect 56 47 57 48
rect 51 47 52 48
rect 50 47 51 48
rect 49 47 50 48
rect 48 47 49 48
rect 47 47 48 48
rect 46 47 47 48
rect 45 47 46 48
rect 44 47 45 48
rect 43 47 44 48
rect 42 47 43 48
rect 41 47 42 48
rect 40 47 41 48
rect 39 47 40 48
rect 38 47 39 48
rect 37 47 38 48
rect 36 47 37 48
rect 35 47 36 48
rect 32 47 33 48
rect 31 47 32 48
rect 30 47 31 48
rect 29 47 30 48
rect 28 47 29 48
rect 27 47 28 48
rect 26 47 27 48
rect 25 47 26 48
rect 24 47 25 48
rect 173 48 174 49
rect 172 48 173 49
rect 171 48 172 49
rect 170 48 171 49
rect 169 48 170 49
rect 168 48 169 49
rect 167 48 168 49
rect 166 48 167 49
rect 165 48 166 49
rect 164 48 165 49
rect 163 48 164 49
rect 113 48 114 49
rect 112 48 113 49
rect 111 48 112 49
rect 110 48 111 49
rect 109 48 110 49
rect 108 48 109 49
rect 107 48 108 49
rect 106 48 107 49
rect 105 48 106 49
rect 104 48 105 49
rect 103 48 104 49
rect 102 48 103 49
rect 101 48 102 49
rect 100 48 101 49
rect 99 48 100 49
rect 98 48 99 49
rect 97 48 98 49
rect 96 48 97 49
rect 95 48 96 49
rect 94 48 95 49
rect 93 48 94 49
rect 92 48 93 49
rect 91 48 92 49
rect 90 48 91 49
rect 89 48 90 49
rect 88 48 89 49
rect 87 48 88 49
rect 86 48 87 49
rect 85 48 86 49
rect 84 48 85 49
rect 83 48 84 49
rect 82 48 83 49
rect 81 48 82 49
rect 80 48 81 49
rect 79 48 80 49
rect 78 48 79 49
rect 77 48 78 49
rect 76 48 77 49
rect 75 48 76 49
rect 67 48 68 49
rect 66 48 67 49
rect 65 48 66 49
rect 64 48 65 49
rect 63 48 64 49
rect 62 48 63 49
rect 61 48 62 49
rect 60 48 61 49
rect 59 48 60 49
rect 58 48 59 49
rect 57 48 58 49
rect 56 48 57 49
rect 51 48 52 49
rect 50 48 51 49
rect 49 48 50 49
rect 48 48 49 49
rect 47 48 48 49
rect 46 48 47 49
rect 45 48 46 49
rect 44 48 45 49
rect 43 48 44 49
rect 42 48 43 49
rect 41 48 42 49
rect 40 48 41 49
rect 39 48 40 49
rect 38 48 39 49
rect 37 48 38 49
rect 36 48 37 49
rect 31 48 32 49
rect 30 48 31 49
rect 29 48 30 49
rect 28 48 29 49
rect 27 48 28 49
rect 26 48 27 49
rect 25 48 26 49
rect 24 48 25 49
rect 23 48 24 49
rect 22 48 23 49
rect 177 49 178 50
rect 176 49 177 50
rect 175 49 176 50
rect 174 49 175 50
rect 173 49 174 50
rect 172 49 173 50
rect 171 49 172 50
rect 170 49 171 50
rect 169 49 170 50
rect 168 49 169 50
rect 167 49 168 50
rect 166 49 167 50
rect 165 49 166 50
rect 164 49 165 50
rect 163 49 164 50
rect 114 49 115 50
rect 113 49 114 50
rect 112 49 113 50
rect 111 49 112 50
rect 110 49 111 50
rect 109 49 110 50
rect 108 49 109 50
rect 107 49 108 50
rect 106 49 107 50
rect 105 49 106 50
rect 104 49 105 50
rect 103 49 104 50
rect 102 49 103 50
rect 101 49 102 50
rect 100 49 101 50
rect 99 49 100 50
rect 98 49 99 50
rect 97 49 98 50
rect 96 49 97 50
rect 95 49 96 50
rect 94 49 95 50
rect 93 49 94 50
rect 92 49 93 50
rect 91 49 92 50
rect 90 49 91 50
rect 89 49 90 50
rect 88 49 89 50
rect 87 49 88 50
rect 86 49 87 50
rect 85 49 86 50
rect 84 49 85 50
rect 83 49 84 50
rect 82 49 83 50
rect 81 49 82 50
rect 80 49 81 50
rect 79 49 80 50
rect 78 49 79 50
rect 77 49 78 50
rect 76 49 77 50
rect 75 49 76 50
rect 67 49 68 50
rect 66 49 67 50
rect 65 49 66 50
rect 64 49 65 50
rect 63 49 64 50
rect 62 49 63 50
rect 61 49 62 50
rect 60 49 61 50
rect 59 49 60 50
rect 58 49 59 50
rect 57 49 58 50
rect 56 49 57 50
rect 55 49 56 50
rect 52 49 53 50
rect 51 49 52 50
rect 50 49 51 50
rect 49 49 50 50
rect 48 49 49 50
rect 47 49 48 50
rect 46 49 47 50
rect 45 49 46 50
rect 44 49 45 50
rect 43 49 44 50
rect 42 49 43 50
rect 41 49 42 50
rect 40 49 41 50
rect 39 49 40 50
rect 38 49 39 50
rect 31 49 32 50
rect 30 49 31 50
rect 29 49 30 50
rect 28 49 29 50
rect 27 49 28 50
rect 26 49 27 50
rect 25 49 26 50
rect 24 49 25 50
rect 23 49 24 50
rect 22 49 23 50
rect 21 49 22 50
rect 179 50 180 51
rect 178 50 179 51
rect 177 50 178 51
rect 176 50 177 51
rect 175 50 176 51
rect 174 50 175 51
rect 173 50 174 51
rect 172 50 173 51
rect 171 50 172 51
rect 170 50 171 51
rect 169 50 170 51
rect 168 50 169 51
rect 167 50 168 51
rect 166 50 167 51
rect 165 50 166 51
rect 164 50 165 51
rect 163 50 164 51
rect 115 50 116 51
rect 114 50 115 51
rect 113 50 114 51
rect 112 50 113 51
rect 111 50 112 51
rect 110 50 111 51
rect 109 50 110 51
rect 108 50 109 51
rect 107 50 108 51
rect 106 50 107 51
rect 105 50 106 51
rect 104 50 105 51
rect 103 50 104 51
rect 102 50 103 51
rect 101 50 102 51
rect 100 50 101 51
rect 99 50 100 51
rect 98 50 99 51
rect 97 50 98 51
rect 96 50 97 51
rect 95 50 96 51
rect 94 50 95 51
rect 93 50 94 51
rect 92 50 93 51
rect 91 50 92 51
rect 90 50 91 51
rect 89 50 90 51
rect 88 50 89 51
rect 87 50 88 51
rect 86 50 87 51
rect 85 50 86 51
rect 84 50 85 51
rect 83 50 84 51
rect 82 50 83 51
rect 81 50 82 51
rect 80 50 81 51
rect 79 50 80 51
rect 78 50 79 51
rect 77 50 78 51
rect 76 50 77 51
rect 75 50 76 51
rect 74 50 75 51
rect 67 50 68 51
rect 66 50 67 51
rect 65 50 66 51
rect 64 50 65 51
rect 63 50 64 51
rect 62 50 63 51
rect 61 50 62 51
rect 60 50 61 51
rect 59 50 60 51
rect 58 50 59 51
rect 57 50 58 51
rect 56 50 57 51
rect 55 50 56 51
rect 54 50 55 51
rect 53 50 54 51
rect 52 50 53 51
rect 51 50 52 51
rect 50 50 51 51
rect 49 50 50 51
rect 48 50 49 51
rect 47 50 48 51
rect 46 50 47 51
rect 45 50 46 51
rect 44 50 45 51
rect 43 50 44 51
rect 42 50 43 51
rect 41 50 42 51
rect 40 50 41 51
rect 39 50 40 51
rect 38 50 39 51
rect 37 50 38 51
rect 30 50 31 51
rect 29 50 30 51
rect 28 50 29 51
rect 27 50 28 51
rect 26 50 27 51
rect 25 50 26 51
rect 24 50 25 51
rect 23 50 24 51
rect 22 50 23 51
rect 21 50 22 51
rect 20 50 21 51
rect 19 50 20 51
rect 197 51 198 52
rect 196 51 197 52
rect 195 51 196 52
rect 194 51 195 52
rect 193 51 194 52
rect 192 51 193 52
rect 191 51 192 52
rect 190 51 191 52
rect 189 51 190 52
rect 180 51 181 52
rect 179 51 180 52
rect 178 51 179 52
rect 177 51 178 52
rect 176 51 177 52
rect 175 51 176 52
rect 174 51 175 52
rect 173 51 174 52
rect 172 51 173 52
rect 171 51 172 52
rect 170 51 171 52
rect 169 51 170 52
rect 168 51 169 52
rect 167 51 168 52
rect 166 51 167 52
rect 165 51 166 52
rect 164 51 165 52
rect 163 51 164 52
rect 110 51 111 52
rect 109 51 110 52
rect 108 51 109 52
rect 107 51 108 52
rect 106 51 107 52
rect 105 51 106 52
rect 104 51 105 52
rect 103 51 104 52
rect 102 51 103 52
rect 101 51 102 52
rect 100 51 101 52
rect 99 51 100 52
rect 98 51 99 52
rect 97 51 98 52
rect 96 51 97 52
rect 95 51 96 52
rect 94 51 95 52
rect 93 51 94 52
rect 92 51 93 52
rect 91 51 92 52
rect 90 51 91 52
rect 89 51 90 52
rect 88 51 89 52
rect 87 51 88 52
rect 86 51 87 52
rect 85 51 86 52
rect 84 51 85 52
rect 83 51 84 52
rect 82 51 83 52
rect 81 51 82 52
rect 80 51 81 52
rect 79 51 80 52
rect 78 51 79 52
rect 77 51 78 52
rect 76 51 77 52
rect 75 51 76 52
rect 74 51 75 52
rect 66 51 67 52
rect 65 51 66 52
rect 64 51 65 52
rect 63 51 64 52
rect 62 51 63 52
rect 61 51 62 52
rect 60 51 61 52
rect 59 51 60 52
rect 58 51 59 52
rect 57 51 58 52
rect 56 51 57 52
rect 55 51 56 52
rect 54 51 55 52
rect 53 51 54 52
rect 52 51 53 52
rect 51 51 52 52
rect 50 51 51 52
rect 49 51 50 52
rect 48 51 49 52
rect 47 51 48 52
rect 46 51 47 52
rect 45 51 46 52
rect 44 51 45 52
rect 43 51 44 52
rect 42 51 43 52
rect 41 51 42 52
rect 40 51 41 52
rect 39 51 40 52
rect 38 51 39 52
rect 37 51 38 52
rect 36 51 37 52
rect 35 51 36 52
rect 30 51 31 52
rect 29 51 30 52
rect 28 51 29 52
rect 27 51 28 52
rect 26 51 27 52
rect 25 51 26 52
rect 24 51 25 52
rect 23 51 24 52
rect 22 51 23 52
rect 21 51 22 52
rect 20 51 21 52
rect 19 51 20 52
rect 18 51 19 52
rect 197 52 198 53
rect 196 52 197 53
rect 191 52 192 53
rect 190 52 191 53
rect 189 52 190 53
rect 180 52 181 53
rect 179 52 180 53
rect 178 52 179 53
rect 177 52 178 53
rect 176 52 177 53
rect 175 52 176 53
rect 174 52 175 53
rect 173 52 174 53
rect 172 52 173 53
rect 171 52 172 53
rect 170 52 171 53
rect 169 52 170 53
rect 168 52 169 53
rect 167 52 168 53
rect 166 52 167 53
rect 165 52 166 53
rect 164 52 165 53
rect 163 52 164 53
rect 104 52 105 53
rect 103 52 104 53
rect 102 52 103 53
rect 101 52 102 53
rect 100 52 101 53
rect 99 52 100 53
rect 98 52 99 53
rect 97 52 98 53
rect 96 52 97 53
rect 95 52 96 53
rect 94 52 95 53
rect 93 52 94 53
rect 92 52 93 53
rect 91 52 92 53
rect 90 52 91 53
rect 89 52 90 53
rect 88 52 89 53
rect 87 52 88 53
rect 86 52 87 53
rect 85 52 86 53
rect 84 52 85 53
rect 83 52 84 53
rect 82 52 83 53
rect 81 52 82 53
rect 80 52 81 53
rect 79 52 80 53
rect 78 52 79 53
rect 77 52 78 53
rect 76 52 77 53
rect 75 52 76 53
rect 74 52 75 53
rect 73 52 74 53
rect 66 52 67 53
rect 65 52 66 53
rect 64 52 65 53
rect 63 52 64 53
rect 62 52 63 53
rect 61 52 62 53
rect 60 52 61 53
rect 59 52 60 53
rect 58 52 59 53
rect 57 52 58 53
rect 56 52 57 53
rect 55 52 56 53
rect 54 52 55 53
rect 53 52 54 53
rect 52 52 53 53
rect 51 52 52 53
rect 50 52 51 53
rect 49 52 50 53
rect 48 52 49 53
rect 47 52 48 53
rect 46 52 47 53
rect 45 52 46 53
rect 44 52 45 53
rect 43 52 44 53
rect 42 52 43 53
rect 41 52 42 53
rect 40 52 41 53
rect 39 52 40 53
rect 38 52 39 53
rect 37 52 38 53
rect 36 52 37 53
rect 35 52 36 53
rect 34 52 35 53
rect 30 52 31 53
rect 29 52 30 53
rect 28 52 29 53
rect 27 52 28 53
rect 26 52 27 53
rect 25 52 26 53
rect 24 52 25 53
rect 23 52 24 53
rect 22 52 23 53
rect 21 52 22 53
rect 20 52 21 53
rect 19 52 20 53
rect 18 52 19 53
rect 192 53 193 54
rect 191 53 192 54
rect 190 53 191 54
rect 189 53 190 54
rect 180 53 181 54
rect 179 53 180 54
rect 178 53 179 54
rect 177 53 178 54
rect 164 53 165 54
rect 163 53 164 54
rect 102 53 103 54
rect 101 53 102 54
rect 100 53 101 54
rect 99 53 100 54
rect 98 53 99 54
rect 97 53 98 54
rect 96 53 97 54
rect 95 53 96 54
rect 94 53 95 54
rect 93 53 94 54
rect 92 53 93 54
rect 91 53 92 54
rect 90 53 91 54
rect 89 53 90 54
rect 88 53 89 54
rect 87 53 88 54
rect 86 53 87 54
rect 85 53 86 54
rect 84 53 85 54
rect 83 53 84 54
rect 82 53 83 54
rect 81 53 82 54
rect 80 53 81 54
rect 79 53 80 54
rect 78 53 79 54
rect 77 53 78 54
rect 76 53 77 54
rect 75 53 76 54
rect 74 53 75 54
rect 73 53 74 54
rect 66 53 67 54
rect 65 53 66 54
rect 64 53 65 54
rect 63 53 64 54
rect 62 53 63 54
rect 61 53 62 54
rect 60 53 61 54
rect 59 53 60 54
rect 58 53 59 54
rect 57 53 58 54
rect 56 53 57 54
rect 55 53 56 54
rect 54 53 55 54
rect 53 53 54 54
rect 52 53 53 54
rect 51 53 52 54
rect 50 53 51 54
rect 49 53 50 54
rect 48 53 49 54
rect 47 53 48 54
rect 46 53 47 54
rect 45 53 46 54
rect 44 53 45 54
rect 43 53 44 54
rect 42 53 43 54
rect 41 53 42 54
rect 40 53 41 54
rect 39 53 40 54
rect 38 53 39 54
rect 37 53 38 54
rect 36 53 37 54
rect 35 53 36 54
rect 34 53 35 54
rect 33 53 34 54
rect 29 53 30 54
rect 28 53 29 54
rect 27 53 28 54
rect 26 53 27 54
rect 25 53 26 54
rect 24 53 25 54
rect 23 53 24 54
rect 22 53 23 54
rect 21 53 22 54
rect 20 53 21 54
rect 19 53 20 54
rect 18 53 19 54
rect 17 53 18 54
rect 193 54 194 55
rect 192 54 193 55
rect 191 54 192 55
rect 181 54 182 55
rect 180 54 181 55
rect 179 54 180 55
rect 178 54 179 55
rect 163 54 164 55
rect 100 54 101 55
rect 99 54 100 55
rect 98 54 99 55
rect 97 54 98 55
rect 96 54 97 55
rect 95 54 96 55
rect 94 54 95 55
rect 93 54 94 55
rect 92 54 93 55
rect 91 54 92 55
rect 90 54 91 55
rect 89 54 90 55
rect 88 54 89 55
rect 87 54 88 55
rect 86 54 87 55
rect 85 54 86 55
rect 84 54 85 55
rect 83 54 84 55
rect 82 54 83 55
rect 81 54 82 55
rect 80 54 81 55
rect 79 54 80 55
rect 78 54 79 55
rect 77 54 78 55
rect 76 54 77 55
rect 75 54 76 55
rect 74 54 75 55
rect 73 54 74 55
rect 72 54 73 55
rect 65 54 66 55
rect 64 54 65 55
rect 63 54 64 55
rect 62 54 63 55
rect 61 54 62 55
rect 60 54 61 55
rect 59 54 60 55
rect 58 54 59 55
rect 57 54 58 55
rect 56 54 57 55
rect 55 54 56 55
rect 54 54 55 55
rect 53 54 54 55
rect 52 54 53 55
rect 51 54 52 55
rect 50 54 51 55
rect 49 54 50 55
rect 48 54 49 55
rect 47 54 48 55
rect 46 54 47 55
rect 45 54 46 55
rect 44 54 45 55
rect 43 54 44 55
rect 42 54 43 55
rect 41 54 42 55
rect 40 54 41 55
rect 39 54 40 55
rect 38 54 39 55
rect 37 54 38 55
rect 36 54 37 55
rect 35 54 36 55
rect 34 54 35 55
rect 33 54 34 55
rect 32 54 33 55
rect 29 54 30 55
rect 28 54 29 55
rect 27 54 28 55
rect 26 54 27 55
rect 25 54 26 55
rect 24 54 25 55
rect 23 54 24 55
rect 22 54 23 55
rect 21 54 22 55
rect 20 54 21 55
rect 19 54 20 55
rect 18 54 19 55
rect 17 54 18 55
rect 194 55 195 56
rect 193 55 194 56
rect 192 55 193 56
rect 181 55 182 56
rect 180 55 181 56
rect 179 55 180 56
rect 122 55 123 56
rect 121 55 122 56
rect 120 55 121 56
rect 119 55 120 56
rect 118 55 119 56
rect 117 55 118 56
rect 116 55 117 56
rect 115 55 116 56
rect 98 55 99 56
rect 97 55 98 56
rect 96 55 97 56
rect 95 55 96 56
rect 94 55 95 56
rect 93 55 94 56
rect 92 55 93 56
rect 91 55 92 56
rect 90 55 91 56
rect 89 55 90 56
rect 88 55 89 56
rect 87 55 88 56
rect 86 55 87 56
rect 85 55 86 56
rect 84 55 85 56
rect 83 55 84 56
rect 82 55 83 56
rect 81 55 82 56
rect 80 55 81 56
rect 79 55 80 56
rect 78 55 79 56
rect 77 55 78 56
rect 76 55 77 56
rect 75 55 76 56
rect 74 55 75 56
rect 73 55 74 56
rect 72 55 73 56
rect 65 55 66 56
rect 64 55 65 56
rect 63 55 64 56
rect 62 55 63 56
rect 61 55 62 56
rect 60 55 61 56
rect 59 55 60 56
rect 58 55 59 56
rect 57 55 58 56
rect 56 55 57 56
rect 55 55 56 56
rect 54 55 55 56
rect 53 55 54 56
rect 52 55 53 56
rect 51 55 52 56
rect 50 55 51 56
rect 49 55 50 56
rect 48 55 49 56
rect 47 55 48 56
rect 46 55 47 56
rect 45 55 46 56
rect 44 55 45 56
rect 43 55 44 56
rect 42 55 43 56
rect 41 55 42 56
rect 40 55 41 56
rect 39 55 40 56
rect 38 55 39 56
rect 37 55 38 56
rect 36 55 37 56
rect 35 55 36 56
rect 34 55 35 56
rect 33 55 34 56
rect 32 55 33 56
rect 29 55 30 56
rect 28 55 29 56
rect 27 55 28 56
rect 26 55 27 56
rect 25 55 26 56
rect 24 55 25 56
rect 23 55 24 56
rect 22 55 23 56
rect 21 55 22 56
rect 20 55 21 56
rect 19 55 20 56
rect 18 55 19 56
rect 17 55 18 56
rect 195 56 196 57
rect 194 56 195 57
rect 193 56 194 57
rect 181 56 182 57
rect 180 56 181 57
rect 179 56 180 57
rect 124 56 125 57
rect 123 56 124 57
rect 122 56 123 57
rect 121 56 122 57
rect 120 56 121 57
rect 119 56 120 57
rect 118 56 119 57
rect 117 56 118 57
rect 116 56 117 57
rect 115 56 116 57
rect 114 56 115 57
rect 113 56 114 57
rect 112 56 113 57
rect 97 56 98 57
rect 96 56 97 57
rect 95 56 96 57
rect 94 56 95 57
rect 93 56 94 57
rect 92 56 93 57
rect 91 56 92 57
rect 90 56 91 57
rect 89 56 90 57
rect 88 56 89 57
rect 87 56 88 57
rect 86 56 87 57
rect 85 56 86 57
rect 84 56 85 57
rect 83 56 84 57
rect 82 56 83 57
rect 81 56 82 57
rect 80 56 81 57
rect 79 56 80 57
rect 78 56 79 57
rect 77 56 78 57
rect 76 56 77 57
rect 75 56 76 57
rect 74 56 75 57
rect 73 56 74 57
rect 72 56 73 57
rect 64 56 65 57
rect 63 56 64 57
rect 62 56 63 57
rect 61 56 62 57
rect 60 56 61 57
rect 59 56 60 57
rect 58 56 59 57
rect 57 56 58 57
rect 56 56 57 57
rect 55 56 56 57
rect 54 56 55 57
rect 53 56 54 57
rect 52 56 53 57
rect 51 56 52 57
rect 50 56 51 57
rect 49 56 50 57
rect 48 56 49 57
rect 47 56 48 57
rect 46 56 47 57
rect 45 56 46 57
rect 44 56 45 57
rect 43 56 44 57
rect 42 56 43 57
rect 41 56 42 57
rect 40 56 41 57
rect 39 56 40 57
rect 38 56 39 57
rect 37 56 38 57
rect 36 56 37 57
rect 35 56 36 57
rect 34 56 35 57
rect 33 56 34 57
rect 32 56 33 57
rect 31 56 32 57
rect 29 56 30 57
rect 28 56 29 57
rect 27 56 28 57
rect 26 56 27 57
rect 25 56 26 57
rect 24 56 25 57
rect 23 56 24 57
rect 22 56 23 57
rect 21 56 22 57
rect 20 56 21 57
rect 19 56 20 57
rect 18 56 19 57
rect 17 56 18 57
rect 197 57 198 58
rect 196 57 197 58
rect 195 57 196 58
rect 194 57 195 58
rect 193 57 194 58
rect 191 57 192 58
rect 190 57 191 58
rect 189 57 190 58
rect 181 57 182 58
rect 180 57 181 58
rect 179 57 180 58
rect 125 57 126 58
rect 124 57 125 58
rect 123 57 124 58
rect 122 57 123 58
rect 121 57 122 58
rect 120 57 121 58
rect 119 57 120 58
rect 118 57 119 58
rect 117 57 118 58
rect 116 57 117 58
rect 115 57 116 58
rect 114 57 115 58
rect 113 57 114 58
rect 112 57 113 58
rect 111 57 112 58
rect 110 57 111 58
rect 97 57 98 58
rect 96 57 97 58
rect 95 57 96 58
rect 94 57 95 58
rect 93 57 94 58
rect 92 57 93 58
rect 91 57 92 58
rect 90 57 91 58
rect 89 57 90 58
rect 88 57 89 58
rect 87 57 88 58
rect 86 57 87 58
rect 85 57 86 58
rect 84 57 85 58
rect 83 57 84 58
rect 82 57 83 58
rect 81 57 82 58
rect 80 57 81 58
rect 79 57 80 58
rect 78 57 79 58
rect 77 57 78 58
rect 76 57 77 58
rect 75 57 76 58
rect 74 57 75 58
rect 73 57 74 58
rect 72 57 73 58
rect 71 57 72 58
rect 64 57 65 58
rect 63 57 64 58
rect 62 57 63 58
rect 61 57 62 58
rect 60 57 61 58
rect 59 57 60 58
rect 58 57 59 58
rect 57 57 58 58
rect 56 57 57 58
rect 55 57 56 58
rect 54 57 55 58
rect 53 57 54 58
rect 52 57 53 58
rect 51 57 52 58
rect 50 57 51 58
rect 49 57 50 58
rect 48 57 49 58
rect 47 57 48 58
rect 46 57 47 58
rect 45 57 46 58
rect 44 57 45 58
rect 43 57 44 58
rect 42 57 43 58
rect 41 57 42 58
rect 40 57 41 58
rect 39 57 40 58
rect 38 57 39 58
rect 37 57 38 58
rect 36 57 37 58
rect 35 57 36 58
rect 34 57 35 58
rect 33 57 34 58
rect 32 57 33 58
rect 31 57 32 58
rect 28 57 29 58
rect 27 57 28 58
rect 26 57 27 58
rect 25 57 26 58
rect 24 57 25 58
rect 23 57 24 58
rect 22 57 23 58
rect 21 57 22 58
rect 20 57 21 58
rect 19 57 20 58
rect 18 57 19 58
rect 17 57 18 58
rect 197 58 198 59
rect 196 58 197 59
rect 195 58 196 59
rect 194 58 195 59
rect 193 58 194 59
rect 192 58 193 59
rect 191 58 192 59
rect 190 58 191 59
rect 189 58 190 59
rect 181 58 182 59
rect 180 58 181 59
rect 179 58 180 59
rect 163 58 164 59
rect 127 58 128 59
rect 126 58 127 59
rect 125 58 126 59
rect 124 58 125 59
rect 123 58 124 59
rect 122 58 123 59
rect 121 58 122 59
rect 120 58 121 59
rect 119 58 120 59
rect 118 58 119 59
rect 117 58 118 59
rect 116 58 117 59
rect 115 58 116 59
rect 114 58 115 59
rect 113 58 114 59
rect 112 58 113 59
rect 111 58 112 59
rect 110 58 111 59
rect 109 58 110 59
rect 108 58 109 59
rect 96 58 97 59
rect 95 58 96 59
rect 94 58 95 59
rect 93 58 94 59
rect 92 58 93 59
rect 91 58 92 59
rect 90 58 91 59
rect 89 58 90 59
rect 88 58 89 59
rect 87 58 88 59
rect 86 58 87 59
rect 85 58 86 59
rect 84 58 85 59
rect 83 58 84 59
rect 82 58 83 59
rect 81 58 82 59
rect 80 58 81 59
rect 79 58 80 59
rect 78 58 79 59
rect 77 58 78 59
rect 76 58 77 59
rect 75 58 76 59
rect 74 58 75 59
rect 73 58 74 59
rect 72 58 73 59
rect 71 58 72 59
rect 63 58 64 59
rect 62 58 63 59
rect 61 58 62 59
rect 60 58 61 59
rect 59 58 60 59
rect 58 58 59 59
rect 57 58 58 59
rect 56 58 57 59
rect 55 58 56 59
rect 54 58 55 59
rect 53 58 54 59
rect 52 58 53 59
rect 51 58 52 59
rect 50 58 51 59
rect 49 58 50 59
rect 48 58 49 59
rect 47 58 48 59
rect 46 58 47 59
rect 45 58 46 59
rect 44 58 45 59
rect 43 58 44 59
rect 42 58 43 59
rect 41 58 42 59
rect 40 58 41 59
rect 39 58 40 59
rect 38 58 39 59
rect 37 58 38 59
rect 36 58 37 59
rect 35 58 36 59
rect 34 58 35 59
rect 33 58 34 59
rect 32 58 33 59
rect 31 58 32 59
rect 30 58 31 59
rect 28 58 29 59
rect 27 58 28 59
rect 26 58 27 59
rect 25 58 26 59
rect 24 58 25 59
rect 23 58 24 59
rect 22 58 23 59
rect 21 58 22 59
rect 20 58 21 59
rect 19 58 20 59
rect 18 58 19 59
rect 180 59 181 60
rect 179 59 180 60
rect 178 59 179 60
rect 163 59 164 60
rect 128 59 129 60
rect 127 59 128 60
rect 126 59 127 60
rect 125 59 126 60
rect 124 59 125 60
rect 123 59 124 60
rect 122 59 123 60
rect 121 59 122 60
rect 120 59 121 60
rect 119 59 120 60
rect 118 59 119 60
rect 117 59 118 60
rect 116 59 117 60
rect 115 59 116 60
rect 114 59 115 60
rect 113 59 114 60
rect 112 59 113 60
rect 111 59 112 60
rect 110 59 111 60
rect 109 59 110 60
rect 108 59 109 60
rect 107 59 108 60
rect 95 59 96 60
rect 94 59 95 60
rect 93 59 94 60
rect 92 59 93 60
rect 91 59 92 60
rect 90 59 91 60
rect 89 59 90 60
rect 88 59 89 60
rect 87 59 88 60
rect 86 59 87 60
rect 85 59 86 60
rect 84 59 85 60
rect 83 59 84 60
rect 82 59 83 60
rect 81 59 82 60
rect 80 59 81 60
rect 79 59 80 60
rect 78 59 79 60
rect 77 59 78 60
rect 76 59 77 60
rect 75 59 76 60
rect 74 59 75 60
rect 73 59 74 60
rect 72 59 73 60
rect 71 59 72 60
rect 70 59 71 60
rect 63 59 64 60
rect 62 59 63 60
rect 61 59 62 60
rect 60 59 61 60
rect 59 59 60 60
rect 58 59 59 60
rect 57 59 58 60
rect 56 59 57 60
rect 55 59 56 60
rect 54 59 55 60
rect 53 59 54 60
rect 52 59 53 60
rect 51 59 52 60
rect 50 59 51 60
rect 49 59 50 60
rect 48 59 49 60
rect 47 59 48 60
rect 46 59 47 60
rect 45 59 46 60
rect 44 59 45 60
rect 43 59 44 60
rect 42 59 43 60
rect 41 59 42 60
rect 40 59 41 60
rect 39 59 40 60
rect 38 59 39 60
rect 37 59 38 60
rect 36 59 37 60
rect 35 59 36 60
rect 34 59 35 60
rect 33 59 34 60
rect 32 59 33 60
rect 31 59 32 60
rect 30 59 31 60
rect 29 59 30 60
rect 28 59 29 60
rect 27 59 28 60
rect 26 59 27 60
rect 25 59 26 60
rect 24 59 25 60
rect 23 59 24 60
rect 22 59 23 60
rect 21 59 22 60
rect 20 59 21 60
rect 19 59 20 60
rect 18 59 19 60
rect 180 60 181 61
rect 179 60 180 61
rect 178 60 179 61
rect 177 60 178 61
rect 164 60 165 61
rect 163 60 164 61
rect 129 60 130 61
rect 128 60 129 61
rect 127 60 128 61
rect 126 60 127 61
rect 125 60 126 61
rect 124 60 125 61
rect 123 60 124 61
rect 122 60 123 61
rect 121 60 122 61
rect 120 60 121 61
rect 119 60 120 61
rect 118 60 119 61
rect 117 60 118 61
rect 116 60 117 61
rect 115 60 116 61
rect 114 60 115 61
rect 113 60 114 61
rect 112 60 113 61
rect 111 60 112 61
rect 110 60 111 61
rect 109 60 110 61
rect 108 60 109 61
rect 107 60 108 61
rect 106 60 107 61
rect 105 60 106 61
rect 95 60 96 61
rect 94 60 95 61
rect 93 60 94 61
rect 92 60 93 61
rect 91 60 92 61
rect 90 60 91 61
rect 89 60 90 61
rect 88 60 89 61
rect 87 60 88 61
rect 86 60 87 61
rect 85 60 86 61
rect 84 60 85 61
rect 83 60 84 61
rect 82 60 83 61
rect 81 60 82 61
rect 80 60 81 61
rect 79 60 80 61
rect 78 60 79 61
rect 77 60 78 61
rect 76 60 77 61
rect 75 60 76 61
rect 74 60 75 61
rect 73 60 74 61
rect 72 60 73 61
rect 71 60 72 61
rect 70 60 71 61
rect 62 60 63 61
rect 61 60 62 61
rect 60 60 61 61
rect 59 60 60 61
rect 58 60 59 61
rect 57 60 58 61
rect 56 60 57 61
rect 55 60 56 61
rect 54 60 55 61
rect 53 60 54 61
rect 52 60 53 61
rect 51 60 52 61
rect 50 60 51 61
rect 49 60 50 61
rect 48 60 49 61
rect 47 60 48 61
rect 46 60 47 61
rect 45 60 46 61
rect 44 60 45 61
rect 43 60 44 61
rect 42 60 43 61
rect 41 60 42 61
rect 40 60 41 61
rect 39 60 40 61
rect 38 60 39 61
rect 37 60 38 61
rect 36 60 37 61
rect 35 60 36 61
rect 34 60 35 61
rect 33 60 34 61
rect 32 60 33 61
rect 31 60 32 61
rect 30 60 31 61
rect 29 60 30 61
rect 28 60 29 61
rect 27 60 28 61
rect 26 60 27 61
rect 25 60 26 61
rect 24 60 25 61
rect 23 60 24 61
rect 22 60 23 61
rect 21 60 22 61
rect 20 60 21 61
rect 19 60 20 61
rect 179 61 180 62
rect 178 61 179 62
rect 177 61 178 62
rect 176 61 177 62
rect 175 61 176 62
rect 174 61 175 62
rect 173 61 174 62
rect 172 61 173 62
rect 171 61 172 62
rect 170 61 171 62
rect 169 61 170 62
rect 168 61 169 62
rect 167 61 168 62
rect 166 61 167 62
rect 165 61 166 62
rect 164 61 165 62
rect 163 61 164 62
rect 130 61 131 62
rect 129 61 130 62
rect 128 61 129 62
rect 127 61 128 62
rect 126 61 127 62
rect 125 61 126 62
rect 124 61 125 62
rect 123 61 124 62
rect 122 61 123 62
rect 121 61 122 62
rect 120 61 121 62
rect 119 61 120 62
rect 118 61 119 62
rect 117 61 118 62
rect 116 61 117 62
rect 115 61 116 62
rect 114 61 115 62
rect 113 61 114 62
rect 112 61 113 62
rect 111 61 112 62
rect 110 61 111 62
rect 109 61 110 62
rect 108 61 109 62
rect 107 61 108 62
rect 106 61 107 62
rect 105 61 106 62
rect 104 61 105 62
rect 94 61 95 62
rect 93 61 94 62
rect 92 61 93 62
rect 91 61 92 62
rect 90 61 91 62
rect 89 61 90 62
rect 88 61 89 62
rect 87 61 88 62
rect 86 61 87 62
rect 85 61 86 62
rect 84 61 85 62
rect 83 61 84 62
rect 82 61 83 62
rect 81 61 82 62
rect 80 61 81 62
rect 79 61 80 62
rect 78 61 79 62
rect 77 61 78 62
rect 76 61 77 62
rect 75 61 76 62
rect 74 61 75 62
rect 73 61 74 62
rect 72 61 73 62
rect 71 61 72 62
rect 70 61 71 62
rect 69 61 70 62
rect 61 61 62 62
rect 60 61 61 62
rect 59 61 60 62
rect 58 61 59 62
rect 57 61 58 62
rect 56 61 57 62
rect 55 61 56 62
rect 54 61 55 62
rect 53 61 54 62
rect 52 61 53 62
rect 51 61 52 62
rect 50 61 51 62
rect 49 61 50 62
rect 48 61 49 62
rect 47 61 48 62
rect 46 61 47 62
rect 45 61 46 62
rect 44 61 45 62
rect 43 61 44 62
rect 42 61 43 62
rect 41 61 42 62
rect 40 61 41 62
rect 39 61 40 62
rect 38 61 39 62
rect 37 61 38 62
rect 36 61 37 62
rect 35 61 36 62
rect 34 61 35 62
rect 33 61 34 62
rect 32 61 33 62
rect 31 61 32 62
rect 30 61 31 62
rect 29 61 30 62
rect 28 61 29 62
rect 27 61 28 62
rect 26 61 27 62
rect 25 61 26 62
rect 24 61 25 62
rect 23 61 24 62
rect 22 61 23 62
rect 21 61 22 62
rect 20 61 21 62
rect 178 62 179 63
rect 177 62 178 63
rect 176 62 177 63
rect 175 62 176 63
rect 174 62 175 63
rect 173 62 174 63
rect 172 62 173 63
rect 171 62 172 63
rect 170 62 171 63
rect 169 62 170 63
rect 168 62 169 63
rect 167 62 168 63
rect 166 62 167 63
rect 165 62 166 63
rect 164 62 165 63
rect 163 62 164 63
rect 130 62 131 63
rect 129 62 130 63
rect 128 62 129 63
rect 127 62 128 63
rect 126 62 127 63
rect 125 62 126 63
rect 124 62 125 63
rect 123 62 124 63
rect 122 62 123 63
rect 121 62 122 63
rect 120 62 121 63
rect 119 62 120 63
rect 118 62 119 63
rect 117 62 118 63
rect 116 62 117 63
rect 115 62 116 63
rect 114 62 115 63
rect 113 62 114 63
rect 112 62 113 63
rect 111 62 112 63
rect 110 62 111 63
rect 109 62 110 63
rect 108 62 109 63
rect 107 62 108 63
rect 106 62 107 63
rect 105 62 106 63
rect 104 62 105 63
rect 103 62 104 63
rect 94 62 95 63
rect 93 62 94 63
rect 92 62 93 63
rect 91 62 92 63
rect 90 62 91 63
rect 89 62 90 63
rect 88 62 89 63
rect 87 62 88 63
rect 86 62 87 63
rect 85 62 86 63
rect 84 62 85 63
rect 83 62 84 63
rect 82 62 83 63
rect 81 62 82 63
rect 80 62 81 63
rect 79 62 80 63
rect 78 62 79 63
rect 77 62 78 63
rect 76 62 77 63
rect 75 62 76 63
rect 74 62 75 63
rect 73 62 74 63
rect 72 62 73 63
rect 71 62 72 63
rect 70 62 71 63
rect 69 62 70 63
rect 60 62 61 63
rect 59 62 60 63
rect 58 62 59 63
rect 57 62 58 63
rect 56 62 57 63
rect 55 62 56 63
rect 54 62 55 63
rect 53 62 54 63
rect 52 62 53 63
rect 51 62 52 63
rect 50 62 51 63
rect 49 62 50 63
rect 48 62 49 63
rect 47 62 48 63
rect 46 62 47 63
rect 45 62 46 63
rect 44 62 45 63
rect 43 62 44 63
rect 42 62 43 63
rect 41 62 42 63
rect 40 62 41 63
rect 39 62 40 63
rect 38 62 39 63
rect 37 62 38 63
rect 36 62 37 63
rect 35 62 36 63
rect 34 62 35 63
rect 33 62 34 63
rect 32 62 33 63
rect 31 62 32 63
rect 30 62 31 63
rect 29 62 30 63
rect 28 62 29 63
rect 27 62 28 63
rect 26 62 27 63
rect 25 62 26 63
rect 24 62 25 63
rect 23 62 24 63
rect 22 62 23 63
rect 21 62 22 63
rect 14 62 15 63
rect 197 63 198 64
rect 196 63 197 64
rect 189 63 190 64
rect 175 63 176 64
rect 167 63 168 64
rect 166 63 167 64
rect 165 63 166 64
rect 164 63 165 64
rect 163 63 164 64
rect 131 63 132 64
rect 130 63 131 64
rect 129 63 130 64
rect 128 63 129 64
rect 127 63 128 64
rect 126 63 127 64
rect 125 63 126 64
rect 124 63 125 64
rect 123 63 124 64
rect 122 63 123 64
rect 121 63 122 64
rect 120 63 121 64
rect 119 63 120 64
rect 118 63 119 64
rect 117 63 118 64
rect 116 63 117 64
rect 115 63 116 64
rect 114 63 115 64
rect 113 63 114 64
rect 112 63 113 64
rect 111 63 112 64
rect 110 63 111 64
rect 109 63 110 64
rect 108 63 109 64
rect 107 63 108 64
rect 106 63 107 64
rect 105 63 106 64
rect 104 63 105 64
rect 103 63 104 64
rect 102 63 103 64
rect 93 63 94 64
rect 92 63 93 64
rect 91 63 92 64
rect 90 63 91 64
rect 89 63 90 64
rect 88 63 89 64
rect 87 63 88 64
rect 86 63 87 64
rect 85 63 86 64
rect 84 63 85 64
rect 83 63 84 64
rect 82 63 83 64
rect 81 63 82 64
rect 80 63 81 64
rect 79 63 80 64
rect 78 63 79 64
rect 77 63 78 64
rect 76 63 77 64
rect 75 63 76 64
rect 74 63 75 64
rect 73 63 74 64
rect 72 63 73 64
rect 71 63 72 64
rect 70 63 71 64
rect 69 63 70 64
rect 68 63 69 64
rect 59 63 60 64
rect 58 63 59 64
rect 57 63 58 64
rect 56 63 57 64
rect 55 63 56 64
rect 54 63 55 64
rect 53 63 54 64
rect 52 63 53 64
rect 51 63 52 64
rect 50 63 51 64
rect 49 63 50 64
rect 48 63 49 64
rect 47 63 48 64
rect 46 63 47 64
rect 45 63 46 64
rect 44 63 45 64
rect 43 63 44 64
rect 42 63 43 64
rect 41 63 42 64
rect 40 63 41 64
rect 39 63 40 64
rect 38 63 39 64
rect 37 63 38 64
rect 36 63 37 64
rect 35 63 36 64
rect 34 63 35 64
rect 33 63 34 64
rect 32 63 33 64
rect 31 63 32 64
rect 30 63 31 64
rect 29 63 30 64
rect 28 63 29 64
rect 27 63 28 64
rect 26 63 27 64
rect 25 63 26 64
rect 24 63 25 64
rect 23 63 24 64
rect 22 63 23 64
rect 21 63 22 64
rect 16 63 17 64
rect 15 63 16 64
rect 14 63 15 64
rect 13 63 14 64
rect 12 63 13 64
rect 196 64 197 65
rect 195 64 196 65
rect 194 64 195 65
rect 193 64 194 65
rect 192 64 193 65
rect 191 64 192 65
rect 190 64 191 65
rect 189 64 190 65
rect 164 64 165 65
rect 163 64 164 65
rect 132 64 133 65
rect 131 64 132 65
rect 130 64 131 65
rect 129 64 130 65
rect 128 64 129 65
rect 127 64 128 65
rect 126 64 127 65
rect 125 64 126 65
rect 124 64 125 65
rect 123 64 124 65
rect 122 64 123 65
rect 121 64 122 65
rect 120 64 121 65
rect 119 64 120 65
rect 118 64 119 65
rect 117 64 118 65
rect 116 64 117 65
rect 115 64 116 65
rect 114 64 115 65
rect 113 64 114 65
rect 112 64 113 65
rect 111 64 112 65
rect 110 64 111 65
rect 109 64 110 65
rect 108 64 109 65
rect 107 64 108 65
rect 106 64 107 65
rect 105 64 106 65
rect 104 64 105 65
rect 103 64 104 65
rect 102 64 103 65
rect 93 64 94 65
rect 92 64 93 65
rect 91 64 92 65
rect 90 64 91 65
rect 89 64 90 65
rect 88 64 89 65
rect 87 64 88 65
rect 86 64 87 65
rect 85 64 86 65
rect 84 64 85 65
rect 83 64 84 65
rect 82 64 83 65
rect 81 64 82 65
rect 80 64 81 65
rect 79 64 80 65
rect 78 64 79 65
rect 77 64 78 65
rect 76 64 77 65
rect 75 64 76 65
rect 74 64 75 65
rect 73 64 74 65
rect 72 64 73 65
rect 71 64 72 65
rect 70 64 71 65
rect 69 64 70 65
rect 68 64 69 65
rect 58 64 59 65
rect 57 64 58 65
rect 56 64 57 65
rect 55 64 56 65
rect 54 64 55 65
rect 53 64 54 65
rect 52 64 53 65
rect 51 64 52 65
rect 50 64 51 65
rect 49 64 50 65
rect 48 64 49 65
rect 47 64 48 65
rect 46 64 47 65
rect 45 64 46 65
rect 44 64 45 65
rect 43 64 44 65
rect 42 64 43 65
rect 41 64 42 65
rect 40 64 41 65
rect 39 64 40 65
rect 38 64 39 65
rect 37 64 38 65
rect 36 64 37 65
rect 35 64 36 65
rect 34 64 35 65
rect 33 64 34 65
rect 32 64 33 65
rect 31 64 32 65
rect 30 64 31 65
rect 29 64 30 65
rect 28 64 29 65
rect 27 64 28 65
rect 26 64 27 65
rect 25 64 26 65
rect 24 64 25 65
rect 23 64 24 65
rect 22 64 23 65
rect 21 64 22 65
rect 16 64 17 65
rect 15 64 16 65
rect 14 64 15 65
rect 13 64 14 65
rect 12 64 13 65
rect 11 64 12 65
rect 10 64 11 65
rect 196 65 197 66
rect 195 65 196 66
rect 194 65 195 66
rect 193 65 194 66
rect 192 65 193 66
rect 191 65 192 66
rect 190 65 191 66
rect 189 65 190 66
rect 163 65 164 66
rect 132 65 133 66
rect 131 65 132 66
rect 130 65 131 66
rect 129 65 130 66
rect 128 65 129 66
rect 127 65 128 66
rect 126 65 127 66
rect 125 65 126 66
rect 124 65 125 66
rect 123 65 124 66
rect 122 65 123 66
rect 121 65 122 66
rect 120 65 121 66
rect 119 65 120 66
rect 118 65 119 66
rect 117 65 118 66
rect 116 65 117 66
rect 115 65 116 66
rect 114 65 115 66
rect 113 65 114 66
rect 112 65 113 66
rect 111 65 112 66
rect 110 65 111 66
rect 109 65 110 66
rect 108 65 109 66
rect 107 65 108 66
rect 106 65 107 66
rect 105 65 106 66
rect 104 65 105 66
rect 103 65 104 66
rect 102 65 103 66
rect 101 65 102 66
rect 92 65 93 66
rect 91 65 92 66
rect 90 65 91 66
rect 89 65 90 66
rect 88 65 89 66
rect 87 65 88 66
rect 86 65 87 66
rect 85 65 86 66
rect 84 65 85 66
rect 83 65 84 66
rect 82 65 83 66
rect 81 65 82 66
rect 80 65 81 66
rect 79 65 80 66
rect 78 65 79 66
rect 77 65 78 66
rect 76 65 77 66
rect 75 65 76 66
rect 74 65 75 66
rect 73 65 74 66
rect 72 65 73 66
rect 71 65 72 66
rect 70 65 71 66
rect 69 65 70 66
rect 68 65 69 66
rect 67 65 68 66
rect 57 65 58 66
rect 56 65 57 66
rect 55 65 56 66
rect 54 65 55 66
rect 53 65 54 66
rect 52 65 53 66
rect 51 65 52 66
rect 50 65 51 66
rect 49 65 50 66
rect 48 65 49 66
rect 47 65 48 66
rect 46 65 47 66
rect 45 65 46 66
rect 44 65 45 66
rect 43 65 44 66
rect 42 65 43 66
rect 41 65 42 66
rect 40 65 41 66
rect 39 65 40 66
rect 38 65 39 66
rect 37 65 38 66
rect 36 65 37 66
rect 35 65 36 66
rect 34 65 35 66
rect 33 65 34 66
rect 32 65 33 66
rect 31 65 32 66
rect 30 65 31 66
rect 29 65 30 66
rect 28 65 29 66
rect 27 65 28 66
rect 26 65 27 66
rect 25 65 26 66
rect 24 65 25 66
rect 23 65 24 66
rect 22 65 23 66
rect 21 65 22 66
rect 17 65 18 66
rect 16 65 17 66
rect 15 65 16 66
rect 14 65 15 66
rect 13 65 14 66
rect 12 65 13 66
rect 11 65 12 66
rect 10 65 11 66
rect 133 66 134 67
rect 132 66 133 67
rect 131 66 132 67
rect 130 66 131 67
rect 129 66 130 67
rect 128 66 129 67
rect 127 66 128 67
rect 126 66 127 67
rect 125 66 126 67
rect 124 66 125 67
rect 123 66 124 67
rect 122 66 123 67
rect 121 66 122 67
rect 120 66 121 67
rect 119 66 120 67
rect 118 66 119 67
rect 117 66 118 67
rect 116 66 117 67
rect 115 66 116 67
rect 114 66 115 67
rect 113 66 114 67
rect 112 66 113 67
rect 111 66 112 67
rect 110 66 111 67
rect 109 66 110 67
rect 108 66 109 67
rect 107 66 108 67
rect 106 66 107 67
rect 105 66 106 67
rect 104 66 105 67
rect 103 66 104 67
rect 102 66 103 67
rect 101 66 102 67
rect 100 66 101 67
rect 92 66 93 67
rect 91 66 92 67
rect 90 66 91 67
rect 89 66 90 67
rect 88 66 89 67
rect 87 66 88 67
rect 86 66 87 67
rect 85 66 86 67
rect 84 66 85 67
rect 83 66 84 67
rect 82 66 83 67
rect 81 66 82 67
rect 80 66 81 67
rect 79 66 80 67
rect 78 66 79 67
rect 77 66 78 67
rect 76 66 77 67
rect 75 66 76 67
rect 74 66 75 67
rect 73 66 74 67
rect 72 66 73 67
rect 71 66 72 67
rect 70 66 71 67
rect 69 66 70 67
rect 68 66 69 67
rect 67 66 68 67
rect 66 66 67 67
rect 55 66 56 67
rect 54 66 55 67
rect 53 66 54 67
rect 52 66 53 67
rect 51 66 52 67
rect 50 66 51 67
rect 49 66 50 67
rect 48 66 49 67
rect 47 66 48 67
rect 46 66 47 67
rect 45 66 46 67
rect 44 66 45 67
rect 43 66 44 67
rect 42 66 43 67
rect 41 66 42 67
rect 40 66 41 67
rect 39 66 40 67
rect 38 66 39 67
rect 37 66 38 67
rect 36 66 37 67
rect 35 66 36 67
rect 34 66 35 67
rect 33 66 34 67
rect 32 66 33 67
rect 31 66 32 67
rect 30 66 31 67
rect 29 66 30 67
rect 28 66 29 67
rect 27 66 28 67
rect 26 66 27 67
rect 25 66 26 67
rect 24 66 25 67
rect 23 66 24 67
rect 22 66 23 67
rect 21 66 22 67
rect 20 66 21 67
rect 16 66 17 67
rect 15 66 16 67
rect 14 66 15 67
rect 13 66 14 67
rect 12 66 13 67
rect 11 66 12 67
rect 10 66 11 67
rect 9 66 10 67
rect 163 67 164 68
rect 134 67 135 68
rect 133 67 134 68
rect 132 67 133 68
rect 131 67 132 68
rect 130 67 131 68
rect 129 67 130 68
rect 128 67 129 68
rect 127 67 128 68
rect 126 67 127 68
rect 125 67 126 68
rect 124 67 125 68
rect 123 67 124 68
rect 122 67 123 68
rect 121 67 122 68
rect 120 67 121 68
rect 119 67 120 68
rect 118 67 119 68
rect 117 67 118 68
rect 116 67 117 68
rect 115 67 116 68
rect 114 67 115 68
rect 113 67 114 68
rect 112 67 113 68
rect 111 67 112 68
rect 110 67 111 68
rect 109 67 110 68
rect 108 67 109 68
rect 107 67 108 68
rect 106 67 107 68
rect 105 67 106 68
rect 104 67 105 68
rect 103 67 104 68
rect 102 67 103 68
rect 101 67 102 68
rect 100 67 101 68
rect 92 67 93 68
rect 91 67 92 68
rect 90 67 91 68
rect 89 67 90 68
rect 88 67 89 68
rect 87 67 88 68
rect 86 67 87 68
rect 85 67 86 68
rect 84 67 85 68
rect 83 67 84 68
rect 82 67 83 68
rect 81 67 82 68
rect 80 67 81 68
rect 79 67 80 68
rect 78 67 79 68
rect 77 67 78 68
rect 76 67 77 68
rect 75 67 76 68
rect 74 67 75 68
rect 73 67 74 68
rect 72 67 73 68
rect 71 67 72 68
rect 70 67 71 68
rect 69 67 70 68
rect 68 67 69 68
rect 67 67 68 68
rect 66 67 67 68
rect 65 67 66 68
rect 54 67 55 68
rect 53 67 54 68
rect 52 67 53 68
rect 51 67 52 68
rect 50 67 51 68
rect 49 67 50 68
rect 48 67 49 68
rect 47 67 48 68
rect 46 67 47 68
rect 45 67 46 68
rect 44 67 45 68
rect 43 67 44 68
rect 42 67 43 68
rect 41 67 42 68
rect 40 67 41 68
rect 39 67 40 68
rect 38 67 39 68
rect 37 67 38 68
rect 36 67 37 68
rect 35 67 36 68
rect 34 67 35 68
rect 33 67 34 68
rect 32 67 33 68
rect 31 67 32 68
rect 30 67 31 68
rect 29 67 30 68
rect 28 67 29 68
rect 27 67 28 68
rect 26 67 27 68
rect 25 67 26 68
rect 24 67 25 68
rect 23 67 24 68
rect 22 67 23 68
rect 21 67 22 68
rect 20 67 21 68
rect 16 67 17 68
rect 15 67 16 68
rect 14 67 15 68
rect 13 67 14 68
rect 12 67 13 68
rect 11 67 12 68
rect 10 67 11 68
rect 9 67 10 68
rect 8 67 9 68
rect 180 68 181 69
rect 163 68 164 69
rect 135 68 136 69
rect 134 68 135 69
rect 133 68 134 69
rect 132 68 133 69
rect 131 68 132 69
rect 130 68 131 69
rect 129 68 130 69
rect 128 68 129 69
rect 127 68 128 69
rect 126 68 127 69
rect 125 68 126 69
rect 124 68 125 69
rect 123 68 124 69
rect 122 68 123 69
rect 121 68 122 69
rect 120 68 121 69
rect 119 68 120 69
rect 118 68 119 69
rect 117 68 118 69
rect 116 68 117 69
rect 115 68 116 69
rect 114 68 115 69
rect 113 68 114 69
rect 112 68 113 69
rect 111 68 112 69
rect 110 68 111 69
rect 109 68 110 69
rect 108 68 109 69
rect 107 68 108 69
rect 106 68 107 69
rect 105 68 106 69
rect 104 68 105 69
rect 103 68 104 69
rect 102 68 103 69
rect 101 68 102 69
rect 100 68 101 69
rect 99 68 100 69
rect 91 68 92 69
rect 90 68 91 69
rect 89 68 90 69
rect 88 68 89 69
rect 87 68 88 69
rect 86 68 87 69
rect 85 68 86 69
rect 84 68 85 69
rect 83 68 84 69
rect 82 68 83 69
rect 81 68 82 69
rect 80 68 81 69
rect 79 68 80 69
rect 78 68 79 69
rect 77 68 78 69
rect 76 68 77 69
rect 75 68 76 69
rect 74 68 75 69
rect 73 68 74 69
rect 72 68 73 69
rect 71 68 72 69
rect 70 68 71 69
rect 69 68 70 69
rect 68 68 69 69
rect 67 68 68 69
rect 66 68 67 69
rect 65 68 66 69
rect 64 68 65 69
rect 52 68 53 69
rect 51 68 52 69
rect 50 68 51 69
rect 49 68 50 69
rect 48 68 49 69
rect 47 68 48 69
rect 46 68 47 69
rect 45 68 46 69
rect 44 68 45 69
rect 43 68 44 69
rect 42 68 43 69
rect 41 68 42 69
rect 40 68 41 69
rect 39 68 40 69
rect 38 68 39 69
rect 37 68 38 69
rect 36 68 37 69
rect 35 68 36 69
rect 34 68 35 69
rect 33 68 34 69
rect 32 68 33 69
rect 31 68 32 69
rect 30 68 31 69
rect 29 68 30 69
rect 28 68 29 69
rect 27 68 28 69
rect 26 68 27 69
rect 25 68 26 69
rect 24 68 25 69
rect 23 68 24 69
rect 22 68 23 69
rect 21 68 22 69
rect 20 68 21 69
rect 19 68 20 69
rect 16 68 17 69
rect 15 68 16 69
rect 14 68 15 69
rect 13 68 14 69
rect 12 68 13 69
rect 11 68 12 69
rect 10 68 11 69
rect 9 68 10 69
rect 8 68 9 69
rect 180 69 181 70
rect 179 69 180 70
rect 164 69 165 70
rect 163 69 164 70
rect 136 69 137 70
rect 135 69 136 70
rect 134 69 135 70
rect 133 69 134 70
rect 122 69 123 70
rect 121 69 122 70
rect 120 69 121 70
rect 119 69 120 70
rect 118 69 119 70
rect 117 69 118 70
rect 116 69 117 70
rect 115 69 116 70
rect 114 69 115 70
rect 113 69 114 70
rect 112 69 113 70
rect 111 69 112 70
rect 110 69 111 70
rect 109 69 110 70
rect 108 69 109 70
rect 107 69 108 70
rect 106 69 107 70
rect 105 69 106 70
rect 104 69 105 70
rect 103 69 104 70
rect 102 69 103 70
rect 101 69 102 70
rect 100 69 101 70
rect 99 69 100 70
rect 98 69 99 70
rect 91 69 92 70
rect 90 69 91 70
rect 89 69 90 70
rect 88 69 89 70
rect 87 69 88 70
rect 86 69 87 70
rect 85 69 86 70
rect 84 69 85 70
rect 83 69 84 70
rect 82 69 83 70
rect 81 69 82 70
rect 80 69 81 70
rect 79 69 80 70
rect 78 69 79 70
rect 77 69 78 70
rect 76 69 77 70
rect 75 69 76 70
rect 74 69 75 70
rect 73 69 74 70
rect 72 69 73 70
rect 71 69 72 70
rect 70 69 71 70
rect 69 69 70 70
rect 68 69 69 70
rect 67 69 68 70
rect 66 69 67 70
rect 65 69 66 70
rect 64 69 65 70
rect 51 69 52 70
rect 50 69 51 70
rect 49 69 50 70
rect 48 69 49 70
rect 47 69 48 70
rect 46 69 47 70
rect 45 69 46 70
rect 44 69 45 70
rect 43 69 44 70
rect 42 69 43 70
rect 41 69 42 70
rect 40 69 41 70
rect 39 69 40 70
rect 38 69 39 70
rect 37 69 38 70
rect 36 69 37 70
rect 35 69 36 70
rect 34 69 35 70
rect 33 69 34 70
rect 32 69 33 70
rect 31 69 32 70
rect 30 69 31 70
rect 29 69 30 70
rect 28 69 29 70
rect 27 69 28 70
rect 26 69 27 70
rect 25 69 26 70
rect 24 69 25 70
rect 23 69 24 70
rect 22 69 23 70
rect 21 69 22 70
rect 20 69 21 70
rect 19 69 20 70
rect 15 69 16 70
rect 14 69 15 70
rect 13 69 14 70
rect 12 69 13 70
rect 11 69 12 70
rect 10 69 11 70
rect 9 69 10 70
rect 8 69 9 70
rect 189 70 190 71
rect 180 70 181 71
rect 179 70 180 71
rect 178 70 179 71
rect 177 70 178 71
rect 176 70 177 71
rect 175 70 176 71
rect 174 70 175 71
rect 173 70 174 71
rect 172 70 173 71
rect 171 70 172 71
rect 170 70 171 71
rect 169 70 170 71
rect 168 70 169 71
rect 167 70 168 71
rect 166 70 167 71
rect 165 70 166 71
rect 164 70 165 71
rect 163 70 164 71
rect 119 70 120 71
rect 118 70 119 71
rect 117 70 118 71
rect 116 70 117 71
rect 115 70 116 71
rect 114 70 115 71
rect 113 70 114 71
rect 112 70 113 71
rect 111 70 112 71
rect 110 70 111 71
rect 109 70 110 71
rect 108 70 109 71
rect 107 70 108 71
rect 106 70 107 71
rect 105 70 106 71
rect 104 70 105 71
rect 103 70 104 71
rect 102 70 103 71
rect 101 70 102 71
rect 100 70 101 71
rect 99 70 100 71
rect 98 70 99 71
rect 90 70 91 71
rect 89 70 90 71
rect 88 70 89 71
rect 87 70 88 71
rect 86 70 87 71
rect 85 70 86 71
rect 84 70 85 71
rect 83 70 84 71
rect 82 70 83 71
rect 81 70 82 71
rect 80 70 81 71
rect 79 70 80 71
rect 78 70 79 71
rect 77 70 78 71
rect 76 70 77 71
rect 75 70 76 71
rect 74 70 75 71
rect 73 70 74 71
rect 72 70 73 71
rect 71 70 72 71
rect 70 70 71 71
rect 69 70 70 71
rect 68 70 69 71
rect 67 70 68 71
rect 66 70 67 71
rect 65 70 66 71
rect 64 70 65 71
rect 63 70 64 71
rect 49 70 50 71
rect 48 70 49 71
rect 47 70 48 71
rect 46 70 47 71
rect 45 70 46 71
rect 44 70 45 71
rect 43 70 44 71
rect 42 70 43 71
rect 41 70 42 71
rect 40 70 41 71
rect 39 70 40 71
rect 38 70 39 71
rect 37 70 38 71
rect 36 70 37 71
rect 35 70 36 71
rect 34 70 35 71
rect 33 70 34 71
rect 32 70 33 71
rect 31 70 32 71
rect 30 70 31 71
rect 29 70 30 71
rect 28 70 29 71
rect 27 70 28 71
rect 26 70 27 71
rect 25 70 26 71
rect 24 70 25 71
rect 23 70 24 71
rect 22 70 23 71
rect 21 70 22 71
rect 20 70 21 71
rect 19 70 20 71
rect 15 70 16 71
rect 14 70 15 71
rect 13 70 14 71
rect 12 70 13 71
rect 11 70 12 71
rect 10 70 11 71
rect 9 70 10 71
rect 8 70 9 71
rect 191 71 192 72
rect 190 71 191 72
rect 189 71 190 72
rect 180 71 181 72
rect 179 71 180 72
rect 178 71 179 72
rect 177 71 178 72
rect 176 71 177 72
rect 175 71 176 72
rect 174 71 175 72
rect 173 71 174 72
rect 172 71 173 72
rect 171 71 172 72
rect 170 71 171 72
rect 169 71 170 72
rect 168 71 169 72
rect 167 71 168 72
rect 166 71 167 72
rect 165 71 166 72
rect 164 71 165 72
rect 163 71 164 72
rect 117 71 118 72
rect 116 71 117 72
rect 115 71 116 72
rect 114 71 115 72
rect 113 71 114 72
rect 112 71 113 72
rect 111 71 112 72
rect 110 71 111 72
rect 109 71 110 72
rect 108 71 109 72
rect 107 71 108 72
rect 106 71 107 72
rect 105 71 106 72
rect 104 71 105 72
rect 103 71 104 72
rect 102 71 103 72
rect 101 71 102 72
rect 100 71 101 72
rect 99 71 100 72
rect 98 71 99 72
rect 97 71 98 72
rect 90 71 91 72
rect 89 71 90 72
rect 88 71 89 72
rect 87 71 88 72
rect 86 71 87 72
rect 85 71 86 72
rect 84 71 85 72
rect 83 71 84 72
rect 82 71 83 72
rect 81 71 82 72
rect 80 71 81 72
rect 79 71 80 72
rect 78 71 79 72
rect 77 71 78 72
rect 76 71 77 72
rect 75 71 76 72
rect 74 71 75 72
rect 73 71 74 72
rect 72 71 73 72
rect 71 71 72 72
rect 70 71 71 72
rect 69 71 70 72
rect 68 71 69 72
rect 67 71 68 72
rect 66 71 67 72
rect 65 71 66 72
rect 64 71 65 72
rect 63 71 64 72
rect 62 71 63 72
rect 61 71 62 72
rect 48 71 49 72
rect 47 71 48 72
rect 46 71 47 72
rect 45 71 46 72
rect 44 71 45 72
rect 43 71 44 72
rect 42 71 43 72
rect 41 71 42 72
rect 40 71 41 72
rect 39 71 40 72
rect 38 71 39 72
rect 37 71 38 72
rect 36 71 37 72
rect 35 71 36 72
rect 34 71 35 72
rect 32 71 33 72
rect 31 71 32 72
rect 30 71 31 72
rect 29 71 30 72
rect 28 71 29 72
rect 27 71 28 72
rect 26 71 27 72
rect 25 71 26 72
rect 24 71 25 72
rect 23 71 24 72
rect 22 71 23 72
rect 21 71 22 72
rect 20 71 21 72
rect 19 71 20 72
rect 18 71 19 72
rect 14 71 15 72
rect 13 71 14 72
rect 12 71 13 72
rect 11 71 12 72
rect 10 71 11 72
rect 9 71 10 72
rect 8 71 9 72
rect 193 72 194 73
rect 192 72 193 73
rect 191 72 192 73
rect 190 72 191 73
rect 189 72 190 73
rect 180 72 181 73
rect 179 72 180 73
rect 168 72 169 73
rect 167 72 168 73
rect 166 72 167 73
rect 165 72 166 73
rect 164 72 165 73
rect 163 72 164 73
rect 115 72 116 73
rect 114 72 115 73
rect 113 72 114 73
rect 112 72 113 73
rect 111 72 112 73
rect 110 72 111 73
rect 109 72 110 73
rect 108 72 109 73
rect 107 72 108 73
rect 106 72 107 73
rect 105 72 106 73
rect 104 72 105 73
rect 103 72 104 73
rect 102 72 103 73
rect 101 72 102 73
rect 100 72 101 73
rect 99 72 100 73
rect 98 72 99 73
rect 97 72 98 73
rect 89 72 90 73
rect 88 72 89 73
rect 87 72 88 73
rect 86 72 87 73
rect 85 72 86 73
rect 84 72 85 73
rect 83 72 84 73
rect 82 72 83 73
rect 81 72 82 73
rect 80 72 81 73
rect 79 72 80 73
rect 78 72 79 73
rect 77 72 78 73
rect 76 72 77 73
rect 75 72 76 73
rect 74 72 75 73
rect 73 72 74 73
rect 72 72 73 73
rect 71 72 72 73
rect 70 72 71 73
rect 69 72 70 73
rect 68 72 69 73
rect 67 72 68 73
rect 66 72 67 73
rect 65 72 66 73
rect 64 72 65 73
rect 63 72 64 73
rect 62 72 63 73
rect 61 72 62 73
rect 60 72 61 73
rect 45 72 46 73
rect 44 72 45 73
rect 43 72 44 73
rect 42 72 43 73
rect 41 72 42 73
rect 40 72 41 73
rect 39 72 40 73
rect 38 72 39 73
rect 30 72 31 73
rect 29 72 30 73
rect 28 72 29 73
rect 27 72 28 73
rect 26 72 27 73
rect 25 72 26 73
rect 24 72 25 73
rect 23 72 24 73
rect 22 72 23 73
rect 21 72 22 73
rect 20 72 21 73
rect 19 72 20 73
rect 18 72 19 73
rect 14 72 15 73
rect 13 72 14 73
rect 12 72 13 73
rect 11 72 12 73
rect 10 72 11 73
rect 9 72 10 73
rect 196 73 197 74
rect 195 73 196 74
rect 194 73 195 74
rect 193 73 194 74
rect 192 73 193 74
rect 191 73 192 74
rect 189 73 190 74
rect 180 73 181 74
rect 169 73 170 74
rect 168 73 169 74
rect 167 73 168 74
rect 166 73 167 74
rect 165 73 166 74
rect 164 73 165 74
rect 114 73 115 74
rect 113 73 114 74
rect 112 73 113 74
rect 111 73 112 74
rect 110 73 111 74
rect 109 73 110 74
rect 108 73 109 74
rect 107 73 108 74
rect 106 73 107 74
rect 105 73 106 74
rect 104 73 105 74
rect 103 73 104 74
rect 102 73 103 74
rect 101 73 102 74
rect 100 73 101 74
rect 99 73 100 74
rect 98 73 99 74
rect 97 73 98 74
rect 96 73 97 74
rect 89 73 90 74
rect 88 73 89 74
rect 87 73 88 74
rect 86 73 87 74
rect 85 73 86 74
rect 84 73 85 74
rect 83 73 84 74
rect 82 73 83 74
rect 81 73 82 74
rect 80 73 81 74
rect 79 73 80 74
rect 78 73 79 74
rect 77 73 78 74
rect 76 73 77 74
rect 75 73 76 74
rect 74 73 75 74
rect 73 73 74 74
rect 72 73 73 74
rect 71 73 72 74
rect 70 73 71 74
rect 69 73 70 74
rect 68 73 69 74
rect 67 73 68 74
rect 66 73 67 74
rect 65 73 66 74
rect 64 73 65 74
rect 63 73 64 74
rect 62 73 63 74
rect 61 73 62 74
rect 60 73 61 74
rect 59 73 60 74
rect 29 73 30 74
rect 28 73 29 74
rect 27 73 28 74
rect 26 73 27 74
rect 25 73 26 74
rect 24 73 25 74
rect 23 73 24 74
rect 22 73 23 74
rect 21 73 22 74
rect 20 73 21 74
rect 19 73 20 74
rect 18 73 19 74
rect 14 73 15 74
rect 13 73 14 74
rect 12 73 13 74
rect 11 73 12 74
rect 10 73 11 74
rect 9 73 10 74
rect 197 74 198 75
rect 196 74 197 75
rect 195 74 196 75
rect 194 74 195 75
rect 180 74 181 75
rect 170 74 171 75
rect 169 74 170 75
rect 168 74 169 75
rect 167 74 168 75
rect 166 74 167 75
rect 165 74 166 75
rect 113 74 114 75
rect 112 74 113 75
rect 111 74 112 75
rect 110 74 111 75
rect 109 74 110 75
rect 108 74 109 75
rect 107 74 108 75
rect 106 74 107 75
rect 105 74 106 75
rect 104 74 105 75
rect 103 74 104 75
rect 102 74 103 75
rect 101 74 102 75
rect 100 74 101 75
rect 99 74 100 75
rect 98 74 99 75
rect 97 74 98 75
rect 96 74 97 75
rect 88 74 89 75
rect 87 74 88 75
rect 86 74 87 75
rect 85 74 86 75
rect 84 74 85 75
rect 83 74 84 75
rect 82 74 83 75
rect 81 74 82 75
rect 80 74 81 75
rect 79 74 80 75
rect 78 74 79 75
rect 77 74 78 75
rect 76 74 77 75
rect 75 74 76 75
rect 74 74 75 75
rect 73 74 74 75
rect 72 74 73 75
rect 71 74 72 75
rect 70 74 71 75
rect 69 74 70 75
rect 68 74 69 75
rect 67 74 68 75
rect 66 74 67 75
rect 65 74 66 75
rect 64 74 65 75
rect 63 74 64 75
rect 62 74 63 75
rect 61 74 62 75
rect 60 74 61 75
rect 59 74 60 75
rect 58 74 59 75
rect 57 74 58 75
rect 28 74 29 75
rect 27 74 28 75
rect 26 74 27 75
rect 25 74 26 75
rect 24 74 25 75
rect 23 74 24 75
rect 22 74 23 75
rect 21 74 22 75
rect 20 74 21 75
rect 19 74 20 75
rect 14 74 15 75
rect 13 74 14 75
rect 12 74 13 75
rect 11 74 12 75
rect 10 74 11 75
rect 9 74 10 75
rect 195 75 196 76
rect 194 75 195 76
rect 193 75 194 76
rect 171 75 172 76
rect 170 75 171 76
rect 169 75 170 76
rect 168 75 169 76
rect 167 75 168 76
rect 166 75 167 76
rect 112 75 113 76
rect 111 75 112 76
rect 110 75 111 76
rect 109 75 110 76
rect 108 75 109 76
rect 107 75 108 76
rect 106 75 107 76
rect 105 75 106 76
rect 104 75 105 76
rect 103 75 104 76
rect 102 75 103 76
rect 101 75 102 76
rect 100 75 101 76
rect 99 75 100 76
rect 98 75 99 76
rect 97 75 98 76
rect 96 75 97 76
rect 95 75 96 76
rect 87 75 88 76
rect 86 75 87 76
rect 85 75 86 76
rect 84 75 85 76
rect 83 75 84 76
rect 82 75 83 76
rect 81 75 82 76
rect 80 75 81 76
rect 79 75 80 76
rect 78 75 79 76
rect 77 75 78 76
rect 76 75 77 76
rect 75 75 76 76
rect 74 75 75 76
rect 73 75 74 76
rect 72 75 73 76
rect 71 75 72 76
rect 70 75 71 76
rect 69 75 70 76
rect 68 75 69 76
rect 67 75 68 76
rect 66 75 67 76
rect 65 75 66 76
rect 64 75 65 76
rect 63 75 64 76
rect 62 75 63 76
rect 61 75 62 76
rect 60 75 61 76
rect 59 75 60 76
rect 58 75 59 76
rect 57 75 58 76
rect 56 75 57 76
rect 28 75 29 76
rect 27 75 28 76
rect 26 75 27 76
rect 25 75 26 76
rect 24 75 25 76
rect 23 75 24 76
rect 22 75 23 76
rect 21 75 22 76
rect 20 75 21 76
rect 19 75 20 76
rect 14 75 15 76
rect 13 75 14 76
rect 12 75 13 76
rect 11 75 12 76
rect 10 75 11 76
rect 193 76 194 77
rect 192 76 193 77
rect 191 76 192 77
rect 190 76 191 77
rect 189 76 190 77
rect 172 76 173 77
rect 171 76 172 77
rect 170 76 171 77
rect 169 76 170 77
rect 168 76 169 77
rect 167 76 168 77
rect 111 76 112 77
rect 110 76 111 77
rect 109 76 110 77
rect 108 76 109 77
rect 107 76 108 77
rect 106 76 107 77
rect 105 76 106 77
rect 104 76 105 77
rect 103 76 104 77
rect 102 76 103 77
rect 101 76 102 77
rect 100 76 101 77
rect 99 76 100 77
rect 98 76 99 77
rect 97 76 98 77
rect 96 76 97 77
rect 95 76 96 77
rect 87 76 88 77
rect 86 76 87 77
rect 85 76 86 77
rect 84 76 85 77
rect 83 76 84 77
rect 82 76 83 77
rect 81 76 82 77
rect 80 76 81 77
rect 79 76 80 77
rect 78 76 79 77
rect 77 76 78 77
rect 76 76 77 77
rect 75 76 76 77
rect 74 76 75 77
rect 73 76 74 77
rect 72 76 73 77
rect 71 76 72 77
rect 70 76 71 77
rect 69 76 70 77
rect 68 76 69 77
rect 67 76 68 77
rect 66 76 67 77
rect 65 76 66 77
rect 64 76 65 77
rect 63 76 64 77
rect 62 76 63 77
rect 61 76 62 77
rect 60 76 61 77
rect 59 76 60 77
rect 58 76 59 77
rect 57 76 58 77
rect 56 76 57 77
rect 55 76 56 77
rect 54 76 55 77
rect 27 76 28 77
rect 26 76 27 77
rect 25 76 26 77
rect 24 76 25 77
rect 23 76 24 77
rect 22 76 23 77
rect 21 76 22 77
rect 20 76 21 77
rect 14 76 15 77
rect 13 76 14 77
rect 12 76 13 77
rect 11 76 12 77
rect 10 76 11 77
rect 190 77 191 78
rect 189 77 190 78
rect 174 77 175 78
rect 173 77 174 78
rect 172 77 173 78
rect 171 77 172 78
rect 170 77 171 78
rect 169 77 170 78
rect 168 77 169 78
rect 131 77 132 78
rect 130 77 131 78
rect 129 77 130 78
rect 128 77 129 78
rect 127 77 128 78
rect 126 77 127 78
rect 110 77 111 78
rect 109 77 110 78
rect 108 77 109 78
rect 107 77 108 78
rect 106 77 107 78
rect 105 77 106 78
rect 104 77 105 78
rect 103 77 104 78
rect 102 77 103 78
rect 101 77 102 78
rect 100 77 101 78
rect 99 77 100 78
rect 98 77 99 78
rect 97 77 98 78
rect 96 77 97 78
rect 95 77 96 78
rect 94 77 95 78
rect 86 77 87 78
rect 85 77 86 78
rect 84 77 85 78
rect 83 77 84 78
rect 82 77 83 78
rect 81 77 82 78
rect 80 77 81 78
rect 79 77 80 78
rect 78 77 79 78
rect 77 77 78 78
rect 76 77 77 78
rect 75 77 76 78
rect 74 77 75 78
rect 73 77 74 78
rect 72 77 73 78
rect 71 77 72 78
rect 70 77 71 78
rect 69 77 70 78
rect 68 77 69 78
rect 67 77 68 78
rect 66 77 67 78
rect 65 77 66 78
rect 64 77 65 78
rect 63 77 64 78
rect 62 77 63 78
rect 61 77 62 78
rect 60 77 61 78
rect 59 77 60 78
rect 58 77 59 78
rect 57 77 58 78
rect 56 77 57 78
rect 55 77 56 78
rect 54 77 55 78
rect 53 77 54 78
rect 52 77 53 78
rect 51 77 52 78
rect 26 77 27 78
rect 25 77 26 78
rect 24 77 25 78
rect 23 77 24 78
rect 22 77 23 78
rect 21 77 22 78
rect 20 77 21 78
rect 14 77 15 78
rect 13 77 14 78
rect 12 77 13 78
rect 11 77 12 78
rect 10 77 11 78
rect 175 78 176 79
rect 174 78 175 79
rect 173 78 174 79
rect 172 78 173 79
rect 171 78 172 79
rect 170 78 171 79
rect 135 78 136 79
rect 134 78 135 79
rect 133 78 134 79
rect 132 78 133 79
rect 131 78 132 79
rect 130 78 131 79
rect 129 78 130 79
rect 128 78 129 79
rect 127 78 128 79
rect 126 78 127 79
rect 125 78 126 79
rect 124 78 125 79
rect 123 78 124 79
rect 122 78 123 79
rect 109 78 110 79
rect 108 78 109 79
rect 107 78 108 79
rect 106 78 107 79
rect 105 78 106 79
rect 104 78 105 79
rect 103 78 104 79
rect 102 78 103 79
rect 101 78 102 79
rect 100 78 101 79
rect 99 78 100 79
rect 98 78 99 79
rect 97 78 98 79
rect 96 78 97 79
rect 95 78 96 79
rect 94 78 95 79
rect 85 78 86 79
rect 84 78 85 79
rect 83 78 84 79
rect 82 78 83 79
rect 81 78 82 79
rect 80 78 81 79
rect 79 78 80 79
rect 78 78 79 79
rect 77 78 78 79
rect 76 78 77 79
rect 75 78 76 79
rect 74 78 75 79
rect 73 78 74 79
rect 72 78 73 79
rect 71 78 72 79
rect 70 78 71 79
rect 69 78 70 79
rect 68 78 69 79
rect 67 78 68 79
rect 66 78 67 79
rect 65 78 66 79
rect 64 78 65 79
rect 63 78 64 79
rect 62 78 63 79
rect 61 78 62 79
rect 60 78 61 79
rect 59 78 60 79
rect 58 78 59 79
rect 57 78 58 79
rect 56 78 57 79
rect 55 78 56 79
rect 54 78 55 79
rect 53 78 54 79
rect 52 78 53 79
rect 51 78 52 79
rect 50 78 51 79
rect 49 78 50 79
rect 48 78 49 79
rect 35 78 36 79
rect 34 78 35 79
rect 33 78 34 79
rect 24 78 25 79
rect 23 78 24 79
rect 22 78 23 79
rect 14 78 15 79
rect 13 78 14 79
rect 12 78 13 79
rect 11 78 12 79
rect 10 78 11 79
rect 176 79 177 80
rect 175 79 176 80
rect 174 79 175 80
rect 173 79 174 80
rect 172 79 173 80
rect 171 79 172 80
rect 137 79 138 80
rect 136 79 137 80
rect 135 79 136 80
rect 134 79 135 80
rect 133 79 134 80
rect 132 79 133 80
rect 131 79 132 80
rect 130 79 131 80
rect 129 79 130 80
rect 128 79 129 80
rect 127 79 128 80
rect 126 79 127 80
rect 125 79 126 80
rect 124 79 125 80
rect 123 79 124 80
rect 122 79 123 80
rect 121 79 122 80
rect 120 79 121 80
rect 119 79 120 80
rect 109 79 110 80
rect 108 79 109 80
rect 107 79 108 80
rect 106 79 107 80
rect 105 79 106 80
rect 104 79 105 80
rect 103 79 104 80
rect 102 79 103 80
rect 101 79 102 80
rect 100 79 101 80
rect 99 79 100 80
rect 98 79 99 80
rect 97 79 98 80
rect 96 79 97 80
rect 95 79 96 80
rect 94 79 95 80
rect 93 79 94 80
rect 84 79 85 80
rect 83 79 84 80
rect 82 79 83 80
rect 81 79 82 80
rect 80 79 81 80
rect 79 79 80 80
rect 78 79 79 80
rect 77 79 78 80
rect 76 79 77 80
rect 75 79 76 80
rect 74 79 75 80
rect 73 79 74 80
rect 72 79 73 80
rect 71 79 72 80
rect 70 79 71 80
rect 69 79 70 80
rect 68 79 69 80
rect 67 79 68 80
rect 66 79 67 80
rect 65 79 66 80
rect 64 79 65 80
rect 63 79 64 80
rect 62 79 63 80
rect 61 79 62 80
rect 60 79 61 80
rect 59 79 60 80
rect 58 79 59 80
rect 57 79 58 80
rect 56 79 57 80
rect 55 79 56 80
rect 54 79 55 80
rect 53 79 54 80
rect 52 79 53 80
rect 51 79 52 80
rect 50 79 51 80
rect 49 79 50 80
rect 48 79 49 80
rect 47 79 48 80
rect 46 79 47 80
rect 45 79 46 80
rect 44 79 45 80
rect 43 79 44 80
rect 42 79 43 80
rect 41 79 42 80
rect 40 79 41 80
rect 38 79 39 80
rect 37 79 38 80
rect 36 79 37 80
rect 35 79 36 80
rect 34 79 35 80
rect 33 79 34 80
rect 15 79 16 80
rect 14 79 15 80
rect 13 79 14 80
rect 12 79 13 80
rect 11 79 12 80
rect 10 79 11 80
rect 177 80 178 81
rect 176 80 177 81
rect 175 80 176 81
rect 174 80 175 81
rect 173 80 174 81
rect 172 80 173 81
rect 163 80 164 81
rect 138 80 139 81
rect 137 80 138 81
rect 136 80 137 81
rect 135 80 136 81
rect 134 80 135 81
rect 133 80 134 81
rect 132 80 133 81
rect 131 80 132 81
rect 130 80 131 81
rect 129 80 130 81
rect 128 80 129 81
rect 127 80 128 81
rect 126 80 127 81
rect 125 80 126 81
rect 124 80 125 81
rect 123 80 124 81
rect 122 80 123 81
rect 121 80 122 81
rect 120 80 121 81
rect 119 80 120 81
rect 118 80 119 81
rect 117 80 118 81
rect 108 80 109 81
rect 107 80 108 81
rect 106 80 107 81
rect 105 80 106 81
rect 104 80 105 81
rect 103 80 104 81
rect 102 80 103 81
rect 101 80 102 81
rect 100 80 101 81
rect 99 80 100 81
rect 98 80 99 81
rect 97 80 98 81
rect 96 80 97 81
rect 95 80 96 81
rect 94 80 95 81
rect 93 80 94 81
rect 92 80 93 81
rect 83 80 84 81
rect 82 80 83 81
rect 81 80 82 81
rect 80 80 81 81
rect 79 80 80 81
rect 78 80 79 81
rect 77 80 78 81
rect 76 80 77 81
rect 75 80 76 81
rect 74 80 75 81
rect 73 80 74 81
rect 72 80 73 81
rect 71 80 72 81
rect 70 80 71 81
rect 69 80 70 81
rect 68 80 69 81
rect 67 80 68 81
rect 66 80 67 81
rect 65 80 66 81
rect 64 80 65 81
rect 63 80 64 81
rect 62 80 63 81
rect 61 80 62 81
rect 60 80 61 81
rect 59 80 60 81
rect 58 80 59 81
rect 57 80 58 81
rect 56 80 57 81
rect 55 80 56 81
rect 54 80 55 81
rect 53 80 54 81
rect 52 80 53 81
rect 51 80 52 81
rect 50 80 51 81
rect 49 80 50 81
rect 48 80 49 81
rect 47 80 48 81
rect 46 80 47 81
rect 45 80 46 81
rect 44 80 45 81
rect 43 80 44 81
rect 42 80 43 81
rect 41 80 42 81
rect 40 80 41 81
rect 39 80 40 81
rect 38 80 39 81
rect 37 80 38 81
rect 36 80 37 81
rect 35 80 36 81
rect 34 80 35 81
rect 33 80 34 81
rect 15 80 16 81
rect 14 80 15 81
rect 13 80 14 81
rect 12 80 13 81
rect 11 80 12 81
rect 10 80 11 81
rect 179 81 180 82
rect 178 81 179 82
rect 177 81 178 82
rect 176 81 177 82
rect 175 81 176 82
rect 174 81 175 82
rect 173 81 174 82
rect 163 81 164 82
rect 140 81 141 82
rect 139 81 140 82
rect 138 81 139 82
rect 137 81 138 82
rect 136 81 137 82
rect 135 81 136 82
rect 134 81 135 82
rect 133 81 134 82
rect 132 81 133 82
rect 131 81 132 82
rect 130 81 131 82
rect 129 81 130 82
rect 128 81 129 82
rect 127 81 128 82
rect 126 81 127 82
rect 125 81 126 82
rect 124 81 125 82
rect 123 81 124 82
rect 122 81 123 82
rect 121 81 122 82
rect 120 81 121 82
rect 119 81 120 82
rect 118 81 119 82
rect 117 81 118 82
rect 116 81 117 82
rect 115 81 116 82
rect 107 81 108 82
rect 106 81 107 82
rect 105 81 106 82
rect 104 81 105 82
rect 103 81 104 82
rect 102 81 103 82
rect 101 81 102 82
rect 100 81 101 82
rect 99 81 100 82
rect 98 81 99 82
rect 97 81 98 82
rect 96 81 97 82
rect 95 81 96 82
rect 94 81 95 82
rect 93 81 94 82
rect 92 81 93 82
rect 82 81 83 82
rect 81 81 82 82
rect 80 81 81 82
rect 79 81 80 82
rect 78 81 79 82
rect 77 81 78 82
rect 76 81 77 82
rect 75 81 76 82
rect 74 81 75 82
rect 73 81 74 82
rect 72 81 73 82
rect 71 81 72 82
rect 70 81 71 82
rect 69 81 70 82
rect 68 81 69 82
rect 67 81 68 82
rect 66 81 67 82
rect 65 81 66 82
rect 64 81 65 82
rect 63 81 64 82
rect 62 81 63 82
rect 61 81 62 82
rect 60 81 61 82
rect 59 81 60 82
rect 58 81 59 82
rect 57 81 58 82
rect 56 81 57 82
rect 55 81 56 82
rect 54 81 55 82
rect 53 81 54 82
rect 52 81 53 82
rect 51 81 52 82
rect 50 81 51 82
rect 49 81 50 82
rect 48 81 49 82
rect 47 81 48 82
rect 46 81 47 82
rect 45 81 46 82
rect 44 81 45 82
rect 43 81 44 82
rect 42 81 43 82
rect 41 81 42 82
rect 40 81 41 82
rect 39 81 40 82
rect 38 81 39 82
rect 37 81 38 82
rect 36 81 37 82
rect 35 81 36 82
rect 34 81 35 82
rect 33 81 34 82
rect 16 81 17 82
rect 15 81 16 82
rect 14 81 15 82
rect 13 81 14 82
rect 12 81 13 82
rect 11 81 12 82
rect 10 81 11 82
rect 197 82 198 83
rect 196 82 197 83
rect 189 82 190 83
rect 180 82 181 83
rect 179 82 180 83
rect 178 82 179 83
rect 177 82 178 83
rect 176 82 177 83
rect 175 82 176 83
rect 174 82 175 83
rect 164 82 165 83
rect 163 82 164 83
rect 141 82 142 83
rect 140 82 141 83
rect 139 82 140 83
rect 138 82 139 83
rect 137 82 138 83
rect 136 82 137 83
rect 135 82 136 83
rect 134 82 135 83
rect 133 82 134 83
rect 132 82 133 83
rect 131 82 132 83
rect 130 82 131 83
rect 129 82 130 83
rect 128 82 129 83
rect 127 82 128 83
rect 126 82 127 83
rect 125 82 126 83
rect 124 82 125 83
rect 123 82 124 83
rect 122 82 123 83
rect 121 82 122 83
rect 120 82 121 83
rect 119 82 120 83
rect 118 82 119 83
rect 117 82 118 83
rect 116 82 117 83
rect 115 82 116 83
rect 114 82 115 83
rect 107 82 108 83
rect 106 82 107 83
rect 105 82 106 83
rect 104 82 105 83
rect 103 82 104 83
rect 102 82 103 83
rect 101 82 102 83
rect 100 82 101 83
rect 99 82 100 83
rect 98 82 99 83
rect 97 82 98 83
rect 96 82 97 83
rect 95 82 96 83
rect 94 82 95 83
rect 93 82 94 83
rect 92 82 93 83
rect 91 82 92 83
rect 81 82 82 83
rect 80 82 81 83
rect 79 82 80 83
rect 78 82 79 83
rect 77 82 78 83
rect 76 82 77 83
rect 75 82 76 83
rect 74 82 75 83
rect 73 82 74 83
rect 72 82 73 83
rect 71 82 72 83
rect 70 82 71 83
rect 69 82 70 83
rect 68 82 69 83
rect 67 82 68 83
rect 66 82 67 83
rect 65 82 66 83
rect 64 82 65 83
rect 63 82 64 83
rect 62 82 63 83
rect 61 82 62 83
rect 60 82 61 83
rect 59 82 60 83
rect 58 82 59 83
rect 57 82 58 83
rect 56 82 57 83
rect 55 82 56 83
rect 54 82 55 83
rect 53 82 54 83
rect 52 82 53 83
rect 51 82 52 83
rect 50 82 51 83
rect 49 82 50 83
rect 48 82 49 83
rect 47 82 48 83
rect 46 82 47 83
rect 45 82 46 83
rect 44 82 45 83
rect 43 82 44 83
rect 42 82 43 83
rect 41 82 42 83
rect 40 82 41 83
rect 39 82 40 83
rect 38 82 39 83
rect 37 82 38 83
rect 36 82 37 83
rect 35 82 36 83
rect 34 82 35 83
rect 33 82 34 83
rect 16 82 17 83
rect 15 82 16 83
rect 14 82 15 83
rect 13 82 14 83
rect 12 82 13 83
rect 11 82 12 83
rect 10 82 11 83
rect 196 83 197 84
rect 195 83 196 84
rect 194 83 195 84
rect 193 83 194 84
rect 192 83 193 84
rect 191 83 192 84
rect 190 83 191 84
rect 189 83 190 84
rect 181 83 182 84
rect 180 83 181 84
rect 179 83 180 84
rect 178 83 179 84
rect 177 83 178 84
rect 176 83 177 84
rect 175 83 176 84
rect 174 83 175 84
rect 173 83 174 84
rect 172 83 173 84
rect 171 83 172 84
rect 170 83 171 84
rect 169 83 170 84
rect 168 83 169 84
rect 167 83 168 84
rect 166 83 167 84
rect 165 83 166 84
rect 164 83 165 84
rect 163 83 164 84
rect 142 83 143 84
rect 141 83 142 84
rect 140 83 141 84
rect 139 83 140 84
rect 138 83 139 84
rect 137 83 138 84
rect 136 83 137 84
rect 135 83 136 84
rect 134 83 135 84
rect 133 83 134 84
rect 132 83 133 84
rect 131 83 132 84
rect 130 83 131 84
rect 129 83 130 84
rect 128 83 129 84
rect 127 83 128 84
rect 126 83 127 84
rect 125 83 126 84
rect 124 83 125 84
rect 123 83 124 84
rect 122 83 123 84
rect 121 83 122 84
rect 120 83 121 84
rect 119 83 120 84
rect 118 83 119 84
rect 117 83 118 84
rect 116 83 117 84
rect 115 83 116 84
rect 114 83 115 84
rect 113 83 114 84
rect 106 83 107 84
rect 105 83 106 84
rect 104 83 105 84
rect 103 83 104 84
rect 102 83 103 84
rect 101 83 102 84
rect 100 83 101 84
rect 99 83 100 84
rect 98 83 99 84
rect 97 83 98 84
rect 96 83 97 84
rect 95 83 96 84
rect 94 83 95 84
rect 93 83 94 84
rect 92 83 93 84
rect 91 83 92 84
rect 90 83 91 84
rect 80 83 81 84
rect 79 83 80 84
rect 78 83 79 84
rect 77 83 78 84
rect 76 83 77 84
rect 75 83 76 84
rect 74 83 75 84
rect 73 83 74 84
rect 72 83 73 84
rect 71 83 72 84
rect 70 83 71 84
rect 69 83 70 84
rect 68 83 69 84
rect 67 83 68 84
rect 66 83 67 84
rect 65 83 66 84
rect 64 83 65 84
rect 63 83 64 84
rect 62 83 63 84
rect 61 83 62 84
rect 60 83 61 84
rect 59 83 60 84
rect 58 83 59 84
rect 57 83 58 84
rect 56 83 57 84
rect 55 83 56 84
rect 54 83 55 84
rect 53 83 54 84
rect 52 83 53 84
rect 51 83 52 84
rect 50 83 51 84
rect 49 83 50 84
rect 48 83 49 84
rect 47 83 48 84
rect 46 83 47 84
rect 45 83 46 84
rect 44 83 45 84
rect 43 83 44 84
rect 42 83 43 84
rect 41 83 42 84
rect 40 83 41 84
rect 39 83 40 84
rect 38 83 39 84
rect 37 83 38 84
rect 36 83 37 84
rect 35 83 36 84
rect 34 83 35 84
rect 33 83 34 84
rect 25 83 26 84
rect 24 83 25 84
rect 23 83 24 84
rect 17 83 18 84
rect 16 83 17 84
rect 15 83 16 84
rect 14 83 15 84
rect 13 83 14 84
rect 12 83 13 84
rect 11 83 12 84
rect 10 83 11 84
rect 197 84 198 85
rect 196 84 197 85
rect 195 84 196 85
rect 194 84 195 85
rect 193 84 194 85
rect 192 84 193 85
rect 191 84 192 85
rect 190 84 191 85
rect 189 84 190 85
rect 180 84 181 85
rect 179 84 180 85
rect 178 84 179 85
rect 177 84 178 85
rect 176 84 177 85
rect 175 84 176 85
rect 174 84 175 85
rect 173 84 174 85
rect 172 84 173 85
rect 171 84 172 85
rect 170 84 171 85
rect 169 84 170 85
rect 168 84 169 85
rect 167 84 168 85
rect 166 84 167 85
rect 165 84 166 85
rect 164 84 165 85
rect 163 84 164 85
rect 143 84 144 85
rect 142 84 143 85
rect 141 84 142 85
rect 140 84 141 85
rect 139 84 140 85
rect 138 84 139 85
rect 137 84 138 85
rect 136 84 137 85
rect 135 84 136 85
rect 134 84 135 85
rect 133 84 134 85
rect 132 84 133 85
rect 131 84 132 85
rect 130 84 131 85
rect 129 84 130 85
rect 128 84 129 85
rect 127 84 128 85
rect 126 84 127 85
rect 125 84 126 85
rect 124 84 125 85
rect 123 84 124 85
rect 122 84 123 85
rect 121 84 122 85
rect 120 84 121 85
rect 119 84 120 85
rect 118 84 119 85
rect 117 84 118 85
rect 116 84 117 85
rect 115 84 116 85
rect 114 84 115 85
rect 113 84 114 85
rect 112 84 113 85
rect 111 84 112 85
rect 106 84 107 85
rect 105 84 106 85
rect 104 84 105 85
rect 103 84 104 85
rect 102 84 103 85
rect 101 84 102 85
rect 100 84 101 85
rect 99 84 100 85
rect 98 84 99 85
rect 97 84 98 85
rect 96 84 97 85
rect 95 84 96 85
rect 94 84 95 85
rect 93 84 94 85
rect 92 84 93 85
rect 91 84 92 85
rect 90 84 91 85
rect 79 84 80 85
rect 78 84 79 85
rect 77 84 78 85
rect 76 84 77 85
rect 75 84 76 85
rect 74 84 75 85
rect 73 84 74 85
rect 72 84 73 85
rect 71 84 72 85
rect 70 84 71 85
rect 69 84 70 85
rect 68 84 69 85
rect 67 84 68 85
rect 66 84 67 85
rect 65 84 66 85
rect 64 84 65 85
rect 63 84 64 85
rect 62 84 63 85
rect 61 84 62 85
rect 60 84 61 85
rect 59 84 60 85
rect 58 84 59 85
rect 57 84 58 85
rect 56 84 57 85
rect 55 84 56 85
rect 54 84 55 85
rect 53 84 54 85
rect 52 84 53 85
rect 51 84 52 85
rect 50 84 51 85
rect 49 84 50 85
rect 48 84 49 85
rect 47 84 48 85
rect 46 84 47 85
rect 45 84 46 85
rect 44 84 45 85
rect 43 84 44 85
rect 42 84 43 85
rect 41 84 42 85
rect 40 84 41 85
rect 39 84 40 85
rect 38 84 39 85
rect 37 84 38 85
rect 36 84 37 85
rect 35 84 36 85
rect 34 84 35 85
rect 33 84 34 85
rect 26 84 27 85
rect 25 84 26 85
rect 24 84 25 85
rect 23 84 24 85
rect 22 84 23 85
rect 21 84 22 85
rect 20 84 21 85
rect 19 84 20 85
rect 18 84 19 85
rect 17 84 18 85
rect 16 84 17 85
rect 15 84 16 85
rect 14 84 15 85
rect 13 84 14 85
rect 12 84 13 85
rect 11 84 12 85
rect 10 84 11 85
rect 197 85 198 86
rect 193 85 194 86
rect 192 85 193 86
rect 164 85 165 86
rect 163 85 164 86
rect 144 85 145 86
rect 143 85 144 86
rect 142 85 143 86
rect 141 85 142 86
rect 140 85 141 86
rect 139 85 140 86
rect 138 85 139 86
rect 137 85 138 86
rect 136 85 137 86
rect 135 85 136 86
rect 134 85 135 86
rect 133 85 134 86
rect 132 85 133 86
rect 131 85 132 86
rect 130 85 131 86
rect 129 85 130 86
rect 128 85 129 86
rect 127 85 128 86
rect 126 85 127 86
rect 125 85 126 86
rect 124 85 125 86
rect 123 85 124 86
rect 122 85 123 86
rect 121 85 122 86
rect 120 85 121 86
rect 119 85 120 86
rect 118 85 119 86
rect 117 85 118 86
rect 116 85 117 86
rect 115 85 116 86
rect 114 85 115 86
rect 113 85 114 86
rect 112 85 113 86
rect 111 85 112 86
rect 110 85 111 86
rect 105 85 106 86
rect 104 85 105 86
rect 103 85 104 86
rect 102 85 103 86
rect 101 85 102 86
rect 100 85 101 86
rect 99 85 100 86
rect 98 85 99 86
rect 97 85 98 86
rect 96 85 97 86
rect 95 85 96 86
rect 94 85 95 86
rect 93 85 94 86
rect 92 85 93 86
rect 91 85 92 86
rect 90 85 91 86
rect 89 85 90 86
rect 78 85 79 86
rect 77 85 78 86
rect 76 85 77 86
rect 75 85 76 86
rect 74 85 75 86
rect 73 85 74 86
rect 72 85 73 86
rect 71 85 72 86
rect 70 85 71 86
rect 69 85 70 86
rect 68 85 69 86
rect 67 85 68 86
rect 66 85 67 86
rect 65 85 66 86
rect 64 85 65 86
rect 63 85 64 86
rect 62 85 63 86
rect 61 85 62 86
rect 60 85 61 86
rect 59 85 60 86
rect 58 85 59 86
rect 57 85 58 86
rect 56 85 57 86
rect 55 85 56 86
rect 54 85 55 86
rect 53 85 54 86
rect 52 85 53 86
rect 51 85 52 86
rect 50 85 51 86
rect 49 85 50 86
rect 48 85 49 86
rect 47 85 48 86
rect 46 85 47 86
rect 45 85 46 86
rect 44 85 45 86
rect 43 85 44 86
rect 42 85 43 86
rect 41 85 42 86
rect 40 85 41 86
rect 39 85 40 86
rect 38 85 39 86
rect 37 85 38 86
rect 36 85 37 86
rect 35 85 36 86
rect 34 85 35 86
rect 27 85 28 86
rect 26 85 27 86
rect 25 85 26 86
rect 24 85 25 86
rect 23 85 24 86
rect 22 85 23 86
rect 21 85 22 86
rect 20 85 21 86
rect 19 85 20 86
rect 18 85 19 86
rect 17 85 18 86
rect 16 85 17 86
rect 15 85 16 86
rect 14 85 15 86
rect 13 85 14 86
rect 12 85 13 86
rect 11 85 12 86
rect 10 85 11 86
rect 193 86 194 87
rect 192 86 193 87
rect 189 86 190 87
rect 163 86 164 87
rect 145 86 146 87
rect 144 86 145 87
rect 143 86 144 87
rect 142 86 143 87
rect 141 86 142 87
rect 140 86 141 87
rect 139 86 140 87
rect 138 86 139 87
rect 137 86 138 87
rect 136 86 137 87
rect 135 86 136 87
rect 134 86 135 87
rect 133 86 134 87
rect 132 86 133 87
rect 131 86 132 87
rect 130 86 131 87
rect 129 86 130 87
rect 128 86 129 87
rect 127 86 128 87
rect 126 86 127 87
rect 125 86 126 87
rect 124 86 125 87
rect 123 86 124 87
rect 122 86 123 87
rect 121 86 122 87
rect 120 86 121 87
rect 119 86 120 87
rect 118 86 119 87
rect 117 86 118 87
rect 116 86 117 87
rect 115 86 116 87
rect 114 86 115 87
rect 113 86 114 87
rect 112 86 113 87
rect 111 86 112 87
rect 110 86 111 87
rect 109 86 110 87
rect 108 86 109 87
rect 104 86 105 87
rect 103 86 104 87
rect 102 86 103 87
rect 101 86 102 87
rect 100 86 101 87
rect 99 86 100 87
rect 98 86 99 87
rect 97 86 98 87
rect 96 86 97 87
rect 95 86 96 87
rect 94 86 95 87
rect 93 86 94 87
rect 92 86 93 87
rect 91 86 92 87
rect 90 86 91 87
rect 89 86 90 87
rect 88 86 89 87
rect 77 86 78 87
rect 76 86 77 87
rect 75 86 76 87
rect 74 86 75 87
rect 73 86 74 87
rect 72 86 73 87
rect 71 86 72 87
rect 70 86 71 87
rect 69 86 70 87
rect 68 86 69 87
rect 67 86 68 87
rect 66 86 67 87
rect 65 86 66 87
rect 64 86 65 87
rect 63 86 64 87
rect 62 86 63 87
rect 61 86 62 87
rect 60 86 61 87
rect 59 86 60 87
rect 58 86 59 87
rect 57 86 58 87
rect 56 86 57 87
rect 55 86 56 87
rect 54 86 55 87
rect 53 86 54 87
rect 52 86 53 87
rect 51 86 52 87
rect 50 86 51 87
rect 49 86 50 87
rect 48 86 49 87
rect 47 86 48 87
rect 46 86 47 87
rect 45 86 46 87
rect 44 86 45 87
rect 43 86 44 87
rect 42 86 43 87
rect 41 86 42 87
rect 40 86 41 87
rect 39 86 40 87
rect 38 86 39 87
rect 37 86 38 87
rect 36 86 37 87
rect 35 86 36 87
rect 34 86 35 87
rect 27 86 28 87
rect 26 86 27 87
rect 25 86 26 87
rect 24 86 25 87
rect 23 86 24 87
rect 22 86 23 87
rect 21 86 22 87
rect 20 86 21 87
rect 19 86 20 87
rect 18 86 19 87
rect 17 86 18 87
rect 16 86 17 87
rect 15 86 16 87
rect 14 86 15 87
rect 13 86 14 87
rect 12 86 13 87
rect 11 86 12 87
rect 10 86 11 87
rect 197 87 198 88
rect 196 87 197 88
rect 193 87 194 88
rect 192 87 193 88
rect 190 87 191 88
rect 189 87 190 88
rect 146 87 147 88
rect 145 87 146 88
rect 144 87 145 88
rect 143 87 144 88
rect 142 87 143 88
rect 141 87 142 88
rect 140 87 141 88
rect 139 87 140 88
rect 138 87 139 88
rect 137 87 138 88
rect 136 87 137 88
rect 135 87 136 88
rect 134 87 135 88
rect 133 87 134 88
rect 132 87 133 88
rect 131 87 132 88
rect 130 87 131 88
rect 129 87 130 88
rect 128 87 129 88
rect 127 87 128 88
rect 126 87 127 88
rect 125 87 126 88
rect 124 87 125 88
rect 123 87 124 88
rect 122 87 123 88
rect 121 87 122 88
rect 120 87 121 88
rect 119 87 120 88
rect 118 87 119 88
rect 117 87 118 88
rect 116 87 117 88
rect 115 87 116 88
rect 114 87 115 88
rect 113 87 114 88
rect 112 87 113 88
rect 111 87 112 88
rect 110 87 111 88
rect 109 87 110 88
rect 108 87 109 88
rect 107 87 108 88
rect 104 87 105 88
rect 103 87 104 88
rect 102 87 103 88
rect 101 87 102 88
rect 100 87 101 88
rect 99 87 100 88
rect 98 87 99 88
rect 97 87 98 88
rect 96 87 97 88
rect 95 87 96 88
rect 94 87 95 88
rect 93 87 94 88
rect 92 87 93 88
rect 91 87 92 88
rect 90 87 91 88
rect 89 87 90 88
rect 88 87 89 88
rect 87 87 88 88
rect 75 87 76 88
rect 74 87 75 88
rect 73 87 74 88
rect 72 87 73 88
rect 71 87 72 88
rect 70 87 71 88
rect 69 87 70 88
rect 68 87 69 88
rect 67 87 68 88
rect 66 87 67 88
rect 65 87 66 88
rect 64 87 65 88
rect 63 87 64 88
rect 62 87 63 88
rect 61 87 62 88
rect 60 87 61 88
rect 59 87 60 88
rect 58 87 59 88
rect 57 87 58 88
rect 56 87 57 88
rect 55 87 56 88
rect 54 87 55 88
rect 53 87 54 88
rect 52 87 53 88
rect 51 87 52 88
rect 50 87 51 88
rect 49 87 50 88
rect 48 87 49 88
rect 47 87 48 88
rect 46 87 47 88
rect 45 87 46 88
rect 44 87 45 88
rect 43 87 44 88
rect 42 87 43 88
rect 41 87 42 88
rect 40 87 41 88
rect 39 87 40 88
rect 38 87 39 88
rect 37 87 38 88
rect 36 87 37 88
rect 35 87 36 88
rect 28 87 29 88
rect 27 87 28 88
rect 26 87 27 88
rect 25 87 26 88
rect 24 87 25 88
rect 23 87 24 88
rect 22 87 23 88
rect 21 87 22 88
rect 20 87 21 88
rect 19 87 20 88
rect 18 87 19 88
rect 17 87 18 88
rect 16 87 17 88
rect 15 87 16 88
rect 14 87 15 88
rect 13 87 14 88
rect 12 87 13 88
rect 11 87 12 88
rect 10 87 11 88
rect 9 87 10 88
rect 196 88 197 89
rect 195 88 196 89
rect 190 88 191 89
rect 173 88 174 89
rect 172 88 173 89
rect 171 88 172 89
rect 170 88 171 89
rect 146 88 147 89
rect 145 88 146 89
rect 144 88 145 89
rect 143 88 144 89
rect 142 88 143 89
rect 141 88 142 89
rect 140 88 141 89
rect 139 88 140 89
rect 138 88 139 89
rect 137 88 138 89
rect 136 88 137 89
rect 135 88 136 89
rect 134 88 135 89
rect 133 88 134 89
rect 132 88 133 89
rect 131 88 132 89
rect 130 88 131 89
rect 129 88 130 89
rect 128 88 129 89
rect 127 88 128 89
rect 126 88 127 89
rect 125 88 126 89
rect 124 88 125 89
rect 123 88 124 89
rect 122 88 123 89
rect 121 88 122 89
rect 120 88 121 89
rect 119 88 120 89
rect 118 88 119 89
rect 117 88 118 89
rect 116 88 117 89
rect 115 88 116 89
rect 114 88 115 89
rect 113 88 114 89
rect 112 88 113 89
rect 111 88 112 89
rect 110 88 111 89
rect 109 88 110 89
rect 108 88 109 89
rect 107 88 108 89
rect 106 88 107 89
rect 105 88 106 89
rect 104 88 105 89
rect 103 88 104 89
rect 102 88 103 89
rect 101 88 102 89
rect 100 88 101 89
rect 99 88 100 89
rect 98 88 99 89
rect 97 88 98 89
rect 96 88 97 89
rect 95 88 96 89
rect 94 88 95 89
rect 93 88 94 89
rect 92 88 93 89
rect 91 88 92 89
rect 90 88 91 89
rect 89 88 90 89
rect 88 88 89 89
rect 87 88 88 89
rect 86 88 87 89
rect 73 88 74 89
rect 72 88 73 89
rect 71 88 72 89
rect 70 88 71 89
rect 69 88 70 89
rect 68 88 69 89
rect 67 88 68 89
rect 66 88 67 89
rect 65 88 66 89
rect 64 88 65 89
rect 63 88 64 89
rect 62 88 63 89
rect 61 88 62 89
rect 60 88 61 89
rect 59 88 60 89
rect 58 88 59 89
rect 57 88 58 89
rect 56 88 57 89
rect 55 88 56 89
rect 54 88 55 89
rect 53 88 54 89
rect 52 88 53 89
rect 51 88 52 89
rect 50 88 51 89
rect 49 88 50 89
rect 48 88 49 89
rect 47 88 48 89
rect 46 88 47 89
rect 45 88 46 89
rect 44 88 45 89
rect 43 88 44 89
rect 42 88 43 89
rect 41 88 42 89
rect 40 88 41 89
rect 39 88 40 89
rect 38 88 39 89
rect 37 88 38 89
rect 36 88 37 89
rect 29 88 30 89
rect 28 88 29 89
rect 27 88 28 89
rect 26 88 27 89
rect 25 88 26 89
rect 24 88 25 89
rect 23 88 24 89
rect 22 88 23 89
rect 21 88 22 89
rect 20 88 21 89
rect 19 88 20 89
rect 18 88 19 89
rect 17 88 18 89
rect 16 88 17 89
rect 15 88 16 89
rect 14 88 15 89
rect 13 88 14 89
rect 12 88 13 89
rect 11 88 12 89
rect 10 88 11 89
rect 9 88 10 89
rect 176 89 177 90
rect 175 89 176 90
rect 174 89 175 90
rect 173 89 174 90
rect 172 89 173 90
rect 171 89 172 90
rect 170 89 171 90
rect 169 89 170 90
rect 168 89 169 90
rect 167 89 168 90
rect 147 89 148 90
rect 146 89 147 90
rect 145 89 146 90
rect 144 89 145 90
rect 143 89 144 90
rect 142 89 143 90
rect 141 89 142 90
rect 140 89 141 90
rect 139 89 140 90
rect 138 89 139 90
rect 137 89 138 90
rect 136 89 137 90
rect 135 89 136 90
rect 134 89 135 90
rect 133 89 134 90
rect 132 89 133 90
rect 131 89 132 90
rect 130 89 131 90
rect 129 89 130 90
rect 128 89 129 90
rect 127 89 128 90
rect 126 89 127 90
rect 125 89 126 90
rect 124 89 125 90
rect 123 89 124 90
rect 122 89 123 90
rect 121 89 122 90
rect 120 89 121 90
rect 119 89 120 90
rect 118 89 119 90
rect 117 89 118 90
rect 116 89 117 90
rect 115 89 116 90
rect 114 89 115 90
rect 113 89 114 90
rect 112 89 113 90
rect 111 89 112 90
rect 110 89 111 90
rect 109 89 110 90
rect 108 89 109 90
rect 107 89 108 90
rect 106 89 107 90
rect 105 89 106 90
rect 104 89 105 90
rect 103 89 104 90
rect 102 89 103 90
rect 101 89 102 90
rect 100 89 101 90
rect 99 89 100 90
rect 98 89 99 90
rect 97 89 98 90
rect 96 89 97 90
rect 95 89 96 90
rect 94 89 95 90
rect 93 89 94 90
rect 92 89 93 90
rect 91 89 92 90
rect 90 89 91 90
rect 89 89 90 90
rect 88 89 89 90
rect 87 89 88 90
rect 86 89 87 90
rect 85 89 86 90
rect 71 89 72 90
rect 70 89 71 90
rect 69 89 70 90
rect 68 89 69 90
rect 67 89 68 90
rect 66 89 67 90
rect 65 89 66 90
rect 64 89 65 90
rect 63 89 64 90
rect 62 89 63 90
rect 61 89 62 90
rect 60 89 61 90
rect 59 89 60 90
rect 58 89 59 90
rect 57 89 58 90
rect 56 89 57 90
rect 55 89 56 90
rect 54 89 55 90
rect 53 89 54 90
rect 52 89 53 90
rect 51 89 52 90
rect 50 89 51 90
rect 49 89 50 90
rect 48 89 49 90
rect 47 89 48 90
rect 46 89 47 90
rect 45 89 46 90
rect 44 89 45 90
rect 43 89 44 90
rect 42 89 43 90
rect 41 89 42 90
rect 40 89 41 90
rect 39 89 40 90
rect 38 89 39 90
rect 29 89 30 90
rect 28 89 29 90
rect 27 89 28 90
rect 26 89 27 90
rect 25 89 26 90
rect 24 89 25 90
rect 23 89 24 90
rect 22 89 23 90
rect 21 89 22 90
rect 20 89 21 90
rect 19 89 20 90
rect 18 89 19 90
rect 17 89 18 90
rect 16 89 17 90
rect 15 89 16 90
rect 14 89 15 90
rect 13 89 14 90
rect 12 89 13 90
rect 11 89 12 90
rect 10 89 11 90
rect 9 89 10 90
rect 177 90 178 91
rect 176 90 177 91
rect 175 90 176 91
rect 174 90 175 91
rect 173 90 174 91
rect 172 90 173 91
rect 171 90 172 91
rect 170 90 171 91
rect 169 90 170 91
rect 168 90 169 91
rect 167 90 168 91
rect 166 90 167 91
rect 147 90 148 91
rect 146 90 147 91
rect 145 90 146 91
rect 144 90 145 91
rect 143 90 144 91
rect 142 90 143 91
rect 141 90 142 91
rect 140 90 141 91
rect 139 90 140 91
rect 138 90 139 91
rect 137 90 138 91
rect 136 90 137 91
rect 135 90 136 91
rect 134 90 135 91
rect 133 90 134 91
rect 132 90 133 91
rect 131 90 132 91
rect 130 90 131 91
rect 129 90 130 91
rect 128 90 129 91
rect 127 90 128 91
rect 126 90 127 91
rect 125 90 126 91
rect 124 90 125 91
rect 123 90 124 91
rect 122 90 123 91
rect 121 90 122 91
rect 120 90 121 91
rect 119 90 120 91
rect 118 90 119 91
rect 117 90 118 91
rect 116 90 117 91
rect 115 90 116 91
rect 114 90 115 91
rect 113 90 114 91
rect 112 90 113 91
rect 111 90 112 91
rect 110 90 111 91
rect 109 90 110 91
rect 108 90 109 91
rect 107 90 108 91
rect 106 90 107 91
rect 105 90 106 91
rect 104 90 105 91
rect 103 90 104 91
rect 102 90 103 91
rect 101 90 102 91
rect 100 90 101 91
rect 99 90 100 91
rect 98 90 99 91
rect 97 90 98 91
rect 96 90 97 91
rect 95 90 96 91
rect 94 90 95 91
rect 93 90 94 91
rect 92 90 93 91
rect 91 90 92 91
rect 90 90 91 91
rect 89 90 90 91
rect 88 90 89 91
rect 87 90 88 91
rect 86 90 87 91
rect 85 90 86 91
rect 84 90 85 91
rect 83 90 84 91
rect 68 90 69 91
rect 67 90 68 91
rect 66 90 67 91
rect 65 90 66 91
rect 64 90 65 91
rect 63 90 64 91
rect 62 90 63 91
rect 61 90 62 91
rect 60 90 61 91
rect 59 90 60 91
rect 58 90 59 91
rect 57 90 58 91
rect 56 90 57 91
rect 55 90 56 91
rect 54 90 55 91
rect 53 90 54 91
rect 52 90 53 91
rect 51 90 52 91
rect 50 90 51 91
rect 49 90 50 91
rect 48 90 49 91
rect 47 90 48 91
rect 46 90 47 91
rect 45 90 46 91
rect 44 90 45 91
rect 43 90 44 91
rect 42 90 43 91
rect 41 90 42 91
rect 40 90 41 91
rect 39 90 40 91
rect 30 90 31 91
rect 29 90 30 91
rect 28 90 29 91
rect 27 90 28 91
rect 26 90 27 91
rect 25 90 26 91
rect 24 90 25 91
rect 23 90 24 91
rect 22 90 23 91
rect 21 90 22 91
rect 20 90 21 91
rect 19 90 20 91
rect 18 90 19 91
rect 17 90 18 91
rect 16 90 17 91
rect 15 90 16 91
rect 14 90 15 91
rect 13 90 14 91
rect 12 90 13 91
rect 11 90 12 91
rect 10 90 11 91
rect 9 90 10 91
rect 178 91 179 92
rect 177 91 178 92
rect 176 91 177 92
rect 175 91 176 92
rect 174 91 175 92
rect 173 91 174 92
rect 172 91 173 92
rect 171 91 172 92
rect 170 91 171 92
rect 169 91 170 92
rect 168 91 169 92
rect 167 91 168 92
rect 166 91 167 92
rect 165 91 166 92
rect 148 91 149 92
rect 147 91 148 92
rect 146 91 147 92
rect 145 91 146 92
rect 144 91 145 92
rect 143 91 144 92
rect 142 91 143 92
rect 141 91 142 92
rect 140 91 141 92
rect 139 91 140 92
rect 138 91 139 92
rect 137 91 138 92
rect 136 91 137 92
rect 135 91 136 92
rect 134 91 135 92
rect 133 91 134 92
rect 132 91 133 92
rect 131 91 132 92
rect 130 91 131 92
rect 129 91 130 92
rect 128 91 129 92
rect 127 91 128 92
rect 126 91 127 92
rect 125 91 126 92
rect 124 91 125 92
rect 123 91 124 92
rect 122 91 123 92
rect 121 91 122 92
rect 120 91 121 92
rect 119 91 120 92
rect 118 91 119 92
rect 117 91 118 92
rect 116 91 117 92
rect 115 91 116 92
rect 114 91 115 92
rect 113 91 114 92
rect 112 91 113 92
rect 111 91 112 92
rect 110 91 111 92
rect 109 91 110 92
rect 108 91 109 92
rect 107 91 108 92
rect 106 91 107 92
rect 105 91 106 92
rect 104 91 105 92
rect 103 91 104 92
rect 102 91 103 92
rect 101 91 102 92
rect 100 91 101 92
rect 99 91 100 92
rect 98 91 99 92
rect 97 91 98 92
rect 96 91 97 92
rect 95 91 96 92
rect 94 91 95 92
rect 93 91 94 92
rect 92 91 93 92
rect 91 91 92 92
rect 90 91 91 92
rect 89 91 90 92
rect 88 91 89 92
rect 87 91 88 92
rect 86 91 87 92
rect 85 91 86 92
rect 84 91 85 92
rect 83 91 84 92
rect 82 91 83 92
rect 65 91 66 92
rect 64 91 65 92
rect 63 91 64 92
rect 62 91 63 92
rect 61 91 62 92
rect 60 91 61 92
rect 59 91 60 92
rect 58 91 59 92
rect 57 91 58 92
rect 56 91 57 92
rect 55 91 56 92
rect 54 91 55 92
rect 53 91 54 92
rect 52 91 53 92
rect 51 91 52 92
rect 50 91 51 92
rect 49 91 50 92
rect 48 91 49 92
rect 47 91 48 92
rect 46 91 47 92
rect 45 91 46 92
rect 44 91 45 92
rect 43 91 44 92
rect 42 91 43 92
rect 41 91 42 92
rect 31 91 32 92
rect 30 91 31 92
rect 29 91 30 92
rect 28 91 29 92
rect 27 91 28 92
rect 26 91 27 92
rect 25 91 26 92
rect 24 91 25 92
rect 23 91 24 92
rect 22 91 23 92
rect 21 91 22 92
rect 20 91 21 92
rect 19 91 20 92
rect 18 91 19 92
rect 17 91 18 92
rect 16 91 17 92
rect 15 91 16 92
rect 14 91 15 92
rect 13 91 14 92
rect 12 91 13 92
rect 11 91 12 92
rect 10 91 11 92
rect 9 91 10 92
rect 8 91 9 92
rect 189 92 190 93
rect 179 92 180 93
rect 178 92 179 93
rect 177 92 178 93
rect 176 92 177 93
rect 175 92 176 93
rect 174 92 175 93
rect 173 92 174 93
rect 172 92 173 93
rect 171 92 172 93
rect 170 92 171 93
rect 169 92 170 93
rect 168 92 169 93
rect 167 92 168 93
rect 166 92 167 93
rect 165 92 166 93
rect 164 92 165 93
rect 148 92 149 93
rect 147 92 148 93
rect 146 92 147 93
rect 145 92 146 93
rect 144 92 145 93
rect 143 92 144 93
rect 142 92 143 93
rect 141 92 142 93
rect 140 92 141 93
rect 126 92 127 93
rect 125 92 126 93
rect 124 92 125 93
rect 123 92 124 93
rect 122 92 123 93
rect 121 92 122 93
rect 120 92 121 93
rect 119 92 120 93
rect 118 92 119 93
rect 117 92 118 93
rect 116 92 117 93
rect 115 92 116 93
rect 114 92 115 93
rect 113 92 114 93
rect 112 92 113 93
rect 111 92 112 93
rect 110 92 111 93
rect 109 92 110 93
rect 108 92 109 93
rect 107 92 108 93
rect 106 92 107 93
rect 105 92 106 93
rect 104 92 105 93
rect 103 92 104 93
rect 102 92 103 93
rect 101 92 102 93
rect 100 92 101 93
rect 99 92 100 93
rect 98 92 99 93
rect 97 92 98 93
rect 96 92 97 93
rect 95 92 96 93
rect 94 92 95 93
rect 93 92 94 93
rect 92 92 93 93
rect 91 92 92 93
rect 90 92 91 93
rect 89 92 90 93
rect 88 92 89 93
rect 87 92 88 93
rect 86 92 87 93
rect 85 92 86 93
rect 84 92 85 93
rect 83 92 84 93
rect 82 92 83 93
rect 81 92 82 93
rect 80 92 81 93
rect 64 92 65 93
rect 63 92 64 93
rect 62 92 63 93
rect 61 92 62 93
rect 60 92 61 93
rect 59 92 60 93
rect 58 92 59 93
rect 57 92 58 93
rect 56 92 57 93
rect 55 92 56 93
rect 54 92 55 93
rect 53 92 54 93
rect 52 92 53 93
rect 51 92 52 93
rect 50 92 51 93
rect 49 92 50 93
rect 48 92 49 93
rect 47 92 48 93
rect 46 92 47 93
rect 45 92 46 93
rect 44 92 45 93
rect 32 92 33 93
rect 31 92 32 93
rect 30 92 31 93
rect 29 92 30 93
rect 28 92 29 93
rect 27 92 28 93
rect 26 92 27 93
rect 25 92 26 93
rect 24 92 25 93
rect 23 92 24 93
rect 22 92 23 93
rect 21 92 22 93
rect 20 92 21 93
rect 19 92 20 93
rect 18 92 19 93
rect 17 92 18 93
rect 16 92 17 93
rect 15 92 16 93
rect 14 92 15 93
rect 13 92 14 93
rect 12 92 13 93
rect 11 92 12 93
rect 10 92 11 93
rect 9 92 10 93
rect 8 92 9 93
rect 197 93 198 94
rect 196 93 197 94
rect 195 93 196 94
rect 194 93 195 94
rect 193 93 194 94
rect 192 93 193 94
rect 191 93 192 94
rect 190 93 191 94
rect 189 93 190 94
rect 180 93 181 94
rect 179 93 180 94
rect 178 93 179 94
rect 177 93 178 94
rect 176 93 177 94
rect 175 93 176 94
rect 167 93 168 94
rect 166 93 167 94
rect 165 93 166 94
rect 164 93 165 94
rect 149 93 150 94
rect 148 93 149 94
rect 147 93 148 94
rect 146 93 147 94
rect 145 93 146 94
rect 144 93 145 94
rect 123 93 124 94
rect 122 93 123 94
rect 121 93 122 94
rect 120 93 121 94
rect 119 93 120 94
rect 118 93 119 94
rect 117 93 118 94
rect 116 93 117 94
rect 115 93 116 94
rect 114 93 115 94
rect 113 93 114 94
rect 112 93 113 94
rect 111 93 112 94
rect 110 93 111 94
rect 109 93 110 94
rect 108 93 109 94
rect 107 93 108 94
rect 106 93 107 94
rect 105 93 106 94
rect 104 93 105 94
rect 103 93 104 94
rect 102 93 103 94
rect 101 93 102 94
rect 100 93 101 94
rect 99 93 100 94
rect 98 93 99 94
rect 97 93 98 94
rect 96 93 97 94
rect 95 93 96 94
rect 94 93 95 94
rect 93 93 94 94
rect 92 93 93 94
rect 91 93 92 94
rect 90 93 91 94
rect 89 93 90 94
rect 88 93 89 94
rect 87 93 88 94
rect 86 93 87 94
rect 85 93 86 94
rect 84 93 85 94
rect 83 93 84 94
rect 82 93 83 94
rect 81 93 82 94
rect 80 93 81 94
rect 79 93 80 94
rect 78 93 79 94
rect 77 93 78 94
rect 63 93 64 94
rect 62 93 63 94
rect 61 93 62 94
rect 60 93 61 94
rect 59 93 60 94
rect 58 93 59 94
rect 57 93 58 94
rect 56 93 57 94
rect 55 93 56 94
rect 54 93 55 94
rect 53 93 54 94
rect 52 93 53 94
rect 51 93 52 94
rect 50 93 51 94
rect 49 93 50 94
rect 48 93 49 94
rect 47 93 48 94
rect 46 93 47 94
rect 33 93 34 94
rect 32 93 33 94
rect 31 93 32 94
rect 30 93 31 94
rect 29 93 30 94
rect 28 93 29 94
rect 27 93 28 94
rect 26 93 27 94
rect 25 93 26 94
rect 24 93 25 94
rect 23 93 24 94
rect 22 93 23 94
rect 21 93 22 94
rect 20 93 21 94
rect 19 93 20 94
rect 18 93 19 94
rect 17 93 18 94
rect 16 93 17 94
rect 15 93 16 94
rect 14 93 15 94
rect 13 93 14 94
rect 12 93 13 94
rect 11 93 12 94
rect 10 93 11 94
rect 9 93 10 94
rect 8 93 9 94
rect 197 94 198 95
rect 196 94 197 95
rect 195 94 196 95
rect 194 94 195 95
rect 193 94 194 95
rect 192 94 193 95
rect 191 94 192 95
rect 190 94 191 95
rect 189 94 190 95
rect 180 94 181 95
rect 179 94 180 95
rect 178 94 179 95
rect 177 94 178 95
rect 165 94 166 95
rect 164 94 165 95
rect 163 94 164 95
rect 149 94 150 95
rect 148 94 149 95
rect 147 94 148 95
rect 121 94 122 95
rect 120 94 121 95
rect 119 94 120 95
rect 118 94 119 95
rect 117 94 118 95
rect 116 94 117 95
rect 115 94 116 95
rect 114 94 115 95
rect 113 94 114 95
rect 112 94 113 95
rect 111 94 112 95
rect 110 94 111 95
rect 109 94 110 95
rect 108 94 109 95
rect 107 94 108 95
rect 106 94 107 95
rect 105 94 106 95
rect 104 94 105 95
rect 103 94 104 95
rect 102 94 103 95
rect 101 94 102 95
rect 100 94 101 95
rect 99 94 100 95
rect 98 94 99 95
rect 97 94 98 95
rect 96 94 97 95
rect 95 94 96 95
rect 94 94 95 95
rect 93 94 94 95
rect 92 94 93 95
rect 91 94 92 95
rect 90 94 91 95
rect 89 94 90 95
rect 88 94 89 95
rect 87 94 88 95
rect 86 94 87 95
rect 85 94 86 95
rect 84 94 85 95
rect 83 94 84 95
rect 82 94 83 95
rect 81 94 82 95
rect 80 94 81 95
rect 79 94 80 95
rect 78 94 79 95
rect 77 94 78 95
rect 76 94 77 95
rect 75 94 76 95
rect 63 94 64 95
rect 62 94 63 95
rect 61 94 62 95
rect 60 94 61 95
rect 59 94 60 95
rect 58 94 59 95
rect 57 94 58 95
rect 56 94 57 95
rect 55 94 56 95
rect 54 94 55 95
rect 53 94 54 95
rect 52 94 53 95
rect 51 94 52 95
rect 50 94 51 95
rect 49 94 50 95
rect 48 94 49 95
rect 47 94 48 95
rect 34 94 35 95
rect 33 94 34 95
rect 32 94 33 95
rect 31 94 32 95
rect 30 94 31 95
rect 29 94 30 95
rect 28 94 29 95
rect 27 94 28 95
rect 26 94 27 95
rect 25 94 26 95
rect 24 94 25 95
rect 23 94 24 95
rect 22 94 23 95
rect 21 94 22 95
rect 20 94 21 95
rect 19 94 20 95
rect 18 94 19 95
rect 17 94 18 95
rect 16 94 17 95
rect 15 94 16 95
rect 14 94 15 95
rect 13 94 14 95
rect 12 94 13 95
rect 11 94 12 95
rect 10 94 11 95
rect 9 94 10 95
rect 8 94 9 95
rect 197 95 198 96
rect 193 95 194 96
rect 189 95 190 96
rect 180 95 181 96
rect 179 95 180 96
rect 164 95 165 96
rect 163 95 164 96
rect 149 95 150 96
rect 119 95 120 96
rect 118 95 119 96
rect 117 95 118 96
rect 116 95 117 96
rect 115 95 116 96
rect 114 95 115 96
rect 113 95 114 96
rect 112 95 113 96
rect 111 95 112 96
rect 110 95 111 96
rect 109 95 110 96
rect 108 95 109 96
rect 107 95 108 96
rect 106 95 107 96
rect 105 95 106 96
rect 104 95 105 96
rect 103 95 104 96
rect 102 95 103 96
rect 101 95 102 96
rect 100 95 101 96
rect 99 95 100 96
rect 98 95 99 96
rect 97 95 98 96
rect 96 95 97 96
rect 95 95 96 96
rect 94 95 95 96
rect 93 95 94 96
rect 92 95 93 96
rect 91 95 92 96
rect 90 95 91 96
rect 89 95 90 96
rect 88 95 89 96
rect 87 95 88 96
rect 86 95 87 96
rect 85 95 86 96
rect 84 95 85 96
rect 83 95 84 96
rect 82 95 83 96
rect 81 95 82 96
rect 80 95 81 96
rect 79 95 80 96
rect 78 95 79 96
rect 77 95 78 96
rect 76 95 77 96
rect 75 95 76 96
rect 74 95 75 96
rect 73 95 74 96
rect 63 95 64 96
rect 62 95 63 96
rect 61 95 62 96
rect 60 95 61 96
rect 59 95 60 96
rect 58 95 59 96
rect 57 95 58 96
rect 56 95 57 96
rect 55 95 56 96
rect 54 95 55 96
rect 53 95 54 96
rect 52 95 53 96
rect 51 95 52 96
rect 50 95 51 96
rect 49 95 50 96
rect 36 95 37 96
rect 35 95 36 96
rect 34 95 35 96
rect 33 95 34 96
rect 32 95 33 96
rect 31 95 32 96
rect 30 95 31 96
rect 29 95 30 96
rect 28 95 29 96
rect 27 95 28 96
rect 26 95 27 96
rect 25 95 26 96
rect 24 95 25 96
rect 23 95 24 96
rect 22 95 23 96
rect 21 95 22 96
rect 20 95 21 96
rect 19 95 20 96
rect 18 95 19 96
rect 17 95 18 96
rect 16 95 17 96
rect 15 95 16 96
rect 14 95 15 96
rect 13 95 14 96
rect 12 95 13 96
rect 11 95 12 96
rect 10 95 11 96
rect 9 95 10 96
rect 8 95 9 96
rect 195 96 196 97
rect 194 96 195 97
rect 193 96 194 97
rect 192 96 193 97
rect 189 96 190 97
rect 181 96 182 97
rect 180 96 181 97
rect 179 96 180 97
rect 164 96 165 97
rect 163 96 164 97
rect 117 96 118 97
rect 116 96 117 97
rect 115 96 116 97
rect 114 96 115 97
rect 113 96 114 97
rect 112 96 113 97
rect 111 96 112 97
rect 110 96 111 97
rect 109 96 110 97
rect 108 96 109 97
rect 107 96 108 97
rect 106 96 107 97
rect 105 96 106 97
rect 104 96 105 97
rect 103 96 104 97
rect 102 96 103 97
rect 101 96 102 97
rect 100 96 101 97
rect 99 96 100 97
rect 98 96 99 97
rect 97 96 98 97
rect 96 96 97 97
rect 95 96 96 97
rect 94 96 95 97
rect 93 96 94 97
rect 92 96 93 97
rect 91 96 92 97
rect 90 96 91 97
rect 89 96 90 97
rect 88 96 89 97
rect 87 96 88 97
rect 86 96 87 97
rect 85 96 86 97
rect 84 96 85 97
rect 83 96 84 97
rect 82 96 83 97
rect 81 96 82 97
rect 80 96 81 97
rect 79 96 80 97
rect 78 96 79 97
rect 77 96 78 97
rect 76 96 77 97
rect 75 96 76 97
rect 74 96 75 97
rect 73 96 74 97
rect 72 96 73 97
rect 71 96 72 97
rect 63 96 64 97
rect 62 96 63 97
rect 61 96 62 97
rect 60 96 61 97
rect 59 96 60 97
rect 58 96 59 97
rect 57 96 58 97
rect 56 96 57 97
rect 55 96 56 97
rect 54 96 55 97
rect 53 96 54 97
rect 52 96 53 97
rect 51 96 52 97
rect 50 96 51 97
rect 37 96 38 97
rect 36 96 37 97
rect 35 96 36 97
rect 34 96 35 97
rect 33 96 34 97
rect 32 96 33 97
rect 31 96 32 97
rect 30 96 31 97
rect 29 96 30 97
rect 28 96 29 97
rect 27 96 28 97
rect 26 96 27 97
rect 25 96 26 97
rect 24 96 25 97
rect 23 96 24 97
rect 22 96 23 97
rect 21 96 22 97
rect 20 96 21 97
rect 19 96 20 97
rect 18 96 19 97
rect 17 96 18 97
rect 16 96 17 97
rect 15 96 16 97
rect 14 96 15 97
rect 13 96 14 97
rect 12 96 13 97
rect 11 96 12 97
rect 10 96 11 97
rect 9 96 10 97
rect 8 96 9 97
rect 7 96 8 97
rect 196 97 197 98
rect 195 97 196 98
rect 194 97 195 98
rect 193 97 194 98
rect 192 97 193 98
rect 191 97 192 98
rect 190 97 191 98
rect 189 97 190 98
rect 181 97 182 98
rect 180 97 181 98
rect 163 97 164 98
rect 162 97 163 98
rect 116 97 117 98
rect 115 97 116 98
rect 114 97 115 98
rect 113 97 114 98
rect 112 97 113 98
rect 111 97 112 98
rect 110 97 111 98
rect 109 97 110 98
rect 108 97 109 98
rect 107 97 108 98
rect 106 97 107 98
rect 105 97 106 98
rect 104 97 105 98
rect 103 97 104 98
rect 102 97 103 98
rect 101 97 102 98
rect 100 97 101 98
rect 99 97 100 98
rect 98 97 99 98
rect 97 97 98 98
rect 96 97 97 98
rect 95 97 96 98
rect 94 97 95 98
rect 93 97 94 98
rect 92 97 93 98
rect 91 97 92 98
rect 90 97 91 98
rect 89 97 90 98
rect 88 97 89 98
rect 87 97 88 98
rect 86 97 87 98
rect 85 97 86 98
rect 84 97 85 98
rect 83 97 84 98
rect 82 97 83 98
rect 81 97 82 98
rect 80 97 81 98
rect 79 97 80 98
rect 78 97 79 98
rect 77 97 78 98
rect 76 97 77 98
rect 75 97 76 98
rect 74 97 75 98
rect 73 97 74 98
rect 72 97 73 98
rect 71 97 72 98
rect 70 97 71 98
rect 63 97 64 98
rect 62 97 63 98
rect 61 97 62 98
rect 60 97 61 98
rect 59 97 60 98
rect 58 97 59 98
rect 57 97 58 98
rect 56 97 57 98
rect 55 97 56 98
rect 54 97 55 98
rect 53 97 54 98
rect 52 97 53 98
rect 51 97 52 98
rect 50 97 51 98
rect 39 97 40 98
rect 38 97 39 98
rect 37 97 38 98
rect 36 97 37 98
rect 35 97 36 98
rect 34 97 35 98
rect 33 97 34 98
rect 32 97 33 98
rect 31 97 32 98
rect 30 97 31 98
rect 29 97 30 98
rect 28 97 29 98
rect 27 97 28 98
rect 26 97 27 98
rect 25 97 26 98
rect 24 97 25 98
rect 23 97 24 98
rect 22 97 23 98
rect 21 97 22 98
rect 20 97 21 98
rect 19 97 20 98
rect 18 97 19 98
rect 17 97 18 98
rect 16 97 17 98
rect 15 97 16 98
rect 14 97 15 98
rect 13 97 14 98
rect 12 97 13 98
rect 11 97 12 98
rect 10 97 11 98
rect 9 97 10 98
rect 8 97 9 98
rect 7 97 8 98
rect 197 98 198 99
rect 196 98 197 99
rect 195 98 196 99
rect 192 98 193 99
rect 191 98 192 99
rect 190 98 191 99
rect 189 98 190 99
rect 181 98 182 99
rect 180 98 181 99
rect 172 98 173 99
rect 163 98 164 99
rect 162 98 163 99
rect 115 98 116 99
rect 114 98 115 99
rect 113 98 114 99
rect 112 98 113 99
rect 111 98 112 99
rect 110 98 111 99
rect 109 98 110 99
rect 108 98 109 99
rect 107 98 108 99
rect 106 98 107 99
rect 105 98 106 99
rect 104 98 105 99
rect 103 98 104 99
rect 102 98 103 99
rect 101 98 102 99
rect 100 98 101 99
rect 99 98 100 99
rect 98 98 99 99
rect 97 98 98 99
rect 96 98 97 99
rect 95 98 96 99
rect 94 98 95 99
rect 93 98 94 99
rect 92 98 93 99
rect 91 98 92 99
rect 90 98 91 99
rect 89 98 90 99
rect 88 98 89 99
rect 87 98 88 99
rect 86 98 87 99
rect 85 98 86 99
rect 84 98 85 99
rect 83 98 84 99
rect 82 98 83 99
rect 81 98 82 99
rect 80 98 81 99
rect 79 98 80 99
rect 78 98 79 99
rect 77 98 78 99
rect 76 98 77 99
rect 75 98 76 99
rect 74 98 75 99
rect 73 98 74 99
rect 72 98 73 99
rect 71 98 72 99
rect 63 98 64 99
rect 62 98 63 99
rect 61 98 62 99
rect 60 98 61 99
rect 59 98 60 99
rect 58 98 59 99
rect 57 98 58 99
rect 56 98 57 99
rect 55 98 56 99
rect 54 98 55 99
rect 53 98 54 99
rect 52 98 53 99
rect 51 98 52 99
rect 41 98 42 99
rect 40 98 41 99
rect 39 98 40 99
rect 38 98 39 99
rect 37 98 38 99
rect 36 98 37 99
rect 35 98 36 99
rect 34 98 35 99
rect 33 98 34 99
rect 32 98 33 99
rect 31 98 32 99
rect 30 98 31 99
rect 29 98 30 99
rect 28 98 29 99
rect 27 98 28 99
rect 26 98 27 99
rect 25 98 26 99
rect 24 98 25 99
rect 23 98 24 99
rect 22 98 23 99
rect 21 98 22 99
rect 20 98 21 99
rect 19 98 20 99
rect 18 98 19 99
rect 17 98 18 99
rect 16 98 17 99
rect 15 98 16 99
rect 14 98 15 99
rect 13 98 14 99
rect 12 98 13 99
rect 11 98 12 99
rect 10 98 11 99
rect 9 98 10 99
rect 8 98 9 99
rect 7 98 8 99
rect 197 99 198 100
rect 196 99 197 100
rect 181 99 182 100
rect 180 99 181 100
rect 173 99 174 100
rect 172 99 173 100
rect 163 99 164 100
rect 162 99 163 100
rect 114 99 115 100
rect 113 99 114 100
rect 112 99 113 100
rect 111 99 112 100
rect 110 99 111 100
rect 109 99 110 100
rect 108 99 109 100
rect 107 99 108 100
rect 106 99 107 100
rect 105 99 106 100
rect 104 99 105 100
rect 103 99 104 100
rect 102 99 103 100
rect 101 99 102 100
rect 100 99 101 100
rect 99 99 100 100
rect 98 99 99 100
rect 97 99 98 100
rect 96 99 97 100
rect 95 99 96 100
rect 94 99 95 100
rect 93 99 94 100
rect 92 99 93 100
rect 91 99 92 100
rect 90 99 91 100
rect 89 99 90 100
rect 88 99 89 100
rect 87 99 88 100
rect 86 99 87 100
rect 85 99 86 100
rect 84 99 85 100
rect 83 99 84 100
rect 82 99 83 100
rect 81 99 82 100
rect 80 99 81 100
rect 79 99 80 100
rect 78 99 79 100
rect 77 99 78 100
rect 76 99 77 100
rect 75 99 76 100
rect 74 99 75 100
rect 73 99 74 100
rect 72 99 73 100
rect 63 99 64 100
rect 62 99 63 100
rect 61 99 62 100
rect 60 99 61 100
rect 59 99 60 100
rect 58 99 59 100
rect 57 99 58 100
rect 56 99 57 100
rect 55 99 56 100
rect 54 99 55 100
rect 53 99 54 100
rect 52 99 53 100
rect 43 99 44 100
rect 42 99 43 100
rect 41 99 42 100
rect 40 99 41 100
rect 39 99 40 100
rect 38 99 39 100
rect 37 99 38 100
rect 36 99 37 100
rect 35 99 36 100
rect 34 99 35 100
rect 33 99 34 100
rect 32 99 33 100
rect 31 99 32 100
rect 30 99 31 100
rect 29 99 30 100
rect 28 99 29 100
rect 27 99 28 100
rect 26 99 27 100
rect 25 99 26 100
rect 24 99 25 100
rect 23 99 24 100
rect 22 99 23 100
rect 21 99 22 100
rect 20 99 21 100
rect 19 99 20 100
rect 18 99 19 100
rect 17 99 18 100
rect 16 99 17 100
rect 14 99 15 100
rect 13 99 14 100
rect 12 99 13 100
rect 11 99 12 100
rect 10 99 11 100
rect 9 99 10 100
rect 8 99 9 100
rect 7 99 8 100
rect 181 100 182 101
rect 180 100 181 101
rect 173 100 174 101
rect 172 100 173 101
rect 163 100 164 101
rect 162 100 163 101
rect 113 100 114 101
rect 112 100 113 101
rect 111 100 112 101
rect 110 100 111 101
rect 109 100 110 101
rect 108 100 109 101
rect 107 100 108 101
rect 106 100 107 101
rect 105 100 106 101
rect 104 100 105 101
rect 103 100 104 101
rect 102 100 103 101
rect 101 100 102 101
rect 100 100 101 101
rect 99 100 100 101
rect 98 100 99 101
rect 97 100 98 101
rect 96 100 97 101
rect 95 100 96 101
rect 94 100 95 101
rect 93 100 94 101
rect 92 100 93 101
rect 91 100 92 101
rect 90 100 91 101
rect 89 100 90 101
rect 88 100 89 101
rect 87 100 88 101
rect 86 100 87 101
rect 85 100 86 101
rect 84 100 85 101
rect 83 100 84 101
rect 82 100 83 101
rect 81 100 82 101
rect 80 100 81 101
rect 79 100 80 101
rect 78 100 79 101
rect 77 100 78 101
rect 76 100 77 101
rect 75 100 76 101
rect 74 100 75 101
rect 64 100 65 101
rect 63 100 64 101
rect 62 100 63 101
rect 61 100 62 101
rect 60 100 61 101
rect 59 100 60 101
rect 58 100 59 101
rect 57 100 58 101
rect 56 100 57 101
rect 55 100 56 101
rect 54 100 55 101
rect 53 100 54 101
rect 52 100 53 101
rect 44 100 45 101
rect 43 100 44 101
rect 42 100 43 101
rect 41 100 42 101
rect 40 100 41 101
rect 39 100 40 101
rect 38 100 39 101
rect 37 100 38 101
rect 36 100 37 101
rect 35 100 36 101
rect 34 100 35 101
rect 33 100 34 101
rect 32 100 33 101
rect 31 100 32 101
rect 30 100 31 101
rect 29 100 30 101
rect 28 100 29 101
rect 27 100 28 101
rect 26 100 27 101
rect 25 100 26 101
rect 24 100 25 101
rect 23 100 24 101
rect 22 100 23 101
rect 21 100 22 101
rect 20 100 21 101
rect 19 100 20 101
rect 18 100 19 101
rect 17 100 18 101
rect 16 100 17 101
rect 13 100 14 101
rect 12 100 13 101
rect 11 100 12 101
rect 10 100 11 101
rect 9 100 10 101
rect 8 100 9 101
rect 7 100 8 101
rect 181 101 182 102
rect 180 101 181 102
rect 179 101 180 102
rect 178 101 179 102
rect 177 101 178 102
rect 176 101 177 102
rect 175 101 176 102
rect 174 101 175 102
rect 173 101 174 102
rect 172 101 173 102
rect 164 101 165 102
rect 163 101 164 102
rect 162 101 163 102
rect 131 101 132 102
rect 130 101 131 102
rect 129 101 130 102
rect 128 101 129 102
rect 127 101 128 102
rect 126 101 127 102
rect 125 101 126 102
rect 124 101 125 102
rect 123 101 124 102
rect 122 101 123 102
rect 121 101 122 102
rect 120 101 121 102
rect 119 101 120 102
rect 112 101 113 102
rect 111 101 112 102
rect 110 101 111 102
rect 109 101 110 102
rect 108 101 109 102
rect 107 101 108 102
rect 106 101 107 102
rect 105 101 106 102
rect 104 101 105 102
rect 103 101 104 102
rect 102 101 103 102
rect 101 101 102 102
rect 100 101 101 102
rect 99 101 100 102
rect 98 101 99 102
rect 97 101 98 102
rect 96 101 97 102
rect 95 101 96 102
rect 94 101 95 102
rect 93 101 94 102
rect 92 101 93 102
rect 91 101 92 102
rect 90 101 91 102
rect 89 101 90 102
rect 88 101 89 102
rect 87 101 88 102
rect 86 101 87 102
rect 85 101 86 102
rect 84 101 85 102
rect 83 101 84 102
rect 82 101 83 102
rect 81 101 82 102
rect 80 101 81 102
rect 79 101 80 102
rect 78 101 79 102
rect 77 101 78 102
rect 76 101 77 102
rect 64 101 65 102
rect 63 101 64 102
rect 62 101 63 102
rect 61 101 62 102
rect 60 101 61 102
rect 59 101 60 102
rect 58 101 59 102
rect 57 101 58 102
rect 56 101 57 102
rect 55 101 56 102
rect 54 101 55 102
rect 53 101 54 102
rect 52 101 53 102
rect 45 101 46 102
rect 44 101 45 102
rect 43 101 44 102
rect 42 101 43 102
rect 41 101 42 102
rect 40 101 41 102
rect 39 101 40 102
rect 38 101 39 102
rect 37 101 38 102
rect 36 101 37 102
rect 35 101 36 102
rect 34 101 35 102
rect 33 101 34 102
rect 32 101 33 102
rect 31 101 32 102
rect 30 101 31 102
rect 29 101 30 102
rect 28 101 29 102
rect 27 101 28 102
rect 26 101 27 102
rect 25 101 26 102
rect 24 101 25 102
rect 23 101 24 102
rect 22 101 23 102
rect 21 101 22 102
rect 20 101 21 102
rect 19 101 20 102
rect 18 101 19 102
rect 17 101 18 102
rect 16 101 17 102
rect 13 101 14 102
rect 12 101 13 102
rect 11 101 12 102
rect 10 101 11 102
rect 9 101 10 102
rect 8 101 9 102
rect 7 101 8 102
rect 180 102 181 103
rect 179 102 180 103
rect 178 102 179 103
rect 177 102 178 103
rect 176 102 177 103
rect 175 102 176 103
rect 174 102 175 103
rect 173 102 174 103
rect 172 102 173 103
rect 165 102 166 103
rect 164 102 165 103
rect 163 102 164 103
rect 135 102 136 103
rect 134 102 135 103
rect 133 102 134 103
rect 132 102 133 103
rect 131 102 132 103
rect 130 102 131 103
rect 129 102 130 103
rect 128 102 129 103
rect 127 102 128 103
rect 126 102 127 103
rect 125 102 126 103
rect 124 102 125 103
rect 123 102 124 103
rect 122 102 123 103
rect 121 102 122 103
rect 120 102 121 103
rect 119 102 120 103
rect 118 102 119 103
rect 117 102 118 103
rect 116 102 117 103
rect 115 102 116 103
rect 112 102 113 103
rect 111 102 112 103
rect 110 102 111 103
rect 109 102 110 103
rect 108 102 109 103
rect 107 102 108 103
rect 106 102 107 103
rect 105 102 106 103
rect 104 102 105 103
rect 103 102 104 103
rect 102 102 103 103
rect 101 102 102 103
rect 100 102 101 103
rect 99 102 100 103
rect 98 102 99 103
rect 97 102 98 103
rect 96 102 97 103
rect 95 102 96 103
rect 94 102 95 103
rect 93 102 94 103
rect 92 102 93 103
rect 91 102 92 103
rect 90 102 91 103
rect 89 102 90 103
rect 88 102 89 103
rect 87 102 88 103
rect 86 102 87 103
rect 85 102 86 103
rect 84 102 85 103
rect 83 102 84 103
rect 82 102 83 103
rect 81 102 82 103
rect 80 102 81 103
rect 79 102 80 103
rect 78 102 79 103
rect 65 102 66 103
rect 64 102 65 103
rect 63 102 64 103
rect 62 102 63 103
rect 61 102 62 103
rect 60 102 61 103
rect 59 102 60 103
rect 58 102 59 103
rect 57 102 58 103
rect 56 102 57 103
rect 55 102 56 103
rect 54 102 55 103
rect 53 102 54 103
rect 46 102 47 103
rect 45 102 46 103
rect 44 102 45 103
rect 43 102 44 103
rect 42 102 43 103
rect 41 102 42 103
rect 40 102 41 103
rect 39 102 40 103
rect 38 102 39 103
rect 37 102 38 103
rect 36 102 37 103
rect 35 102 36 103
rect 34 102 35 103
rect 33 102 34 103
rect 32 102 33 103
rect 31 102 32 103
rect 30 102 31 103
rect 29 102 30 103
rect 28 102 29 103
rect 27 102 28 103
rect 26 102 27 103
rect 25 102 26 103
rect 24 102 25 103
rect 23 102 24 103
rect 22 102 23 103
rect 21 102 22 103
rect 20 102 21 103
rect 19 102 20 103
rect 18 102 19 103
rect 17 102 18 103
rect 13 102 14 103
rect 12 102 13 103
rect 11 102 12 103
rect 10 102 11 103
rect 9 102 10 103
rect 8 102 9 103
rect 7 102 8 103
rect 6 102 7 103
rect 196 103 197 104
rect 195 103 196 104
rect 191 103 192 104
rect 190 103 191 104
rect 180 103 181 104
rect 179 103 180 104
rect 178 103 179 104
rect 177 103 178 104
rect 176 103 177 104
rect 175 103 176 104
rect 174 103 175 104
rect 173 103 174 104
rect 172 103 173 104
rect 166 103 167 104
rect 165 103 166 104
rect 164 103 165 104
rect 163 103 164 104
rect 135 103 136 104
rect 134 103 135 104
rect 133 103 134 104
rect 132 103 133 104
rect 131 103 132 104
rect 130 103 131 104
rect 129 103 130 104
rect 128 103 129 104
rect 127 103 128 104
rect 126 103 127 104
rect 125 103 126 104
rect 124 103 125 104
rect 123 103 124 104
rect 122 103 123 104
rect 121 103 122 104
rect 120 103 121 104
rect 119 103 120 104
rect 118 103 119 104
rect 117 103 118 104
rect 116 103 117 104
rect 115 103 116 104
rect 114 103 115 104
rect 113 103 114 104
rect 111 103 112 104
rect 110 103 111 104
rect 109 103 110 104
rect 108 103 109 104
rect 107 103 108 104
rect 106 103 107 104
rect 105 103 106 104
rect 104 103 105 104
rect 103 103 104 104
rect 102 103 103 104
rect 101 103 102 104
rect 100 103 101 104
rect 99 103 100 104
rect 98 103 99 104
rect 93 103 94 104
rect 92 103 93 104
rect 91 103 92 104
rect 90 103 91 104
rect 89 103 90 104
rect 88 103 89 104
rect 87 103 88 104
rect 86 103 87 104
rect 85 103 86 104
rect 84 103 85 104
rect 83 103 84 104
rect 82 103 83 104
rect 81 103 82 104
rect 66 103 67 104
rect 65 103 66 104
rect 64 103 65 104
rect 63 103 64 104
rect 62 103 63 104
rect 61 103 62 104
rect 60 103 61 104
rect 59 103 60 104
rect 58 103 59 104
rect 57 103 58 104
rect 56 103 57 104
rect 55 103 56 104
rect 54 103 55 104
rect 53 103 54 104
rect 47 103 48 104
rect 46 103 47 104
rect 45 103 46 104
rect 44 103 45 104
rect 43 103 44 104
rect 42 103 43 104
rect 41 103 42 104
rect 40 103 41 104
rect 39 103 40 104
rect 38 103 39 104
rect 37 103 38 104
rect 36 103 37 104
rect 35 103 36 104
rect 34 103 35 104
rect 33 103 34 104
rect 32 103 33 104
rect 31 103 32 104
rect 30 103 31 104
rect 29 103 30 104
rect 28 103 29 104
rect 27 103 28 104
rect 26 103 27 104
rect 25 103 26 104
rect 24 103 25 104
rect 23 103 24 104
rect 22 103 23 104
rect 21 103 22 104
rect 20 103 21 104
rect 19 103 20 104
rect 18 103 19 104
rect 17 103 18 104
rect 13 103 14 104
rect 12 103 13 104
rect 11 103 12 104
rect 10 103 11 104
rect 9 103 10 104
rect 8 103 9 104
rect 7 103 8 104
rect 197 104 198 105
rect 196 104 197 105
rect 192 104 193 105
rect 191 104 192 105
rect 190 104 191 105
rect 189 104 190 105
rect 180 104 181 105
rect 179 104 180 105
rect 178 104 179 105
rect 177 104 178 105
rect 176 104 177 105
rect 175 104 176 105
rect 174 104 175 105
rect 173 104 174 105
rect 172 104 173 105
rect 167 104 168 105
rect 166 104 167 105
rect 165 104 166 105
rect 164 104 165 105
rect 163 104 164 105
rect 133 104 134 105
rect 132 104 133 105
rect 131 104 132 105
rect 130 104 131 105
rect 129 104 130 105
rect 128 104 129 105
rect 127 104 128 105
rect 126 104 127 105
rect 125 104 126 105
rect 124 104 125 105
rect 123 104 124 105
rect 122 104 123 105
rect 121 104 122 105
rect 120 104 121 105
rect 119 104 120 105
rect 118 104 119 105
rect 117 104 118 105
rect 116 104 117 105
rect 115 104 116 105
rect 114 104 115 105
rect 113 104 114 105
rect 112 104 113 105
rect 111 104 112 105
rect 110 104 111 105
rect 109 104 110 105
rect 108 104 109 105
rect 107 104 108 105
rect 106 104 107 105
rect 105 104 106 105
rect 104 104 105 105
rect 103 104 104 105
rect 102 104 103 105
rect 101 104 102 105
rect 100 104 101 105
rect 99 104 100 105
rect 98 104 99 105
rect 67 104 68 105
rect 66 104 67 105
rect 65 104 66 105
rect 64 104 65 105
rect 63 104 64 105
rect 62 104 63 105
rect 61 104 62 105
rect 60 104 61 105
rect 59 104 60 105
rect 58 104 59 105
rect 57 104 58 105
rect 56 104 57 105
rect 55 104 56 105
rect 54 104 55 105
rect 53 104 54 105
rect 47 104 48 105
rect 46 104 47 105
rect 45 104 46 105
rect 44 104 45 105
rect 43 104 44 105
rect 42 104 43 105
rect 41 104 42 105
rect 40 104 41 105
rect 39 104 40 105
rect 38 104 39 105
rect 37 104 38 105
rect 36 104 37 105
rect 35 104 36 105
rect 34 104 35 105
rect 33 104 34 105
rect 32 104 33 105
rect 31 104 32 105
rect 30 104 31 105
rect 29 104 30 105
rect 28 104 29 105
rect 27 104 28 105
rect 26 104 27 105
rect 25 104 26 105
rect 24 104 25 105
rect 23 104 24 105
rect 22 104 23 105
rect 21 104 22 105
rect 20 104 21 105
rect 19 104 20 105
rect 18 104 19 105
rect 17 104 18 105
rect 13 104 14 105
rect 12 104 13 105
rect 11 104 12 105
rect 10 104 11 105
rect 9 104 10 105
rect 8 104 9 105
rect 7 104 8 105
rect 6 104 7 105
rect 197 105 198 106
rect 193 105 194 106
rect 192 105 193 106
rect 191 105 192 106
rect 189 105 190 106
rect 188 105 189 106
rect 173 105 174 106
rect 172 105 173 106
rect 132 105 133 106
rect 131 105 132 106
rect 130 105 131 106
rect 129 105 130 106
rect 128 105 129 106
rect 127 105 128 106
rect 126 105 127 106
rect 125 105 126 106
rect 124 105 125 106
rect 123 105 124 106
rect 122 105 123 106
rect 121 105 122 106
rect 120 105 121 106
rect 119 105 120 106
rect 118 105 119 106
rect 117 105 118 106
rect 116 105 117 106
rect 115 105 116 106
rect 114 105 115 106
rect 113 105 114 106
rect 112 105 113 106
rect 111 105 112 106
rect 110 105 111 106
rect 109 105 110 106
rect 108 105 109 106
rect 107 105 108 106
rect 106 105 107 106
rect 105 105 106 106
rect 104 105 105 106
rect 103 105 104 106
rect 102 105 103 106
rect 101 105 102 106
rect 100 105 101 106
rect 99 105 100 106
rect 98 105 99 106
rect 97 105 98 106
rect 68 105 69 106
rect 67 105 68 106
rect 66 105 67 106
rect 65 105 66 106
rect 64 105 65 106
rect 63 105 64 106
rect 62 105 63 106
rect 61 105 62 106
rect 60 105 61 106
rect 59 105 60 106
rect 58 105 59 106
rect 57 105 58 106
rect 56 105 57 106
rect 55 105 56 106
rect 54 105 55 106
rect 53 105 54 106
rect 48 105 49 106
rect 47 105 48 106
rect 46 105 47 106
rect 45 105 46 106
rect 44 105 45 106
rect 43 105 44 106
rect 42 105 43 106
rect 41 105 42 106
rect 40 105 41 106
rect 39 105 40 106
rect 38 105 39 106
rect 37 105 38 106
rect 36 105 37 106
rect 35 105 36 106
rect 34 105 35 106
rect 33 105 34 106
rect 32 105 33 106
rect 31 105 32 106
rect 30 105 31 106
rect 29 105 30 106
rect 28 105 29 106
rect 27 105 28 106
rect 26 105 27 106
rect 25 105 26 106
rect 24 105 25 106
rect 23 105 24 106
rect 22 105 23 106
rect 21 105 22 106
rect 20 105 21 106
rect 19 105 20 106
rect 18 105 19 106
rect 13 105 14 106
rect 12 105 13 106
rect 11 105 12 106
rect 10 105 11 106
rect 9 105 10 106
rect 8 105 9 106
rect 7 105 8 106
rect 6 105 7 106
rect 197 106 198 107
rect 194 106 195 107
rect 193 106 194 107
rect 192 106 193 107
rect 189 106 190 107
rect 188 106 189 107
rect 173 106 174 107
rect 172 106 173 107
rect 130 106 131 107
rect 129 106 130 107
rect 128 106 129 107
rect 127 106 128 107
rect 126 106 127 107
rect 125 106 126 107
rect 124 106 125 107
rect 123 106 124 107
rect 122 106 123 107
rect 121 106 122 107
rect 120 106 121 107
rect 119 106 120 107
rect 118 106 119 107
rect 117 106 118 107
rect 116 106 117 107
rect 115 106 116 107
rect 114 106 115 107
rect 113 106 114 107
rect 112 106 113 107
rect 111 106 112 107
rect 110 106 111 107
rect 109 106 110 107
rect 108 106 109 107
rect 107 106 108 107
rect 106 106 107 107
rect 105 106 106 107
rect 104 106 105 107
rect 103 106 104 107
rect 102 106 103 107
rect 101 106 102 107
rect 100 106 101 107
rect 99 106 100 107
rect 98 106 99 107
rect 97 106 98 107
rect 69 106 70 107
rect 68 106 69 107
rect 67 106 68 107
rect 66 106 67 107
rect 65 106 66 107
rect 64 106 65 107
rect 63 106 64 107
rect 62 106 63 107
rect 61 106 62 107
rect 60 106 61 107
rect 59 106 60 107
rect 58 106 59 107
rect 57 106 58 107
rect 56 106 57 107
rect 55 106 56 107
rect 54 106 55 107
rect 48 106 49 107
rect 47 106 48 107
rect 46 106 47 107
rect 45 106 46 107
rect 44 106 45 107
rect 43 106 44 107
rect 42 106 43 107
rect 41 106 42 107
rect 40 106 41 107
rect 39 106 40 107
rect 38 106 39 107
rect 37 106 38 107
rect 36 106 37 107
rect 35 106 36 107
rect 34 106 35 107
rect 33 106 34 107
rect 32 106 33 107
rect 31 106 32 107
rect 30 106 31 107
rect 29 106 30 107
rect 28 106 29 107
rect 27 106 28 107
rect 26 106 27 107
rect 25 106 26 107
rect 24 106 25 107
rect 23 106 24 107
rect 22 106 23 107
rect 21 106 22 107
rect 20 106 21 107
rect 19 106 20 107
rect 18 106 19 107
rect 13 106 14 107
rect 12 106 13 107
rect 11 106 12 107
rect 10 106 11 107
rect 9 106 10 107
rect 8 106 9 107
rect 7 106 8 107
rect 6 106 7 107
rect 196 107 197 108
rect 195 107 196 108
rect 194 107 195 108
rect 193 107 194 108
rect 192 107 193 108
rect 189 107 190 108
rect 188 107 189 108
rect 129 107 130 108
rect 128 107 129 108
rect 127 107 128 108
rect 126 107 127 108
rect 125 107 126 108
rect 124 107 125 108
rect 123 107 124 108
rect 122 107 123 108
rect 121 107 122 108
rect 120 107 121 108
rect 119 107 120 108
rect 118 107 119 108
rect 117 107 118 108
rect 116 107 117 108
rect 115 107 116 108
rect 114 107 115 108
rect 113 107 114 108
rect 112 107 113 108
rect 111 107 112 108
rect 110 107 111 108
rect 109 107 110 108
rect 108 107 109 108
rect 107 107 108 108
rect 106 107 107 108
rect 105 107 106 108
rect 104 107 105 108
rect 103 107 104 108
rect 102 107 103 108
rect 101 107 102 108
rect 100 107 101 108
rect 99 107 100 108
rect 98 107 99 108
rect 97 107 98 108
rect 71 107 72 108
rect 70 107 71 108
rect 69 107 70 108
rect 68 107 69 108
rect 67 107 68 108
rect 66 107 67 108
rect 65 107 66 108
rect 64 107 65 108
rect 63 107 64 108
rect 62 107 63 108
rect 61 107 62 108
rect 60 107 61 108
rect 59 107 60 108
rect 58 107 59 108
rect 57 107 58 108
rect 56 107 57 108
rect 55 107 56 108
rect 54 107 55 108
rect 48 107 49 108
rect 47 107 48 108
rect 46 107 47 108
rect 45 107 46 108
rect 44 107 45 108
rect 43 107 44 108
rect 42 107 43 108
rect 41 107 42 108
rect 40 107 41 108
rect 39 107 40 108
rect 38 107 39 108
rect 37 107 38 108
rect 36 107 37 108
rect 35 107 36 108
rect 34 107 35 108
rect 33 107 34 108
rect 32 107 33 108
rect 31 107 32 108
rect 30 107 31 108
rect 29 107 30 108
rect 27 107 28 108
rect 26 107 27 108
rect 25 107 26 108
rect 24 107 25 108
rect 23 107 24 108
rect 22 107 23 108
rect 21 107 22 108
rect 20 107 21 108
rect 19 107 20 108
rect 18 107 19 108
rect 14 107 15 108
rect 13 107 14 108
rect 12 107 13 108
rect 11 107 12 108
rect 10 107 11 108
rect 9 107 10 108
rect 8 107 9 108
rect 7 107 8 108
rect 6 107 7 108
rect 195 108 196 109
rect 194 108 195 109
rect 193 108 194 109
rect 190 108 191 109
rect 189 108 190 109
rect 128 108 129 109
rect 127 108 128 109
rect 126 108 127 109
rect 125 108 126 109
rect 124 108 125 109
rect 123 108 124 109
rect 122 108 123 109
rect 121 108 122 109
rect 120 108 121 109
rect 119 108 120 109
rect 118 108 119 109
rect 117 108 118 109
rect 116 108 117 109
rect 115 108 116 109
rect 114 108 115 109
rect 113 108 114 109
rect 112 108 113 109
rect 111 108 112 109
rect 110 108 111 109
rect 109 108 110 109
rect 108 108 109 109
rect 107 108 108 109
rect 106 108 107 109
rect 105 108 106 109
rect 104 108 105 109
rect 103 108 104 109
rect 102 108 103 109
rect 101 108 102 109
rect 100 108 101 109
rect 99 108 100 109
rect 98 108 99 109
rect 97 108 98 109
rect 73 108 74 109
rect 72 108 73 109
rect 71 108 72 109
rect 70 108 71 109
rect 69 108 70 109
rect 68 108 69 109
rect 67 108 68 109
rect 66 108 67 109
rect 65 108 66 109
rect 64 108 65 109
rect 63 108 64 109
rect 62 108 63 109
rect 61 108 62 109
rect 60 108 61 109
rect 59 108 60 109
rect 58 108 59 109
rect 57 108 58 109
rect 56 108 57 109
rect 55 108 56 109
rect 54 108 55 109
rect 49 108 50 109
rect 48 108 49 109
rect 47 108 48 109
rect 46 108 47 109
rect 45 108 46 109
rect 44 108 45 109
rect 43 108 44 109
rect 42 108 43 109
rect 41 108 42 109
rect 40 108 41 109
rect 39 108 40 109
rect 38 108 39 109
rect 37 108 38 109
rect 36 108 37 109
rect 35 108 36 109
rect 34 108 35 109
rect 33 108 34 109
rect 32 108 33 109
rect 27 108 28 109
rect 26 108 27 109
rect 25 108 26 109
rect 24 108 25 109
rect 23 108 24 109
rect 22 108 23 109
rect 21 108 22 109
rect 20 108 21 109
rect 19 108 20 109
rect 14 108 15 109
rect 13 108 14 109
rect 12 108 13 109
rect 11 108 12 109
rect 10 108 11 109
rect 9 108 10 109
rect 8 108 9 109
rect 7 108 8 109
rect 6 108 7 109
rect 127 109 128 110
rect 126 109 127 110
rect 125 109 126 110
rect 124 109 125 110
rect 123 109 124 110
rect 122 109 123 110
rect 121 109 122 110
rect 120 109 121 110
rect 119 109 120 110
rect 118 109 119 110
rect 117 109 118 110
rect 116 109 117 110
rect 115 109 116 110
rect 114 109 115 110
rect 113 109 114 110
rect 112 109 113 110
rect 111 109 112 110
rect 110 109 111 110
rect 109 109 110 110
rect 108 109 109 110
rect 107 109 108 110
rect 106 109 107 110
rect 105 109 106 110
rect 104 109 105 110
rect 103 109 104 110
rect 102 109 103 110
rect 101 109 102 110
rect 100 109 101 110
rect 99 109 100 110
rect 98 109 99 110
rect 97 109 98 110
rect 96 109 97 110
rect 77 109 78 110
rect 76 109 77 110
rect 75 109 76 110
rect 74 109 75 110
rect 73 109 74 110
rect 72 109 73 110
rect 71 109 72 110
rect 70 109 71 110
rect 69 109 70 110
rect 68 109 69 110
rect 67 109 68 110
rect 66 109 67 110
rect 65 109 66 110
rect 64 109 65 110
rect 63 109 64 110
rect 62 109 63 110
rect 61 109 62 110
rect 60 109 61 110
rect 59 109 60 110
rect 58 109 59 110
rect 57 109 58 110
rect 56 109 57 110
rect 55 109 56 110
rect 54 109 55 110
rect 49 109 50 110
rect 48 109 49 110
rect 47 109 48 110
rect 46 109 47 110
rect 45 109 46 110
rect 44 109 45 110
rect 43 109 44 110
rect 42 109 43 110
rect 41 109 42 110
rect 40 109 41 110
rect 39 109 40 110
rect 38 109 39 110
rect 37 109 38 110
rect 36 109 37 110
rect 35 109 36 110
rect 34 109 35 110
rect 33 109 34 110
rect 27 109 28 110
rect 26 109 27 110
rect 25 109 26 110
rect 24 109 25 110
rect 23 109 24 110
rect 22 109 23 110
rect 21 109 22 110
rect 20 109 21 110
rect 19 109 20 110
rect 14 109 15 110
rect 13 109 14 110
rect 12 109 13 110
rect 11 109 12 110
rect 10 109 11 110
rect 9 109 10 110
rect 8 109 9 110
rect 7 109 8 110
rect 6 109 7 110
rect 126 110 127 111
rect 125 110 126 111
rect 124 110 125 111
rect 123 110 124 111
rect 122 110 123 111
rect 121 110 122 111
rect 120 110 121 111
rect 119 110 120 111
rect 118 110 119 111
rect 117 110 118 111
rect 116 110 117 111
rect 115 110 116 111
rect 114 110 115 111
rect 113 110 114 111
rect 112 110 113 111
rect 111 110 112 111
rect 110 110 111 111
rect 109 110 110 111
rect 108 110 109 111
rect 107 110 108 111
rect 106 110 107 111
rect 105 110 106 111
rect 104 110 105 111
rect 103 110 104 111
rect 102 110 103 111
rect 101 110 102 111
rect 100 110 101 111
rect 99 110 100 111
rect 98 110 99 111
rect 97 110 98 111
rect 96 110 97 111
rect 87 110 88 111
rect 86 110 87 111
rect 82 110 83 111
rect 81 110 82 111
rect 80 110 81 111
rect 79 110 80 111
rect 78 110 79 111
rect 77 110 78 111
rect 76 110 77 111
rect 75 110 76 111
rect 74 110 75 111
rect 73 110 74 111
rect 72 110 73 111
rect 71 110 72 111
rect 70 110 71 111
rect 69 110 70 111
rect 68 110 69 111
rect 67 110 68 111
rect 66 110 67 111
rect 65 110 66 111
rect 64 110 65 111
rect 63 110 64 111
rect 62 110 63 111
rect 61 110 62 111
rect 60 110 61 111
rect 59 110 60 111
rect 58 110 59 111
rect 57 110 58 111
rect 56 110 57 111
rect 55 110 56 111
rect 54 110 55 111
rect 49 110 50 111
rect 48 110 49 111
rect 47 110 48 111
rect 46 110 47 111
rect 45 110 46 111
rect 44 110 45 111
rect 43 110 44 111
rect 42 110 43 111
rect 41 110 42 111
rect 40 110 41 111
rect 39 110 40 111
rect 38 110 39 111
rect 37 110 38 111
rect 36 110 37 111
rect 35 110 36 111
rect 34 110 35 111
rect 27 110 28 111
rect 26 110 27 111
rect 25 110 26 111
rect 24 110 25 111
rect 23 110 24 111
rect 22 110 23 111
rect 21 110 22 111
rect 20 110 21 111
rect 19 110 20 111
rect 15 110 16 111
rect 14 110 15 111
rect 13 110 14 111
rect 12 110 13 111
rect 11 110 12 111
rect 10 110 11 111
rect 9 110 10 111
rect 8 110 9 111
rect 7 110 8 111
rect 6 110 7 111
rect 125 111 126 112
rect 124 111 125 112
rect 123 111 124 112
rect 122 111 123 112
rect 121 111 122 112
rect 120 111 121 112
rect 119 111 120 112
rect 118 111 119 112
rect 117 111 118 112
rect 116 111 117 112
rect 115 111 116 112
rect 114 111 115 112
rect 113 111 114 112
rect 112 111 113 112
rect 111 111 112 112
rect 110 111 111 112
rect 109 111 110 112
rect 108 111 109 112
rect 107 111 108 112
rect 106 111 107 112
rect 105 111 106 112
rect 104 111 105 112
rect 103 111 104 112
rect 102 111 103 112
rect 101 111 102 112
rect 100 111 101 112
rect 99 111 100 112
rect 98 111 99 112
rect 97 111 98 112
rect 96 111 97 112
rect 87 111 88 112
rect 86 111 87 112
rect 85 111 86 112
rect 84 111 85 112
rect 83 111 84 112
rect 82 111 83 112
rect 81 111 82 112
rect 80 111 81 112
rect 79 111 80 112
rect 78 111 79 112
rect 77 111 78 112
rect 76 111 77 112
rect 75 111 76 112
rect 74 111 75 112
rect 73 111 74 112
rect 72 111 73 112
rect 71 111 72 112
rect 70 111 71 112
rect 69 111 70 112
rect 68 111 69 112
rect 67 111 68 112
rect 66 111 67 112
rect 65 111 66 112
rect 64 111 65 112
rect 63 111 64 112
rect 62 111 63 112
rect 61 111 62 112
rect 60 111 61 112
rect 59 111 60 112
rect 58 111 59 112
rect 57 111 58 112
rect 56 111 57 112
rect 55 111 56 112
rect 49 111 50 112
rect 48 111 49 112
rect 47 111 48 112
rect 46 111 47 112
rect 45 111 46 112
rect 44 111 45 112
rect 43 111 44 112
rect 42 111 43 112
rect 41 111 42 112
rect 40 111 41 112
rect 39 111 40 112
rect 38 111 39 112
rect 37 111 38 112
rect 36 111 37 112
rect 35 111 36 112
rect 34 111 35 112
rect 28 111 29 112
rect 27 111 28 112
rect 26 111 27 112
rect 25 111 26 112
rect 24 111 25 112
rect 23 111 24 112
rect 22 111 23 112
rect 21 111 22 112
rect 20 111 21 112
rect 19 111 20 112
rect 15 111 16 112
rect 14 111 15 112
rect 13 111 14 112
rect 12 111 13 112
rect 11 111 12 112
rect 10 111 11 112
rect 9 111 10 112
rect 8 111 9 112
rect 7 111 8 112
rect 6 111 7 112
rect 189 112 190 113
rect 124 112 125 113
rect 123 112 124 113
rect 122 112 123 113
rect 121 112 122 113
rect 120 112 121 113
rect 119 112 120 113
rect 118 112 119 113
rect 117 112 118 113
rect 116 112 117 113
rect 115 112 116 113
rect 114 112 115 113
rect 113 112 114 113
rect 112 112 113 113
rect 111 112 112 113
rect 110 112 111 113
rect 109 112 110 113
rect 108 112 109 113
rect 107 112 108 113
rect 106 112 107 113
rect 105 112 106 113
rect 104 112 105 113
rect 103 112 104 113
rect 102 112 103 113
rect 101 112 102 113
rect 100 112 101 113
rect 99 112 100 113
rect 98 112 99 113
rect 97 112 98 113
rect 96 112 97 113
rect 95 112 96 113
rect 87 112 88 113
rect 86 112 87 113
rect 85 112 86 113
rect 84 112 85 113
rect 83 112 84 113
rect 82 112 83 113
rect 81 112 82 113
rect 80 112 81 113
rect 79 112 80 113
rect 78 112 79 113
rect 77 112 78 113
rect 76 112 77 113
rect 75 112 76 113
rect 74 112 75 113
rect 73 112 74 113
rect 72 112 73 113
rect 71 112 72 113
rect 70 112 71 113
rect 69 112 70 113
rect 68 112 69 113
rect 67 112 68 113
rect 66 112 67 113
rect 65 112 66 113
rect 64 112 65 113
rect 63 112 64 113
rect 62 112 63 113
rect 61 112 62 113
rect 60 112 61 113
rect 59 112 60 113
rect 58 112 59 113
rect 57 112 58 113
rect 56 112 57 113
rect 55 112 56 113
rect 49 112 50 113
rect 48 112 49 113
rect 47 112 48 113
rect 46 112 47 113
rect 45 112 46 113
rect 44 112 45 113
rect 43 112 44 113
rect 42 112 43 113
rect 41 112 42 113
rect 40 112 41 113
rect 39 112 40 113
rect 38 112 39 113
rect 37 112 38 113
rect 36 112 37 113
rect 35 112 36 113
rect 28 112 29 113
rect 27 112 28 113
rect 26 112 27 113
rect 25 112 26 113
rect 24 112 25 113
rect 23 112 24 113
rect 22 112 23 113
rect 21 112 22 113
rect 20 112 21 113
rect 15 112 16 113
rect 14 112 15 113
rect 13 112 14 113
rect 12 112 13 113
rect 11 112 12 113
rect 10 112 11 113
rect 9 112 10 113
rect 8 112 9 113
rect 7 112 8 113
rect 6 112 7 113
rect 197 113 198 114
rect 196 113 197 114
rect 195 113 196 114
rect 194 113 195 114
rect 193 113 194 114
rect 192 113 193 114
rect 191 113 192 114
rect 190 113 191 114
rect 189 113 190 114
rect 124 113 125 114
rect 123 113 124 114
rect 122 113 123 114
rect 121 113 122 114
rect 120 113 121 114
rect 119 113 120 114
rect 118 113 119 114
rect 117 113 118 114
rect 116 113 117 114
rect 115 113 116 114
rect 114 113 115 114
rect 113 113 114 114
rect 112 113 113 114
rect 111 113 112 114
rect 110 113 111 114
rect 109 113 110 114
rect 108 113 109 114
rect 107 113 108 114
rect 106 113 107 114
rect 105 113 106 114
rect 104 113 105 114
rect 103 113 104 114
rect 102 113 103 114
rect 101 113 102 114
rect 100 113 101 114
rect 99 113 100 114
rect 98 113 99 114
rect 97 113 98 114
rect 96 113 97 114
rect 95 113 96 114
rect 86 113 87 114
rect 85 113 86 114
rect 84 113 85 114
rect 83 113 84 114
rect 82 113 83 114
rect 81 113 82 114
rect 80 113 81 114
rect 79 113 80 114
rect 78 113 79 114
rect 77 113 78 114
rect 76 113 77 114
rect 75 113 76 114
rect 74 113 75 114
rect 73 113 74 114
rect 72 113 73 114
rect 71 113 72 114
rect 70 113 71 114
rect 69 113 70 114
rect 68 113 69 114
rect 67 113 68 114
rect 66 113 67 114
rect 65 113 66 114
rect 64 113 65 114
rect 63 113 64 114
rect 62 113 63 114
rect 61 113 62 114
rect 60 113 61 114
rect 59 113 60 114
rect 58 113 59 114
rect 57 113 58 114
rect 56 113 57 114
rect 55 113 56 114
rect 49 113 50 114
rect 48 113 49 114
rect 47 113 48 114
rect 46 113 47 114
rect 45 113 46 114
rect 44 113 45 114
rect 43 113 44 114
rect 42 113 43 114
rect 41 113 42 114
rect 40 113 41 114
rect 39 113 40 114
rect 38 113 39 114
rect 37 113 38 114
rect 36 113 37 114
rect 29 113 30 114
rect 28 113 29 114
rect 27 113 28 114
rect 26 113 27 114
rect 25 113 26 114
rect 24 113 25 114
rect 23 113 24 114
rect 22 113 23 114
rect 21 113 22 114
rect 20 113 21 114
rect 15 113 16 114
rect 14 113 15 114
rect 13 113 14 114
rect 12 113 13 114
rect 11 113 12 114
rect 10 113 11 114
rect 9 113 10 114
rect 8 113 9 114
rect 7 113 8 114
rect 6 113 7 114
rect 197 114 198 115
rect 196 114 197 115
rect 195 114 196 115
rect 194 114 195 115
rect 193 114 194 115
rect 192 114 193 115
rect 191 114 192 115
rect 190 114 191 115
rect 189 114 190 115
rect 123 114 124 115
rect 122 114 123 115
rect 121 114 122 115
rect 120 114 121 115
rect 119 114 120 115
rect 118 114 119 115
rect 117 114 118 115
rect 116 114 117 115
rect 115 114 116 115
rect 114 114 115 115
rect 113 114 114 115
rect 112 114 113 115
rect 111 114 112 115
rect 110 114 111 115
rect 109 114 110 115
rect 108 114 109 115
rect 107 114 108 115
rect 106 114 107 115
rect 105 114 106 115
rect 104 114 105 115
rect 103 114 104 115
rect 102 114 103 115
rect 101 114 102 115
rect 100 114 101 115
rect 99 114 100 115
rect 98 114 99 115
rect 97 114 98 115
rect 96 114 97 115
rect 95 114 96 115
rect 86 114 87 115
rect 85 114 86 115
rect 84 114 85 115
rect 83 114 84 115
rect 82 114 83 115
rect 81 114 82 115
rect 80 114 81 115
rect 79 114 80 115
rect 78 114 79 115
rect 77 114 78 115
rect 76 114 77 115
rect 75 114 76 115
rect 74 114 75 115
rect 73 114 74 115
rect 72 114 73 115
rect 71 114 72 115
rect 70 114 71 115
rect 69 114 70 115
rect 68 114 69 115
rect 67 114 68 115
rect 66 114 67 115
rect 65 114 66 115
rect 64 114 65 115
rect 63 114 64 115
rect 62 114 63 115
rect 61 114 62 115
rect 60 114 61 115
rect 59 114 60 115
rect 58 114 59 115
rect 57 114 58 115
rect 56 114 57 115
rect 50 114 51 115
rect 49 114 50 115
rect 48 114 49 115
rect 47 114 48 115
rect 46 114 47 115
rect 45 114 46 115
rect 44 114 45 115
rect 43 114 44 115
rect 42 114 43 115
rect 41 114 42 115
rect 40 114 41 115
rect 39 114 40 115
rect 38 114 39 115
rect 37 114 38 115
rect 36 114 37 115
rect 29 114 30 115
rect 28 114 29 115
rect 27 114 28 115
rect 26 114 27 115
rect 25 114 26 115
rect 24 114 25 115
rect 23 114 24 115
rect 22 114 23 115
rect 21 114 22 115
rect 20 114 21 115
rect 15 114 16 115
rect 14 114 15 115
rect 13 114 14 115
rect 12 114 13 115
rect 11 114 12 115
rect 10 114 11 115
rect 9 114 10 115
rect 8 114 9 115
rect 7 114 8 115
rect 6 114 7 115
rect 196 115 197 116
rect 189 115 190 116
rect 180 115 181 116
rect 163 115 164 116
rect 122 115 123 116
rect 121 115 122 116
rect 120 115 121 116
rect 119 115 120 116
rect 118 115 119 116
rect 117 115 118 116
rect 116 115 117 116
rect 115 115 116 116
rect 114 115 115 116
rect 113 115 114 116
rect 112 115 113 116
rect 111 115 112 116
rect 110 115 111 116
rect 109 115 110 116
rect 108 115 109 116
rect 107 115 108 116
rect 106 115 107 116
rect 105 115 106 116
rect 104 115 105 116
rect 103 115 104 116
rect 102 115 103 116
rect 101 115 102 116
rect 100 115 101 116
rect 99 115 100 116
rect 98 115 99 116
rect 97 115 98 116
rect 96 115 97 116
rect 95 115 96 116
rect 94 115 95 116
rect 85 115 86 116
rect 84 115 85 116
rect 83 115 84 116
rect 82 115 83 116
rect 81 115 82 116
rect 80 115 81 116
rect 79 115 80 116
rect 78 115 79 116
rect 77 115 78 116
rect 76 115 77 116
rect 75 115 76 116
rect 74 115 75 116
rect 73 115 74 116
rect 72 115 73 116
rect 71 115 72 116
rect 70 115 71 116
rect 69 115 70 116
rect 68 115 69 116
rect 67 115 68 116
rect 66 115 67 116
rect 65 115 66 116
rect 64 115 65 116
rect 63 115 64 116
rect 62 115 63 116
rect 61 115 62 116
rect 60 115 61 116
rect 59 115 60 116
rect 58 115 59 116
rect 57 115 58 116
rect 56 115 57 116
rect 50 115 51 116
rect 49 115 50 116
rect 48 115 49 116
rect 47 115 48 116
rect 46 115 47 116
rect 45 115 46 116
rect 44 115 45 116
rect 43 115 44 116
rect 42 115 43 116
rect 41 115 42 116
rect 40 115 41 116
rect 39 115 40 116
rect 38 115 39 116
rect 37 115 38 116
rect 30 115 31 116
rect 29 115 30 116
rect 28 115 29 116
rect 27 115 28 116
rect 26 115 27 116
rect 25 115 26 116
rect 24 115 25 116
rect 23 115 24 116
rect 22 115 23 116
rect 21 115 22 116
rect 20 115 21 116
rect 16 115 17 116
rect 15 115 16 116
rect 14 115 15 116
rect 13 115 14 116
rect 12 115 13 116
rect 11 115 12 116
rect 10 115 11 116
rect 9 115 10 116
rect 8 115 9 116
rect 7 115 8 116
rect 6 115 7 116
rect 180 116 181 117
rect 164 116 165 117
rect 163 116 164 117
rect 121 116 122 117
rect 120 116 121 117
rect 119 116 120 117
rect 118 116 119 117
rect 117 116 118 117
rect 116 116 117 117
rect 115 116 116 117
rect 114 116 115 117
rect 113 116 114 117
rect 112 116 113 117
rect 111 116 112 117
rect 110 116 111 117
rect 109 116 110 117
rect 108 116 109 117
rect 107 116 108 117
rect 106 116 107 117
rect 105 116 106 117
rect 104 116 105 117
rect 103 116 104 117
rect 102 116 103 117
rect 101 116 102 117
rect 100 116 101 117
rect 99 116 100 117
rect 98 116 99 117
rect 97 116 98 117
rect 96 116 97 117
rect 95 116 96 117
rect 94 116 95 117
rect 85 116 86 117
rect 84 116 85 117
rect 83 116 84 117
rect 82 116 83 117
rect 81 116 82 117
rect 80 116 81 117
rect 79 116 80 117
rect 78 116 79 117
rect 77 116 78 117
rect 76 116 77 117
rect 75 116 76 117
rect 74 116 75 117
rect 73 116 74 117
rect 72 116 73 117
rect 71 116 72 117
rect 70 116 71 117
rect 69 116 70 117
rect 68 116 69 117
rect 67 116 68 117
rect 66 116 67 117
rect 65 116 66 117
rect 64 116 65 117
rect 63 116 64 117
rect 62 116 63 117
rect 61 116 62 117
rect 60 116 61 117
rect 59 116 60 117
rect 58 116 59 117
rect 57 116 58 117
rect 56 116 57 117
rect 50 116 51 117
rect 49 116 50 117
rect 48 116 49 117
rect 47 116 48 117
rect 46 116 47 117
rect 45 116 46 117
rect 44 116 45 117
rect 43 116 44 117
rect 42 116 43 117
rect 41 116 42 117
rect 40 116 41 117
rect 39 116 40 117
rect 38 116 39 117
rect 37 116 38 117
rect 30 116 31 117
rect 29 116 30 117
rect 28 116 29 117
rect 27 116 28 117
rect 26 116 27 117
rect 25 116 26 117
rect 24 116 25 117
rect 23 116 24 117
rect 22 116 23 117
rect 21 116 22 117
rect 20 116 21 117
rect 16 116 17 117
rect 15 116 16 117
rect 14 116 15 117
rect 13 116 14 117
rect 12 116 13 117
rect 11 116 12 117
rect 10 116 11 117
rect 9 116 10 117
rect 8 116 9 117
rect 7 116 8 117
rect 6 116 7 117
rect 180 117 181 118
rect 179 117 180 118
rect 178 117 179 118
rect 177 117 178 118
rect 176 117 177 118
rect 175 117 176 118
rect 174 117 175 118
rect 173 117 174 118
rect 172 117 173 118
rect 171 117 172 118
rect 170 117 171 118
rect 169 117 170 118
rect 168 117 169 118
rect 167 117 168 118
rect 166 117 167 118
rect 165 117 166 118
rect 164 117 165 118
rect 163 117 164 118
rect 121 117 122 118
rect 120 117 121 118
rect 119 117 120 118
rect 118 117 119 118
rect 117 117 118 118
rect 116 117 117 118
rect 115 117 116 118
rect 114 117 115 118
rect 113 117 114 118
rect 112 117 113 118
rect 111 117 112 118
rect 110 117 111 118
rect 109 117 110 118
rect 108 117 109 118
rect 107 117 108 118
rect 106 117 107 118
rect 105 117 106 118
rect 104 117 105 118
rect 103 117 104 118
rect 102 117 103 118
rect 101 117 102 118
rect 100 117 101 118
rect 99 117 100 118
rect 98 117 99 118
rect 97 117 98 118
rect 96 117 97 118
rect 95 117 96 118
rect 94 117 95 118
rect 93 117 94 118
rect 84 117 85 118
rect 83 117 84 118
rect 82 117 83 118
rect 81 117 82 118
rect 80 117 81 118
rect 79 117 80 118
rect 78 117 79 118
rect 77 117 78 118
rect 76 117 77 118
rect 75 117 76 118
rect 74 117 75 118
rect 73 117 74 118
rect 72 117 73 118
rect 71 117 72 118
rect 70 117 71 118
rect 69 117 70 118
rect 68 117 69 118
rect 67 117 68 118
rect 66 117 67 118
rect 65 117 66 118
rect 64 117 65 118
rect 63 117 64 118
rect 62 117 63 118
rect 61 117 62 118
rect 60 117 61 118
rect 59 117 60 118
rect 58 117 59 118
rect 57 117 58 118
rect 50 117 51 118
rect 49 117 50 118
rect 48 117 49 118
rect 47 117 48 118
rect 46 117 47 118
rect 45 117 46 118
rect 44 117 45 118
rect 43 117 44 118
rect 42 117 43 118
rect 41 117 42 118
rect 40 117 41 118
rect 39 117 40 118
rect 38 117 39 118
rect 37 117 38 118
rect 30 117 31 118
rect 29 117 30 118
rect 28 117 29 118
rect 27 117 28 118
rect 26 117 27 118
rect 25 117 26 118
rect 24 117 25 118
rect 23 117 24 118
rect 22 117 23 118
rect 21 117 22 118
rect 20 117 21 118
rect 16 117 17 118
rect 15 117 16 118
rect 14 117 15 118
rect 13 117 14 118
rect 12 117 13 118
rect 11 117 12 118
rect 10 117 11 118
rect 9 117 10 118
rect 8 117 9 118
rect 7 117 8 118
rect 6 117 7 118
rect 180 118 181 119
rect 179 118 180 119
rect 178 118 179 119
rect 177 118 178 119
rect 176 118 177 119
rect 175 118 176 119
rect 174 118 175 119
rect 173 118 174 119
rect 172 118 173 119
rect 171 118 172 119
rect 170 118 171 119
rect 169 118 170 119
rect 168 118 169 119
rect 167 118 168 119
rect 166 118 167 119
rect 165 118 166 119
rect 164 118 165 119
rect 163 118 164 119
rect 120 118 121 119
rect 119 118 120 119
rect 118 118 119 119
rect 117 118 118 119
rect 116 118 117 119
rect 115 118 116 119
rect 114 118 115 119
rect 113 118 114 119
rect 112 118 113 119
rect 111 118 112 119
rect 110 118 111 119
rect 109 118 110 119
rect 108 118 109 119
rect 107 118 108 119
rect 106 118 107 119
rect 105 118 106 119
rect 104 118 105 119
rect 103 118 104 119
rect 102 118 103 119
rect 101 118 102 119
rect 100 118 101 119
rect 99 118 100 119
rect 98 118 99 119
rect 97 118 98 119
rect 96 118 97 119
rect 95 118 96 119
rect 94 118 95 119
rect 93 118 94 119
rect 84 118 85 119
rect 83 118 84 119
rect 82 118 83 119
rect 81 118 82 119
rect 80 118 81 119
rect 79 118 80 119
rect 78 118 79 119
rect 77 118 78 119
rect 76 118 77 119
rect 75 118 76 119
rect 74 118 75 119
rect 73 118 74 119
rect 72 118 73 119
rect 71 118 72 119
rect 70 118 71 119
rect 69 118 70 119
rect 68 118 69 119
rect 67 118 68 119
rect 66 118 67 119
rect 65 118 66 119
rect 64 118 65 119
rect 63 118 64 119
rect 62 118 63 119
rect 61 118 62 119
rect 60 118 61 119
rect 59 118 60 119
rect 58 118 59 119
rect 57 118 58 119
rect 51 118 52 119
rect 50 118 51 119
rect 49 118 50 119
rect 48 118 49 119
rect 47 118 48 119
rect 46 118 47 119
rect 45 118 46 119
rect 44 118 45 119
rect 43 118 44 119
rect 42 118 43 119
rect 41 118 42 119
rect 40 118 41 119
rect 39 118 40 119
rect 38 118 39 119
rect 37 118 38 119
rect 31 118 32 119
rect 30 118 31 119
rect 29 118 30 119
rect 28 118 29 119
rect 27 118 28 119
rect 26 118 27 119
rect 25 118 26 119
rect 24 118 25 119
rect 23 118 24 119
rect 22 118 23 119
rect 21 118 22 119
rect 20 118 21 119
rect 16 118 17 119
rect 15 118 16 119
rect 14 118 15 119
rect 13 118 14 119
rect 12 118 13 119
rect 11 118 12 119
rect 10 118 11 119
rect 9 118 10 119
rect 8 118 9 119
rect 7 118 8 119
rect 6 118 7 119
rect 190 119 191 120
rect 189 119 190 120
rect 180 119 181 120
rect 179 119 180 120
rect 178 119 179 120
rect 177 119 178 120
rect 176 119 177 120
rect 175 119 176 120
rect 174 119 175 120
rect 173 119 174 120
rect 172 119 173 120
rect 171 119 172 120
rect 170 119 171 120
rect 169 119 170 120
rect 168 119 169 120
rect 167 119 168 120
rect 166 119 167 120
rect 165 119 166 120
rect 164 119 165 120
rect 163 119 164 120
rect 119 119 120 120
rect 118 119 119 120
rect 117 119 118 120
rect 116 119 117 120
rect 115 119 116 120
rect 114 119 115 120
rect 113 119 114 120
rect 112 119 113 120
rect 111 119 112 120
rect 110 119 111 120
rect 109 119 110 120
rect 108 119 109 120
rect 107 119 108 120
rect 106 119 107 120
rect 105 119 106 120
rect 104 119 105 120
rect 103 119 104 120
rect 102 119 103 120
rect 101 119 102 120
rect 100 119 101 120
rect 99 119 100 120
rect 98 119 99 120
rect 97 119 98 120
rect 96 119 97 120
rect 95 119 96 120
rect 94 119 95 120
rect 93 119 94 120
rect 92 119 93 120
rect 83 119 84 120
rect 82 119 83 120
rect 81 119 82 120
rect 80 119 81 120
rect 79 119 80 120
rect 78 119 79 120
rect 77 119 78 120
rect 76 119 77 120
rect 75 119 76 120
rect 74 119 75 120
rect 73 119 74 120
rect 72 119 73 120
rect 71 119 72 120
rect 70 119 71 120
rect 69 119 70 120
rect 68 119 69 120
rect 67 119 68 120
rect 66 119 67 120
rect 65 119 66 120
rect 64 119 65 120
rect 63 119 64 120
rect 62 119 63 120
rect 61 119 62 120
rect 60 119 61 120
rect 59 119 60 120
rect 58 119 59 120
rect 51 119 52 120
rect 50 119 51 120
rect 49 119 50 120
rect 48 119 49 120
rect 47 119 48 120
rect 46 119 47 120
rect 45 119 46 120
rect 44 119 45 120
rect 43 119 44 120
rect 42 119 43 120
rect 41 119 42 120
rect 40 119 41 120
rect 39 119 40 120
rect 38 119 39 120
rect 31 119 32 120
rect 30 119 31 120
rect 29 119 30 120
rect 28 119 29 120
rect 27 119 28 120
rect 26 119 27 120
rect 25 119 26 120
rect 24 119 25 120
rect 23 119 24 120
rect 22 119 23 120
rect 21 119 22 120
rect 20 119 21 120
rect 16 119 17 120
rect 15 119 16 120
rect 14 119 15 120
rect 13 119 14 120
rect 12 119 13 120
rect 11 119 12 120
rect 10 119 11 120
rect 9 119 10 120
rect 8 119 9 120
rect 7 119 8 120
rect 6 119 7 120
rect 189 120 190 121
rect 180 120 181 121
rect 179 120 180 121
rect 178 120 179 121
rect 177 120 178 121
rect 176 120 177 121
rect 175 120 176 121
rect 174 120 175 121
rect 173 120 174 121
rect 172 120 173 121
rect 171 120 172 121
rect 170 120 171 121
rect 169 120 170 121
rect 168 120 169 121
rect 167 120 168 121
rect 166 120 167 121
rect 165 120 166 121
rect 164 120 165 121
rect 163 120 164 121
rect 118 120 119 121
rect 117 120 118 121
rect 116 120 117 121
rect 115 120 116 121
rect 114 120 115 121
rect 113 120 114 121
rect 112 120 113 121
rect 111 120 112 121
rect 110 120 111 121
rect 109 120 110 121
rect 108 120 109 121
rect 107 120 108 121
rect 106 120 107 121
rect 105 120 106 121
rect 104 120 105 121
rect 103 120 104 121
rect 102 120 103 121
rect 101 120 102 121
rect 100 120 101 121
rect 99 120 100 121
rect 98 120 99 121
rect 97 120 98 121
rect 96 120 97 121
rect 95 120 96 121
rect 94 120 95 121
rect 93 120 94 121
rect 92 120 93 121
rect 82 120 83 121
rect 81 120 82 121
rect 80 120 81 121
rect 79 120 80 121
rect 78 120 79 121
rect 77 120 78 121
rect 76 120 77 121
rect 75 120 76 121
rect 74 120 75 121
rect 73 120 74 121
rect 72 120 73 121
rect 71 120 72 121
rect 70 120 71 121
rect 69 120 70 121
rect 68 120 69 121
rect 67 120 68 121
rect 66 120 67 121
rect 65 120 66 121
rect 64 120 65 121
rect 63 120 64 121
rect 62 120 63 121
rect 61 120 62 121
rect 60 120 61 121
rect 59 120 60 121
rect 58 120 59 121
rect 51 120 52 121
rect 50 120 51 121
rect 49 120 50 121
rect 48 120 49 121
rect 47 120 48 121
rect 46 120 47 121
rect 45 120 46 121
rect 44 120 45 121
rect 43 120 44 121
rect 42 120 43 121
rect 41 120 42 121
rect 40 120 41 121
rect 39 120 40 121
rect 38 120 39 121
rect 31 120 32 121
rect 30 120 31 121
rect 29 120 30 121
rect 28 120 29 121
rect 27 120 28 121
rect 26 120 27 121
rect 25 120 26 121
rect 24 120 25 121
rect 23 120 24 121
rect 22 120 23 121
rect 21 120 22 121
rect 20 120 21 121
rect 17 120 18 121
rect 16 120 17 121
rect 15 120 16 121
rect 14 120 15 121
rect 13 120 14 121
rect 12 120 13 121
rect 11 120 12 121
rect 10 120 11 121
rect 9 120 10 121
rect 8 120 9 121
rect 7 120 8 121
rect 6 120 7 121
rect 180 121 181 122
rect 179 121 180 122
rect 172 121 173 122
rect 171 121 172 122
rect 170 121 171 122
rect 165 121 166 122
rect 164 121 165 122
rect 163 121 164 122
rect 117 121 118 122
rect 116 121 117 122
rect 115 121 116 122
rect 114 121 115 122
rect 113 121 114 122
rect 112 121 113 122
rect 111 121 112 122
rect 110 121 111 122
rect 109 121 110 122
rect 108 121 109 122
rect 107 121 108 122
rect 106 121 107 122
rect 105 121 106 122
rect 104 121 105 122
rect 103 121 104 122
rect 102 121 103 122
rect 101 121 102 122
rect 100 121 101 122
rect 99 121 100 122
rect 98 121 99 122
rect 97 121 98 122
rect 96 121 97 122
rect 95 121 96 122
rect 94 121 95 122
rect 93 121 94 122
rect 92 121 93 122
rect 91 121 92 122
rect 82 121 83 122
rect 81 121 82 122
rect 80 121 81 122
rect 79 121 80 122
rect 78 121 79 122
rect 77 121 78 122
rect 76 121 77 122
rect 75 121 76 122
rect 74 121 75 122
rect 73 121 74 122
rect 72 121 73 122
rect 71 121 72 122
rect 70 121 71 122
rect 69 121 70 122
rect 68 121 69 122
rect 67 121 68 122
rect 66 121 67 122
rect 65 121 66 122
rect 64 121 65 122
rect 63 121 64 122
rect 62 121 63 122
rect 61 121 62 122
rect 60 121 61 122
rect 59 121 60 122
rect 52 121 53 122
rect 51 121 52 122
rect 50 121 51 122
rect 49 121 50 122
rect 48 121 49 122
rect 47 121 48 122
rect 46 121 47 122
rect 45 121 46 122
rect 44 121 45 122
rect 43 121 44 122
rect 42 121 43 122
rect 41 121 42 122
rect 40 121 41 122
rect 39 121 40 122
rect 38 121 39 122
rect 32 121 33 122
rect 31 121 32 122
rect 30 121 31 122
rect 29 121 30 122
rect 28 121 29 122
rect 27 121 28 122
rect 26 121 27 122
rect 25 121 26 122
rect 24 121 25 122
rect 23 121 24 122
rect 22 121 23 122
rect 21 121 22 122
rect 20 121 21 122
rect 17 121 18 122
rect 16 121 17 122
rect 15 121 16 122
rect 14 121 15 122
rect 13 121 14 122
rect 12 121 13 122
rect 11 121 12 122
rect 10 121 11 122
rect 9 121 10 122
rect 8 121 9 122
rect 7 121 8 122
rect 6 121 7 122
rect 197 122 198 123
rect 196 122 197 123
rect 195 122 196 123
rect 194 122 195 123
rect 193 122 194 123
rect 192 122 193 123
rect 191 122 192 123
rect 190 122 191 123
rect 189 122 190 123
rect 180 122 181 123
rect 171 122 172 123
rect 170 122 171 123
rect 163 122 164 123
rect 116 122 117 123
rect 115 122 116 123
rect 114 122 115 123
rect 113 122 114 123
rect 112 122 113 123
rect 111 122 112 123
rect 110 122 111 123
rect 109 122 110 123
rect 108 122 109 123
rect 107 122 108 123
rect 106 122 107 123
rect 105 122 106 123
rect 104 122 105 123
rect 103 122 104 123
rect 102 122 103 123
rect 101 122 102 123
rect 100 122 101 123
rect 99 122 100 123
rect 98 122 99 123
rect 97 122 98 123
rect 96 122 97 123
rect 95 122 96 123
rect 94 122 95 123
rect 93 122 94 123
rect 92 122 93 123
rect 91 122 92 123
rect 90 122 91 123
rect 81 122 82 123
rect 80 122 81 123
rect 79 122 80 123
rect 78 122 79 123
rect 77 122 78 123
rect 76 122 77 123
rect 75 122 76 123
rect 74 122 75 123
rect 73 122 74 123
rect 72 122 73 123
rect 71 122 72 123
rect 70 122 71 123
rect 69 122 70 123
rect 68 122 69 123
rect 67 122 68 123
rect 66 122 67 123
rect 65 122 66 123
rect 64 122 65 123
rect 63 122 64 123
rect 62 122 63 123
rect 61 122 62 123
rect 60 122 61 123
rect 59 122 60 123
rect 52 122 53 123
rect 51 122 52 123
rect 50 122 51 123
rect 49 122 50 123
rect 48 122 49 123
rect 47 122 48 123
rect 46 122 47 123
rect 45 122 46 123
rect 44 122 45 123
rect 43 122 44 123
rect 42 122 43 123
rect 41 122 42 123
rect 40 122 41 123
rect 39 122 40 123
rect 38 122 39 123
rect 32 122 33 123
rect 31 122 32 123
rect 30 122 31 123
rect 29 122 30 123
rect 28 122 29 123
rect 27 122 28 123
rect 26 122 27 123
rect 25 122 26 123
rect 24 122 25 123
rect 23 122 24 123
rect 22 122 23 123
rect 21 122 22 123
rect 17 122 18 123
rect 16 122 17 123
rect 15 122 16 123
rect 14 122 15 123
rect 13 122 14 123
rect 12 122 13 123
rect 11 122 12 123
rect 10 122 11 123
rect 9 122 10 123
rect 8 122 9 123
rect 7 122 8 123
rect 6 122 7 123
rect 196 123 197 124
rect 195 123 196 124
rect 194 123 195 124
rect 193 123 194 124
rect 192 123 193 124
rect 191 123 192 124
rect 190 123 191 124
rect 189 123 190 124
rect 180 123 181 124
rect 171 123 172 124
rect 170 123 171 124
rect 163 123 164 124
rect 115 123 116 124
rect 114 123 115 124
rect 113 123 114 124
rect 112 123 113 124
rect 111 123 112 124
rect 110 123 111 124
rect 109 123 110 124
rect 108 123 109 124
rect 107 123 108 124
rect 106 123 107 124
rect 105 123 106 124
rect 104 123 105 124
rect 103 123 104 124
rect 102 123 103 124
rect 101 123 102 124
rect 100 123 101 124
rect 99 123 100 124
rect 98 123 99 124
rect 97 123 98 124
rect 96 123 97 124
rect 95 123 96 124
rect 94 123 95 124
rect 93 123 94 124
rect 92 123 93 124
rect 91 123 92 124
rect 90 123 91 124
rect 80 123 81 124
rect 79 123 80 124
rect 78 123 79 124
rect 77 123 78 124
rect 76 123 77 124
rect 75 123 76 124
rect 74 123 75 124
rect 73 123 74 124
rect 72 123 73 124
rect 71 123 72 124
rect 70 123 71 124
rect 69 123 70 124
rect 68 123 69 124
rect 67 123 68 124
rect 66 123 67 124
rect 65 123 66 124
rect 64 123 65 124
rect 63 123 64 124
rect 62 123 63 124
rect 61 123 62 124
rect 60 123 61 124
rect 53 123 54 124
rect 52 123 53 124
rect 51 123 52 124
rect 50 123 51 124
rect 49 123 50 124
rect 48 123 49 124
rect 47 123 48 124
rect 46 123 47 124
rect 45 123 46 124
rect 44 123 45 124
rect 43 123 44 124
rect 42 123 43 124
rect 41 123 42 124
rect 40 123 41 124
rect 39 123 40 124
rect 32 123 33 124
rect 31 123 32 124
rect 30 123 31 124
rect 29 123 30 124
rect 28 123 29 124
rect 27 123 28 124
rect 26 123 27 124
rect 25 123 26 124
rect 24 123 25 124
rect 23 123 24 124
rect 22 123 23 124
rect 21 123 22 124
rect 17 123 18 124
rect 16 123 17 124
rect 15 123 16 124
rect 14 123 15 124
rect 13 123 14 124
rect 12 123 13 124
rect 11 123 12 124
rect 10 123 11 124
rect 9 123 10 124
rect 8 123 9 124
rect 7 123 8 124
rect 196 124 197 125
rect 194 124 195 125
rect 193 124 194 125
rect 192 124 193 125
rect 191 124 192 125
rect 189 124 190 125
rect 171 124 172 125
rect 170 124 171 125
rect 114 124 115 125
rect 113 124 114 125
rect 112 124 113 125
rect 111 124 112 125
rect 110 124 111 125
rect 109 124 110 125
rect 108 124 109 125
rect 107 124 108 125
rect 106 124 107 125
rect 105 124 106 125
rect 104 124 105 125
rect 103 124 104 125
rect 102 124 103 125
rect 101 124 102 125
rect 100 124 101 125
rect 99 124 100 125
rect 98 124 99 125
rect 97 124 98 125
rect 96 124 97 125
rect 95 124 96 125
rect 94 124 95 125
rect 93 124 94 125
rect 92 124 93 125
rect 91 124 92 125
rect 90 124 91 125
rect 89 124 90 125
rect 79 124 80 125
rect 78 124 79 125
rect 77 124 78 125
rect 76 124 77 125
rect 75 124 76 125
rect 74 124 75 125
rect 73 124 74 125
rect 72 124 73 125
rect 71 124 72 125
rect 70 124 71 125
rect 69 124 70 125
rect 68 124 69 125
rect 67 124 68 125
rect 66 124 67 125
rect 65 124 66 125
rect 64 124 65 125
rect 63 124 64 125
rect 62 124 63 125
rect 61 124 62 125
rect 53 124 54 125
rect 52 124 53 125
rect 51 124 52 125
rect 50 124 51 125
rect 49 124 50 125
rect 48 124 49 125
rect 47 124 48 125
rect 46 124 47 125
rect 45 124 46 125
rect 44 124 45 125
rect 43 124 44 125
rect 42 124 43 125
rect 41 124 42 125
rect 40 124 41 125
rect 39 124 40 125
rect 32 124 33 125
rect 31 124 32 125
rect 30 124 31 125
rect 29 124 30 125
rect 28 124 29 125
rect 27 124 28 125
rect 26 124 27 125
rect 25 124 26 125
rect 24 124 25 125
rect 23 124 24 125
rect 22 124 23 125
rect 21 124 22 125
rect 17 124 18 125
rect 16 124 17 125
rect 15 124 16 125
rect 14 124 15 125
rect 13 124 14 125
rect 12 124 13 125
rect 11 124 12 125
rect 10 124 11 125
rect 9 124 10 125
rect 8 124 9 125
rect 7 124 8 125
rect 189 125 190 126
rect 171 125 172 126
rect 170 125 171 126
rect 113 125 114 126
rect 112 125 113 126
rect 111 125 112 126
rect 110 125 111 126
rect 109 125 110 126
rect 108 125 109 126
rect 107 125 108 126
rect 106 125 107 126
rect 105 125 106 126
rect 104 125 105 126
rect 103 125 104 126
rect 102 125 103 126
rect 101 125 102 126
rect 100 125 101 126
rect 99 125 100 126
rect 98 125 99 126
rect 97 125 98 126
rect 96 125 97 126
rect 95 125 96 126
rect 94 125 95 126
rect 93 125 94 126
rect 92 125 93 126
rect 91 125 92 126
rect 90 125 91 126
rect 89 125 90 126
rect 88 125 89 126
rect 78 125 79 126
rect 77 125 78 126
rect 76 125 77 126
rect 75 125 76 126
rect 74 125 75 126
rect 73 125 74 126
rect 72 125 73 126
rect 71 125 72 126
rect 70 125 71 126
rect 69 125 70 126
rect 68 125 69 126
rect 67 125 68 126
rect 66 125 67 126
rect 65 125 66 126
rect 64 125 65 126
rect 63 125 64 126
rect 62 125 63 126
rect 53 125 54 126
rect 52 125 53 126
rect 51 125 52 126
rect 50 125 51 126
rect 49 125 50 126
rect 48 125 49 126
rect 47 125 48 126
rect 46 125 47 126
rect 45 125 46 126
rect 44 125 45 126
rect 43 125 44 126
rect 42 125 43 126
rect 41 125 42 126
rect 40 125 41 126
rect 39 125 40 126
rect 33 125 34 126
rect 32 125 33 126
rect 31 125 32 126
rect 30 125 31 126
rect 29 125 30 126
rect 28 125 29 126
rect 27 125 28 126
rect 26 125 27 126
rect 25 125 26 126
rect 24 125 25 126
rect 23 125 24 126
rect 22 125 23 126
rect 21 125 22 126
rect 17 125 18 126
rect 16 125 17 126
rect 15 125 16 126
rect 14 125 15 126
rect 13 125 14 126
rect 12 125 13 126
rect 11 125 12 126
rect 10 125 11 126
rect 9 125 10 126
rect 8 125 9 126
rect 7 125 8 126
rect 190 126 191 127
rect 189 126 190 127
rect 188 126 189 127
rect 180 126 181 127
rect 171 126 172 127
rect 170 126 171 127
rect 163 126 164 127
rect 111 126 112 127
rect 110 126 111 127
rect 109 126 110 127
rect 108 126 109 127
rect 107 126 108 127
rect 106 126 107 127
rect 105 126 106 127
rect 104 126 105 127
rect 103 126 104 127
rect 102 126 103 127
rect 101 126 102 127
rect 100 126 101 127
rect 99 126 100 127
rect 98 126 99 127
rect 97 126 98 127
rect 96 126 97 127
rect 95 126 96 127
rect 94 126 95 127
rect 93 126 94 127
rect 92 126 93 127
rect 91 126 92 127
rect 90 126 91 127
rect 89 126 90 127
rect 88 126 89 127
rect 76 126 77 127
rect 75 126 76 127
rect 74 126 75 127
rect 73 126 74 127
rect 72 126 73 127
rect 71 126 72 127
rect 70 126 71 127
rect 69 126 70 127
rect 68 126 69 127
rect 67 126 68 127
rect 66 126 67 127
rect 65 126 66 127
rect 64 126 65 127
rect 54 126 55 127
rect 53 126 54 127
rect 52 126 53 127
rect 51 126 52 127
rect 50 126 51 127
rect 49 126 50 127
rect 48 126 49 127
rect 47 126 48 127
rect 46 126 47 127
rect 45 126 46 127
rect 44 126 45 127
rect 43 126 44 127
rect 42 126 43 127
rect 41 126 42 127
rect 40 126 41 127
rect 39 126 40 127
rect 33 126 34 127
rect 32 126 33 127
rect 31 126 32 127
rect 30 126 31 127
rect 29 126 30 127
rect 28 126 29 127
rect 27 126 28 127
rect 26 126 27 127
rect 25 126 26 127
rect 24 126 25 127
rect 23 126 24 127
rect 22 126 23 127
rect 17 126 18 127
rect 16 126 17 127
rect 15 126 16 127
rect 14 126 15 127
rect 13 126 14 127
rect 12 126 13 127
rect 11 126 12 127
rect 10 126 11 127
rect 9 126 10 127
rect 8 126 9 127
rect 180 127 181 128
rect 171 127 172 128
rect 170 127 171 128
rect 163 127 164 128
rect 110 127 111 128
rect 109 127 110 128
rect 108 127 109 128
rect 107 127 108 128
rect 106 127 107 128
rect 105 127 106 128
rect 104 127 105 128
rect 103 127 104 128
rect 102 127 103 128
rect 101 127 102 128
rect 100 127 101 128
rect 99 127 100 128
rect 98 127 99 128
rect 97 127 98 128
rect 96 127 97 128
rect 95 127 96 128
rect 94 127 95 128
rect 93 127 94 128
rect 92 127 93 128
rect 91 127 92 128
rect 90 127 91 128
rect 89 127 90 128
rect 88 127 89 128
rect 87 127 88 128
rect 75 127 76 128
rect 74 127 75 128
rect 73 127 74 128
rect 72 127 73 128
rect 71 127 72 128
rect 70 127 71 128
rect 69 127 70 128
rect 68 127 69 128
rect 67 127 68 128
rect 66 127 67 128
rect 54 127 55 128
rect 53 127 54 128
rect 52 127 53 128
rect 51 127 52 128
rect 50 127 51 128
rect 49 127 50 128
rect 48 127 49 128
rect 47 127 48 128
rect 46 127 47 128
rect 45 127 46 128
rect 44 127 45 128
rect 43 127 44 128
rect 42 127 43 128
rect 41 127 42 128
rect 40 127 41 128
rect 33 127 34 128
rect 32 127 33 128
rect 31 127 32 128
rect 30 127 31 128
rect 29 127 30 128
rect 28 127 29 128
rect 27 127 28 128
rect 26 127 27 128
rect 25 127 26 128
rect 24 127 25 128
rect 23 127 24 128
rect 22 127 23 128
rect 17 127 18 128
rect 16 127 17 128
rect 15 127 16 128
rect 14 127 15 128
rect 13 127 14 128
rect 12 127 13 128
rect 11 127 12 128
rect 10 127 11 128
rect 9 127 10 128
rect 8 127 9 128
rect 180 128 181 129
rect 179 128 180 129
rect 172 128 173 129
rect 171 128 172 129
rect 170 128 171 129
rect 164 128 165 129
rect 163 128 164 129
rect 109 128 110 129
rect 108 128 109 129
rect 107 128 108 129
rect 106 128 107 129
rect 105 128 106 129
rect 104 128 105 129
rect 103 128 104 129
rect 102 128 103 129
rect 101 128 102 129
rect 100 128 101 129
rect 99 128 100 129
rect 98 128 99 129
rect 97 128 98 129
rect 96 128 97 129
rect 95 128 96 129
rect 94 128 95 129
rect 93 128 94 129
rect 92 128 93 129
rect 91 128 92 129
rect 90 128 91 129
rect 89 128 90 129
rect 88 128 89 129
rect 87 128 88 129
rect 86 128 87 129
rect 72 128 73 129
rect 71 128 72 129
rect 70 128 71 129
rect 69 128 70 129
rect 68 128 69 129
rect 55 128 56 129
rect 54 128 55 129
rect 53 128 54 129
rect 52 128 53 129
rect 51 128 52 129
rect 50 128 51 129
rect 49 128 50 129
rect 48 128 49 129
rect 47 128 48 129
rect 46 128 47 129
rect 45 128 46 129
rect 44 128 45 129
rect 43 128 44 129
rect 42 128 43 129
rect 41 128 42 129
rect 40 128 41 129
rect 34 128 35 129
rect 33 128 34 129
rect 32 128 33 129
rect 31 128 32 129
rect 30 128 31 129
rect 29 128 30 129
rect 28 128 29 129
rect 27 128 28 129
rect 26 128 27 129
rect 25 128 26 129
rect 24 128 25 129
rect 23 128 24 129
rect 22 128 23 129
rect 18 128 19 129
rect 17 128 18 129
rect 16 128 17 129
rect 15 128 16 129
rect 14 128 15 129
rect 13 128 14 129
rect 12 128 13 129
rect 11 128 12 129
rect 10 128 11 129
rect 9 128 10 129
rect 180 129 181 130
rect 179 129 180 130
rect 178 129 179 130
rect 177 129 178 130
rect 176 129 177 130
rect 175 129 176 130
rect 174 129 175 130
rect 173 129 174 130
rect 172 129 173 130
rect 171 129 172 130
rect 170 129 171 130
rect 169 129 170 130
rect 168 129 169 130
rect 167 129 168 130
rect 166 129 167 130
rect 165 129 166 130
rect 164 129 165 130
rect 163 129 164 130
rect 107 129 108 130
rect 106 129 107 130
rect 105 129 106 130
rect 104 129 105 130
rect 103 129 104 130
rect 102 129 103 130
rect 101 129 102 130
rect 100 129 101 130
rect 99 129 100 130
rect 98 129 99 130
rect 97 129 98 130
rect 96 129 97 130
rect 95 129 96 130
rect 94 129 95 130
rect 93 129 94 130
rect 92 129 93 130
rect 91 129 92 130
rect 90 129 91 130
rect 89 129 90 130
rect 88 129 89 130
rect 87 129 88 130
rect 86 129 87 130
rect 85 129 86 130
rect 56 129 57 130
rect 55 129 56 130
rect 54 129 55 130
rect 53 129 54 130
rect 52 129 53 130
rect 51 129 52 130
rect 50 129 51 130
rect 49 129 50 130
rect 48 129 49 130
rect 47 129 48 130
rect 46 129 47 130
rect 45 129 46 130
rect 44 129 45 130
rect 43 129 44 130
rect 42 129 43 130
rect 41 129 42 130
rect 34 129 35 130
rect 33 129 34 130
rect 32 129 33 130
rect 31 129 32 130
rect 30 129 31 130
rect 29 129 30 130
rect 28 129 29 130
rect 27 129 28 130
rect 26 129 27 130
rect 25 129 26 130
rect 24 129 25 130
rect 23 129 24 130
rect 18 129 19 130
rect 17 129 18 130
rect 16 129 17 130
rect 15 129 16 130
rect 14 129 15 130
rect 13 129 14 130
rect 12 129 13 130
rect 11 129 12 130
rect 10 129 11 130
rect 9 129 10 130
rect 180 130 181 131
rect 179 130 180 131
rect 178 130 179 131
rect 177 130 178 131
rect 176 130 177 131
rect 175 130 176 131
rect 174 130 175 131
rect 173 130 174 131
rect 172 130 173 131
rect 171 130 172 131
rect 170 130 171 131
rect 169 130 170 131
rect 168 130 169 131
rect 167 130 168 131
rect 166 130 167 131
rect 165 130 166 131
rect 164 130 165 131
rect 163 130 164 131
rect 105 130 106 131
rect 104 130 105 131
rect 103 130 104 131
rect 102 130 103 131
rect 101 130 102 131
rect 100 130 101 131
rect 99 130 100 131
rect 98 130 99 131
rect 97 130 98 131
rect 96 130 97 131
rect 95 130 96 131
rect 94 130 95 131
rect 93 130 94 131
rect 92 130 93 131
rect 91 130 92 131
rect 90 130 91 131
rect 89 130 90 131
rect 88 130 89 131
rect 87 130 88 131
rect 86 130 87 131
rect 85 130 86 131
rect 84 130 85 131
rect 57 130 58 131
rect 56 130 57 131
rect 55 130 56 131
rect 54 130 55 131
rect 53 130 54 131
rect 52 130 53 131
rect 51 130 52 131
rect 50 130 51 131
rect 49 130 50 131
rect 48 130 49 131
rect 47 130 48 131
rect 46 130 47 131
rect 45 130 46 131
rect 44 130 45 131
rect 43 130 44 131
rect 42 130 43 131
rect 41 130 42 131
rect 34 130 35 131
rect 33 130 34 131
rect 32 130 33 131
rect 31 130 32 131
rect 30 130 31 131
rect 29 130 30 131
rect 28 130 29 131
rect 27 130 28 131
rect 26 130 27 131
rect 25 130 26 131
rect 24 130 25 131
rect 23 130 24 131
rect 18 130 19 131
rect 17 130 18 131
rect 16 130 17 131
rect 15 130 16 131
rect 14 130 15 131
rect 13 130 14 131
rect 12 130 13 131
rect 11 130 12 131
rect 10 130 11 131
rect 189 131 190 132
rect 180 131 181 132
rect 179 131 180 132
rect 178 131 179 132
rect 177 131 178 132
rect 176 131 177 132
rect 175 131 176 132
rect 174 131 175 132
rect 173 131 174 132
rect 172 131 173 132
rect 171 131 172 132
rect 170 131 171 132
rect 169 131 170 132
rect 168 131 169 132
rect 167 131 168 132
rect 166 131 167 132
rect 165 131 166 132
rect 164 131 165 132
rect 163 131 164 132
rect 103 131 104 132
rect 102 131 103 132
rect 101 131 102 132
rect 100 131 101 132
rect 99 131 100 132
rect 98 131 99 132
rect 97 131 98 132
rect 96 131 97 132
rect 95 131 96 132
rect 94 131 95 132
rect 93 131 94 132
rect 92 131 93 132
rect 91 131 92 132
rect 90 131 91 132
rect 89 131 90 132
rect 88 131 89 132
rect 87 131 88 132
rect 86 131 87 132
rect 85 131 86 132
rect 84 131 85 132
rect 83 131 84 132
rect 58 131 59 132
rect 57 131 58 132
rect 56 131 57 132
rect 55 131 56 132
rect 54 131 55 132
rect 53 131 54 132
rect 52 131 53 132
rect 51 131 52 132
rect 50 131 51 132
rect 49 131 50 132
rect 48 131 49 132
rect 47 131 48 132
rect 46 131 47 132
rect 45 131 46 132
rect 44 131 45 132
rect 43 131 44 132
rect 42 131 43 132
rect 35 131 36 132
rect 34 131 35 132
rect 33 131 34 132
rect 32 131 33 132
rect 31 131 32 132
rect 30 131 31 132
rect 29 131 30 132
rect 28 131 29 132
rect 27 131 28 132
rect 26 131 27 132
rect 25 131 26 132
rect 24 131 25 132
rect 23 131 24 132
rect 18 131 19 132
rect 17 131 18 132
rect 16 131 17 132
rect 15 131 16 132
rect 14 131 15 132
rect 13 131 14 132
rect 12 131 13 132
rect 11 131 12 132
rect 10 131 11 132
rect 191 132 192 133
rect 190 132 191 133
rect 189 132 190 133
rect 180 132 181 133
rect 179 132 180 133
rect 178 132 179 133
rect 177 132 178 133
rect 176 132 177 133
rect 175 132 176 133
rect 174 132 175 133
rect 173 132 174 133
rect 172 132 173 133
rect 171 132 172 133
rect 170 132 171 133
rect 169 132 170 133
rect 168 132 169 133
rect 167 132 168 133
rect 166 132 167 133
rect 165 132 166 133
rect 164 132 165 133
rect 163 132 164 133
rect 101 132 102 133
rect 100 132 101 133
rect 99 132 100 133
rect 98 132 99 133
rect 97 132 98 133
rect 96 132 97 133
rect 95 132 96 133
rect 94 132 95 133
rect 93 132 94 133
rect 92 132 93 133
rect 91 132 92 133
rect 90 132 91 133
rect 89 132 90 133
rect 88 132 89 133
rect 87 132 88 133
rect 86 132 87 133
rect 85 132 86 133
rect 84 132 85 133
rect 83 132 84 133
rect 82 132 83 133
rect 59 132 60 133
rect 58 132 59 133
rect 57 132 58 133
rect 56 132 57 133
rect 55 132 56 133
rect 54 132 55 133
rect 53 132 54 133
rect 52 132 53 133
rect 51 132 52 133
rect 50 132 51 133
rect 49 132 50 133
rect 48 132 49 133
rect 47 132 48 133
rect 46 132 47 133
rect 45 132 46 133
rect 44 132 45 133
rect 43 132 44 133
rect 35 132 36 133
rect 34 132 35 133
rect 33 132 34 133
rect 32 132 33 133
rect 31 132 32 133
rect 30 132 31 133
rect 29 132 30 133
rect 28 132 29 133
rect 27 132 28 133
rect 26 132 27 133
rect 25 132 26 133
rect 24 132 25 133
rect 19 132 20 133
rect 18 132 19 133
rect 17 132 18 133
rect 16 132 17 133
rect 15 132 16 133
rect 14 132 15 133
rect 13 132 14 133
rect 12 132 13 133
rect 11 132 12 133
rect 197 133 198 134
rect 196 133 197 134
rect 195 133 196 134
rect 194 133 195 134
rect 193 133 194 134
rect 192 133 193 134
rect 191 133 192 134
rect 190 133 191 134
rect 189 133 190 134
rect 180 133 181 134
rect 179 133 180 134
rect 163 133 164 134
rect 98 133 99 134
rect 97 133 98 134
rect 96 133 97 134
rect 95 133 96 134
rect 94 133 95 134
rect 93 133 94 134
rect 92 133 93 134
rect 91 133 92 134
rect 90 133 91 134
rect 89 133 90 134
rect 88 133 89 134
rect 87 133 88 134
rect 86 133 87 134
rect 85 133 86 134
rect 84 133 85 134
rect 83 133 84 134
rect 82 133 83 134
rect 81 133 82 134
rect 61 133 62 134
rect 60 133 61 134
rect 59 133 60 134
rect 58 133 59 134
rect 57 133 58 134
rect 56 133 57 134
rect 55 133 56 134
rect 54 133 55 134
rect 53 133 54 134
rect 52 133 53 134
rect 51 133 52 134
rect 50 133 51 134
rect 49 133 50 134
rect 48 133 49 134
rect 47 133 48 134
rect 46 133 47 134
rect 45 133 46 134
rect 44 133 45 134
rect 43 133 44 134
rect 36 133 37 134
rect 35 133 36 134
rect 34 133 35 134
rect 33 133 34 134
rect 32 133 33 134
rect 31 133 32 134
rect 30 133 31 134
rect 29 133 30 134
rect 28 133 29 134
rect 27 133 28 134
rect 26 133 27 134
rect 25 133 26 134
rect 24 133 25 134
rect 19 133 20 134
rect 18 133 19 134
rect 17 133 18 134
rect 16 133 17 134
rect 15 133 16 134
rect 14 133 15 134
rect 13 133 14 134
rect 12 133 13 134
rect 196 134 197 135
rect 195 134 196 135
rect 194 134 195 135
rect 193 134 194 135
rect 192 134 193 135
rect 180 134 181 135
rect 163 134 164 135
rect 93 134 94 135
rect 92 134 93 135
rect 91 134 92 135
rect 90 134 91 135
rect 89 134 90 135
rect 88 134 89 135
rect 87 134 88 135
rect 86 134 87 135
rect 85 134 86 135
rect 83 134 84 135
rect 62 134 63 135
rect 61 134 62 135
rect 60 134 61 135
rect 59 134 60 135
rect 58 134 59 135
rect 57 134 58 135
rect 56 134 57 135
rect 55 134 56 135
rect 54 134 55 135
rect 53 134 54 135
rect 52 134 53 135
rect 51 134 52 135
rect 50 134 51 135
rect 49 134 50 135
rect 48 134 49 135
rect 47 134 48 135
rect 46 134 47 135
rect 45 134 46 135
rect 44 134 45 135
rect 36 134 37 135
rect 35 134 36 135
rect 34 134 35 135
rect 33 134 34 135
rect 32 134 33 135
rect 31 134 32 135
rect 30 134 31 135
rect 29 134 30 135
rect 28 134 29 135
rect 27 134 28 135
rect 26 134 27 135
rect 25 134 26 135
rect 24 134 25 135
rect 19 134 20 135
rect 18 134 19 135
rect 17 134 18 135
rect 16 134 17 135
rect 15 134 16 135
rect 14 134 15 135
rect 13 134 14 135
rect 196 135 197 136
rect 195 135 196 136
rect 194 135 195 136
rect 193 135 194 136
rect 192 135 193 136
rect 191 135 192 136
rect 64 135 65 136
rect 63 135 64 136
rect 62 135 63 136
rect 61 135 62 136
rect 60 135 61 136
rect 59 135 60 136
rect 58 135 59 136
rect 57 135 58 136
rect 56 135 57 136
rect 55 135 56 136
rect 54 135 55 136
rect 53 135 54 136
rect 52 135 53 136
rect 51 135 52 136
rect 50 135 51 136
rect 49 135 50 136
rect 48 135 49 136
rect 47 135 48 136
rect 46 135 47 136
rect 45 135 46 136
rect 37 135 38 136
rect 36 135 37 136
rect 35 135 36 136
rect 34 135 35 136
rect 33 135 34 136
rect 32 135 33 136
rect 31 135 32 136
rect 30 135 31 136
rect 29 135 30 136
rect 28 135 29 136
rect 27 135 28 136
rect 26 135 27 136
rect 25 135 26 136
rect 20 135 21 136
rect 19 135 20 136
rect 18 135 19 136
rect 17 135 18 136
rect 16 135 17 136
rect 15 135 16 136
rect 14 135 15 136
rect 13 135 14 136
rect 191 136 192 137
rect 190 136 191 137
rect 189 136 190 137
rect 66 136 67 137
rect 65 136 66 137
rect 64 136 65 137
rect 63 136 64 137
rect 62 136 63 137
rect 61 136 62 137
rect 60 136 61 137
rect 59 136 60 137
rect 58 136 59 137
rect 57 136 58 137
rect 56 136 57 137
rect 55 136 56 137
rect 54 136 55 137
rect 53 136 54 137
rect 52 136 53 137
rect 51 136 52 137
rect 50 136 51 137
rect 49 136 50 137
rect 48 136 49 137
rect 47 136 48 137
rect 46 136 47 137
rect 38 136 39 137
rect 37 136 38 137
rect 36 136 37 137
rect 35 136 36 137
rect 34 136 35 137
rect 33 136 34 137
rect 32 136 33 137
rect 31 136 32 137
rect 30 136 31 137
rect 29 136 30 137
rect 28 136 29 137
rect 27 136 28 137
rect 26 136 27 137
rect 25 136 26 137
rect 20 136 21 137
rect 19 136 20 137
rect 18 136 19 137
rect 17 136 18 137
rect 16 136 17 137
rect 15 136 16 137
rect 14 136 15 137
rect 189 137 190 138
rect 69 137 70 138
rect 68 137 69 138
rect 67 137 68 138
rect 66 137 67 138
rect 65 137 66 138
rect 64 137 65 138
rect 63 137 64 138
rect 62 137 63 138
rect 61 137 62 138
rect 60 137 61 138
rect 59 137 60 138
rect 58 137 59 138
rect 57 137 58 138
rect 56 137 57 138
rect 55 137 56 138
rect 54 137 55 138
rect 53 137 54 138
rect 52 137 53 138
rect 51 137 52 138
rect 50 137 51 138
rect 49 137 50 138
rect 48 137 49 138
rect 47 137 48 138
rect 38 137 39 138
rect 37 137 38 138
rect 36 137 37 138
rect 35 137 36 138
rect 34 137 35 138
rect 33 137 34 138
rect 32 137 33 138
rect 31 137 32 138
rect 30 137 31 138
rect 29 137 30 138
rect 28 137 29 138
rect 27 137 28 138
rect 26 137 27 138
rect 25 137 26 138
rect 20 137 21 138
rect 19 137 20 138
rect 18 137 19 138
rect 17 137 18 138
rect 16 137 17 138
rect 15 137 16 138
rect 180 138 181 139
rect 163 138 164 139
rect 72 138 73 139
rect 71 138 72 139
rect 70 138 71 139
rect 69 138 70 139
rect 68 138 69 139
rect 67 138 68 139
rect 66 138 67 139
rect 65 138 66 139
rect 64 138 65 139
rect 63 138 64 139
rect 62 138 63 139
rect 61 138 62 139
rect 60 138 61 139
rect 59 138 60 139
rect 58 138 59 139
rect 57 138 58 139
rect 56 138 57 139
rect 55 138 56 139
rect 54 138 55 139
rect 53 138 54 139
rect 52 138 53 139
rect 51 138 52 139
rect 50 138 51 139
rect 49 138 50 139
rect 48 138 49 139
rect 47 138 48 139
rect 39 138 40 139
rect 38 138 39 139
rect 37 138 38 139
rect 36 138 37 139
rect 35 138 36 139
rect 34 138 35 139
rect 33 138 34 139
rect 32 138 33 139
rect 31 138 32 139
rect 30 138 31 139
rect 29 138 30 139
rect 28 138 29 139
rect 27 138 28 139
rect 26 138 27 139
rect 21 138 22 139
rect 20 138 21 139
rect 19 138 20 139
rect 18 138 19 139
rect 17 138 18 139
rect 16 138 17 139
rect 180 139 181 140
rect 163 139 164 140
rect 76 139 77 140
rect 75 139 76 140
rect 74 139 75 140
rect 73 139 74 140
rect 72 139 73 140
rect 71 139 72 140
rect 70 139 71 140
rect 69 139 70 140
rect 68 139 69 140
rect 67 139 68 140
rect 66 139 67 140
rect 65 139 66 140
rect 64 139 65 140
rect 63 139 64 140
rect 62 139 63 140
rect 61 139 62 140
rect 60 139 61 140
rect 59 139 60 140
rect 58 139 59 140
rect 57 139 58 140
rect 56 139 57 140
rect 55 139 56 140
rect 54 139 55 140
rect 53 139 54 140
rect 52 139 53 140
rect 51 139 52 140
rect 50 139 51 140
rect 49 139 50 140
rect 48 139 49 140
rect 40 139 41 140
rect 39 139 40 140
rect 38 139 39 140
rect 37 139 38 140
rect 36 139 37 140
rect 35 139 36 140
rect 34 139 35 140
rect 33 139 34 140
rect 32 139 33 140
rect 31 139 32 140
rect 30 139 31 140
rect 29 139 30 140
rect 28 139 29 140
rect 27 139 28 140
rect 26 139 27 140
rect 21 139 22 140
rect 20 139 21 140
rect 19 139 20 140
rect 18 139 19 140
rect 17 139 18 140
rect 180 140 181 141
rect 179 140 180 141
rect 178 140 179 141
rect 177 140 178 141
rect 176 140 177 141
rect 175 140 176 141
rect 174 140 175 141
rect 173 140 174 141
rect 172 140 173 141
rect 171 140 172 141
rect 170 140 171 141
rect 169 140 170 141
rect 168 140 169 141
rect 167 140 168 141
rect 166 140 167 141
rect 165 140 166 141
rect 164 140 165 141
rect 163 140 164 141
rect 75 140 76 141
rect 74 140 75 141
rect 73 140 74 141
rect 72 140 73 141
rect 71 140 72 141
rect 70 140 71 141
rect 69 140 70 141
rect 68 140 69 141
rect 67 140 68 141
rect 66 140 67 141
rect 65 140 66 141
rect 64 140 65 141
rect 63 140 64 141
rect 62 140 63 141
rect 61 140 62 141
rect 60 140 61 141
rect 59 140 60 141
rect 58 140 59 141
rect 57 140 58 141
rect 56 140 57 141
rect 55 140 56 141
rect 54 140 55 141
rect 53 140 54 141
rect 52 140 53 141
rect 51 140 52 141
rect 50 140 51 141
rect 49 140 50 141
rect 41 140 42 141
rect 40 140 41 141
rect 39 140 40 141
rect 38 140 39 141
rect 37 140 38 141
rect 36 140 37 141
rect 35 140 36 141
rect 34 140 35 141
rect 33 140 34 141
rect 32 140 33 141
rect 31 140 32 141
rect 30 140 31 141
rect 29 140 30 141
rect 28 140 29 141
rect 27 140 28 141
rect 22 140 23 141
rect 21 140 22 141
rect 20 140 21 141
rect 19 140 20 141
rect 18 140 19 141
rect 180 141 181 142
rect 179 141 180 142
rect 178 141 179 142
rect 177 141 178 142
rect 176 141 177 142
rect 175 141 176 142
rect 174 141 175 142
rect 173 141 174 142
rect 172 141 173 142
rect 171 141 172 142
rect 170 141 171 142
rect 169 141 170 142
rect 168 141 169 142
rect 167 141 168 142
rect 166 141 167 142
rect 165 141 166 142
rect 164 141 165 142
rect 163 141 164 142
rect 74 141 75 142
rect 73 141 74 142
rect 72 141 73 142
rect 71 141 72 142
rect 70 141 71 142
rect 69 141 70 142
rect 68 141 69 142
rect 67 141 68 142
rect 66 141 67 142
rect 65 141 66 142
rect 64 141 65 142
rect 63 141 64 142
rect 62 141 63 142
rect 61 141 62 142
rect 60 141 61 142
rect 59 141 60 142
rect 58 141 59 142
rect 57 141 58 142
rect 56 141 57 142
rect 55 141 56 142
rect 54 141 55 142
rect 53 141 54 142
rect 52 141 53 142
rect 51 141 52 142
rect 50 141 51 142
rect 41 141 42 142
rect 40 141 41 142
rect 39 141 40 142
rect 38 141 39 142
rect 37 141 38 142
rect 36 141 37 142
rect 35 141 36 142
rect 34 141 35 142
rect 33 141 34 142
rect 32 141 33 142
rect 31 141 32 142
rect 30 141 31 142
rect 29 141 30 142
rect 28 141 29 142
rect 27 141 28 142
rect 22 141 23 142
rect 21 141 22 142
rect 20 141 21 142
rect 19 141 20 142
rect 180 142 181 143
rect 179 142 180 143
rect 178 142 179 143
rect 177 142 178 143
rect 176 142 177 143
rect 175 142 176 143
rect 174 142 175 143
rect 173 142 174 143
rect 172 142 173 143
rect 171 142 172 143
rect 170 142 171 143
rect 169 142 170 143
rect 168 142 169 143
rect 167 142 168 143
rect 166 142 167 143
rect 165 142 166 143
rect 164 142 165 143
rect 163 142 164 143
rect 72 142 73 143
rect 71 142 72 143
rect 70 142 71 143
rect 69 142 70 143
rect 68 142 69 143
rect 67 142 68 143
rect 66 142 67 143
rect 65 142 66 143
rect 64 142 65 143
rect 63 142 64 143
rect 62 142 63 143
rect 61 142 62 143
rect 60 142 61 143
rect 59 142 60 143
rect 58 142 59 143
rect 57 142 58 143
rect 56 142 57 143
rect 55 142 56 143
rect 54 142 55 143
rect 53 142 54 143
rect 52 142 53 143
rect 51 142 52 143
rect 42 142 43 143
rect 41 142 42 143
rect 40 142 41 143
rect 39 142 40 143
rect 38 142 39 143
rect 37 142 38 143
rect 36 142 37 143
rect 35 142 36 143
rect 34 142 35 143
rect 33 142 34 143
rect 32 142 33 143
rect 31 142 32 143
rect 30 142 31 143
rect 29 142 30 143
rect 28 142 29 143
rect 27 142 28 143
rect 23 142 24 143
rect 22 142 23 143
rect 21 142 22 143
rect 20 142 21 143
rect 180 143 181 144
rect 179 143 180 144
rect 178 143 179 144
rect 177 143 178 144
rect 176 143 177 144
rect 175 143 176 144
rect 174 143 175 144
rect 173 143 174 144
rect 172 143 173 144
rect 171 143 172 144
rect 170 143 171 144
rect 169 143 170 144
rect 168 143 169 144
rect 167 143 168 144
rect 166 143 167 144
rect 165 143 166 144
rect 164 143 165 144
rect 163 143 164 144
rect 70 143 71 144
rect 69 143 70 144
rect 68 143 69 144
rect 67 143 68 144
rect 66 143 67 144
rect 65 143 66 144
rect 64 143 65 144
rect 63 143 64 144
rect 62 143 63 144
rect 61 143 62 144
rect 60 143 61 144
rect 59 143 60 144
rect 58 143 59 144
rect 57 143 58 144
rect 56 143 57 144
rect 55 143 56 144
rect 54 143 55 144
rect 53 143 54 144
rect 43 143 44 144
rect 42 143 43 144
rect 41 143 42 144
rect 40 143 41 144
rect 39 143 40 144
rect 38 143 39 144
rect 37 143 38 144
rect 36 143 37 144
rect 35 143 36 144
rect 34 143 35 144
rect 33 143 34 144
rect 32 143 33 144
rect 31 143 32 144
rect 30 143 31 144
rect 29 143 30 144
rect 28 143 29 144
rect 23 143 24 144
rect 180 144 181 145
rect 179 144 180 145
rect 172 144 173 145
rect 171 144 172 145
rect 170 144 171 145
rect 164 144 165 145
rect 163 144 164 145
rect 65 144 66 145
rect 64 144 65 145
rect 63 144 64 145
rect 62 144 63 145
rect 61 144 62 145
rect 60 144 61 145
rect 59 144 60 145
rect 58 144 59 145
rect 57 144 58 145
rect 56 144 57 145
rect 44 144 45 145
rect 43 144 44 145
rect 42 144 43 145
rect 41 144 42 145
rect 40 144 41 145
rect 39 144 40 145
rect 38 144 39 145
rect 37 144 38 145
rect 36 144 37 145
rect 35 144 36 145
rect 34 144 35 145
rect 33 144 34 145
rect 32 144 33 145
rect 31 144 32 145
rect 30 144 31 145
rect 29 144 30 145
rect 28 144 29 145
rect 180 145 181 146
rect 172 145 173 146
rect 171 145 172 146
rect 163 145 164 146
rect 45 145 46 146
rect 44 145 45 146
rect 43 145 44 146
rect 42 145 43 146
rect 41 145 42 146
rect 40 145 41 146
rect 39 145 40 146
rect 38 145 39 146
rect 37 145 38 146
rect 36 145 37 146
rect 35 145 36 146
rect 34 145 35 146
rect 33 145 34 146
rect 32 145 33 146
rect 31 145 32 146
rect 30 145 31 146
rect 29 145 30 146
rect 180 146 181 147
rect 172 146 173 147
rect 171 146 172 147
rect 163 146 164 147
rect 47 146 48 147
rect 46 146 47 147
rect 45 146 46 147
rect 44 146 45 147
rect 43 146 44 147
rect 42 146 43 147
rect 41 146 42 147
rect 40 146 41 147
rect 39 146 40 147
rect 38 146 39 147
rect 37 146 38 147
rect 36 146 37 147
rect 35 146 36 147
rect 34 146 35 147
rect 33 146 34 147
rect 32 146 33 147
rect 31 146 32 147
rect 30 146 31 147
rect 180 147 181 148
rect 172 147 173 148
rect 171 147 172 148
rect 163 147 164 148
rect 48 147 49 148
rect 47 147 48 148
rect 46 147 47 148
rect 45 147 46 148
rect 44 147 45 148
rect 43 147 44 148
rect 42 147 43 148
rect 41 147 42 148
rect 40 147 41 148
rect 39 147 40 148
rect 38 147 39 148
rect 37 147 38 148
rect 36 147 37 148
rect 35 147 36 148
rect 34 147 35 148
rect 33 147 34 148
rect 32 147 33 148
rect 31 147 32 148
rect 180 148 181 149
rect 173 148 174 149
rect 172 148 173 149
rect 171 148 172 149
rect 170 148 171 149
rect 164 148 165 149
rect 163 148 164 149
rect 50 148 51 149
rect 49 148 50 149
rect 48 148 49 149
rect 47 148 48 149
rect 46 148 47 149
rect 45 148 46 149
rect 44 148 45 149
rect 43 148 44 149
rect 42 148 43 149
rect 41 148 42 149
rect 40 148 41 149
rect 39 148 40 149
rect 38 148 39 149
rect 37 148 38 149
rect 36 148 37 149
rect 35 148 36 149
rect 34 148 35 149
rect 33 148 34 149
rect 32 148 33 149
rect 180 149 181 150
rect 179 149 180 150
rect 174 149 175 150
rect 173 149 174 150
rect 172 149 173 150
rect 171 149 172 150
rect 170 149 171 150
rect 169 149 170 150
rect 164 149 165 150
rect 163 149 164 150
rect 51 149 52 150
rect 50 149 51 150
rect 49 149 50 150
rect 48 149 49 150
rect 47 149 48 150
rect 46 149 47 150
rect 45 149 46 150
rect 44 149 45 150
rect 43 149 44 150
rect 42 149 43 150
rect 41 149 42 150
rect 40 149 41 150
rect 39 149 40 150
rect 38 149 39 150
rect 37 149 38 150
rect 36 149 37 150
rect 35 149 36 150
rect 34 149 35 150
rect 180 150 181 151
rect 179 150 180 151
rect 178 150 179 151
rect 167 150 168 151
rect 166 150 167 151
rect 165 150 166 151
rect 164 150 165 151
rect 163 150 164 151
rect 51 150 52 151
rect 50 150 51 151
rect 49 150 50 151
rect 48 150 49 151
rect 47 150 48 151
rect 46 150 47 151
rect 45 150 46 151
rect 44 150 45 151
rect 43 150 44 151
rect 42 150 43 151
rect 41 150 42 151
rect 40 150 41 151
rect 39 150 40 151
rect 38 150 39 151
rect 37 150 38 151
rect 180 151 181 152
rect 179 151 180 152
rect 178 151 179 152
rect 177 151 178 152
rect 176 151 177 152
rect 166 151 167 152
rect 165 151 166 152
rect 164 151 165 152
rect 47 151 48 152
rect 46 151 47 152
rect 45 151 46 152
rect 44 151 45 152
rect 43 151 44 152
rect 42 151 43 152
rect 178 152 179 153
rect 177 152 178 153
rect 176 152 177 153
rect 180 155 181 156
rect 163 155 164 156
rect 180 156 181 157
rect 163 156 164 157
rect 180 157 181 158
rect 179 157 180 158
rect 178 157 179 158
rect 177 157 178 158
rect 176 157 177 158
rect 175 157 176 158
rect 174 157 175 158
rect 173 157 174 158
rect 172 157 173 158
rect 171 157 172 158
rect 170 157 171 158
rect 169 157 170 158
rect 168 157 169 158
rect 167 157 168 158
rect 166 157 167 158
rect 165 157 166 158
rect 164 157 165 158
rect 163 157 164 158
rect 180 158 181 159
rect 179 158 180 159
rect 178 158 179 159
rect 177 158 178 159
rect 176 158 177 159
rect 175 158 176 159
rect 174 158 175 159
rect 173 158 174 159
rect 172 158 173 159
rect 171 158 172 159
rect 170 158 171 159
rect 169 158 170 159
rect 168 158 169 159
rect 167 158 168 159
rect 166 158 167 159
rect 165 158 166 159
rect 164 158 165 159
rect 163 158 164 159
rect 180 159 181 160
rect 179 159 180 160
rect 178 159 179 160
rect 177 159 178 160
rect 176 159 177 160
rect 175 159 176 160
rect 174 159 175 160
rect 173 159 174 160
rect 172 159 173 160
rect 171 159 172 160
rect 170 159 171 160
rect 169 159 170 160
rect 168 159 169 160
rect 167 159 168 160
rect 166 159 167 160
rect 165 159 166 160
rect 164 159 165 160
rect 163 159 164 160
rect 180 160 181 161
rect 179 160 180 161
rect 178 160 179 161
rect 177 160 178 161
rect 176 160 177 161
rect 175 160 176 161
rect 174 160 175 161
rect 173 160 174 161
rect 172 160 173 161
rect 171 160 172 161
rect 170 160 171 161
rect 169 160 170 161
rect 168 160 169 161
rect 167 160 168 161
rect 166 160 167 161
rect 165 160 166 161
rect 164 160 165 161
rect 163 160 164 161
rect 180 161 181 162
rect 179 161 180 162
rect 178 161 179 162
rect 177 161 178 162
rect 176 161 177 162
rect 175 161 176 162
rect 174 161 175 162
rect 173 161 174 162
rect 172 161 173 162
rect 171 161 172 162
rect 170 161 171 162
rect 169 161 170 162
rect 168 161 169 162
rect 167 161 168 162
rect 166 161 167 162
rect 165 161 166 162
rect 164 161 165 162
rect 163 161 164 162
rect 180 162 181 163
rect 179 162 180 163
rect 172 162 173 163
rect 171 162 172 163
rect 163 162 164 163
rect 180 163 181 164
rect 172 163 173 164
rect 171 163 172 164
rect 163 163 164 164
rect 180 164 181 165
rect 172 164 173 165
rect 171 164 172 165
rect 163 164 164 165
rect 180 165 181 166
rect 172 165 173 166
rect 171 165 172 166
rect 170 165 171 166
rect 164 165 165 166
rect 163 165 164 166
rect 180 166 181 167
rect 179 166 180 167
rect 174 166 175 167
rect 173 166 174 167
rect 172 166 173 167
rect 171 166 172 167
rect 170 166 171 167
rect 169 166 170 167
rect 164 166 165 167
rect 163 166 164 167
rect 180 167 181 168
rect 179 167 180 168
rect 178 167 179 168
rect 173 167 174 168
rect 172 167 173 168
rect 171 167 172 168
rect 170 167 171 168
rect 169 167 170 168
rect 166 167 167 168
rect 165 167 166 168
rect 164 167 165 168
rect 163 167 164 168
rect 180 168 181 169
rect 179 168 180 169
rect 178 168 179 169
rect 177 168 178 169
rect 166 168 167 169
rect 165 168 166 169
rect 164 168 165 169
rect 163 168 164 169
rect 179 169 180 170
rect 178 169 179 170
rect 177 169 178 170
rect 176 169 177 170
rect 143 176 144 177
rect 142 176 143 177
rect 141 176 142 177
rect 140 176 141 177
rect 139 176 140 177
rect 138 176 139 177
rect 137 176 138 177
rect 136 176 137 177
rect 135 176 136 177
rect 134 176 135 177
rect 133 176 134 177
rect 132 176 133 177
rect 131 176 132 177
rect 130 176 131 177
rect 129 176 130 177
rect 128 176 129 177
rect 127 176 128 177
rect 126 176 127 177
rect 125 176 126 177
rect 124 176 125 177
rect 123 176 124 177
rect 122 176 123 177
rect 121 176 122 177
rect 120 176 121 177
rect 119 176 120 177
rect 118 176 119 177
rect 117 176 118 177
rect 116 176 117 177
rect 115 176 116 177
rect 114 176 115 177
rect 113 176 114 177
rect 112 176 113 177
rect 111 176 112 177
rect 110 176 111 177
rect 109 176 110 177
rect 108 176 109 177
rect 107 176 108 177
rect 106 176 107 177
rect 105 176 106 177
rect 104 176 105 177
rect 103 176 104 177
rect 102 176 103 177
rect 145 177 146 178
rect 144 177 145 178
rect 143 177 144 178
rect 142 177 143 178
rect 141 177 142 178
rect 140 177 141 178
rect 139 177 140 178
rect 138 177 139 178
rect 137 177 138 178
rect 136 177 137 178
rect 135 177 136 178
rect 134 177 135 178
rect 133 177 134 178
rect 132 177 133 178
rect 131 177 132 178
rect 130 177 131 178
rect 129 177 130 178
rect 128 177 129 178
rect 127 177 128 178
rect 126 177 127 178
rect 125 177 126 178
rect 124 177 125 178
rect 123 177 124 178
rect 122 177 123 178
rect 121 177 122 178
rect 120 177 121 178
rect 119 177 120 178
rect 118 177 119 178
rect 117 177 118 178
rect 116 177 117 178
rect 115 177 116 178
rect 114 177 115 178
rect 113 177 114 178
rect 112 177 113 178
rect 111 177 112 178
rect 110 177 111 178
rect 109 177 110 178
rect 108 177 109 178
rect 107 177 108 178
rect 106 177 107 178
rect 105 177 106 178
rect 104 177 105 178
rect 103 177 104 178
rect 102 177 103 178
rect 196 178 197 179
rect 195 178 196 179
rect 194 178 195 179
rect 193 178 194 179
rect 192 178 193 179
rect 191 178 192 179
rect 190 178 191 179
rect 189 178 190 179
rect 172 178 173 179
rect 167 178 168 179
rect 166 178 167 179
rect 165 178 166 179
rect 146 178 147 179
rect 145 178 146 179
rect 144 178 145 179
rect 143 178 144 179
rect 142 178 143 179
rect 141 178 142 179
rect 140 178 141 179
rect 139 178 140 179
rect 138 178 139 179
rect 137 178 138 179
rect 136 178 137 179
rect 135 178 136 179
rect 134 178 135 179
rect 133 178 134 179
rect 132 178 133 179
rect 131 178 132 179
rect 130 178 131 179
rect 129 178 130 179
rect 128 178 129 179
rect 127 178 128 179
rect 126 178 127 179
rect 125 178 126 179
rect 124 178 125 179
rect 123 178 124 179
rect 122 178 123 179
rect 121 178 122 179
rect 120 178 121 179
rect 119 178 120 179
rect 118 178 119 179
rect 117 178 118 179
rect 116 178 117 179
rect 115 178 116 179
rect 114 178 115 179
rect 113 178 114 179
rect 112 178 113 179
rect 111 178 112 179
rect 110 178 111 179
rect 109 178 110 179
rect 108 178 109 179
rect 107 178 108 179
rect 106 178 107 179
rect 105 178 106 179
rect 104 178 105 179
rect 103 178 104 179
rect 102 178 103 179
rect 197 179 198 180
rect 196 179 197 180
rect 195 179 196 180
rect 194 179 195 180
rect 193 179 194 180
rect 192 179 193 180
rect 191 179 192 180
rect 190 179 191 180
rect 189 179 190 180
rect 174 179 175 180
rect 173 179 174 180
rect 172 179 173 180
rect 171 179 172 180
rect 170 179 171 180
rect 167 179 168 180
rect 166 179 167 180
rect 165 179 166 180
rect 147 179 148 180
rect 146 179 147 180
rect 145 179 146 180
rect 144 179 145 180
rect 143 179 144 180
rect 142 179 143 180
rect 141 179 142 180
rect 140 179 141 180
rect 139 179 140 180
rect 138 179 139 180
rect 137 179 138 180
rect 136 179 137 180
rect 135 179 136 180
rect 134 179 135 180
rect 133 179 134 180
rect 132 179 133 180
rect 131 179 132 180
rect 130 179 131 180
rect 129 179 130 180
rect 128 179 129 180
rect 127 179 128 180
rect 126 179 127 180
rect 125 179 126 180
rect 124 179 125 180
rect 123 179 124 180
rect 122 179 123 180
rect 121 179 122 180
rect 120 179 121 180
rect 119 179 120 180
rect 118 179 119 180
rect 117 179 118 180
rect 116 179 117 180
rect 115 179 116 180
rect 114 179 115 180
rect 113 179 114 180
rect 112 179 113 180
rect 111 179 112 180
rect 110 179 111 180
rect 109 179 110 180
rect 108 179 109 180
rect 107 179 108 180
rect 106 179 107 180
rect 105 179 106 180
rect 104 179 105 180
rect 103 179 104 180
rect 102 179 103 180
rect 196 180 197 181
rect 195 180 196 181
rect 194 180 195 181
rect 193 180 194 181
rect 192 180 193 181
rect 191 180 192 181
rect 190 180 191 181
rect 189 180 190 181
rect 174 180 175 181
rect 173 180 174 181
rect 172 180 173 181
rect 171 180 172 181
rect 170 180 171 181
rect 169 180 170 181
rect 167 180 168 181
rect 166 180 167 181
rect 165 180 166 181
rect 148 180 149 181
rect 147 180 148 181
rect 146 180 147 181
rect 145 180 146 181
rect 144 180 145 181
rect 143 180 144 181
rect 142 180 143 181
rect 141 180 142 181
rect 140 180 141 181
rect 139 180 140 181
rect 138 180 139 181
rect 137 180 138 181
rect 136 180 137 181
rect 135 180 136 181
rect 134 180 135 181
rect 133 180 134 181
rect 132 180 133 181
rect 131 180 132 181
rect 130 180 131 181
rect 129 180 130 181
rect 128 180 129 181
rect 127 180 128 181
rect 126 180 127 181
rect 125 180 126 181
rect 124 180 125 181
rect 123 180 124 181
rect 122 180 123 181
rect 121 180 122 181
rect 120 180 121 181
rect 119 180 120 181
rect 118 180 119 181
rect 117 180 118 181
rect 116 180 117 181
rect 115 180 116 181
rect 114 180 115 181
rect 113 180 114 181
rect 112 180 113 181
rect 111 180 112 181
rect 110 180 111 181
rect 109 180 110 181
rect 108 180 109 181
rect 107 180 108 181
rect 106 180 107 181
rect 105 180 106 181
rect 104 180 105 181
rect 103 180 104 181
rect 102 180 103 181
rect 196 181 197 182
rect 193 181 194 182
rect 192 181 193 182
rect 189 181 190 182
rect 182 181 183 182
rect 181 181 182 182
rect 180 181 181 182
rect 179 181 180 182
rect 178 181 179 182
rect 175 181 176 182
rect 174 181 175 182
rect 173 181 174 182
rect 172 181 173 182
rect 171 181 172 182
rect 170 181 171 182
rect 169 181 170 182
rect 167 181 168 182
rect 166 181 167 182
rect 165 181 166 182
rect 163 181 164 182
rect 162 181 163 182
rect 148 181 149 182
rect 147 181 148 182
rect 146 181 147 182
rect 145 181 146 182
rect 144 181 145 182
rect 143 181 144 182
rect 142 181 143 182
rect 141 181 142 182
rect 140 181 141 182
rect 139 181 140 182
rect 138 181 139 182
rect 137 181 138 182
rect 136 181 137 182
rect 135 181 136 182
rect 134 181 135 182
rect 133 181 134 182
rect 132 181 133 182
rect 131 181 132 182
rect 130 181 131 182
rect 129 181 130 182
rect 128 181 129 182
rect 127 181 128 182
rect 126 181 127 182
rect 125 181 126 182
rect 124 181 125 182
rect 123 181 124 182
rect 122 181 123 182
rect 121 181 122 182
rect 120 181 121 182
rect 119 181 120 182
rect 118 181 119 182
rect 117 181 118 182
rect 116 181 117 182
rect 115 181 116 182
rect 114 181 115 182
rect 113 181 114 182
rect 112 181 113 182
rect 111 181 112 182
rect 110 181 111 182
rect 109 181 110 182
rect 108 181 109 182
rect 107 181 108 182
rect 106 181 107 182
rect 105 181 106 182
rect 104 181 105 182
rect 103 181 104 182
rect 102 181 103 182
rect 196 182 197 183
rect 193 182 194 183
rect 192 182 193 183
rect 189 182 190 183
rect 183 182 184 183
rect 182 182 183 183
rect 181 182 182 183
rect 180 182 181 183
rect 179 182 180 183
rect 178 182 179 183
rect 177 182 178 183
rect 175 182 176 183
rect 174 182 175 183
rect 173 182 174 183
rect 172 182 173 183
rect 171 182 172 183
rect 170 182 171 183
rect 169 182 170 183
rect 167 182 168 183
rect 166 182 167 183
rect 165 182 166 183
rect 163 182 164 183
rect 162 182 163 183
rect 149 182 150 183
rect 148 182 149 183
rect 147 182 148 183
rect 146 182 147 183
rect 145 182 146 183
rect 144 182 145 183
rect 143 182 144 183
rect 142 182 143 183
rect 141 182 142 183
rect 140 182 141 183
rect 139 182 140 183
rect 138 182 139 183
rect 137 182 138 183
rect 136 182 137 183
rect 135 182 136 183
rect 134 182 135 183
rect 133 182 134 183
rect 132 182 133 183
rect 131 182 132 183
rect 130 182 131 183
rect 129 182 130 183
rect 128 182 129 183
rect 127 182 128 183
rect 126 182 127 183
rect 125 182 126 183
rect 124 182 125 183
rect 123 182 124 183
rect 122 182 123 183
rect 121 182 122 183
rect 120 182 121 183
rect 119 182 120 183
rect 118 182 119 183
rect 117 182 118 183
rect 116 182 117 183
rect 115 182 116 183
rect 114 182 115 183
rect 113 182 114 183
rect 112 182 113 183
rect 111 182 112 183
rect 110 182 111 183
rect 109 182 110 183
rect 108 182 109 183
rect 107 182 108 183
rect 106 182 107 183
rect 105 182 106 183
rect 104 182 105 183
rect 103 182 104 183
rect 102 182 103 183
rect 62 182 63 183
rect 61 182 62 183
rect 60 182 61 183
rect 59 182 60 183
rect 197 183 198 184
rect 196 183 197 184
rect 193 183 194 184
rect 192 183 193 184
rect 189 183 190 184
rect 183 183 184 184
rect 182 183 183 184
rect 181 183 182 184
rect 180 183 181 184
rect 179 183 180 184
rect 178 183 179 184
rect 177 183 178 184
rect 175 183 176 184
rect 174 183 175 184
rect 173 183 174 184
rect 171 183 172 184
rect 170 183 171 184
rect 169 183 170 184
rect 168 183 169 184
rect 167 183 168 184
rect 166 183 167 184
rect 165 183 166 184
rect 163 183 164 184
rect 162 183 163 184
rect 149 183 150 184
rect 148 183 149 184
rect 147 183 148 184
rect 146 183 147 184
rect 145 183 146 184
rect 144 183 145 184
rect 143 183 144 184
rect 142 183 143 184
rect 141 183 142 184
rect 140 183 141 184
rect 139 183 140 184
rect 138 183 139 184
rect 137 183 138 184
rect 136 183 137 184
rect 135 183 136 184
rect 134 183 135 184
rect 133 183 134 184
rect 132 183 133 184
rect 131 183 132 184
rect 130 183 131 184
rect 129 183 130 184
rect 128 183 129 184
rect 127 183 128 184
rect 126 183 127 184
rect 125 183 126 184
rect 124 183 125 184
rect 123 183 124 184
rect 122 183 123 184
rect 121 183 122 184
rect 120 183 121 184
rect 119 183 120 184
rect 118 183 119 184
rect 117 183 118 184
rect 116 183 117 184
rect 115 183 116 184
rect 114 183 115 184
rect 113 183 114 184
rect 112 183 113 184
rect 111 183 112 184
rect 110 183 111 184
rect 109 183 110 184
rect 108 183 109 184
rect 107 183 108 184
rect 106 183 107 184
rect 105 183 106 184
rect 104 183 105 184
rect 103 183 104 184
rect 102 183 103 184
rect 62 183 63 184
rect 61 183 62 184
rect 60 183 61 184
rect 59 183 60 184
rect 29 183 30 184
rect 28 183 29 184
rect 183 184 184 185
rect 182 184 183 185
rect 181 184 182 185
rect 180 184 181 185
rect 179 184 180 185
rect 178 184 179 185
rect 177 184 178 185
rect 175 184 176 185
rect 174 184 175 185
rect 170 184 171 185
rect 169 184 170 185
rect 168 184 169 185
rect 167 184 168 185
rect 166 184 167 185
rect 165 184 166 185
rect 163 184 164 185
rect 162 184 163 185
rect 149 184 150 185
rect 148 184 149 185
rect 147 184 148 185
rect 146 184 147 185
rect 145 184 146 185
rect 144 184 145 185
rect 143 184 144 185
rect 142 184 143 185
rect 141 184 142 185
rect 140 184 141 185
rect 139 184 140 185
rect 138 184 139 185
rect 137 184 138 185
rect 136 184 137 185
rect 135 184 136 185
rect 134 184 135 185
rect 133 184 134 185
rect 132 184 133 185
rect 131 184 132 185
rect 130 184 131 185
rect 129 184 130 185
rect 128 184 129 185
rect 127 184 128 185
rect 126 184 127 185
rect 125 184 126 185
rect 124 184 125 185
rect 123 184 124 185
rect 122 184 123 185
rect 121 184 122 185
rect 120 184 121 185
rect 119 184 120 185
rect 118 184 119 185
rect 117 184 118 185
rect 116 184 117 185
rect 115 184 116 185
rect 114 184 115 185
rect 113 184 114 185
rect 112 184 113 185
rect 111 184 112 185
rect 110 184 111 185
rect 109 184 110 185
rect 108 184 109 185
rect 107 184 108 185
rect 106 184 107 185
rect 105 184 106 185
rect 104 184 105 185
rect 103 184 104 185
rect 102 184 103 185
rect 62 184 63 185
rect 61 184 62 185
rect 60 184 61 185
rect 59 184 60 185
rect 29 184 30 185
rect 28 184 29 185
rect 27 184 28 185
rect 26 184 27 185
rect 18 184 19 185
rect 196 185 197 186
rect 195 185 196 186
rect 194 185 195 186
rect 193 185 194 186
rect 192 185 193 186
rect 191 185 192 186
rect 190 185 191 186
rect 189 185 190 186
rect 188 185 189 186
rect 183 185 184 186
rect 182 185 183 186
rect 181 185 182 186
rect 180 185 181 186
rect 179 185 180 186
rect 178 185 179 186
rect 175 185 176 186
rect 174 185 175 186
rect 170 185 171 186
rect 169 185 170 186
rect 168 185 169 186
rect 167 185 168 186
rect 166 185 167 186
rect 165 185 166 186
rect 163 185 164 186
rect 162 185 163 186
rect 149 185 150 186
rect 148 185 149 186
rect 147 185 148 186
rect 146 185 147 186
rect 145 185 146 186
rect 144 185 145 186
rect 143 185 144 186
rect 142 185 143 186
rect 141 185 142 186
rect 140 185 141 186
rect 139 185 140 186
rect 138 185 139 186
rect 137 185 138 186
rect 136 185 137 186
rect 135 185 136 186
rect 134 185 135 186
rect 133 185 134 186
rect 132 185 133 186
rect 131 185 132 186
rect 130 185 131 186
rect 129 185 130 186
rect 128 185 129 186
rect 127 185 128 186
rect 126 185 127 186
rect 125 185 126 186
rect 124 185 125 186
rect 123 185 124 186
rect 122 185 123 186
rect 121 185 122 186
rect 120 185 121 186
rect 119 185 120 186
rect 118 185 119 186
rect 117 185 118 186
rect 116 185 117 186
rect 115 185 116 186
rect 114 185 115 186
rect 113 185 114 186
rect 112 185 113 186
rect 111 185 112 186
rect 110 185 111 186
rect 109 185 110 186
rect 108 185 109 186
rect 107 185 108 186
rect 106 185 107 186
rect 105 185 106 186
rect 104 185 105 186
rect 103 185 104 186
rect 102 185 103 186
rect 78 185 79 186
rect 77 185 78 186
rect 76 185 77 186
rect 75 185 76 186
rect 74 185 75 186
rect 73 185 74 186
rect 72 185 73 186
rect 71 185 72 186
rect 70 185 71 186
rect 69 185 70 186
rect 68 185 69 186
rect 67 185 68 186
rect 66 185 67 186
rect 65 185 66 186
rect 64 185 65 186
rect 63 185 64 186
rect 62 185 63 186
rect 61 185 62 186
rect 60 185 61 186
rect 59 185 60 186
rect 58 185 59 186
rect 57 185 58 186
rect 56 185 57 186
rect 55 185 56 186
rect 54 185 55 186
rect 29 185 30 186
rect 28 185 29 186
rect 27 185 28 186
rect 26 185 27 186
rect 25 185 26 186
rect 19 185 20 186
rect 18 185 19 186
rect 17 185 18 186
rect 196 186 197 187
rect 195 186 196 187
rect 194 186 195 187
rect 193 186 194 187
rect 192 186 193 187
rect 191 186 192 187
rect 190 186 191 187
rect 189 186 190 187
rect 188 186 189 187
rect 183 186 184 187
rect 182 186 183 187
rect 181 186 182 187
rect 180 186 181 187
rect 175 186 176 187
rect 174 186 175 187
rect 170 186 171 187
rect 169 186 170 187
rect 168 186 169 187
rect 167 186 168 187
rect 166 186 167 187
rect 165 186 166 187
rect 163 186 164 187
rect 162 186 163 187
rect 149 186 150 187
rect 148 186 149 187
rect 147 186 148 187
rect 146 186 147 187
rect 145 186 146 187
rect 144 186 145 187
rect 143 186 144 187
rect 142 186 143 187
rect 141 186 142 187
rect 140 186 141 187
rect 139 186 140 187
rect 138 186 139 187
rect 137 186 138 187
rect 136 186 137 187
rect 135 186 136 187
rect 134 186 135 187
rect 133 186 134 187
rect 132 186 133 187
rect 131 186 132 187
rect 130 186 131 187
rect 129 186 130 187
rect 128 186 129 187
rect 127 186 128 187
rect 126 186 127 187
rect 125 186 126 187
rect 124 186 125 187
rect 123 186 124 187
rect 122 186 123 187
rect 121 186 122 187
rect 120 186 121 187
rect 119 186 120 187
rect 118 186 119 187
rect 117 186 118 187
rect 116 186 117 187
rect 115 186 116 187
rect 114 186 115 187
rect 113 186 114 187
rect 112 186 113 187
rect 111 186 112 187
rect 110 186 111 187
rect 109 186 110 187
rect 108 186 109 187
rect 107 186 108 187
rect 106 186 107 187
rect 105 186 106 187
rect 104 186 105 187
rect 103 186 104 187
rect 102 186 103 187
rect 78 186 79 187
rect 77 186 78 187
rect 76 186 77 187
rect 75 186 76 187
rect 74 186 75 187
rect 73 186 74 187
rect 72 186 73 187
rect 71 186 72 187
rect 70 186 71 187
rect 69 186 70 187
rect 68 186 69 187
rect 67 186 68 187
rect 66 186 67 187
rect 65 186 66 187
rect 64 186 65 187
rect 63 186 64 187
rect 62 186 63 187
rect 61 186 62 187
rect 60 186 61 187
rect 59 186 60 187
rect 58 186 59 187
rect 57 186 58 187
rect 56 186 57 187
rect 55 186 56 187
rect 54 186 55 187
rect 53 186 54 187
rect 52 186 53 187
rect 29 186 30 187
rect 28 186 29 187
rect 27 186 28 187
rect 26 186 27 187
rect 25 186 26 187
rect 24 186 25 187
rect 19 186 20 187
rect 18 186 19 187
rect 17 186 18 187
rect 16 186 17 187
rect 183 187 184 188
rect 182 187 183 188
rect 181 187 182 188
rect 180 187 181 188
rect 175 187 176 188
rect 174 187 175 188
rect 173 187 174 188
rect 171 187 172 188
rect 170 187 171 188
rect 169 187 170 188
rect 168 187 169 188
rect 167 187 168 188
rect 166 187 167 188
rect 165 187 166 188
rect 163 187 164 188
rect 162 187 163 188
rect 149 187 150 188
rect 148 187 149 188
rect 147 187 148 188
rect 146 187 147 188
rect 145 187 146 188
rect 144 187 145 188
rect 143 187 144 188
rect 142 187 143 188
rect 141 187 142 188
rect 140 187 141 188
rect 139 187 140 188
rect 138 187 139 188
rect 137 187 138 188
rect 136 187 137 188
rect 135 187 136 188
rect 134 187 135 188
rect 133 187 134 188
rect 132 187 133 188
rect 131 187 132 188
rect 130 187 131 188
rect 129 187 130 188
rect 128 187 129 188
rect 127 187 128 188
rect 126 187 127 188
rect 125 187 126 188
rect 124 187 125 188
rect 123 187 124 188
rect 122 187 123 188
rect 121 187 122 188
rect 120 187 121 188
rect 119 187 120 188
rect 118 187 119 188
rect 117 187 118 188
rect 116 187 117 188
rect 115 187 116 188
rect 114 187 115 188
rect 113 187 114 188
rect 112 187 113 188
rect 111 187 112 188
rect 110 187 111 188
rect 109 187 110 188
rect 108 187 109 188
rect 107 187 108 188
rect 106 187 107 188
rect 105 187 106 188
rect 104 187 105 188
rect 103 187 104 188
rect 102 187 103 188
rect 78 187 79 188
rect 77 187 78 188
rect 76 187 77 188
rect 75 187 76 188
rect 74 187 75 188
rect 73 187 74 188
rect 72 187 73 188
rect 71 187 72 188
rect 70 187 71 188
rect 69 187 70 188
rect 68 187 69 188
rect 67 187 68 188
rect 66 187 67 188
rect 65 187 66 188
rect 64 187 65 188
rect 63 187 64 188
rect 62 187 63 188
rect 61 187 62 188
rect 60 187 61 188
rect 59 187 60 188
rect 58 187 59 188
rect 57 187 58 188
rect 56 187 57 188
rect 55 187 56 188
rect 54 187 55 188
rect 53 187 54 188
rect 52 187 53 188
rect 29 187 30 188
rect 28 187 29 188
rect 27 187 28 188
rect 26 187 27 188
rect 25 187 26 188
rect 24 187 25 188
rect 23 187 24 188
rect 19 187 20 188
rect 18 187 19 188
rect 17 187 18 188
rect 16 187 17 188
rect 15 187 16 188
rect 196 188 197 189
rect 195 188 196 189
rect 194 188 195 189
rect 193 188 194 189
rect 192 188 193 189
rect 183 188 184 189
rect 182 188 183 189
rect 181 188 182 189
rect 180 188 181 189
rect 175 188 176 189
rect 174 188 175 189
rect 173 188 174 189
rect 171 188 172 189
rect 170 188 171 189
rect 169 188 170 189
rect 168 188 169 189
rect 167 188 168 189
rect 166 188 167 189
rect 165 188 166 189
rect 163 188 164 189
rect 162 188 163 189
rect 149 188 150 189
rect 148 188 149 189
rect 147 188 148 189
rect 146 188 147 189
rect 145 188 146 189
rect 144 188 145 189
rect 143 188 144 189
rect 142 188 143 189
rect 141 188 142 189
rect 140 188 141 189
rect 139 188 140 189
rect 138 188 139 189
rect 137 188 138 189
rect 136 188 137 189
rect 135 188 136 189
rect 134 188 135 189
rect 133 188 134 189
rect 132 188 133 189
rect 131 188 132 189
rect 130 188 131 189
rect 129 188 130 189
rect 128 188 129 189
rect 127 188 128 189
rect 126 188 127 189
rect 125 188 126 189
rect 124 188 125 189
rect 123 188 124 189
rect 122 188 123 189
rect 121 188 122 189
rect 120 188 121 189
rect 119 188 120 189
rect 118 188 119 189
rect 117 188 118 189
rect 116 188 117 189
rect 115 188 116 189
rect 114 188 115 189
rect 113 188 114 189
rect 112 188 113 189
rect 111 188 112 189
rect 110 188 111 189
rect 109 188 110 189
rect 108 188 109 189
rect 107 188 108 189
rect 106 188 107 189
rect 105 188 106 189
rect 104 188 105 189
rect 103 188 104 189
rect 102 188 103 189
rect 78 188 79 189
rect 77 188 78 189
rect 76 188 77 189
rect 75 188 76 189
rect 74 188 75 189
rect 73 188 74 189
rect 72 188 73 189
rect 71 188 72 189
rect 70 188 71 189
rect 69 188 70 189
rect 68 188 69 189
rect 67 188 68 189
rect 66 188 67 189
rect 65 188 66 189
rect 64 188 65 189
rect 63 188 64 189
rect 62 188 63 189
rect 61 188 62 189
rect 60 188 61 189
rect 59 188 60 189
rect 58 188 59 189
rect 57 188 58 189
rect 56 188 57 189
rect 55 188 56 189
rect 54 188 55 189
rect 53 188 54 189
rect 52 188 53 189
rect 51 188 52 189
rect 29 188 30 189
rect 28 188 29 189
rect 27 188 28 189
rect 25 188 26 189
rect 24 188 25 189
rect 23 188 24 189
rect 22 188 23 189
rect 17 188 18 189
rect 16 188 17 189
rect 15 188 16 189
rect 196 189 197 190
rect 195 189 196 190
rect 194 189 195 190
rect 193 189 194 190
rect 192 189 193 190
rect 191 189 192 190
rect 183 189 184 190
rect 182 189 183 190
rect 181 189 182 190
rect 180 189 181 190
rect 175 189 176 190
rect 174 189 175 190
rect 173 189 174 190
rect 172 189 173 190
rect 171 189 172 190
rect 170 189 171 190
rect 169 189 170 190
rect 167 189 168 190
rect 166 189 167 190
rect 165 189 166 190
rect 163 189 164 190
rect 162 189 163 190
rect 149 189 150 190
rect 148 189 149 190
rect 147 189 148 190
rect 146 189 147 190
rect 145 189 146 190
rect 144 189 145 190
rect 143 189 144 190
rect 142 189 143 190
rect 141 189 142 190
rect 140 189 141 190
rect 139 189 140 190
rect 138 189 139 190
rect 137 189 138 190
rect 136 189 137 190
rect 135 189 136 190
rect 134 189 135 190
rect 133 189 134 190
rect 132 189 133 190
rect 131 189 132 190
rect 130 189 131 190
rect 129 189 130 190
rect 128 189 129 190
rect 127 189 128 190
rect 126 189 127 190
rect 125 189 126 190
rect 124 189 125 190
rect 123 189 124 190
rect 122 189 123 190
rect 121 189 122 190
rect 120 189 121 190
rect 119 189 120 190
rect 118 189 119 190
rect 117 189 118 190
rect 116 189 117 190
rect 115 189 116 190
rect 114 189 115 190
rect 113 189 114 190
rect 112 189 113 190
rect 111 189 112 190
rect 110 189 111 190
rect 109 189 110 190
rect 108 189 109 190
rect 107 189 108 190
rect 106 189 107 190
rect 105 189 106 190
rect 104 189 105 190
rect 103 189 104 190
rect 102 189 103 190
rect 78 189 79 190
rect 77 189 78 190
rect 76 189 77 190
rect 75 189 76 190
rect 74 189 75 190
rect 73 189 74 190
rect 72 189 73 190
rect 71 189 72 190
rect 70 189 71 190
rect 69 189 70 190
rect 68 189 69 190
rect 67 189 68 190
rect 66 189 67 190
rect 65 189 66 190
rect 64 189 65 190
rect 63 189 64 190
rect 62 189 63 190
rect 61 189 62 190
rect 60 189 61 190
rect 59 189 60 190
rect 58 189 59 190
rect 57 189 58 190
rect 56 189 57 190
rect 55 189 56 190
rect 54 189 55 190
rect 53 189 54 190
rect 52 189 53 190
rect 51 189 52 190
rect 29 189 30 190
rect 28 189 29 190
rect 27 189 28 190
rect 24 189 25 190
rect 23 189 24 190
rect 22 189 23 190
rect 21 189 22 190
rect 17 189 18 190
rect 16 189 17 190
rect 15 189 16 190
rect 197 190 198 191
rect 196 190 197 191
rect 194 190 195 191
rect 192 190 193 191
rect 191 190 192 191
rect 183 190 184 191
rect 182 190 183 191
rect 181 190 182 191
rect 180 190 181 191
rect 175 190 176 191
rect 174 190 175 191
rect 173 190 174 191
rect 172 190 173 191
rect 171 190 172 191
rect 170 190 171 191
rect 169 190 170 191
rect 167 190 168 191
rect 166 190 167 191
rect 165 190 166 191
rect 149 190 150 191
rect 148 190 149 191
rect 147 190 148 191
rect 146 190 147 191
rect 145 190 146 191
rect 144 190 145 191
rect 143 190 144 191
rect 142 190 143 191
rect 141 190 142 191
rect 140 190 141 191
rect 139 190 140 191
rect 138 190 139 191
rect 137 190 138 191
rect 136 190 137 191
rect 135 190 136 191
rect 134 190 135 191
rect 133 190 134 191
rect 132 190 133 191
rect 131 190 132 191
rect 130 190 131 191
rect 129 190 130 191
rect 128 190 129 191
rect 127 190 128 191
rect 126 190 127 191
rect 125 190 126 191
rect 124 190 125 191
rect 123 190 124 191
rect 122 190 123 191
rect 121 190 122 191
rect 120 190 121 191
rect 119 190 120 191
rect 118 190 119 191
rect 117 190 118 191
rect 116 190 117 191
rect 115 190 116 191
rect 114 190 115 191
rect 113 190 114 191
rect 112 190 113 191
rect 111 190 112 191
rect 110 190 111 191
rect 109 190 110 191
rect 108 190 109 191
rect 107 190 108 191
rect 106 190 107 191
rect 105 190 106 191
rect 104 190 105 191
rect 103 190 104 191
rect 102 190 103 191
rect 78 190 79 191
rect 77 190 78 191
rect 76 190 77 191
rect 75 190 76 191
rect 74 190 75 191
rect 73 190 74 191
rect 72 190 73 191
rect 71 190 72 191
rect 70 190 71 191
rect 69 190 70 191
rect 68 190 69 191
rect 67 190 68 191
rect 66 190 67 191
rect 65 190 66 191
rect 64 190 65 191
rect 63 190 64 191
rect 62 190 63 191
rect 61 190 62 191
rect 60 190 61 191
rect 59 190 60 191
rect 58 190 59 191
rect 57 190 58 191
rect 56 190 57 191
rect 55 190 56 191
rect 54 190 55 191
rect 53 190 54 191
rect 52 190 53 191
rect 51 190 52 191
rect 29 190 30 191
rect 28 190 29 191
rect 27 190 28 191
rect 23 190 24 191
rect 22 190 23 191
rect 21 190 22 191
rect 20 190 21 191
rect 17 190 18 191
rect 16 190 17 191
rect 15 190 16 191
rect 197 191 198 192
rect 196 191 197 192
rect 194 191 195 192
rect 193 191 194 192
rect 192 191 193 192
rect 191 191 192 192
rect 183 191 184 192
rect 182 191 183 192
rect 181 191 182 192
rect 180 191 181 192
rect 174 191 175 192
rect 173 191 174 192
rect 172 191 173 192
rect 171 191 172 192
rect 170 191 171 192
rect 167 191 168 192
rect 166 191 167 192
rect 165 191 166 192
rect 149 191 150 192
rect 148 191 149 192
rect 147 191 148 192
rect 146 191 147 192
rect 145 191 146 192
rect 144 191 145 192
rect 143 191 144 192
rect 142 191 143 192
rect 141 191 142 192
rect 140 191 141 192
rect 139 191 140 192
rect 138 191 139 192
rect 137 191 138 192
rect 136 191 137 192
rect 135 191 136 192
rect 134 191 135 192
rect 133 191 134 192
rect 132 191 133 192
rect 131 191 132 192
rect 130 191 131 192
rect 129 191 130 192
rect 128 191 129 192
rect 127 191 128 192
rect 126 191 127 192
rect 125 191 126 192
rect 124 191 125 192
rect 123 191 124 192
rect 122 191 123 192
rect 121 191 122 192
rect 120 191 121 192
rect 119 191 120 192
rect 118 191 119 192
rect 117 191 118 192
rect 116 191 117 192
rect 115 191 116 192
rect 114 191 115 192
rect 113 191 114 192
rect 112 191 113 192
rect 111 191 112 192
rect 110 191 111 192
rect 109 191 110 192
rect 108 191 109 192
rect 107 191 108 192
rect 106 191 107 192
rect 105 191 106 192
rect 104 191 105 192
rect 103 191 104 192
rect 102 191 103 192
rect 62 191 63 192
rect 61 191 62 192
rect 60 191 61 192
rect 59 191 60 192
rect 54 191 55 192
rect 53 191 54 192
rect 52 191 53 192
rect 51 191 52 192
rect 29 191 30 192
rect 28 191 29 192
rect 27 191 28 192
rect 22 191 23 192
rect 21 191 22 192
rect 20 191 21 192
rect 19 191 20 192
rect 18 191 19 192
rect 17 191 18 192
rect 16 191 17 192
rect 15 191 16 192
rect 196 192 197 193
rect 194 192 195 193
rect 193 192 194 193
rect 192 192 193 193
rect 191 192 192 193
rect 183 192 184 193
rect 182 192 183 193
rect 181 192 182 193
rect 180 192 181 193
rect 173 192 174 193
rect 172 192 173 193
rect 171 192 172 193
rect 167 192 168 193
rect 166 192 167 193
rect 165 192 166 193
rect 149 192 150 193
rect 148 192 149 193
rect 147 192 148 193
rect 146 192 147 193
rect 145 192 146 193
rect 144 192 145 193
rect 143 192 144 193
rect 142 192 143 193
rect 141 192 142 193
rect 140 192 141 193
rect 139 192 140 193
rect 138 192 139 193
rect 137 192 138 193
rect 136 192 137 193
rect 135 192 136 193
rect 134 192 135 193
rect 133 192 134 193
rect 132 192 133 193
rect 131 192 132 193
rect 130 192 131 193
rect 129 192 130 193
rect 128 192 129 193
rect 127 192 128 193
rect 126 192 127 193
rect 125 192 126 193
rect 124 192 125 193
rect 123 192 124 193
rect 122 192 123 193
rect 121 192 122 193
rect 120 192 121 193
rect 119 192 120 193
rect 118 192 119 193
rect 117 192 118 193
rect 116 192 117 193
rect 115 192 116 193
rect 114 192 115 193
rect 113 192 114 193
rect 112 192 113 193
rect 111 192 112 193
rect 110 192 111 193
rect 109 192 110 193
rect 108 192 109 193
rect 107 192 108 193
rect 106 192 107 193
rect 105 192 106 193
rect 104 192 105 193
rect 103 192 104 193
rect 102 192 103 193
rect 62 192 63 193
rect 61 192 62 193
rect 60 192 61 193
rect 59 192 60 193
rect 54 192 55 193
rect 53 192 54 193
rect 52 192 53 193
rect 51 192 52 193
rect 28 192 29 193
rect 27 192 28 193
rect 21 192 22 193
rect 20 192 21 193
rect 19 192 20 193
rect 18 192 19 193
rect 17 192 18 193
rect 16 192 17 193
rect 196 193 197 194
rect 194 193 195 194
rect 193 193 194 194
rect 183 193 184 194
rect 182 193 183 194
rect 181 193 182 194
rect 180 193 181 194
rect 166 193 167 194
rect 165 193 166 194
rect 149 193 150 194
rect 148 193 149 194
rect 147 193 148 194
rect 146 193 147 194
rect 145 193 146 194
rect 144 193 145 194
rect 143 193 144 194
rect 142 193 143 194
rect 141 193 142 194
rect 140 193 141 194
rect 139 193 140 194
rect 138 193 139 194
rect 137 193 138 194
rect 136 193 137 194
rect 135 193 136 194
rect 134 193 135 194
rect 133 193 134 194
rect 132 193 133 194
rect 131 193 132 194
rect 130 193 131 194
rect 129 193 130 194
rect 128 193 129 194
rect 127 193 128 194
rect 126 193 127 194
rect 125 193 126 194
rect 124 193 125 194
rect 123 193 124 194
rect 122 193 123 194
rect 121 193 122 194
rect 120 193 121 194
rect 119 193 120 194
rect 118 193 119 194
rect 117 193 118 194
rect 116 193 117 194
rect 115 193 116 194
rect 114 193 115 194
rect 113 193 114 194
rect 112 193 113 194
rect 111 193 112 194
rect 110 193 111 194
rect 109 193 110 194
rect 108 193 109 194
rect 107 193 108 194
rect 106 193 107 194
rect 105 193 106 194
rect 104 193 105 194
rect 103 193 104 194
rect 102 193 103 194
rect 62 193 63 194
rect 61 193 62 194
rect 60 193 61 194
rect 59 193 60 194
rect 54 193 55 194
rect 53 193 54 194
rect 52 193 53 194
rect 51 193 52 194
rect 20 193 21 194
rect 19 193 20 194
rect 18 193 19 194
rect 17 193 18 194
rect 195 194 196 195
rect 194 194 195 195
rect 193 194 194 195
rect 183 194 184 195
rect 182 194 183 195
rect 181 194 182 195
rect 180 194 181 195
rect 149 194 150 195
rect 148 194 149 195
rect 147 194 148 195
rect 146 194 147 195
rect 145 194 146 195
rect 144 194 145 195
rect 143 194 144 195
rect 142 194 143 195
rect 141 194 142 195
rect 140 194 141 195
rect 139 194 140 195
rect 138 194 139 195
rect 137 194 138 195
rect 136 194 137 195
rect 135 194 136 195
rect 134 194 135 195
rect 133 194 134 195
rect 132 194 133 195
rect 131 194 132 195
rect 130 194 131 195
rect 129 194 130 195
rect 128 194 129 195
rect 127 194 128 195
rect 126 194 127 195
rect 125 194 126 195
rect 124 194 125 195
rect 123 194 124 195
rect 122 194 123 195
rect 121 194 122 195
rect 120 194 121 195
rect 119 194 120 195
rect 118 194 119 195
rect 117 194 118 195
rect 116 194 117 195
rect 115 194 116 195
rect 114 194 115 195
rect 113 194 114 195
rect 112 194 113 195
rect 111 194 112 195
rect 110 194 111 195
rect 109 194 110 195
rect 108 194 109 195
rect 107 194 108 195
rect 106 194 107 195
rect 105 194 106 195
rect 104 194 105 195
rect 103 194 104 195
rect 102 194 103 195
rect 62 194 63 195
rect 61 194 62 195
rect 60 194 61 195
rect 59 194 60 195
rect 54 194 55 195
rect 53 194 54 195
rect 52 194 53 195
rect 51 194 52 195
rect 196 195 197 196
rect 195 195 196 196
rect 194 195 195 196
rect 193 195 194 196
rect 192 195 193 196
rect 191 195 192 196
rect 183 195 184 196
rect 182 195 183 196
rect 181 195 182 196
rect 180 195 181 196
rect 149 195 150 196
rect 148 195 149 196
rect 147 195 148 196
rect 146 195 147 196
rect 145 195 146 196
rect 144 195 145 196
rect 143 195 144 196
rect 142 195 143 196
rect 141 195 142 196
rect 140 195 141 196
rect 139 195 140 196
rect 138 195 139 196
rect 137 195 138 196
rect 136 195 137 196
rect 135 195 136 196
rect 134 195 135 196
rect 133 195 134 196
rect 132 195 133 196
rect 131 195 132 196
rect 130 195 131 196
rect 129 195 130 196
rect 128 195 129 196
rect 127 195 128 196
rect 126 195 127 196
rect 125 195 126 196
rect 124 195 125 196
rect 123 195 124 196
rect 122 195 123 196
rect 121 195 122 196
rect 120 195 121 196
rect 119 195 120 196
rect 118 195 119 196
rect 117 195 118 196
rect 116 195 117 196
rect 115 195 116 196
rect 114 195 115 196
rect 113 195 114 196
rect 112 195 113 196
rect 111 195 112 196
rect 110 195 111 196
rect 109 195 110 196
rect 108 195 109 196
rect 107 195 108 196
rect 106 195 107 196
rect 105 195 106 196
rect 104 195 105 196
rect 103 195 104 196
rect 102 195 103 196
rect 53 195 54 196
rect 52 195 53 196
rect 51 195 52 196
rect 27 195 28 196
rect 26 195 27 196
rect 25 195 26 196
rect 24 195 25 196
rect 23 195 24 196
rect 22 195 23 196
rect 21 195 22 196
rect 196 196 197 197
rect 195 196 196 197
rect 192 196 193 197
rect 191 196 192 197
rect 183 196 184 197
rect 182 196 183 197
rect 181 196 182 197
rect 180 196 181 197
rect 177 196 178 197
rect 176 196 177 197
rect 175 196 176 197
rect 174 196 175 197
rect 173 196 174 197
rect 172 196 173 197
rect 171 196 172 197
rect 170 196 171 197
rect 169 196 170 197
rect 168 196 169 197
rect 167 196 168 197
rect 166 196 167 197
rect 165 196 166 197
rect 164 196 165 197
rect 163 196 164 197
rect 162 196 163 197
rect 149 196 150 197
rect 148 196 149 197
rect 147 196 148 197
rect 146 196 147 197
rect 145 196 146 197
rect 144 196 145 197
rect 143 196 144 197
rect 142 196 143 197
rect 141 196 142 197
rect 140 196 141 197
rect 139 196 140 197
rect 138 196 139 197
rect 137 196 138 197
rect 136 196 137 197
rect 135 196 136 197
rect 134 196 135 197
rect 133 196 134 197
rect 132 196 133 197
rect 131 196 132 197
rect 130 196 131 197
rect 129 196 130 197
rect 128 196 129 197
rect 127 196 128 197
rect 126 196 127 197
rect 125 196 126 197
rect 124 196 125 197
rect 123 196 124 197
rect 122 196 123 197
rect 121 196 122 197
rect 120 196 121 197
rect 119 196 120 197
rect 118 196 119 197
rect 117 196 118 197
rect 116 196 117 197
rect 115 196 116 197
rect 114 196 115 197
rect 113 196 114 197
rect 112 196 113 197
rect 111 196 112 197
rect 110 196 111 197
rect 109 196 110 197
rect 108 196 109 197
rect 107 196 108 197
rect 106 196 107 197
rect 105 196 106 197
rect 104 196 105 197
rect 103 196 104 197
rect 102 196 103 197
rect 28 196 29 197
rect 27 196 28 197
rect 26 196 27 197
rect 25 196 26 197
rect 24 196 25 197
rect 23 196 24 197
rect 22 196 23 197
rect 21 196 22 197
rect 20 196 21 197
rect 19 196 20 197
rect 18 196 19 197
rect 197 197 198 198
rect 196 197 197 198
rect 192 197 193 198
rect 191 197 192 198
rect 183 197 184 198
rect 182 197 183 198
rect 181 197 182 198
rect 180 197 181 198
rect 177 197 178 198
rect 176 197 177 198
rect 175 197 176 198
rect 174 197 175 198
rect 173 197 174 198
rect 172 197 173 198
rect 171 197 172 198
rect 170 197 171 198
rect 169 197 170 198
rect 168 197 169 198
rect 167 197 168 198
rect 166 197 167 198
rect 165 197 166 198
rect 164 197 165 198
rect 163 197 164 198
rect 162 197 163 198
rect 149 197 150 198
rect 148 197 149 198
rect 147 197 148 198
rect 146 197 147 198
rect 145 197 146 198
rect 144 197 145 198
rect 143 197 144 198
rect 142 197 143 198
rect 141 197 142 198
rect 140 197 141 198
rect 139 197 140 198
rect 138 197 139 198
rect 137 197 138 198
rect 136 197 137 198
rect 135 197 136 198
rect 134 197 135 198
rect 133 197 134 198
rect 132 197 133 198
rect 131 197 132 198
rect 130 197 131 198
rect 129 197 130 198
rect 128 197 129 198
rect 127 197 128 198
rect 126 197 127 198
rect 125 197 126 198
rect 124 197 125 198
rect 123 197 124 198
rect 122 197 123 198
rect 121 197 122 198
rect 120 197 121 198
rect 119 197 120 198
rect 118 197 119 198
rect 117 197 118 198
rect 116 197 117 198
rect 115 197 116 198
rect 114 197 115 198
rect 113 197 114 198
rect 112 197 113 198
rect 111 197 112 198
rect 110 197 111 198
rect 109 197 110 198
rect 108 197 109 198
rect 107 197 108 198
rect 106 197 107 198
rect 105 197 106 198
rect 104 197 105 198
rect 103 197 104 198
rect 102 197 103 198
rect 78 197 79 198
rect 77 197 78 198
rect 76 197 77 198
rect 75 197 76 198
rect 74 197 75 198
rect 73 197 74 198
rect 72 197 73 198
rect 71 197 72 198
rect 70 197 71 198
rect 69 197 70 198
rect 68 197 69 198
rect 67 197 68 198
rect 66 197 67 198
rect 65 197 66 198
rect 64 197 65 198
rect 63 197 64 198
rect 62 197 63 198
rect 61 197 62 198
rect 60 197 61 198
rect 59 197 60 198
rect 55 197 56 198
rect 54 197 55 198
rect 53 197 54 198
rect 52 197 53 198
rect 51 197 52 198
rect 29 197 30 198
rect 28 197 29 198
rect 27 197 28 198
rect 26 197 27 198
rect 25 197 26 198
rect 24 197 25 198
rect 23 197 24 198
rect 22 197 23 198
rect 21 197 22 198
rect 20 197 21 198
rect 19 197 20 198
rect 18 197 19 198
rect 17 197 18 198
rect 197 198 198 199
rect 196 198 197 199
rect 192 198 193 199
rect 191 198 192 199
rect 183 198 184 199
rect 182 198 183 199
rect 181 198 182 199
rect 180 198 181 199
rect 177 198 178 199
rect 176 198 177 199
rect 175 198 176 199
rect 174 198 175 199
rect 173 198 174 199
rect 172 198 173 199
rect 171 198 172 199
rect 170 198 171 199
rect 169 198 170 199
rect 168 198 169 199
rect 167 198 168 199
rect 166 198 167 199
rect 165 198 166 199
rect 164 198 165 199
rect 163 198 164 199
rect 162 198 163 199
rect 149 198 150 199
rect 148 198 149 199
rect 147 198 148 199
rect 146 198 147 199
rect 145 198 146 199
rect 144 198 145 199
rect 143 198 144 199
rect 142 198 143 199
rect 141 198 142 199
rect 140 198 141 199
rect 139 198 140 199
rect 138 198 139 199
rect 137 198 138 199
rect 136 198 137 199
rect 135 198 136 199
rect 134 198 135 199
rect 133 198 134 199
rect 132 198 133 199
rect 131 198 132 199
rect 130 198 131 199
rect 129 198 130 199
rect 128 198 129 199
rect 127 198 128 199
rect 126 198 127 199
rect 125 198 126 199
rect 124 198 125 199
rect 123 198 124 199
rect 122 198 123 199
rect 121 198 122 199
rect 120 198 121 199
rect 119 198 120 199
rect 118 198 119 199
rect 117 198 118 199
rect 116 198 117 199
rect 115 198 116 199
rect 114 198 115 199
rect 113 198 114 199
rect 112 198 113 199
rect 111 198 112 199
rect 110 198 111 199
rect 109 198 110 199
rect 108 198 109 199
rect 107 198 108 199
rect 106 198 107 199
rect 105 198 106 199
rect 104 198 105 199
rect 103 198 104 199
rect 102 198 103 199
rect 78 198 79 199
rect 77 198 78 199
rect 76 198 77 199
rect 75 198 76 199
rect 74 198 75 199
rect 73 198 74 199
rect 72 198 73 199
rect 71 198 72 199
rect 70 198 71 199
rect 69 198 70 199
rect 68 198 69 199
rect 67 198 68 199
rect 66 198 67 199
rect 65 198 66 199
rect 64 198 65 199
rect 63 198 64 199
rect 62 198 63 199
rect 61 198 62 199
rect 60 198 61 199
rect 59 198 60 199
rect 55 198 56 199
rect 54 198 55 199
rect 53 198 54 199
rect 52 198 53 199
rect 51 198 52 199
rect 29 198 30 199
rect 28 198 29 199
rect 27 198 28 199
rect 21 198 22 199
rect 20 198 21 199
rect 19 198 20 199
rect 18 198 19 199
rect 17 198 18 199
rect 16 198 17 199
rect 191 199 192 200
rect 182 199 183 200
rect 181 199 182 200
rect 170 199 171 200
rect 169 199 170 200
rect 168 199 169 200
rect 149 199 150 200
rect 148 199 149 200
rect 147 199 148 200
rect 146 199 147 200
rect 145 199 146 200
rect 144 199 145 200
rect 143 199 144 200
rect 142 199 143 200
rect 141 199 142 200
rect 140 199 141 200
rect 139 199 140 200
rect 137 199 138 200
rect 136 199 137 200
rect 135 199 136 200
rect 134 199 135 200
rect 133 199 134 200
rect 132 199 133 200
rect 131 199 132 200
rect 130 199 131 200
rect 129 199 130 200
rect 128 199 129 200
rect 127 199 128 200
rect 126 199 127 200
rect 125 199 126 200
rect 124 199 125 200
rect 123 199 124 200
rect 122 199 123 200
rect 121 199 122 200
rect 120 199 121 200
rect 118 199 119 200
rect 117 199 118 200
rect 116 199 117 200
rect 115 199 116 200
rect 114 199 115 200
rect 112 199 113 200
rect 111 199 112 200
rect 110 199 111 200
rect 109 199 110 200
rect 108 199 109 200
rect 107 199 108 200
rect 106 199 107 200
rect 105 199 106 200
rect 104 199 105 200
rect 103 199 104 200
rect 102 199 103 200
rect 78 199 79 200
rect 77 199 78 200
rect 76 199 77 200
rect 75 199 76 200
rect 74 199 75 200
rect 73 199 74 200
rect 72 199 73 200
rect 71 199 72 200
rect 70 199 71 200
rect 69 199 70 200
rect 68 199 69 200
rect 67 199 68 200
rect 66 199 67 200
rect 65 199 66 200
rect 64 199 65 200
rect 63 199 64 200
rect 62 199 63 200
rect 61 199 62 200
rect 60 199 61 200
rect 59 199 60 200
rect 55 199 56 200
rect 54 199 55 200
rect 53 199 54 200
rect 52 199 53 200
rect 51 199 52 200
rect 29 199 30 200
rect 28 199 29 200
rect 27 199 28 200
rect 18 199 19 200
rect 17 199 18 200
rect 16 199 17 200
rect 15 199 16 200
rect 195 200 196 201
rect 194 200 195 201
rect 193 200 194 201
rect 192 200 193 201
rect 191 200 192 201
rect 190 200 191 201
rect 170 200 171 201
rect 169 200 170 201
rect 168 200 169 201
rect 149 200 150 201
rect 148 200 149 201
rect 147 200 148 201
rect 146 200 147 201
rect 145 200 146 201
rect 144 200 145 201
rect 143 200 144 201
rect 142 200 143 201
rect 141 200 142 201
rect 140 200 141 201
rect 131 200 132 201
rect 130 200 131 201
rect 129 200 130 201
rect 128 200 129 201
rect 127 200 128 201
rect 126 200 127 201
rect 125 200 126 201
rect 124 200 125 201
rect 123 200 124 201
rect 122 200 123 201
rect 121 200 122 201
rect 112 200 113 201
rect 111 200 112 201
rect 110 200 111 201
rect 109 200 110 201
rect 108 200 109 201
rect 107 200 108 201
rect 106 200 107 201
rect 105 200 106 201
rect 104 200 105 201
rect 103 200 104 201
rect 102 200 103 201
rect 78 200 79 201
rect 77 200 78 201
rect 76 200 77 201
rect 75 200 76 201
rect 74 200 75 201
rect 73 200 74 201
rect 72 200 73 201
rect 71 200 72 201
rect 70 200 71 201
rect 69 200 70 201
rect 68 200 69 201
rect 67 200 68 201
rect 66 200 67 201
rect 65 200 66 201
rect 64 200 65 201
rect 63 200 64 201
rect 62 200 63 201
rect 61 200 62 201
rect 60 200 61 201
rect 59 200 60 201
rect 55 200 56 201
rect 54 200 55 201
rect 53 200 54 201
rect 52 200 53 201
rect 51 200 52 201
rect 29 200 30 201
rect 28 200 29 201
rect 27 200 28 201
rect 17 200 18 201
rect 16 200 17 201
rect 15 200 16 201
rect 196 201 197 202
rect 195 201 196 202
rect 194 201 195 202
rect 193 201 194 202
rect 192 201 193 202
rect 191 201 192 202
rect 190 201 191 202
rect 189 201 190 202
rect 170 201 171 202
rect 169 201 170 202
rect 168 201 169 202
rect 149 201 150 202
rect 148 201 149 202
rect 147 201 148 202
rect 146 201 147 202
rect 145 201 146 202
rect 144 201 145 202
rect 143 201 144 202
rect 142 201 143 202
rect 141 201 142 202
rect 140 201 141 202
rect 130 201 131 202
rect 129 201 130 202
rect 128 201 129 202
rect 127 201 128 202
rect 126 201 127 202
rect 125 201 126 202
rect 124 201 125 202
rect 123 201 124 202
rect 122 201 123 202
rect 121 201 122 202
rect 112 201 113 202
rect 111 201 112 202
rect 110 201 111 202
rect 109 201 110 202
rect 108 201 109 202
rect 107 201 108 202
rect 106 201 107 202
rect 105 201 106 202
rect 104 201 105 202
rect 103 201 104 202
rect 102 201 103 202
rect 78 201 79 202
rect 77 201 78 202
rect 76 201 77 202
rect 75 201 76 202
rect 74 201 75 202
rect 73 201 74 202
rect 72 201 73 202
rect 71 201 72 202
rect 70 201 71 202
rect 69 201 70 202
rect 68 201 69 202
rect 67 201 68 202
rect 66 201 67 202
rect 65 201 66 202
rect 64 201 65 202
rect 63 201 64 202
rect 62 201 63 202
rect 61 201 62 202
rect 60 201 61 202
rect 59 201 60 202
rect 55 201 56 202
rect 54 201 55 202
rect 53 201 54 202
rect 52 201 53 202
rect 51 201 52 202
rect 28 201 29 202
rect 27 201 28 202
rect 26 201 27 202
rect 25 201 26 202
rect 17 201 18 202
rect 16 201 17 202
rect 15 201 16 202
rect 196 202 197 203
rect 195 202 196 203
rect 194 202 195 203
rect 193 202 194 203
rect 192 202 193 203
rect 191 202 192 203
rect 190 202 191 203
rect 189 202 190 203
rect 149 202 150 203
rect 148 202 149 203
rect 147 202 148 203
rect 146 202 147 203
rect 145 202 146 203
rect 144 202 145 203
rect 143 202 144 203
rect 142 202 143 203
rect 141 202 142 203
rect 140 202 141 203
rect 130 202 131 203
rect 129 202 130 203
rect 128 202 129 203
rect 127 202 128 203
rect 126 202 127 203
rect 125 202 126 203
rect 124 202 125 203
rect 123 202 124 203
rect 122 202 123 203
rect 121 202 122 203
rect 112 202 113 203
rect 111 202 112 203
rect 110 202 111 203
rect 109 202 110 203
rect 108 202 109 203
rect 107 202 108 203
rect 106 202 107 203
rect 105 202 106 203
rect 104 202 105 203
rect 103 202 104 203
rect 102 202 103 203
rect 78 202 79 203
rect 77 202 78 203
rect 76 202 77 203
rect 75 202 76 203
rect 74 202 75 203
rect 73 202 74 203
rect 72 202 73 203
rect 71 202 72 203
rect 70 202 71 203
rect 69 202 70 203
rect 68 202 69 203
rect 67 202 68 203
rect 66 202 67 203
rect 65 202 66 203
rect 64 202 65 203
rect 63 202 64 203
rect 62 202 63 203
rect 61 202 62 203
rect 60 202 61 203
rect 59 202 60 203
rect 55 202 56 203
rect 54 202 55 203
rect 53 202 54 203
rect 52 202 53 203
rect 51 202 52 203
rect 28 202 29 203
rect 27 202 28 203
rect 26 202 27 203
rect 25 202 26 203
rect 24 202 25 203
rect 23 202 24 203
rect 22 202 23 203
rect 21 202 22 203
rect 17 202 18 203
rect 16 202 17 203
rect 15 202 16 203
rect 196 203 197 204
rect 191 203 192 204
rect 149 203 150 204
rect 148 203 149 204
rect 147 203 148 204
rect 146 203 147 204
rect 145 203 146 204
rect 144 203 145 204
rect 143 203 144 204
rect 142 203 143 204
rect 141 203 142 204
rect 140 203 141 204
rect 130 203 131 204
rect 129 203 130 204
rect 128 203 129 204
rect 127 203 128 204
rect 126 203 127 204
rect 125 203 126 204
rect 124 203 125 204
rect 123 203 124 204
rect 122 203 123 204
rect 121 203 122 204
rect 112 203 113 204
rect 111 203 112 204
rect 110 203 111 204
rect 109 203 110 204
rect 108 203 109 204
rect 107 203 108 204
rect 106 203 107 204
rect 105 203 106 204
rect 104 203 105 204
rect 103 203 104 204
rect 102 203 103 204
rect 27 203 28 204
rect 26 203 27 204
rect 25 203 26 204
rect 24 203 25 204
rect 23 203 24 204
rect 22 203 23 204
rect 21 203 22 204
rect 20 203 21 204
rect 19 203 20 204
rect 18 203 19 204
rect 17 203 18 204
rect 16 203 17 204
rect 15 203 16 204
rect 196 204 197 205
rect 195 204 196 205
rect 194 204 195 205
rect 193 204 194 205
rect 192 204 193 205
rect 191 204 192 205
rect 149 204 150 205
rect 148 204 149 205
rect 147 204 148 205
rect 146 204 147 205
rect 145 204 146 205
rect 144 204 145 205
rect 143 204 144 205
rect 142 204 143 205
rect 141 204 142 205
rect 140 204 141 205
rect 130 204 131 205
rect 129 204 130 205
rect 128 204 129 205
rect 127 204 128 205
rect 126 204 127 205
rect 125 204 126 205
rect 124 204 125 205
rect 123 204 124 205
rect 122 204 123 205
rect 121 204 122 205
rect 112 204 113 205
rect 111 204 112 205
rect 110 204 111 205
rect 109 204 110 205
rect 108 204 109 205
rect 107 204 108 205
rect 106 204 107 205
rect 105 204 106 205
rect 104 204 105 205
rect 103 204 104 205
rect 102 204 103 205
rect 25 204 26 205
rect 24 204 25 205
rect 23 204 24 205
rect 22 204 23 205
rect 21 204 22 205
rect 20 204 21 205
rect 19 204 20 205
rect 18 204 19 205
rect 17 204 18 205
rect 16 204 17 205
rect 197 205 198 206
rect 196 205 197 206
rect 195 205 196 206
rect 194 205 195 206
rect 193 205 194 206
rect 192 205 193 206
rect 191 205 192 206
rect 149 205 150 206
rect 148 205 149 206
rect 147 205 148 206
rect 146 205 147 206
rect 145 205 146 206
rect 144 205 145 206
rect 143 205 144 206
rect 142 205 143 206
rect 141 205 142 206
rect 140 205 141 206
rect 130 205 131 206
rect 129 205 130 206
rect 128 205 129 206
rect 127 205 128 206
rect 126 205 127 206
rect 125 205 126 206
rect 124 205 125 206
rect 123 205 124 206
rect 122 205 123 206
rect 121 205 122 206
rect 112 205 113 206
rect 111 205 112 206
rect 110 205 111 206
rect 109 205 110 206
rect 108 205 109 206
rect 107 205 108 206
rect 106 205 107 206
rect 105 205 106 206
rect 104 205 105 206
rect 103 205 104 206
rect 102 205 103 206
rect 22 205 23 206
rect 21 205 22 206
rect 20 205 21 206
rect 19 205 20 206
rect 18 205 19 206
rect 196 206 197 207
rect 195 206 196 207
rect 194 206 195 207
rect 193 206 194 207
rect 192 206 193 207
rect 191 206 192 207
rect 149 206 150 207
rect 148 206 149 207
rect 147 206 148 207
rect 146 206 147 207
rect 145 206 146 207
rect 144 206 145 207
rect 143 206 144 207
rect 142 206 143 207
rect 141 206 142 207
rect 140 206 141 207
rect 130 206 131 207
rect 129 206 130 207
rect 128 206 129 207
rect 127 206 128 207
rect 126 206 127 207
rect 125 206 126 207
rect 124 206 125 207
rect 123 206 124 207
rect 122 206 123 207
rect 121 206 122 207
rect 112 206 113 207
rect 111 206 112 207
rect 110 206 111 207
rect 109 206 110 207
rect 108 206 109 207
rect 107 206 108 207
rect 106 206 107 207
rect 105 206 106 207
rect 104 206 105 207
rect 103 206 104 207
rect 102 206 103 207
rect 192 207 193 208
rect 191 207 192 208
rect 149 207 150 208
rect 148 207 149 208
rect 147 207 148 208
rect 146 207 147 208
rect 145 207 146 208
rect 144 207 145 208
rect 143 207 144 208
rect 142 207 143 208
rect 141 207 142 208
rect 140 207 141 208
rect 130 207 131 208
rect 129 207 130 208
rect 128 207 129 208
rect 127 207 128 208
rect 126 207 127 208
rect 125 207 126 208
rect 124 207 125 208
rect 123 207 124 208
rect 122 207 123 208
rect 121 207 122 208
rect 112 207 113 208
rect 111 207 112 208
rect 110 207 111 208
rect 109 207 110 208
rect 108 207 109 208
rect 107 207 108 208
rect 106 207 107 208
rect 105 207 106 208
rect 104 207 105 208
rect 103 207 104 208
rect 102 207 103 208
rect 29 207 30 208
rect 28 207 29 208
rect 27 207 28 208
rect 195 208 196 209
rect 194 208 195 209
rect 193 208 194 209
rect 192 208 193 209
rect 191 208 192 209
rect 149 208 150 209
rect 148 208 149 209
rect 147 208 148 209
rect 146 208 147 209
rect 145 208 146 209
rect 144 208 145 209
rect 143 208 144 209
rect 142 208 143 209
rect 141 208 142 209
rect 140 208 141 209
rect 130 208 131 209
rect 129 208 130 209
rect 128 208 129 209
rect 127 208 128 209
rect 126 208 127 209
rect 125 208 126 209
rect 124 208 125 209
rect 123 208 124 209
rect 122 208 123 209
rect 121 208 122 209
rect 112 208 113 209
rect 111 208 112 209
rect 110 208 111 209
rect 109 208 110 209
rect 108 208 109 209
rect 107 208 108 209
rect 106 208 107 209
rect 105 208 106 209
rect 104 208 105 209
rect 103 208 104 209
rect 102 208 103 209
rect 78 208 79 209
rect 77 208 78 209
rect 76 208 77 209
rect 75 208 76 209
rect 74 208 75 209
rect 73 208 74 209
rect 72 208 73 209
rect 71 208 72 209
rect 70 208 71 209
rect 69 208 70 209
rect 68 208 69 209
rect 67 208 68 209
rect 66 208 67 209
rect 65 208 66 209
rect 64 208 65 209
rect 63 208 64 209
rect 62 208 63 209
rect 61 208 62 209
rect 60 208 61 209
rect 59 208 60 209
rect 29 208 30 209
rect 28 208 29 209
rect 27 208 28 209
rect 26 208 27 209
rect 19 208 20 209
rect 18 208 19 209
rect 196 209 197 210
rect 195 209 196 210
rect 194 209 195 210
rect 193 209 194 210
rect 192 209 193 210
rect 149 209 150 210
rect 148 209 149 210
rect 147 209 148 210
rect 146 209 147 210
rect 145 209 146 210
rect 144 209 145 210
rect 143 209 144 210
rect 142 209 143 210
rect 141 209 142 210
rect 140 209 141 210
rect 130 209 131 210
rect 129 209 130 210
rect 128 209 129 210
rect 127 209 128 210
rect 126 209 127 210
rect 125 209 126 210
rect 124 209 125 210
rect 123 209 124 210
rect 122 209 123 210
rect 121 209 122 210
rect 112 209 113 210
rect 111 209 112 210
rect 110 209 111 210
rect 109 209 110 210
rect 108 209 109 210
rect 107 209 108 210
rect 106 209 107 210
rect 105 209 106 210
rect 104 209 105 210
rect 103 209 104 210
rect 102 209 103 210
rect 78 209 79 210
rect 77 209 78 210
rect 76 209 77 210
rect 75 209 76 210
rect 74 209 75 210
rect 73 209 74 210
rect 72 209 73 210
rect 71 209 72 210
rect 70 209 71 210
rect 69 209 70 210
rect 68 209 69 210
rect 67 209 68 210
rect 66 209 67 210
rect 65 209 66 210
rect 64 209 65 210
rect 63 209 64 210
rect 62 209 63 210
rect 61 209 62 210
rect 60 209 61 210
rect 59 209 60 210
rect 29 209 30 210
rect 28 209 29 210
rect 27 209 28 210
rect 26 209 27 210
rect 25 209 26 210
rect 19 209 20 210
rect 18 209 19 210
rect 17 209 18 210
rect 16 209 17 210
rect 196 210 197 211
rect 195 210 196 211
rect 194 210 195 211
rect 193 210 194 211
rect 192 210 193 211
rect 191 210 192 211
rect 149 210 150 211
rect 148 210 149 211
rect 147 210 148 211
rect 146 210 147 211
rect 145 210 146 211
rect 144 210 145 211
rect 143 210 144 211
rect 142 210 143 211
rect 141 210 142 211
rect 140 210 141 211
rect 130 210 131 211
rect 129 210 130 211
rect 128 210 129 211
rect 127 210 128 211
rect 126 210 127 211
rect 125 210 126 211
rect 124 210 125 211
rect 123 210 124 211
rect 122 210 123 211
rect 121 210 122 211
rect 112 210 113 211
rect 111 210 112 211
rect 110 210 111 211
rect 109 210 110 211
rect 108 210 109 211
rect 107 210 108 211
rect 106 210 107 211
rect 105 210 106 211
rect 104 210 105 211
rect 103 210 104 211
rect 102 210 103 211
rect 78 210 79 211
rect 77 210 78 211
rect 76 210 77 211
rect 75 210 76 211
rect 74 210 75 211
rect 73 210 74 211
rect 72 210 73 211
rect 71 210 72 211
rect 70 210 71 211
rect 69 210 70 211
rect 68 210 69 211
rect 67 210 68 211
rect 66 210 67 211
rect 65 210 66 211
rect 64 210 65 211
rect 63 210 64 211
rect 62 210 63 211
rect 61 210 62 211
rect 60 210 61 211
rect 59 210 60 211
rect 29 210 30 211
rect 28 210 29 211
rect 27 210 28 211
rect 26 210 27 211
rect 25 210 26 211
rect 24 210 25 211
rect 19 210 20 211
rect 18 210 19 211
rect 17 210 18 211
rect 16 210 17 211
rect 15 210 16 211
rect 197 211 198 212
rect 196 211 197 212
rect 192 211 193 212
rect 191 211 192 212
rect 171 211 172 212
rect 149 211 150 212
rect 148 211 149 212
rect 147 211 148 212
rect 146 211 147 212
rect 145 211 146 212
rect 144 211 145 212
rect 143 211 144 212
rect 142 211 143 212
rect 141 211 142 212
rect 140 211 141 212
rect 130 211 131 212
rect 129 211 130 212
rect 128 211 129 212
rect 127 211 128 212
rect 126 211 127 212
rect 125 211 126 212
rect 124 211 125 212
rect 123 211 124 212
rect 122 211 123 212
rect 121 211 122 212
rect 112 211 113 212
rect 111 211 112 212
rect 110 211 111 212
rect 109 211 110 212
rect 108 211 109 212
rect 107 211 108 212
rect 106 211 107 212
rect 105 211 106 212
rect 104 211 105 212
rect 103 211 104 212
rect 102 211 103 212
rect 78 211 79 212
rect 77 211 78 212
rect 76 211 77 212
rect 75 211 76 212
rect 74 211 75 212
rect 73 211 74 212
rect 72 211 73 212
rect 71 211 72 212
rect 70 211 71 212
rect 69 211 70 212
rect 68 211 69 212
rect 67 211 68 212
rect 66 211 67 212
rect 65 211 66 212
rect 64 211 65 212
rect 63 211 64 212
rect 62 211 63 212
rect 61 211 62 212
rect 60 211 61 212
rect 59 211 60 212
rect 29 211 30 212
rect 28 211 29 212
rect 27 211 28 212
rect 26 211 27 212
rect 25 211 26 212
rect 24 211 25 212
rect 23 211 24 212
rect 18 211 19 212
rect 17 211 18 212
rect 16 211 17 212
rect 15 211 16 212
rect 197 212 198 213
rect 196 212 197 213
rect 192 212 193 213
rect 191 212 192 213
rect 173 212 174 213
rect 172 212 173 213
rect 171 212 172 213
rect 170 212 171 213
rect 149 212 150 213
rect 148 212 149 213
rect 147 212 148 213
rect 146 212 147 213
rect 145 212 146 213
rect 144 212 145 213
rect 143 212 144 213
rect 142 212 143 213
rect 141 212 142 213
rect 140 212 141 213
rect 130 212 131 213
rect 129 212 130 213
rect 128 212 129 213
rect 127 212 128 213
rect 126 212 127 213
rect 125 212 126 213
rect 124 212 125 213
rect 123 212 124 213
rect 122 212 123 213
rect 121 212 122 213
rect 112 212 113 213
rect 111 212 112 213
rect 110 212 111 213
rect 109 212 110 213
rect 108 212 109 213
rect 107 212 108 213
rect 106 212 107 213
rect 105 212 106 213
rect 104 212 105 213
rect 103 212 104 213
rect 102 212 103 213
rect 78 212 79 213
rect 77 212 78 213
rect 76 212 77 213
rect 75 212 76 213
rect 74 212 75 213
rect 73 212 74 213
rect 72 212 73 213
rect 71 212 72 213
rect 70 212 71 213
rect 69 212 70 213
rect 68 212 69 213
rect 67 212 68 213
rect 66 212 67 213
rect 65 212 66 213
rect 64 212 65 213
rect 63 212 64 213
rect 62 212 63 213
rect 61 212 62 213
rect 60 212 61 213
rect 59 212 60 213
rect 29 212 30 213
rect 28 212 29 213
rect 27 212 28 213
rect 25 212 26 213
rect 24 212 25 213
rect 23 212 24 213
rect 22 212 23 213
rect 17 212 18 213
rect 16 212 17 213
rect 15 212 16 213
rect 196 213 197 214
rect 195 213 196 214
rect 194 213 195 214
rect 193 213 194 214
rect 192 213 193 214
rect 191 213 192 214
rect 173 213 174 214
rect 172 213 173 214
rect 171 213 172 214
rect 170 213 171 214
rect 149 213 150 214
rect 148 213 149 214
rect 147 213 148 214
rect 146 213 147 214
rect 145 213 146 214
rect 144 213 145 214
rect 143 213 144 214
rect 142 213 143 214
rect 141 213 142 214
rect 140 213 141 214
rect 130 213 131 214
rect 129 213 130 214
rect 128 213 129 214
rect 127 213 128 214
rect 126 213 127 214
rect 125 213 126 214
rect 124 213 125 214
rect 123 213 124 214
rect 122 213 123 214
rect 121 213 122 214
rect 112 213 113 214
rect 111 213 112 214
rect 110 213 111 214
rect 109 213 110 214
rect 108 213 109 214
rect 107 213 108 214
rect 106 213 107 214
rect 105 213 106 214
rect 104 213 105 214
rect 103 213 104 214
rect 102 213 103 214
rect 66 213 67 214
rect 65 213 66 214
rect 64 213 65 214
rect 63 213 64 214
rect 62 213 63 214
rect 61 213 62 214
rect 60 213 61 214
rect 29 213 30 214
rect 28 213 29 214
rect 27 213 28 214
rect 24 213 25 214
rect 23 213 24 214
rect 22 213 23 214
rect 21 213 22 214
rect 17 213 18 214
rect 16 213 17 214
rect 15 213 16 214
rect 196 214 197 215
rect 195 214 196 215
rect 194 214 195 215
rect 193 214 194 215
rect 192 214 193 215
rect 178 214 179 215
rect 177 214 178 215
rect 173 214 174 215
rect 172 214 173 215
rect 171 214 172 215
rect 170 214 171 215
rect 164 214 165 215
rect 163 214 164 215
rect 149 214 150 215
rect 148 214 149 215
rect 147 214 148 215
rect 146 214 147 215
rect 145 214 146 215
rect 144 214 145 215
rect 143 214 144 215
rect 142 214 143 215
rect 141 214 142 215
rect 140 214 141 215
rect 130 214 131 215
rect 129 214 130 215
rect 128 214 129 215
rect 127 214 128 215
rect 126 214 127 215
rect 125 214 126 215
rect 124 214 125 215
rect 123 214 124 215
rect 122 214 123 215
rect 121 214 122 215
rect 112 214 113 215
rect 111 214 112 215
rect 110 214 111 215
rect 109 214 110 215
rect 108 214 109 215
rect 107 214 108 215
rect 106 214 107 215
rect 105 214 106 215
rect 104 214 105 215
rect 103 214 104 215
rect 102 214 103 215
rect 64 214 65 215
rect 63 214 64 215
rect 62 214 63 215
rect 61 214 62 215
rect 60 214 61 215
rect 59 214 60 215
rect 29 214 30 215
rect 28 214 29 215
rect 27 214 28 215
rect 23 214 24 215
rect 22 214 23 215
rect 21 214 22 215
rect 20 214 21 215
rect 19 214 20 215
rect 18 214 19 215
rect 17 214 18 215
rect 16 214 17 215
rect 15 214 16 215
rect 179 215 180 216
rect 178 215 179 216
rect 177 215 178 216
rect 176 215 177 216
rect 173 215 174 216
rect 172 215 173 216
rect 171 215 172 216
rect 170 215 171 216
rect 165 215 166 216
rect 164 215 165 216
rect 163 215 164 216
rect 162 215 163 216
rect 149 215 150 216
rect 148 215 149 216
rect 147 215 148 216
rect 146 215 147 216
rect 145 215 146 216
rect 144 215 145 216
rect 143 215 144 216
rect 142 215 143 216
rect 141 215 142 216
rect 140 215 141 216
rect 130 215 131 216
rect 129 215 130 216
rect 128 215 129 216
rect 127 215 128 216
rect 126 215 127 216
rect 125 215 126 216
rect 124 215 125 216
rect 123 215 124 216
rect 122 215 123 216
rect 121 215 122 216
rect 112 215 113 216
rect 111 215 112 216
rect 110 215 111 216
rect 109 215 110 216
rect 108 215 109 216
rect 107 215 108 216
rect 106 215 107 216
rect 105 215 106 216
rect 104 215 105 216
rect 103 215 104 216
rect 102 215 103 216
rect 63 215 64 216
rect 62 215 63 216
rect 61 215 62 216
rect 60 215 61 216
rect 59 215 60 216
rect 29 215 30 216
rect 28 215 29 216
rect 27 215 28 216
rect 22 215 23 216
rect 21 215 22 216
rect 20 215 21 216
rect 19 215 20 216
rect 18 215 19 216
rect 17 215 18 216
rect 16 215 17 216
rect 15 215 16 216
rect 196 216 197 217
rect 195 216 196 217
rect 194 216 195 217
rect 193 216 194 217
rect 192 216 193 217
rect 191 216 192 217
rect 179 216 180 217
rect 178 216 179 217
rect 177 216 178 217
rect 176 216 177 217
rect 173 216 174 217
rect 172 216 173 217
rect 171 216 172 217
rect 170 216 171 217
rect 165 216 166 217
rect 164 216 165 217
rect 163 216 164 217
rect 162 216 163 217
rect 149 216 150 217
rect 148 216 149 217
rect 147 216 148 217
rect 146 216 147 217
rect 145 216 146 217
rect 144 216 145 217
rect 143 216 144 217
rect 142 216 143 217
rect 141 216 142 217
rect 140 216 141 217
rect 130 216 131 217
rect 129 216 130 217
rect 128 216 129 217
rect 127 216 128 217
rect 126 216 127 217
rect 125 216 126 217
rect 124 216 125 217
rect 123 216 124 217
rect 122 216 123 217
rect 121 216 122 217
rect 112 216 113 217
rect 111 216 112 217
rect 110 216 111 217
rect 109 216 110 217
rect 108 216 109 217
rect 107 216 108 217
rect 106 216 107 217
rect 105 216 106 217
rect 104 216 105 217
rect 103 216 104 217
rect 102 216 103 217
rect 63 216 64 217
rect 62 216 63 217
rect 61 216 62 217
rect 60 216 61 217
rect 59 216 60 217
rect 58 216 59 217
rect 21 216 22 217
rect 20 216 21 217
rect 19 216 20 217
rect 18 216 19 217
rect 17 216 18 217
rect 16 216 17 217
rect 197 217 198 218
rect 196 217 197 218
rect 195 217 196 218
rect 194 217 195 218
rect 193 217 194 218
rect 192 217 193 218
rect 191 217 192 218
rect 179 217 180 218
rect 178 217 179 218
rect 177 217 178 218
rect 176 217 177 218
rect 173 217 174 218
rect 172 217 173 218
rect 171 217 172 218
rect 170 217 171 218
rect 165 217 166 218
rect 164 217 165 218
rect 163 217 164 218
rect 162 217 163 218
rect 149 217 150 218
rect 148 217 149 218
rect 147 217 148 218
rect 146 217 147 218
rect 145 217 146 218
rect 144 217 145 218
rect 143 217 144 218
rect 142 217 143 218
rect 141 217 142 218
rect 140 217 141 218
rect 130 217 131 218
rect 129 217 130 218
rect 128 217 129 218
rect 127 217 128 218
rect 126 217 127 218
rect 125 217 126 218
rect 124 217 125 218
rect 123 217 124 218
rect 122 217 123 218
rect 121 217 122 218
rect 112 217 113 218
rect 111 217 112 218
rect 110 217 111 218
rect 109 217 110 218
rect 108 217 109 218
rect 107 217 108 218
rect 106 217 107 218
rect 105 217 106 218
rect 104 217 105 218
rect 103 217 104 218
rect 102 217 103 218
rect 63 217 64 218
rect 62 217 63 218
rect 61 217 62 218
rect 60 217 61 218
rect 59 217 60 218
rect 58 217 59 218
rect 19 217 20 218
rect 18 217 19 218
rect 192 218 193 219
rect 191 218 192 219
rect 179 218 180 219
rect 178 218 179 219
rect 177 218 178 219
rect 176 218 177 219
rect 173 218 174 219
rect 172 218 173 219
rect 171 218 172 219
rect 170 218 171 219
rect 165 218 166 219
rect 164 218 165 219
rect 163 218 164 219
rect 162 218 163 219
rect 149 218 150 219
rect 148 218 149 219
rect 147 218 148 219
rect 146 218 147 219
rect 145 218 146 219
rect 144 218 145 219
rect 143 218 144 219
rect 142 218 143 219
rect 141 218 142 219
rect 140 218 141 219
rect 130 218 131 219
rect 129 218 130 219
rect 128 218 129 219
rect 127 218 128 219
rect 126 218 127 219
rect 125 218 126 219
rect 124 218 125 219
rect 123 218 124 219
rect 122 218 123 219
rect 121 218 122 219
rect 112 218 113 219
rect 111 218 112 219
rect 110 218 111 219
rect 109 218 110 219
rect 108 218 109 219
rect 107 218 108 219
rect 106 218 107 219
rect 105 218 106 219
rect 104 218 105 219
rect 103 218 104 219
rect 102 218 103 219
rect 63 218 64 219
rect 62 218 63 219
rect 61 218 62 219
rect 60 218 61 219
rect 59 218 60 219
rect 26 218 27 219
rect 25 218 26 219
rect 24 218 25 219
rect 192 219 193 220
rect 191 219 192 220
rect 179 219 180 220
rect 178 219 179 220
rect 177 219 178 220
rect 176 219 177 220
rect 173 219 174 220
rect 172 219 173 220
rect 171 219 172 220
rect 170 219 171 220
rect 165 219 166 220
rect 164 219 165 220
rect 163 219 164 220
rect 162 219 163 220
rect 149 219 150 220
rect 148 219 149 220
rect 147 219 148 220
rect 146 219 147 220
rect 145 219 146 220
rect 144 219 145 220
rect 143 219 144 220
rect 142 219 143 220
rect 141 219 142 220
rect 140 219 141 220
rect 130 219 131 220
rect 129 219 130 220
rect 128 219 129 220
rect 127 219 128 220
rect 126 219 127 220
rect 125 219 126 220
rect 124 219 125 220
rect 123 219 124 220
rect 122 219 123 220
rect 121 219 122 220
rect 112 219 113 220
rect 111 219 112 220
rect 110 219 111 220
rect 109 219 110 220
rect 108 219 109 220
rect 107 219 108 220
rect 106 219 107 220
rect 105 219 106 220
rect 104 219 105 220
rect 103 219 104 220
rect 102 219 103 220
rect 85 219 86 220
rect 84 219 85 220
rect 83 219 84 220
rect 63 219 64 220
rect 62 219 63 220
rect 61 219 62 220
rect 60 219 61 220
rect 59 219 60 220
rect 26 219 27 220
rect 25 219 26 220
rect 24 219 25 220
rect 23 219 24 220
rect 196 220 197 221
rect 195 220 196 221
rect 194 220 195 221
rect 193 220 194 221
rect 192 220 193 221
rect 191 220 192 221
rect 179 220 180 221
rect 178 220 179 221
rect 177 220 178 221
rect 176 220 177 221
rect 173 220 174 221
rect 172 220 173 221
rect 171 220 172 221
rect 170 220 171 221
rect 165 220 166 221
rect 164 220 165 221
rect 163 220 164 221
rect 162 220 163 221
rect 149 220 150 221
rect 148 220 149 221
rect 147 220 148 221
rect 146 220 147 221
rect 145 220 146 221
rect 144 220 145 221
rect 143 220 144 221
rect 142 220 143 221
rect 141 220 142 221
rect 140 220 141 221
rect 130 220 131 221
rect 129 220 130 221
rect 128 220 129 221
rect 127 220 128 221
rect 126 220 127 221
rect 125 220 126 221
rect 124 220 125 221
rect 123 220 124 221
rect 122 220 123 221
rect 121 220 122 221
rect 112 220 113 221
rect 111 220 112 221
rect 110 220 111 221
rect 109 220 110 221
rect 108 220 109 221
rect 107 220 108 221
rect 106 220 107 221
rect 105 220 106 221
rect 104 220 105 221
rect 103 220 104 221
rect 102 220 103 221
rect 86 220 87 221
rect 85 220 86 221
rect 84 220 85 221
rect 83 220 84 221
rect 60 220 61 221
rect 59 220 60 221
rect 26 220 27 221
rect 25 220 26 221
rect 24 220 25 221
rect 23 220 24 221
rect 22 220 23 221
rect 197 221 198 222
rect 196 221 197 222
rect 195 221 196 222
rect 194 221 195 222
rect 193 221 194 222
rect 192 221 193 222
rect 191 221 192 222
rect 179 221 180 222
rect 178 221 179 222
rect 177 221 178 222
rect 176 221 177 222
rect 173 221 174 222
rect 172 221 173 222
rect 171 221 172 222
rect 170 221 171 222
rect 165 221 166 222
rect 164 221 165 222
rect 163 221 164 222
rect 162 221 163 222
rect 149 221 150 222
rect 148 221 149 222
rect 147 221 148 222
rect 146 221 147 222
rect 145 221 146 222
rect 144 221 145 222
rect 143 221 144 222
rect 142 221 143 222
rect 141 221 142 222
rect 140 221 141 222
rect 130 221 131 222
rect 129 221 130 222
rect 128 221 129 222
rect 127 221 128 222
rect 126 221 127 222
rect 125 221 126 222
rect 124 221 125 222
rect 123 221 124 222
rect 122 221 123 222
rect 121 221 122 222
rect 112 221 113 222
rect 111 221 112 222
rect 110 221 111 222
rect 109 221 110 222
rect 108 221 109 222
rect 107 221 108 222
rect 106 221 107 222
rect 105 221 106 222
rect 104 221 105 222
rect 103 221 104 222
rect 102 221 103 222
rect 86 221 87 222
rect 85 221 86 222
rect 84 221 85 222
rect 83 221 84 222
rect 26 221 27 222
rect 25 221 26 222
rect 24 221 25 222
rect 23 221 24 222
rect 22 221 23 222
rect 21 221 22 222
rect 179 222 180 223
rect 178 222 179 223
rect 177 222 178 223
rect 176 222 177 223
rect 175 222 176 223
rect 174 222 175 223
rect 173 222 174 223
rect 172 222 173 223
rect 171 222 172 223
rect 170 222 171 223
rect 165 222 166 223
rect 164 222 165 223
rect 163 222 164 223
rect 162 222 163 223
rect 149 222 150 223
rect 148 222 149 223
rect 147 222 148 223
rect 146 222 147 223
rect 145 222 146 223
rect 144 222 145 223
rect 143 222 144 223
rect 142 222 143 223
rect 141 222 142 223
rect 140 222 141 223
rect 130 222 131 223
rect 129 222 130 223
rect 128 222 129 223
rect 127 222 128 223
rect 126 222 127 223
rect 125 222 126 223
rect 124 222 125 223
rect 123 222 124 223
rect 122 222 123 223
rect 121 222 122 223
rect 112 222 113 223
rect 111 222 112 223
rect 110 222 111 223
rect 109 222 110 223
rect 108 222 109 223
rect 107 222 108 223
rect 106 222 107 223
rect 105 222 106 223
rect 104 222 105 223
rect 103 222 104 223
rect 102 222 103 223
rect 86 222 87 223
rect 85 222 86 223
rect 84 222 85 223
rect 83 222 84 223
rect 26 222 27 223
rect 25 222 26 223
rect 24 222 25 223
rect 22 222 23 223
rect 21 222 22 223
rect 20 222 21 223
rect 196 223 197 224
rect 195 223 196 224
rect 194 223 195 224
rect 193 223 194 224
rect 192 223 193 224
rect 191 223 192 224
rect 189 223 190 224
rect 188 223 189 224
rect 179 223 180 224
rect 178 223 179 224
rect 177 223 178 224
rect 176 223 177 224
rect 175 223 176 224
rect 174 223 175 224
rect 173 223 174 224
rect 172 223 173 224
rect 171 223 172 224
rect 170 223 171 224
rect 165 223 166 224
rect 164 223 165 224
rect 163 223 164 224
rect 162 223 163 224
rect 149 223 150 224
rect 148 223 149 224
rect 147 223 148 224
rect 146 223 147 224
rect 145 223 146 224
rect 144 223 145 224
rect 143 223 144 224
rect 142 223 143 224
rect 141 223 142 224
rect 140 223 141 224
rect 130 223 131 224
rect 129 223 130 224
rect 128 223 129 224
rect 127 223 128 224
rect 126 223 127 224
rect 125 223 126 224
rect 124 223 125 224
rect 123 223 124 224
rect 122 223 123 224
rect 121 223 122 224
rect 112 223 113 224
rect 111 223 112 224
rect 110 223 111 224
rect 109 223 110 224
rect 108 223 109 224
rect 107 223 108 224
rect 106 223 107 224
rect 105 223 106 224
rect 104 223 105 224
rect 103 223 104 224
rect 102 223 103 224
rect 86 223 87 224
rect 85 223 86 224
rect 84 223 85 224
rect 83 223 84 224
rect 29 223 30 224
rect 28 223 29 224
rect 26 223 27 224
rect 25 223 26 224
rect 24 223 25 224
rect 21 223 22 224
rect 20 223 21 224
rect 19 223 20 224
rect 18 223 19 224
rect 196 224 197 225
rect 195 224 196 225
rect 194 224 195 225
rect 193 224 194 225
rect 192 224 193 225
rect 191 224 192 225
rect 189 224 190 225
rect 188 224 189 225
rect 179 224 180 225
rect 178 224 179 225
rect 177 224 178 225
rect 176 224 177 225
rect 175 224 176 225
rect 174 224 175 225
rect 173 224 174 225
rect 172 224 173 225
rect 171 224 172 225
rect 170 224 171 225
rect 165 224 166 225
rect 164 224 165 225
rect 163 224 164 225
rect 162 224 163 225
rect 149 224 150 225
rect 148 224 149 225
rect 147 224 148 225
rect 146 224 147 225
rect 145 224 146 225
rect 144 224 145 225
rect 143 224 144 225
rect 142 224 143 225
rect 141 224 142 225
rect 140 224 141 225
rect 130 224 131 225
rect 129 224 130 225
rect 128 224 129 225
rect 127 224 128 225
rect 126 224 127 225
rect 125 224 126 225
rect 124 224 125 225
rect 123 224 124 225
rect 122 224 123 225
rect 121 224 122 225
rect 112 224 113 225
rect 111 224 112 225
rect 110 224 111 225
rect 109 224 110 225
rect 108 224 109 225
rect 107 224 108 225
rect 106 224 107 225
rect 105 224 106 225
rect 104 224 105 225
rect 103 224 104 225
rect 102 224 103 225
rect 86 224 87 225
rect 85 224 86 225
rect 84 224 85 225
rect 83 224 84 225
rect 29 224 30 225
rect 28 224 29 225
rect 27 224 28 225
rect 26 224 27 225
rect 25 224 26 225
rect 24 224 25 225
rect 23 224 24 225
rect 20 224 21 225
rect 19 224 20 225
rect 18 224 19 225
rect 17 224 18 225
rect 179 225 180 226
rect 178 225 179 226
rect 177 225 178 226
rect 176 225 177 226
rect 173 225 174 226
rect 172 225 173 226
rect 171 225 172 226
rect 170 225 171 226
rect 165 225 166 226
rect 164 225 165 226
rect 163 225 164 226
rect 162 225 163 226
rect 149 225 150 226
rect 148 225 149 226
rect 147 225 148 226
rect 146 225 147 226
rect 145 225 146 226
rect 144 225 145 226
rect 143 225 144 226
rect 142 225 143 226
rect 141 225 142 226
rect 140 225 141 226
rect 130 225 131 226
rect 129 225 130 226
rect 128 225 129 226
rect 127 225 128 226
rect 126 225 127 226
rect 125 225 126 226
rect 124 225 125 226
rect 123 225 124 226
rect 122 225 123 226
rect 121 225 122 226
rect 112 225 113 226
rect 111 225 112 226
rect 110 225 111 226
rect 109 225 110 226
rect 108 225 109 226
rect 107 225 108 226
rect 106 225 107 226
rect 105 225 106 226
rect 104 225 105 226
rect 103 225 104 226
rect 102 225 103 226
rect 86 225 87 226
rect 85 225 86 226
rect 84 225 85 226
rect 83 225 84 226
rect 29 225 30 226
rect 28 225 29 226
rect 27 225 28 226
rect 26 225 27 226
rect 25 225 26 226
rect 24 225 25 226
rect 23 225 24 226
rect 22 225 23 226
rect 21 225 22 226
rect 20 225 21 226
rect 19 225 20 226
rect 18 225 19 226
rect 17 225 18 226
rect 16 225 17 226
rect 195 226 196 227
rect 194 226 195 227
rect 193 226 194 227
rect 192 226 193 227
rect 179 226 180 227
rect 178 226 179 227
rect 177 226 178 227
rect 176 226 177 227
rect 173 226 174 227
rect 172 226 173 227
rect 171 226 172 227
rect 170 226 171 227
rect 165 226 166 227
rect 164 226 165 227
rect 163 226 164 227
rect 162 226 163 227
rect 149 226 150 227
rect 148 226 149 227
rect 147 226 148 227
rect 146 226 147 227
rect 145 226 146 227
rect 144 226 145 227
rect 143 226 144 227
rect 142 226 143 227
rect 141 226 142 227
rect 140 226 141 227
rect 130 226 131 227
rect 129 226 130 227
rect 128 226 129 227
rect 127 226 128 227
rect 126 226 127 227
rect 125 226 126 227
rect 124 226 125 227
rect 123 226 124 227
rect 122 226 123 227
rect 121 226 122 227
rect 112 226 113 227
rect 111 226 112 227
rect 110 226 111 227
rect 109 226 110 227
rect 108 226 109 227
rect 107 226 108 227
rect 106 226 107 227
rect 105 226 106 227
rect 104 226 105 227
rect 103 226 104 227
rect 102 226 103 227
rect 86 226 87 227
rect 85 226 86 227
rect 84 226 85 227
rect 83 226 84 227
rect 27 226 28 227
rect 26 226 27 227
rect 25 226 26 227
rect 24 226 25 227
rect 23 226 24 227
rect 22 226 23 227
rect 21 226 22 227
rect 20 226 21 227
rect 19 226 20 227
rect 18 226 19 227
rect 17 226 18 227
rect 16 226 17 227
rect 15 226 16 227
rect 196 227 197 228
rect 195 227 196 228
rect 194 227 195 228
rect 193 227 194 228
rect 192 227 193 228
rect 191 227 192 228
rect 179 227 180 228
rect 178 227 179 228
rect 177 227 178 228
rect 176 227 177 228
rect 173 227 174 228
rect 172 227 173 228
rect 171 227 172 228
rect 170 227 171 228
rect 165 227 166 228
rect 164 227 165 228
rect 163 227 164 228
rect 162 227 163 228
rect 149 227 150 228
rect 148 227 149 228
rect 147 227 148 228
rect 146 227 147 228
rect 145 227 146 228
rect 144 227 145 228
rect 143 227 144 228
rect 142 227 143 228
rect 141 227 142 228
rect 140 227 141 228
rect 130 227 131 228
rect 129 227 130 228
rect 128 227 129 228
rect 127 227 128 228
rect 126 227 127 228
rect 125 227 126 228
rect 124 227 125 228
rect 123 227 124 228
rect 122 227 123 228
rect 121 227 122 228
rect 112 227 113 228
rect 111 227 112 228
rect 110 227 111 228
rect 109 227 110 228
rect 108 227 109 228
rect 107 227 108 228
rect 106 227 107 228
rect 105 227 106 228
rect 104 227 105 228
rect 103 227 104 228
rect 102 227 103 228
rect 86 227 87 228
rect 85 227 86 228
rect 84 227 85 228
rect 83 227 84 228
rect 26 227 27 228
rect 25 227 26 228
rect 24 227 25 228
rect 22 227 23 228
rect 21 227 22 228
rect 20 227 21 228
rect 19 227 20 228
rect 18 227 19 228
rect 17 227 18 228
rect 16 227 17 228
rect 15 227 16 228
rect 196 228 197 229
rect 195 228 196 229
rect 192 228 193 229
rect 191 228 192 229
rect 179 228 180 229
rect 178 228 179 229
rect 177 228 178 229
rect 176 228 177 229
rect 173 228 174 229
rect 172 228 173 229
rect 171 228 172 229
rect 170 228 171 229
rect 165 228 166 229
rect 164 228 165 229
rect 163 228 164 229
rect 162 228 163 229
rect 149 228 150 229
rect 148 228 149 229
rect 147 228 148 229
rect 146 228 147 229
rect 145 228 146 229
rect 144 228 145 229
rect 143 228 144 229
rect 142 228 143 229
rect 141 228 142 229
rect 140 228 141 229
rect 130 228 131 229
rect 129 228 130 229
rect 128 228 129 229
rect 127 228 128 229
rect 126 228 127 229
rect 125 228 126 229
rect 124 228 125 229
rect 123 228 124 229
rect 122 228 123 229
rect 121 228 122 229
rect 112 228 113 229
rect 111 228 112 229
rect 110 228 111 229
rect 109 228 110 229
rect 108 228 109 229
rect 107 228 108 229
rect 106 228 107 229
rect 105 228 106 229
rect 104 228 105 229
rect 103 228 104 229
rect 102 228 103 229
rect 86 228 87 229
rect 85 228 86 229
rect 84 228 85 229
rect 83 228 84 229
rect 25 228 26 229
rect 24 228 25 229
rect 18 228 19 229
rect 17 228 18 229
rect 16 228 17 229
rect 15 228 16 229
rect 197 229 198 230
rect 196 229 197 230
rect 192 229 193 230
rect 191 229 192 230
rect 183 229 184 230
rect 182 229 183 230
rect 181 229 182 230
rect 180 229 181 230
rect 179 229 180 230
rect 178 229 179 230
rect 177 229 178 230
rect 176 229 177 230
rect 173 229 174 230
rect 172 229 173 230
rect 171 229 172 230
rect 170 229 171 230
rect 169 229 170 230
rect 168 229 169 230
rect 167 229 168 230
rect 166 229 167 230
rect 165 229 166 230
rect 164 229 165 230
rect 163 229 164 230
rect 162 229 163 230
rect 149 229 150 230
rect 148 229 149 230
rect 147 229 148 230
rect 146 229 147 230
rect 145 229 146 230
rect 144 229 145 230
rect 143 229 144 230
rect 142 229 143 230
rect 141 229 142 230
rect 140 229 141 230
rect 130 229 131 230
rect 129 229 130 230
rect 128 229 129 230
rect 127 229 128 230
rect 126 229 127 230
rect 125 229 126 230
rect 124 229 125 230
rect 123 229 124 230
rect 122 229 123 230
rect 121 229 122 230
rect 112 229 113 230
rect 111 229 112 230
rect 110 229 111 230
rect 109 229 110 230
rect 108 229 109 230
rect 107 229 108 230
rect 106 229 107 230
rect 105 229 106 230
rect 104 229 105 230
rect 103 229 104 230
rect 102 229 103 230
rect 86 229 87 230
rect 85 229 86 230
rect 84 229 85 230
rect 83 229 84 230
rect 196 230 197 231
rect 191 230 192 231
rect 183 230 184 231
rect 182 230 183 231
rect 181 230 182 231
rect 180 230 181 231
rect 179 230 180 231
rect 178 230 179 231
rect 177 230 178 231
rect 176 230 177 231
rect 173 230 174 231
rect 172 230 173 231
rect 171 230 172 231
rect 170 230 171 231
rect 169 230 170 231
rect 168 230 169 231
rect 167 230 168 231
rect 166 230 167 231
rect 165 230 166 231
rect 164 230 165 231
rect 163 230 164 231
rect 162 230 163 231
rect 149 230 150 231
rect 148 230 149 231
rect 147 230 148 231
rect 146 230 147 231
rect 145 230 146 231
rect 144 230 145 231
rect 143 230 144 231
rect 142 230 143 231
rect 141 230 142 231
rect 140 230 141 231
rect 130 230 131 231
rect 129 230 130 231
rect 128 230 129 231
rect 127 230 128 231
rect 126 230 127 231
rect 125 230 126 231
rect 124 230 125 231
rect 123 230 124 231
rect 122 230 123 231
rect 121 230 122 231
rect 112 230 113 231
rect 111 230 112 231
rect 110 230 111 231
rect 109 230 110 231
rect 108 230 109 231
rect 107 230 108 231
rect 106 230 107 231
rect 105 230 106 231
rect 104 230 105 231
rect 103 230 104 231
rect 102 230 103 231
rect 86 230 87 231
rect 85 230 86 231
rect 84 230 85 231
rect 83 230 84 231
rect 25 230 26 231
rect 24 230 25 231
rect 23 230 24 231
rect 196 231 197 232
rect 193 231 194 232
rect 192 231 193 232
rect 183 231 184 232
rect 182 231 183 232
rect 181 231 182 232
rect 180 231 181 232
rect 179 231 180 232
rect 178 231 179 232
rect 177 231 178 232
rect 176 231 177 232
rect 173 231 174 232
rect 172 231 173 232
rect 171 231 172 232
rect 170 231 171 232
rect 169 231 170 232
rect 168 231 169 232
rect 167 231 168 232
rect 166 231 167 232
rect 165 231 166 232
rect 164 231 165 232
rect 163 231 164 232
rect 162 231 163 232
rect 149 231 150 232
rect 148 231 149 232
rect 147 231 148 232
rect 146 231 147 232
rect 145 231 146 232
rect 144 231 145 232
rect 143 231 144 232
rect 142 231 143 232
rect 141 231 142 232
rect 140 231 141 232
rect 130 231 131 232
rect 129 231 130 232
rect 128 231 129 232
rect 127 231 128 232
rect 126 231 127 232
rect 125 231 126 232
rect 124 231 125 232
rect 123 231 124 232
rect 122 231 123 232
rect 121 231 122 232
rect 112 231 113 232
rect 111 231 112 232
rect 110 231 111 232
rect 109 231 110 232
rect 108 231 109 232
rect 107 231 108 232
rect 106 231 107 232
rect 105 231 106 232
rect 104 231 105 232
rect 103 231 104 232
rect 102 231 103 232
rect 86 231 87 232
rect 85 231 86 232
rect 84 231 85 232
rect 83 231 84 232
rect 25 231 26 232
rect 24 231 25 232
rect 23 231 24 232
rect 197 232 198 233
rect 196 232 197 233
rect 194 232 195 233
rect 193 232 194 233
rect 192 232 193 233
rect 191 232 192 233
rect 183 232 184 233
rect 182 232 183 233
rect 181 232 182 233
rect 180 232 181 233
rect 179 232 180 233
rect 178 232 179 233
rect 177 232 178 233
rect 176 232 177 233
rect 173 232 174 233
rect 172 232 173 233
rect 171 232 172 233
rect 170 232 171 233
rect 169 232 170 233
rect 168 232 169 233
rect 167 232 168 233
rect 166 232 167 233
rect 165 232 166 233
rect 164 232 165 233
rect 163 232 164 233
rect 162 232 163 233
rect 149 232 150 233
rect 148 232 149 233
rect 147 232 148 233
rect 146 232 147 233
rect 145 232 146 233
rect 144 232 145 233
rect 143 232 144 233
rect 142 232 143 233
rect 141 232 142 233
rect 140 232 141 233
rect 130 232 131 233
rect 129 232 130 233
rect 128 232 129 233
rect 127 232 128 233
rect 126 232 127 233
rect 125 232 126 233
rect 124 232 125 233
rect 123 232 124 233
rect 122 232 123 233
rect 121 232 122 233
rect 112 232 113 233
rect 111 232 112 233
rect 110 232 111 233
rect 109 232 110 233
rect 108 232 109 233
rect 107 232 108 233
rect 106 232 107 233
rect 105 232 106 233
rect 104 232 105 233
rect 103 232 104 233
rect 102 232 103 233
rect 86 232 87 233
rect 85 232 86 233
rect 84 232 85 233
rect 83 232 84 233
rect 25 232 26 233
rect 24 232 25 233
rect 23 232 24 233
rect 197 233 198 234
rect 196 233 197 234
rect 194 233 195 234
rect 193 233 194 234
rect 192 233 193 234
rect 191 233 192 234
rect 173 233 174 234
rect 172 233 173 234
rect 171 233 172 234
rect 170 233 171 234
rect 164 233 165 234
rect 163 233 164 234
rect 149 233 150 234
rect 148 233 149 234
rect 147 233 148 234
rect 146 233 147 234
rect 145 233 146 234
rect 144 233 145 234
rect 143 233 144 234
rect 142 233 143 234
rect 141 233 142 234
rect 140 233 141 234
rect 130 233 131 234
rect 129 233 130 234
rect 128 233 129 234
rect 127 233 128 234
rect 126 233 127 234
rect 125 233 126 234
rect 124 233 125 234
rect 123 233 124 234
rect 122 233 123 234
rect 121 233 122 234
rect 112 233 113 234
rect 111 233 112 234
rect 110 233 111 234
rect 109 233 110 234
rect 108 233 109 234
rect 107 233 108 234
rect 106 233 107 234
rect 105 233 106 234
rect 104 233 105 234
rect 103 233 104 234
rect 102 233 103 234
rect 86 233 87 234
rect 85 233 86 234
rect 84 233 85 234
rect 83 233 84 234
rect 25 233 26 234
rect 24 233 25 234
rect 23 233 24 234
rect 197 234 198 235
rect 196 234 197 235
rect 195 234 196 235
rect 194 234 195 235
rect 192 234 193 235
rect 191 234 192 235
rect 173 234 174 235
rect 172 234 173 235
rect 171 234 172 235
rect 170 234 171 235
rect 149 234 150 235
rect 148 234 149 235
rect 147 234 148 235
rect 146 234 147 235
rect 145 234 146 235
rect 144 234 145 235
rect 143 234 144 235
rect 142 234 143 235
rect 141 234 142 235
rect 140 234 141 235
rect 130 234 131 235
rect 129 234 130 235
rect 128 234 129 235
rect 127 234 128 235
rect 126 234 127 235
rect 125 234 126 235
rect 124 234 125 235
rect 123 234 124 235
rect 122 234 123 235
rect 121 234 122 235
rect 112 234 113 235
rect 111 234 112 235
rect 110 234 111 235
rect 109 234 110 235
rect 108 234 109 235
rect 107 234 108 235
rect 106 234 107 235
rect 105 234 106 235
rect 104 234 105 235
rect 103 234 104 235
rect 102 234 103 235
rect 86 234 87 235
rect 85 234 86 235
rect 84 234 85 235
rect 83 234 84 235
rect 25 234 26 235
rect 24 234 25 235
rect 23 234 24 235
rect 196 235 197 236
rect 195 235 196 236
rect 194 235 195 236
rect 192 235 193 236
rect 191 235 192 236
rect 173 235 174 236
rect 172 235 173 236
rect 171 235 172 236
rect 170 235 171 236
rect 149 235 150 236
rect 148 235 149 236
rect 147 235 148 236
rect 146 235 147 236
rect 145 235 146 236
rect 144 235 145 236
rect 143 235 144 236
rect 142 235 143 236
rect 141 235 142 236
rect 140 235 141 236
rect 130 235 131 236
rect 129 235 130 236
rect 128 235 129 236
rect 127 235 128 236
rect 126 235 127 236
rect 125 235 126 236
rect 124 235 125 236
rect 123 235 124 236
rect 122 235 123 236
rect 121 235 122 236
rect 112 235 113 236
rect 111 235 112 236
rect 110 235 111 236
rect 109 235 110 236
rect 108 235 109 236
rect 107 235 108 236
rect 106 235 107 236
rect 105 235 106 236
rect 104 235 105 236
rect 103 235 104 236
rect 102 235 103 236
rect 86 235 87 236
rect 85 235 86 236
rect 84 235 85 236
rect 83 235 84 236
rect 25 235 26 236
rect 24 235 25 236
rect 23 235 24 236
rect 172 236 173 237
rect 171 236 172 237
rect 149 236 150 237
rect 148 236 149 237
rect 147 236 148 237
rect 146 236 147 237
rect 145 236 146 237
rect 144 236 145 237
rect 143 236 144 237
rect 142 236 143 237
rect 141 236 142 237
rect 140 236 141 237
rect 130 236 131 237
rect 129 236 130 237
rect 128 236 129 237
rect 127 236 128 237
rect 126 236 127 237
rect 125 236 126 237
rect 124 236 125 237
rect 123 236 124 237
rect 122 236 123 237
rect 121 236 122 237
rect 112 236 113 237
rect 111 236 112 237
rect 110 236 111 237
rect 109 236 110 237
rect 108 236 109 237
rect 107 236 108 237
rect 106 236 107 237
rect 105 236 106 237
rect 104 236 105 237
rect 103 236 104 237
rect 102 236 103 237
rect 86 236 87 237
rect 85 236 86 237
rect 84 236 85 237
rect 83 236 84 237
rect 149 237 150 238
rect 148 237 149 238
rect 147 237 148 238
rect 146 237 147 238
rect 145 237 146 238
rect 144 237 145 238
rect 143 237 144 238
rect 142 237 143 238
rect 141 237 142 238
rect 140 237 141 238
rect 130 237 131 238
rect 129 237 130 238
rect 128 237 129 238
rect 127 237 128 238
rect 126 237 127 238
rect 125 237 126 238
rect 124 237 125 238
rect 123 237 124 238
rect 122 237 123 238
rect 121 237 122 238
rect 112 237 113 238
rect 111 237 112 238
rect 110 237 111 238
rect 109 237 110 238
rect 108 237 109 238
rect 107 237 108 238
rect 106 237 107 238
rect 105 237 106 238
rect 104 237 105 238
rect 103 237 104 238
rect 102 237 103 238
rect 86 237 87 238
rect 85 237 86 238
rect 84 237 85 238
rect 83 237 84 238
rect 26 237 27 238
rect 25 237 26 238
rect 149 238 150 239
rect 148 238 149 239
rect 147 238 148 239
rect 146 238 147 239
rect 145 238 146 239
rect 144 238 145 239
rect 143 238 144 239
rect 142 238 143 239
rect 141 238 142 239
rect 140 238 141 239
rect 130 238 131 239
rect 129 238 130 239
rect 128 238 129 239
rect 127 238 128 239
rect 126 238 127 239
rect 125 238 126 239
rect 124 238 125 239
rect 123 238 124 239
rect 122 238 123 239
rect 121 238 122 239
rect 112 238 113 239
rect 111 238 112 239
rect 110 238 111 239
rect 109 238 110 239
rect 108 238 109 239
rect 107 238 108 239
rect 106 238 107 239
rect 105 238 106 239
rect 104 238 105 239
rect 103 238 104 239
rect 102 238 103 239
rect 86 238 87 239
rect 85 238 86 239
rect 84 238 85 239
rect 83 238 84 239
rect 28 238 29 239
rect 27 238 28 239
rect 26 238 27 239
rect 25 238 26 239
rect 149 239 150 240
rect 148 239 149 240
rect 147 239 148 240
rect 146 239 147 240
rect 145 239 146 240
rect 144 239 145 240
rect 143 239 144 240
rect 142 239 143 240
rect 141 239 142 240
rect 140 239 141 240
rect 130 239 131 240
rect 129 239 130 240
rect 128 239 129 240
rect 127 239 128 240
rect 126 239 127 240
rect 125 239 126 240
rect 124 239 125 240
rect 123 239 124 240
rect 122 239 123 240
rect 121 239 122 240
rect 112 239 113 240
rect 111 239 112 240
rect 110 239 111 240
rect 109 239 110 240
rect 108 239 109 240
rect 107 239 108 240
rect 106 239 107 240
rect 105 239 106 240
rect 104 239 105 240
rect 103 239 104 240
rect 102 239 103 240
rect 86 239 87 240
rect 85 239 86 240
rect 84 239 85 240
rect 83 239 84 240
rect 28 239 29 240
rect 27 239 28 240
rect 26 239 27 240
rect 25 239 26 240
rect 19 239 20 240
rect 18 239 19 240
rect 17 239 18 240
rect 196 240 197 241
rect 195 240 196 241
rect 194 240 195 241
rect 192 240 193 241
rect 191 240 192 241
rect 149 240 150 241
rect 148 240 149 241
rect 147 240 148 241
rect 146 240 147 241
rect 145 240 146 241
rect 144 240 145 241
rect 143 240 144 241
rect 142 240 143 241
rect 141 240 142 241
rect 140 240 141 241
rect 130 240 131 241
rect 129 240 130 241
rect 128 240 129 241
rect 127 240 128 241
rect 126 240 127 241
rect 125 240 126 241
rect 124 240 125 241
rect 123 240 124 241
rect 122 240 123 241
rect 121 240 122 241
rect 112 240 113 241
rect 111 240 112 241
rect 110 240 111 241
rect 109 240 110 241
rect 108 240 109 241
rect 107 240 108 241
rect 106 240 107 241
rect 105 240 106 241
rect 104 240 105 241
rect 103 240 104 241
rect 102 240 103 241
rect 86 240 87 241
rect 85 240 86 241
rect 84 240 85 241
rect 83 240 84 241
rect 29 240 30 241
rect 28 240 29 241
rect 27 240 28 241
rect 26 240 27 241
rect 19 240 20 241
rect 18 240 19 241
rect 17 240 18 241
rect 16 240 17 241
rect 196 241 197 242
rect 195 241 196 242
rect 194 241 195 242
rect 193 241 194 242
rect 192 241 193 242
rect 191 241 192 242
rect 149 241 150 242
rect 148 241 149 242
rect 147 241 148 242
rect 146 241 147 242
rect 145 241 146 242
rect 144 241 145 242
rect 143 241 144 242
rect 142 241 143 242
rect 141 241 142 242
rect 140 241 141 242
rect 130 241 131 242
rect 129 241 130 242
rect 128 241 129 242
rect 127 241 128 242
rect 126 241 127 242
rect 125 241 126 242
rect 124 241 125 242
rect 123 241 124 242
rect 122 241 123 242
rect 121 241 122 242
rect 112 241 113 242
rect 111 241 112 242
rect 110 241 111 242
rect 109 241 110 242
rect 108 241 109 242
rect 107 241 108 242
rect 106 241 107 242
rect 105 241 106 242
rect 104 241 105 242
rect 103 241 104 242
rect 102 241 103 242
rect 85 241 86 242
rect 84 241 85 242
rect 83 241 84 242
rect 29 241 30 242
rect 28 241 29 242
rect 27 241 28 242
rect 19 241 20 242
rect 18 241 19 242
rect 17 241 18 242
rect 16 241 17 242
rect 15 241 16 242
rect 197 242 198 243
rect 196 242 197 243
rect 194 242 195 243
rect 193 242 194 243
rect 192 242 193 243
rect 191 242 192 243
rect 149 242 150 243
rect 148 242 149 243
rect 147 242 148 243
rect 146 242 147 243
rect 145 242 146 243
rect 144 242 145 243
rect 143 242 144 243
rect 142 242 143 243
rect 141 242 142 243
rect 140 242 141 243
rect 130 242 131 243
rect 129 242 130 243
rect 128 242 129 243
rect 127 242 128 243
rect 126 242 127 243
rect 125 242 126 243
rect 124 242 125 243
rect 123 242 124 243
rect 122 242 123 243
rect 121 242 122 243
rect 112 242 113 243
rect 111 242 112 243
rect 110 242 111 243
rect 109 242 110 243
rect 108 242 109 243
rect 107 242 108 243
rect 106 242 107 243
rect 105 242 106 243
rect 104 242 105 243
rect 103 242 104 243
rect 102 242 103 243
rect 29 242 30 243
rect 28 242 29 243
rect 27 242 28 243
rect 22 242 23 243
rect 21 242 22 243
rect 17 242 18 243
rect 16 242 17 243
rect 15 242 16 243
rect 196 243 197 244
rect 195 243 196 244
rect 194 243 195 244
rect 193 243 194 244
rect 192 243 193 244
rect 191 243 192 244
rect 149 243 150 244
rect 148 243 149 244
rect 147 243 148 244
rect 146 243 147 244
rect 145 243 146 244
rect 144 243 145 244
rect 143 243 144 244
rect 142 243 143 244
rect 141 243 142 244
rect 140 243 141 244
rect 130 243 131 244
rect 129 243 130 244
rect 128 243 129 244
rect 127 243 128 244
rect 126 243 127 244
rect 125 243 126 244
rect 124 243 125 244
rect 123 243 124 244
rect 122 243 123 244
rect 121 243 122 244
rect 112 243 113 244
rect 111 243 112 244
rect 110 243 111 244
rect 109 243 110 244
rect 108 243 109 244
rect 107 243 108 244
rect 106 243 107 244
rect 105 243 106 244
rect 104 243 105 244
rect 103 243 104 244
rect 102 243 103 244
rect 29 243 30 244
rect 28 243 29 244
rect 27 243 28 244
rect 23 243 24 244
rect 22 243 23 244
rect 21 243 22 244
rect 20 243 21 244
rect 17 243 18 244
rect 16 243 17 244
rect 15 243 16 244
rect 197 244 198 245
rect 196 244 197 245
rect 195 244 196 245
rect 194 244 195 245
rect 193 244 194 245
rect 192 244 193 245
rect 191 244 192 245
rect 149 244 150 245
rect 148 244 149 245
rect 147 244 148 245
rect 146 244 147 245
rect 145 244 146 245
rect 144 244 145 245
rect 143 244 144 245
rect 142 244 143 245
rect 141 244 142 245
rect 140 244 141 245
rect 130 244 131 245
rect 129 244 130 245
rect 128 244 129 245
rect 127 244 128 245
rect 126 244 127 245
rect 125 244 126 245
rect 124 244 125 245
rect 123 244 124 245
rect 122 244 123 245
rect 121 244 122 245
rect 112 244 113 245
rect 111 244 112 245
rect 110 244 111 245
rect 109 244 110 245
rect 108 244 109 245
rect 107 244 108 245
rect 106 244 107 245
rect 105 244 106 245
rect 104 244 105 245
rect 103 244 104 245
rect 102 244 103 245
rect 86 244 87 245
rect 85 244 86 245
rect 84 244 85 245
rect 83 244 84 245
rect 82 244 83 245
rect 81 244 82 245
rect 80 244 81 245
rect 79 244 80 245
rect 78 244 79 245
rect 77 244 78 245
rect 76 244 77 245
rect 75 244 76 245
rect 74 244 75 245
rect 73 244 74 245
rect 72 244 73 245
rect 71 244 72 245
rect 70 244 71 245
rect 69 244 70 245
rect 68 244 69 245
rect 67 244 68 245
rect 66 244 67 245
rect 65 244 66 245
rect 64 244 65 245
rect 63 244 64 245
rect 62 244 63 245
rect 61 244 62 245
rect 60 244 61 245
rect 59 244 60 245
rect 28 244 29 245
rect 27 244 28 245
rect 26 244 27 245
rect 25 244 26 245
rect 24 244 25 245
rect 23 244 24 245
rect 22 244 23 245
rect 21 244 22 245
rect 20 244 21 245
rect 17 244 18 245
rect 16 244 17 245
rect 15 244 16 245
rect 196 245 197 246
rect 195 245 196 246
rect 194 245 195 246
rect 193 245 194 246
rect 192 245 193 246
rect 149 245 150 246
rect 148 245 149 246
rect 147 245 148 246
rect 146 245 147 246
rect 145 245 146 246
rect 144 245 145 246
rect 143 245 144 246
rect 142 245 143 246
rect 141 245 142 246
rect 140 245 141 246
rect 130 245 131 246
rect 129 245 130 246
rect 128 245 129 246
rect 127 245 128 246
rect 126 245 127 246
rect 125 245 126 246
rect 124 245 125 246
rect 123 245 124 246
rect 122 245 123 246
rect 121 245 122 246
rect 112 245 113 246
rect 111 245 112 246
rect 110 245 111 246
rect 109 245 110 246
rect 108 245 109 246
rect 107 245 108 246
rect 106 245 107 246
rect 105 245 106 246
rect 104 245 105 246
rect 103 245 104 246
rect 102 245 103 246
rect 86 245 87 246
rect 85 245 86 246
rect 84 245 85 246
rect 83 245 84 246
rect 82 245 83 246
rect 81 245 82 246
rect 80 245 81 246
rect 79 245 80 246
rect 78 245 79 246
rect 77 245 78 246
rect 76 245 77 246
rect 75 245 76 246
rect 74 245 75 246
rect 73 245 74 246
rect 72 245 73 246
rect 71 245 72 246
rect 70 245 71 246
rect 69 245 70 246
rect 68 245 69 246
rect 67 245 68 246
rect 66 245 67 246
rect 65 245 66 246
rect 64 245 65 246
rect 63 245 64 246
rect 62 245 63 246
rect 61 245 62 246
rect 60 245 61 246
rect 59 245 60 246
rect 28 245 29 246
rect 27 245 28 246
rect 26 245 27 246
rect 25 245 26 246
rect 24 245 25 246
rect 23 245 24 246
rect 22 245 23 246
rect 21 245 22 246
rect 20 245 21 246
rect 19 245 20 246
rect 18 245 19 246
rect 17 245 18 246
rect 16 245 17 246
rect 15 245 16 246
rect 149 246 150 247
rect 148 246 149 247
rect 147 246 148 247
rect 146 246 147 247
rect 145 246 146 247
rect 144 246 145 247
rect 143 246 144 247
rect 142 246 143 247
rect 141 246 142 247
rect 140 246 141 247
rect 130 246 131 247
rect 129 246 130 247
rect 128 246 129 247
rect 127 246 128 247
rect 126 246 127 247
rect 125 246 126 247
rect 124 246 125 247
rect 123 246 124 247
rect 122 246 123 247
rect 121 246 122 247
rect 112 246 113 247
rect 111 246 112 247
rect 110 246 111 247
rect 109 246 110 247
rect 108 246 109 247
rect 107 246 108 247
rect 106 246 107 247
rect 105 246 106 247
rect 104 246 105 247
rect 103 246 104 247
rect 102 246 103 247
rect 86 246 87 247
rect 85 246 86 247
rect 84 246 85 247
rect 83 246 84 247
rect 82 246 83 247
rect 81 246 82 247
rect 80 246 81 247
rect 79 246 80 247
rect 78 246 79 247
rect 77 246 78 247
rect 76 246 77 247
rect 75 246 76 247
rect 74 246 75 247
rect 73 246 74 247
rect 72 246 73 247
rect 71 246 72 247
rect 70 246 71 247
rect 69 246 70 247
rect 68 246 69 247
rect 67 246 68 247
rect 66 246 67 247
rect 65 246 66 247
rect 64 246 65 247
rect 63 246 64 247
rect 62 246 63 247
rect 61 246 62 247
rect 60 246 61 247
rect 59 246 60 247
rect 27 246 28 247
rect 26 246 27 247
rect 25 246 26 247
rect 24 246 25 247
rect 23 246 24 247
rect 21 246 22 247
rect 20 246 21 247
rect 19 246 20 247
rect 18 246 19 247
rect 17 246 18 247
rect 16 246 17 247
rect 197 247 198 248
rect 196 247 197 248
rect 195 247 196 248
rect 194 247 195 248
rect 193 247 194 248
rect 192 247 193 248
rect 191 247 192 248
rect 173 247 174 248
rect 172 247 173 248
rect 149 247 150 248
rect 148 247 149 248
rect 147 247 148 248
rect 146 247 147 248
rect 145 247 146 248
rect 144 247 145 248
rect 143 247 144 248
rect 142 247 143 248
rect 141 247 142 248
rect 140 247 141 248
rect 130 247 131 248
rect 129 247 130 248
rect 128 247 129 248
rect 127 247 128 248
rect 126 247 127 248
rect 125 247 126 248
rect 124 247 125 248
rect 123 247 124 248
rect 122 247 123 248
rect 121 247 122 248
rect 112 247 113 248
rect 111 247 112 248
rect 110 247 111 248
rect 109 247 110 248
rect 108 247 109 248
rect 107 247 108 248
rect 106 247 107 248
rect 105 247 106 248
rect 104 247 105 248
rect 103 247 104 248
rect 102 247 103 248
rect 86 247 87 248
rect 85 247 86 248
rect 84 247 85 248
rect 83 247 84 248
rect 82 247 83 248
rect 81 247 82 248
rect 80 247 81 248
rect 79 247 80 248
rect 78 247 79 248
rect 77 247 78 248
rect 76 247 77 248
rect 75 247 76 248
rect 74 247 75 248
rect 73 247 74 248
rect 72 247 73 248
rect 71 247 72 248
rect 70 247 71 248
rect 69 247 70 248
rect 68 247 69 248
rect 67 247 68 248
rect 66 247 67 248
rect 65 247 66 248
rect 64 247 65 248
rect 63 247 64 248
rect 62 247 63 248
rect 61 247 62 248
rect 60 247 61 248
rect 59 247 60 248
rect 25 247 26 248
rect 24 247 25 248
rect 20 247 21 248
rect 19 247 20 248
rect 18 247 19 248
rect 17 247 18 248
rect 196 248 197 249
rect 195 248 196 249
rect 194 248 195 249
rect 193 248 194 249
rect 192 248 193 249
rect 191 248 192 249
rect 174 248 175 249
rect 173 248 174 249
rect 172 248 173 249
rect 165 248 166 249
rect 164 248 165 249
rect 163 248 164 249
rect 149 248 150 249
rect 148 248 149 249
rect 147 248 148 249
rect 146 248 147 249
rect 145 248 146 249
rect 144 248 145 249
rect 143 248 144 249
rect 142 248 143 249
rect 141 248 142 249
rect 140 248 141 249
rect 130 248 131 249
rect 129 248 130 249
rect 128 248 129 249
rect 127 248 128 249
rect 126 248 127 249
rect 125 248 126 249
rect 124 248 125 249
rect 123 248 124 249
rect 122 248 123 249
rect 121 248 122 249
rect 112 248 113 249
rect 111 248 112 249
rect 110 248 111 249
rect 109 248 110 249
rect 108 248 109 249
rect 107 248 108 249
rect 106 248 107 249
rect 105 248 106 249
rect 104 248 105 249
rect 103 248 104 249
rect 102 248 103 249
rect 86 248 87 249
rect 85 248 86 249
rect 84 248 85 249
rect 83 248 84 249
rect 82 248 83 249
rect 81 248 82 249
rect 80 248 81 249
rect 79 248 80 249
rect 78 248 79 249
rect 77 248 78 249
rect 76 248 77 249
rect 75 248 76 249
rect 74 248 75 249
rect 73 248 74 249
rect 72 248 73 249
rect 71 248 72 249
rect 70 248 71 249
rect 69 248 70 249
rect 68 248 69 249
rect 67 248 68 249
rect 66 248 67 249
rect 65 248 66 249
rect 64 248 65 249
rect 63 248 64 249
rect 62 248 63 249
rect 61 248 62 249
rect 60 248 61 249
rect 59 248 60 249
rect 192 249 193 250
rect 191 249 192 250
rect 174 249 175 250
rect 173 249 174 250
rect 172 249 173 250
rect 171 249 172 250
rect 165 249 166 250
rect 164 249 165 250
rect 163 249 164 250
rect 149 249 150 250
rect 148 249 149 250
rect 147 249 148 250
rect 146 249 147 250
rect 145 249 146 250
rect 144 249 145 250
rect 143 249 144 250
rect 142 249 143 250
rect 141 249 142 250
rect 140 249 141 250
rect 130 249 131 250
rect 129 249 130 250
rect 128 249 129 250
rect 127 249 128 250
rect 126 249 127 250
rect 125 249 126 250
rect 124 249 125 250
rect 123 249 124 250
rect 122 249 123 250
rect 121 249 122 250
rect 112 249 113 250
rect 111 249 112 250
rect 110 249 111 250
rect 109 249 110 250
rect 108 249 109 250
rect 107 249 108 250
rect 106 249 107 250
rect 105 249 106 250
rect 104 249 105 250
rect 103 249 104 250
rect 102 249 103 250
rect 76 249 77 250
rect 75 249 76 250
rect 74 249 75 250
rect 73 249 74 250
rect 72 249 73 250
rect 71 249 72 250
rect 70 249 71 250
rect 66 249 67 250
rect 65 249 66 250
rect 64 249 65 250
rect 63 249 64 250
rect 62 249 63 250
rect 61 249 62 250
rect 196 250 197 251
rect 195 250 196 251
rect 194 250 195 251
rect 193 250 194 251
rect 192 250 193 251
rect 191 250 192 251
rect 174 250 175 251
rect 173 250 174 251
rect 172 250 173 251
rect 171 250 172 251
rect 170 250 171 251
rect 165 250 166 251
rect 164 250 165 251
rect 163 250 164 251
rect 149 250 150 251
rect 148 250 149 251
rect 147 250 148 251
rect 146 250 147 251
rect 145 250 146 251
rect 144 250 145 251
rect 143 250 144 251
rect 142 250 143 251
rect 141 250 142 251
rect 140 250 141 251
rect 130 250 131 251
rect 129 250 130 251
rect 128 250 129 251
rect 127 250 128 251
rect 126 250 127 251
rect 125 250 126 251
rect 124 250 125 251
rect 123 250 124 251
rect 122 250 123 251
rect 121 250 122 251
rect 112 250 113 251
rect 111 250 112 251
rect 110 250 111 251
rect 109 250 110 251
rect 108 250 109 251
rect 107 250 108 251
rect 106 250 107 251
rect 105 250 106 251
rect 104 250 105 251
rect 103 250 104 251
rect 102 250 103 251
rect 77 250 78 251
rect 76 250 77 251
rect 75 250 76 251
rect 74 250 75 251
rect 73 250 74 251
rect 63 250 64 251
rect 62 250 63 251
rect 61 250 62 251
rect 60 250 61 251
rect 197 251 198 252
rect 196 251 197 252
rect 195 251 196 252
rect 194 251 195 252
rect 193 251 194 252
rect 192 251 193 252
rect 191 251 192 252
rect 182 251 183 252
rect 181 251 182 252
rect 180 251 181 252
rect 179 251 180 252
rect 178 251 179 252
rect 177 251 178 252
rect 176 251 177 252
rect 173 251 174 252
rect 172 251 173 252
rect 171 251 172 252
rect 170 251 171 252
rect 169 251 170 252
rect 165 251 166 252
rect 164 251 165 252
rect 163 251 164 252
rect 149 251 150 252
rect 148 251 149 252
rect 147 251 148 252
rect 146 251 147 252
rect 145 251 146 252
rect 144 251 145 252
rect 143 251 144 252
rect 142 251 143 252
rect 141 251 142 252
rect 140 251 141 252
rect 130 251 131 252
rect 129 251 130 252
rect 128 251 129 252
rect 127 251 128 252
rect 126 251 127 252
rect 125 251 126 252
rect 124 251 125 252
rect 123 251 124 252
rect 122 251 123 252
rect 121 251 122 252
rect 112 251 113 252
rect 111 251 112 252
rect 110 251 111 252
rect 109 251 110 252
rect 108 251 109 252
rect 107 251 108 252
rect 106 251 107 252
rect 105 251 106 252
rect 104 251 105 252
rect 103 251 104 252
rect 102 251 103 252
rect 77 251 78 252
rect 76 251 77 252
rect 75 251 76 252
rect 74 251 75 252
rect 62 251 63 252
rect 61 251 62 252
rect 60 251 61 252
rect 59 251 60 252
rect 196 252 197 253
rect 195 252 196 253
rect 194 252 195 253
rect 193 252 194 253
rect 192 252 193 253
rect 183 252 184 253
rect 182 252 183 253
rect 181 252 182 253
rect 180 252 181 253
rect 179 252 180 253
rect 178 252 179 253
rect 177 252 178 253
rect 176 252 177 253
rect 173 252 174 253
rect 172 252 173 253
rect 171 252 172 253
rect 170 252 171 253
rect 169 252 170 253
rect 168 252 169 253
rect 165 252 166 253
rect 164 252 165 253
rect 163 252 164 253
rect 78 252 79 253
rect 77 252 78 253
rect 76 252 77 253
rect 75 252 76 253
rect 62 252 63 253
rect 61 252 62 253
rect 60 252 61 253
rect 59 252 60 253
rect 195 253 196 254
rect 194 253 195 254
rect 193 253 194 254
rect 183 253 184 254
rect 182 253 183 254
rect 181 253 182 254
rect 180 253 181 254
rect 179 253 180 254
rect 178 253 179 254
rect 177 253 178 254
rect 176 253 177 254
rect 172 253 173 254
rect 171 253 172 254
rect 170 253 171 254
rect 169 253 170 254
rect 168 253 169 254
rect 167 253 168 254
rect 166 253 167 254
rect 165 253 166 254
rect 164 253 165 254
rect 163 253 164 254
rect 78 253 79 254
rect 77 253 78 254
rect 76 253 77 254
rect 75 253 76 254
rect 62 253 63 254
rect 61 253 62 254
rect 60 253 61 254
rect 59 253 60 254
rect 196 254 197 255
rect 195 254 196 255
rect 194 254 195 255
rect 193 254 194 255
rect 192 254 193 255
rect 191 254 192 255
rect 183 254 184 255
rect 182 254 183 255
rect 181 254 182 255
rect 180 254 181 255
rect 179 254 180 255
rect 178 254 179 255
rect 177 254 178 255
rect 176 254 177 255
rect 171 254 172 255
rect 170 254 171 255
rect 169 254 170 255
rect 168 254 169 255
rect 167 254 168 255
rect 166 254 167 255
rect 165 254 166 255
rect 164 254 165 255
rect 163 254 164 255
rect 78 254 79 255
rect 77 254 78 255
rect 76 254 77 255
rect 75 254 76 255
rect 62 254 63 255
rect 61 254 62 255
rect 60 254 61 255
rect 59 254 60 255
rect 58 254 59 255
rect 196 255 197 256
rect 195 255 196 256
rect 194 255 195 256
rect 193 255 194 256
rect 192 255 193 256
rect 191 255 192 256
rect 183 255 184 256
rect 182 255 183 256
rect 181 255 182 256
rect 180 255 181 256
rect 171 255 172 256
rect 170 255 171 256
rect 169 255 170 256
rect 168 255 169 256
rect 167 255 168 256
rect 166 255 167 256
rect 165 255 166 256
rect 164 255 165 256
rect 163 255 164 256
rect 78 255 79 256
rect 77 255 78 256
rect 76 255 77 256
rect 75 255 76 256
rect 62 255 63 256
rect 61 255 62 256
rect 60 255 61 256
rect 59 255 60 256
rect 58 255 59 256
rect 29 255 30 256
rect 28 255 29 256
rect 27 255 28 256
rect 26 255 27 256
rect 197 256 198 257
rect 196 256 197 257
rect 192 256 193 257
rect 191 256 192 257
rect 183 256 184 257
rect 182 256 183 257
rect 181 256 182 257
rect 180 256 181 257
rect 172 256 173 257
rect 171 256 172 257
rect 170 256 171 257
rect 169 256 170 257
rect 168 256 169 257
rect 167 256 168 257
rect 166 256 167 257
rect 165 256 166 257
rect 164 256 165 257
rect 163 256 164 257
rect 78 256 79 257
rect 77 256 78 257
rect 76 256 77 257
rect 75 256 76 257
rect 74 256 75 257
rect 63 256 64 257
rect 62 256 63 257
rect 61 256 62 257
rect 60 256 61 257
rect 59 256 60 257
rect 58 256 59 257
rect 29 256 30 257
rect 28 256 29 257
rect 27 256 28 257
rect 26 256 27 257
rect 25 256 26 257
rect 24 256 25 257
rect 23 256 24 257
rect 22 256 23 257
rect 21 256 22 257
rect 197 257 198 258
rect 196 257 197 258
rect 195 257 196 258
rect 194 257 195 258
rect 193 257 194 258
rect 192 257 193 258
rect 191 257 192 258
rect 190 257 191 258
rect 189 257 190 258
rect 188 257 189 258
rect 183 257 184 258
rect 182 257 183 258
rect 181 257 182 258
rect 180 257 181 258
rect 172 257 173 258
rect 171 257 172 258
rect 170 257 171 258
rect 169 257 170 258
rect 168 257 169 258
rect 165 257 166 258
rect 164 257 165 258
rect 163 257 164 258
rect 78 257 79 258
rect 77 257 78 258
rect 76 257 77 258
rect 75 257 76 258
rect 74 257 75 258
rect 73 257 74 258
rect 72 257 73 258
rect 65 257 66 258
rect 64 257 65 258
rect 63 257 64 258
rect 62 257 63 258
rect 61 257 62 258
rect 60 257 61 258
rect 59 257 60 258
rect 29 257 30 258
rect 28 257 29 258
rect 27 257 28 258
rect 26 257 27 258
rect 25 257 26 258
rect 24 257 25 258
rect 23 257 24 258
rect 22 257 23 258
rect 21 257 22 258
rect 20 257 21 258
rect 19 257 20 258
rect 18 257 19 258
rect 17 257 18 258
rect 16 257 17 258
rect 197 258 198 259
rect 196 258 197 259
rect 195 258 196 259
rect 194 258 195 259
rect 193 258 194 259
rect 192 258 193 259
rect 191 258 192 259
rect 190 258 191 259
rect 189 258 190 259
rect 188 258 189 259
rect 183 258 184 259
rect 182 258 183 259
rect 181 258 182 259
rect 180 258 181 259
rect 173 258 174 259
rect 172 258 173 259
rect 171 258 172 259
rect 170 258 171 259
rect 165 258 166 259
rect 164 258 165 259
rect 163 258 164 259
rect 78 258 79 259
rect 77 258 78 259
rect 76 258 77 259
rect 75 258 76 259
rect 74 258 75 259
rect 73 258 74 259
rect 72 258 73 259
rect 71 258 72 259
rect 70 258 71 259
rect 69 258 70 259
rect 68 258 69 259
rect 67 258 68 259
rect 66 258 67 259
rect 65 258 66 259
rect 64 258 65 259
rect 63 258 64 259
rect 62 258 63 259
rect 61 258 62 259
rect 60 258 61 259
rect 59 258 60 259
rect 26 258 27 259
rect 25 258 26 259
rect 24 258 25 259
rect 23 258 24 259
rect 22 258 23 259
rect 21 258 22 259
rect 20 258 21 259
rect 19 258 20 259
rect 18 258 19 259
rect 17 258 18 259
rect 16 258 17 259
rect 15 258 16 259
rect 14 258 15 259
rect 196 259 197 260
rect 195 259 196 260
rect 194 259 195 260
rect 193 259 194 260
rect 192 259 193 260
rect 191 259 192 260
rect 190 259 191 260
rect 189 259 190 260
rect 188 259 189 260
rect 183 259 184 260
rect 182 259 183 260
rect 181 259 182 260
rect 180 259 181 260
rect 173 259 174 260
rect 172 259 173 260
rect 171 259 172 260
rect 170 259 171 260
rect 165 259 166 260
rect 164 259 165 260
rect 163 259 164 260
rect 77 259 78 260
rect 76 259 77 260
rect 75 259 76 260
rect 74 259 75 260
rect 73 259 74 260
rect 72 259 73 260
rect 71 259 72 260
rect 70 259 71 260
rect 69 259 70 260
rect 68 259 69 260
rect 67 259 68 260
rect 66 259 67 260
rect 65 259 66 260
rect 64 259 65 260
rect 63 259 64 260
rect 62 259 63 260
rect 61 259 62 260
rect 60 259 61 260
rect 20 259 21 260
rect 19 259 20 260
rect 18 259 19 260
rect 17 259 18 260
rect 16 259 17 260
rect 15 259 16 260
rect 14 259 15 260
rect 183 260 184 261
rect 182 260 183 261
rect 181 260 182 261
rect 180 260 181 261
rect 174 260 175 261
rect 173 260 174 261
rect 172 260 173 261
rect 171 260 172 261
rect 165 260 166 261
rect 164 260 165 261
rect 163 260 164 261
rect 76 260 77 261
rect 75 260 76 261
rect 74 260 75 261
rect 73 260 74 261
rect 72 260 73 261
rect 71 260 72 261
rect 70 260 71 261
rect 69 260 70 261
rect 68 260 69 261
rect 67 260 68 261
rect 66 260 67 261
rect 65 260 66 261
rect 64 260 65 261
rect 63 260 64 261
rect 62 260 63 261
rect 61 260 62 261
rect 29 260 30 261
rect 28 260 29 261
rect 27 260 28 261
rect 26 260 27 261
rect 25 260 26 261
rect 24 260 25 261
rect 23 260 24 261
rect 22 260 23 261
rect 21 260 22 261
rect 20 260 21 261
rect 19 260 20 261
rect 18 260 19 261
rect 17 260 18 261
rect 16 260 17 261
rect 15 260 16 261
rect 14 260 15 261
rect 183 261 184 262
rect 182 261 183 262
rect 181 261 182 262
rect 180 261 181 262
rect 173 261 174 262
rect 172 261 173 262
rect 169 261 170 262
rect 168 261 169 262
rect 167 261 168 262
rect 166 261 167 262
rect 165 261 166 262
rect 164 261 165 262
rect 163 261 164 262
rect 75 261 76 262
rect 74 261 75 262
rect 73 261 74 262
rect 72 261 73 262
rect 71 261 72 262
rect 70 261 71 262
rect 69 261 70 262
rect 68 261 69 262
rect 67 261 68 262
rect 66 261 67 262
rect 65 261 66 262
rect 64 261 65 262
rect 63 261 64 262
rect 62 261 63 262
rect 29 261 30 262
rect 28 261 29 262
rect 27 261 28 262
rect 26 261 27 262
rect 25 261 26 262
rect 24 261 25 262
rect 23 261 24 262
rect 22 261 23 262
rect 21 261 22 262
rect 20 261 21 262
rect 19 261 20 262
rect 18 261 19 262
rect 17 261 18 262
rect 16 261 17 262
rect 15 261 16 262
rect 14 261 15 262
rect 183 262 184 263
rect 182 262 183 263
rect 181 262 182 263
rect 180 262 181 263
rect 172 262 173 263
rect 169 262 170 263
rect 168 262 169 263
rect 167 262 168 263
rect 166 262 167 263
rect 73 262 74 263
rect 72 262 73 263
rect 71 262 72 263
rect 70 262 71 263
rect 69 262 70 263
rect 68 262 69 263
rect 67 262 68 263
rect 66 262 67 263
rect 65 262 66 263
rect 64 262 65 263
rect 63 262 64 263
rect 29 262 30 263
rect 28 262 29 263
rect 27 262 28 263
rect 26 262 27 263
rect 25 262 26 263
rect 24 262 25 263
rect 23 262 24 263
rect 22 262 23 263
rect 21 262 22 263
rect 20 262 21 263
rect 19 262 20 263
rect 18 262 19 263
rect 17 262 18 263
rect 16 262 17 263
rect 15 262 16 263
rect 189 263 190 264
rect 183 263 184 264
rect 182 263 183 264
rect 181 263 182 264
rect 180 263 181 264
rect 169 263 170 264
rect 168 263 169 264
rect 167 263 168 264
rect 166 263 167 264
rect 69 263 70 264
rect 68 263 69 264
rect 67 263 68 264
rect 29 263 30 264
rect 28 263 29 264
rect 27 263 28 264
rect 26 263 27 264
rect 25 263 26 264
rect 24 263 25 264
rect 23 263 24 264
rect 189 264 190 265
rect 183 264 184 265
rect 182 264 183 265
rect 181 264 182 265
rect 180 264 181 265
rect 169 264 170 265
rect 168 264 169 265
rect 167 264 168 265
rect 166 264 167 265
rect 27 264 28 265
rect 26 264 27 265
rect 25 264 26 265
rect 24 264 25 265
rect 23 264 24 265
rect 22 264 23 265
rect 21 264 22 265
rect 190 265 191 266
rect 189 265 190 266
rect 183 265 184 266
rect 182 265 183 266
rect 181 265 182 266
rect 180 265 181 266
rect 177 265 178 266
rect 176 265 177 266
rect 175 265 176 266
rect 174 265 175 266
rect 173 265 174 266
rect 172 265 173 266
rect 171 265 172 266
rect 170 265 171 266
rect 169 265 170 266
rect 168 265 169 266
rect 167 265 168 266
rect 166 265 167 266
rect 165 265 166 266
rect 164 265 165 266
rect 163 265 164 266
rect 162 265 163 266
rect 112 265 113 266
rect 111 265 112 266
rect 110 265 111 266
rect 109 265 110 266
rect 108 265 109 266
rect 107 265 108 266
rect 106 265 107 266
rect 105 265 106 266
rect 104 265 105 266
rect 103 265 104 266
rect 102 265 103 266
rect 25 265 26 266
rect 24 265 25 266
rect 23 265 24 266
rect 22 265 23 266
rect 21 265 22 266
rect 20 265 21 266
rect 19 265 20 266
rect 197 266 198 267
rect 196 266 197 267
rect 195 266 196 267
rect 194 266 195 267
rect 193 266 194 267
rect 192 266 193 267
rect 191 266 192 267
rect 190 266 191 267
rect 189 266 190 267
rect 183 266 184 267
rect 182 266 183 267
rect 181 266 182 267
rect 180 266 181 267
rect 177 266 178 267
rect 176 266 177 267
rect 175 266 176 267
rect 174 266 175 267
rect 173 266 174 267
rect 172 266 173 267
rect 171 266 172 267
rect 170 266 171 267
rect 169 266 170 267
rect 168 266 169 267
rect 167 266 168 267
rect 166 266 167 267
rect 165 266 166 267
rect 164 266 165 267
rect 163 266 164 267
rect 162 266 163 267
rect 112 266 113 267
rect 111 266 112 267
rect 110 266 111 267
rect 109 266 110 267
rect 108 266 109 267
rect 107 266 108 267
rect 106 266 107 267
rect 105 266 106 267
rect 104 266 105 267
rect 103 266 104 267
rect 102 266 103 267
rect 73 266 74 267
rect 72 266 73 267
rect 71 266 72 267
rect 70 266 71 267
rect 69 266 70 267
rect 68 266 69 267
rect 67 266 68 267
rect 66 266 67 267
rect 65 266 66 267
rect 64 266 65 267
rect 29 266 30 267
rect 22 266 23 267
rect 21 266 22 267
rect 20 266 21 267
rect 19 266 20 267
rect 18 266 19 267
rect 17 266 18 267
rect 196 267 197 268
rect 195 267 196 268
rect 194 267 195 268
rect 193 267 194 268
rect 192 267 193 268
rect 191 267 192 268
rect 190 267 191 268
rect 189 267 190 268
rect 183 267 184 268
rect 182 267 183 268
rect 181 267 182 268
rect 180 267 181 268
rect 177 267 178 268
rect 176 267 177 268
rect 175 267 176 268
rect 174 267 175 268
rect 173 267 174 268
rect 172 267 173 268
rect 171 267 172 268
rect 170 267 171 268
rect 169 267 170 268
rect 168 267 169 268
rect 167 267 168 268
rect 166 267 167 268
rect 165 267 166 268
rect 164 267 165 268
rect 163 267 164 268
rect 162 267 163 268
rect 112 267 113 268
rect 111 267 112 268
rect 110 267 111 268
rect 109 267 110 268
rect 108 267 109 268
rect 107 267 108 268
rect 106 267 107 268
rect 105 267 106 268
rect 104 267 105 268
rect 103 267 104 268
rect 102 267 103 268
rect 75 267 76 268
rect 74 267 75 268
rect 73 267 74 268
rect 72 267 73 268
rect 71 267 72 268
rect 70 267 71 268
rect 69 267 70 268
rect 68 267 69 268
rect 67 267 68 268
rect 66 267 67 268
rect 65 267 66 268
rect 64 267 65 268
rect 63 267 64 268
rect 62 267 63 268
rect 29 267 30 268
rect 28 267 29 268
rect 27 267 28 268
rect 26 267 27 268
rect 25 267 26 268
rect 24 267 25 268
rect 20 267 21 268
rect 19 267 20 268
rect 18 267 19 268
rect 17 267 18 268
rect 16 267 17 268
rect 15 267 16 268
rect 189 268 190 269
rect 183 268 184 269
rect 182 268 183 269
rect 181 268 182 269
rect 180 268 181 269
rect 177 268 178 269
rect 176 268 177 269
rect 175 268 176 269
rect 174 268 175 269
rect 173 268 174 269
rect 172 268 173 269
rect 171 268 172 269
rect 170 268 171 269
rect 169 268 170 269
rect 168 268 169 269
rect 167 268 168 269
rect 166 268 167 269
rect 165 268 166 269
rect 164 268 165 269
rect 163 268 164 269
rect 162 268 163 269
rect 112 268 113 269
rect 111 268 112 269
rect 110 268 111 269
rect 109 268 110 269
rect 108 268 109 269
rect 107 268 108 269
rect 106 268 107 269
rect 105 268 106 269
rect 104 268 105 269
rect 103 268 104 269
rect 102 268 103 269
rect 76 268 77 269
rect 75 268 76 269
rect 74 268 75 269
rect 73 268 74 269
rect 72 268 73 269
rect 71 268 72 269
rect 70 268 71 269
rect 69 268 70 269
rect 68 268 69 269
rect 67 268 68 269
rect 66 268 67 269
rect 65 268 66 269
rect 64 268 65 269
rect 63 268 64 269
rect 62 268 63 269
rect 61 268 62 269
rect 29 268 30 269
rect 28 268 29 269
rect 27 268 28 269
rect 26 268 27 269
rect 25 268 26 269
rect 24 268 25 269
rect 23 268 24 269
rect 22 268 23 269
rect 21 268 22 269
rect 20 268 21 269
rect 19 268 20 269
rect 18 268 19 269
rect 17 268 18 269
rect 16 268 17 269
rect 15 268 16 269
rect 14 268 15 269
rect 195 269 196 270
rect 194 269 195 270
rect 193 269 194 270
rect 192 269 193 270
rect 189 269 190 270
rect 182 269 183 270
rect 181 269 182 270
rect 112 269 113 270
rect 111 269 112 270
rect 110 269 111 270
rect 109 269 110 270
rect 108 269 109 270
rect 107 269 108 270
rect 106 269 107 270
rect 105 269 106 270
rect 104 269 105 270
rect 103 269 104 270
rect 102 269 103 270
rect 77 269 78 270
rect 76 269 77 270
rect 75 269 76 270
rect 74 269 75 270
rect 73 269 74 270
rect 72 269 73 270
rect 71 269 72 270
rect 70 269 71 270
rect 69 269 70 270
rect 68 269 69 270
rect 67 269 68 270
rect 66 269 67 270
rect 65 269 66 270
rect 64 269 65 270
rect 63 269 64 270
rect 62 269 63 270
rect 61 269 62 270
rect 60 269 61 270
rect 28 269 29 270
rect 27 269 28 270
rect 26 269 27 270
rect 25 269 26 270
rect 24 269 25 270
rect 23 269 24 270
rect 22 269 23 270
rect 21 269 22 270
rect 20 269 21 270
rect 19 269 20 270
rect 18 269 19 270
rect 17 269 18 270
rect 16 269 17 270
rect 15 269 16 270
rect 14 269 15 270
rect 196 270 197 271
rect 195 270 196 271
rect 194 270 195 271
rect 193 270 194 271
rect 192 270 193 271
rect 191 270 192 271
rect 112 270 113 271
rect 111 270 112 271
rect 110 270 111 271
rect 109 270 110 271
rect 108 270 109 271
rect 107 270 108 271
rect 106 270 107 271
rect 105 270 106 271
rect 104 270 105 271
rect 103 270 104 271
rect 102 270 103 271
rect 77 270 78 271
rect 76 270 77 271
rect 75 270 76 271
rect 74 270 75 271
rect 73 270 74 271
rect 72 270 73 271
rect 71 270 72 271
rect 70 270 71 271
rect 69 270 70 271
rect 68 270 69 271
rect 67 270 68 271
rect 66 270 67 271
rect 65 270 66 271
rect 64 270 65 271
rect 63 270 64 271
rect 62 270 63 271
rect 61 270 62 271
rect 60 270 61 271
rect 23 270 24 271
rect 22 270 23 271
rect 21 270 22 271
rect 20 270 21 271
rect 19 270 20 271
rect 18 270 19 271
rect 17 270 18 271
rect 16 270 17 271
rect 15 270 16 271
rect 14 270 15 271
rect 197 271 198 272
rect 196 271 197 272
rect 195 271 196 272
rect 194 271 195 272
rect 193 271 194 272
rect 192 271 193 272
rect 191 271 192 272
rect 112 271 113 272
rect 111 271 112 272
rect 110 271 111 272
rect 109 271 110 272
rect 108 271 109 272
rect 107 271 108 272
rect 106 271 107 272
rect 105 271 106 272
rect 104 271 105 272
rect 103 271 104 272
rect 102 271 103 272
rect 78 271 79 272
rect 77 271 78 272
rect 76 271 77 272
rect 75 271 76 272
rect 74 271 75 272
rect 73 271 74 272
rect 72 271 73 272
rect 71 271 72 272
rect 70 271 71 272
rect 69 271 70 272
rect 68 271 69 272
rect 67 271 68 272
rect 66 271 67 272
rect 65 271 66 272
rect 64 271 65 272
rect 63 271 64 272
rect 62 271 63 272
rect 61 271 62 272
rect 60 271 61 272
rect 59 271 60 272
rect 18 271 19 272
rect 17 271 18 272
rect 16 271 17 272
rect 15 271 16 272
rect 14 271 15 272
rect 197 272 198 273
rect 196 272 197 273
rect 194 272 195 273
rect 192 272 193 273
rect 191 272 192 273
rect 112 272 113 273
rect 111 272 112 273
rect 110 272 111 273
rect 109 272 110 273
rect 108 272 109 273
rect 107 272 108 273
rect 106 272 107 273
rect 105 272 106 273
rect 104 272 105 273
rect 103 272 104 273
rect 102 272 103 273
rect 78 272 79 273
rect 77 272 78 273
rect 76 272 77 273
rect 75 272 76 273
rect 74 272 75 273
rect 70 272 71 273
rect 69 272 70 273
rect 68 272 69 273
rect 67 272 68 273
rect 63 272 64 273
rect 62 272 63 273
rect 61 272 62 273
rect 60 272 61 273
rect 59 272 60 273
rect 33 272 34 273
rect 32 272 33 273
rect 197 273 198 274
rect 196 273 197 274
rect 194 273 195 274
rect 193 273 194 274
rect 192 273 193 274
rect 191 273 192 274
rect 112 273 113 274
rect 111 273 112 274
rect 110 273 111 274
rect 109 273 110 274
rect 108 273 109 274
rect 107 273 108 274
rect 106 273 107 274
rect 105 273 106 274
rect 104 273 105 274
rect 103 273 104 274
rect 102 273 103 274
rect 78 273 79 274
rect 77 273 78 274
rect 76 273 77 274
rect 75 273 76 274
rect 74 273 75 274
rect 70 273 71 274
rect 69 273 70 274
rect 68 273 69 274
rect 67 273 68 274
rect 62 273 63 274
rect 61 273 62 274
rect 60 273 61 274
rect 59 273 60 274
rect 58 273 59 274
rect 33 273 34 274
rect 32 273 33 274
rect 19 273 20 274
rect 196 274 197 275
rect 194 274 195 275
rect 193 274 194 275
rect 192 274 193 275
rect 112 274 113 275
rect 111 274 112 275
rect 110 274 111 275
rect 109 274 110 275
rect 108 274 109 275
rect 107 274 108 275
rect 106 274 107 275
rect 105 274 106 275
rect 104 274 105 275
rect 103 274 104 275
rect 102 274 103 275
rect 78 274 79 275
rect 77 274 78 275
rect 76 274 77 275
rect 75 274 76 275
rect 70 274 71 275
rect 69 274 70 275
rect 68 274 69 275
rect 67 274 68 275
rect 62 274 63 275
rect 61 274 62 275
rect 60 274 61 275
rect 59 274 60 275
rect 58 274 59 275
rect 33 274 34 275
rect 32 274 33 275
rect 31 274 32 275
rect 25 274 26 275
rect 24 274 25 275
rect 23 274 24 275
rect 22 274 23 275
rect 21 274 22 275
rect 20 274 21 275
rect 19 274 20 275
rect 18 274 19 275
rect 112 275 113 276
rect 111 275 112 276
rect 110 275 111 276
rect 109 275 110 276
rect 108 275 109 276
rect 107 275 108 276
rect 106 275 107 276
rect 105 275 106 276
rect 104 275 105 276
rect 103 275 104 276
rect 102 275 103 276
rect 78 275 79 276
rect 77 275 78 276
rect 76 275 77 276
rect 75 275 76 276
rect 70 275 71 276
rect 69 275 70 276
rect 68 275 69 276
rect 67 275 68 276
rect 62 275 63 276
rect 61 275 62 276
rect 60 275 61 276
rect 59 275 60 276
rect 58 275 59 276
rect 33 275 34 276
rect 32 275 33 276
rect 31 275 32 276
rect 30 275 31 276
rect 29 275 30 276
rect 28 275 29 276
rect 27 275 28 276
rect 26 275 27 276
rect 25 275 26 276
rect 24 275 25 276
rect 23 275 24 276
rect 22 275 23 276
rect 21 275 22 276
rect 20 275 21 276
rect 19 275 20 276
rect 18 275 19 276
rect 196 276 197 277
rect 195 276 196 277
rect 194 276 195 277
rect 193 276 194 277
rect 192 276 193 277
rect 191 276 192 277
rect 190 276 191 277
rect 189 276 190 277
rect 188 276 189 277
rect 112 276 113 277
rect 111 276 112 277
rect 110 276 111 277
rect 109 276 110 277
rect 108 276 109 277
rect 107 276 108 277
rect 106 276 107 277
rect 105 276 106 277
rect 104 276 105 277
rect 103 276 104 277
rect 102 276 103 277
rect 78 276 79 277
rect 77 276 78 277
rect 76 276 77 277
rect 75 276 76 277
rect 70 276 71 277
rect 69 276 70 277
rect 68 276 69 277
rect 67 276 68 277
rect 62 276 63 277
rect 61 276 62 277
rect 60 276 61 277
rect 59 276 60 277
rect 58 276 59 277
rect 32 276 33 277
rect 31 276 32 277
rect 30 276 31 277
rect 29 276 30 277
rect 28 276 29 277
rect 27 276 28 277
rect 26 276 27 277
rect 25 276 26 277
rect 24 276 25 277
rect 23 276 24 277
rect 22 276 23 277
rect 21 276 22 277
rect 20 276 21 277
rect 19 276 20 277
rect 196 277 197 278
rect 195 277 196 278
rect 194 277 195 278
rect 193 277 194 278
rect 192 277 193 278
rect 191 277 192 278
rect 190 277 191 278
rect 189 277 190 278
rect 188 277 189 278
rect 112 277 113 278
rect 111 277 112 278
rect 110 277 111 278
rect 109 277 110 278
rect 108 277 109 278
rect 107 277 108 278
rect 106 277 107 278
rect 105 277 106 278
rect 104 277 105 278
rect 103 277 104 278
rect 102 277 103 278
rect 78 277 79 278
rect 77 277 78 278
rect 76 277 77 278
rect 75 277 76 278
rect 70 277 71 278
rect 69 277 70 278
rect 68 277 69 278
rect 67 277 68 278
rect 62 277 63 278
rect 61 277 62 278
rect 60 277 61 278
rect 59 277 60 278
rect 31 277 32 278
rect 30 277 31 278
rect 29 277 30 278
rect 28 277 29 278
rect 27 277 28 278
rect 26 277 27 278
rect 25 277 26 278
rect 112 278 113 279
rect 111 278 112 279
rect 110 278 111 279
rect 109 278 110 279
rect 108 278 109 279
rect 107 278 108 279
rect 106 278 107 279
rect 105 278 106 279
rect 104 278 105 279
rect 103 278 104 279
rect 102 278 103 279
rect 78 278 79 279
rect 77 278 78 279
rect 76 278 77 279
rect 75 278 76 279
rect 74 278 75 279
rect 73 278 74 279
rect 70 278 71 279
rect 69 278 70 279
rect 68 278 69 279
rect 67 278 68 279
rect 64 278 65 279
rect 63 278 64 279
rect 62 278 63 279
rect 61 278 62 279
rect 60 278 61 279
rect 59 278 60 279
rect 29 278 30 279
rect 28 278 29 279
rect 27 278 28 279
rect 26 278 27 279
rect 25 278 26 279
rect 24 278 25 279
rect 196 279 197 280
rect 195 279 196 280
rect 194 279 195 280
rect 193 279 194 280
rect 192 279 193 280
rect 112 279 113 280
rect 111 279 112 280
rect 110 279 111 280
rect 109 279 110 280
rect 108 279 109 280
rect 107 279 108 280
rect 106 279 107 280
rect 105 279 106 280
rect 104 279 105 280
rect 103 279 104 280
rect 102 279 103 280
rect 78 279 79 280
rect 77 279 78 280
rect 76 279 77 280
rect 75 279 76 280
rect 74 279 75 280
rect 73 279 74 280
rect 72 279 73 280
rect 70 279 71 280
rect 69 279 70 280
rect 68 279 69 280
rect 67 279 68 280
rect 66 279 67 280
rect 65 279 66 280
rect 64 279 65 280
rect 63 279 64 280
rect 62 279 63 280
rect 61 279 62 280
rect 60 279 61 280
rect 59 279 60 280
rect 28 279 29 280
rect 27 279 28 280
rect 26 279 27 280
rect 25 279 26 280
rect 24 279 25 280
rect 23 279 24 280
rect 22 279 23 280
rect 196 280 197 281
rect 195 280 196 281
rect 194 280 195 281
rect 193 280 194 281
rect 192 280 193 281
rect 191 280 192 281
rect 178 280 179 281
rect 112 280 113 281
rect 111 280 112 281
rect 110 280 111 281
rect 109 280 110 281
rect 108 280 109 281
rect 107 280 108 281
rect 106 280 107 281
rect 105 280 106 281
rect 104 280 105 281
rect 103 280 104 281
rect 102 280 103 281
rect 77 280 78 281
rect 76 280 77 281
rect 75 280 76 281
rect 74 280 75 281
rect 73 280 74 281
rect 70 280 71 281
rect 69 280 70 281
rect 68 280 69 281
rect 67 280 68 281
rect 66 280 67 281
rect 65 280 66 281
rect 64 280 65 281
rect 63 280 64 281
rect 62 280 63 281
rect 61 280 62 281
rect 60 280 61 281
rect 26 280 27 281
rect 25 280 26 281
rect 24 280 25 281
rect 23 280 24 281
rect 22 280 23 281
rect 21 280 22 281
rect 20 280 21 281
rect 197 281 198 282
rect 196 281 197 282
rect 194 281 195 282
rect 193 281 194 282
rect 192 281 193 282
rect 191 281 192 282
rect 179 281 180 282
rect 178 281 179 282
rect 177 281 178 282
rect 166 281 167 282
rect 112 281 113 282
rect 111 281 112 282
rect 110 281 111 282
rect 109 281 110 282
rect 108 281 109 282
rect 107 281 108 282
rect 106 281 107 282
rect 105 281 106 282
rect 104 281 105 282
rect 103 281 104 282
rect 102 281 103 282
rect 77 281 78 282
rect 76 281 77 282
rect 75 281 76 282
rect 74 281 75 282
rect 73 281 74 282
rect 70 281 71 282
rect 69 281 70 282
rect 68 281 69 282
rect 67 281 68 282
rect 66 281 67 282
rect 65 281 66 282
rect 64 281 65 282
rect 63 281 64 282
rect 62 281 63 282
rect 61 281 62 282
rect 24 281 25 282
rect 23 281 24 282
rect 22 281 23 282
rect 21 281 22 282
rect 20 281 21 282
rect 19 281 20 282
rect 197 282 198 283
rect 196 282 197 283
rect 194 282 195 283
rect 192 282 193 283
rect 191 282 192 283
rect 179 282 180 283
rect 178 282 179 283
rect 177 282 178 283
rect 176 282 177 283
rect 166 282 167 283
rect 165 282 166 283
rect 164 282 165 283
rect 112 282 113 283
rect 111 282 112 283
rect 110 282 111 283
rect 109 282 110 283
rect 108 282 109 283
rect 107 282 108 283
rect 106 282 107 283
rect 105 282 106 283
rect 104 282 105 283
rect 103 282 104 283
rect 102 282 103 283
rect 76 282 77 283
rect 75 282 76 283
rect 74 282 75 283
rect 73 282 74 283
rect 70 282 71 283
rect 69 282 70 283
rect 68 282 69 283
rect 67 282 68 283
rect 66 282 67 283
rect 65 282 66 283
rect 64 282 65 283
rect 63 282 64 283
rect 62 282 63 283
rect 22 282 23 283
rect 21 282 22 283
rect 20 282 21 283
rect 19 282 20 283
rect 18 282 19 283
rect 196 283 197 284
rect 194 283 195 284
rect 193 283 194 284
rect 192 283 193 284
rect 191 283 192 284
rect 179 283 180 284
rect 178 283 179 284
rect 177 283 178 284
rect 176 283 177 284
rect 175 283 176 284
rect 166 283 167 284
rect 165 283 166 284
rect 164 283 165 284
rect 112 283 113 284
rect 111 283 112 284
rect 110 283 111 284
rect 109 283 110 284
rect 108 283 109 284
rect 107 283 108 284
rect 106 283 107 284
rect 105 283 106 284
rect 104 283 105 284
rect 103 283 104 284
rect 102 283 103 284
rect 74 283 75 284
rect 73 283 74 284
rect 70 283 71 284
rect 69 283 70 284
rect 68 283 69 284
rect 67 283 68 284
rect 66 283 67 284
rect 65 283 66 284
rect 64 283 65 284
rect 63 283 64 284
rect 20 283 21 284
rect 19 283 20 284
rect 18 283 19 284
rect 196 284 197 285
rect 194 284 195 285
rect 193 284 194 285
rect 192 284 193 285
rect 179 284 180 285
rect 178 284 179 285
rect 177 284 178 285
rect 176 284 177 285
rect 175 284 176 285
rect 174 284 175 285
rect 166 284 167 285
rect 165 284 166 285
rect 164 284 165 285
rect 112 284 113 285
rect 111 284 112 285
rect 110 284 111 285
rect 109 284 110 285
rect 108 284 109 285
rect 107 284 108 285
rect 106 284 107 285
rect 105 284 106 285
rect 104 284 105 285
rect 103 284 104 285
rect 102 284 103 285
rect 69 284 70 285
rect 68 284 69 285
rect 67 284 68 285
rect 195 285 196 286
rect 194 285 195 286
rect 193 285 194 286
rect 178 285 179 286
rect 177 285 178 286
rect 176 285 177 286
rect 175 285 176 286
rect 174 285 175 286
rect 173 285 174 286
rect 166 285 167 286
rect 165 285 166 286
rect 164 285 165 286
rect 112 285 113 286
rect 111 285 112 286
rect 110 285 111 286
rect 109 285 110 286
rect 108 285 109 286
rect 107 285 108 286
rect 106 285 107 286
rect 105 285 106 286
rect 104 285 105 286
rect 103 285 104 286
rect 102 285 103 286
rect 196 286 197 287
rect 195 286 196 287
rect 194 286 195 287
rect 193 286 194 287
rect 192 286 193 287
rect 191 286 192 287
rect 177 286 178 287
rect 176 286 177 287
rect 175 286 176 287
rect 174 286 175 287
rect 173 286 174 287
rect 172 286 173 287
rect 171 286 172 287
rect 170 286 171 287
rect 169 286 170 287
rect 166 286 167 287
rect 165 286 166 287
rect 164 286 165 287
rect 112 286 113 287
rect 111 286 112 287
rect 110 286 111 287
rect 109 286 110 287
rect 108 286 109 287
rect 107 286 108 287
rect 106 286 107 287
rect 105 286 106 287
rect 104 286 105 287
rect 103 286 104 287
rect 102 286 103 287
rect 196 287 197 288
rect 195 287 196 288
rect 194 287 195 288
rect 193 287 194 288
rect 192 287 193 288
rect 191 287 192 288
rect 176 287 177 288
rect 175 287 176 288
rect 174 287 175 288
rect 173 287 174 288
rect 172 287 173 288
rect 171 287 172 288
rect 170 287 171 288
rect 169 287 170 288
rect 168 287 169 288
rect 167 287 168 288
rect 166 287 167 288
rect 165 287 166 288
rect 164 287 165 288
rect 112 287 113 288
rect 111 287 112 288
rect 110 287 111 288
rect 109 287 110 288
rect 108 287 109 288
rect 107 287 108 288
rect 106 287 107 288
rect 105 287 106 288
rect 104 287 105 288
rect 103 287 104 288
rect 102 287 103 288
rect 197 288 198 289
rect 196 288 197 289
rect 192 288 193 289
rect 191 288 192 289
rect 174 288 175 289
rect 173 288 174 289
rect 172 288 173 289
rect 171 288 172 289
rect 170 288 171 289
rect 169 288 170 289
rect 168 288 169 289
rect 167 288 168 289
rect 166 288 167 289
rect 165 288 166 289
rect 164 288 165 289
rect 112 288 113 289
rect 111 288 112 289
rect 110 288 111 289
rect 109 288 110 289
rect 108 288 109 289
rect 107 288 108 289
rect 106 288 107 289
rect 105 288 106 289
rect 104 288 105 289
rect 103 288 104 289
rect 102 288 103 289
rect 197 289 198 290
rect 196 289 197 290
rect 192 289 193 290
rect 191 289 192 290
rect 174 289 175 290
rect 173 289 174 290
rect 172 289 173 290
rect 171 289 172 290
rect 170 289 171 290
rect 169 289 170 290
rect 168 289 169 290
rect 167 289 168 290
rect 166 289 167 290
rect 165 289 166 290
rect 164 289 165 290
rect 112 289 113 290
rect 111 289 112 290
rect 110 289 111 290
rect 109 289 110 290
rect 108 289 109 290
rect 107 289 108 290
rect 106 289 107 290
rect 105 289 106 290
rect 104 289 105 290
rect 103 289 104 290
rect 102 289 103 290
rect 196 290 197 291
rect 195 290 196 291
rect 193 290 194 291
rect 176 290 177 291
rect 175 290 176 291
rect 174 290 175 291
rect 173 290 174 291
rect 172 290 173 291
rect 171 290 172 291
rect 170 290 171 291
rect 169 290 170 291
rect 168 290 169 291
rect 167 290 168 291
rect 166 290 167 291
rect 165 290 166 291
rect 164 290 165 291
rect 112 290 113 291
rect 111 290 112 291
rect 110 290 111 291
rect 109 290 110 291
rect 108 290 109 291
rect 107 290 108 291
rect 106 290 107 291
rect 105 290 106 291
rect 104 290 105 291
rect 103 290 104 291
rect 102 290 103 291
rect 196 291 197 292
rect 195 291 196 292
rect 194 291 195 292
rect 193 291 194 292
rect 192 291 193 292
rect 177 291 178 292
rect 176 291 177 292
rect 175 291 176 292
rect 174 291 175 292
rect 173 291 174 292
rect 172 291 173 292
rect 171 291 172 292
rect 166 291 167 292
rect 165 291 166 292
rect 164 291 165 292
rect 112 291 113 292
rect 111 291 112 292
rect 110 291 111 292
rect 109 291 110 292
rect 108 291 109 292
rect 107 291 108 292
rect 106 291 107 292
rect 105 291 106 292
rect 104 291 105 292
rect 103 291 104 292
rect 102 291 103 292
rect 25 291 26 292
rect 24 291 25 292
rect 23 291 24 292
rect 22 291 23 292
rect 21 291 22 292
rect 196 292 197 293
rect 195 292 196 293
rect 194 292 195 293
rect 193 292 194 293
rect 192 292 193 293
rect 191 292 192 293
rect 177 292 178 293
rect 176 292 177 293
rect 175 292 176 293
rect 174 292 175 293
rect 173 292 174 293
rect 166 292 167 293
rect 165 292 166 293
rect 164 292 165 293
rect 149 292 150 293
rect 148 292 149 293
rect 147 292 148 293
rect 146 292 147 293
rect 145 292 146 293
rect 144 292 145 293
rect 143 292 144 293
rect 142 292 143 293
rect 141 292 142 293
rect 140 292 141 293
rect 139 292 140 293
rect 138 292 139 293
rect 137 292 138 293
rect 136 292 137 293
rect 135 292 136 293
rect 134 292 135 293
rect 133 292 134 293
rect 132 292 133 293
rect 131 292 132 293
rect 130 292 131 293
rect 129 292 130 293
rect 128 292 129 293
rect 127 292 128 293
rect 126 292 127 293
rect 125 292 126 293
rect 124 292 125 293
rect 123 292 124 293
rect 122 292 123 293
rect 121 292 122 293
rect 120 292 121 293
rect 119 292 120 293
rect 118 292 119 293
rect 117 292 118 293
rect 116 292 117 293
rect 115 292 116 293
rect 114 292 115 293
rect 113 292 114 293
rect 112 292 113 293
rect 111 292 112 293
rect 110 292 111 293
rect 109 292 110 293
rect 108 292 109 293
rect 107 292 108 293
rect 106 292 107 293
rect 105 292 106 293
rect 104 292 105 293
rect 103 292 104 293
rect 102 292 103 293
rect 27 292 28 293
rect 26 292 27 293
rect 25 292 26 293
rect 24 292 25 293
rect 23 292 24 293
rect 22 292 23 293
rect 21 292 22 293
rect 20 292 21 293
rect 19 292 20 293
rect 18 292 19 293
rect 197 293 198 294
rect 196 293 197 294
rect 192 293 193 294
rect 191 293 192 294
rect 178 293 179 294
rect 177 293 178 294
rect 176 293 177 294
rect 175 293 176 294
rect 166 293 167 294
rect 165 293 166 294
rect 164 293 165 294
rect 149 293 150 294
rect 148 293 149 294
rect 147 293 148 294
rect 146 293 147 294
rect 145 293 146 294
rect 144 293 145 294
rect 143 293 144 294
rect 142 293 143 294
rect 141 293 142 294
rect 140 293 141 294
rect 139 293 140 294
rect 138 293 139 294
rect 137 293 138 294
rect 136 293 137 294
rect 135 293 136 294
rect 134 293 135 294
rect 133 293 134 294
rect 132 293 133 294
rect 131 293 132 294
rect 130 293 131 294
rect 129 293 130 294
rect 128 293 129 294
rect 127 293 128 294
rect 126 293 127 294
rect 125 293 126 294
rect 124 293 125 294
rect 123 293 124 294
rect 122 293 123 294
rect 121 293 122 294
rect 120 293 121 294
rect 119 293 120 294
rect 118 293 119 294
rect 117 293 118 294
rect 116 293 117 294
rect 115 293 116 294
rect 114 293 115 294
rect 113 293 114 294
rect 112 293 113 294
rect 111 293 112 294
rect 110 293 111 294
rect 109 293 110 294
rect 108 293 109 294
rect 107 293 108 294
rect 106 293 107 294
rect 105 293 106 294
rect 104 293 105 294
rect 103 293 104 294
rect 102 293 103 294
rect 28 293 29 294
rect 27 293 28 294
rect 26 293 27 294
rect 25 293 26 294
rect 24 293 25 294
rect 23 293 24 294
rect 22 293 23 294
rect 21 293 22 294
rect 20 293 21 294
rect 19 293 20 294
rect 18 293 19 294
rect 17 293 18 294
rect 197 294 198 295
rect 196 294 197 295
rect 192 294 193 295
rect 191 294 192 295
rect 179 294 180 295
rect 178 294 179 295
rect 177 294 178 295
rect 176 294 177 295
rect 175 294 176 295
rect 166 294 167 295
rect 165 294 166 295
rect 164 294 165 295
rect 149 294 150 295
rect 148 294 149 295
rect 147 294 148 295
rect 146 294 147 295
rect 145 294 146 295
rect 144 294 145 295
rect 143 294 144 295
rect 142 294 143 295
rect 141 294 142 295
rect 140 294 141 295
rect 139 294 140 295
rect 138 294 139 295
rect 137 294 138 295
rect 136 294 137 295
rect 135 294 136 295
rect 134 294 135 295
rect 133 294 134 295
rect 132 294 133 295
rect 131 294 132 295
rect 130 294 131 295
rect 129 294 130 295
rect 128 294 129 295
rect 127 294 128 295
rect 126 294 127 295
rect 125 294 126 295
rect 124 294 125 295
rect 123 294 124 295
rect 122 294 123 295
rect 121 294 122 295
rect 120 294 121 295
rect 119 294 120 295
rect 118 294 119 295
rect 117 294 118 295
rect 116 294 117 295
rect 115 294 116 295
rect 114 294 115 295
rect 113 294 114 295
rect 112 294 113 295
rect 111 294 112 295
rect 110 294 111 295
rect 109 294 110 295
rect 108 294 109 295
rect 107 294 108 295
rect 106 294 107 295
rect 105 294 106 295
rect 104 294 105 295
rect 103 294 104 295
rect 102 294 103 295
rect 29 294 30 295
rect 28 294 29 295
rect 27 294 28 295
rect 26 294 27 295
rect 25 294 26 295
rect 24 294 25 295
rect 23 294 24 295
rect 22 294 23 295
rect 21 294 22 295
rect 20 294 21 295
rect 19 294 20 295
rect 18 294 19 295
rect 17 294 18 295
rect 16 294 17 295
rect 196 295 197 296
rect 195 295 196 296
rect 194 295 195 296
rect 193 295 194 296
rect 192 295 193 296
rect 191 295 192 296
rect 178 295 179 296
rect 177 295 178 296
rect 176 295 177 296
rect 166 295 167 296
rect 165 295 166 296
rect 164 295 165 296
rect 149 295 150 296
rect 148 295 149 296
rect 147 295 148 296
rect 146 295 147 296
rect 145 295 146 296
rect 144 295 145 296
rect 143 295 144 296
rect 142 295 143 296
rect 141 295 142 296
rect 140 295 141 296
rect 139 295 140 296
rect 138 295 139 296
rect 137 295 138 296
rect 136 295 137 296
rect 135 295 136 296
rect 134 295 135 296
rect 133 295 134 296
rect 132 295 133 296
rect 131 295 132 296
rect 130 295 131 296
rect 129 295 130 296
rect 128 295 129 296
rect 127 295 128 296
rect 126 295 127 296
rect 125 295 126 296
rect 124 295 125 296
rect 123 295 124 296
rect 122 295 123 296
rect 121 295 122 296
rect 120 295 121 296
rect 119 295 120 296
rect 118 295 119 296
rect 117 295 118 296
rect 116 295 117 296
rect 115 295 116 296
rect 114 295 115 296
rect 113 295 114 296
rect 112 295 113 296
rect 111 295 112 296
rect 110 295 111 296
rect 109 295 110 296
rect 108 295 109 296
rect 107 295 108 296
rect 106 295 107 296
rect 105 295 106 296
rect 104 295 105 296
rect 103 295 104 296
rect 102 295 103 296
rect 29 295 30 296
rect 28 295 29 296
rect 27 295 28 296
rect 26 295 27 296
rect 19 295 20 296
rect 18 295 19 296
rect 17 295 18 296
rect 16 295 17 296
rect 15 295 16 296
rect 196 296 197 297
rect 195 296 196 297
rect 194 296 195 297
rect 193 296 194 297
rect 192 296 193 297
rect 177 296 178 297
rect 149 296 150 297
rect 148 296 149 297
rect 147 296 148 297
rect 146 296 147 297
rect 145 296 146 297
rect 144 296 145 297
rect 143 296 144 297
rect 142 296 143 297
rect 141 296 142 297
rect 140 296 141 297
rect 139 296 140 297
rect 138 296 139 297
rect 137 296 138 297
rect 136 296 137 297
rect 135 296 136 297
rect 134 296 135 297
rect 133 296 134 297
rect 132 296 133 297
rect 131 296 132 297
rect 130 296 131 297
rect 129 296 130 297
rect 128 296 129 297
rect 127 296 128 297
rect 126 296 127 297
rect 125 296 126 297
rect 124 296 125 297
rect 123 296 124 297
rect 122 296 123 297
rect 121 296 122 297
rect 120 296 121 297
rect 119 296 120 297
rect 118 296 119 297
rect 117 296 118 297
rect 116 296 117 297
rect 115 296 116 297
rect 114 296 115 297
rect 113 296 114 297
rect 112 296 113 297
rect 111 296 112 297
rect 110 296 111 297
rect 109 296 110 297
rect 108 296 109 297
rect 107 296 108 297
rect 106 296 107 297
rect 105 296 106 297
rect 104 296 105 297
rect 103 296 104 297
rect 102 296 103 297
rect 29 296 30 297
rect 28 296 29 297
rect 27 296 28 297
rect 17 296 18 297
rect 16 296 17 297
rect 15 296 16 297
rect 194 297 195 298
rect 149 297 150 298
rect 148 297 149 298
rect 147 297 148 298
rect 146 297 147 298
rect 145 297 146 298
rect 144 297 145 298
rect 143 297 144 298
rect 142 297 143 298
rect 141 297 142 298
rect 140 297 141 298
rect 139 297 140 298
rect 138 297 139 298
rect 137 297 138 298
rect 136 297 137 298
rect 135 297 136 298
rect 134 297 135 298
rect 133 297 134 298
rect 132 297 133 298
rect 131 297 132 298
rect 130 297 131 298
rect 129 297 130 298
rect 128 297 129 298
rect 127 297 128 298
rect 126 297 127 298
rect 125 297 126 298
rect 124 297 125 298
rect 123 297 124 298
rect 122 297 123 298
rect 121 297 122 298
rect 120 297 121 298
rect 119 297 120 298
rect 118 297 119 298
rect 117 297 118 298
rect 116 297 117 298
rect 115 297 116 298
rect 114 297 115 298
rect 113 297 114 298
rect 112 297 113 298
rect 111 297 112 298
rect 110 297 111 298
rect 109 297 110 298
rect 108 297 109 298
rect 107 297 108 298
rect 106 297 107 298
rect 105 297 106 298
rect 104 297 105 298
rect 103 297 104 298
rect 102 297 103 298
rect 29 297 30 298
rect 28 297 29 298
rect 27 297 28 298
rect 17 297 18 298
rect 16 297 17 298
rect 15 297 16 298
rect 14 297 15 298
rect 196 298 197 299
rect 195 298 196 299
rect 194 298 195 299
rect 193 298 194 299
rect 192 298 193 299
rect 191 298 192 299
rect 182 298 183 299
rect 181 298 182 299
rect 180 298 181 299
rect 179 298 180 299
rect 178 298 179 299
rect 177 298 178 299
rect 176 298 177 299
rect 175 298 176 299
rect 174 298 175 299
rect 173 298 174 299
rect 172 298 173 299
rect 171 298 172 299
rect 170 298 171 299
rect 169 298 170 299
rect 168 298 169 299
rect 167 298 168 299
rect 166 298 167 299
rect 165 298 166 299
rect 164 298 165 299
rect 163 298 164 299
rect 149 298 150 299
rect 148 298 149 299
rect 147 298 148 299
rect 146 298 147 299
rect 145 298 146 299
rect 144 298 145 299
rect 143 298 144 299
rect 142 298 143 299
rect 141 298 142 299
rect 140 298 141 299
rect 139 298 140 299
rect 138 298 139 299
rect 137 298 138 299
rect 136 298 137 299
rect 135 298 136 299
rect 134 298 135 299
rect 133 298 134 299
rect 132 298 133 299
rect 131 298 132 299
rect 130 298 131 299
rect 129 298 130 299
rect 128 298 129 299
rect 127 298 128 299
rect 126 298 127 299
rect 125 298 126 299
rect 124 298 125 299
rect 123 298 124 299
rect 122 298 123 299
rect 121 298 122 299
rect 120 298 121 299
rect 119 298 120 299
rect 118 298 119 299
rect 117 298 118 299
rect 116 298 117 299
rect 115 298 116 299
rect 114 298 115 299
rect 113 298 114 299
rect 112 298 113 299
rect 111 298 112 299
rect 110 298 111 299
rect 109 298 110 299
rect 108 298 109 299
rect 107 298 108 299
rect 106 298 107 299
rect 105 298 106 299
rect 104 298 105 299
rect 103 298 104 299
rect 102 298 103 299
rect 69 298 70 299
rect 68 298 69 299
rect 67 298 68 299
rect 29 298 30 299
rect 28 298 29 299
rect 27 298 28 299
rect 16 298 17 299
rect 15 298 16 299
rect 14 298 15 299
rect 197 299 198 300
rect 196 299 197 300
rect 195 299 196 300
rect 194 299 195 300
rect 193 299 194 300
rect 192 299 193 300
rect 191 299 192 300
rect 183 299 184 300
rect 182 299 183 300
rect 181 299 182 300
rect 180 299 181 300
rect 179 299 180 300
rect 178 299 179 300
rect 177 299 178 300
rect 176 299 177 300
rect 175 299 176 300
rect 174 299 175 300
rect 173 299 174 300
rect 172 299 173 300
rect 171 299 172 300
rect 170 299 171 300
rect 169 299 170 300
rect 168 299 169 300
rect 167 299 168 300
rect 166 299 167 300
rect 165 299 166 300
rect 164 299 165 300
rect 163 299 164 300
rect 162 299 163 300
rect 149 299 150 300
rect 148 299 149 300
rect 147 299 148 300
rect 146 299 147 300
rect 145 299 146 300
rect 144 299 145 300
rect 143 299 144 300
rect 142 299 143 300
rect 141 299 142 300
rect 140 299 141 300
rect 139 299 140 300
rect 138 299 139 300
rect 137 299 138 300
rect 136 299 137 300
rect 135 299 136 300
rect 134 299 135 300
rect 133 299 134 300
rect 132 299 133 300
rect 131 299 132 300
rect 130 299 131 300
rect 129 299 130 300
rect 128 299 129 300
rect 127 299 128 300
rect 126 299 127 300
rect 125 299 126 300
rect 124 299 125 300
rect 123 299 124 300
rect 122 299 123 300
rect 121 299 122 300
rect 120 299 121 300
rect 119 299 120 300
rect 118 299 119 300
rect 117 299 118 300
rect 116 299 117 300
rect 115 299 116 300
rect 114 299 115 300
rect 113 299 114 300
rect 112 299 113 300
rect 111 299 112 300
rect 110 299 111 300
rect 109 299 110 300
rect 108 299 109 300
rect 107 299 108 300
rect 106 299 107 300
rect 105 299 106 300
rect 104 299 105 300
rect 103 299 104 300
rect 102 299 103 300
rect 75 299 76 300
rect 74 299 75 300
rect 73 299 74 300
rect 72 299 73 300
rect 71 299 72 300
rect 70 299 71 300
rect 69 299 70 300
rect 68 299 69 300
rect 67 299 68 300
rect 66 299 67 300
rect 65 299 66 300
rect 64 299 65 300
rect 63 299 64 300
rect 62 299 63 300
rect 61 299 62 300
rect 29 299 30 300
rect 28 299 29 300
rect 27 299 28 300
rect 16 299 17 300
rect 15 299 16 300
rect 14 299 15 300
rect 192 300 193 301
rect 191 300 192 301
rect 183 300 184 301
rect 182 300 183 301
rect 181 300 182 301
rect 180 300 181 301
rect 179 300 180 301
rect 178 300 179 301
rect 177 300 178 301
rect 176 300 177 301
rect 175 300 176 301
rect 174 300 175 301
rect 173 300 174 301
rect 172 300 173 301
rect 171 300 172 301
rect 170 300 171 301
rect 169 300 170 301
rect 168 300 169 301
rect 167 300 168 301
rect 166 300 167 301
rect 165 300 166 301
rect 164 300 165 301
rect 163 300 164 301
rect 162 300 163 301
rect 149 300 150 301
rect 148 300 149 301
rect 147 300 148 301
rect 146 300 147 301
rect 145 300 146 301
rect 144 300 145 301
rect 143 300 144 301
rect 142 300 143 301
rect 141 300 142 301
rect 140 300 141 301
rect 139 300 140 301
rect 138 300 139 301
rect 137 300 138 301
rect 136 300 137 301
rect 135 300 136 301
rect 134 300 135 301
rect 133 300 134 301
rect 132 300 133 301
rect 131 300 132 301
rect 130 300 131 301
rect 129 300 130 301
rect 128 300 129 301
rect 127 300 128 301
rect 126 300 127 301
rect 125 300 126 301
rect 124 300 125 301
rect 123 300 124 301
rect 122 300 123 301
rect 121 300 122 301
rect 120 300 121 301
rect 119 300 120 301
rect 118 300 119 301
rect 117 300 118 301
rect 116 300 117 301
rect 115 300 116 301
rect 114 300 115 301
rect 113 300 114 301
rect 112 300 113 301
rect 111 300 112 301
rect 110 300 111 301
rect 109 300 110 301
rect 108 300 109 301
rect 107 300 108 301
rect 106 300 107 301
rect 105 300 106 301
rect 104 300 105 301
rect 103 300 104 301
rect 102 300 103 301
rect 78 300 79 301
rect 77 300 78 301
rect 76 300 77 301
rect 75 300 76 301
rect 74 300 75 301
rect 73 300 74 301
rect 72 300 73 301
rect 71 300 72 301
rect 70 300 71 301
rect 69 300 70 301
rect 68 300 69 301
rect 67 300 68 301
rect 66 300 67 301
rect 65 300 66 301
rect 64 300 65 301
rect 63 300 64 301
rect 62 300 63 301
rect 61 300 62 301
rect 60 300 61 301
rect 59 300 60 301
rect 58 300 59 301
rect 29 300 30 301
rect 28 300 29 301
rect 27 300 28 301
rect 26 300 27 301
rect 16 300 17 301
rect 15 300 16 301
rect 14 300 15 301
rect 192 301 193 302
rect 191 301 192 302
rect 183 301 184 302
rect 182 301 183 302
rect 181 301 182 302
rect 180 301 181 302
rect 179 301 180 302
rect 178 301 179 302
rect 177 301 178 302
rect 176 301 177 302
rect 175 301 176 302
rect 174 301 175 302
rect 173 301 174 302
rect 172 301 173 302
rect 171 301 172 302
rect 170 301 171 302
rect 169 301 170 302
rect 168 301 169 302
rect 167 301 168 302
rect 166 301 167 302
rect 165 301 166 302
rect 164 301 165 302
rect 163 301 164 302
rect 162 301 163 302
rect 149 301 150 302
rect 148 301 149 302
rect 147 301 148 302
rect 146 301 147 302
rect 145 301 146 302
rect 144 301 145 302
rect 143 301 144 302
rect 142 301 143 302
rect 141 301 142 302
rect 140 301 141 302
rect 139 301 140 302
rect 138 301 139 302
rect 137 301 138 302
rect 136 301 137 302
rect 135 301 136 302
rect 134 301 135 302
rect 133 301 134 302
rect 132 301 133 302
rect 131 301 132 302
rect 130 301 131 302
rect 129 301 130 302
rect 128 301 129 302
rect 127 301 128 302
rect 126 301 127 302
rect 125 301 126 302
rect 124 301 125 302
rect 123 301 124 302
rect 122 301 123 302
rect 121 301 122 302
rect 120 301 121 302
rect 119 301 120 302
rect 118 301 119 302
rect 117 301 118 302
rect 116 301 117 302
rect 115 301 116 302
rect 114 301 115 302
rect 113 301 114 302
rect 112 301 113 302
rect 111 301 112 302
rect 110 301 111 302
rect 109 301 110 302
rect 108 301 109 302
rect 107 301 108 302
rect 106 301 107 302
rect 105 301 106 302
rect 104 301 105 302
rect 103 301 104 302
rect 102 301 103 302
rect 81 301 82 302
rect 80 301 81 302
rect 79 301 80 302
rect 78 301 79 302
rect 77 301 78 302
rect 76 301 77 302
rect 75 301 76 302
rect 74 301 75 302
rect 73 301 74 302
rect 72 301 73 302
rect 71 301 72 302
rect 70 301 71 302
rect 69 301 70 302
rect 68 301 69 302
rect 67 301 68 302
rect 66 301 67 302
rect 65 301 66 302
rect 64 301 65 302
rect 63 301 64 302
rect 62 301 63 302
rect 61 301 62 302
rect 60 301 61 302
rect 59 301 60 302
rect 58 301 59 302
rect 57 301 58 302
rect 56 301 57 302
rect 28 301 29 302
rect 27 301 28 302
rect 26 301 27 302
rect 25 301 26 302
rect 17 301 18 302
rect 16 301 17 302
rect 15 301 16 302
rect 14 301 15 302
rect 197 302 198 303
rect 196 302 197 303
rect 195 302 196 303
rect 194 302 195 303
rect 193 302 194 303
rect 192 302 193 303
rect 191 302 192 303
rect 173 302 174 303
rect 172 302 173 303
rect 171 302 172 303
rect 170 302 171 303
rect 149 302 150 303
rect 148 302 149 303
rect 147 302 148 303
rect 146 302 147 303
rect 145 302 146 303
rect 144 302 145 303
rect 143 302 144 303
rect 142 302 143 303
rect 141 302 142 303
rect 140 302 141 303
rect 139 302 140 303
rect 138 302 139 303
rect 137 302 138 303
rect 136 302 137 303
rect 135 302 136 303
rect 134 302 135 303
rect 133 302 134 303
rect 132 302 133 303
rect 131 302 132 303
rect 130 302 131 303
rect 129 302 130 303
rect 128 302 129 303
rect 127 302 128 303
rect 126 302 127 303
rect 125 302 126 303
rect 124 302 125 303
rect 123 302 124 303
rect 122 302 123 303
rect 121 302 122 303
rect 120 302 121 303
rect 119 302 120 303
rect 118 302 119 303
rect 117 302 118 303
rect 116 302 117 303
rect 115 302 116 303
rect 114 302 115 303
rect 113 302 114 303
rect 112 302 113 303
rect 111 302 112 303
rect 110 302 111 303
rect 109 302 110 303
rect 108 302 109 303
rect 107 302 108 303
rect 106 302 107 303
rect 105 302 106 303
rect 104 302 105 303
rect 103 302 104 303
rect 102 302 103 303
rect 82 302 83 303
rect 81 302 82 303
rect 80 302 81 303
rect 79 302 80 303
rect 78 302 79 303
rect 77 302 78 303
rect 76 302 77 303
rect 75 302 76 303
rect 74 302 75 303
rect 73 302 74 303
rect 72 302 73 303
rect 71 302 72 303
rect 70 302 71 303
rect 69 302 70 303
rect 68 302 69 303
rect 67 302 68 303
rect 66 302 67 303
rect 65 302 66 303
rect 64 302 65 303
rect 63 302 64 303
rect 62 302 63 303
rect 61 302 62 303
rect 60 302 61 303
rect 59 302 60 303
rect 58 302 59 303
rect 57 302 58 303
rect 56 302 57 303
rect 55 302 56 303
rect 54 302 55 303
rect 27 302 28 303
rect 26 302 27 303
rect 25 302 26 303
rect 19 302 20 303
rect 18 302 19 303
rect 17 302 18 303
rect 16 302 17 303
rect 15 302 16 303
rect 196 303 197 304
rect 195 303 196 304
rect 194 303 195 304
rect 193 303 194 304
rect 192 303 193 304
rect 191 303 192 304
rect 173 303 174 304
rect 172 303 173 304
rect 171 303 172 304
rect 170 303 171 304
rect 149 303 150 304
rect 148 303 149 304
rect 147 303 148 304
rect 146 303 147 304
rect 145 303 146 304
rect 144 303 145 304
rect 143 303 144 304
rect 142 303 143 304
rect 141 303 142 304
rect 140 303 141 304
rect 139 303 140 304
rect 138 303 139 304
rect 137 303 138 304
rect 136 303 137 304
rect 135 303 136 304
rect 134 303 135 304
rect 133 303 134 304
rect 132 303 133 304
rect 131 303 132 304
rect 130 303 131 304
rect 129 303 130 304
rect 128 303 129 304
rect 127 303 128 304
rect 126 303 127 304
rect 125 303 126 304
rect 124 303 125 304
rect 123 303 124 304
rect 122 303 123 304
rect 121 303 122 304
rect 120 303 121 304
rect 119 303 120 304
rect 118 303 119 304
rect 117 303 118 304
rect 116 303 117 304
rect 115 303 116 304
rect 114 303 115 304
rect 113 303 114 304
rect 112 303 113 304
rect 111 303 112 304
rect 110 303 111 304
rect 109 303 110 304
rect 108 303 109 304
rect 107 303 108 304
rect 106 303 107 304
rect 105 303 106 304
rect 104 303 105 304
rect 103 303 104 304
rect 102 303 103 304
rect 84 303 85 304
rect 83 303 84 304
rect 82 303 83 304
rect 81 303 82 304
rect 80 303 81 304
rect 79 303 80 304
rect 78 303 79 304
rect 77 303 78 304
rect 76 303 77 304
rect 75 303 76 304
rect 74 303 75 304
rect 73 303 74 304
rect 72 303 73 304
rect 71 303 72 304
rect 70 303 71 304
rect 69 303 70 304
rect 68 303 69 304
rect 67 303 68 304
rect 66 303 67 304
rect 65 303 66 304
rect 64 303 65 304
rect 63 303 64 304
rect 62 303 63 304
rect 61 303 62 304
rect 60 303 61 304
rect 59 303 60 304
rect 58 303 59 304
rect 57 303 58 304
rect 56 303 57 304
rect 55 303 56 304
rect 54 303 55 304
rect 53 303 54 304
rect 26 303 27 304
rect 25 303 26 304
rect 19 303 20 304
rect 18 303 19 304
rect 17 303 18 304
rect 16 303 17 304
rect 192 304 193 305
rect 191 304 192 305
rect 173 304 174 305
rect 172 304 173 305
rect 171 304 172 305
rect 170 304 171 305
rect 149 304 150 305
rect 148 304 149 305
rect 147 304 148 305
rect 146 304 147 305
rect 145 304 146 305
rect 144 304 145 305
rect 143 304 144 305
rect 142 304 143 305
rect 141 304 142 305
rect 140 304 141 305
rect 139 304 140 305
rect 138 304 139 305
rect 137 304 138 305
rect 136 304 137 305
rect 135 304 136 305
rect 134 304 135 305
rect 133 304 134 305
rect 132 304 133 305
rect 131 304 132 305
rect 130 304 131 305
rect 129 304 130 305
rect 128 304 129 305
rect 127 304 128 305
rect 126 304 127 305
rect 125 304 126 305
rect 124 304 125 305
rect 123 304 124 305
rect 122 304 123 305
rect 121 304 122 305
rect 120 304 121 305
rect 119 304 120 305
rect 118 304 119 305
rect 117 304 118 305
rect 116 304 117 305
rect 115 304 116 305
rect 114 304 115 305
rect 113 304 114 305
rect 112 304 113 305
rect 111 304 112 305
rect 110 304 111 305
rect 109 304 110 305
rect 108 304 109 305
rect 107 304 108 305
rect 106 304 107 305
rect 105 304 106 305
rect 104 304 105 305
rect 103 304 104 305
rect 102 304 103 305
rect 85 304 86 305
rect 84 304 85 305
rect 83 304 84 305
rect 82 304 83 305
rect 81 304 82 305
rect 80 304 81 305
rect 79 304 80 305
rect 78 304 79 305
rect 77 304 78 305
rect 76 304 77 305
rect 75 304 76 305
rect 61 304 62 305
rect 60 304 61 305
rect 59 304 60 305
rect 58 304 59 305
rect 57 304 58 305
rect 56 304 57 305
rect 55 304 56 305
rect 54 304 55 305
rect 53 304 54 305
rect 52 304 53 305
rect 51 304 52 305
rect 18 304 19 305
rect 17 304 18 305
rect 196 305 197 306
rect 195 305 196 306
rect 194 305 195 306
rect 193 305 194 306
rect 192 305 193 306
rect 191 305 192 306
rect 172 305 173 306
rect 171 305 172 306
rect 149 305 150 306
rect 148 305 149 306
rect 147 305 148 306
rect 146 305 147 306
rect 145 305 146 306
rect 144 305 145 306
rect 143 305 144 306
rect 142 305 143 306
rect 141 305 142 306
rect 140 305 141 306
rect 139 305 140 306
rect 138 305 139 306
rect 137 305 138 306
rect 136 305 137 306
rect 135 305 136 306
rect 134 305 135 306
rect 133 305 134 306
rect 132 305 133 306
rect 131 305 132 306
rect 130 305 131 306
rect 129 305 130 306
rect 128 305 129 306
rect 127 305 128 306
rect 126 305 127 306
rect 125 305 126 306
rect 124 305 125 306
rect 123 305 124 306
rect 122 305 123 306
rect 121 305 122 306
rect 120 305 121 306
rect 119 305 120 306
rect 118 305 119 306
rect 117 305 118 306
rect 116 305 117 306
rect 115 305 116 306
rect 114 305 115 306
rect 113 305 114 306
rect 112 305 113 306
rect 111 305 112 306
rect 110 305 111 306
rect 109 305 110 306
rect 108 305 109 306
rect 107 305 108 306
rect 106 305 107 306
rect 105 305 106 306
rect 104 305 105 306
rect 103 305 104 306
rect 102 305 103 306
rect 86 305 87 306
rect 85 305 86 306
rect 84 305 85 306
rect 83 305 84 306
rect 82 305 83 306
rect 81 305 82 306
rect 80 305 81 306
rect 57 305 58 306
rect 56 305 57 306
rect 55 305 56 306
rect 54 305 55 306
rect 53 305 54 306
rect 52 305 53 306
rect 51 305 52 306
rect 197 306 198 307
rect 196 306 197 307
rect 195 306 196 307
rect 194 306 195 307
rect 193 306 194 307
rect 192 306 193 307
rect 191 306 192 307
rect 149 306 150 307
rect 148 306 149 307
rect 147 306 148 307
rect 146 306 147 307
rect 145 306 146 307
rect 144 306 145 307
rect 143 306 144 307
rect 142 306 143 307
rect 141 306 142 307
rect 140 306 141 307
rect 139 306 140 307
rect 138 306 139 307
rect 137 306 138 307
rect 136 306 137 307
rect 135 306 136 307
rect 134 306 135 307
rect 133 306 134 307
rect 132 306 133 307
rect 131 306 132 307
rect 130 306 131 307
rect 129 306 130 307
rect 128 306 129 307
rect 127 306 128 307
rect 126 306 127 307
rect 125 306 126 307
rect 124 306 125 307
rect 123 306 124 307
rect 122 306 123 307
rect 121 306 122 307
rect 120 306 121 307
rect 119 306 120 307
rect 118 306 119 307
rect 117 306 118 307
rect 116 306 117 307
rect 115 306 116 307
rect 114 306 115 307
rect 113 306 114 307
rect 112 306 113 307
rect 111 306 112 307
rect 110 306 111 307
rect 109 306 110 307
rect 108 306 109 307
rect 107 306 108 307
rect 106 306 107 307
rect 105 306 106 307
rect 104 306 105 307
rect 103 306 104 307
rect 102 306 103 307
rect 86 306 87 307
rect 85 306 86 307
rect 84 306 85 307
rect 83 306 84 307
rect 82 306 83 307
rect 55 306 56 307
rect 54 306 55 307
rect 53 306 54 307
rect 52 306 53 307
rect 51 306 52 307
rect 29 306 30 307
rect 28 306 29 307
rect 27 306 28 307
rect 26 306 27 307
rect 25 306 26 307
rect 196 307 197 308
rect 195 307 196 308
rect 194 307 195 308
rect 193 307 194 308
rect 192 307 193 308
rect 149 307 150 308
rect 148 307 149 308
rect 147 307 148 308
rect 146 307 147 308
rect 145 307 146 308
rect 144 307 145 308
rect 143 307 144 308
rect 142 307 143 308
rect 141 307 142 308
rect 140 307 141 308
rect 139 307 140 308
rect 138 307 139 308
rect 137 307 138 308
rect 136 307 137 308
rect 135 307 136 308
rect 134 307 135 308
rect 133 307 134 308
rect 132 307 133 308
rect 131 307 132 308
rect 130 307 131 308
rect 129 307 130 308
rect 128 307 129 308
rect 127 307 128 308
rect 126 307 127 308
rect 125 307 126 308
rect 124 307 125 308
rect 123 307 124 308
rect 122 307 123 308
rect 121 307 122 308
rect 120 307 121 308
rect 119 307 120 308
rect 118 307 119 308
rect 117 307 118 308
rect 116 307 117 308
rect 115 307 116 308
rect 114 307 115 308
rect 113 307 114 308
rect 112 307 113 308
rect 111 307 112 308
rect 110 307 111 308
rect 109 307 110 308
rect 108 307 109 308
rect 107 307 108 308
rect 106 307 107 308
rect 105 307 106 308
rect 104 307 105 308
rect 103 307 104 308
rect 102 307 103 308
rect 86 307 87 308
rect 85 307 86 308
rect 52 307 53 308
rect 51 307 52 308
rect 29 307 30 308
rect 28 307 29 308
rect 27 307 28 308
rect 26 307 27 308
rect 25 307 26 308
rect 24 307 25 308
rect 23 307 24 308
rect 22 307 23 308
rect 21 307 22 308
rect 20 307 21 308
rect 196 308 197 309
rect 192 308 193 309
rect 149 308 150 309
rect 148 308 149 309
rect 147 308 148 309
rect 146 308 147 309
rect 145 308 146 309
rect 144 308 145 309
rect 143 308 144 309
rect 142 308 143 309
rect 141 308 142 309
rect 140 308 141 309
rect 139 308 140 309
rect 138 308 139 309
rect 137 308 138 309
rect 136 308 137 309
rect 135 308 136 309
rect 134 308 135 309
rect 133 308 134 309
rect 132 308 133 309
rect 131 308 132 309
rect 130 308 131 309
rect 129 308 130 309
rect 128 308 129 309
rect 127 308 128 309
rect 126 308 127 309
rect 125 308 126 309
rect 124 308 125 309
rect 123 308 124 309
rect 122 308 123 309
rect 121 308 122 309
rect 120 308 121 309
rect 119 308 120 309
rect 118 308 119 309
rect 117 308 118 309
rect 116 308 117 309
rect 115 308 116 309
rect 114 308 115 309
rect 113 308 114 309
rect 112 308 113 309
rect 111 308 112 309
rect 110 308 111 309
rect 109 308 110 309
rect 108 308 109 309
rect 107 308 108 309
rect 106 308 107 309
rect 105 308 106 309
rect 104 308 105 309
rect 103 308 104 309
rect 102 308 103 309
rect 29 308 30 309
rect 28 308 29 309
rect 27 308 28 309
rect 26 308 27 309
rect 25 308 26 309
rect 24 308 25 309
rect 23 308 24 309
rect 22 308 23 309
rect 21 308 22 309
rect 20 308 21 309
rect 19 308 20 309
rect 18 308 19 309
rect 17 308 18 309
rect 16 308 17 309
rect 15 308 16 309
rect 197 309 198 310
rect 196 309 197 310
rect 195 309 196 310
rect 194 309 195 310
rect 193 309 194 310
rect 192 309 193 310
rect 191 309 192 310
rect 149 309 150 310
rect 148 309 149 310
rect 147 309 148 310
rect 146 309 147 310
rect 145 309 146 310
rect 144 309 145 310
rect 143 309 144 310
rect 142 309 143 310
rect 141 309 142 310
rect 140 309 141 310
rect 139 309 140 310
rect 138 309 139 310
rect 137 309 138 310
rect 136 309 137 310
rect 135 309 136 310
rect 134 309 135 310
rect 133 309 134 310
rect 132 309 133 310
rect 131 309 132 310
rect 130 309 131 310
rect 129 309 130 310
rect 128 309 129 310
rect 127 309 128 310
rect 126 309 127 310
rect 125 309 126 310
rect 124 309 125 310
rect 123 309 124 310
rect 122 309 123 310
rect 121 309 122 310
rect 120 309 121 310
rect 119 309 120 310
rect 118 309 119 310
rect 117 309 118 310
rect 116 309 117 310
rect 115 309 116 310
rect 114 309 115 310
rect 113 309 114 310
rect 112 309 113 310
rect 111 309 112 310
rect 110 309 111 310
rect 109 309 110 310
rect 108 309 109 310
rect 107 309 108 310
rect 106 309 107 310
rect 105 309 106 310
rect 104 309 105 310
rect 103 309 104 310
rect 102 309 103 310
rect 25 309 26 310
rect 24 309 25 310
rect 23 309 24 310
rect 22 309 23 310
rect 21 309 22 310
rect 20 309 21 310
rect 19 309 20 310
rect 18 309 19 310
rect 17 309 18 310
rect 16 309 17 310
rect 15 309 16 310
rect 14 309 15 310
rect 196 310 197 311
rect 195 310 196 311
rect 194 310 195 311
rect 193 310 194 311
rect 192 310 193 311
rect 191 310 192 311
rect 149 310 150 311
rect 148 310 149 311
rect 147 310 148 311
rect 146 310 147 311
rect 145 310 146 311
rect 144 310 145 311
rect 143 310 144 311
rect 142 310 143 311
rect 141 310 142 311
rect 140 310 141 311
rect 139 310 140 311
rect 138 310 139 311
rect 137 310 138 311
rect 136 310 137 311
rect 135 310 136 311
rect 134 310 135 311
rect 133 310 134 311
rect 132 310 133 311
rect 131 310 132 311
rect 130 310 131 311
rect 129 310 130 311
rect 128 310 129 311
rect 127 310 128 311
rect 126 310 127 311
rect 125 310 126 311
rect 124 310 125 311
rect 123 310 124 311
rect 122 310 123 311
rect 121 310 122 311
rect 120 310 121 311
rect 119 310 120 311
rect 118 310 119 311
rect 117 310 118 311
rect 116 310 117 311
rect 115 310 116 311
rect 114 310 115 311
rect 113 310 114 311
rect 112 310 113 311
rect 111 310 112 311
rect 110 310 111 311
rect 109 310 110 311
rect 108 310 109 311
rect 107 310 108 311
rect 106 310 107 311
rect 105 310 106 311
rect 104 310 105 311
rect 103 310 104 311
rect 102 310 103 311
rect 21 310 22 311
rect 20 310 21 311
rect 19 310 20 311
rect 18 310 19 311
rect 17 310 18 311
rect 16 310 17 311
rect 15 310 16 311
rect 14 310 15 311
rect 192 311 193 312
rect 191 311 192 312
rect 149 311 150 312
rect 148 311 149 312
rect 147 311 148 312
rect 146 311 147 312
rect 145 311 146 312
rect 144 311 145 312
rect 143 311 144 312
rect 142 311 143 312
rect 141 311 142 312
rect 140 311 141 312
rect 139 311 140 312
rect 138 311 139 312
rect 137 311 138 312
rect 136 311 137 312
rect 135 311 136 312
rect 134 311 135 312
rect 133 311 134 312
rect 132 311 133 312
rect 131 311 132 312
rect 130 311 131 312
rect 129 311 130 312
rect 128 311 129 312
rect 127 311 128 312
rect 126 311 127 312
rect 125 311 126 312
rect 124 311 125 312
rect 123 311 124 312
rect 122 311 123 312
rect 121 311 122 312
rect 120 311 121 312
rect 119 311 120 312
rect 118 311 119 312
rect 117 311 118 312
rect 116 311 117 312
rect 115 311 116 312
rect 114 311 115 312
rect 113 311 114 312
rect 112 311 113 312
rect 111 311 112 312
rect 110 311 111 312
rect 109 311 110 312
rect 108 311 109 312
rect 107 311 108 312
rect 106 311 107 312
rect 105 311 106 312
rect 104 311 105 312
rect 103 311 104 312
rect 102 311 103 312
rect 20 311 21 312
rect 19 311 20 312
rect 16 311 17 312
rect 15 311 16 312
rect 196 312 197 313
rect 195 312 196 313
rect 194 312 195 313
rect 193 312 194 313
rect 192 312 193 313
rect 191 312 192 313
rect 149 312 150 313
rect 148 312 149 313
rect 147 312 148 313
rect 146 312 147 313
rect 145 312 146 313
rect 144 312 145 313
rect 143 312 144 313
rect 142 312 143 313
rect 141 312 142 313
rect 140 312 141 313
rect 139 312 140 313
rect 138 312 139 313
rect 137 312 138 313
rect 136 312 137 313
rect 135 312 136 313
rect 134 312 135 313
rect 133 312 134 313
rect 132 312 133 313
rect 131 312 132 313
rect 130 312 131 313
rect 129 312 130 313
rect 128 312 129 313
rect 127 312 128 313
rect 126 312 127 313
rect 125 312 126 313
rect 124 312 125 313
rect 123 312 124 313
rect 122 312 123 313
rect 121 312 122 313
rect 120 312 121 313
rect 119 312 120 313
rect 118 312 119 313
rect 117 312 118 313
rect 116 312 117 313
rect 115 312 116 313
rect 114 312 115 313
rect 113 312 114 313
rect 112 312 113 313
rect 111 312 112 313
rect 110 312 111 313
rect 109 312 110 313
rect 108 312 109 313
rect 107 312 108 313
rect 106 312 107 313
rect 105 312 106 313
rect 104 312 105 313
rect 103 312 104 313
rect 102 312 103 313
rect 78 312 79 313
rect 77 312 78 313
rect 76 312 77 313
rect 75 312 76 313
rect 74 312 75 313
rect 73 312 74 313
rect 72 312 73 313
rect 71 312 72 313
rect 70 312 71 313
rect 69 312 70 313
rect 68 312 69 313
rect 67 312 68 313
rect 66 312 67 313
rect 65 312 66 313
rect 64 312 65 313
rect 63 312 64 313
rect 62 312 63 313
rect 61 312 62 313
rect 60 312 61 313
rect 59 312 60 313
rect 58 312 59 313
rect 57 312 58 313
rect 56 312 57 313
rect 55 312 56 313
rect 54 312 55 313
rect 53 312 54 313
rect 52 312 53 313
rect 51 312 52 313
rect 20 312 21 313
rect 19 312 20 313
rect 197 313 198 314
rect 196 313 197 314
rect 195 313 196 314
rect 194 313 195 314
rect 193 313 194 314
rect 192 313 193 314
rect 191 313 192 314
rect 149 313 150 314
rect 148 313 149 314
rect 147 313 148 314
rect 146 313 147 314
rect 145 313 146 314
rect 144 313 145 314
rect 143 313 144 314
rect 142 313 143 314
rect 141 313 142 314
rect 140 313 141 314
rect 139 313 140 314
rect 138 313 139 314
rect 137 313 138 314
rect 136 313 137 314
rect 135 313 136 314
rect 134 313 135 314
rect 133 313 134 314
rect 132 313 133 314
rect 131 313 132 314
rect 130 313 131 314
rect 129 313 130 314
rect 128 313 129 314
rect 127 313 128 314
rect 126 313 127 314
rect 125 313 126 314
rect 124 313 125 314
rect 123 313 124 314
rect 122 313 123 314
rect 121 313 122 314
rect 120 313 121 314
rect 119 313 120 314
rect 118 313 119 314
rect 117 313 118 314
rect 116 313 117 314
rect 115 313 116 314
rect 114 313 115 314
rect 113 313 114 314
rect 112 313 113 314
rect 111 313 112 314
rect 110 313 111 314
rect 109 313 110 314
rect 108 313 109 314
rect 107 313 108 314
rect 106 313 107 314
rect 105 313 106 314
rect 104 313 105 314
rect 103 313 104 314
rect 102 313 103 314
rect 78 313 79 314
rect 77 313 78 314
rect 76 313 77 314
rect 75 313 76 314
rect 74 313 75 314
rect 73 313 74 314
rect 72 313 73 314
rect 71 313 72 314
rect 70 313 71 314
rect 69 313 70 314
rect 68 313 69 314
rect 67 313 68 314
rect 66 313 67 314
rect 65 313 66 314
rect 64 313 65 314
rect 63 313 64 314
rect 62 313 63 314
rect 61 313 62 314
rect 60 313 61 314
rect 59 313 60 314
rect 58 313 59 314
rect 57 313 58 314
rect 56 313 57 314
rect 55 313 56 314
rect 54 313 55 314
rect 53 313 54 314
rect 52 313 53 314
rect 51 313 52 314
rect 29 313 30 314
rect 28 313 29 314
rect 27 313 28 314
rect 26 313 27 314
rect 25 313 26 314
rect 20 313 21 314
rect 19 313 20 314
rect 18 313 19 314
rect 192 314 193 315
rect 191 314 192 315
rect 174 314 175 315
rect 149 314 150 315
rect 148 314 149 315
rect 147 314 148 315
rect 146 314 147 315
rect 145 314 146 315
rect 144 314 145 315
rect 143 314 144 315
rect 142 314 143 315
rect 141 314 142 315
rect 140 314 141 315
rect 139 314 140 315
rect 138 314 139 315
rect 137 314 138 315
rect 136 314 137 315
rect 135 314 136 315
rect 134 314 135 315
rect 133 314 134 315
rect 132 314 133 315
rect 131 314 132 315
rect 130 314 131 315
rect 129 314 130 315
rect 128 314 129 315
rect 127 314 128 315
rect 126 314 127 315
rect 125 314 126 315
rect 124 314 125 315
rect 123 314 124 315
rect 122 314 123 315
rect 121 314 122 315
rect 120 314 121 315
rect 119 314 120 315
rect 118 314 119 315
rect 117 314 118 315
rect 116 314 117 315
rect 115 314 116 315
rect 114 314 115 315
rect 113 314 114 315
rect 112 314 113 315
rect 111 314 112 315
rect 110 314 111 315
rect 109 314 110 315
rect 108 314 109 315
rect 107 314 108 315
rect 106 314 107 315
rect 105 314 106 315
rect 104 314 105 315
rect 103 314 104 315
rect 102 314 103 315
rect 78 314 79 315
rect 77 314 78 315
rect 76 314 77 315
rect 75 314 76 315
rect 74 314 75 315
rect 73 314 74 315
rect 72 314 73 315
rect 71 314 72 315
rect 70 314 71 315
rect 69 314 70 315
rect 68 314 69 315
rect 67 314 68 315
rect 66 314 67 315
rect 65 314 66 315
rect 64 314 65 315
rect 63 314 64 315
rect 62 314 63 315
rect 61 314 62 315
rect 60 314 61 315
rect 59 314 60 315
rect 58 314 59 315
rect 57 314 58 315
rect 56 314 57 315
rect 55 314 56 315
rect 54 314 55 315
rect 53 314 54 315
rect 52 314 53 315
rect 51 314 52 315
rect 29 314 30 315
rect 28 314 29 315
rect 27 314 28 315
rect 26 314 27 315
rect 25 314 26 315
rect 24 314 25 315
rect 23 314 24 315
rect 22 314 23 315
rect 21 314 22 315
rect 20 314 21 315
rect 19 314 20 315
rect 18 314 19 315
rect 192 315 193 316
rect 191 315 192 316
rect 175 315 176 316
rect 174 315 175 316
rect 173 315 174 316
rect 149 315 150 316
rect 148 315 149 316
rect 147 315 148 316
rect 146 315 147 316
rect 145 315 146 316
rect 144 315 145 316
rect 143 315 144 316
rect 142 315 143 316
rect 141 315 142 316
rect 140 315 141 316
rect 139 315 140 316
rect 138 315 139 316
rect 137 315 138 316
rect 136 315 137 316
rect 135 315 136 316
rect 134 315 135 316
rect 133 315 134 316
rect 132 315 133 316
rect 131 315 132 316
rect 130 315 131 316
rect 129 315 130 316
rect 128 315 129 316
rect 127 315 128 316
rect 126 315 127 316
rect 125 315 126 316
rect 124 315 125 316
rect 123 315 124 316
rect 122 315 123 316
rect 121 315 122 316
rect 120 315 121 316
rect 119 315 120 316
rect 118 315 119 316
rect 117 315 118 316
rect 116 315 117 316
rect 115 315 116 316
rect 114 315 115 316
rect 113 315 114 316
rect 112 315 113 316
rect 111 315 112 316
rect 110 315 111 316
rect 109 315 110 316
rect 108 315 109 316
rect 107 315 108 316
rect 106 315 107 316
rect 105 315 106 316
rect 104 315 105 316
rect 103 315 104 316
rect 102 315 103 316
rect 78 315 79 316
rect 77 315 78 316
rect 76 315 77 316
rect 75 315 76 316
rect 74 315 75 316
rect 73 315 74 316
rect 72 315 73 316
rect 71 315 72 316
rect 70 315 71 316
rect 69 315 70 316
rect 68 315 69 316
rect 67 315 68 316
rect 66 315 67 316
rect 65 315 66 316
rect 64 315 65 316
rect 63 315 64 316
rect 62 315 63 316
rect 61 315 62 316
rect 60 315 61 316
rect 59 315 60 316
rect 58 315 59 316
rect 57 315 58 316
rect 56 315 57 316
rect 55 315 56 316
rect 54 315 55 316
rect 53 315 54 316
rect 52 315 53 316
rect 51 315 52 316
rect 29 315 30 316
rect 28 315 29 316
rect 27 315 28 316
rect 26 315 27 316
rect 25 315 26 316
rect 24 315 25 316
rect 23 315 24 316
rect 22 315 23 316
rect 21 315 22 316
rect 20 315 21 316
rect 19 315 20 316
rect 18 315 19 316
rect 196 316 197 317
rect 195 316 196 317
rect 194 316 195 317
rect 193 316 194 317
rect 192 316 193 317
rect 191 316 192 317
rect 175 316 176 317
rect 174 316 175 317
rect 173 316 174 317
rect 112 316 113 317
rect 111 316 112 317
rect 110 316 111 317
rect 109 316 110 317
rect 108 316 109 317
rect 107 316 108 317
rect 106 316 107 317
rect 105 316 106 317
rect 104 316 105 317
rect 103 316 104 317
rect 102 316 103 317
rect 78 316 79 317
rect 77 316 78 317
rect 76 316 77 317
rect 75 316 76 317
rect 74 316 75 317
rect 73 316 74 317
rect 72 316 73 317
rect 71 316 72 317
rect 70 316 71 317
rect 69 316 70 317
rect 68 316 69 317
rect 67 316 68 317
rect 66 316 67 317
rect 65 316 66 317
rect 64 316 65 317
rect 63 316 64 317
rect 62 316 63 317
rect 61 316 62 317
rect 60 316 61 317
rect 59 316 60 317
rect 58 316 59 317
rect 57 316 58 317
rect 56 316 57 317
rect 55 316 56 317
rect 54 316 55 317
rect 53 316 54 317
rect 52 316 53 317
rect 51 316 52 317
rect 26 316 27 317
rect 25 316 26 317
rect 24 316 25 317
rect 23 316 24 317
rect 22 316 23 317
rect 21 316 22 317
rect 20 316 21 317
rect 19 316 20 317
rect 196 317 197 318
rect 195 317 196 318
rect 194 317 195 318
rect 193 317 194 318
rect 192 317 193 318
rect 181 317 182 318
rect 180 317 181 318
rect 179 317 180 318
rect 175 317 176 318
rect 174 317 175 318
rect 173 317 174 318
rect 112 317 113 318
rect 111 317 112 318
rect 110 317 111 318
rect 109 317 110 318
rect 108 317 109 318
rect 107 317 108 318
rect 106 317 107 318
rect 105 317 106 318
rect 104 317 105 318
rect 103 317 104 318
rect 102 317 103 318
rect 78 317 79 318
rect 77 317 78 318
rect 76 317 77 318
rect 75 317 76 318
rect 74 317 75 318
rect 73 317 74 318
rect 72 317 73 318
rect 71 317 72 318
rect 70 317 71 318
rect 69 317 70 318
rect 68 317 69 318
rect 67 317 68 318
rect 66 317 67 318
rect 65 317 66 318
rect 64 317 65 318
rect 63 317 64 318
rect 62 317 63 318
rect 61 317 62 318
rect 60 317 61 318
rect 59 317 60 318
rect 58 317 59 318
rect 57 317 58 318
rect 56 317 57 318
rect 55 317 56 318
rect 54 317 55 318
rect 53 317 54 318
rect 52 317 53 318
rect 51 317 52 318
rect 21 317 22 318
rect 182 318 183 319
rect 181 318 182 319
rect 180 318 181 319
rect 179 318 180 319
rect 178 318 179 319
rect 175 318 176 319
rect 174 318 175 319
rect 173 318 174 319
rect 171 318 172 319
rect 170 318 171 319
rect 169 318 170 319
rect 168 318 169 319
rect 167 318 168 319
rect 166 318 167 319
rect 165 318 166 319
rect 164 318 165 319
rect 163 318 164 319
rect 162 318 163 319
rect 112 318 113 319
rect 111 318 112 319
rect 110 318 111 319
rect 109 318 110 319
rect 108 318 109 319
rect 107 318 108 319
rect 106 318 107 319
rect 105 318 106 319
rect 104 318 105 319
rect 103 318 104 319
rect 102 318 103 319
rect 66 318 67 319
rect 65 318 66 319
rect 64 318 65 319
rect 63 318 64 319
rect 62 318 63 319
rect 55 318 56 319
rect 54 318 55 319
rect 53 318 54 319
rect 52 318 53 319
rect 51 318 52 319
rect 196 319 197 320
rect 195 319 196 320
rect 194 319 195 320
rect 193 319 194 320
rect 192 319 193 320
rect 191 319 192 320
rect 182 319 183 320
rect 181 319 182 320
rect 180 319 181 320
rect 179 319 180 320
rect 178 319 179 320
rect 177 319 178 320
rect 175 319 176 320
rect 174 319 175 320
rect 173 319 174 320
rect 171 319 172 320
rect 170 319 171 320
rect 169 319 170 320
rect 168 319 169 320
rect 167 319 168 320
rect 166 319 167 320
rect 165 319 166 320
rect 164 319 165 320
rect 163 319 164 320
rect 162 319 163 320
rect 112 319 113 320
rect 111 319 112 320
rect 110 319 111 320
rect 109 319 110 320
rect 108 319 109 320
rect 107 319 108 320
rect 106 319 107 320
rect 105 319 106 320
rect 104 319 105 320
rect 103 319 104 320
rect 102 319 103 320
rect 66 319 67 320
rect 65 319 66 320
rect 64 319 65 320
rect 63 319 64 320
rect 62 319 63 320
rect 55 319 56 320
rect 54 319 55 320
rect 53 319 54 320
rect 52 319 53 320
rect 51 319 52 320
rect 29 319 30 320
rect 28 319 29 320
rect 27 319 28 320
rect 26 319 27 320
rect 25 319 26 320
rect 197 320 198 321
rect 196 320 197 321
rect 195 320 196 321
rect 194 320 195 321
rect 193 320 194 321
rect 192 320 193 321
rect 191 320 192 321
rect 183 320 184 321
rect 182 320 183 321
rect 181 320 182 321
rect 180 320 181 321
rect 179 320 180 321
rect 178 320 179 321
rect 177 320 178 321
rect 175 320 176 321
rect 174 320 175 321
rect 173 320 174 321
rect 171 320 172 321
rect 170 320 171 321
rect 169 320 170 321
rect 168 320 169 321
rect 167 320 168 321
rect 166 320 167 321
rect 165 320 166 321
rect 164 320 165 321
rect 163 320 164 321
rect 162 320 163 321
rect 112 320 113 321
rect 111 320 112 321
rect 110 320 111 321
rect 109 320 110 321
rect 108 320 109 321
rect 107 320 108 321
rect 106 320 107 321
rect 105 320 106 321
rect 104 320 105 321
rect 103 320 104 321
rect 102 320 103 321
rect 66 320 67 321
rect 65 320 66 321
rect 64 320 65 321
rect 63 320 64 321
rect 62 320 63 321
rect 55 320 56 321
rect 54 320 55 321
rect 53 320 54 321
rect 52 320 53 321
rect 51 320 52 321
rect 29 320 30 321
rect 28 320 29 321
rect 27 320 28 321
rect 26 320 27 321
rect 25 320 26 321
rect 24 320 25 321
rect 23 320 24 321
rect 22 320 23 321
rect 21 320 22 321
rect 20 320 21 321
rect 196 321 197 322
rect 183 321 184 322
rect 182 321 183 322
rect 181 321 182 322
rect 180 321 181 322
rect 179 321 180 322
rect 178 321 179 322
rect 177 321 178 322
rect 175 321 176 322
rect 174 321 175 322
rect 173 321 174 322
rect 171 321 172 322
rect 170 321 171 322
rect 169 321 170 322
rect 168 321 169 322
rect 167 321 168 322
rect 166 321 167 322
rect 165 321 166 322
rect 164 321 165 322
rect 163 321 164 322
rect 162 321 163 322
rect 112 321 113 322
rect 111 321 112 322
rect 110 321 111 322
rect 109 321 110 322
rect 108 321 109 322
rect 107 321 108 322
rect 106 321 107 322
rect 105 321 106 322
rect 104 321 105 322
rect 103 321 104 322
rect 102 321 103 322
rect 66 321 67 322
rect 65 321 66 322
rect 64 321 65 322
rect 63 321 64 322
rect 62 321 63 322
rect 55 321 56 322
rect 54 321 55 322
rect 53 321 54 322
rect 52 321 53 322
rect 51 321 52 322
rect 29 321 30 322
rect 28 321 29 322
rect 27 321 28 322
rect 26 321 27 322
rect 25 321 26 322
rect 24 321 25 322
rect 23 321 24 322
rect 22 321 23 322
rect 21 321 22 322
rect 20 321 21 322
rect 19 321 20 322
rect 16 321 17 322
rect 15 321 16 322
rect 196 322 197 323
rect 183 322 184 323
rect 182 322 183 323
rect 181 322 182 323
rect 179 322 180 323
rect 178 322 179 323
rect 177 322 178 323
rect 175 322 176 323
rect 174 322 175 323
rect 173 322 174 323
rect 171 322 172 323
rect 170 322 171 323
rect 169 322 170 323
rect 167 322 168 323
rect 166 322 167 323
rect 164 322 165 323
rect 163 322 164 323
rect 162 322 163 323
rect 112 322 113 323
rect 111 322 112 323
rect 110 322 111 323
rect 109 322 110 323
rect 108 322 109 323
rect 107 322 108 323
rect 106 322 107 323
rect 105 322 106 323
rect 104 322 105 323
rect 103 322 104 323
rect 102 322 103 323
rect 66 322 67 323
rect 65 322 66 323
rect 64 322 65 323
rect 63 322 64 323
rect 62 322 63 323
rect 55 322 56 323
rect 54 322 55 323
rect 53 322 54 323
rect 52 322 53 323
rect 51 322 52 323
rect 25 322 26 323
rect 24 322 25 323
rect 23 322 24 323
rect 22 322 23 323
rect 21 322 22 323
rect 20 322 21 323
rect 19 322 20 323
rect 18 322 19 323
rect 16 322 17 323
rect 15 322 16 323
rect 14 322 15 323
rect 197 323 198 324
rect 196 323 197 324
rect 195 323 196 324
rect 194 323 195 324
rect 193 323 194 324
rect 192 323 193 324
rect 191 323 192 324
rect 183 323 184 324
rect 182 323 183 324
rect 178 323 179 324
rect 177 323 178 324
rect 175 323 176 324
rect 174 323 175 324
rect 173 323 174 324
rect 171 323 172 324
rect 170 323 171 324
rect 169 323 170 324
rect 167 323 168 324
rect 166 323 167 324
rect 164 323 165 324
rect 163 323 164 324
rect 162 323 163 324
rect 112 323 113 324
rect 111 323 112 324
rect 110 323 111 324
rect 109 323 110 324
rect 108 323 109 324
rect 107 323 108 324
rect 106 323 107 324
rect 105 323 106 324
rect 104 323 105 324
rect 103 323 104 324
rect 102 323 103 324
rect 66 323 67 324
rect 65 323 66 324
rect 64 323 65 324
rect 63 323 64 324
rect 62 323 63 324
rect 55 323 56 324
rect 54 323 55 324
rect 53 323 54 324
rect 52 323 53 324
rect 51 323 52 324
rect 21 323 22 324
rect 20 323 21 324
rect 19 323 20 324
rect 16 323 17 324
rect 15 323 16 324
rect 14 323 15 324
rect 196 324 197 325
rect 195 324 196 325
rect 194 324 195 325
rect 193 324 194 325
rect 192 324 193 325
rect 191 324 192 325
rect 184 324 185 325
rect 183 324 184 325
rect 182 324 183 325
rect 178 324 179 325
rect 177 324 178 325
rect 176 324 177 325
rect 175 324 176 325
rect 174 324 175 325
rect 173 324 174 325
rect 171 324 172 325
rect 170 324 171 325
rect 169 324 170 325
rect 167 324 168 325
rect 166 324 167 325
rect 164 324 165 325
rect 163 324 164 325
rect 162 324 163 325
rect 112 324 113 325
rect 111 324 112 325
rect 110 324 111 325
rect 109 324 110 325
rect 108 324 109 325
rect 107 324 108 325
rect 106 324 107 325
rect 105 324 106 325
rect 104 324 105 325
rect 103 324 104 325
rect 102 324 103 325
rect 66 324 67 325
rect 65 324 66 325
rect 64 324 65 325
rect 63 324 64 325
rect 62 324 63 325
rect 55 324 56 325
rect 54 324 55 325
rect 53 324 54 325
rect 52 324 53 325
rect 51 324 52 325
rect 33 324 34 325
rect 32 324 33 325
rect 31 324 32 325
rect 30 324 31 325
rect 29 324 30 325
rect 28 324 29 325
rect 16 324 17 325
rect 15 324 16 325
rect 184 325 185 326
rect 183 325 184 326
rect 182 325 183 326
rect 178 325 179 326
rect 177 325 178 326
rect 176 325 177 326
rect 175 325 176 326
rect 174 325 175 326
rect 173 325 174 326
rect 172 325 173 326
rect 171 325 172 326
rect 170 325 171 326
rect 169 325 170 326
rect 167 325 168 326
rect 166 325 167 326
rect 164 325 165 326
rect 163 325 164 326
rect 162 325 163 326
rect 112 325 113 326
rect 111 325 112 326
rect 110 325 111 326
rect 109 325 110 326
rect 108 325 109 326
rect 107 325 108 326
rect 106 325 107 326
rect 105 325 106 326
rect 104 325 105 326
rect 103 325 104 326
rect 102 325 103 326
rect 66 325 67 326
rect 65 325 66 326
rect 64 325 65 326
rect 63 325 64 326
rect 62 325 63 326
rect 55 325 56 326
rect 54 325 55 326
rect 53 325 54 326
rect 52 325 53 326
rect 51 325 52 326
rect 33 325 34 326
rect 32 325 33 326
rect 31 325 32 326
rect 30 325 31 326
rect 29 325 30 326
rect 28 325 29 326
rect 27 325 28 326
rect 26 325 27 326
rect 25 325 26 326
rect 24 325 25 326
rect 196 326 197 327
rect 195 326 196 327
rect 194 326 195 327
rect 193 326 194 327
rect 192 326 193 327
rect 191 326 192 327
rect 184 326 185 327
rect 183 326 184 327
rect 182 326 183 327
rect 178 326 179 327
rect 177 326 178 327
rect 176 326 177 327
rect 175 326 176 327
rect 174 326 175 327
rect 173 326 174 327
rect 172 326 173 327
rect 171 326 172 327
rect 170 326 171 327
rect 169 326 170 327
rect 167 326 168 327
rect 166 326 167 327
rect 164 326 165 327
rect 163 326 164 327
rect 162 326 163 327
rect 112 326 113 327
rect 111 326 112 327
rect 110 326 111 327
rect 109 326 110 327
rect 108 326 109 327
rect 107 326 108 327
rect 106 326 107 327
rect 105 326 106 327
rect 104 326 105 327
rect 103 326 104 327
rect 102 326 103 327
rect 66 326 67 327
rect 65 326 66 327
rect 64 326 65 327
rect 63 326 64 327
rect 62 326 63 327
rect 55 326 56 327
rect 54 326 55 327
rect 53 326 54 327
rect 52 326 53 327
rect 51 326 52 327
rect 33 326 34 327
rect 32 326 33 327
rect 31 326 32 327
rect 30 326 31 327
rect 29 326 30 327
rect 28 326 29 327
rect 27 326 28 327
rect 26 326 27 327
rect 25 326 26 327
rect 24 326 25 327
rect 23 326 24 327
rect 22 326 23 327
rect 21 326 22 327
rect 20 326 21 327
rect 19 326 20 327
rect 197 327 198 328
rect 196 327 197 328
rect 195 327 196 328
rect 194 327 195 328
rect 193 327 194 328
rect 192 327 193 328
rect 191 327 192 328
rect 184 327 185 328
rect 183 327 184 328
rect 182 327 183 328
rect 178 327 179 328
rect 177 327 178 328
rect 176 327 177 328
rect 175 327 176 328
rect 174 327 175 328
rect 173 327 174 328
rect 172 327 173 328
rect 171 327 172 328
rect 170 327 171 328
rect 169 327 170 328
rect 167 327 168 328
rect 166 327 167 328
rect 164 327 165 328
rect 163 327 164 328
rect 162 327 163 328
rect 112 327 113 328
rect 111 327 112 328
rect 110 327 111 328
rect 109 327 110 328
rect 108 327 109 328
rect 107 327 108 328
rect 106 327 107 328
rect 105 327 106 328
rect 104 327 105 328
rect 103 327 104 328
rect 102 327 103 328
rect 66 327 67 328
rect 65 327 66 328
rect 64 327 65 328
rect 63 327 64 328
rect 62 327 63 328
rect 55 327 56 328
rect 54 327 55 328
rect 53 327 54 328
rect 52 327 53 328
rect 51 327 52 328
rect 29 327 30 328
rect 28 327 29 328
rect 27 327 28 328
rect 26 327 27 328
rect 25 327 26 328
rect 24 327 25 328
rect 23 327 24 328
rect 22 327 23 328
rect 21 327 22 328
rect 20 327 21 328
rect 19 327 20 328
rect 18 327 19 328
rect 196 328 197 329
rect 193 328 194 329
rect 192 328 193 329
rect 191 328 192 329
rect 184 328 185 329
rect 183 328 184 329
rect 182 328 183 329
rect 178 328 179 329
rect 177 328 178 329
rect 176 328 177 329
rect 175 328 176 329
rect 174 328 175 329
rect 173 328 174 329
rect 172 328 173 329
rect 171 328 172 329
rect 170 328 171 329
rect 169 328 170 329
rect 167 328 168 329
rect 166 328 167 329
rect 164 328 165 329
rect 163 328 164 329
rect 162 328 163 329
rect 112 328 113 329
rect 111 328 112 329
rect 110 328 111 329
rect 109 328 110 329
rect 108 328 109 329
rect 107 328 108 329
rect 106 328 107 329
rect 105 328 106 329
rect 104 328 105 329
rect 103 328 104 329
rect 102 328 103 329
rect 66 328 67 329
rect 65 328 66 329
rect 64 328 65 329
rect 63 328 64 329
rect 62 328 63 329
rect 55 328 56 329
rect 54 328 55 329
rect 53 328 54 329
rect 52 328 53 329
rect 51 328 52 329
rect 28 328 29 329
rect 27 328 28 329
rect 26 328 27 329
rect 25 328 26 329
rect 24 328 25 329
rect 23 328 24 329
rect 22 328 23 329
rect 21 328 22 329
rect 20 328 21 329
rect 19 328 20 329
rect 18 328 19 329
rect 192 329 193 330
rect 191 329 192 330
rect 184 329 185 330
rect 183 329 184 330
rect 182 329 183 330
rect 178 329 179 330
rect 177 329 178 330
rect 176 329 177 330
rect 175 329 176 330
rect 174 329 175 330
rect 173 329 174 330
rect 171 329 172 330
rect 170 329 171 330
rect 169 329 170 330
rect 167 329 168 330
rect 166 329 167 330
rect 164 329 165 330
rect 163 329 164 330
rect 162 329 163 330
rect 112 329 113 330
rect 111 329 112 330
rect 110 329 111 330
rect 109 329 110 330
rect 108 329 109 330
rect 107 329 108 330
rect 106 329 107 330
rect 105 329 106 330
rect 104 329 105 330
rect 103 329 104 330
rect 102 329 103 330
rect 55 329 56 330
rect 54 329 55 330
rect 53 329 54 330
rect 52 329 53 330
rect 51 329 52 330
rect 29 329 30 330
rect 28 329 29 330
rect 27 329 28 330
rect 21 329 22 330
rect 20 329 21 330
rect 19 329 20 330
rect 196 330 197 331
rect 195 330 196 331
rect 194 330 195 331
rect 193 330 194 331
rect 192 330 193 331
rect 191 330 192 331
rect 184 330 185 331
rect 183 330 184 331
rect 182 330 183 331
rect 179 330 180 331
rect 178 330 179 331
rect 177 330 178 331
rect 175 330 176 331
rect 174 330 175 331
rect 173 330 174 331
rect 171 330 172 331
rect 170 330 171 331
rect 169 330 170 331
rect 167 330 168 331
rect 166 330 167 331
rect 164 330 165 331
rect 163 330 164 331
rect 162 330 163 331
rect 112 330 113 331
rect 111 330 112 331
rect 110 330 111 331
rect 109 330 110 331
rect 108 330 109 331
rect 107 330 108 331
rect 106 330 107 331
rect 105 330 106 331
rect 104 330 105 331
rect 103 330 104 331
rect 102 330 103 331
rect 55 330 56 331
rect 54 330 55 331
rect 53 330 54 331
rect 52 330 53 331
rect 51 330 52 331
rect 29 330 30 331
rect 28 330 29 331
rect 20 330 21 331
rect 19 330 20 331
rect 197 331 198 332
rect 196 331 197 332
rect 195 331 196 332
rect 194 331 195 332
rect 193 331 194 332
rect 192 331 193 332
rect 191 331 192 332
rect 183 331 184 332
rect 182 331 183 332
rect 181 331 182 332
rect 179 331 180 332
rect 178 331 179 332
rect 177 331 178 332
rect 175 331 176 332
rect 174 331 175 332
rect 173 331 174 332
rect 171 331 172 332
rect 170 331 171 332
rect 169 331 170 332
rect 167 331 168 332
rect 166 331 167 332
rect 164 331 165 332
rect 163 331 164 332
rect 162 331 163 332
rect 112 331 113 332
rect 111 331 112 332
rect 110 331 111 332
rect 109 331 110 332
rect 108 331 109 332
rect 107 331 108 332
rect 106 331 107 332
rect 105 331 106 332
rect 104 331 105 332
rect 103 331 104 332
rect 102 331 103 332
rect 29 331 30 332
rect 28 331 29 332
rect 27 331 28 332
rect 19 331 20 332
rect 18 331 19 332
rect 183 332 184 333
rect 182 332 183 333
rect 181 332 182 333
rect 179 332 180 333
rect 178 332 179 333
rect 177 332 178 333
rect 175 332 176 333
rect 174 332 175 333
rect 173 332 174 333
rect 171 332 172 333
rect 170 332 171 333
rect 169 332 170 333
rect 167 332 168 333
rect 166 332 167 333
rect 164 332 165 333
rect 163 332 164 333
rect 162 332 163 333
rect 112 332 113 333
rect 111 332 112 333
rect 110 332 111 333
rect 109 332 110 333
rect 108 332 109 333
rect 107 332 108 333
rect 106 332 107 333
rect 105 332 106 333
rect 104 332 105 333
rect 103 332 104 333
rect 102 332 103 333
rect 29 332 30 333
rect 28 332 29 333
rect 27 332 28 333
rect 26 332 27 333
rect 20 332 21 333
rect 19 332 20 333
rect 18 332 19 333
rect 196 333 197 334
rect 195 333 196 334
rect 194 333 195 334
rect 193 333 194 334
rect 192 333 193 334
rect 191 333 192 334
rect 189 333 190 334
rect 188 333 189 334
rect 183 333 184 334
rect 182 333 183 334
rect 181 333 182 334
rect 180 333 181 334
rect 179 333 180 334
rect 178 333 179 334
rect 177 333 178 334
rect 175 333 176 334
rect 174 333 175 334
rect 173 333 174 334
rect 171 333 172 334
rect 170 333 171 334
rect 169 333 170 334
rect 167 333 168 334
rect 166 333 167 334
rect 164 333 165 334
rect 163 333 164 334
rect 162 333 163 334
rect 112 333 113 334
rect 111 333 112 334
rect 110 333 111 334
rect 109 333 110 334
rect 108 333 109 334
rect 107 333 108 334
rect 106 333 107 334
rect 105 333 106 334
rect 104 333 105 334
rect 103 333 104 334
rect 102 333 103 334
rect 28 333 29 334
rect 27 333 28 334
rect 26 333 27 334
rect 25 333 26 334
rect 24 333 25 334
rect 23 333 24 334
rect 22 333 23 334
rect 21 333 22 334
rect 20 333 21 334
rect 19 333 20 334
rect 18 333 19 334
rect 197 334 198 335
rect 196 334 197 335
rect 195 334 196 335
rect 194 334 195 335
rect 193 334 194 335
rect 192 334 193 335
rect 191 334 192 335
rect 189 334 190 335
rect 188 334 189 335
rect 183 334 184 335
rect 182 334 183 335
rect 181 334 182 335
rect 180 334 181 335
rect 179 334 180 335
rect 178 334 179 335
rect 175 334 176 335
rect 174 334 175 335
rect 173 334 174 335
rect 171 334 172 335
rect 170 334 171 335
rect 169 334 170 335
rect 167 334 168 335
rect 166 334 167 335
rect 164 334 165 335
rect 163 334 164 335
rect 162 334 163 335
rect 112 334 113 335
rect 111 334 112 335
rect 110 334 111 335
rect 109 334 110 335
rect 108 334 109 335
rect 107 334 108 335
rect 106 334 107 335
rect 105 334 106 335
rect 104 334 105 335
rect 103 334 104 335
rect 102 334 103 335
rect 27 334 28 335
rect 26 334 27 335
rect 25 334 26 335
rect 24 334 25 335
rect 23 334 24 335
rect 22 334 23 335
rect 21 334 22 335
rect 20 334 21 335
rect 19 334 20 335
rect 196 335 197 336
rect 194 335 195 336
rect 189 335 190 336
rect 182 335 183 336
rect 181 335 182 336
rect 180 335 181 336
rect 179 335 180 336
rect 178 335 179 336
rect 175 335 176 336
rect 174 335 175 336
rect 173 335 174 336
rect 171 335 172 336
rect 170 335 171 336
rect 169 335 170 336
rect 167 335 168 336
rect 166 335 167 336
rect 164 335 165 336
rect 163 335 164 336
rect 162 335 163 336
rect 112 335 113 336
rect 111 335 112 336
rect 110 335 111 336
rect 109 335 110 336
rect 108 335 109 336
rect 107 335 108 336
rect 106 335 107 336
rect 105 335 106 336
rect 104 335 105 336
rect 103 335 104 336
rect 102 335 103 336
rect 78 335 79 336
rect 77 335 78 336
rect 76 335 77 336
rect 75 335 76 336
rect 74 335 75 336
rect 73 335 74 336
rect 72 335 73 336
rect 71 335 72 336
rect 70 335 71 336
rect 69 335 70 336
rect 68 335 69 336
rect 67 335 68 336
rect 66 335 67 336
rect 65 335 66 336
rect 64 335 65 336
rect 63 335 64 336
rect 62 335 63 336
rect 61 335 62 336
rect 60 335 61 336
rect 59 335 60 336
rect 58 335 59 336
rect 57 335 58 336
rect 56 335 57 336
rect 55 335 56 336
rect 54 335 55 336
rect 53 335 54 336
rect 52 335 53 336
rect 51 335 52 336
rect 26 335 27 336
rect 25 335 26 336
rect 24 335 25 336
rect 23 335 24 336
rect 22 335 23 336
rect 21 335 22 336
rect 20 335 21 336
rect 19 335 20 336
rect 195 336 196 337
rect 194 336 195 337
rect 193 336 194 337
rect 192 336 193 337
rect 181 336 182 337
rect 180 336 181 337
rect 179 336 180 337
rect 175 336 176 337
rect 174 336 175 337
rect 173 336 174 337
rect 170 336 171 337
rect 169 336 170 337
rect 112 336 113 337
rect 111 336 112 337
rect 110 336 111 337
rect 109 336 110 337
rect 108 336 109 337
rect 107 336 108 337
rect 106 336 107 337
rect 105 336 106 337
rect 104 336 105 337
rect 103 336 104 337
rect 102 336 103 337
rect 78 336 79 337
rect 77 336 78 337
rect 76 336 77 337
rect 75 336 76 337
rect 74 336 75 337
rect 73 336 74 337
rect 72 336 73 337
rect 71 336 72 337
rect 70 336 71 337
rect 69 336 70 337
rect 68 336 69 337
rect 67 336 68 337
rect 66 336 67 337
rect 65 336 66 337
rect 64 336 65 337
rect 63 336 64 337
rect 62 336 63 337
rect 61 336 62 337
rect 60 336 61 337
rect 59 336 60 337
rect 58 336 59 337
rect 57 336 58 337
rect 56 336 57 337
rect 55 336 56 337
rect 54 336 55 337
rect 53 336 54 337
rect 52 336 53 337
rect 51 336 52 337
rect 24 336 25 337
rect 23 336 24 337
rect 22 336 23 337
rect 21 336 22 337
rect 196 337 197 338
rect 195 337 196 338
rect 194 337 195 338
rect 193 337 194 338
rect 192 337 193 338
rect 191 337 192 338
rect 175 337 176 338
rect 174 337 175 338
rect 173 337 174 338
rect 112 337 113 338
rect 111 337 112 338
rect 110 337 111 338
rect 109 337 110 338
rect 108 337 109 338
rect 107 337 108 338
rect 106 337 107 338
rect 105 337 106 338
rect 104 337 105 338
rect 103 337 104 338
rect 102 337 103 338
rect 78 337 79 338
rect 77 337 78 338
rect 76 337 77 338
rect 75 337 76 338
rect 74 337 75 338
rect 73 337 74 338
rect 72 337 73 338
rect 71 337 72 338
rect 70 337 71 338
rect 69 337 70 338
rect 68 337 69 338
rect 67 337 68 338
rect 66 337 67 338
rect 65 337 66 338
rect 64 337 65 338
rect 63 337 64 338
rect 62 337 63 338
rect 61 337 62 338
rect 60 337 61 338
rect 59 337 60 338
rect 58 337 59 338
rect 57 337 58 338
rect 56 337 57 338
rect 55 337 56 338
rect 54 337 55 338
rect 53 337 54 338
rect 52 337 53 338
rect 51 337 52 338
rect 196 338 197 339
rect 195 338 196 339
rect 192 338 193 339
rect 191 338 192 339
rect 175 338 176 339
rect 174 338 175 339
rect 173 338 174 339
rect 112 338 113 339
rect 111 338 112 339
rect 110 338 111 339
rect 109 338 110 339
rect 108 338 109 339
rect 107 338 108 339
rect 106 338 107 339
rect 105 338 106 339
rect 104 338 105 339
rect 103 338 104 339
rect 102 338 103 339
rect 78 338 79 339
rect 77 338 78 339
rect 76 338 77 339
rect 75 338 76 339
rect 74 338 75 339
rect 73 338 74 339
rect 72 338 73 339
rect 71 338 72 339
rect 70 338 71 339
rect 69 338 70 339
rect 68 338 69 339
rect 67 338 68 339
rect 66 338 67 339
rect 65 338 66 339
rect 64 338 65 339
rect 63 338 64 339
rect 62 338 63 339
rect 61 338 62 339
rect 60 338 61 339
rect 59 338 60 339
rect 58 338 59 339
rect 57 338 58 339
rect 56 338 57 339
rect 55 338 56 339
rect 54 338 55 339
rect 53 338 54 339
rect 52 338 53 339
rect 51 338 52 339
rect 197 339 198 340
rect 196 339 197 340
rect 192 339 193 340
rect 191 339 192 340
rect 174 339 175 340
rect 112 339 113 340
rect 111 339 112 340
rect 110 339 111 340
rect 109 339 110 340
rect 108 339 109 340
rect 107 339 108 340
rect 106 339 107 340
rect 105 339 106 340
rect 104 339 105 340
rect 103 339 104 340
rect 102 339 103 340
rect 78 339 79 340
rect 77 339 78 340
rect 76 339 77 340
rect 75 339 76 340
rect 74 339 75 340
rect 73 339 74 340
rect 72 339 73 340
rect 71 339 72 340
rect 70 339 71 340
rect 69 339 70 340
rect 68 339 69 340
rect 67 339 68 340
rect 66 339 67 340
rect 65 339 66 340
rect 64 339 65 340
rect 63 339 64 340
rect 62 339 63 340
rect 61 339 62 340
rect 60 339 61 340
rect 59 339 60 340
rect 58 339 59 340
rect 57 339 58 340
rect 56 339 57 340
rect 55 339 56 340
rect 54 339 55 340
rect 53 339 54 340
rect 52 339 53 340
rect 51 339 52 340
rect 196 340 197 341
rect 192 340 193 341
rect 191 340 192 341
rect 112 340 113 341
rect 111 340 112 341
rect 110 340 111 341
rect 109 340 110 341
rect 108 340 109 341
rect 107 340 108 341
rect 106 340 107 341
rect 105 340 106 341
rect 104 340 105 341
rect 103 340 104 341
rect 102 340 103 341
rect 78 340 79 341
rect 77 340 78 341
rect 76 340 77 341
rect 75 340 76 341
rect 74 340 75 341
rect 73 340 74 341
rect 72 340 73 341
rect 71 340 72 341
rect 70 340 71 341
rect 69 340 70 341
rect 68 340 69 341
rect 67 340 68 341
rect 66 340 67 341
rect 65 340 66 341
rect 64 340 65 341
rect 63 340 64 341
rect 62 340 63 341
rect 61 340 62 341
rect 60 340 61 341
rect 59 340 60 341
rect 58 340 59 341
rect 57 340 58 341
rect 56 340 57 341
rect 55 340 56 341
rect 54 340 55 341
rect 53 340 54 341
rect 52 340 53 341
rect 51 340 52 341
rect 195 341 196 342
rect 112 341 113 342
rect 111 341 112 342
rect 110 341 111 342
rect 109 341 110 342
rect 108 341 109 342
rect 107 341 108 342
rect 106 341 107 342
rect 105 341 106 342
rect 104 341 105 342
rect 103 341 104 342
rect 102 341 103 342
rect 196 342 197 343
rect 195 342 196 343
rect 194 342 195 343
rect 192 342 193 343
rect 191 342 192 343
rect 112 342 113 343
rect 111 342 112 343
rect 110 342 111 343
rect 109 342 110 343
rect 108 342 109 343
rect 107 342 108 343
rect 106 342 107 343
rect 105 342 106 343
rect 104 342 105 343
rect 103 342 104 343
rect 102 342 103 343
rect 197 343 198 344
rect 196 343 197 344
rect 195 343 196 344
rect 194 343 195 344
rect 193 343 194 344
rect 192 343 193 344
rect 191 343 192 344
rect 29 343 30 344
rect 28 343 29 344
rect 197 344 198 345
rect 196 344 197 345
rect 194 344 195 345
rect 193 344 194 345
rect 192 344 193 345
rect 191 344 192 345
rect 29 344 30 345
rect 28 344 29 345
rect 27 344 28 345
rect 26 344 27 345
rect 25 344 26 345
rect 24 344 25 345
rect 196 345 197 346
rect 195 345 196 346
rect 194 345 195 346
rect 193 345 194 346
rect 192 345 193 346
rect 191 345 192 346
rect 29 345 30 346
rect 28 345 29 346
rect 27 345 28 346
rect 26 345 27 346
rect 25 345 26 346
rect 24 345 25 346
rect 23 345 24 346
rect 22 345 23 346
rect 21 345 22 346
rect 20 345 21 346
rect 19 345 20 346
rect 197 346 198 347
rect 196 346 197 347
rect 195 346 196 347
rect 194 346 195 347
rect 193 346 194 347
rect 192 346 193 347
rect 191 346 192 347
rect 78 346 79 347
rect 77 346 78 347
rect 76 346 77 347
rect 75 346 76 347
rect 74 346 75 347
rect 73 346 74 347
rect 72 346 73 347
rect 71 346 72 347
rect 70 346 71 347
rect 69 346 70 347
rect 68 346 69 347
rect 67 346 68 347
rect 66 346 67 347
rect 65 346 66 347
rect 64 346 65 347
rect 63 346 64 347
rect 62 346 63 347
rect 61 346 62 347
rect 60 346 61 347
rect 59 346 60 347
rect 58 346 59 347
rect 57 346 58 347
rect 56 346 57 347
rect 55 346 56 347
rect 54 346 55 347
rect 53 346 54 347
rect 52 346 53 347
rect 51 346 52 347
rect 28 346 29 347
rect 27 346 28 347
rect 26 346 27 347
rect 25 346 26 347
rect 24 346 25 347
rect 23 346 24 347
rect 22 346 23 347
rect 21 346 22 347
rect 20 346 21 347
rect 19 346 20 347
rect 18 346 19 347
rect 17 346 18 347
rect 16 346 17 347
rect 15 346 16 347
rect 196 347 197 348
rect 78 347 79 348
rect 77 347 78 348
rect 76 347 77 348
rect 75 347 76 348
rect 74 347 75 348
rect 73 347 74 348
rect 72 347 73 348
rect 71 347 72 348
rect 70 347 71 348
rect 69 347 70 348
rect 68 347 69 348
rect 67 347 68 348
rect 66 347 67 348
rect 65 347 66 348
rect 64 347 65 348
rect 63 347 64 348
rect 62 347 63 348
rect 61 347 62 348
rect 60 347 61 348
rect 59 347 60 348
rect 58 347 59 348
rect 57 347 58 348
rect 56 347 57 348
rect 55 347 56 348
rect 54 347 55 348
rect 53 347 54 348
rect 52 347 53 348
rect 51 347 52 348
rect 23 347 24 348
rect 22 347 23 348
rect 21 347 22 348
rect 20 347 21 348
rect 19 347 20 348
rect 18 347 19 348
rect 17 347 18 348
rect 16 347 17 348
rect 15 347 16 348
rect 14 347 15 348
rect 192 348 193 349
rect 191 348 192 349
rect 78 348 79 349
rect 77 348 78 349
rect 76 348 77 349
rect 75 348 76 349
rect 74 348 75 349
rect 73 348 74 349
rect 72 348 73 349
rect 71 348 72 349
rect 70 348 71 349
rect 69 348 70 349
rect 68 348 69 349
rect 67 348 68 349
rect 66 348 67 349
rect 65 348 66 349
rect 64 348 65 349
rect 63 348 64 349
rect 62 348 63 349
rect 61 348 62 349
rect 60 348 61 349
rect 59 348 60 349
rect 58 348 59 349
rect 57 348 58 349
rect 56 348 57 349
rect 55 348 56 349
rect 54 348 55 349
rect 53 348 54 349
rect 52 348 53 349
rect 51 348 52 349
rect 20 348 21 349
rect 19 348 20 349
rect 18 348 19 349
rect 17 348 18 349
rect 16 348 17 349
rect 15 348 16 349
rect 14 348 15 349
rect 196 349 197 350
rect 195 349 196 350
rect 194 349 195 350
rect 193 349 194 350
rect 192 349 193 350
rect 191 349 192 350
rect 190 349 191 350
rect 189 349 190 350
rect 173 349 174 350
rect 78 349 79 350
rect 77 349 78 350
rect 76 349 77 350
rect 75 349 76 350
rect 74 349 75 350
rect 73 349 74 350
rect 72 349 73 350
rect 71 349 72 350
rect 70 349 71 350
rect 69 349 70 350
rect 68 349 69 350
rect 67 349 68 350
rect 66 349 67 350
rect 65 349 66 350
rect 64 349 65 350
rect 63 349 64 350
rect 62 349 63 350
rect 61 349 62 350
rect 60 349 61 350
rect 59 349 60 350
rect 58 349 59 350
rect 57 349 58 350
rect 56 349 57 350
rect 55 349 56 350
rect 54 349 55 350
rect 53 349 54 350
rect 52 349 53 350
rect 51 349 52 350
rect 29 349 30 350
rect 28 349 29 350
rect 27 349 28 350
rect 26 349 27 350
rect 25 349 26 350
rect 24 349 25 350
rect 23 349 24 350
rect 22 349 23 350
rect 21 349 22 350
rect 20 349 21 350
rect 19 349 20 350
rect 18 349 19 350
rect 17 349 18 350
rect 16 349 17 350
rect 15 349 16 350
rect 14 349 15 350
rect 196 350 197 351
rect 195 350 196 351
rect 194 350 195 351
rect 193 350 194 351
rect 192 350 193 351
rect 191 350 192 351
rect 190 350 191 351
rect 189 350 190 351
rect 174 350 175 351
rect 173 350 174 351
rect 172 350 173 351
rect 78 350 79 351
rect 77 350 78 351
rect 76 350 77 351
rect 75 350 76 351
rect 74 350 75 351
rect 73 350 74 351
rect 72 350 73 351
rect 71 350 72 351
rect 70 350 71 351
rect 69 350 70 351
rect 68 350 69 351
rect 67 350 68 351
rect 66 350 67 351
rect 65 350 66 351
rect 64 350 65 351
rect 63 350 64 351
rect 62 350 63 351
rect 61 350 62 351
rect 60 350 61 351
rect 59 350 60 351
rect 58 350 59 351
rect 57 350 58 351
rect 56 350 57 351
rect 55 350 56 351
rect 54 350 55 351
rect 53 350 54 351
rect 52 350 53 351
rect 51 350 52 351
rect 29 350 30 351
rect 28 350 29 351
rect 27 350 28 351
rect 26 350 27 351
rect 25 350 26 351
rect 24 350 25 351
rect 23 350 24 351
rect 22 350 23 351
rect 21 350 22 351
rect 20 350 21 351
rect 19 350 20 351
rect 18 350 19 351
rect 17 350 18 351
rect 16 350 17 351
rect 15 350 16 351
rect 197 351 198 352
rect 196 351 197 352
rect 192 351 193 352
rect 191 351 192 352
rect 174 351 175 352
rect 173 351 174 352
rect 172 351 173 352
rect 78 351 79 352
rect 77 351 78 352
rect 76 351 77 352
rect 75 351 76 352
rect 74 351 75 352
rect 73 351 74 352
rect 72 351 73 352
rect 71 351 72 352
rect 70 351 71 352
rect 69 351 70 352
rect 68 351 69 352
rect 67 351 68 352
rect 66 351 67 352
rect 65 351 66 352
rect 64 351 65 352
rect 63 351 64 352
rect 62 351 63 352
rect 61 351 62 352
rect 60 351 61 352
rect 59 351 60 352
rect 58 351 59 352
rect 57 351 58 352
rect 56 351 57 352
rect 55 351 56 352
rect 54 351 55 352
rect 53 351 54 352
rect 52 351 53 352
rect 51 351 52 352
rect 29 351 30 352
rect 28 351 29 352
rect 27 351 28 352
rect 26 351 27 352
rect 25 351 26 352
rect 24 351 25 352
rect 196 352 197 353
rect 191 352 192 353
rect 174 352 175 353
rect 173 352 174 353
rect 172 352 173 353
rect 171 352 172 353
rect 67 352 68 353
rect 66 352 67 353
rect 65 352 66 353
rect 64 352 65 353
rect 63 352 64 353
rect 62 352 63 353
rect 55 352 56 353
rect 54 352 55 353
rect 53 352 54 353
rect 52 352 53 353
rect 51 352 52 353
rect 28 352 29 353
rect 27 352 28 353
rect 26 352 27 353
rect 25 352 26 353
rect 24 352 25 353
rect 23 352 24 353
rect 22 352 23 353
rect 196 353 197 354
rect 195 353 196 354
rect 194 353 195 354
rect 193 353 194 354
rect 192 353 193 354
rect 191 353 192 354
rect 189 353 190 354
rect 188 353 189 354
rect 173 353 174 354
rect 172 353 173 354
rect 171 353 172 354
rect 170 353 171 354
rect 66 353 67 354
rect 65 353 66 354
rect 64 353 65 354
rect 63 353 64 354
rect 62 353 63 354
rect 55 353 56 354
rect 54 353 55 354
rect 53 353 54 354
rect 52 353 53 354
rect 51 353 52 354
rect 26 353 27 354
rect 25 353 26 354
rect 24 353 25 354
rect 23 353 24 354
rect 22 353 23 354
rect 21 353 22 354
rect 20 353 21 354
rect 196 354 197 355
rect 195 354 196 355
rect 194 354 195 355
rect 193 354 194 355
rect 192 354 193 355
rect 191 354 192 355
rect 189 354 190 355
rect 188 354 189 355
rect 182 354 183 355
rect 181 354 182 355
rect 180 354 181 355
rect 179 354 180 355
rect 178 354 179 355
rect 177 354 178 355
rect 176 354 177 355
rect 173 354 174 355
rect 172 354 173 355
rect 171 354 172 355
rect 170 354 171 355
rect 169 354 170 355
rect 149 354 150 355
rect 148 354 149 355
rect 147 354 148 355
rect 146 354 147 355
rect 145 354 146 355
rect 144 354 145 355
rect 143 354 144 355
rect 142 354 143 355
rect 141 354 142 355
rect 140 354 141 355
rect 139 354 140 355
rect 138 354 139 355
rect 137 354 138 355
rect 136 354 137 355
rect 135 354 136 355
rect 134 354 135 355
rect 133 354 134 355
rect 132 354 133 355
rect 131 354 132 355
rect 130 354 131 355
rect 129 354 130 355
rect 128 354 129 355
rect 127 354 128 355
rect 126 354 127 355
rect 125 354 126 355
rect 124 354 125 355
rect 123 354 124 355
rect 122 354 123 355
rect 121 354 122 355
rect 120 354 121 355
rect 119 354 120 355
rect 118 354 119 355
rect 117 354 118 355
rect 116 354 117 355
rect 115 354 116 355
rect 114 354 115 355
rect 113 354 114 355
rect 112 354 113 355
rect 111 354 112 355
rect 110 354 111 355
rect 109 354 110 355
rect 108 354 109 355
rect 107 354 108 355
rect 106 354 107 355
rect 105 354 106 355
rect 104 354 105 355
rect 103 354 104 355
rect 102 354 103 355
rect 67 354 68 355
rect 66 354 67 355
rect 65 354 66 355
rect 64 354 65 355
rect 63 354 64 355
rect 62 354 63 355
rect 55 354 56 355
rect 54 354 55 355
rect 53 354 54 355
rect 52 354 53 355
rect 51 354 52 355
rect 24 354 25 355
rect 23 354 24 355
rect 22 354 23 355
rect 21 354 22 355
rect 20 354 21 355
rect 19 354 20 355
rect 18 354 19 355
rect 183 355 184 356
rect 182 355 183 356
rect 181 355 182 356
rect 180 355 181 356
rect 179 355 180 356
rect 178 355 179 356
rect 177 355 178 356
rect 176 355 177 356
rect 172 355 173 356
rect 171 355 172 356
rect 170 355 171 356
rect 169 355 170 356
rect 168 355 169 356
rect 167 355 168 356
rect 166 355 167 356
rect 149 355 150 356
rect 148 355 149 356
rect 147 355 148 356
rect 146 355 147 356
rect 145 355 146 356
rect 144 355 145 356
rect 143 355 144 356
rect 142 355 143 356
rect 141 355 142 356
rect 140 355 141 356
rect 139 355 140 356
rect 138 355 139 356
rect 137 355 138 356
rect 136 355 137 356
rect 135 355 136 356
rect 134 355 135 356
rect 133 355 134 356
rect 132 355 133 356
rect 131 355 132 356
rect 130 355 131 356
rect 129 355 130 356
rect 128 355 129 356
rect 127 355 128 356
rect 126 355 127 356
rect 125 355 126 356
rect 124 355 125 356
rect 123 355 124 356
rect 122 355 123 356
rect 121 355 122 356
rect 120 355 121 356
rect 119 355 120 356
rect 118 355 119 356
rect 117 355 118 356
rect 116 355 117 356
rect 115 355 116 356
rect 114 355 115 356
rect 113 355 114 356
rect 112 355 113 356
rect 111 355 112 356
rect 110 355 111 356
rect 109 355 110 356
rect 108 355 109 356
rect 107 355 108 356
rect 106 355 107 356
rect 105 355 106 356
rect 104 355 105 356
rect 103 355 104 356
rect 102 355 103 356
rect 67 355 68 356
rect 66 355 67 356
rect 65 355 66 356
rect 64 355 65 356
rect 63 355 64 356
rect 62 355 63 356
rect 55 355 56 356
rect 54 355 55 356
rect 53 355 54 356
rect 52 355 53 356
rect 51 355 52 356
rect 29 355 30 356
rect 28 355 29 356
rect 27 355 28 356
rect 21 355 22 356
rect 20 355 21 356
rect 19 355 20 356
rect 18 355 19 356
rect 17 355 18 356
rect 16 355 17 356
rect 196 356 197 357
rect 195 356 196 357
rect 194 356 195 357
rect 193 356 194 357
rect 192 356 193 357
rect 183 356 184 357
rect 182 356 183 357
rect 181 356 182 357
rect 180 356 181 357
rect 179 356 180 357
rect 178 356 179 357
rect 177 356 178 357
rect 176 356 177 357
rect 171 356 172 357
rect 170 356 171 357
rect 169 356 170 357
rect 168 356 169 357
rect 167 356 168 357
rect 166 356 167 357
rect 165 356 166 357
rect 164 356 165 357
rect 163 356 164 357
rect 162 356 163 357
rect 149 356 150 357
rect 148 356 149 357
rect 147 356 148 357
rect 146 356 147 357
rect 145 356 146 357
rect 144 356 145 357
rect 143 356 144 357
rect 142 356 143 357
rect 141 356 142 357
rect 140 356 141 357
rect 139 356 140 357
rect 138 356 139 357
rect 137 356 138 357
rect 136 356 137 357
rect 135 356 136 357
rect 134 356 135 357
rect 133 356 134 357
rect 132 356 133 357
rect 131 356 132 357
rect 130 356 131 357
rect 129 356 130 357
rect 128 356 129 357
rect 127 356 128 357
rect 126 356 127 357
rect 125 356 126 357
rect 124 356 125 357
rect 123 356 124 357
rect 122 356 123 357
rect 121 356 122 357
rect 120 356 121 357
rect 119 356 120 357
rect 118 356 119 357
rect 117 356 118 357
rect 116 356 117 357
rect 115 356 116 357
rect 114 356 115 357
rect 113 356 114 357
rect 112 356 113 357
rect 111 356 112 357
rect 110 356 111 357
rect 109 356 110 357
rect 108 356 109 357
rect 107 356 108 357
rect 106 356 107 357
rect 105 356 106 357
rect 104 356 105 357
rect 103 356 104 357
rect 102 356 103 357
rect 67 356 68 357
rect 66 356 67 357
rect 65 356 66 357
rect 64 356 65 357
rect 63 356 64 357
rect 62 356 63 357
rect 55 356 56 357
rect 54 356 55 357
rect 53 356 54 357
rect 52 356 53 357
rect 51 356 52 357
rect 29 356 30 357
rect 28 356 29 357
rect 27 356 28 357
rect 26 356 27 357
rect 25 356 26 357
rect 24 356 25 357
rect 23 356 24 357
rect 22 356 23 357
rect 20 356 21 357
rect 19 356 20 357
rect 18 356 19 357
rect 17 356 18 357
rect 16 356 17 357
rect 15 356 16 357
rect 196 357 197 358
rect 195 357 196 358
rect 194 357 195 358
rect 193 357 194 358
rect 192 357 193 358
rect 191 357 192 358
rect 183 357 184 358
rect 182 357 183 358
rect 181 357 182 358
rect 180 357 181 358
rect 170 357 171 358
rect 169 357 170 358
rect 168 357 169 358
rect 167 357 168 358
rect 166 357 167 358
rect 165 357 166 358
rect 164 357 165 358
rect 163 357 164 358
rect 162 357 163 358
rect 149 357 150 358
rect 148 357 149 358
rect 147 357 148 358
rect 146 357 147 358
rect 145 357 146 358
rect 144 357 145 358
rect 143 357 144 358
rect 142 357 143 358
rect 141 357 142 358
rect 140 357 141 358
rect 139 357 140 358
rect 138 357 139 358
rect 137 357 138 358
rect 136 357 137 358
rect 135 357 136 358
rect 134 357 135 358
rect 133 357 134 358
rect 132 357 133 358
rect 131 357 132 358
rect 130 357 131 358
rect 129 357 130 358
rect 128 357 129 358
rect 127 357 128 358
rect 126 357 127 358
rect 125 357 126 358
rect 124 357 125 358
rect 123 357 124 358
rect 122 357 123 358
rect 121 357 122 358
rect 120 357 121 358
rect 119 357 120 358
rect 118 357 119 358
rect 117 357 118 358
rect 116 357 117 358
rect 115 357 116 358
rect 114 357 115 358
rect 113 357 114 358
rect 112 357 113 358
rect 111 357 112 358
rect 110 357 111 358
rect 109 357 110 358
rect 108 357 109 358
rect 107 357 108 358
rect 106 357 107 358
rect 105 357 106 358
rect 104 357 105 358
rect 103 357 104 358
rect 102 357 103 358
rect 68 357 69 358
rect 67 357 68 358
rect 66 357 67 358
rect 65 357 66 358
rect 64 357 65 358
rect 63 357 64 358
rect 62 357 63 358
rect 55 357 56 358
rect 54 357 55 358
rect 53 357 54 358
rect 52 357 53 358
rect 51 357 52 358
rect 29 357 30 358
rect 28 357 29 358
rect 27 357 28 358
rect 26 357 27 358
rect 25 357 26 358
rect 24 357 25 358
rect 23 357 24 358
rect 22 357 23 358
rect 21 357 22 358
rect 20 357 21 358
rect 19 357 20 358
rect 18 357 19 358
rect 17 357 18 358
rect 16 357 17 358
rect 15 357 16 358
rect 14 357 15 358
rect 196 358 197 359
rect 192 358 193 359
rect 191 358 192 359
rect 183 358 184 359
rect 182 358 183 359
rect 181 358 182 359
rect 180 358 181 359
rect 171 358 172 359
rect 170 358 171 359
rect 169 358 170 359
rect 168 358 169 359
rect 167 358 168 359
rect 166 358 167 359
rect 165 358 166 359
rect 164 358 165 359
rect 163 358 164 359
rect 162 358 163 359
rect 149 358 150 359
rect 148 358 149 359
rect 147 358 148 359
rect 146 358 147 359
rect 145 358 146 359
rect 144 358 145 359
rect 143 358 144 359
rect 142 358 143 359
rect 141 358 142 359
rect 140 358 141 359
rect 139 358 140 359
rect 138 358 139 359
rect 137 358 138 359
rect 136 358 137 359
rect 135 358 136 359
rect 134 358 135 359
rect 133 358 134 359
rect 132 358 133 359
rect 131 358 132 359
rect 130 358 131 359
rect 129 358 130 359
rect 128 358 129 359
rect 127 358 128 359
rect 126 358 127 359
rect 125 358 126 359
rect 124 358 125 359
rect 123 358 124 359
rect 122 358 123 359
rect 121 358 122 359
rect 120 358 121 359
rect 119 358 120 359
rect 118 358 119 359
rect 117 358 118 359
rect 116 358 117 359
rect 115 358 116 359
rect 114 358 115 359
rect 113 358 114 359
rect 112 358 113 359
rect 111 358 112 359
rect 110 358 111 359
rect 109 358 110 359
rect 108 358 109 359
rect 107 358 108 359
rect 106 358 107 359
rect 105 358 106 359
rect 104 358 105 359
rect 103 358 104 359
rect 102 358 103 359
rect 70 358 71 359
rect 69 358 70 359
rect 68 358 69 359
rect 67 358 68 359
rect 66 358 67 359
rect 65 358 66 359
rect 64 358 65 359
rect 63 358 64 359
rect 62 358 63 359
rect 55 358 56 359
rect 54 358 55 359
rect 53 358 54 359
rect 52 358 53 359
rect 51 358 52 359
rect 26 358 27 359
rect 25 358 26 359
rect 24 358 25 359
rect 23 358 24 359
rect 22 358 23 359
rect 21 358 22 359
rect 20 358 21 359
rect 19 358 20 359
rect 18 358 19 359
rect 17 358 18 359
rect 16 358 17 359
rect 15 358 16 359
rect 14 358 15 359
rect 197 359 198 360
rect 196 359 197 360
rect 192 359 193 360
rect 191 359 192 360
rect 183 359 184 360
rect 182 359 183 360
rect 181 359 182 360
rect 180 359 181 360
rect 171 359 172 360
rect 170 359 171 360
rect 169 359 170 360
rect 168 359 169 360
rect 167 359 168 360
rect 166 359 167 360
rect 165 359 166 360
rect 164 359 165 360
rect 163 359 164 360
rect 162 359 163 360
rect 149 359 150 360
rect 148 359 149 360
rect 147 359 148 360
rect 146 359 147 360
rect 145 359 146 360
rect 144 359 145 360
rect 143 359 144 360
rect 142 359 143 360
rect 141 359 142 360
rect 140 359 141 360
rect 139 359 140 360
rect 138 359 139 360
rect 137 359 138 360
rect 136 359 137 360
rect 135 359 136 360
rect 134 359 135 360
rect 133 359 134 360
rect 132 359 133 360
rect 131 359 132 360
rect 130 359 131 360
rect 129 359 130 360
rect 128 359 129 360
rect 127 359 128 360
rect 126 359 127 360
rect 125 359 126 360
rect 124 359 125 360
rect 123 359 124 360
rect 122 359 123 360
rect 121 359 122 360
rect 120 359 121 360
rect 119 359 120 360
rect 118 359 119 360
rect 117 359 118 360
rect 116 359 117 360
rect 115 359 116 360
rect 114 359 115 360
rect 113 359 114 360
rect 112 359 113 360
rect 111 359 112 360
rect 110 359 111 360
rect 109 359 110 360
rect 108 359 109 360
rect 107 359 108 360
rect 106 359 107 360
rect 105 359 106 360
rect 104 359 105 360
rect 103 359 104 360
rect 102 359 103 360
rect 71 359 72 360
rect 70 359 71 360
rect 69 359 70 360
rect 68 359 69 360
rect 67 359 68 360
rect 66 359 67 360
rect 65 359 66 360
rect 64 359 65 360
rect 63 359 64 360
rect 62 359 63 360
rect 55 359 56 360
rect 54 359 55 360
rect 53 359 54 360
rect 52 359 53 360
rect 51 359 52 360
rect 21 359 22 360
rect 20 359 21 360
rect 19 359 20 360
rect 18 359 19 360
rect 17 359 18 360
rect 16 359 17 360
rect 15 359 16 360
rect 14 359 15 360
rect 196 360 197 361
rect 195 360 196 361
rect 194 360 195 361
rect 193 360 194 361
rect 192 360 193 361
rect 191 360 192 361
rect 183 360 184 361
rect 182 360 183 361
rect 181 360 182 361
rect 180 360 181 361
rect 172 360 173 361
rect 171 360 172 361
rect 170 360 171 361
rect 169 360 170 361
rect 168 360 169 361
rect 149 360 150 361
rect 148 360 149 361
rect 147 360 148 361
rect 146 360 147 361
rect 145 360 146 361
rect 144 360 145 361
rect 143 360 144 361
rect 142 360 143 361
rect 141 360 142 361
rect 140 360 141 361
rect 139 360 140 361
rect 138 360 139 361
rect 137 360 138 361
rect 136 360 137 361
rect 135 360 136 361
rect 134 360 135 361
rect 133 360 134 361
rect 132 360 133 361
rect 131 360 132 361
rect 130 360 131 361
rect 129 360 130 361
rect 128 360 129 361
rect 127 360 128 361
rect 126 360 127 361
rect 125 360 126 361
rect 124 360 125 361
rect 123 360 124 361
rect 122 360 123 361
rect 121 360 122 361
rect 120 360 121 361
rect 119 360 120 361
rect 118 360 119 361
rect 117 360 118 361
rect 116 360 117 361
rect 115 360 116 361
rect 114 360 115 361
rect 113 360 114 361
rect 112 360 113 361
rect 111 360 112 361
rect 110 360 111 361
rect 109 360 110 361
rect 108 360 109 361
rect 107 360 108 361
rect 106 360 107 361
rect 105 360 106 361
rect 104 360 105 361
rect 103 360 104 361
rect 102 360 103 361
rect 73 360 74 361
rect 72 360 73 361
rect 71 360 72 361
rect 70 360 71 361
rect 69 360 70 361
rect 68 360 69 361
rect 67 360 68 361
rect 66 360 67 361
rect 65 360 66 361
rect 64 360 65 361
rect 63 360 64 361
rect 62 360 63 361
rect 56 360 57 361
rect 55 360 56 361
rect 54 360 55 361
rect 53 360 54 361
rect 52 360 53 361
rect 51 360 52 361
rect 15 360 16 361
rect 196 361 197 362
rect 195 361 196 362
rect 194 361 195 362
rect 193 361 194 362
rect 192 361 193 362
rect 191 361 192 362
rect 183 361 184 362
rect 182 361 183 362
rect 181 361 182 362
rect 180 361 181 362
rect 173 361 174 362
rect 172 361 173 362
rect 171 361 172 362
rect 170 361 171 362
rect 169 361 170 362
rect 149 361 150 362
rect 148 361 149 362
rect 147 361 148 362
rect 146 361 147 362
rect 145 361 146 362
rect 144 361 145 362
rect 143 361 144 362
rect 142 361 143 362
rect 141 361 142 362
rect 140 361 141 362
rect 139 361 140 362
rect 138 361 139 362
rect 137 361 138 362
rect 136 361 137 362
rect 135 361 136 362
rect 134 361 135 362
rect 133 361 134 362
rect 132 361 133 362
rect 131 361 132 362
rect 130 361 131 362
rect 129 361 130 362
rect 128 361 129 362
rect 127 361 128 362
rect 126 361 127 362
rect 125 361 126 362
rect 124 361 125 362
rect 123 361 124 362
rect 122 361 123 362
rect 121 361 122 362
rect 120 361 121 362
rect 119 361 120 362
rect 118 361 119 362
rect 117 361 118 362
rect 116 361 117 362
rect 115 361 116 362
rect 114 361 115 362
rect 113 361 114 362
rect 112 361 113 362
rect 111 361 112 362
rect 110 361 111 362
rect 109 361 110 362
rect 108 361 109 362
rect 107 361 108 362
rect 106 361 107 362
rect 105 361 106 362
rect 104 361 105 362
rect 103 361 104 362
rect 102 361 103 362
rect 74 361 75 362
rect 73 361 74 362
rect 72 361 73 362
rect 71 361 72 362
rect 70 361 71 362
rect 69 361 70 362
rect 68 361 69 362
rect 67 361 68 362
rect 66 361 67 362
rect 65 361 66 362
rect 64 361 65 362
rect 63 361 64 362
rect 62 361 63 362
rect 56 361 57 362
rect 55 361 56 362
rect 54 361 55 362
rect 53 361 54 362
rect 52 361 53 362
rect 51 361 52 362
rect 29 361 30 362
rect 28 361 29 362
rect 27 361 28 362
rect 194 362 195 363
rect 183 362 184 363
rect 182 362 183 363
rect 181 362 182 363
rect 180 362 181 363
rect 173 362 174 363
rect 172 362 173 363
rect 171 362 172 363
rect 170 362 171 363
rect 149 362 150 363
rect 148 362 149 363
rect 147 362 148 363
rect 146 362 147 363
rect 145 362 146 363
rect 144 362 145 363
rect 143 362 144 363
rect 142 362 143 363
rect 141 362 142 363
rect 140 362 141 363
rect 139 362 140 363
rect 138 362 139 363
rect 137 362 138 363
rect 136 362 137 363
rect 135 362 136 363
rect 134 362 135 363
rect 133 362 134 363
rect 132 362 133 363
rect 131 362 132 363
rect 130 362 131 363
rect 129 362 130 363
rect 128 362 129 363
rect 127 362 128 363
rect 126 362 127 363
rect 125 362 126 363
rect 124 362 125 363
rect 123 362 124 363
rect 122 362 123 363
rect 121 362 122 363
rect 120 362 121 363
rect 119 362 120 363
rect 118 362 119 363
rect 117 362 118 363
rect 116 362 117 363
rect 115 362 116 363
rect 114 362 115 363
rect 113 362 114 363
rect 112 362 113 363
rect 111 362 112 363
rect 110 362 111 363
rect 109 362 110 363
rect 108 362 109 363
rect 107 362 108 363
rect 106 362 107 363
rect 105 362 106 363
rect 104 362 105 363
rect 103 362 104 363
rect 102 362 103 363
rect 75 362 76 363
rect 74 362 75 363
rect 73 362 74 363
rect 72 362 73 363
rect 71 362 72 363
rect 70 362 71 363
rect 69 362 70 363
rect 68 362 69 363
rect 67 362 68 363
rect 66 362 67 363
rect 65 362 66 363
rect 64 362 65 363
rect 63 362 64 363
rect 62 362 63 363
rect 61 362 62 363
rect 57 362 58 363
rect 56 362 57 363
rect 55 362 56 363
rect 54 362 55 363
rect 53 362 54 363
rect 52 362 53 363
rect 51 362 52 363
rect 29 362 30 363
rect 28 362 29 363
rect 27 362 28 363
rect 26 362 27 363
rect 25 362 26 363
rect 24 362 25 363
rect 23 362 24 363
rect 196 363 197 364
rect 195 363 196 364
rect 193 363 194 364
rect 192 363 193 364
rect 191 363 192 364
rect 183 363 184 364
rect 182 363 183 364
rect 181 363 182 364
rect 180 363 181 364
rect 174 363 175 364
rect 173 363 174 364
rect 172 363 173 364
rect 171 363 172 364
rect 149 363 150 364
rect 148 363 149 364
rect 147 363 148 364
rect 146 363 147 364
rect 145 363 146 364
rect 144 363 145 364
rect 143 363 144 364
rect 142 363 143 364
rect 141 363 142 364
rect 140 363 141 364
rect 139 363 140 364
rect 138 363 139 364
rect 137 363 138 364
rect 136 363 137 364
rect 135 363 136 364
rect 134 363 135 364
rect 133 363 134 364
rect 132 363 133 364
rect 131 363 132 364
rect 130 363 131 364
rect 129 363 130 364
rect 128 363 129 364
rect 127 363 128 364
rect 126 363 127 364
rect 125 363 126 364
rect 124 363 125 364
rect 123 363 124 364
rect 122 363 123 364
rect 121 363 122 364
rect 120 363 121 364
rect 119 363 120 364
rect 118 363 119 364
rect 117 363 118 364
rect 116 363 117 364
rect 115 363 116 364
rect 114 363 115 364
rect 113 363 114 364
rect 112 363 113 364
rect 111 363 112 364
rect 110 363 111 364
rect 109 363 110 364
rect 108 363 109 364
rect 107 363 108 364
rect 106 363 107 364
rect 105 363 106 364
rect 104 363 105 364
rect 103 363 104 364
rect 102 363 103 364
rect 77 363 78 364
rect 76 363 77 364
rect 75 363 76 364
rect 74 363 75 364
rect 73 363 74 364
rect 72 363 73 364
rect 71 363 72 364
rect 70 363 71 364
rect 69 363 70 364
rect 68 363 69 364
rect 65 363 66 364
rect 64 363 65 364
rect 63 363 64 364
rect 62 363 63 364
rect 61 363 62 364
rect 60 363 61 364
rect 59 363 60 364
rect 58 363 59 364
rect 57 363 58 364
rect 56 363 57 364
rect 55 363 56 364
rect 54 363 55 364
rect 53 363 54 364
rect 52 363 53 364
rect 29 363 30 364
rect 28 363 29 364
rect 27 363 28 364
rect 26 363 27 364
rect 25 363 26 364
rect 24 363 25 364
rect 23 363 24 364
rect 22 363 23 364
rect 21 363 22 364
rect 20 363 21 364
rect 19 363 20 364
rect 18 363 19 364
rect 197 364 198 365
rect 196 364 197 365
rect 195 364 196 365
rect 194 364 195 365
rect 193 364 194 365
rect 192 364 193 365
rect 191 364 192 365
rect 183 364 184 365
rect 182 364 183 365
rect 181 364 182 365
rect 180 364 181 365
rect 174 364 175 365
rect 173 364 174 365
rect 172 364 173 365
rect 171 364 172 365
rect 149 364 150 365
rect 148 364 149 365
rect 147 364 148 365
rect 146 364 147 365
rect 145 364 146 365
rect 144 364 145 365
rect 143 364 144 365
rect 142 364 143 365
rect 141 364 142 365
rect 140 364 141 365
rect 139 364 140 365
rect 138 364 139 365
rect 137 364 138 365
rect 136 364 137 365
rect 135 364 136 365
rect 134 364 135 365
rect 133 364 134 365
rect 132 364 133 365
rect 131 364 132 365
rect 130 364 131 365
rect 129 364 130 365
rect 128 364 129 365
rect 127 364 128 365
rect 126 364 127 365
rect 125 364 126 365
rect 124 364 125 365
rect 123 364 124 365
rect 122 364 123 365
rect 121 364 122 365
rect 120 364 121 365
rect 119 364 120 365
rect 118 364 119 365
rect 117 364 118 365
rect 116 364 117 365
rect 115 364 116 365
rect 114 364 115 365
rect 113 364 114 365
rect 112 364 113 365
rect 111 364 112 365
rect 110 364 111 365
rect 109 364 110 365
rect 108 364 109 365
rect 107 364 108 365
rect 106 364 107 365
rect 105 364 106 365
rect 104 364 105 365
rect 103 364 104 365
rect 102 364 103 365
rect 78 364 79 365
rect 77 364 78 365
rect 76 364 77 365
rect 75 364 76 365
rect 74 364 75 365
rect 73 364 74 365
rect 72 364 73 365
rect 71 364 72 365
rect 70 364 71 365
rect 69 364 70 365
rect 65 364 66 365
rect 64 364 65 365
rect 63 364 64 365
rect 62 364 63 365
rect 61 364 62 365
rect 60 364 61 365
rect 59 364 60 365
rect 58 364 59 365
rect 57 364 58 365
rect 56 364 57 365
rect 55 364 56 365
rect 54 364 55 365
rect 53 364 54 365
rect 52 364 53 365
rect 28 364 29 365
rect 27 364 28 365
rect 26 364 27 365
rect 25 364 26 365
rect 24 364 25 365
rect 23 364 24 365
rect 22 364 23 365
rect 21 364 22 365
rect 20 364 21 365
rect 19 364 20 365
rect 18 364 19 365
rect 17 364 18 365
rect 16 364 17 365
rect 15 364 16 365
rect 196 365 197 366
rect 193 365 194 366
rect 192 365 193 366
rect 191 365 192 366
rect 183 365 184 366
rect 182 365 183 366
rect 181 365 182 366
rect 180 365 181 366
rect 172 365 173 366
rect 149 365 150 366
rect 148 365 149 366
rect 147 365 148 366
rect 146 365 147 366
rect 145 365 146 366
rect 144 365 145 366
rect 143 365 144 366
rect 142 365 143 366
rect 141 365 142 366
rect 140 365 141 366
rect 139 365 140 366
rect 138 365 139 366
rect 137 365 138 366
rect 136 365 137 366
rect 135 365 136 366
rect 134 365 135 366
rect 133 365 134 366
rect 132 365 133 366
rect 131 365 132 366
rect 130 365 131 366
rect 129 365 130 366
rect 128 365 129 366
rect 127 365 128 366
rect 126 365 127 366
rect 125 365 126 366
rect 124 365 125 366
rect 123 365 124 366
rect 122 365 123 366
rect 121 365 122 366
rect 120 365 121 366
rect 119 365 120 366
rect 118 365 119 366
rect 117 365 118 366
rect 116 365 117 366
rect 115 365 116 366
rect 114 365 115 366
rect 113 365 114 366
rect 112 365 113 366
rect 111 365 112 366
rect 110 365 111 366
rect 109 365 110 366
rect 108 365 109 366
rect 107 365 108 366
rect 106 365 107 366
rect 105 365 106 366
rect 104 365 105 366
rect 103 365 104 366
rect 102 365 103 366
rect 78 365 79 366
rect 77 365 78 366
rect 76 365 77 366
rect 75 365 76 366
rect 74 365 75 366
rect 73 365 74 366
rect 72 365 73 366
rect 71 365 72 366
rect 70 365 71 366
rect 64 365 65 366
rect 63 365 64 366
rect 62 365 63 366
rect 61 365 62 366
rect 60 365 61 366
rect 59 365 60 366
rect 58 365 59 366
rect 57 365 58 366
rect 56 365 57 366
rect 55 365 56 366
rect 54 365 55 366
rect 53 365 54 366
rect 24 365 25 366
rect 23 365 24 366
rect 22 365 23 366
rect 21 365 22 366
rect 20 365 21 366
rect 19 365 20 366
rect 18 365 19 366
rect 17 365 18 366
rect 16 365 17 366
rect 15 365 16 366
rect 14 365 15 366
rect 192 366 193 367
rect 191 366 192 367
rect 183 366 184 367
rect 182 366 183 367
rect 181 366 182 367
rect 180 366 181 367
rect 149 366 150 367
rect 148 366 149 367
rect 147 366 148 367
rect 146 366 147 367
rect 145 366 146 367
rect 144 366 145 367
rect 143 366 144 367
rect 142 366 143 367
rect 141 366 142 367
rect 140 366 141 367
rect 139 366 140 367
rect 138 366 139 367
rect 137 366 138 367
rect 136 366 137 367
rect 135 366 136 367
rect 134 366 135 367
rect 133 366 134 367
rect 132 366 133 367
rect 131 366 132 367
rect 130 366 131 367
rect 129 366 130 367
rect 128 366 129 367
rect 127 366 128 367
rect 126 366 127 367
rect 125 366 126 367
rect 124 366 125 367
rect 123 366 124 367
rect 122 366 123 367
rect 121 366 122 367
rect 120 366 121 367
rect 119 366 120 367
rect 118 366 119 367
rect 117 366 118 367
rect 116 366 117 367
rect 115 366 116 367
rect 114 366 115 367
rect 113 366 114 367
rect 112 366 113 367
rect 111 366 112 367
rect 110 366 111 367
rect 109 366 110 367
rect 108 366 109 367
rect 107 366 108 367
rect 106 366 107 367
rect 105 366 106 367
rect 104 366 105 367
rect 103 366 104 367
rect 102 366 103 367
rect 78 366 79 367
rect 77 366 78 367
rect 76 366 77 367
rect 75 366 76 367
rect 74 366 75 367
rect 73 366 74 367
rect 72 366 73 367
rect 71 366 72 367
rect 64 366 65 367
rect 63 366 64 367
rect 62 366 63 367
rect 61 366 62 367
rect 60 366 61 367
rect 59 366 60 367
rect 58 366 59 367
rect 57 366 58 367
rect 56 366 57 367
rect 55 366 56 367
rect 54 366 55 367
rect 53 366 54 367
rect 23 366 24 367
rect 22 366 23 367
rect 21 366 22 367
rect 19 366 20 367
rect 18 366 19 367
rect 17 366 18 367
rect 16 366 17 367
rect 15 366 16 367
rect 14 366 15 367
rect 196 367 197 368
rect 195 367 196 368
rect 194 367 195 368
rect 193 367 194 368
rect 192 367 193 368
rect 191 367 192 368
rect 183 367 184 368
rect 182 367 183 368
rect 181 367 182 368
rect 180 367 181 368
rect 149 367 150 368
rect 148 367 149 368
rect 147 367 148 368
rect 146 367 147 368
rect 145 367 146 368
rect 144 367 145 368
rect 143 367 144 368
rect 142 367 143 368
rect 141 367 142 368
rect 140 367 141 368
rect 139 367 140 368
rect 138 367 139 368
rect 137 367 138 368
rect 136 367 137 368
rect 135 367 136 368
rect 134 367 135 368
rect 133 367 134 368
rect 132 367 133 368
rect 131 367 132 368
rect 130 367 131 368
rect 129 367 130 368
rect 128 367 129 368
rect 127 367 128 368
rect 126 367 127 368
rect 125 367 126 368
rect 124 367 125 368
rect 123 367 124 368
rect 122 367 123 368
rect 121 367 122 368
rect 120 367 121 368
rect 119 367 120 368
rect 118 367 119 368
rect 117 367 118 368
rect 116 367 117 368
rect 115 367 116 368
rect 114 367 115 368
rect 113 367 114 368
rect 112 367 113 368
rect 111 367 112 368
rect 110 367 111 368
rect 109 367 110 368
rect 108 367 109 368
rect 107 367 108 368
rect 106 367 107 368
rect 105 367 106 368
rect 104 367 105 368
rect 103 367 104 368
rect 102 367 103 368
rect 78 367 79 368
rect 77 367 78 368
rect 76 367 77 368
rect 75 367 76 368
rect 74 367 75 368
rect 73 367 74 368
rect 63 367 64 368
rect 62 367 63 368
rect 61 367 62 368
rect 60 367 61 368
rect 59 367 60 368
rect 58 367 59 368
rect 57 367 58 368
rect 56 367 57 368
rect 55 367 56 368
rect 54 367 55 368
rect 23 367 24 368
rect 22 367 23 368
rect 21 367 22 368
rect 16 367 17 368
rect 15 367 16 368
rect 14 367 15 368
rect 197 368 198 369
rect 196 368 197 369
rect 195 368 196 369
rect 194 368 195 369
rect 193 368 194 369
rect 192 368 193 369
rect 191 368 192 369
rect 183 368 184 369
rect 182 368 183 369
rect 181 368 182 369
rect 180 368 181 369
rect 177 368 178 369
rect 176 368 177 369
rect 175 368 176 369
rect 174 368 175 369
rect 173 368 174 369
rect 172 368 173 369
rect 171 368 172 369
rect 170 368 171 369
rect 169 368 170 369
rect 168 368 169 369
rect 167 368 168 369
rect 166 368 167 369
rect 165 368 166 369
rect 164 368 165 369
rect 163 368 164 369
rect 162 368 163 369
rect 149 368 150 369
rect 148 368 149 369
rect 147 368 148 369
rect 146 368 147 369
rect 145 368 146 369
rect 144 368 145 369
rect 143 368 144 369
rect 142 368 143 369
rect 141 368 142 369
rect 140 368 141 369
rect 139 368 140 369
rect 138 368 139 369
rect 137 368 138 369
rect 136 368 137 369
rect 135 368 136 369
rect 134 368 135 369
rect 133 368 134 369
rect 132 368 133 369
rect 131 368 132 369
rect 130 368 131 369
rect 129 368 130 369
rect 128 368 129 369
rect 127 368 128 369
rect 126 368 127 369
rect 125 368 126 369
rect 124 368 125 369
rect 123 368 124 369
rect 122 368 123 369
rect 121 368 122 369
rect 120 368 121 369
rect 119 368 120 369
rect 118 368 119 369
rect 117 368 118 369
rect 116 368 117 369
rect 115 368 116 369
rect 114 368 115 369
rect 113 368 114 369
rect 112 368 113 369
rect 111 368 112 369
rect 110 368 111 369
rect 109 368 110 369
rect 108 368 109 369
rect 107 368 108 369
rect 106 368 107 369
rect 105 368 106 369
rect 104 368 105 369
rect 103 368 104 369
rect 102 368 103 369
rect 78 368 79 369
rect 77 368 78 369
rect 76 368 77 369
rect 75 368 76 369
rect 61 368 62 369
rect 60 368 61 369
rect 59 368 60 369
rect 58 368 59 369
rect 57 368 58 369
rect 56 368 57 369
rect 23 368 24 369
rect 22 368 23 369
rect 21 368 22 369
rect 16 368 17 369
rect 15 368 16 369
rect 14 368 15 369
rect 183 369 184 370
rect 182 369 183 370
rect 181 369 182 370
rect 180 369 181 370
rect 177 369 178 370
rect 176 369 177 370
rect 175 369 176 370
rect 174 369 175 370
rect 173 369 174 370
rect 172 369 173 370
rect 171 369 172 370
rect 170 369 171 370
rect 169 369 170 370
rect 168 369 169 370
rect 167 369 168 370
rect 166 369 167 370
rect 165 369 166 370
rect 164 369 165 370
rect 163 369 164 370
rect 162 369 163 370
rect 149 369 150 370
rect 148 369 149 370
rect 147 369 148 370
rect 146 369 147 370
rect 145 369 146 370
rect 144 369 145 370
rect 143 369 144 370
rect 142 369 143 370
rect 141 369 142 370
rect 140 369 141 370
rect 139 369 140 370
rect 138 369 139 370
rect 137 369 138 370
rect 136 369 137 370
rect 135 369 136 370
rect 134 369 135 370
rect 133 369 134 370
rect 132 369 133 370
rect 131 369 132 370
rect 130 369 131 370
rect 129 369 130 370
rect 128 369 129 370
rect 127 369 128 370
rect 126 369 127 370
rect 125 369 126 370
rect 124 369 125 370
rect 123 369 124 370
rect 122 369 123 370
rect 121 369 122 370
rect 120 369 121 370
rect 119 369 120 370
rect 118 369 119 370
rect 117 369 118 370
rect 116 369 117 370
rect 115 369 116 370
rect 114 369 115 370
rect 113 369 114 370
rect 112 369 113 370
rect 111 369 112 370
rect 110 369 111 370
rect 109 369 110 370
rect 108 369 109 370
rect 107 369 108 370
rect 106 369 107 370
rect 105 369 106 370
rect 104 369 105 370
rect 103 369 104 370
rect 102 369 103 370
rect 78 369 79 370
rect 77 369 78 370
rect 76 369 77 370
rect 23 369 24 370
rect 22 369 23 370
rect 21 369 22 370
rect 16 369 17 370
rect 15 369 16 370
rect 14 369 15 370
rect 196 370 197 371
rect 193 370 194 371
rect 192 370 193 371
rect 183 370 184 371
rect 182 370 183 371
rect 181 370 182 371
rect 180 370 181 371
rect 177 370 178 371
rect 176 370 177 371
rect 175 370 176 371
rect 174 370 175 371
rect 173 370 174 371
rect 172 370 173 371
rect 171 370 172 371
rect 170 370 171 371
rect 169 370 170 371
rect 168 370 169 371
rect 167 370 168 371
rect 166 370 167 371
rect 165 370 166 371
rect 164 370 165 371
rect 163 370 164 371
rect 162 370 163 371
rect 149 370 150 371
rect 148 370 149 371
rect 147 370 148 371
rect 146 370 147 371
rect 145 370 146 371
rect 144 370 145 371
rect 143 370 144 371
rect 142 370 143 371
rect 141 370 142 371
rect 140 370 141 371
rect 139 370 140 371
rect 138 370 139 371
rect 137 370 138 371
rect 136 370 137 371
rect 135 370 136 371
rect 134 370 135 371
rect 133 370 134 371
rect 132 370 133 371
rect 131 370 132 371
rect 130 370 131 371
rect 129 370 130 371
rect 128 370 129 371
rect 127 370 128 371
rect 126 370 127 371
rect 125 370 126 371
rect 124 370 125 371
rect 123 370 124 371
rect 122 370 123 371
rect 121 370 122 371
rect 120 370 121 371
rect 119 370 120 371
rect 118 370 119 371
rect 117 370 118 371
rect 116 370 117 371
rect 115 370 116 371
rect 114 370 115 371
rect 113 370 114 371
rect 112 370 113 371
rect 111 370 112 371
rect 110 370 111 371
rect 109 370 110 371
rect 108 370 109 371
rect 107 370 108 371
rect 106 370 107 371
rect 105 370 106 371
rect 104 370 105 371
rect 103 370 104 371
rect 102 370 103 371
rect 78 370 79 371
rect 23 370 24 371
rect 22 370 23 371
rect 21 370 22 371
rect 16 370 17 371
rect 15 370 16 371
rect 14 370 15 371
rect 197 371 198 372
rect 196 371 197 372
rect 194 371 195 372
rect 193 371 194 372
rect 192 371 193 372
rect 191 371 192 372
rect 183 371 184 372
rect 182 371 183 372
rect 181 371 182 372
rect 180 371 181 372
rect 177 371 178 372
rect 176 371 177 372
rect 175 371 176 372
rect 174 371 175 372
rect 173 371 174 372
rect 172 371 173 372
rect 171 371 172 372
rect 170 371 171 372
rect 169 371 170 372
rect 168 371 169 372
rect 167 371 168 372
rect 166 371 167 372
rect 165 371 166 372
rect 164 371 165 372
rect 163 371 164 372
rect 162 371 163 372
rect 149 371 150 372
rect 148 371 149 372
rect 147 371 148 372
rect 146 371 147 372
rect 145 371 146 372
rect 144 371 145 372
rect 143 371 144 372
rect 142 371 143 372
rect 141 371 142 372
rect 140 371 141 372
rect 139 371 140 372
rect 138 371 139 372
rect 137 371 138 372
rect 136 371 137 372
rect 135 371 136 372
rect 134 371 135 372
rect 133 371 134 372
rect 132 371 133 372
rect 131 371 132 372
rect 130 371 131 372
rect 129 371 130 372
rect 128 371 129 372
rect 127 371 128 372
rect 126 371 127 372
rect 125 371 126 372
rect 124 371 125 372
rect 123 371 124 372
rect 122 371 123 372
rect 121 371 122 372
rect 120 371 121 372
rect 119 371 120 372
rect 118 371 119 372
rect 117 371 118 372
rect 116 371 117 372
rect 115 371 116 372
rect 114 371 115 372
rect 113 371 114 372
rect 112 371 113 372
rect 111 371 112 372
rect 110 371 111 372
rect 109 371 110 372
rect 108 371 109 372
rect 107 371 108 372
rect 106 371 107 372
rect 105 371 106 372
rect 104 371 105 372
rect 103 371 104 372
rect 102 371 103 372
rect 23 371 24 372
rect 22 371 23 372
rect 21 371 22 372
rect 20 371 21 372
rect 17 371 18 372
rect 16 371 17 372
rect 15 371 16 372
rect 197 372 198 373
rect 196 372 197 373
rect 195 372 196 373
rect 194 372 195 373
rect 193 372 194 373
rect 192 372 193 373
rect 191 372 192 373
rect 182 372 183 373
rect 181 372 182 373
rect 149 372 150 373
rect 148 372 149 373
rect 147 372 148 373
rect 146 372 147 373
rect 145 372 146 373
rect 144 372 145 373
rect 143 372 144 373
rect 142 372 143 373
rect 141 372 142 373
rect 140 372 141 373
rect 139 372 140 373
rect 138 372 139 373
rect 137 372 138 373
rect 136 372 137 373
rect 135 372 136 373
rect 134 372 135 373
rect 133 372 134 373
rect 132 372 133 373
rect 131 372 132 373
rect 130 372 131 373
rect 129 372 130 373
rect 128 372 129 373
rect 127 372 128 373
rect 126 372 127 373
rect 125 372 126 373
rect 124 372 125 373
rect 123 372 124 373
rect 122 372 123 373
rect 121 372 122 373
rect 120 372 121 373
rect 119 372 120 373
rect 118 372 119 373
rect 117 372 118 373
rect 116 372 117 373
rect 115 372 116 373
rect 114 372 115 373
rect 113 372 114 373
rect 112 372 113 373
rect 111 372 112 373
rect 110 372 111 373
rect 109 372 110 373
rect 108 372 109 373
rect 107 372 108 373
rect 106 372 107 373
rect 105 372 106 373
rect 104 372 105 373
rect 103 372 104 373
rect 102 372 103 373
rect 22 372 23 373
rect 21 372 22 373
rect 20 372 21 373
rect 19 372 20 373
rect 18 372 19 373
rect 17 372 18 373
rect 16 372 17 373
rect 15 372 16 373
rect 196 373 197 374
rect 195 373 196 374
rect 194 373 195 374
rect 192 373 193 374
rect 191 373 192 374
rect 149 373 150 374
rect 148 373 149 374
rect 147 373 148 374
rect 146 373 147 374
rect 145 373 146 374
rect 144 373 145 374
rect 143 373 144 374
rect 142 373 143 374
rect 141 373 142 374
rect 140 373 141 374
rect 139 373 140 374
rect 138 373 139 374
rect 137 373 138 374
rect 136 373 137 374
rect 135 373 136 374
rect 134 373 135 374
rect 133 373 134 374
rect 132 373 133 374
rect 131 373 132 374
rect 130 373 131 374
rect 129 373 130 374
rect 128 373 129 374
rect 127 373 128 374
rect 126 373 127 374
rect 125 373 126 374
rect 124 373 125 374
rect 123 373 124 374
rect 122 373 123 374
rect 121 373 122 374
rect 120 373 121 374
rect 119 373 120 374
rect 118 373 119 374
rect 117 373 118 374
rect 116 373 117 374
rect 115 373 116 374
rect 114 373 115 374
rect 113 373 114 374
rect 112 373 113 374
rect 111 373 112 374
rect 110 373 111 374
rect 109 373 110 374
rect 108 373 109 374
rect 107 373 108 374
rect 106 373 107 374
rect 105 373 106 374
rect 104 373 105 374
rect 103 373 104 374
rect 102 373 103 374
rect 74 373 75 374
rect 73 373 74 374
rect 72 373 73 374
rect 71 373 72 374
rect 70 373 71 374
rect 69 373 70 374
rect 68 373 69 374
rect 67 373 68 374
rect 59 373 60 374
rect 58 373 59 374
rect 57 373 58 374
rect 56 373 57 374
rect 22 373 23 374
rect 21 373 22 374
rect 20 373 21 374
rect 19 373 20 374
rect 18 373 19 374
rect 17 373 18 374
rect 16 373 17 374
rect 15 373 16 374
rect 196 374 197 375
rect 195 374 196 375
rect 194 374 195 375
rect 191 374 192 375
rect 149 374 150 375
rect 148 374 149 375
rect 147 374 148 375
rect 146 374 147 375
rect 145 374 146 375
rect 144 374 145 375
rect 143 374 144 375
rect 142 374 143 375
rect 141 374 142 375
rect 140 374 141 375
rect 139 374 140 375
rect 138 374 139 375
rect 137 374 138 375
rect 136 374 137 375
rect 135 374 136 375
rect 134 374 135 375
rect 133 374 134 375
rect 132 374 133 375
rect 131 374 132 375
rect 130 374 131 375
rect 129 374 130 375
rect 128 374 129 375
rect 127 374 128 375
rect 126 374 127 375
rect 125 374 126 375
rect 124 374 125 375
rect 123 374 124 375
rect 122 374 123 375
rect 121 374 122 375
rect 120 374 121 375
rect 119 374 120 375
rect 118 374 119 375
rect 117 374 118 375
rect 116 374 117 375
rect 115 374 116 375
rect 114 374 115 375
rect 113 374 114 375
rect 112 374 113 375
rect 111 374 112 375
rect 110 374 111 375
rect 109 374 110 375
rect 108 374 109 375
rect 107 374 108 375
rect 106 374 107 375
rect 105 374 106 375
rect 104 374 105 375
rect 103 374 104 375
rect 102 374 103 375
rect 75 374 76 375
rect 74 374 75 375
rect 73 374 74 375
rect 72 374 73 375
rect 71 374 72 375
rect 70 374 71 375
rect 69 374 70 375
rect 68 374 69 375
rect 67 374 68 375
rect 66 374 67 375
rect 61 374 62 375
rect 60 374 61 375
rect 59 374 60 375
rect 58 374 59 375
rect 57 374 58 375
rect 56 374 57 375
rect 55 374 56 375
rect 54 374 55 375
rect 20 374 21 375
rect 19 374 20 375
rect 18 374 19 375
rect 17 374 18 375
rect 16 374 17 375
rect 149 375 150 376
rect 148 375 149 376
rect 147 375 148 376
rect 146 375 147 376
rect 145 375 146 376
rect 144 375 145 376
rect 143 375 144 376
rect 142 375 143 376
rect 141 375 142 376
rect 140 375 141 376
rect 139 375 140 376
rect 138 375 139 376
rect 137 375 138 376
rect 136 375 137 376
rect 135 375 136 376
rect 134 375 135 376
rect 133 375 134 376
rect 132 375 133 376
rect 131 375 132 376
rect 130 375 131 376
rect 129 375 130 376
rect 128 375 129 376
rect 127 375 128 376
rect 126 375 127 376
rect 125 375 126 376
rect 124 375 125 376
rect 123 375 124 376
rect 122 375 123 376
rect 121 375 122 376
rect 120 375 121 376
rect 119 375 120 376
rect 118 375 119 376
rect 117 375 118 376
rect 116 375 117 376
rect 115 375 116 376
rect 114 375 115 376
rect 113 375 114 376
rect 112 375 113 376
rect 111 375 112 376
rect 110 375 111 376
rect 109 375 110 376
rect 108 375 109 376
rect 107 375 108 376
rect 106 375 107 376
rect 105 375 106 376
rect 104 375 105 376
rect 103 375 104 376
rect 102 375 103 376
rect 76 375 77 376
rect 75 375 76 376
rect 74 375 75 376
rect 73 375 74 376
rect 72 375 73 376
rect 71 375 72 376
rect 70 375 71 376
rect 69 375 70 376
rect 68 375 69 376
rect 67 375 68 376
rect 66 375 67 376
rect 65 375 66 376
rect 62 375 63 376
rect 61 375 62 376
rect 60 375 61 376
rect 59 375 60 376
rect 58 375 59 376
rect 57 375 58 376
rect 56 375 57 376
rect 55 375 56 376
rect 54 375 55 376
rect 53 375 54 376
rect 149 376 150 377
rect 148 376 149 377
rect 147 376 148 377
rect 146 376 147 377
rect 145 376 146 377
rect 144 376 145 377
rect 143 376 144 377
rect 142 376 143 377
rect 141 376 142 377
rect 140 376 141 377
rect 139 376 140 377
rect 138 376 139 377
rect 137 376 138 377
rect 136 376 137 377
rect 135 376 136 377
rect 134 376 135 377
rect 133 376 134 377
rect 132 376 133 377
rect 131 376 132 377
rect 130 376 131 377
rect 129 376 130 377
rect 128 376 129 377
rect 127 376 128 377
rect 126 376 127 377
rect 125 376 126 377
rect 124 376 125 377
rect 123 376 124 377
rect 122 376 123 377
rect 121 376 122 377
rect 120 376 121 377
rect 119 376 120 377
rect 118 376 119 377
rect 117 376 118 377
rect 116 376 117 377
rect 115 376 116 377
rect 114 376 115 377
rect 113 376 114 377
rect 112 376 113 377
rect 111 376 112 377
rect 110 376 111 377
rect 109 376 110 377
rect 108 376 109 377
rect 107 376 108 377
rect 106 376 107 377
rect 105 376 106 377
rect 104 376 105 377
rect 103 376 104 377
rect 102 376 103 377
rect 77 376 78 377
rect 76 376 77 377
rect 75 376 76 377
rect 74 376 75 377
rect 73 376 74 377
rect 72 376 73 377
rect 71 376 72 377
rect 70 376 71 377
rect 69 376 70 377
rect 68 376 69 377
rect 67 376 68 377
rect 66 376 67 377
rect 65 376 66 377
rect 64 376 65 377
rect 63 376 64 377
rect 62 376 63 377
rect 61 376 62 377
rect 60 376 61 377
rect 59 376 60 377
rect 58 376 59 377
rect 57 376 58 377
rect 56 376 57 377
rect 55 376 56 377
rect 54 376 55 377
rect 53 376 54 377
rect 52 376 53 377
rect 149 377 150 378
rect 148 377 149 378
rect 147 377 148 378
rect 146 377 147 378
rect 145 377 146 378
rect 144 377 145 378
rect 143 377 144 378
rect 142 377 143 378
rect 141 377 142 378
rect 140 377 141 378
rect 139 377 140 378
rect 138 377 139 378
rect 137 377 138 378
rect 136 377 137 378
rect 135 377 136 378
rect 134 377 135 378
rect 133 377 134 378
rect 132 377 133 378
rect 131 377 132 378
rect 130 377 131 378
rect 129 377 130 378
rect 128 377 129 378
rect 127 377 128 378
rect 126 377 127 378
rect 125 377 126 378
rect 124 377 125 378
rect 123 377 124 378
rect 122 377 123 378
rect 121 377 122 378
rect 120 377 121 378
rect 119 377 120 378
rect 118 377 119 378
rect 117 377 118 378
rect 116 377 117 378
rect 115 377 116 378
rect 114 377 115 378
rect 113 377 114 378
rect 112 377 113 378
rect 111 377 112 378
rect 110 377 111 378
rect 109 377 110 378
rect 108 377 109 378
rect 107 377 108 378
rect 106 377 107 378
rect 105 377 106 378
rect 104 377 105 378
rect 103 377 104 378
rect 102 377 103 378
rect 78 377 79 378
rect 77 377 78 378
rect 76 377 77 378
rect 75 377 76 378
rect 74 377 75 378
rect 73 377 74 378
rect 72 377 73 378
rect 71 377 72 378
rect 70 377 71 378
rect 69 377 70 378
rect 68 377 69 378
rect 67 377 68 378
rect 66 377 67 378
rect 65 377 66 378
rect 64 377 65 378
rect 63 377 64 378
rect 62 377 63 378
rect 61 377 62 378
rect 60 377 61 378
rect 59 377 60 378
rect 58 377 59 378
rect 57 377 58 378
rect 56 377 57 378
rect 55 377 56 378
rect 54 377 55 378
rect 53 377 54 378
rect 52 377 53 378
rect 29 377 30 378
rect 28 377 29 378
rect 27 377 28 378
rect 26 377 27 378
rect 25 377 26 378
rect 24 377 25 378
rect 23 377 24 378
rect 22 377 23 378
rect 21 377 22 378
rect 20 377 21 378
rect 19 377 20 378
rect 18 377 19 378
rect 17 377 18 378
rect 16 377 17 378
rect 15 377 16 378
rect 14 377 15 378
rect 112 378 113 379
rect 111 378 112 379
rect 110 378 111 379
rect 109 378 110 379
rect 108 378 109 379
rect 107 378 108 379
rect 106 378 107 379
rect 105 378 106 379
rect 104 378 105 379
rect 103 378 104 379
rect 102 378 103 379
rect 78 378 79 379
rect 77 378 78 379
rect 76 378 77 379
rect 75 378 76 379
rect 74 378 75 379
rect 73 378 74 379
rect 67 378 68 379
rect 66 378 67 379
rect 65 378 66 379
rect 64 378 65 379
rect 63 378 64 379
rect 62 378 63 379
rect 61 378 62 379
rect 60 378 61 379
rect 59 378 60 379
rect 58 378 59 379
rect 57 378 58 379
rect 56 378 57 379
rect 55 378 56 379
rect 54 378 55 379
rect 53 378 54 379
rect 52 378 53 379
rect 29 378 30 379
rect 28 378 29 379
rect 27 378 28 379
rect 26 378 27 379
rect 25 378 26 379
rect 24 378 25 379
rect 23 378 24 379
rect 22 378 23 379
rect 21 378 22 379
rect 20 378 21 379
rect 19 378 20 379
rect 18 378 19 379
rect 17 378 18 379
rect 16 378 17 379
rect 15 378 16 379
rect 14 378 15 379
rect 197 379 198 380
rect 196 379 197 380
rect 195 379 196 380
rect 194 379 195 380
rect 193 379 194 380
rect 192 379 193 380
rect 191 379 192 380
rect 190 379 191 380
rect 189 379 190 380
rect 112 379 113 380
rect 111 379 112 380
rect 110 379 111 380
rect 109 379 110 380
rect 108 379 109 380
rect 107 379 108 380
rect 106 379 107 380
rect 105 379 106 380
rect 104 379 105 380
rect 103 379 104 380
rect 102 379 103 380
rect 78 379 79 380
rect 77 379 78 380
rect 76 379 77 380
rect 75 379 76 380
rect 74 379 75 380
rect 66 379 67 380
rect 65 379 66 380
rect 64 379 65 380
rect 63 379 64 380
rect 62 379 63 380
rect 61 379 62 380
rect 55 379 56 380
rect 54 379 55 380
rect 53 379 54 380
rect 52 379 53 380
rect 51 379 52 380
rect 29 379 30 380
rect 28 379 29 380
rect 27 379 28 380
rect 26 379 27 380
rect 25 379 26 380
rect 24 379 25 380
rect 23 379 24 380
rect 22 379 23 380
rect 21 379 22 380
rect 20 379 21 380
rect 19 379 20 380
rect 18 379 19 380
rect 17 379 18 380
rect 16 379 17 380
rect 15 379 16 380
rect 196 380 197 381
rect 195 380 196 381
rect 194 380 195 381
rect 193 380 194 381
rect 192 380 193 381
rect 191 380 192 381
rect 190 380 191 381
rect 189 380 190 381
rect 112 380 113 381
rect 111 380 112 381
rect 110 380 111 381
rect 109 380 110 381
rect 108 380 109 381
rect 107 380 108 381
rect 106 380 107 381
rect 105 380 106 381
rect 104 380 105 381
rect 103 380 104 381
rect 102 380 103 381
rect 78 380 79 381
rect 77 380 78 381
rect 76 380 77 381
rect 75 380 76 381
rect 65 380 66 381
rect 64 380 65 381
rect 63 380 64 381
rect 62 380 63 381
rect 55 380 56 381
rect 54 380 55 381
rect 53 380 54 381
rect 52 380 53 381
rect 51 380 52 381
rect 29 380 30 381
rect 28 380 29 381
rect 27 380 28 381
rect 26 380 27 381
rect 25 380 26 381
rect 24 380 25 381
rect 193 381 194 382
rect 192 381 193 382
rect 189 381 190 382
rect 112 381 113 382
rect 111 381 112 382
rect 110 381 111 382
rect 109 381 110 382
rect 108 381 109 382
rect 107 381 108 382
rect 106 381 107 382
rect 105 381 106 382
rect 104 381 105 382
rect 103 381 104 382
rect 102 381 103 382
rect 78 381 79 382
rect 77 381 78 382
rect 76 381 77 382
rect 75 381 76 382
rect 65 381 66 382
rect 64 381 65 382
rect 63 381 64 382
rect 62 381 63 382
rect 55 381 56 382
rect 54 381 55 382
rect 53 381 54 382
rect 52 381 53 382
rect 51 381 52 382
rect 28 381 29 382
rect 27 381 28 382
rect 26 381 27 382
rect 25 381 26 382
rect 24 381 25 382
rect 23 381 24 382
rect 22 381 23 382
rect 194 382 195 383
rect 193 382 194 383
rect 192 382 193 383
rect 190 382 191 383
rect 189 382 190 383
rect 112 382 113 383
rect 111 382 112 383
rect 110 382 111 383
rect 109 382 110 383
rect 108 382 109 383
rect 107 382 108 383
rect 106 382 107 383
rect 105 382 106 383
rect 104 382 105 383
rect 103 382 104 383
rect 102 382 103 383
rect 78 382 79 383
rect 77 382 78 383
rect 76 382 77 383
rect 75 382 76 383
rect 65 382 66 383
rect 64 382 65 383
rect 63 382 64 383
rect 62 382 63 383
rect 55 382 56 383
rect 54 382 55 383
rect 53 382 54 383
rect 52 382 53 383
rect 51 382 52 383
rect 26 382 27 383
rect 25 382 26 383
rect 24 382 25 383
rect 23 382 24 383
rect 22 382 23 383
rect 21 382 22 383
rect 20 382 21 383
rect 196 383 197 384
rect 195 383 196 384
rect 194 383 195 384
rect 193 383 194 384
rect 192 383 193 384
rect 191 383 192 384
rect 190 383 191 384
rect 189 383 190 384
rect 112 383 113 384
rect 111 383 112 384
rect 110 383 111 384
rect 109 383 110 384
rect 108 383 109 384
rect 107 383 108 384
rect 106 383 107 384
rect 105 383 106 384
rect 104 383 105 384
rect 103 383 104 384
rect 102 383 103 384
rect 78 383 79 384
rect 77 383 78 384
rect 76 383 77 384
rect 75 383 76 384
rect 66 383 67 384
rect 65 383 66 384
rect 64 383 65 384
rect 63 383 64 384
rect 62 383 63 384
rect 61 383 62 384
rect 55 383 56 384
rect 54 383 55 384
rect 53 383 54 384
rect 52 383 53 384
rect 51 383 52 384
rect 24 383 25 384
rect 23 383 24 384
rect 22 383 23 384
rect 21 383 22 384
rect 20 383 21 384
rect 19 383 20 384
rect 18 383 19 384
rect 196 384 197 385
rect 195 384 196 385
rect 194 384 195 385
rect 192 384 193 385
rect 191 384 192 385
rect 190 384 191 385
rect 189 384 190 385
rect 112 384 113 385
rect 111 384 112 385
rect 110 384 111 385
rect 109 384 110 385
rect 108 384 109 385
rect 107 384 108 385
rect 106 384 107 385
rect 105 384 106 385
rect 104 384 105 385
rect 103 384 104 385
rect 102 384 103 385
rect 78 384 79 385
rect 77 384 78 385
rect 76 384 77 385
rect 75 384 76 385
rect 74 384 75 385
rect 67 384 68 385
rect 66 384 67 385
rect 65 384 66 385
rect 64 384 65 385
rect 63 384 64 385
rect 62 384 63 385
rect 61 384 62 385
rect 60 384 61 385
rect 56 384 57 385
rect 55 384 56 385
rect 54 384 55 385
rect 53 384 54 385
rect 52 384 53 385
rect 51 384 52 385
rect 22 384 23 385
rect 21 384 22 385
rect 20 384 21 385
rect 19 384 20 385
rect 18 384 19 385
rect 17 384 18 385
rect 16 384 17 385
rect 196 385 197 386
rect 194 385 195 386
rect 170 385 171 386
rect 169 385 170 386
rect 168 385 169 386
rect 167 385 168 386
rect 166 385 167 386
rect 165 385 166 386
rect 112 385 113 386
rect 111 385 112 386
rect 110 385 111 386
rect 109 385 110 386
rect 108 385 109 386
rect 107 385 108 386
rect 106 385 107 386
rect 105 385 106 386
rect 104 385 105 386
rect 103 385 104 386
rect 102 385 103 386
rect 78 385 79 386
rect 77 385 78 386
rect 76 385 77 386
rect 75 385 76 386
rect 74 385 75 386
rect 73 385 74 386
rect 72 385 73 386
rect 71 385 72 386
rect 70 385 71 386
rect 69 385 70 386
rect 68 385 69 386
rect 67 385 68 386
rect 66 385 67 386
rect 65 385 66 386
rect 64 385 65 386
rect 63 385 64 386
rect 62 385 63 386
rect 61 385 62 386
rect 60 385 61 386
rect 59 385 60 386
rect 58 385 59 386
rect 57 385 58 386
rect 56 385 57 386
rect 55 385 56 386
rect 54 385 55 386
rect 53 385 54 386
rect 52 385 53 386
rect 19 385 20 386
rect 18 385 19 386
rect 17 385 18 386
rect 16 385 17 386
rect 15 385 16 386
rect 196 386 197 387
rect 195 386 196 387
rect 194 386 195 387
rect 193 386 194 387
rect 192 386 193 387
rect 171 386 172 387
rect 170 386 171 387
rect 169 386 170 387
rect 168 386 169 387
rect 167 386 168 387
rect 166 386 167 387
rect 165 386 166 387
rect 164 386 165 387
rect 128 386 129 387
rect 112 386 113 387
rect 111 386 112 387
rect 110 386 111 387
rect 109 386 110 387
rect 108 386 109 387
rect 107 386 108 387
rect 106 386 107 387
rect 105 386 106 387
rect 104 386 105 387
rect 103 386 104 387
rect 102 386 103 387
rect 77 386 78 387
rect 76 386 77 387
rect 75 386 76 387
rect 74 386 75 387
rect 73 386 74 387
rect 72 386 73 387
rect 71 386 72 387
rect 70 386 71 387
rect 69 386 70 387
rect 68 386 69 387
rect 67 386 68 387
rect 66 386 67 387
rect 65 386 66 387
rect 64 386 65 387
rect 63 386 64 387
rect 62 386 63 387
rect 61 386 62 387
rect 60 386 61 387
rect 59 386 60 387
rect 58 386 59 387
rect 57 386 58 387
rect 56 386 57 387
rect 55 386 56 387
rect 54 386 55 387
rect 53 386 54 387
rect 52 386 53 387
rect 29 386 30 387
rect 28 386 29 387
rect 27 386 28 387
rect 26 386 27 387
rect 25 386 26 387
rect 24 386 25 387
rect 23 386 24 387
rect 22 386 23 387
rect 21 386 22 387
rect 20 386 21 387
rect 19 386 20 387
rect 18 386 19 387
rect 17 386 18 387
rect 16 386 17 387
rect 15 386 16 387
rect 14 386 15 387
rect 196 387 197 388
rect 195 387 196 388
rect 194 387 195 388
rect 193 387 194 388
rect 192 387 193 388
rect 191 387 192 388
rect 172 387 173 388
rect 171 387 172 388
rect 170 387 171 388
rect 169 387 170 388
rect 168 387 169 388
rect 167 387 168 388
rect 166 387 167 388
rect 165 387 166 388
rect 164 387 165 388
rect 163 387 164 388
rect 129 387 130 388
rect 128 387 129 388
rect 127 387 128 388
rect 112 387 113 388
rect 111 387 112 388
rect 110 387 111 388
rect 109 387 110 388
rect 108 387 109 388
rect 107 387 108 388
rect 106 387 107 388
rect 105 387 106 388
rect 104 387 105 388
rect 103 387 104 388
rect 102 387 103 388
rect 77 387 78 388
rect 76 387 77 388
rect 75 387 76 388
rect 74 387 75 388
rect 73 387 74 388
rect 72 387 73 388
rect 71 387 72 388
rect 70 387 71 388
rect 69 387 70 388
rect 68 387 69 388
rect 67 387 68 388
rect 66 387 67 388
rect 65 387 66 388
rect 62 387 63 388
rect 61 387 62 388
rect 60 387 61 388
rect 59 387 60 388
rect 58 387 59 388
rect 57 387 58 388
rect 56 387 57 388
rect 55 387 56 388
rect 54 387 55 388
rect 53 387 54 388
rect 29 387 30 388
rect 28 387 29 388
rect 27 387 28 388
rect 26 387 27 388
rect 25 387 26 388
rect 24 387 25 388
rect 23 387 24 388
rect 22 387 23 388
rect 21 387 22 388
rect 20 387 21 388
rect 19 387 20 388
rect 18 387 19 388
rect 17 387 18 388
rect 16 387 17 388
rect 15 387 16 388
rect 14 387 15 388
rect 197 388 198 389
rect 196 388 197 389
rect 194 388 195 389
rect 192 388 193 389
rect 191 388 192 389
rect 183 388 184 389
rect 182 388 183 389
rect 181 388 182 389
rect 180 388 181 389
rect 179 388 180 389
rect 178 388 179 389
rect 177 388 178 389
rect 176 388 177 389
rect 173 388 174 389
rect 172 388 173 389
rect 171 388 172 389
rect 170 388 171 389
rect 169 388 170 389
rect 166 388 167 389
rect 165 388 166 389
rect 164 388 165 389
rect 163 388 164 389
rect 130 388 131 389
rect 129 388 130 389
rect 128 388 129 389
rect 127 388 128 389
rect 112 388 113 389
rect 111 388 112 389
rect 110 388 111 389
rect 109 388 110 389
rect 108 388 109 389
rect 107 388 108 389
rect 106 388 107 389
rect 105 388 106 389
rect 104 388 105 389
rect 103 388 104 389
rect 102 388 103 389
rect 76 388 77 389
rect 75 388 76 389
rect 74 388 75 389
rect 73 388 74 389
rect 72 388 73 389
rect 71 388 72 389
rect 70 388 71 389
rect 69 388 70 389
rect 68 388 69 389
rect 67 388 68 389
rect 66 388 67 389
rect 65 388 66 389
rect 61 388 62 389
rect 60 388 61 389
rect 59 388 60 389
rect 58 388 59 389
rect 57 388 58 389
rect 56 388 57 389
rect 55 388 56 389
rect 54 388 55 389
rect 29 388 30 389
rect 28 388 29 389
rect 27 388 28 389
rect 26 388 27 389
rect 25 388 26 389
rect 24 388 25 389
rect 23 388 24 389
rect 22 388 23 389
rect 21 388 22 389
rect 20 388 21 389
rect 19 388 20 389
rect 18 388 19 389
rect 17 388 18 389
rect 16 388 17 389
rect 15 388 16 389
rect 197 389 198 390
rect 196 389 197 390
rect 194 389 195 390
rect 192 389 193 390
rect 191 389 192 390
rect 183 389 184 390
rect 182 389 183 390
rect 181 389 182 390
rect 180 389 181 390
rect 179 389 180 390
rect 178 389 179 390
rect 177 389 178 390
rect 176 389 177 390
rect 173 389 174 390
rect 172 389 173 390
rect 171 389 172 390
rect 170 389 171 390
rect 165 389 166 390
rect 164 389 165 390
rect 163 389 164 390
rect 131 389 132 390
rect 130 389 131 390
rect 129 389 130 390
rect 128 389 129 390
rect 127 389 128 390
rect 112 389 113 390
rect 111 389 112 390
rect 110 389 111 390
rect 109 389 110 390
rect 108 389 109 390
rect 107 389 108 390
rect 106 389 107 390
rect 105 389 106 390
rect 104 389 105 390
rect 103 389 104 390
rect 102 389 103 390
rect 75 389 76 390
rect 74 389 75 390
rect 73 389 74 390
rect 72 389 73 390
rect 71 389 72 390
rect 70 389 71 390
rect 69 389 70 390
rect 68 389 69 390
rect 67 389 68 390
rect 66 389 67 390
rect 60 389 61 390
rect 59 389 60 390
rect 58 389 59 390
rect 57 389 58 390
rect 56 389 57 390
rect 29 389 30 390
rect 28 389 29 390
rect 27 389 28 390
rect 26 389 27 390
rect 25 389 26 390
rect 24 389 25 390
rect 197 390 198 391
rect 196 390 197 391
rect 194 390 195 391
rect 193 390 194 391
rect 192 390 193 391
rect 191 390 192 391
rect 183 390 184 391
rect 182 390 183 391
rect 181 390 182 391
rect 180 390 181 391
rect 179 390 180 391
rect 178 390 179 391
rect 177 390 178 391
rect 176 390 177 391
rect 173 390 174 391
rect 172 390 173 391
rect 171 390 172 391
rect 165 390 166 391
rect 164 390 165 391
rect 163 390 164 391
rect 162 390 163 391
rect 131 390 132 391
rect 130 390 131 391
rect 129 390 130 391
rect 128 390 129 391
rect 127 390 128 391
rect 112 390 113 391
rect 111 390 112 391
rect 110 390 111 391
rect 109 390 110 391
rect 108 390 109 391
rect 107 390 108 391
rect 106 390 107 391
rect 105 390 106 391
rect 104 390 105 391
rect 103 390 104 391
rect 102 390 103 391
rect 73 390 74 391
rect 72 390 73 391
rect 71 390 72 391
rect 70 390 71 391
rect 69 390 70 391
rect 68 390 69 391
rect 27 390 28 391
rect 26 390 27 391
rect 25 390 26 391
rect 24 390 25 391
rect 23 390 24 391
rect 22 390 23 391
rect 196 391 197 392
rect 194 391 195 392
rect 193 391 194 392
rect 192 391 193 392
rect 183 391 184 392
rect 182 391 183 392
rect 181 391 182 392
rect 180 391 181 392
rect 179 391 180 392
rect 178 391 179 392
rect 177 391 178 392
rect 176 391 177 392
rect 173 391 174 392
rect 172 391 173 392
rect 171 391 172 392
rect 164 391 165 392
rect 163 391 164 392
rect 162 391 163 392
rect 132 391 133 392
rect 131 391 132 392
rect 130 391 131 392
rect 129 391 130 392
rect 128 391 129 392
rect 127 391 128 392
rect 112 391 113 392
rect 111 391 112 392
rect 110 391 111 392
rect 109 391 110 392
rect 108 391 109 392
rect 107 391 108 392
rect 106 391 107 392
rect 105 391 106 392
rect 104 391 105 392
rect 103 391 104 392
rect 102 391 103 392
rect 25 391 26 392
rect 24 391 25 392
rect 23 391 24 392
rect 22 391 23 392
rect 21 391 22 392
rect 20 391 21 392
rect 196 392 197 393
rect 193 392 194 393
rect 183 392 184 393
rect 182 392 183 393
rect 181 392 182 393
rect 180 392 181 393
rect 173 392 174 393
rect 172 392 173 393
rect 171 392 172 393
rect 165 392 166 393
rect 164 392 165 393
rect 163 392 164 393
rect 162 392 163 393
rect 133 392 134 393
rect 132 392 133 393
rect 131 392 132 393
rect 130 392 131 393
rect 129 392 130 393
rect 128 392 129 393
rect 127 392 128 393
rect 112 392 113 393
rect 111 392 112 393
rect 110 392 111 393
rect 109 392 110 393
rect 108 392 109 393
rect 107 392 108 393
rect 106 392 107 393
rect 105 392 106 393
rect 104 392 105 393
rect 103 392 104 393
rect 102 392 103 393
rect 23 392 24 393
rect 22 392 23 393
rect 21 392 22 393
rect 20 392 21 393
rect 19 392 20 393
rect 18 392 19 393
rect 17 392 18 393
rect 197 393 198 394
rect 196 393 197 394
rect 194 393 195 394
rect 193 393 194 394
rect 192 393 193 394
rect 191 393 192 394
rect 183 393 184 394
rect 182 393 183 394
rect 181 393 182 394
rect 180 393 181 394
rect 173 393 174 394
rect 172 393 173 394
rect 171 393 172 394
rect 170 393 171 394
rect 165 393 166 394
rect 164 393 165 394
rect 163 393 164 394
rect 134 393 135 394
rect 133 393 134 394
rect 132 393 133 394
rect 131 393 132 394
rect 130 393 131 394
rect 129 393 130 394
rect 128 393 129 394
rect 127 393 128 394
rect 112 393 113 394
rect 111 393 112 394
rect 110 393 111 394
rect 109 393 110 394
rect 108 393 109 394
rect 107 393 108 394
rect 106 393 107 394
rect 105 393 106 394
rect 104 393 105 394
rect 103 393 104 394
rect 102 393 103 394
rect 21 393 22 394
rect 20 393 21 394
rect 19 393 20 394
rect 18 393 19 394
rect 17 393 18 394
rect 16 393 17 394
rect 15 393 16 394
rect 197 394 198 395
rect 196 394 197 395
rect 194 394 195 395
rect 193 394 194 395
rect 192 394 193 395
rect 191 394 192 395
rect 183 394 184 395
rect 182 394 183 395
rect 181 394 182 395
rect 180 394 181 395
rect 173 394 174 395
rect 172 394 173 395
rect 171 394 172 395
rect 170 394 171 395
rect 169 394 170 395
rect 166 394 167 395
rect 165 394 166 395
rect 164 394 165 395
rect 163 394 164 395
rect 135 394 136 395
rect 134 394 135 395
rect 133 394 134 395
rect 132 394 133 395
rect 131 394 132 395
rect 130 394 131 395
rect 129 394 130 395
rect 128 394 129 395
rect 127 394 128 395
rect 112 394 113 395
rect 111 394 112 395
rect 110 394 111 395
rect 109 394 110 395
rect 108 394 109 395
rect 107 394 108 395
rect 106 394 107 395
rect 105 394 106 395
rect 104 394 105 395
rect 103 394 104 395
rect 102 394 103 395
rect 86 394 87 395
rect 85 394 86 395
rect 84 394 85 395
rect 53 394 54 395
rect 52 394 53 395
rect 51 394 52 395
rect 19 394 20 395
rect 18 394 19 395
rect 17 394 18 395
rect 16 394 17 395
rect 15 394 16 395
rect 14 394 15 395
rect 197 395 198 396
rect 196 395 197 396
rect 195 395 196 396
rect 194 395 195 396
rect 192 395 193 396
rect 191 395 192 396
rect 183 395 184 396
rect 182 395 183 396
rect 181 395 182 396
rect 180 395 181 396
rect 172 395 173 396
rect 171 395 172 396
rect 170 395 171 396
rect 169 395 170 396
rect 168 395 169 396
rect 167 395 168 396
rect 166 395 167 396
rect 165 395 166 396
rect 164 395 165 396
rect 163 395 164 396
rect 136 395 137 396
rect 135 395 136 396
rect 134 395 135 396
rect 133 395 134 396
rect 132 395 133 396
rect 131 395 132 396
rect 130 395 131 396
rect 129 395 130 396
rect 128 395 129 396
rect 127 395 128 396
rect 112 395 113 396
rect 111 395 112 396
rect 110 395 111 396
rect 109 395 110 396
rect 108 395 109 396
rect 107 395 108 396
rect 106 395 107 396
rect 105 395 106 396
rect 104 395 105 396
rect 103 395 104 396
rect 102 395 103 396
rect 86 395 87 396
rect 85 395 86 396
rect 84 395 85 396
rect 83 395 84 396
rect 82 395 83 396
rect 55 395 56 396
rect 54 395 55 396
rect 53 395 54 396
rect 52 395 53 396
rect 51 395 52 396
rect 17 395 18 396
rect 16 395 17 396
rect 15 395 16 396
rect 14 395 15 396
rect 196 396 197 397
rect 195 396 196 397
rect 194 396 195 397
rect 191 396 192 397
rect 183 396 184 397
rect 182 396 183 397
rect 181 396 182 397
rect 180 396 181 397
rect 172 396 173 397
rect 171 396 172 397
rect 170 396 171 397
rect 169 396 170 397
rect 168 396 169 397
rect 167 396 168 397
rect 166 396 167 397
rect 165 396 166 397
rect 164 396 165 397
rect 136 396 137 397
rect 135 396 136 397
rect 134 396 135 397
rect 133 396 134 397
rect 132 396 133 397
rect 131 396 132 397
rect 130 396 131 397
rect 129 396 130 397
rect 128 396 129 397
rect 127 396 128 397
rect 112 396 113 397
rect 111 396 112 397
rect 110 396 111 397
rect 109 396 110 397
rect 108 396 109 397
rect 107 396 108 397
rect 106 396 107 397
rect 105 396 106 397
rect 104 396 105 397
rect 103 396 104 397
rect 102 396 103 397
rect 86 396 87 397
rect 85 396 86 397
rect 84 396 85 397
rect 83 396 84 397
rect 82 396 83 397
rect 81 396 82 397
rect 80 396 81 397
rect 79 396 80 397
rect 58 396 59 397
rect 57 396 58 397
rect 56 396 57 397
rect 55 396 56 397
rect 54 396 55 397
rect 53 396 54 397
rect 52 396 53 397
rect 51 396 52 397
rect 15 396 16 397
rect 195 397 196 398
rect 194 397 195 398
rect 193 397 194 398
rect 183 397 184 398
rect 182 397 183 398
rect 181 397 182 398
rect 180 397 181 398
rect 171 397 172 398
rect 170 397 171 398
rect 169 397 170 398
rect 168 397 169 398
rect 167 397 168 398
rect 166 397 167 398
rect 165 397 166 398
rect 164 397 165 398
rect 137 397 138 398
rect 136 397 137 398
rect 135 397 136 398
rect 134 397 135 398
rect 133 397 134 398
rect 132 397 133 398
rect 131 397 132 398
rect 130 397 131 398
rect 129 397 130 398
rect 128 397 129 398
rect 127 397 128 398
rect 112 397 113 398
rect 111 397 112 398
rect 110 397 111 398
rect 109 397 110 398
rect 108 397 109 398
rect 107 397 108 398
rect 106 397 107 398
rect 105 397 106 398
rect 104 397 105 398
rect 103 397 104 398
rect 102 397 103 398
rect 85 397 86 398
rect 84 397 85 398
rect 83 397 84 398
rect 82 397 83 398
rect 81 397 82 398
rect 80 397 81 398
rect 79 397 80 398
rect 78 397 79 398
rect 77 397 78 398
rect 76 397 77 398
rect 75 397 76 398
rect 74 397 75 398
rect 63 397 64 398
rect 62 397 63 398
rect 61 397 62 398
rect 60 397 61 398
rect 59 397 60 398
rect 58 397 59 398
rect 57 397 58 398
rect 56 397 57 398
rect 55 397 56 398
rect 54 397 55 398
rect 53 397 54 398
rect 52 397 53 398
rect 196 398 197 399
rect 195 398 196 399
rect 194 398 195 399
rect 193 398 194 399
rect 192 398 193 399
rect 191 398 192 399
rect 183 398 184 399
rect 182 398 183 399
rect 181 398 182 399
rect 180 398 181 399
rect 171 398 172 399
rect 170 398 171 399
rect 169 398 170 399
rect 168 398 169 399
rect 167 398 168 399
rect 166 398 167 399
rect 165 398 166 399
rect 164 398 165 399
rect 138 398 139 399
rect 137 398 138 399
rect 136 398 137 399
rect 135 398 136 399
rect 134 398 135 399
rect 133 398 134 399
rect 132 398 133 399
rect 131 398 132 399
rect 130 398 131 399
rect 129 398 130 399
rect 128 398 129 399
rect 127 398 128 399
rect 112 398 113 399
rect 111 398 112 399
rect 110 398 111 399
rect 109 398 110 399
rect 108 398 109 399
rect 107 398 108 399
rect 106 398 107 399
rect 105 398 106 399
rect 104 398 105 399
rect 103 398 104 399
rect 102 398 103 399
rect 84 398 85 399
rect 83 398 84 399
rect 82 398 83 399
rect 81 398 82 399
rect 80 398 81 399
rect 79 398 80 399
rect 78 398 79 399
rect 77 398 78 399
rect 76 398 77 399
rect 75 398 76 399
rect 74 398 75 399
rect 73 398 74 399
rect 72 398 73 399
rect 71 398 72 399
rect 70 398 71 399
rect 69 398 70 399
rect 68 398 69 399
rect 67 398 68 399
rect 66 398 67 399
rect 65 398 66 399
rect 64 398 65 399
rect 63 398 64 399
rect 62 398 63 399
rect 61 398 62 399
rect 60 398 61 399
rect 59 398 60 399
rect 58 398 59 399
rect 57 398 58 399
rect 56 398 57 399
rect 55 398 56 399
rect 54 398 55 399
rect 53 398 54 399
rect 197 399 198 400
rect 196 399 197 400
rect 195 399 196 400
rect 194 399 195 400
rect 193 399 194 400
rect 192 399 193 400
rect 191 399 192 400
rect 183 399 184 400
rect 182 399 183 400
rect 181 399 182 400
rect 180 399 181 400
rect 171 399 172 400
rect 170 399 171 400
rect 169 399 170 400
rect 167 399 168 400
rect 166 399 167 400
rect 165 399 166 400
rect 164 399 165 400
rect 139 399 140 400
rect 138 399 139 400
rect 137 399 138 400
rect 136 399 137 400
rect 135 399 136 400
rect 134 399 135 400
rect 133 399 134 400
rect 132 399 133 400
rect 131 399 132 400
rect 130 399 131 400
rect 129 399 130 400
rect 128 399 129 400
rect 127 399 128 400
rect 112 399 113 400
rect 111 399 112 400
rect 110 399 111 400
rect 109 399 110 400
rect 108 399 109 400
rect 107 399 108 400
rect 106 399 107 400
rect 105 399 106 400
rect 104 399 105 400
rect 103 399 104 400
rect 102 399 103 400
rect 82 399 83 400
rect 81 399 82 400
rect 80 399 81 400
rect 79 399 80 400
rect 78 399 79 400
rect 77 399 78 400
rect 76 399 77 400
rect 75 399 76 400
rect 74 399 75 400
rect 73 399 74 400
rect 72 399 73 400
rect 71 399 72 400
rect 70 399 71 400
rect 69 399 70 400
rect 68 399 69 400
rect 67 399 68 400
rect 66 399 67 400
rect 65 399 66 400
rect 64 399 65 400
rect 63 399 64 400
rect 62 399 63 400
rect 61 399 62 400
rect 60 399 61 400
rect 59 399 60 400
rect 58 399 59 400
rect 57 399 58 400
rect 56 399 57 400
rect 55 399 56 400
rect 197 400 198 401
rect 196 400 197 401
rect 194 400 195 401
rect 192 400 193 401
rect 191 400 192 401
rect 183 400 184 401
rect 182 400 183 401
rect 181 400 182 401
rect 180 400 181 401
rect 171 400 172 401
rect 170 400 171 401
rect 169 400 170 401
rect 167 400 168 401
rect 166 400 167 401
rect 165 400 166 401
rect 164 400 165 401
rect 140 400 141 401
rect 139 400 140 401
rect 138 400 139 401
rect 137 400 138 401
rect 136 400 137 401
rect 135 400 136 401
rect 134 400 135 401
rect 133 400 134 401
rect 132 400 133 401
rect 131 400 132 401
rect 130 400 131 401
rect 129 400 130 401
rect 128 400 129 401
rect 127 400 128 401
rect 112 400 113 401
rect 111 400 112 401
rect 110 400 111 401
rect 109 400 110 401
rect 108 400 109 401
rect 107 400 108 401
rect 106 400 107 401
rect 105 400 106 401
rect 104 400 105 401
rect 103 400 104 401
rect 102 400 103 401
rect 80 400 81 401
rect 79 400 80 401
rect 78 400 79 401
rect 77 400 78 401
rect 76 400 77 401
rect 75 400 76 401
rect 74 400 75 401
rect 73 400 74 401
rect 72 400 73 401
rect 71 400 72 401
rect 70 400 71 401
rect 69 400 70 401
rect 68 400 69 401
rect 67 400 68 401
rect 66 400 67 401
rect 65 400 66 401
rect 64 400 65 401
rect 63 400 64 401
rect 62 400 63 401
rect 61 400 62 401
rect 60 400 61 401
rect 59 400 60 401
rect 58 400 59 401
rect 57 400 58 401
rect 197 401 198 402
rect 196 401 197 402
rect 194 401 195 402
rect 193 401 194 402
rect 192 401 193 402
rect 191 401 192 402
rect 183 401 184 402
rect 182 401 183 402
rect 181 401 182 402
rect 180 401 181 402
rect 171 401 172 402
rect 170 401 171 402
rect 169 401 170 402
rect 167 401 168 402
rect 166 401 167 402
rect 165 401 166 402
rect 164 401 165 402
rect 140 401 141 402
rect 139 401 140 402
rect 138 401 139 402
rect 137 401 138 402
rect 136 401 137 402
rect 135 401 136 402
rect 134 401 135 402
rect 133 401 134 402
rect 132 401 133 402
rect 131 401 132 402
rect 130 401 131 402
rect 129 401 130 402
rect 128 401 129 402
rect 127 401 128 402
rect 112 401 113 402
rect 111 401 112 402
rect 110 401 111 402
rect 109 401 110 402
rect 108 401 109 402
rect 107 401 108 402
rect 106 401 107 402
rect 105 401 106 402
rect 104 401 105 402
rect 103 401 104 402
rect 102 401 103 402
rect 78 401 79 402
rect 77 401 78 402
rect 76 401 77 402
rect 75 401 76 402
rect 74 401 75 402
rect 73 401 74 402
rect 72 401 73 402
rect 71 401 72 402
rect 70 401 71 402
rect 69 401 70 402
rect 68 401 69 402
rect 67 401 68 402
rect 66 401 67 402
rect 65 401 66 402
rect 64 401 65 402
rect 63 401 64 402
rect 62 401 63 402
rect 61 401 62 402
rect 60 401 61 402
rect 59 401 60 402
rect 196 402 197 403
rect 194 402 195 403
rect 193 402 194 403
rect 192 402 193 403
rect 191 402 192 403
rect 183 402 184 403
rect 182 402 183 403
rect 181 402 182 403
rect 180 402 181 403
rect 177 402 178 403
rect 176 402 177 403
rect 175 402 176 403
rect 174 402 175 403
rect 173 402 174 403
rect 172 402 173 403
rect 171 402 172 403
rect 170 402 171 403
rect 169 402 170 403
rect 168 402 169 403
rect 167 402 168 403
rect 166 402 167 403
rect 165 402 166 403
rect 164 402 165 403
rect 163 402 164 403
rect 162 402 163 403
rect 141 402 142 403
rect 140 402 141 403
rect 139 402 140 403
rect 138 402 139 403
rect 137 402 138 403
rect 136 402 137 403
rect 135 402 136 403
rect 134 402 135 403
rect 133 402 134 403
rect 132 402 133 403
rect 131 402 132 403
rect 130 402 131 403
rect 129 402 130 403
rect 128 402 129 403
rect 127 402 128 403
rect 112 402 113 403
rect 111 402 112 403
rect 110 402 111 403
rect 109 402 110 403
rect 108 402 109 403
rect 107 402 108 403
rect 106 402 107 403
rect 105 402 106 403
rect 104 402 105 403
rect 103 402 104 403
rect 102 402 103 403
rect 74 402 75 403
rect 73 402 74 403
rect 72 402 73 403
rect 71 402 72 403
rect 70 402 71 403
rect 69 402 70 403
rect 68 402 69 403
rect 67 402 68 403
rect 66 402 67 403
rect 65 402 66 403
rect 64 402 65 403
rect 63 402 64 403
rect 62 402 63 403
rect 194 403 195 404
rect 193 403 194 404
rect 183 403 184 404
rect 182 403 183 404
rect 181 403 182 404
rect 180 403 181 404
rect 177 403 178 404
rect 176 403 177 404
rect 175 403 176 404
rect 174 403 175 404
rect 173 403 174 404
rect 172 403 173 404
rect 171 403 172 404
rect 170 403 171 404
rect 169 403 170 404
rect 168 403 169 404
rect 167 403 168 404
rect 166 403 167 404
rect 165 403 166 404
rect 164 403 165 404
rect 163 403 164 404
rect 162 403 163 404
rect 142 403 143 404
rect 141 403 142 404
rect 140 403 141 404
rect 139 403 140 404
rect 138 403 139 404
rect 137 403 138 404
rect 136 403 137 404
rect 135 403 136 404
rect 134 403 135 404
rect 133 403 134 404
rect 132 403 133 404
rect 131 403 132 404
rect 130 403 131 404
rect 129 403 130 404
rect 128 403 129 404
rect 127 403 128 404
rect 112 403 113 404
rect 111 403 112 404
rect 110 403 111 404
rect 109 403 110 404
rect 108 403 109 404
rect 107 403 108 404
rect 106 403 107 404
rect 105 403 106 404
rect 104 403 105 404
rect 103 403 104 404
rect 102 403 103 404
rect 196 404 197 405
rect 195 404 196 405
rect 194 404 195 405
rect 183 404 184 405
rect 182 404 183 405
rect 181 404 182 405
rect 180 404 181 405
rect 177 404 178 405
rect 176 404 177 405
rect 175 404 176 405
rect 174 404 175 405
rect 173 404 174 405
rect 172 404 173 405
rect 171 404 172 405
rect 170 404 171 405
rect 169 404 170 405
rect 168 404 169 405
rect 167 404 168 405
rect 166 404 167 405
rect 165 404 166 405
rect 164 404 165 405
rect 163 404 164 405
rect 162 404 163 405
rect 143 404 144 405
rect 142 404 143 405
rect 141 404 142 405
rect 140 404 141 405
rect 139 404 140 405
rect 138 404 139 405
rect 137 404 138 405
rect 136 404 137 405
rect 135 404 136 405
rect 134 404 135 405
rect 133 404 134 405
rect 132 404 133 405
rect 131 404 132 405
rect 130 404 131 405
rect 129 404 130 405
rect 128 404 129 405
rect 127 404 128 405
rect 112 404 113 405
rect 111 404 112 405
rect 110 404 111 405
rect 109 404 110 405
rect 108 404 109 405
rect 107 404 108 405
rect 106 404 107 405
rect 105 404 106 405
rect 104 404 105 405
rect 103 404 104 405
rect 102 404 103 405
rect 197 405 198 406
rect 196 405 197 406
rect 195 405 196 406
rect 194 405 195 406
rect 192 405 193 406
rect 191 405 192 406
rect 183 405 184 406
rect 182 405 183 406
rect 181 405 182 406
rect 180 405 181 406
rect 177 405 178 406
rect 176 405 177 406
rect 175 405 176 406
rect 174 405 175 406
rect 173 405 174 406
rect 172 405 173 406
rect 171 405 172 406
rect 170 405 171 406
rect 169 405 170 406
rect 168 405 169 406
rect 167 405 168 406
rect 166 405 167 406
rect 165 405 166 406
rect 164 405 165 406
rect 163 405 164 406
rect 162 405 163 406
rect 144 405 145 406
rect 143 405 144 406
rect 142 405 143 406
rect 141 405 142 406
rect 140 405 141 406
rect 139 405 140 406
rect 138 405 139 406
rect 137 405 138 406
rect 136 405 137 406
rect 135 405 136 406
rect 134 405 135 406
rect 133 405 134 406
rect 132 405 133 406
rect 131 405 132 406
rect 130 405 131 406
rect 129 405 130 406
rect 128 405 129 406
rect 127 405 128 406
rect 112 405 113 406
rect 111 405 112 406
rect 110 405 111 406
rect 109 405 110 406
rect 108 405 109 406
rect 107 405 108 406
rect 106 405 107 406
rect 105 405 106 406
rect 104 405 105 406
rect 103 405 104 406
rect 102 405 103 406
rect 197 406 198 407
rect 196 406 197 407
rect 194 406 195 407
rect 193 406 194 407
rect 192 406 193 407
rect 191 406 192 407
rect 182 406 183 407
rect 181 406 182 407
rect 180 406 181 407
rect 176 406 177 407
rect 175 406 176 407
rect 174 406 175 407
rect 173 406 174 407
rect 172 406 173 407
rect 171 406 172 407
rect 170 406 171 407
rect 169 406 170 407
rect 168 406 169 407
rect 167 406 168 407
rect 166 406 167 407
rect 165 406 166 407
rect 164 406 165 407
rect 163 406 164 407
rect 144 406 145 407
rect 143 406 144 407
rect 142 406 143 407
rect 141 406 142 407
rect 140 406 141 407
rect 139 406 140 407
rect 138 406 139 407
rect 137 406 138 407
rect 136 406 137 407
rect 135 406 136 407
rect 134 406 135 407
rect 133 406 134 407
rect 132 406 133 407
rect 131 406 132 407
rect 130 406 131 407
rect 129 406 130 407
rect 128 406 129 407
rect 127 406 128 407
rect 112 406 113 407
rect 111 406 112 407
rect 110 406 111 407
rect 109 406 110 407
rect 108 406 109 407
rect 107 406 108 407
rect 106 406 107 407
rect 105 406 106 407
rect 104 406 105 407
rect 103 406 104 407
rect 102 406 103 407
rect 196 407 197 408
rect 194 407 195 408
rect 193 407 194 408
rect 192 407 193 408
rect 191 407 192 408
rect 145 407 146 408
rect 144 407 145 408
rect 143 407 144 408
rect 142 407 143 408
rect 141 407 142 408
rect 140 407 141 408
rect 139 407 140 408
rect 138 407 139 408
rect 137 407 138 408
rect 136 407 137 408
rect 135 407 136 408
rect 134 407 135 408
rect 133 407 134 408
rect 132 407 133 408
rect 131 407 132 408
rect 130 407 131 408
rect 129 407 130 408
rect 128 407 129 408
rect 127 407 128 408
rect 112 407 113 408
rect 111 407 112 408
rect 110 407 111 408
rect 109 407 110 408
rect 108 407 109 408
rect 107 407 108 408
rect 106 407 107 408
rect 105 407 106 408
rect 104 407 105 408
rect 103 407 104 408
rect 102 407 103 408
rect 197 408 198 409
rect 196 408 197 409
rect 195 408 196 409
rect 194 408 195 409
rect 193 408 194 409
rect 192 408 193 409
rect 191 408 192 409
rect 146 408 147 409
rect 145 408 146 409
rect 144 408 145 409
rect 143 408 144 409
rect 142 408 143 409
rect 141 408 142 409
rect 140 408 141 409
rect 139 408 140 409
rect 138 408 139 409
rect 137 408 138 409
rect 136 408 137 409
rect 135 408 136 409
rect 134 408 135 409
rect 133 408 134 409
rect 132 408 133 409
rect 131 408 132 409
rect 130 408 131 409
rect 129 408 130 409
rect 128 408 129 409
rect 127 408 128 409
rect 112 408 113 409
rect 111 408 112 409
rect 110 408 111 409
rect 109 408 110 409
rect 108 408 109 409
rect 107 408 108 409
rect 106 408 107 409
rect 105 408 106 409
rect 104 408 105 409
rect 103 408 104 409
rect 102 408 103 409
rect 196 409 197 410
rect 195 409 196 410
rect 194 409 195 410
rect 193 409 194 410
rect 192 409 193 410
rect 191 409 192 410
rect 147 409 148 410
rect 146 409 147 410
rect 145 409 146 410
rect 144 409 145 410
rect 143 409 144 410
rect 142 409 143 410
rect 141 409 142 410
rect 140 409 141 410
rect 139 409 140 410
rect 138 409 139 410
rect 137 409 138 410
rect 136 409 137 410
rect 135 409 136 410
rect 134 409 135 410
rect 133 409 134 410
rect 132 409 133 410
rect 131 409 132 410
rect 130 409 131 410
rect 129 409 130 410
rect 128 409 129 410
rect 127 409 128 410
rect 112 409 113 410
rect 111 409 112 410
rect 110 409 111 410
rect 109 409 110 410
rect 108 409 109 410
rect 107 409 108 410
rect 106 409 107 410
rect 105 409 106 410
rect 104 409 105 410
rect 103 409 104 410
rect 102 409 103 410
rect 148 410 149 411
rect 147 410 148 411
rect 146 410 147 411
rect 145 410 146 411
rect 144 410 145 411
rect 143 410 144 411
rect 142 410 143 411
rect 141 410 142 411
rect 140 410 141 411
rect 139 410 140 411
rect 138 410 139 411
rect 137 410 138 411
rect 136 410 137 411
rect 135 410 136 411
rect 134 410 135 411
rect 133 410 134 411
rect 132 410 133 411
rect 131 410 132 411
rect 130 410 131 411
rect 129 410 130 411
rect 128 410 129 411
rect 127 410 128 411
rect 112 410 113 411
rect 111 410 112 411
rect 110 410 111 411
rect 109 410 110 411
rect 108 410 109 411
rect 107 410 108 411
rect 106 410 107 411
rect 105 410 106 411
rect 104 410 105 411
rect 103 410 104 411
rect 102 410 103 411
rect 196 411 197 412
rect 195 411 196 412
rect 194 411 195 412
rect 193 411 194 412
rect 192 411 193 412
rect 191 411 192 412
rect 149 411 150 412
rect 148 411 149 412
rect 147 411 148 412
rect 146 411 147 412
rect 145 411 146 412
rect 144 411 145 412
rect 143 411 144 412
rect 142 411 143 412
rect 141 411 142 412
rect 140 411 141 412
rect 139 411 140 412
rect 138 411 139 412
rect 137 411 138 412
rect 136 411 137 412
rect 135 411 136 412
rect 134 411 135 412
rect 133 411 134 412
rect 132 411 133 412
rect 131 411 132 412
rect 130 411 131 412
rect 129 411 130 412
rect 128 411 129 412
rect 127 411 128 412
rect 112 411 113 412
rect 111 411 112 412
rect 110 411 111 412
rect 109 411 110 412
rect 108 411 109 412
rect 107 411 108 412
rect 106 411 107 412
rect 105 411 106 412
rect 104 411 105 412
rect 103 411 104 412
rect 102 411 103 412
rect 197 412 198 413
rect 196 412 197 413
rect 195 412 196 413
rect 194 412 195 413
rect 193 412 194 413
rect 192 412 193 413
rect 191 412 192 413
rect 149 412 150 413
rect 148 412 149 413
rect 147 412 148 413
rect 146 412 147 413
rect 145 412 146 413
rect 144 412 145 413
rect 143 412 144 413
rect 142 412 143 413
rect 141 412 142 413
rect 140 412 141 413
rect 139 412 140 413
rect 138 412 139 413
rect 137 412 138 413
rect 136 412 137 413
rect 135 412 136 413
rect 134 412 135 413
rect 133 412 134 413
rect 132 412 133 413
rect 131 412 132 413
rect 130 412 131 413
rect 129 412 130 413
rect 128 412 129 413
rect 127 412 128 413
rect 126 412 127 413
rect 125 412 126 413
rect 124 412 125 413
rect 123 412 124 413
rect 122 412 123 413
rect 121 412 122 413
rect 120 412 121 413
rect 119 412 120 413
rect 118 412 119 413
rect 117 412 118 413
rect 116 412 117 413
rect 115 412 116 413
rect 114 412 115 413
rect 113 412 114 413
rect 112 412 113 413
rect 111 412 112 413
rect 110 412 111 413
rect 109 412 110 413
rect 108 412 109 413
rect 107 412 108 413
rect 106 412 107 413
rect 105 412 106 413
rect 104 412 105 413
rect 103 412 104 413
rect 102 412 103 413
rect 192 413 193 414
rect 191 413 192 414
rect 150 413 151 414
rect 149 413 150 414
rect 148 413 149 414
rect 147 413 148 414
rect 146 413 147 414
rect 145 413 146 414
rect 144 413 145 414
rect 143 413 144 414
rect 142 413 143 414
rect 141 413 142 414
rect 140 413 141 414
rect 139 413 140 414
rect 138 413 139 414
rect 137 413 138 414
rect 136 413 137 414
rect 135 413 136 414
rect 134 413 135 414
rect 133 413 134 414
rect 132 413 133 414
rect 131 413 132 414
rect 130 413 131 414
rect 129 413 130 414
rect 128 413 129 414
rect 127 413 128 414
rect 126 413 127 414
rect 125 413 126 414
rect 124 413 125 414
rect 123 413 124 414
rect 122 413 123 414
rect 121 413 122 414
rect 120 413 121 414
rect 119 413 120 414
rect 118 413 119 414
rect 117 413 118 414
rect 116 413 117 414
rect 115 413 116 414
rect 114 413 115 414
rect 113 413 114 414
rect 112 413 113 414
rect 111 413 112 414
rect 110 413 111 414
rect 109 413 110 414
rect 108 413 109 414
rect 107 413 108 414
rect 106 413 107 414
rect 105 413 106 414
rect 104 413 105 414
rect 103 413 104 414
rect 102 413 103 414
rect 192 414 193 415
rect 191 414 192 415
rect 151 414 152 415
rect 150 414 151 415
rect 149 414 150 415
rect 148 414 149 415
rect 147 414 148 415
rect 146 414 147 415
rect 145 414 146 415
rect 144 414 145 415
rect 143 414 144 415
rect 142 414 143 415
rect 141 414 142 415
rect 140 414 141 415
rect 139 414 140 415
rect 138 414 139 415
rect 137 414 138 415
rect 136 414 137 415
rect 135 414 136 415
rect 134 414 135 415
rect 133 414 134 415
rect 132 414 133 415
rect 131 414 132 415
rect 130 414 131 415
rect 129 414 130 415
rect 127 414 128 415
rect 126 414 127 415
rect 125 414 126 415
rect 124 414 125 415
rect 123 414 124 415
rect 122 414 123 415
rect 121 414 122 415
rect 120 414 121 415
rect 119 414 120 415
rect 118 414 119 415
rect 117 414 118 415
rect 116 414 117 415
rect 115 414 116 415
rect 114 414 115 415
rect 113 414 114 415
rect 112 414 113 415
rect 111 414 112 415
rect 110 414 111 415
rect 109 414 110 415
rect 108 414 109 415
rect 107 414 108 415
rect 106 414 107 415
rect 105 414 106 415
rect 104 414 105 415
rect 103 414 104 415
rect 102 414 103 415
rect 196 415 197 416
rect 195 415 196 416
rect 194 415 195 416
rect 193 415 194 416
rect 192 415 193 416
rect 152 415 153 416
rect 151 415 152 416
rect 150 415 151 416
rect 149 415 150 416
rect 148 415 149 416
rect 147 415 148 416
rect 146 415 147 416
rect 145 415 146 416
rect 144 415 145 416
rect 143 415 144 416
rect 142 415 143 416
rect 141 415 142 416
rect 140 415 141 416
rect 139 415 140 416
rect 138 415 139 416
rect 137 415 138 416
rect 136 415 137 416
rect 135 415 136 416
rect 134 415 135 416
rect 133 415 134 416
rect 132 415 133 416
rect 131 415 132 416
rect 130 415 131 416
rect 127 415 128 416
rect 126 415 127 416
rect 125 415 126 416
rect 124 415 125 416
rect 123 415 124 416
rect 122 415 123 416
rect 121 415 122 416
rect 120 415 121 416
rect 119 415 120 416
rect 118 415 119 416
rect 117 415 118 416
rect 116 415 117 416
rect 115 415 116 416
rect 114 415 115 416
rect 113 415 114 416
rect 112 415 113 416
rect 111 415 112 416
rect 110 415 111 416
rect 109 415 110 416
rect 108 415 109 416
rect 107 415 108 416
rect 106 415 107 416
rect 105 415 106 416
rect 104 415 105 416
rect 103 415 104 416
rect 102 415 103 416
rect 196 416 197 417
rect 195 416 196 417
rect 194 416 195 417
rect 193 416 194 417
rect 192 416 193 417
rect 191 416 192 417
rect 153 416 154 417
rect 152 416 153 417
rect 151 416 152 417
rect 150 416 151 417
rect 149 416 150 417
rect 148 416 149 417
rect 147 416 148 417
rect 146 416 147 417
rect 145 416 146 417
rect 144 416 145 417
rect 143 416 144 417
rect 142 416 143 417
rect 141 416 142 417
rect 140 416 141 417
rect 139 416 140 417
rect 138 416 139 417
rect 137 416 138 417
rect 136 416 137 417
rect 135 416 136 417
rect 134 416 135 417
rect 133 416 134 417
rect 132 416 133 417
rect 131 416 132 417
rect 127 416 128 417
rect 126 416 127 417
rect 125 416 126 417
rect 124 416 125 417
rect 123 416 124 417
rect 122 416 123 417
rect 121 416 122 417
rect 120 416 121 417
rect 119 416 120 417
rect 118 416 119 417
rect 117 416 118 417
rect 116 416 117 417
rect 115 416 116 417
rect 114 416 115 417
rect 113 416 114 417
rect 112 416 113 417
rect 111 416 112 417
rect 110 416 111 417
rect 109 416 110 417
rect 108 416 109 417
rect 107 416 108 417
rect 106 416 107 417
rect 105 416 106 417
rect 104 416 105 417
rect 103 416 104 417
rect 102 416 103 417
rect 196 417 197 418
rect 195 417 196 418
rect 192 417 193 418
rect 191 417 192 418
rect 153 417 154 418
rect 152 417 153 418
rect 151 417 152 418
rect 150 417 151 418
rect 149 417 150 418
rect 148 417 149 418
rect 147 417 148 418
rect 146 417 147 418
rect 145 417 146 418
rect 144 417 145 418
rect 143 417 144 418
rect 142 417 143 418
rect 141 417 142 418
rect 140 417 141 418
rect 139 417 140 418
rect 138 417 139 418
rect 137 417 138 418
rect 136 417 137 418
rect 135 417 136 418
rect 134 417 135 418
rect 133 417 134 418
rect 132 417 133 418
rect 131 417 132 418
rect 127 417 128 418
rect 126 417 127 418
rect 125 417 126 418
rect 124 417 125 418
rect 123 417 124 418
rect 122 417 123 418
rect 121 417 122 418
rect 120 417 121 418
rect 119 417 120 418
rect 118 417 119 418
rect 117 417 118 418
rect 116 417 117 418
rect 115 417 116 418
rect 114 417 115 418
rect 113 417 114 418
rect 112 417 113 418
rect 111 417 112 418
rect 110 417 111 418
rect 109 417 110 418
rect 108 417 109 418
rect 107 417 108 418
rect 106 417 107 418
rect 105 417 106 418
rect 104 417 105 418
rect 103 417 104 418
rect 102 417 103 418
rect 197 418 198 419
rect 196 418 197 419
rect 192 418 193 419
rect 191 418 192 419
rect 174 418 175 419
rect 173 418 174 419
rect 172 418 173 419
rect 153 418 154 419
rect 152 418 153 419
rect 151 418 152 419
rect 150 418 151 419
rect 149 418 150 419
rect 148 418 149 419
rect 147 418 148 419
rect 146 418 147 419
rect 145 418 146 419
rect 144 418 145 419
rect 143 418 144 419
rect 142 418 143 419
rect 141 418 142 419
rect 140 418 141 419
rect 139 418 140 419
rect 138 418 139 419
rect 137 418 138 419
rect 136 418 137 419
rect 135 418 136 419
rect 134 418 135 419
rect 133 418 134 419
rect 132 418 133 419
rect 127 418 128 419
rect 126 418 127 419
rect 125 418 126 419
rect 124 418 125 419
rect 123 418 124 419
rect 122 418 123 419
rect 121 418 122 419
rect 120 418 121 419
rect 119 418 120 419
rect 118 418 119 419
rect 117 418 118 419
rect 116 418 117 419
rect 115 418 116 419
rect 114 418 115 419
rect 113 418 114 419
rect 112 418 113 419
rect 111 418 112 419
rect 110 418 111 419
rect 109 418 110 419
rect 108 418 109 419
rect 107 418 108 419
rect 106 418 107 419
rect 105 418 106 419
rect 104 418 105 419
rect 103 418 104 419
rect 102 418 103 419
rect 196 419 197 420
rect 191 419 192 420
rect 174 419 175 420
rect 173 419 174 420
rect 172 419 173 420
rect 153 419 154 420
rect 152 419 153 420
rect 151 419 152 420
rect 150 419 151 420
rect 149 419 150 420
rect 148 419 149 420
rect 147 419 148 420
rect 146 419 147 420
rect 145 419 146 420
rect 144 419 145 420
rect 143 419 144 420
rect 142 419 143 420
rect 141 419 142 420
rect 140 419 141 420
rect 139 419 140 420
rect 138 419 139 420
rect 137 419 138 420
rect 136 419 137 420
rect 135 419 136 420
rect 134 419 135 420
rect 133 419 134 420
rect 127 419 128 420
rect 126 419 127 420
rect 125 419 126 420
rect 124 419 125 420
rect 123 419 124 420
rect 122 419 123 420
rect 121 419 122 420
rect 120 419 121 420
rect 119 419 120 420
rect 118 419 119 420
rect 117 419 118 420
rect 116 419 117 420
rect 115 419 116 420
rect 114 419 115 420
rect 113 419 114 420
rect 112 419 113 420
rect 111 419 112 420
rect 110 419 111 420
rect 109 419 110 420
rect 108 419 109 420
rect 107 419 108 420
rect 106 419 107 420
rect 105 419 106 420
rect 104 419 105 420
rect 103 419 104 420
rect 102 419 103 420
rect 174 420 175 421
rect 173 420 174 421
rect 172 420 173 421
rect 164 420 165 421
rect 153 420 154 421
rect 152 420 153 421
rect 151 420 152 421
rect 150 420 151 421
rect 149 420 150 421
rect 148 420 149 421
rect 147 420 148 421
rect 146 420 147 421
rect 145 420 146 421
rect 144 420 145 421
rect 143 420 144 421
rect 142 420 143 421
rect 141 420 142 421
rect 140 420 141 421
rect 139 420 140 421
rect 138 420 139 421
rect 137 420 138 421
rect 136 420 137 421
rect 135 420 136 421
rect 134 420 135 421
rect 127 420 128 421
rect 126 420 127 421
rect 125 420 126 421
rect 124 420 125 421
rect 123 420 124 421
rect 122 420 123 421
rect 121 420 122 421
rect 120 420 121 421
rect 119 420 120 421
rect 118 420 119 421
rect 117 420 118 421
rect 116 420 117 421
rect 115 420 116 421
rect 114 420 115 421
rect 113 420 114 421
rect 112 420 113 421
rect 111 420 112 421
rect 110 420 111 421
rect 109 420 110 421
rect 108 420 109 421
rect 107 420 108 421
rect 106 420 107 421
rect 105 420 106 421
rect 104 420 105 421
rect 103 420 104 421
rect 102 420 103 421
rect 197 421 198 422
rect 196 421 197 422
rect 195 421 196 422
rect 194 421 195 422
rect 193 421 194 422
rect 192 421 193 422
rect 191 421 192 422
rect 190 421 191 422
rect 189 421 190 422
rect 188 421 189 422
rect 174 421 175 422
rect 173 421 174 422
rect 172 421 173 422
rect 165 421 166 422
rect 164 421 165 422
rect 163 421 164 422
rect 153 421 154 422
rect 152 421 153 422
rect 151 421 152 422
rect 150 421 151 422
rect 149 421 150 422
rect 148 421 149 422
rect 147 421 148 422
rect 146 421 147 422
rect 145 421 146 422
rect 144 421 145 422
rect 143 421 144 422
rect 142 421 143 422
rect 141 421 142 422
rect 140 421 141 422
rect 139 421 140 422
rect 138 421 139 422
rect 137 421 138 422
rect 136 421 137 422
rect 135 421 136 422
rect 127 421 128 422
rect 126 421 127 422
rect 125 421 126 422
rect 124 421 125 422
rect 123 421 124 422
rect 122 421 123 422
rect 121 421 122 422
rect 120 421 121 422
rect 119 421 120 422
rect 118 421 119 422
rect 117 421 118 422
rect 116 421 117 422
rect 115 421 116 422
rect 114 421 115 422
rect 113 421 114 422
rect 112 421 113 422
rect 111 421 112 422
rect 110 421 111 422
rect 109 421 110 422
rect 108 421 109 422
rect 107 421 108 422
rect 106 421 107 422
rect 105 421 106 422
rect 104 421 105 422
rect 103 421 104 422
rect 102 421 103 422
rect 196 422 197 423
rect 195 422 196 423
rect 194 422 195 423
rect 193 422 194 423
rect 192 422 193 423
rect 191 422 192 423
rect 190 422 191 423
rect 189 422 190 423
rect 188 422 189 423
rect 174 422 175 423
rect 173 422 174 423
rect 172 422 173 423
rect 165 422 166 423
rect 164 422 165 423
rect 163 422 164 423
rect 153 422 154 423
rect 152 422 153 423
rect 151 422 152 423
rect 150 422 151 423
rect 149 422 150 423
rect 148 422 149 423
rect 147 422 148 423
rect 146 422 147 423
rect 145 422 146 423
rect 144 422 145 423
rect 143 422 144 423
rect 142 422 143 423
rect 141 422 142 423
rect 140 422 141 423
rect 139 422 140 423
rect 138 422 139 423
rect 137 422 138 423
rect 136 422 137 423
rect 127 422 128 423
rect 126 422 127 423
rect 125 422 126 423
rect 124 422 125 423
rect 123 422 124 423
rect 122 422 123 423
rect 121 422 122 423
rect 120 422 121 423
rect 119 422 120 423
rect 118 422 119 423
rect 117 422 118 423
rect 116 422 117 423
rect 115 422 116 423
rect 114 422 115 423
rect 113 422 114 423
rect 112 422 113 423
rect 111 422 112 423
rect 110 422 111 423
rect 109 422 110 423
rect 108 422 109 423
rect 107 422 108 423
rect 106 422 107 423
rect 105 422 106 423
rect 104 422 105 423
rect 103 422 104 423
rect 102 422 103 423
rect 192 423 193 424
rect 191 423 192 424
rect 174 423 175 424
rect 173 423 174 424
rect 172 423 173 424
rect 165 423 166 424
rect 164 423 165 424
rect 163 423 164 424
rect 153 423 154 424
rect 152 423 153 424
rect 151 423 152 424
rect 150 423 151 424
rect 149 423 150 424
rect 148 423 149 424
rect 147 423 148 424
rect 146 423 147 424
rect 145 423 146 424
rect 144 423 145 424
rect 143 423 144 424
rect 142 423 143 424
rect 141 423 142 424
rect 140 423 141 424
rect 139 423 140 424
rect 138 423 139 424
rect 137 423 138 424
rect 136 423 137 424
rect 127 423 128 424
rect 126 423 127 424
rect 125 423 126 424
rect 124 423 125 424
rect 123 423 124 424
rect 122 423 123 424
rect 121 423 122 424
rect 120 423 121 424
rect 119 423 120 424
rect 118 423 119 424
rect 117 423 118 424
rect 116 423 117 424
rect 115 423 116 424
rect 114 423 115 424
rect 113 423 114 424
rect 112 423 113 424
rect 111 423 112 424
rect 110 423 111 424
rect 109 423 110 424
rect 108 423 109 424
rect 107 423 108 424
rect 106 423 107 424
rect 105 423 106 424
rect 104 423 105 424
rect 103 423 104 424
rect 102 423 103 424
rect 196 424 197 425
rect 195 424 196 425
rect 194 424 195 425
rect 192 424 193 425
rect 191 424 192 425
rect 174 424 175 425
rect 173 424 174 425
rect 172 424 173 425
rect 165 424 166 425
rect 164 424 165 425
rect 163 424 164 425
rect 153 424 154 425
rect 152 424 153 425
rect 151 424 152 425
rect 150 424 151 425
rect 149 424 150 425
rect 148 424 149 425
rect 147 424 148 425
rect 146 424 147 425
rect 145 424 146 425
rect 144 424 145 425
rect 143 424 144 425
rect 142 424 143 425
rect 141 424 142 425
rect 140 424 141 425
rect 139 424 140 425
rect 138 424 139 425
rect 137 424 138 425
rect 127 424 128 425
rect 126 424 127 425
rect 125 424 126 425
rect 124 424 125 425
rect 123 424 124 425
rect 122 424 123 425
rect 121 424 122 425
rect 120 424 121 425
rect 119 424 120 425
rect 118 424 119 425
rect 117 424 118 425
rect 116 424 117 425
rect 115 424 116 425
rect 114 424 115 425
rect 113 424 114 425
rect 112 424 113 425
rect 111 424 112 425
rect 110 424 111 425
rect 109 424 110 425
rect 108 424 109 425
rect 107 424 108 425
rect 106 424 107 425
rect 105 424 106 425
rect 104 424 105 425
rect 103 424 104 425
rect 102 424 103 425
rect 197 425 198 426
rect 196 425 197 426
rect 195 425 196 426
rect 194 425 195 426
rect 193 425 194 426
rect 192 425 193 426
rect 191 425 192 426
rect 174 425 175 426
rect 173 425 174 426
rect 172 425 173 426
rect 165 425 166 426
rect 164 425 165 426
rect 163 425 164 426
rect 153 425 154 426
rect 152 425 153 426
rect 151 425 152 426
rect 150 425 151 426
rect 149 425 150 426
rect 148 425 149 426
rect 147 425 148 426
rect 146 425 147 426
rect 145 425 146 426
rect 144 425 145 426
rect 143 425 144 426
rect 142 425 143 426
rect 141 425 142 426
rect 140 425 141 426
rect 139 425 140 426
rect 138 425 139 426
rect 127 425 128 426
rect 126 425 127 426
rect 125 425 126 426
rect 124 425 125 426
rect 123 425 124 426
rect 122 425 123 426
rect 121 425 122 426
rect 120 425 121 426
rect 119 425 120 426
rect 118 425 119 426
rect 117 425 118 426
rect 116 425 117 426
rect 115 425 116 426
rect 114 425 115 426
rect 113 425 114 426
rect 112 425 113 426
rect 111 425 112 426
rect 110 425 111 426
rect 109 425 110 426
rect 108 425 109 426
rect 107 425 108 426
rect 106 425 107 426
rect 105 425 106 426
rect 104 425 105 426
rect 103 425 104 426
rect 102 425 103 426
rect 174 426 175 427
rect 173 426 174 427
rect 172 426 173 427
rect 165 426 166 427
rect 164 426 165 427
rect 163 426 164 427
rect 153 426 154 427
rect 152 426 153 427
rect 151 426 152 427
rect 150 426 151 427
rect 149 426 150 427
rect 148 426 149 427
rect 147 426 148 427
rect 146 426 147 427
rect 145 426 146 427
rect 144 426 145 427
rect 143 426 144 427
rect 142 426 143 427
rect 141 426 142 427
rect 140 426 141 427
rect 139 426 140 427
rect 127 426 128 427
rect 126 426 127 427
rect 125 426 126 427
rect 124 426 125 427
rect 123 426 124 427
rect 122 426 123 427
rect 121 426 122 427
rect 120 426 121 427
rect 119 426 120 427
rect 118 426 119 427
rect 117 426 118 427
rect 116 426 117 427
rect 115 426 116 427
rect 114 426 115 427
rect 113 426 114 427
rect 112 426 113 427
rect 111 426 112 427
rect 110 426 111 427
rect 109 426 110 427
rect 108 426 109 427
rect 107 426 108 427
rect 106 426 107 427
rect 105 426 106 427
rect 104 426 105 427
rect 103 426 104 427
rect 102 426 103 427
rect 174 427 175 428
rect 173 427 174 428
rect 172 427 173 428
rect 165 427 166 428
rect 164 427 165 428
rect 163 427 164 428
rect 153 427 154 428
rect 152 427 153 428
rect 151 427 152 428
rect 150 427 151 428
rect 149 427 150 428
rect 148 427 149 428
rect 147 427 148 428
rect 146 427 147 428
rect 145 427 146 428
rect 144 427 145 428
rect 143 427 144 428
rect 142 427 143 428
rect 141 427 142 428
rect 140 427 141 428
rect 127 427 128 428
rect 126 427 127 428
rect 125 427 126 428
rect 124 427 125 428
rect 123 427 124 428
rect 122 427 123 428
rect 121 427 122 428
rect 120 427 121 428
rect 119 427 120 428
rect 118 427 119 428
rect 117 427 118 428
rect 116 427 117 428
rect 115 427 116 428
rect 114 427 115 428
rect 113 427 114 428
rect 112 427 113 428
rect 111 427 112 428
rect 110 427 111 428
rect 109 427 110 428
rect 108 427 109 428
rect 107 427 108 428
rect 106 427 107 428
rect 105 427 106 428
rect 104 427 105 428
rect 103 427 104 428
rect 102 427 103 428
rect 183 428 184 429
rect 182 428 183 429
rect 181 428 182 429
rect 180 428 181 429
rect 179 428 180 429
rect 178 428 179 429
rect 177 428 178 429
rect 176 428 177 429
rect 175 428 176 429
rect 174 428 175 429
rect 173 428 174 429
rect 172 428 173 429
rect 165 428 166 429
rect 164 428 165 429
rect 163 428 164 429
rect 153 428 154 429
rect 152 428 153 429
rect 151 428 152 429
rect 150 428 151 429
rect 149 428 150 429
rect 148 428 149 429
rect 147 428 148 429
rect 146 428 147 429
rect 145 428 146 429
rect 144 428 145 429
rect 143 428 144 429
rect 142 428 143 429
rect 141 428 142 429
rect 140 428 141 429
rect 127 428 128 429
rect 126 428 127 429
rect 125 428 126 429
rect 124 428 125 429
rect 123 428 124 429
rect 122 428 123 429
rect 121 428 122 429
rect 120 428 121 429
rect 119 428 120 429
rect 118 428 119 429
rect 117 428 118 429
rect 116 428 117 429
rect 115 428 116 429
rect 114 428 115 429
rect 113 428 114 429
rect 112 428 113 429
rect 111 428 112 429
rect 110 428 111 429
rect 109 428 110 429
rect 108 428 109 429
rect 107 428 108 429
rect 106 428 107 429
rect 105 428 106 429
rect 104 428 105 429
rect 103 428 104 429
rect 183 429 184 430
rect 182 429 183 430
rect 181 429 182 430
rect 180 429 181 430
rect 179 429 180 430
rect 178 429 179 430
rect 177 429 178 430
rect 176 429 177 430
rect 175 429 176 430
rect 174 429 175 430
rect 173 429 174 430
rect 172 429 173 430
rect 165 429 166 430
rect 164 429 165 430
rect 163 429 164 430
rect 153 429 154 430
rect 152 429 153 430
rect 151 429 152 430
rect 150 429 151 430
rect 149 429 150 430
rect 148 429 149 430
rect 147 429 148 430
rect 146 429 147 430
rect 145 429 146 430
rect 144 429 145 430
rect 143 429 144 430
rect 142 429 143 430
rect 141 429 142 430
rect 127 429 128 430
rect 126 429 127 430
rect 125 429 126 430
rect 124 429 125 430
rect 123 429 124 430
rect 122 429 123 430
rect 121 429 122 430
rect 120 429 121 430
rect 119 429 120 430
rect 118 429 119 430
rect 117 429 118 430
rect 116 429 117 430
rect 115 429 116 430
rect 114 429 115 430
rect 113 429 114 430
rect 112 429 113 430
rect 111 429 112 430
rect 110 429 111 430
rect 109 429 110 430
rect 108 429 109 430
rect 107 429 108 430
rect 106 429 107 430
rect 105 429 106 430
rect 104 429 105 430
rect 103 429 104 430
rect 196 430 197 431
rect 195 430 196 431
rect 194 430 195 431
rect 193 430 194 431
rect 192 430 193 431
rect 191 430 192 431
rect 190 430 191 431
rect 189 430 190 431
rect 183 430 184 431
rect 182 430 183 431
rect 181 430 182 431
rect 180 430 181 431
rect 179 430 180 431
rect 178 430 179 431
rect 177 430 178 431
rect 176 430 177 431
rect 175 430 176 431
rect 174 430 175 431
rect 173 430 174 431
rect 172 430 173 431
rect 165 430 166 431
rect 164 430 165 431
rect 163 430 164 431
rect 153 430 154 431
rect 152 430 153 431
rect 151 430 152 431
rect 150 430 151 431
rect 149 430 150 431
rect 148 430 149 431
rect 147 430 148 431
rect 146 430 147 431
rect 145 430 146 431
rect 144 430 145 431
rect 143 430 144 431
rect 142 430 143 431
rect 127 430 128 431
rect 126 430 127 431
rect 125 430 126 431
rect 124 430 125 431
rect 123 430 124 431
rect 122 430 123 431
rect 121 430 122 431
rect 120 430 121 431
rect 119 430 120 431
rect 118 430 119 431
rect 117 430 118 431
rect 116 430 117 431
rect 115 430 116 431
rect 114 430 115 431
rect 113 430 114 431
rect 112 430 113 431
rect 111 430 112 431
rect 110 430 111 431
rect 109 430 110 431
rect 108 430 109 431
rect 107 430 108 431
rect 106 430 107 431
rect 105 430 106 431
rect 104 430 105 431
rect 103 430 104 431
rect 197 431 198 432
rect 196 431 197 432
rect 195 431 196 432
rect 194 431 195 432
rect 193 431 194 432
rect 192 431 193 432
rect 191 431 192 432
rect 190 431 191 432
rect 189 431 190 432
rect 183 431 184 432
rect 182 431 183 432
rect 181 431 182 432
rect 180 431 181 432
rect 179 431 180 432
rect 178 431 179 432
rect 177 431 178 432
rect 176 431 177 432
rect 175 431 176 432
rect 174 431 175 432
rect 173 431 174 432
rect 172 431 173 432
rect 165 431 166 432
rect 164 431 165 432
rect 163 431 164 432
rect 153 431 154 432
rect 152 431 153 432
rect 151 431 152 432
rect 150 431 151 432
rect 149 431 150 432
rect 148 431 149 432
rect 147 431 148 432
rect 146 431 147 432
rect 145 431 146 432
rect 144 431 145 432
rect 143 431 144 432
rect 127 431 128 432
rect 126 431 127 432
rect 125 431 126 432
rect 124 431 125 432
rect 123 431 124 432
rect 122 431 123 432
rect 121 431 122 432
rect 120 431 121 432
rect 119 431 120 432
rect 118 431 119 432
rect 117 431 118 432
rect 116 431 117 432
rect 115 431 116 432
rect 114 431 115 432
rect 113 431 114 432
rect 112 431 113 432
rect 111 431 112 432
rect 110 431 111 432
rect 109 431 110 432
rect 108 431 109 432
rect 107 431 108 432
rect 106 431 107 432
rect 105 431 106 432
rect 104 431 105 432
rect 196 432 197 433
rect 195 432 196 433
rect 194 432 195 433
rect 193 432 194 433
rect 192 432 193 433
rect 191 432 192 433
rect 190 432 191 433
rect 189 432 190 433
rect 174 432 175 433
rect 173 432 174 433
rect 172 432 173 433
rect 165 432 166 433
rect 164 432 165 433
rect 163 432 164 433
rect 153 432 154 433
rect 152 432 153 433
rect 151 432 152 433
rect 150 432 151 433
rect 149 432 150 433
rect 148 432 149 433
rect 147 432 148 433
rect 146 432 147 433
rect 145 432 146 433
rect 144 432 145 433
rect 127 432 128 433
rect 126 432 127 433
rect 125 432 126 433
rect 124 432 125 433
rect 123 432 124 433
rect 122 432 123 433
rect 121 432 122 433
rect 120 432 121 433
rect 119 432 120 433
rect 118 432 119 433
rect 117 432 118 433
rect 116 432 117 433
rect 115 432 116 433
rect 114 432 115 433
rect 113 432 114 433
rect 112 432 113 433
rect 111 432 112 433
rect 110 432 111 433
rect 109 432 110 433
rect 108 432 109 433
rect 107 432 108 433
rect 106 432 107 433
rect 105 432 106 433
rect 174 433 175 434
rect 173 433 174 434
rect 172 433 173 434
rect 165 433 166 434
rect 164 433 165 434
rect 163 433 164 434
rect 153 433 154 434
rect 152 433 153 434
rect 151 433 152 434
rect 150 433 151 434
rect 149 433 150 434
rect 148 433 149 434
rect 147 433 148 434
rect 146 433 147 434
rect 145 433 146 434
rect 144 433 145 434
rect 127 433 128 434
rect 126 433 127 434
rect 125 433 126 434
rect 124 433 125 434
rect 123 433 124 434
rect 122 433 123 434
rect 121 433 122 434
rect 120 433 121 434
rect 119 433 120 434
rect 118 433 119 434
rect 117 433 118 434
rect 116 433 117 434
rect 115 433 116 434
rect 114 433 115 434
rect 113 433 114 434
rect 112 433 113 434
rect 111 433 112 434
rect 110 433 111 434
rect 109 433 110 434
rect 108 433 109 434
rect 107 433 108 434
rect 106 433 107 434
rect 196 434 197 435
rect 195 434 196 435
rect 194 434 195 435
rect 193 434 194 435
rect 192 434 193 435
rect 191 434 192 435
rect 174 434 175 435
rect 173 434 174 435
rect 172 434 173 435
rect 165 434 166 435
rect 164 434 165 435
rect 163 434 164 435
rect 153 434 154 435
rect 152 434 153 435
rect 151 434 152 435
rect 150 434 151 435
rect 149 434 150 435
rect 148 434 149 435
rect 147 434 148 435
rect 146 434 147 435
rect 145 434 146 435
rect 127 434 128 435
rect 126 434 127 435
rect 125 434 126 435
rect 124 434 125 435
rect 123 434 124 435
rect 122 434 123 435
rect 121 434 122 435
rect 120 434 121 435
rect 119 434 120 435
rect 118 434 119 435
rect 117 434 118 435
rect 116 434 117 435
rect 115 434 116 435
rect 114 434 115 435
rect 113 434 114 435
rect 112 434 113 435
rect 111 434 112 435
rect 110 434 111 435
rect 109 434 110 435
rect 108 434 109 435
rect 107 434 108 435
rect 197 435 198 436
rect 196 435 197 436
rect 195 435 196 436
rect 194 435 195 436
rect 193 435 194 436
rect 192 435 193 436
rect 191 435 192 436
rect 174 435 175 436
rect 173 435 174 436
rect 172 435 173 436
rect 171 435 172 436
rect 170 435 171 436
rect 169 435 170 436
rect 168 435 169 436
rect 167 435 168 436
rect 166 435 167 436
rect 165 435 166 436
rect 164 435 165 436
rect 163 435 164 436
rect 153 435 154 436
rect 152 435 153 436
rect 151 435 152 436
rect 150 435 151 436
rect 149 435 150 436
rect 148 435 149 436
rect 147 435 148 436
rect 146 435 147 436
rect 127 435 128 436
rect 126 435 127 436
rect 125 435 126 436
rect 124 435 125 436
rect 123 435 124 436
rect 122 435 123 436
rect 121 435 122 436
rect 120 435 121 436
rect 119 435 120 436
rect 118 435 119 436
rect 117 435 118 436
rect 116 435 117 436
rect 115 435 116 436
rect 114 435 115 436
rect 113 435 114 436
rect 112 435 113 436
rect 111 435 112 436
rect 110 435 111 436
rect 109 435 110 436
rect 108 435 109 436
rect 192 436 193 437
rect 191 436 192 437
rect 174 436 175 437
rect 173 436 174 437
rect 172 436 173 437
rect 171 436 172 437
rect 170 436 171 437
rect 169 436 170 437
rect 168 436 169 437
rect 167 436 168 437
rect 166 436 167 437
rect 165 436 166 437
rect 164 436 165 437
rect 163 436 164 437
rect 153 436 154 437
rect 152 436 153 437
rect 151 436 152 437
rect 150 436 151 437
rect 149 436 150 437
rect 148 436 149 437
rect 147 436 148 437
rect 192 437 193 438
rect 191 437 192 438
rect 174 437 175 438
rect 173 437 174 438
rect 172 437 173 438
rect 171 437 172 438
rect 170 437 171 438
rect 169 437 170 438
rect 168 437 169 438
rect 167 437 168 438
rect 166 437 167 438
rect 165 437 166 438
rect 164 437 165 438
rect 163 437 164 438
rect 153 437 154 438
rect 152 437 153 438
rect 151 437 152 438
rect 150 437 151 438
rect 149 437 150 438
rect 148 437 149 438
rect 196 438 197 439
rect 195 438 196 439
rect 194 438 195 439
rect 193 438 194 439
rect 192 438 193 439
rect 191 438 192 439
rect 174 438 175 439
rect 173 438 174 439
rect 172 438 173 439
rect 170 438 171 439
rect 169 438 170 439
rect 168 438 169 439
rect 167 438 168 439
rect 166 438 167 439
rect 165 438 166 439
rect 164 438 165 439
rect 163 438 164 439
rect 153 438 154 439
rect 152 438 153 439
rect 151 438 152 439
rect 150 438 151 439
rect 149 438 150 439
rect 197 439 198 440
rect 196 439 197 440
rect 195 439 196 440
rect 194 439 195 440
rect 193 439 194 440
rect 192 439 193 440
rect 191 439 192 440
rect 174 439 175 440
rect 173 439 174 440
rect 172 439 173 440
rect 167 439 168 440
rect 166 439 167 440
rect 165 439 166 440
rect 164 439 165 440
rect 163 439 164 440
rect 153 439 154 440
rect 152 439 153 440
rect 151 439 152 440
rect 150 439 151 440
rect 149 439 150 440
rect 192 440 193 441
rect 174 440 175 441
rect 173 440 174 441
rect 172 440 173 441
rect 153 440 154 441
rect 152 440 153 441
rect 151 440 152 441
rect 150 440 151 441
rect 196 441 197 442
rect 193 441 194 442
rect 192 441 193 442
rect 174 441 175 442
rect 173 441 174 442
rect 172 441 173 442
rect 153 441 154 442
rect 152 441 153 442
rect 151 441 152 442
rect 197 442 198 443
rect 196 442 197 443
rect 194 442 195 443
rect 193 442 194 443
rect 192 442 193 443
rect 191 442 192 443
rect 174 442 175 443
rect 173 442 174 443
rect 172 442 173 443
rect 153 442 154 443
rect 152 442 153 443
rect 197 443 198 444
rect 196 443 197 444
rect 195 443 196 444
rect 194 443 195 444
rect 193 443 194 444
rect 192 443 193 444
rect 191 443 192 444
rect 153 443 154 444
rect 152 443 153 444
rect 196 444 197 445
rect 195 444 196 445
rect 194 444 195 445
rect 192 444 193 445
rect 191 444 192 445
rect 196 445 197 446
rect 195 445 196 446
rect 194 445 195 446
rect 192 446 193 447
rect 191 446 192 447
rect 196 447 197 448
rect 195 447 196 448
rect 194 447 195 448
rect 193 447 194 448
rect 192 447 193 448
rect 191 447 192 448
rect 190 447 191 448
rect 197 448 198 449
rect 196 448 197 449
rect 195 448 196 449
rect 194 448 195 449
rect 193 448 194 449
rect 192 448 193 449
rect 191 448 192 449
rect 190 448 191 449
rect 189 448 190 449
rect 197 449 198 450
rect 196 449 197 450
rect 192 449 193 450
rect 191 449 192 450
rect 196 450 197 451
rect 196 451 197 452
rect 195 451 196 452
rect 194 451 195 452
rect 193 451 194 452
rect 192 451 193 452
rect 191 451 192 452
rect 189 451 190 452
rect 188 451 189 452
rect 197 452 198 453
rect 196 452 197 453
rect 195 452 196 453
rect 194 452 195 453
rect 193 452 194 453
rect 192 452 193 453
rect 191 452 192 453
rect 189 452 190 453
rect 188 452 189 453
rect 173 453 174 454
rect 172 453 173 454
rect 171 453 172 454
rect 149 453 150 454
rect 148 453 149 454
rect 147 453 148 454
rect 146 453 147 454
rect 145 453 146 454
rect 144 453 145 454
rect 143 453 144 454
rect 142 453 143 454
rect 141 453 142 454
rect 140 453 141 454
rect 139 453 140 454
rect 138 453 139 454
rect 137 453 138 454
rect 136 453 137 454
rect 135 453 136 454
rect 134 453 135 454
rect 133 453 134 454
rect 132 453 133 454
rect 131 453 132 454
rect 130 453 131 454
rect 129 453 130 454
rect 128 453 129 454
rect 127 453 128 454
rect 126 453 127 454
rect 125 453 126 454
rect 124 453 125 454
rect 123 453 124 454
rect 122 453 123 454
rect 121 453 122 454
rect 120 453 121 454
rect 119 453 120 454
rect 118 453 119 454
rect 117 453 118 454
rect 116 453 117 454
rect 115 453 116 454
rect 114 453 115 454
rect 113 453 114 454
rect 112 453 113 454
rect 111 453 112 454
rect 110 453 111 454
rect 109 453 110 454
rect 108 453 109 454
rect 107 453 108 454
rect 106 453 107 454
rect 105 453 106 454
rect 104 453 105 454
rect 103 453 104 454
rect 102 453 103 454
rect 192 454 193 455
rect 191 454 192 455
rect 173 454 174 455
rect 172 454 173 455
rect 171 454 172 455
rect 170 454 171 455
rect 149 454 150 455
rect 148 454 149 455
rect 147 454 148 455
rect 146 454 147 455
rect 145 454 146 455
rect 144 454 145 455
rect 143 454 144 455
rect 142 454 143 455
rect 141 454 142 455
rect 140 454 141 455
rect 139 454 140 455
rect 138 454 139 455
rect 137 454 138 455
rect 136 454 137 455
rect 135 454 136 455
rect 134 454 135 455
rect 133 454 134 455
rect 132 454 133 455
rect 131 454 132 455
rect 130 454 131 455
rect 129 454 130 455
rect 128 454 129 455
rect 127 454 128 455
rect 126 454 127 455
rect 125 454 126 455
rect 124 454 125 455
rect 123 454 124 455
rect 122 454 123 455
rect 121 454 122 455
rect 120 454 121 455
rect 119 454 120 455
rect 118 454 119 455
rect 117 454 118 455
rect 116 454 117 455
rect 115 454 116 455
rect 114 454 115 455
rect 113 454 114 455
rect 112 454 113 455
rect 111 454 112 455
rect 110 454 111 455
rect 109 454 110 455
rect 108 454 109 455
rect 107 454 108 455
rect 106 454 107 455
rect 105 454 106 455
rect 104 454 105 455
rect 103 454 104 455
rect 102 454 103 455
rect 196 455 197 456
rect 195 455 196 456
rect 194 455 195 456
rect 193 455 194 456
rect 192 455 193 456
rect 191 455 192 456
rect 190 455 191 456
rect 189 455 190 456
rect 173 455 174 456
rect 172 455 173 456
rect 171 455 172 456
rect 170 455 171 456
rect 167 455 168 456
rect 166 455 167 456
rect 165 455 166 456
rect 164 455 165 456
rect 149 455 150 456
rect 148 455 149 456
rect 147 455 148 456
rect 146 455 147 456
rect 145 455 146 456
rect 144 455 145 456
rect 143 455 144 456
rect 142 455 143 456
rect 141 455 142 456
rect 140 455 141 456
rect 139 455 140 456
rect 138 455 139 456
rect 137 455 138 456
rect 136 455 137 456
rect 135 455 136 456
rect 134 455 135 456
rect 133 455 134 456
rect 132 455 133 456
rect 131 455 132 456
rect 130 455 131 456
rect 129 455 130 456
rect 128 455 129 456
rect 127 455 128 456
rect 126 455 127 456
rect 125 455 126 456
rect 124 455 125 456
rect 123 455 124 456
rect 122 455 123 456
rect 121 455 122 456
rect 120 455 121 456
rect 119 455 120 456
rect 118 455 119 456
rect 117 455 118 456
rect 116 455 117 456
rect 115 455 116 456
rect 114 455 115 456
rect 113 455 114 456
rect 112 455 113 456
rect 111 455 112 456
rect 110 455 111 456
rect 109 455 110 456
rect 108 455 109 456
rect 107 455 108 456
rect 106 455 107 456
rect 105 455 106 456
rect 104 455 105 456
rect 103 455 104 456
rect 102 455 103 456
rect 197 456 198 457
rect 196 456 197 457
rect 195 456 196 457
rect 194 456 195 457
rect 193 456 194 457
rect 192 456 193 457
rect 191 456 192 457
rect 190 456 191 457
rect 189 456 190 457
rect 173 456 174 457
rect 172 456 173 457
rect 171 456 172 457
rect 170 456 171 457
rect 168 456 169 457
rect 167 456 168 457
rect 166 456 167 457
rect 165 456 166 457
rect 164 456 165 457
rect 163 456 164 457
rect 149 456 150 457
rect 148 456 149 457
rect 147 456 148 457
rect 146 456 147 457
rect 145 456 146 457
rect 144 456 145 457
rect 143 456 144 457
rect 142 456 143 457
rect 141 456 142 457
rect 140 456 141 457
rect 139 456 140 457
rect 138 456 139 457
rect 137 456 138 457
rect 136 456 137 457
rect 135 456 136 457
rect 134 456 135 457
rect 133 456 134 457
rect 132 456 133 457
rect 131 456 132 457
rect 130 456 131 457
rect 129 456 130 457
rect 128 456 129 457
rect 127 456 128 457
rect 126 456 127 457
rect 125 456 126 457
rect 124 456 125 457
rect 123 456 124 457
rect 122 456 123 457
rect 121 456 122 457
rect 120 456 121 457
rect 119 456 120 457
rect 118 456 119 457
rect 117 456 118 457
rect 116 456 117 457
rect 115 456 116 457
rect 114 456 115 457
rect 113 456 114 457
rect 112 456 113 457
rect 111 456 112 457
rect 110 456 111 457
rect 109 456 110 457
rect 108 456 109 457
rect 107 456 108 457
rect 106 456 107 457
rect 105 456 106 457
rect 104 456 105 457
rect 103 456 104 457
rect 102 456 103 457
rect 197 457 198 458
rect 196 457 197 458
rect 192 457 193 458
rect 191 457 192 458
rect 183 457 184 458
rect 182 457 183 458
rect 181 457 182 458
rect 180 457 181 458
rect 179 457 180 458
rect 178 457 179 458
rect 173 457 174 458
rect 172 457 173 458
rect 171 457 172 458
rect 170 457 171 458
rect 168 457 169 458
rect 167 457 168 458
rect 166 457 167 458
rect 165 457 166 458
rect 164 457 165 458
rect 163 457 164 458
rect 162 457 163 458
rect 149 457 150 458
rect 148 457 149 458
rect 147 457 148 458
rect 146 457 147 458
rect 145 457 146 458
rect 144 457 145 458
rect 143 457 144 458
rect 142 457 143 458
rect 141 457 142 458
rect 140 457 141 458
rect 139 457 140 458
rect 138 457 139 458
rect 137 457 138 458
rect 136 457 137 458
rect 135 457 136 458
rect 134 457 135 458
rect 133 457 134 458
rect 132 457 133 458
rect 131 457 132 458
rect 130 457 131 458
rect 129 457 130 458
rect 128 457 129 458
rect 127 457 128 458
rect 126 457 127 458
rect 125 457 126 458
rect 124 457 125 458
rect 123 457 124 458
rect 122 457 123 458
rect 121 457 122 458
rect 120 457 121 458
rect 119 457 120 458
rect 118 457 119 458
rect 117 457 118 458
rect 116 457 117 458
rect 115 457 116 458
rect 114 457 115 458
rect 113 457 114 458
rect 112 457 113 458
rect 111 457 112 458
rect 110 457 111 458
rect 109 457 110 458
rect 108 457 109 458
rect 107 457 108 458
rect 106 457 107 458
rect 105 457 106 458
rect 104 457 105 458
rect 103 457 104 458
rect 102 457 103 458
rect 196 458 197 459
rect 183 458 184 459
rect 182 458 183 459
rect 181 458 182 459
rect 180 458 181 459
rect 179 458 180 459
rect 178 458 179 459
rect 173 458 174 459
rect 172 458 173 459
rect 171 458 172 459
rect 170 458 171 459
rect 169 458 170 459
rect 168 458 169 459
rect 167 458 168 459
rect 166 458 167 459
rect 165 458 166 459
rect 164 458 165 459
rect 163 458 164 459
rect 162 458 163 459
rect 149 458 150 459
rect 148 458 149 459
rect 147 458 148 459
rect 146 458 147 459
rect 145 458 146 459
rect 144 458 145 459
rect 143 458 144 459
rect 142 458 143 459
rect 141 458 142 459
rect 140 458 141 459
rect 139 458 140 459
rect 138 458 139 459
rect 137 458 138 459
rect 136 458 137 459
rect 135 458 136 459
rect 134 458 135 459
rect 133 458 134 459
rect 132 458 133 459
rect 131 458 132 459
rect 130 458 131 459
rect 129 458 130 459
rect 128 458 129 459
rect 127 458 128 459
rect 126 458 127 459
rect 125 458 126 459
rect 124 458 125 459
rect 123 458 124 459
rect 122 458 123 459
rect 121 458 122 459
rect 120 458 121 459
rect 119 458 120 459
rect 118 458 119 459
rect 117 458 118 459
rect 116 458 117 459
rect 115 458 116 459
rect 114 458 115 459
rect 113 458 114 459
rect 112 458 113 459
rect 111 458 112 459
rect 110 458 111 459
rect 109 458 110 459
rect 108 458 109 459
rect 107 458 108 459
rect 106 458 107 459
rect 105 458 106 459
rect 104 458 105 459
rect 103 458 104 459
rect 102 458 103 459
rect 196 459 197 460
rect 195 459 196 460
rect 194 459 195 460
rect 193 459 194 460
rect 192 459 193 460
rect 191 459 192 460
rect 183 459 184 460
rect 182 459 183 460
rect 181 459 182 460
rect 180 459 181 460
rect 179 459 180 460
rect 178 459 179 460
rect 177 459 178 460
rect 176 459 177 460
rect 175 459 176 460
rect 174 459 175 460
rect 173 459 174 460
rect 172 459 173 460
rect 171 459 172 460
rect 170 459 171 460
rect 169 459 170 460
rect 168 459 169 460
rect 167 459 168 460
rect 166 459 167 460
rect 164 459 165 460
rect 163 459 164 460
rect 162 459 163 460
rect 161 459 162 460
rect 149 459 150 460
rect 148 459 149 460
rect 147 459 148 460
rect 146 459 147 460
rect 145 459 146 460
rect 144 459 145 460
rect 143 459 144 460
rect 142 459 143 460
rect 141 459 142 460
rect 140 459 141 460
rect 139 459 140 460
rect 138 459 139 460
rect 137 459 138 460
rect 136 459 137 460
rect 135 459 136 460
rect 134 459 135 460
rect 133 459 134 460
rect 132 459 133 460
rect 131 459 132 460
rect 130 459 131 460
rect 129 459 130 460
rect 128 459 129 460
rect 127 459 128 460
rect 126 459 127 460
rect 125 459 126 460
rect 124 459 125 460
rect 123 459 124 460
rect 122 459 123 460
rect 121 459 122 460
rect 120 459 121 460
rect 119 459 120 460
rect 118 459 119 460
rect 117 459 118 460
rect 116 459 117 460
rect 115 459 116 460
rect 114 459 115 460
rect 113 459 114 460
rect 112 459 113 460
rect 111 459 112 460
rect 110 459 111 460
rect 109 459 110 460
rect 108 459 109 460
rect 107 459 108 460
rect 106 459 107 460
rect 105 459 106 460
rect 104 459 105 460
rect 103 459 104 460
rect 102 459 103 460
rect 197 460 198 461
rect 196 460 197 461
rect 195 460 196 461
rect 194 460 195 461
rect 193 460 194 461
rect 192 460 193 461
rect 191 460 192 461
rect 183 460 184 461
rect 182 460 183 461
rect 181 460 182 461
rect 180 460 181 461
rect 179 460 180 461
rect 178 460 179 461
rect 177 460 178 461
rect 176 460 177 461
rect 175 460 176 461
rect 174 460 175 461
rect 173 460 174 461
rect 172 460 173 461
rect 171 460 172 461
rect 170 460 171 461
rect 169 460 170 461
rect 168 460 169 461
rect 167 460 168 461
rect 163 460 164 461
rect 162 460 163 461
rect 161 460 162 461
rect 149 460 150 461
rect 148 460 149 461
rect 147 460 148 461
rect 146 460 147 461
rect 145 460 146 461
rect 144 460 145 461
rect 143 460 144 461
rect 142 460 143 461
rect 141 460 142 461
rect 140 460 141 461
rect 139 460 140 461
rect 138 460 139 461
rect 137 460 138 461
rect 136 460 137 461
rect 135 460 136 461
rect 134 460 135 461
rect 133 460 134 461
rect 132 460 133 461
rect 131 460 132 461
rect 130 460 131 461
rect 129 460 130 461
rect 128 460 129 461
rect 127 460 128 461
rect 126 460 127 461
rect 125 460 126 461
rect 124 460 125 461
rect 123 460 124 461
rect 122 460 123 461
rect 121 460 122 461
rect 120 460 121 461
rect 119 460 120 461
rect 118 460 119 461
rect 117 460 118 461
rect 116 460 117 461
rect 115 460 116 461
rect 114 460 115 461
rect 113 460 114 461
rect 112 460 113 461
rect 111 460 112 461
rect 110 460 111 461
rect 109 460 110 461
rect 108 460 109 461
rect 107 460 108 461
rect 106 460 107 461
rect 105 460 106 461
rect 104 460 105 461
rect 103 460 104 461
rect 102 460 103 461
rect 197 461 198 462
rect 196 461 197 462
rect 183 461 184 462
rect 182 461 183 462
rect 181 461 182 462
rect 180 461 181 462
rect 176 461 177 462
rect 175 461 176 462
rect 174 461 175 462
rect 173 461 174 462
rect 172 461 173 462
rect 171 461 172 462
rect 170 461 171 462
rect 169 461 170 462
rect 168 461 169 462
rect 167 461 168 462
rect 163 461 164 462
rect 162 461 163 462
rect 161 461 162 462
rect 149 461 150 462
rect 148 461 149 462
rect 147 461 148 462
rect 146 461 147 462
rect 145 461 146 462
rect 144 461 145 462
rect 143 461 144 462
rect 142 461 143 462
rect 141 461 142 462
rect 140 461 141 462
rect 139 461 140 462
rect 138 461 139 462
rect 137 461 138 462
rect 136 461 137 462
rect 135 461 136 462
rect 134 461 135 462
rect 133 461 134 462
rect 132 461 133 462
rect 131 461 132 462
rect 130 461 131 462
rect 129 461 130 462
rect 128 461 129 462
rect 127 461 128 462
rect 126 461 127 462
rect 125 461 126 462
rect 124 461 125 462
rect 123 461 124 462
rect 122 461 123 462
rect 121 461 122 462
rect 120 461 121 462
rect 119 461 120 462
rect 118 461 119 462
rect 117 461 118 462
rect 116 461 117 462
rect 115 461 116 462
rect 114 461 115 462
rect 113 461 114 462
rect 112 461 113 462
rect 111 461 112 462
rect 110 461 111 462
rect 109 461 110 462
rect 108 461 109 462
rect 107 461 108 462
rect 106 461 107 462
rect 105 461 106 462
rect 104 461 105 462
rect 103 461 104 462
rect 102 461 103 462
rect 196 462 197 463
rect 183 462 184 463
rect 182 462 183 463
rect 181 462 182 463
rect 180 462 181 463
rect 173 462 174 463
rect 172 462 173 463
rect 171 462 172 463
rect 170 462 171 463
rect 169 462 170 463
rect 168 462 169 463
rect 167 462 168 463
rect 163 462 164 463
rect 162 462 163 463
rect 161 462 162 463
rect 149 462 150 463
rect 148 462 149 463
rect 147 462 148 463
rect 146 462 147 463
rect 145 462 146 463
rect 144 462 145 463
rect 143 462 144 463
rect 142 462 143 463
rect 141 462 142 463
rect 140 462 141 463
rect 139 462 140 463
rect 138 462 139 463
rect 137 462 138 463
rect 136 462 137 463
rect 135 462 136 463
rect 134 462 135 463
rect 133 462 134 463
rect 132 462 133 463
rect 131 462 132 463
rect 130 462 131 463
rect 129 462 130 463
rect 128 462 129 463
rect 127 462 128 463
rect 126 462 127 463
rect 125 462 126 463
rect 124 462 125 463
rect 123 462 124 463
rect 122 462 123 463
rect 121 462 122 463
rect 120 462 121 463
rect 119 462 120 463
rect 118 462 119 463
rect 117 462 118 463
rect 116 462 117 463
rect 115 462 116 463
rect 114 462 115 463
rect 113 462 114 463
rect 112 462 113 463
rect 111 462 112 463
rect 110 462 111 463
rect 109 462 110 463
rect 108 462 109 463
rect 107 462 108 463
rect 106 462 107 463
rect 105 462 106 463
rect 104 462 105 463
rect 103 462 104 463
rect 102 462 103 463
rect 197 463 198 464
rect 196 463 197 464
rect 195 463 196 464
rect 194 463 195 464
rect 193 463 194 464
rect 192 463 193 464
rect 191 463 192 464
rect 183 463 184 464
rect 182 463 183 464
rect 181 463 182 464
rect 180 463 181 464
rect 173 463 174 464
rect 172 463 173 464
rect 171 463 172 464
rect 170 463 171 464
rect 169 463 170 464
rect 168 463 169 464
rect 167 463 168 464
rect 163 463 164 464
rect 162 463 163 464
rect 161 463 162 464
rect 149 463 150 464
rect 148 463 149 464
rect 147 463 148 464
rect 146 463 147 464
rect 145 463 146 464
rect 144 463 145 464
rect 143 463 144 464
rect 142 463 143 464
rect 141 463 142 464
rect 140 463 141 464
rect 139 463 140 464
rect 138 463 139 464
rect 137 463 138 464
rect 136 463 137 464
rect 135 463 136 464
rect 134 463 135 464
rect 133 463 134 464
rect 132 463 133 464
rect 131 463 132 464
rect 130 463 131 464
rect 129 463 130 464
rect 128 463 129 464
rect 127 463 128 464
rect 126 463 127 464
rect 125 463 126 464
rect 124 463 125 464
rect 123 463 124 464
rect 122 463 123 464
rect 121 463 122 464
rect 120 463 121 464
rect 119 463 120 464
rect 118 463 119 464
rect 117 463 118 464
rect 116 463 117 464
rect 115 463 116 464
rect 114 463 115 464
rect 113 463 114 464
rect 112 463 113 464
rect 111 463 112 464
rect 110 463 111 464
rect 109 463 110 464
rect 108 463 109 464
rect 107 463 108 464
rect 106 463 107 464
rect 105 463 106 464
rect 104 463 105 464
rect 103 463 104 464
rect 102 463 103 464
rect 196 464 197 465
rect 195 464 196 465
rect 194 464 195 465
rect 193 464 194 465
rect 192 464 193 465
rect 191 464 192 465
rect 183 464 184 465
rect 182 464 183 465
rect 181 464 182 465
rect 180 464 181 465
rect 173 464 174 465
rect 172 464 173 465
rect 171 464 172 465
rect 170 464 171 465
rect 169 464 170 465
rect 168 464 169 465
rect 167 464 168 465
rect 166 464 167 465
rect 164 464 165 465
rect 163 464 164 465
rect 162 464 163 465
rect 149 464 150 465
rect 148 464 149 465
rect 147 464 148 465
rect 146 464 147 465
rect 145 464 146 465
rect 144 464 145 465
rect 143 464 144 465
rect 142 464 143 465
rect 141 464 142 465
rect 140 464 141 465
rect 139 464 140 465
rect 138 464 139 465
rect 137 464 138 465
rect 136 464 137 465
rect 135 464 136 465
rect 134 464 135 465
rect 133 464 134 465
rect 132 464 133 465
rect 131 464 132 465
rect 130 464 131 465
rect 129 464 130 465
rect 128 464 129 465
rect 127 464 128 465
rect 126 464 127 465
rect 125 464 126 465
rect 124 464 125 465
rect 123 464 124 465
rect 122 464 123 465
rect 121 464 122 465
rect 120 464 121 465
rect 119 464 120 465
rect 118 464 119 465
rect 117 464 118 465
rect 116 464 117 465
rect 115 464 116 465
rect 114 464 115 465
rect 113 464 114 465
rect 112 464 113 465
rect 111 464 112 465
rect 110 464 111 465
rect 109 464 110 465
rect 108 464 109 465
rect 107 464 108 465
rect 106 464 107 465
rect 105 464 106 465
rect 104 464 105 465
rect 103 464 104 465
rect 102 464 103 465
rect 183 465 184 466
rect 182 465 183 466
rect 181 465 182 466
rect 180 465 181 466
rect 173 465 174 466
rect 172 465 173 466
rect 171 465 172 466
rect 170 465 171 466
rect 168 465 169 466
rect 167 465 168 466
rect 166 465 167 466
rect 165 465 166 466
rect 164 465 165 466
rect 163 465 164 466
rect 162 465 163 466
rect 149 465 150 466
rect 148 465 149 466
rect 147 465 148 466
rect 146 465 147 466
rect 145 465 146 466
rect 144 465 145 466
rect 143 465 144 466
rect 142 465 143 466
rect 141 465 142 466
rect 140 465 141 466
rect 139 465 140 466
rect 138 465 139 466
rect 137 465 138 466
rect 136 465 137 466
rect 135 465 136 466
rect 134 465 135 466
rect 133 465 134 466
rect 132 465 133 466
rect 131 465 132 466
rect 130 465 131 466
rect 129 465 130 466
rect 128 465 129 466
rect 127 465 128 466
rect 126 465 127 466
rect 125 465 126 466
rect 124 465 125 466
rect 123 465 124 466
rect 122 465 123 466
rect 121 465 122 466
rect 120 465 121 466
rect 119 465 120 466
rect 118 465 119 466
rect 117 465 118 466
rect 116 465 117 466
rect 115 465 116 466
rect 114 465 115 466
rect 113 465 114 466
rect 112 465 113 466
rect 111 465 112 466
rect 110 465 111 466
rect 109 465 110 466
rect 108 465 109 466
rect 107 465 108 466
rect 106 465 107 466
rect 105 465 106 466
rect 104 465 105 466
rect 103 465 104 466
rect 102 465 103 466
rect 195 466 196 467
rect 194 466 195 467
rect 193 466 194 467
rect 192 466 193 467
rect 191 466 192 467
rect 190 466 191 467
rect 183 466 184 467
rect 182 466 183 467
rect 181 466 182 467
rect 180 466 181 467
rect 176 466 177 467
rect 175 466 176 467
rect 174 466 175 467
rect 173 466 174 467
rect 172 466 173 467
rect 171 466 172 467
rect 170 466 171 467
rect 168 466 169 467
rect 167 466 168 467
rect 166 466 167 467
rect 165 466 166 467
rect 164 466 165 467
rect 163 466 164 467
rect 149 466 150 467
rect 148 466 149 467
rect 147 466 148 467
rect 146 466 147 467
rect 145 466 146 467
rect 144 466 145 467
rect 143 466 144 467
rect 142 466 143 467
rect 141 466 142 467
rect 140 466 141 467
rect 139 466 140 467
rect 138 466 139 467
rect 137 466 138 467
rect 136 466 137 467
rect 135 466 136 467
rect 134 466 135 467
rect 133 466 134 467
rect 132 466 133 467
rect 131 466 132 467
rect 130 466 131 467
rect 129 466 130 467
rect 128 466 129 467
rect 127 466 128 467
rect 126 466 127 467
rect 125 466 126 467
rect 124 466 125 467
rect 123 466 124 467
rect 122 466 123 467
rect 121 466 122 467
rect 120 466 121 467
rect 119 466 120 467
rect 118 466 119 467
rect 117 466 118 467
rect 116 466 117 467
rect 115 466 116 467
rect 114 466 115 467
rect 113 466 114 467
rect 112 466 113 467
rect 111 466 112 467
rect 110 466 111 467
rect 109 466 110 467
rect 108 466 109 467
rect 107 466 108 467
rect 106 466 107 467
rect 105 466 106 467
rect 104 466 105 467
rect 103 466 104 467
rect 102 466 103 467
rect 196 467 197 468
rect 195 467 196 468
rect 194 467 195 468
rect 193 467 194 468
rect 192 467 193 468
rect 191 467 192 468
rect 190 467 191 468
rect 189 467 190 468
rect 183 467 184 468
rect 182 467 183 468
rect 181 467 182 468
rect 180 467 181 468
rect 176 467 177 468
rect 175 467 176 468
rect 174 467 175 468
rect 173 467 174 468
rect 172 467 173 468
rect 171 467 172 468
rect 170 467 171 468
rect 167 467 168 468
rect 166 467 167 468
rect 165 467 166 468
rect 164 467 165 468
rect 163 467 164 468
rect 149 467 150 468
rect 148 467 149 468
rect 147 467 148 468
rect 146 467 147 468
rect 145 467 146 468
rect 144 467 145 468
rect 143 467 144 468
rect 142 467 143 468
rect 141 467 142 468
rect 140 467 141 468
rect 139 467 140 468
rect 138 467 139 468
rect 137 467 138 468
rect 136 467 137 468
rect 135 467 136 468
rect 134 467 135 468
rect 133 467 134 468
rect 132 467 133 468
rect 131 467 132 468
rect 130 467 131 468
rect 129 467 130 468
rect 128 467 129 468
rect 127 467 128 468
rect 126 467 127 468
rect 125 467 126 468
rect 124 467 125 468
rect 123 467 124 468
rect 122 467 123 468
rect 121 467 122 468
rect 120 467 121 468
rect 119 467 120 468
rect 118 467 119 468
rect 117 467 118 468
rect 116 467 117 468
rect 115 467 116 468
rect 114 467 115 468
rect 113 467 114 468
rect 112 467 113 468
rect 111 467 112 468
rect 110 467 111 468
rect 109 467 110 468
rect 108 467 109 468
rect 107 467 108 468
rect 106 467 107 468
rect 105 467 106 468
rect 104 467 105 468
rect 103 467 104 468
rect 102 467 103 468
rect 196 468 197 469
rect 195 468 196 469
rect 194 468 195 469
rect 193 468 194 469
rect 192 468 193 469
rect 191 468 192 469
rect 190 468 191 469
rect 189 468 190 469
rect 183 468 184 469
rect 182 468 183 469
rect 181 468 182 469
rect 180 468 181 469
rect 176 468 177 469
rect 175 468 176 469
rect 174 468 175 469
rect 173 468 174 469
rect 172 468 173 469
rect 171 468 172 469
rect 170 468 171 469
rect 166 468 167 469
rect 165 468 166 469
rect 164 468 165 469
rect 149 468 150 469
rect 148 468 149 469
rect 147 468 148 469
rect 146 468 147 469
rect 145 468 146 469
rect 144 468 145 469
rect 143 468 144 469
rect 142 468 143 469
rect 141 468 142 469
rect 140 468 141 469
rect 139 468 140 469
rect 138 468 139 469
rect 137 468 138 469
rect 136 468 137 469
rect 135 468 136 469
rect 134 468 135 469
rect 133 468 134 469
rect 132 468 133 469
rect 131 468 132 469
rect 130 468 131 469
rect 129 468 130 469
rect 128 468 129 469
rect 127 468 128 469
rect 126 468 127 469
rect 125 468 126 469
rect 124 468 125 469
rect 123 468 124 469
rect 122 468 123 469
rect 121 468 122 469
rect 120 468 121 469
rect 119 468 120 469
rect 118 468 119 469
rect 117 468 118 469
rect 116 468 117 469
rect 115 468 116 469
rect 114 468 115 469
rect 113 468 114 469
rect 112 468 113 469
rect 111 468 112 469
rect 110 468 111 469
rect 109 468 110 469
rect 108 468 109 469
rect 107 468 108 469
rect 106 468 107 469
rect 105 468 106 469
rect 104 468 105 469
rect 103 468 104 469
rect 102 468 103 469
rect 197 469 198 470
rect 196 469 197 470
rect 192 469 193 470
rect 191 469 192 470
rect 183 469 184 470
rect 182 469 183 470
rect 181 469 182 470
rect 180 469 181 470
rect 176 469 177 470
rect 175 469 176 470
rect 174 469 175 470
rect 172 469 173 470
rect 171 469 172 470
rect 170 469 171 470
rect 149 469 150 470
rect 148 469 149 470
rect 147 469 148 470
rect 146 469 147 470
rect 145 469 146 470
rect 144 469 145 470
rect 143 469 144 470
rect 142 469 143 470
rect 141 469 142 470
rect 140 469 141 470
rect 139 469 140 470
rect 138 469 139 470
rect 137 469 138 470
rect 136 469 137 470
rect 135 469 136 470
rect 134 469 135 470
rect 133 469 134 470
rect 132 469 133 470
rect 131 469 132 470
rect 130 469 131 470
rect 129 469 130 470
rect 128 469 129 470
rect 127 469 128 470
rect 126 469 127 470
rect 125 469 126 470
rect 124 469 125 470
rect 123 469 124 470
rect 122 469 123 470
rect 121 469 122 470
rect 120 469 121 470
rect 119 469 120 470
rect 118 469 119 470
rect 117 469 118 470
rect 116 469 117 470
rect 115 469 116 470
rect 114 469 115 470
rect 113 469 114 470
rect 112 469 113 470
rect 111 469 112 470
rect 110 469 111 470
rect 109 469 110 470
rect 108 469 109 470
rect 107 469 108 470
rect 106 469 107 470
rect 105 469 106 470
rect 104 469 105 470
rect 103 469 104 470
rect 102 469 103 470
rect 195 470 196 471
rect 194 470 195 471
rect 193 470 194 471
rect 183 470 184 471
rect 182 470 183 471
rect 181 470 182 471
rect 180 470 181 471
rect 176 470 177 471
rect 175 470 176 471
rect 174 470 175 471
rect 172 470 173 471
rect 171 470 172 471
rect 170 470 171 471
rect 149 470 150 471
rect 148 470 149 471
rect 147 470 148 471
rect 146 470 147 471
rect 145 470 146 471
rect 144 470 145 471
rect 143 470 144 471
rect 142 470 143 471
rect 141 470 142 471
rect 140 470 141 471
rect 139 470 140 471
rect 138 470 139 471
rect 137 470 138 471
rect 136 470 137 471
rect 135 470 136 471
rect 134 470 135 471
rect 133 470 134 471
rect 132 470 133 471
rect 131 470 132 471
rect 130 470 131 471
rect 129 470 130 471
rect 128 470 129 471
rect 127 470 128 471
rect 126 470 127 471
rect 125 470 126 471
rect 124 470 125 471
rect 123 470 124 471
rect 122 470 123 471
rect 121 470 122 471
rect 120 470 121 471
rect 119 470 120 471
rect 118 470 119 471
rect 117 470 118 471
rect 116 470 117 471
rect 115 470 116 471
rect 114 470 115 471
rect 113 470 114 471
rect 112 470 113 471
rect 111 470 112 471
rect 110 470 111 471
rect 109 470 110 471
rect 108 470 109 471
rect 107 470 108 471
rect 106 470 107 471
rect 105 470 106 471
rect 104 470 105 471
rect 103 470 104 471
rect 102 470 103 471
rect 196 471 197 472
rect 195 471 196 472
rect 194 471 195 472
rect 193 471 194 472
rect 192 471 193 472
rect 191 471 192 472
rect 183 471 184 472
rect 182 471 183 472
rect 181 471 182 472
rect 180 471 181 472
rect 176 471 177 472
rect 175 471 176 472
rect 174 471 175 472
rect 173 471 174 472
rect 149 471 150 472
rect 148 471 149 472
rect 147 471 148 472
rect 146 471 147 472
rect 145 471 146 472
rect 144 471 145 472
rect 143 471 144 472
rect 142 471 143 472
rect 141 471 142 472
rect 140 471 141 472
rect 139 471 140 472
rect 138 471 139 472
rect 137 471 138 472
rect 136 471 137 472
rect 135 471 136 472
rect 134 471 135 472
rect 133 471 134 472
rect 132 471 133 472
rect 131 471 132 472
rect 130 471 131 472
rect 129 471 130 472
rect 128 471 129 472
rect 127 471 128 472
rect 126 471 127 472
rect 125 471 126 472
rect 124 471 125 472
rect 123 471 124 472
rect 122 471 123 472
rect 121 471 122 472
rect 120 471 121 472
rect 119 471 120 472
rect 118 471 119 472
rect 117 471 118 472
rect 116 471 117 472
rect 115 471 116 472
rect 114 471 115 472
rect 113 471 114 472
rect 112 471 113 472
rect 111 471 112 472
rect 110 471 111 472
rect 109 471 110 472
rect 108 471 109 472
rect 107 471 108 472
rect 106 471 107 472
rect 105 471 106 472
rect 104 471 105 472
rect 103 471 104 472
rect 102 471 103 472
rect 196 472 197 473
rect 195 472 196 473
rect 194 472 195 473
rect 193 472 194 473
rect 192 472 193 473
rect 191 472 192 473
rect 183 472 184 473
rect 182 472 183 473
rect 181 472 182 473
rect 180 472 181 473
rect 178 472 179 473
rect 177 472 178 473
rect 176 472 177 473
rect 175 472 176 473
rect 174 472 175 473
rect 173 472 174 473
rect 172 472 173 473
rect 171 472 172 473
rect 170 472 171 473
rect 169 472 170 473
rect 168 472 169 473
rect 167 472 168 473
rect 166 472 167 473
rect 165 472 166 473
rect 164 472 165 473
rect 163 472 164 473
rect 162 472 163 473
rect 149 472 150 473
rect 148 472 149 473
rect 147 472 148 473
rect 146 472 147 473
rect 145 472 146 473
rect 144 472 145 473
rect 143 472 144 473
rect 142 472 143 473
rect 141 472 142 473
rect 140 472 141 473
rect 139 472 140 473
rect 138 472 139 473
rect 137 472 138 473
rect 136 472 137 473
rect 135 472 136 473
rect 134 472 135 473
rect 133 472 134 473
rect 132 472 133 473
rect 131 472 132 473
rect 130 472 131 473
rect 129 472 130 473
rect 128 472 129 473
rect 127 472 128 473
rect 126 472 127 473
rect 125 472 126 473
rect 124 472 125 473
rect 123 472 124 473
rect 122 472 123 473
rect 121 472 122 473
rect 120 472 121 473
rect 119 472 120 473
rect 118 472 119 473
rect 117 472 118 473
rect 116 472 117 473
rect 115 472 116 473
rect 114 472 115 473
rect 113 472 114 473
rect 112 472 113 473
rect 111 472 112 473
rect 110 472 111 473
rect 109 472 110 473
rect 108 472 109 473
rect 107 472 108 473
rect 106 472 107 473
rect 105 472 106 473
rect 104 472 105 473
rect 103 472 104 473
rect 102 472 103 473
rect 197 473 198 474
rect 196 473 197 474
rect 194 473 195 474
rect 192 473 193 474
rect 191 473 192 474
rect 183 473 184 474
rect 182 473 183 474
rect 181 473 182 474
rect 180 473 181 474
rect 178 473 179 474
rect 177 473 178 474
rect 176 473 177 474
rect 175 473 176 474
rect 174 473 175 474
rect 173 473 174 474
rect 172 473 173 474
rect 171 473 172 474
rect 170 473 171 474
rect 169 473 170 474
rect 168 473 169 474
rect 167 473 168 474
rect 166 473 167 474
rect 165 473 166 474
rect 164 473 165 474
rect 163 473 164 474
rect 162 473 163 474
rect 149 473 150 474
rect 148 473 149 474
rect 147 473 148 474
rect 146 473 147 474
rect 145 473 146 474
rect 144 473 145 474
rect 143 473 144 474
rect 142 473 143 474
rect 141 473 142 474
rect 140 473 141 474
rect 139 473 140 474
rect 138 473 139 474
rect 137 473 138 474
rect 136 473 137 474
rect 135 473 136 474
rect 134 473 135 474
rect 133 473 134 474
rect 132 473 133 474
rect 131 473 132 474
rect 130 473 131 474
rect 129 473 130 474
rect 128 473 129 474
rect 127 473 128 474
rect 126 473 127 474
rect 125 473 126 474
rect 124 473 125 474
rect 123 473 124 474
rect 122 473 123 474
rect 121 473 122 474
rect 120 473 121 474
rect 119 473 120 474
rect 118 473 119 474
rect 117 473 118 474
rect 116 473 117 474
rect 115 473 116 474
rect 114 473 115 474
rect 113 473 114 474
rect 112 473 113 474
rect 111 473 112 474
rect 110 473 111 474
rect 109 473 110 474
rect 108 473 109 474
rect 107 473 108 474
rect 106 473 107 474
rect 105 473 106 474
rect 104 473 105 474
rect 103 473 104 474
rect 102 473 103 474
rect 197 474 198 475
rect 196 474 197 475
rect 194 474 195 475
rect 193 474 194 475
rect 192 474 193 475
rect 191 474 192 475
rect 183 474 184 475
rect 182 474 183 475
rect 181 474 182 475
rect 180 474 181 475
rect 178 474 179 475
rect 177 474 178 475
rect 176 474 177 475
rect 175 474 176 475
rect 174 474 175 475
rect 173 474 174 475
rect 172 474 173 475
rect 171 474 172 475
rect 170 474 171 475
rect 169 474 170 475
rect 168 474 169 475
rect 167 474 168 475
rect 166 474 167 475
rect 165 474 166 475
rect 164 474 165 475
rect 163 474 164 475
rect 162 474 163 475
rect 149 474 150 475
rect 148 474 149 475
rect 147 474 148 475
rect 146 474 147 475
rect 145 474 146 475
rect 144 474 145 475
rect 143 474 144 475
rect 142 474 143 475
rect 141 474 142 475
rect 140 474 141 475
rect 139 474 140 475
rect 138 474 139 475
rect 137 474 138 475
rect 136 474 137 475
rect 135 474 136 475
rect 134 474 135 475
rect 133 474 134 475
rect 132 474 133 475
rect 131 474 132 475
rect 130 474 131 475
rect 129 474 130 475
rect 128 474 129 475
rect 127 474 128 475
rect 126 474 127 475
rect 125 474 126 475
rect 124 474 125 475
rect 123 474 124 475
rect 122 474 123 475
rect 121 474 122 475
rect 120 474 121 475
rect 119 474 120 475
rect 118 474 119 475
rect 117 474 118 475
rect 116 474 117 475
rect 115 474 116 475
rect 114 474 115 475
rect 113 474 114 475
rect 112 474 113 475
rect 111 474 112 475
rect 110 474 111 475
rect 109 474 110 475
rect 108 474 109 475
rect 107 474 108 475
rect 106 474 107 475
rect 105 474 106 475
rect 104 474 105 475
rect 103 474 104 475
rect 102 474 103 475
rect 196 475 197 476
rect 194 475 195 476
rect 193 475 194 476
rect 192 475 193 476
rect 191 475 192 476
rect 182 475 183 476
rect 181 475 182 476
rect 180 475 181 476
rect 177 475 178 476
rect 176 475 177 476
rect 175 475 176 476
rect 174 475 175 476
rect 173 475 174 476
rect 172 475 173 476
rect 171 475 172 476
rect 170 475 171 476
rect 169 475 170 476
rect 168 475 169 476
rect 167 475 168 476
rect 166 475 167 476
rect 165 475 166 476
rect 164 475 165 476
rect 163 475 164 476
rect 162 475 163 476
rect 149 475 150 476
rect 148 475 149 476
rect 147 475 148 476
rect 146 475 147 476
rect 145 475 146 476
rect 144 475 145 476
rect 143 475 144 476
rect 142 475 143 476
rect 141 475 142 476
rect 140 475 141 476
rect 139 475 140 476
rect 138 475 139 476
rect 137 475 138 476
rect 136 475 137 476
rect 135 475 136 476
rect 134 475 135 476
rect 133 475 134 476
rect 132 475 133 476
rect 131 475 132 476
rect 130 475 131 476
rect 129 475 130 476
rect 128 475 129 476
rect 127 475 128 476
rect 126 475 127 476
rect 125 475 126 476
rect 124 475 125 476
rect 123 475 124 476
rect 122 475 123 476
rect 121 475 122 476
rect 120 475 121 476
rect 119 475 120 476
rect 118 475 119 476
rect 117 475 118 476
rect 116 475 117 476
rect 115 475 116 476
rect 114 475 115 476
rect 113 475 114 476
rect 112 475 113 476
rect 111 475 112 476
rect 110 475 111 476
rect 109 475 110 476
rect 108 475 109 476
rect 107 475 108 476
rect 106 475 107 476
rect 105 475 106 476
rect 104 475 105 476
rect 103 475 104 476
rect 102 475 103 476
rect 194 476 195 477
rect 149 476 150 477
rect 148 476 149 477
rect 147 476 148 477
rect 146 476 147 477
rect 145 476 146 477
rect 144 476 145 477
rect 143 476 144 477
rect 142 476 143 477
rect 141 476 142 477
rect 140 476 141 477
rect 139 476 140 477
rect 138 476 139 477
rect 137 476 138 477
rect 136 476 137 477
rect 135 476 136 477
rect 134 476 135 477
rect 133 476 134 477
rect 132 476 133 477
rect 131 476 132 477
rect 130 476 131 477
rect 129 476 130 477
rect 128 476 129 477
rect 127 476 128 477
rect 126 476 127 477
rect 125 476 126 477
rect 124 476 125 477
rect 123 476 124 477
rect 122 476 123 477
rect 121 476 122 477
rect 120 476 121 477
rect 119 476 120 477
rect 118 476 119 477
rect 117 476 118 477
rect 116 476 117 477
rect 115 476 116 477
rect 114 476 115 477
rect 113 476 114 477
rect 112 476 113 477
rect 111 476 112 477
rect 110 476 111 477
rect 109 476 110 477
rect 108 476 109 477
rect 107 476 108 477
rect 106 476 107 477
rect 105 476 106 477
rect 104 476 105 477
rect 103 476 104 477
rect 102 476 103 477
<< metal3 >>
rect 182 9 183 10
rect 165 9 166 10
rect 182 10 183 11
rect 181 10 182 11
rect 166 10 167 11
rect 165 10 166 11
rect 182 11 183 12
rect 181 11 182 12
rect 180 11 181 12
rect 179 11 180 12
rect 178 11 179 12
rect 177 11 178 12
rect 176 11 177 12
rect 175 11 176 12
rect 174 11 175 12
rect 173 11 174 12
rect 172 11 173 12
rect 171 11 172 12
rect 170 11 171 12
rect 169 11 170 12
rect 168 11 169 12
rect 167 11 168 12
rect 166 11 167 12
rect 165 11 166 12
rect 182 12 183 13
rect 181 12 182 13
rect 180 12 181 13
rect 179 12 180 13
rect 178 12 179 13
rect 177 12 178 13
rect 176 12 177 13
rect 175 12 176 13
rect 174 12 175 13
rect 173 12 174 13
rect 172 12 173 13
rect 171 12 172 13
rect 170 12 171 13
rect 169 12 170 13
rect 168 12 169 13
rect 167 12 168 13
rect 166 12 167 13
rect 165 12 166 13
rect 182 13 183 14
rect 181 13 182 14
rect 180 13 181 14
rect 179 13 180 14
rect 178 13 179 14
rect 177 13 178 14
rect 176 13 177 14
rect 175 13 176 14
rect 174 13 175 14
rect 173 13 174 14
rect 172 13 173 14
rect 171 13 172 14
rect 170 13 171 14
rect 169 13 170 14
rect 168 13 169 14
rect 167 13 168 14
rect 166 13 167 14
rect 165 13 166 14
rect 182 14 183 15
rect 181 14 182 15
rect 180 14 181 15
rect 179 14 180 15
rect 178 14 179 15
rect 177 14 178 15
rect 176 14 177 15
rect 175 14 176 15
rect 174 14 175 15
rect 173 14 174 15
rect 172 14 173 15
rect 171 14 172 15
rect 170 14 171 15
rect 169 14 170 15
rect 168 14 169 15
rect 167 14 168 15
rect 166 14 167 15
rect 165 14 166 15
rect 182 15 183 16
rect 181 15 182 16
rect 174 15 175 16
rect 173 15 174 16
rect 166 15 167 16
rect 165 15 166 16
rect 182 16 183 17
rect 175 16 176 17
rect 174 16 175 17
rect 173 16 174 17
rect 172 16 173 17
rect 165 16 166 17
rect 177 17 178 18
rect 176 17 177 18
rect 175 17 176 18
rect 174 17 175 18
rect 173 17 174 18
rect 172 17 173 18
rect 171 17 172 18
rect 178 18 179 19
rect 177 18 178 19
rect 176 18 177 19
rect 175 18 176 19
rect 174 18 175 19
rect 173 18 174 19
rect 172 18 173 19
rect 171 18 172 19
rect 170 18 171 19
rect 180 19 181 20
rect 179 19 180 20
rect 178 19 179 20
rect 177 19 178 20
rect 176 19 177 20
rect 175 19 176 20
rect 174 19 175 20
rect 173 19 174 20
rect 170 19 171 20
rect 169 19 170 20
rect 165 19 166 20
rect 181 20 182 21
rect 180 20 181 21
rect 179 20 180 21
rect 178 20 179 21
rect 177 20 178 21
rect 176 20 177 21
rect 175 20 176 21
rect 169 20 170 21
rect 168 20 169 21
rect 167 20 168 21
rect 165 20 166 21
rect 182 21 183 22
rect 181 21 182 22
rect 180 21 181 22
rect 179 21 180 22
rect 178 21 179 22
rect 177 21 178 22
rect 176 21 177 22
rect 168 21 169 22
rect 167 21 168 22
rect 166 21 167 22
rect 165 21 166 22
rect 182 22 183 23
rect 181 22 182 23
rect 180 22 181 23
rect 179 22 180 23
rect 178 22 179 23
rect 167 22 168 23
rect 166 22 167 23
rect 165 22 166 23
rect 182 23 183 24
rect 181 23 182 24
rect 180 23 181 24
rect 179 23 180 24
rect 166 23 167 24
rect 165 23 166 24
rect 182 24 183 25
rect 181 24 182 25
rect 180 24 181 25
rect 166 24 167 25
rect 165 24 166 25
rect 182 25 183 26
rect 181 25 182 26
rect 165 25 166 26
rect 182 26 183 27
rect 165 26 166 27
rect 43 27 44 28
rect 42 27 43 28
rect 45 28 46 29
rect 44 28 45 29
rect 43 28 44 29
rect 42 28 43 29
rect 41 28 42 29
rect 40 28 41 29
rect 165 29 166 30
rect 45 29 46 30
rect 44 29 45 30
rect 43 29 44 30
rect 42 29 43 30
rect 41 29 42 30
rect 40 29 41 30
rect 39 29 40 30
rect 166 30 167 31
rect 165 30 166 31
rect 50 30 51 31
rect 49 30 50 31
rect 45 30 46 31
rect 44 30 45 31
rect 43 30 44 31
rect 42 30 43 31
rect 41 30 42 31
rect 40 30 41 31
rect 39 30 40 31
rect 38 30 39 31
rect 167 31 168 32
rect 166 31 167 32
rect 165 31 166 32
rect 52 31 53 32
rect 51 31 52 32
rect 50 31 51 32
rect 49 31 50 32
rect 48 31 49 32
rect 45 31 46 32
rect 44 31 45 32
rect 43 31 44 32
rect 42 31 43 32
rect 41 31 42 32
rect 40 31 41 32
rect 39 31 40 32
rect 38 31 39 32
rect 169 32 170 33
rect 168 32 169 33
rect 167 32 168 33
rect 166 32 167 33
rect 165 32 166 33
rect 54 32 55 33
rect 53 32 54 33
rect 52 32 53 33
rect 51 32 52 33
rect 50 32 51 33
rect 49 32 50 33
rect 48 32 49 33
rect 47 32 48 33
rect 44 32 45 33
rect 43 32 44 33
rect 42 32 43 33
rect 41 32 42 33
rect 40 32 41 33
rect 39 32 40 33
rect 38 32 39 33
rect 37 32 38 33
rect 182 33 183 34
rect 171 33 172 34
rect 170 33 171 34
rect 169 33 170 34
rect 168 33 169 34
rect 167 33 168 34
rect 166 33 167 34
rect 165 33 166 34
rect 55 33 56 34
rect 54 33 55 34
rect 53 33 54 34
rect 52 33 53 34
rect 51 33 52 34
rect 50 33 51 34
rect 49 33 50 34
rect 48 33 49 34
rect 47 33 48 34
rect 46 33 47 34
rect 44 33 45 34
rect 43 33 44 34
rect 42 33 43 34
rect 41 33 42 34
rect 40 33 41 34
rect 39 33 40 34
rect 38 33 39 34
rect 37 33 38 34
rect 182 34 183 35
rect 173 34 174 35
rect 172 34 173 35
rect 171 34 172 35
rect 170 34 171 35
rect 169 34 170 35
rect 168 34 169 35
rect 167 34 168 35
rect 166 34 167 35
rect 165 34 166 35
rect 56 34 57 35
rect 55 34 56 35
rect 54 34 55 35
rect 53 34 54 35
rect 52 34 53 35
rect 51 34 52 35
rect 50 34 51 35
rect 49 34 50 35
rect 48 34 49 35
rect 47 34 48 35
rect 46 34 47 35
rect 45 34 46 35
rect 43 34 44 35
rect 42 34 43 35
rect 41 34 42 35
rect 40 34 41 35
rect 39 34 40 35
rect 38 34 39 35
rect 37 34 38 35
rect 36 34 37 35
rect 182 35 183 36
rect 181 35 182 36
rect 180 35 181 36
rect 179 35 180 36
rect 178 35 179 36
rect 177 35 178 36
rect 176 35 177 36
rect 175 35 176 36
rect 174 35 175 36
rect 173 35 174 36
rect 172 35 173 36
rect 171 35 172 36
rect 170 35 171 36
rect 169 35 170 36
rect 168 35 169 36
rect 167 35 168 36
rect 166 35 167 36
rect 165 35 166 36
rect 56 35 57 36
rect 55 35 56 36
rect 54 35 55 36
rect 53 35 54 36
rect 52 35 53 36
rect 51 35 52 36
rect 50 35 51 36
rect 49 35 50 36
rect 48 35 49 36
rect 47 35 48 36
rect 46 35 47 36
rect 45 35 46 36
rect 44 35 45 36
rect 43 35 44 36
rect 42 35 43 36
rect 41 35 42 36
rect 40 35 41 36
rect 39 35 40 36
rect 38 35 39 36
rect 37 35 38 36
rect 36 35 37 36
rect 182 36 183 37
rect 181 36 182 37
rect 180 36 181 37
rect 179 36 180 37
rect 178 36 179 37
rect 177 36 178 37
rect 176 36 177 37
rect 175 36 176 37
rect 174 36 175 37
rect 173 36 174 37
rect 172 36 173 37
rect 171 36 172 37
rect 170 36 171 37
rect 169 36 170 37
rect 165 36 166 37
rect 63 36 64 37
rect 62 36 63 37
rect 61 36 62 37
rect 60 36 61 37
rect 57 36 58 37
rect 56 36 57 37
rect 55 36 56 37
rect 54 36 55 37
rect 53 36 54 37
rect 52 36 53 37
rect 51 36 52 37
rect 50 36 51 37
rect 49 36 50 37
rect 48 36 49 37
rect 47 36 48 37
rect 46 36 47 37
rect 45 36 46 37
rect 44 36 45 37
rect 43 36 44 37
rect 42 36 43 37
rect 41 36 42 37
rect 40 36 41 37
rect 39 36 40 37
rect 38 36 39 37
rect 37 36 38 37
rect 36 36 37 37
rect 35 36 36 37
rect 182 37 183 38
rect 181 37 182 38
rect 180 37 181 38
rect 179 37 180 38
rect 178 37 179 38
rect 177 37 178 38
rect 176 37 177 38
rect 175 37 176 38
rect 174 37 175 38
rect 173 37 174 38
rect 172 37 173 38
rect 171 37 172 38
rect 65 37 66 38
rect 64 37 65 38
rect 63 37 64 38
rect 62 37 63 38
rect 61 37 62 38
rect 60 37 61 38
rect 57 37 58 38
rect 56 37 57 38
rect 55 37 56 38
rect 54 37 55 38
rect 53 37 54 38
rect 52 37 53 38
rect 51 37 52 38
rect 50 37 51 38
rect 49 37 50 38
rect 48 37 49 38
rect 47 37 48 38
rect 46 37 47 38
rect 45 37 46 38
rect 44 37 45 38
rect 43 37 44 38
rect 42 37 43 38
rect 41 37 42 38
rect 40 37 41 38
rect 39 37 40 38
rect 38 37 39 38
rect 37 37 38 38
rect 36 37 37 38
rect 35 37 36 38
rect 182 38 183 39
rect 181 38 182 39
rect 180 38 181 39
rect 179 38 180 39
rect 178 38 179 39
rect 177 38 178 39
rect 176 38 177 39
rect 175 38 176 39
rect 174 38 175 39
rect 173 38 174 39
rect 67 38 68 39
rect 66 38 67 39
rect 65 38 66 39
rect 64 38 65 39
rect 63 38 64 39
rect 62 38 63 39
rect 61 38 62 39
rect 60 38 61 39
rect 57 38 58 39
rect 56 38 57 39
rect 55 38 56 39
rect 54 38 55 39
rect 53 38 54 39
rect 52 38 53 39
rect 51 38 52 39
rect 50 38 51 39
rect 49 38 50 39
rect 48 38 49 39
rect 47 38 48 39
rect 46 38 47 39
rect 45 38 46 39
rect 44 38 45 39
rect 43 38 44 39
rect 42 38 43 39
rect 41 38 42 39
rect 40 38 41 39
rect 39 38 40 39
rect 38 38 39 39
rect 37 38 38 39
rect 36 38 37 39
rect 35 38 36 39
rect 34 38 35 39
rect 182 39 183 40
rect 181 39 182 40
rect 180 39 181 40
rect 179 39 180 40
rect 178 39 179 40
rect 177 39 178 40
rect 176 39 177 40
rect 175 39 176 40
rect 174 39 175 40
rect 173 39 174 40
rect 172 39 173 40
rect 171 39 172 40
rect 69 39 70 40
rect 68 39 69 40
rect 67 39 68 40
rect 66 39 67 40
rect 65 39 66 40
rect 64 39 65 40
rect 63 39 64 40
rect 62 39 63 40
rect 61 39 62 40
rect 60 39 61 40
rect 57 39 58 40
rect 56 39 57 40
rect 55 39 56 40
rect 54 39 55 40
rect 53 39 54 40
rect 52 39 53 40
rect 51 39 52 40
rect 50 39 51 40
rect 49 39 50 40
rect 48 39 49 40
rect 47 39 48 40
rect 46 39 47 40
rect 45 39 46 40
rect 44 39 45 40
rect 43 39 44 40
rect 42 39 43 40
rect 41 39 42 40
rect 40 39 41 40
rect 39 39 40 40
rect 38 39 39 40
rect 37 39 38 40
rect 36 39 37 40
rect 35 39 36 40
rect 34 39 35 40
rect 182 40 183 41
rect 172 40 173 41
rect 171 40 172 41
rect 170 40 171 41
rect 169 40 170 41
rect 165 40 166 41
rect 71 40 72 41
rect 70 40 71 41
rect 69 40 70 41
rect 68 40 69 41
rect 67 40 68 41
rect 66 40 67 41
rect 65 40 66 41
rect 64 40 65 41
rect 63 40 64 41
rect 62 40 63 41
rect 61 40 62 41
rect 60 40 61 41
rect 57 40 58 41
rect 56 40 57 41
rect 55 40 56 41
rect 54 40 55 41
rect 53 40 54 41
rect 52 40 53 41
rect 51 40 52 41
rect 50 40 51 41
rect 49 40 50 41
rect 48 40 49 41
rect 47 40 48 41
rect 46 40 47 41
rect 45 40 46 41
rect 44 40 45 41
rect 43 40 44 41
rect 42 40 43 41
rect 41 40 42 41
rect 40 40 41 41
rect 39 40 40 41
rect 38 40 39 41
rect 37 40 38 41
rect 36 40 37 41
rect 35 40 36 41
rect 34 40 35 41
rect 33 40 34 41
rect 197 41 198 42
rect 196 41 197 42
rect 195 41 196 42
rect 194 41 195 42
rect 193 41 194 42
rect 192 41 193 42
rect 191 41 192 42
rect 182 41 183 42
rect 170 41 171 42
rect 169 41 170 42
rect 168 41 169 42
rect 167 41 168 42
rect 166 41 167 42
rect 165 41 166 42
rect 99 41 100 42
rect 98 41 99 42
rect 97 41 98 42
rect 96 41 97 42
rect 95 41 96 42
rect 94 41 95 42
rect 93 41 94 42
rect 92 41 93 42
rect 91 41 92 42
rect 90 41 91 42
rect 89 41 90 42
rect 72 41 73 42
rect 71 41 72 42
rect 70 41 71 42
rect 69 41 70 42
rect 68 41 69 42
rect 67 41 68 42
rect 66 41 67 42
rect 65 41 66 42
rect 64 41 65 42
rect 63 41 64 42
rect 62 41 63 42
rect 61 41 62 42
rect 60 41 61 42
rect 59 41 60 42
rect 56 41 57 42
rect 55 41 56 42
rect 54 41 55 42
rect 53 41 54 42
rect 52 41 53 42
rect 51 41 52 42
rect 50 41 51 42
rect 49 41 50 42
rect 48 41 49 42
rect 47 41 48 42
rect 46 41 47 42
rect 45 41 46 42
rect 44 41 45 42
rect 43 41 44 42
rect 42 41 43 42
rect 41 41 42 42
rect 40 41 41 42
rect 39 41 40 42
rect 38 41 39 42
rect 37 41 38 42
rect 36 41 37 42
rect 35 41 36 42
rect 34 41 35 42
rect 33 41 34 42
rect 32 41 33 42
rect 198 42 199 43
rect 197 42 198 43
rect 196 42 197 43
rect 195 42 196 43
rect 194 42 195 43
rect 193 42 194 43
rect 192 42 193 43
rect 191 42 192 43
rect 168 42 169 43
rect 167 42 168 43
rect 166 42 167 43
rect 165 42 166 43
rect 103 42 104 43
rect 102 42 103 43
rect 101 42 102 43
rect 100 42 101 43
rect 99 42 100 43
rect 98 42 99 43
rect 97 42 98 43
rect 96 42 97 43
rect 95 42 96 43
rect 94 42 95 43
rect 93 42 94 43
rect 92 42 93 43
rect 91 42 92 43
rect 90 42 91 43
rect 89 42 90 43
rect 88 42 89 43
rect 87 42 88 43
rect 86 42 87 43
rect 72 42 73 43
rect 71 42 72 43
rect 70 42 71 43
rect 69 42 70 43
rect 68 42 69 43
rect 67 42 68 43
rect 66 42 67 43
rect 65 42 66 43
rect 64 42 65 43
rect 63 42 64 43
rect 62 42 63 43
rect 61 42 62 43
rect 60 42 61 43
rect 59 42 60 43
rect 56 42 57 43
rect 55 42 56 43
rect 54 42 55 43
rect 53 42 54 43
rect 52 42 53 43
rect 51 42 52 43
rect 50 42 51 43
rect 49 42 50 43
rect 48 42 49 43
rect 47 42 48 43
rect 46 42 47 43
rect 45 42 46 43
rect 44 42 45 43
rect 43 42 44 43
rect 42 42 43 43
rect 41 42 42 43
rect 40 42 41 43
rect 39 42 40 43
rect 38 42 39 43
rect 37 42 38 43
rect 36 42 37 43
rect 35 42 36 43
rect 34 42 35 43
rect 33 42 34 43
rect 32 42 33 43
rect 199 43 200 44
rect 198 43 199 44
rect 197 43 198 44
rect 191 43 192 44
rect 167 43 168 44
rect 166 43 167 44
rect 165 43 166 44
rect 105 43 106 44
rect 104 43 105 44
rect 103 43 104 44
rect 102 43 103 44
rect 101 43 102 44
rect 100 43 101 44
rect 99 43 100 44
rect 98 43 99 44
rect 97 43 98 44
rect 96 43 97 44
rect 95 43 96 44
rect 94 43 95 44
rect 93 43 94 44
rect 92 43 93 44
rect 91 43 92 44
rect 90 43 91 44
rect 89 43 90 44
rect 88 43 89 44
rect 87 43 88 44
rect 86 43 87 44
rect 85 43 86 44
rect 84 43 85 44
rect 72 43 73 44
rect 71 43 72 44
rect 70 43 71 44
rect 69 43 70 44
rect 68 43 69 44
rect 67 43 68 44
rect 66 43 67 44
rect 65 43 66 44
rect 64 43 65 44
rect 63 43 64 44
rect 62 43 63 44
rect 61 43 62 44
rect 60 43 61 44
rect 59 43 60 44
rect 56 43 57 44
rect 55 43 56 44
rect 54 43 55 44
rect 53 43 54 44
rect 52 43 53 44
rect 51 43 52 44
rect 50 43 51 44
rect 49 43 50 44
rect 48 43 49 44
rect 47 43 48 44
rect 46 43 47 44
rect 45 43 46 44
rect 44 43 45 44
rect 43 43 44 44
rect 42 43 43 44
rect 41 43 42 44
rect 40 43 41 44
rect 39 43 40 44
rect 38 43 39 44
rect 37 43 38 44
rect 36 43 37 44
rect 35 43 36 44
rect 34 43 35 44
rect 33 43 34 44
rect 32 43 33 44
rect 31 43 32 44
rect 199 44 200 45
rect 198 44 199 45
rect 166 44 167 45
rect 165 44 166 45
rect 107 44 108 45
rect 106 44 107 45
rect 105 44 106 45
rect 104 44 105 45
rect 103 44 104 45
rect 102 44 103 45
rect 101 44 102 45
rect 100 44 101 45
rect 99 44 100 45
rect 98 44 99 45
rect 97 44 98 45
rect 96 44 97 45
rect 95 44 96 45
rect 94 44 95 45
rect 93 44 94 45
rect 92 44 93 45
rect 91 44 92 45
rect 90 44 91 45
rect 89 44 90 45
rect 88 44 89 45
rect 87 44 88 45
rect 86 44 87 45
rect 85 44 86 45
rect 84 44 85 45
rect 83 44 84 45
rect 82 44 83 45
rect 71 44 72 45
rect 70 44 71 45
rect 69 44 70 45
rect 68 44 69 45
rect 67 44 68 45
rect 66 44 67 45
rect 65 44 66 45
rect 64 44 65 45
rect 63 44 64 45
rect 62 44 63 45
rect 61 44 62 45
rect 60 44 61 45
rect 59 44 60 45
rect 56 44 57 45
rect 55 44 56 45
rect 54 44 55 45
rect 53 44 54 45
rect 52 44 53 45
rect 51 44 52 45
rect 50 44 51 45
rect 49 44 50 45
rect 48 44 49 45
rect 47 44 48 45
rect 46 44 47 45
rect 45 44 46 45
rect 44 44 45 45
rect 43 44 44 45
rect 42 44 43 45
rect 41 44 42 45
rect 40 44 41 45
rect 39 44 40 45
rect 38 44 39 45
rect 37 44 38 45
rect 36 44 37 45
rect 35 44 36 45
rect 34 44 35 45
rect 33 44 34 45
rect 32 44 33 45
rect 31 44 32 45
rect 30 44 31 45
rect 199 45 200 46
rect 165 45 166 46
rect 109 45 110 46
rect 108 45 109 46
rect 107 45 108 46
rect 106 45 107 46
rect 105 45 106 46
rect 104 45 105 46
rect 103 45 104 46
rect 102 45 103 46
rect 101 45 102 46
rect 100 45 101 46
rect 99 45 100 46
rect 98 45 99 46
rect 97 45 98 46
rect 96 45 97 46
rect 95 45 96 46
rect 94 45 95 46
rect 93 45 94 46
rect 92 45 93 46
rect 91 45 92 46
rect 90 45 91 46
rect 89 45 90 46
rect 88 45 89 46
rect 87 45 88 46
rect 86 45 87 46
rect 85 45 86 46
rect 84 45 85 46
rect 83 45 84 46
rect 82 45 83 46
rect 81 45 82 46
rect 71 45 72 46
rect 70 45 71 46
rect 69 45 70 46
rect 68 45 69 46
rect 67 45 68 46
rect 66 45 67 46
rect 65 45 66 46
rect 64 45 65 46
rect 63 45 64 46
rect 62 45 63 46
rect 61 45 62 46
rect 60 45 61 46
rect 59 45 60 46
rect 56 45 57 46
rect 55 45 56 46
rect 54 45 55 46
rect 53 45 54 46
rect 52 45 53 46
rect 51 45 52 46
rect 50 45 51 46
rect 49 45 50 46
rect 48 45 49 46
rect 47 45 48 46
rect 46 45 47 46
rect 45 45 46 46
rect 44 45 45 46
rect 43 45 44 46
rect 42 45 43 46
rect 41 45 42 46
rect 40 45 41 46
rect 39 45 40 46
rect 38 45 39 46
rect 37 45 38 46
rect 36 45 37 46
rect 35 45 36 46
rect 34 45 35 46
rect 33 45 34 46
rect 32 45 33 46
rect 31 45 32 46
rect 30 45 31 46
rect 199 46 200 47
rect 198 46 199 47
rect 111 46 112 47
rect 110 46 111 47
rect 109 46 110 47
rect 108 46 109 47
rect 107 46 108 47
rect 106 46 107 47
rect 105 46 106 47
rect 104 46 105 47
rect 103 46 104 47
rect 102 46 103 47
rect 101 46 102 47
rect 100 46 101 47
rect 99 46 100 47
rect 98 46 99 47
rect 97 46 98 47
rect 96 46 97 47
rect 95 46 96 47
rect 94 46 95 47
rect 93 46 94 47
rect 92 46 93 47
rect 91 46 92 47
rect 90 46 91 47
rect 89 46 90 47
rect 88 46 89 47
rect 87 46 88 47
rect 86 46 87 47
rect 85 46 86 47
rect 84 46 85 47
rect 83 46 84 47
rect 82 46 83 47
rect 81 46 82 47
rect 80 46 81 47
rect 71 46 72 47
rect 70 46 71 47
rect 69 46 70 47
rect 68 46 69 47
rect 67 46 68 47
rect 66 46 67 47
rect 65 46 66 47
rect 64 46 65 47
rect 63 46 64 47
rect 62 46 63 47
rect 61 46 62 47
rect 60 46 61 47
rect 59 46 60 47
rect 55 46 56 47
rect 54 46 55 47
rect 53 46 54 47
rect 52 46 53 47
rect 51 46 52 47
rect 50 46 51 47
rect 49 46 50 47
rect 48 46 49 47
rect 47 46 48 47
rect 46 46 47 47
rect 45 46 46 47
rect 44 46 45 47
rect 43 46 44 47
rect 42 46 43 47
rect 41 46 42 47
rect 40 46 41 47
rect 39 46 40 47
rect 38 46 39 47
rect 37 46 38 47
rect 36 46 37 47
rect 35 46 36 47
rect 34 46 35 47
rect 33 46 34 47
rect 32 46 33 47
rect 31 46 32 47
rect 30 46 31 47
rect 29 46 30 47
rect 198 47 199 48
rect 197 47 198 48
rect 196 47 197 48
rect 195 47 196 48
rect 194 47 195 48
rect 193 47 194 48
rect 192 47 193 48
rect 191 47 192 48
rect 112 47 113 48
rect 111 47 112 48
rect 110 47 111 48
rect 109 47 110 48
rect 108 47 109 48
rect 107 47 108 48
rect 106 47 107 48
rect 105 47 106 48
rect 104 47 105 48
rect 103 47 104 48
rect 102 47 103 48
rect 101 47 102 48
rect 100 47 101 48
rect 99 47 100 48
rect 98 47 99 48
rect 97 47 98 48
rect 96 47 97 48
rect 95 47 96 48
rect 94 47 95 48
rect 93 47 94 48
rect 92 47 93 48
rect 91 47 92 48
rect 90 47 91 48
rect 89 47 90 48
rect 88 47 89 48
rect 87 47 88 48
rect 86 47 87 48
rect 85 47 86 48
rect 84 47 85 48
rect 83 47 84 48
rect 82 47 83 48
rect 81 47 82 48
rect 80 47 81 48
rect 79 47 80 48
rect 70 47 71 48
rect 69 47 70 48
rect 68 47 69 48
rect 67 47 68 48
rect 66 47 67 48
rect 65 47 66 48
rect 64 47 65 48
rect 63 47 64 48
rect 62 47 63 48
rect 61 47 62 48
rect 60 47 61 48
rect 59 47 60 48
rect 58 47 59 48
rect 55 47 56 48
rect 54 47 55 48
rect 53 47 54 48
rect 52 47 53 48
rect 51 47 52 48
rect 50 47 51 48
rect 49 47 50 48
rect 48 47 49 48
rect 47 47 48 48
rect 46 47 47 48
rect 45 47 46 48
rect 44 47 45 48
rect 43 47 44 48
rect 42 47 43 48
rect 41 47 42 48
rect 40 47 41 48
rect 39 47 40 48
rect 38 47 39 48
rect 37 47 38 48
rect 35 47 36 48
rect 34 47 35 48
rect 33 47 34 48
rect 32 47 33 48
rect 31 47 32 48
rect 30 47 31 48
rect 29 47 30 48
rect 28 47 29 48
rect 192 48 193 49
rect 191 48 192 49
rect 165 48 166 49
rect 113 48 114 49
rect 112 48 113 49
rect 111 48 112 49
rect 110 48 111 49
rect 109 48 110 49
rect 108 48 109 49
rect 107 48 108 49
rect 106 48 107 49
rect 105 48 106 49
rect 104 48 105 49
rect 103 48 104 49
rect 102 48 103 49
rect 101 48 102 49
rect 100 48 101 49
rect 99 48 100 49
rect 98 48 99 49
rect 97 48 98 49
rect 96 48 97 49
rect 95 48 96 49
rect 94 48 95 49
rect 93 48 94 49
rect 92 48 93 49
rect 91 48 92 49
rect 90 48 91 49
rect 89 48 90 49
rect 88 48 89 49
rect 87 48 88 49
rect 86 48 87 49
rect 85 48 86 49
rect 84 48 85 49
rect 83 48 84 49
rect 82 48 83 49
rect 81 48 82 49
rect 80 48 81 49
rect 79 48 80 49
rect 78 48 79 49
rect 70 48 71 49
rect 69 48 70 49
rect 68 48 69 49
rect 67 48 68 49
rect 66 48 67 49
rect 65 48 66 49
rect 64 48 65 49
rect 63 48 64 49
rect 62 48 63 49
rect 61 48 62 49
rect 60 48 61 49
rect 59 48 60 49
rect 58 48 59 49
rect 54 48 55 49
rect 53 48 54 49
rect 52 48 53 49
rect 51 48 52 49
rect 50 48 51 49
rect 49 48 50 49
rect 48 48 49 49
rect 47 48 48 49
rect 46 48 47 49
rect 45 48 46 49
rect 44 48 45 49
rect 43 48 44 49
rect 42 48 43 49
rect 41 48 42 49
rect 40 48 41 49
rect 39 48 40 49
rect 38 48 39 49
rect 37 48 38 49
rect 34 48 35 49
rect 33 48 34 49
rect 32 48 33 49
rect 31 48 32 49
rect 30 48 31 49
rect 29 48 30 49
rect 28 48 29 49
rect 27 48 28 49
rect 165 49 166 50
rect 114 49 115 50
rect 113 49 114 50
rect 112 49 113 50
rect 111 49 112 50
rect 110 49 111 50
rect 109 49 110 50
rect 108 49 109 50
rect 107 49 108 50
rect 106 49 107 50
rect 105 49 106 50
rect 104 49 105 50
rect 103 49 104 50
rect 102 49 103 50
rect 101 49 102 50
rect 100 49 101 50
rect 99 49 100 50
rect 98 49 99 50
rect 97 49 98 50
rect 96 49 97 50
rect 95 49 96 50
rect 94 49 95 50
rect 93 49 94 50
rect 92 49 93 50
rect 91 49 92 50
rect 90 49 91 50
rect 89 49 90 50
rect 88 49 89 50
rect 87 49 88 50
rect 86 49 87 50
rect 85 49 86 50
rect 84 49 85 50
rect 83 49 84 50
rect 82 49 83 50
rect 81 49 82 50
rect 80 49 81 50
rect 79 49 80 50
rect 78 49 79 50
rect 70 49 71 50
rect 69 49 70 50
rect 68 49 69 50
rect 67 49 68 50
rect 66 49 67 50
rect 65 49 66 50
rect 64 49 65 50
rect 63 49 64 50
rect 62 49 63 50
rect 61 49 62 50
rect 60 49 61 50
rect 59 49 60 50
rect 58 49 59 50
rect 53 49 54 50
rect 52 49 53 50
rect 51 49 52 50
rect 50 49 51 50
rect 49 49 50 50
rect 48 49 49 50
rect 47 49 48 50
rect 46 49 47 50
rect 45 49 46 50
rect 44 49 45 50
rect 43 49 44 50
rect 42 49 43 50
rect 41 49 42 50
rect 40 49 41 50
rect 39 49 40 50
rect 38 49 39 50
rect 37 49 38 50
rect 34 49 35 50
rect 33 49 34 50
rect 32 49 33 50
rect 31 49 32 50
rect 30 49 31 50
rect 29 49 30 50
rect 28 49 29 50
rect 27 49 28 50
rect 26 49 27 50
rect 175 50 176 51
rect 174 50 175 51
rect 173 50 174 51
rect 172 50 173 51
rect 171 50 172 51
rect 170 50 171 51
rect 169 50 170 51
rect 168 50 169 51
rect 167 50 168 51
rect 166 50 167 51
rect 165 50 166 51
rect 115 50 116 51
rect 114 50 115 51
rect 113 50 114 51
rect 112 50 113 51
rect 111 50 112 51
rect 110 50 111 51
rect 109 50 110 51
rect 108 50 109 51
rect 107 50 108 51
rect 106 50 107 51
rect 105 50 106 51
rect 104 50 105 51
rect 103 50 104 51
rect 102 50 103 51
rect 101 50 102 51
rect 100 50 101 51
rect 99 50 100 51
rect 98 50 99 51
rect 97 50 98 51
rect 96 50 97 51
rect 95 50 96 51
rect 94 50 95 51
rect 93 50 94 51
rect 92 50 93 51
rect 91 50 92 51
rect 90 50 91 51
rect 89 50 90 51
rect 88 50 89 51
rect 87 50 88 51
rect 86 50 87 51
rect 85 50 86 51
rect 84 50 85 51
rect 83 50 84 51
rect 82 50 83 51
rect 81 50 82 51
rect 80 50 81 51
rect 79 50 80 51
rect 78 50 79 51
rect 77 50 78 51
rect 69 50 70 51
rect 68 50 69 51
rect 67 50 68 51
rect 66 50 67 51
rect 65 50 66 51
rect 64 50 65 51
rect 63 50 64 51
rect 62 50 63 51
rect 61 50 62 51
rect 60 50 61 51
rect 59 50 60 51
rect 58 50 59 51
rect 53 50 54 51
rect 52 50 53 51
rect 51 50 52 51
rect 50 50 51 51
rect 49 50 50 51
rect 48 50 49 51
rect 47 50 48 51
rect 46 50 47 51
rect 45 50 46 51
rect 44 50 45 51
rect 43 50 44 51
rect 42 50 43 51
rect 41 50 42 51
rect 40 50 41 51
rect 39 50 40 51
rect 38 50 39 51
rect 33 50 34 51
rect 32 50 33 51
rect 31 50 32 51
rect 30 50 31 51
rect 29 50 30 51
rect 28 50 29 51
rect 27 50 28 51
rect 26 50 27 51
rect 25 50 26 51
rect 24 50 25 51
rect 179 51 180 52
rect 178 51 179 52
rect 177 51 178 52
rect 176 51 177 52
rect 175 51 176 52
rect 174 51 175 52
rect 173 51 174 52
rect 172 51 173 52
rect 171 51 172 52
rect 170 51 171 52
rect 169 51 170 52
rect 168 51 169 52
rect 167 51 168 52
rect 166 51 167 52
rect 165 51 166 52
rect 116 51 117 52
rect 115 51 116 52
rect 114 51 115 52
rect 113 51 114 52
rect 112 51 113 52
rect 111 51 112 52
rect 110 51 111 52
rect 109 51 110 52
rect 108 51 109 52
rect 107 51 108 52
rect 106 51 107 52
rect 105 51 106 52
rect 104 51 105 52
rect 103 51 104 52
rect 102 51 103 52
rect 101 51 102 52
rect 100 51 101 52
rect 99 51 100 52
rect 98 51 99 52
rect 97 51 98 52
rect 96 51 97 52
rect 95 51 96 52
rect 94 51 95 52
rect 93 51 94 52
rect 92 51 93 52
rect 91 51 92 52
rect 90 51 91 52
rect 89 51 90 52
rect 88 51 89 52
rect 87 51 88 52
rect 86 51 87 52
rect 85 51 86 52
rect 84 51 85 52
rect 83 51 84 52
rect 82 51 83 52
rect 81 51 82 52
rect 80 51 81 52
rect 79 51 80 52
rect 78 51 79 52
rect 77 51 78 52
rect 69 51 70 52
rect 68 51 69 52
rect 67 51 68 52
rect 66 51 67 52
rect 65 51 66 52
rect 64 51 65 52
rect 63 51 64 52
rect 62 51 63 52
rect 61 51 62 52
rect 60 51 61 52
rect 59 51 60 52
rect 58 51 59 52
rect 57 51 58 52
rect 54 51 55 52
rect 53 51 54 52
rect 52 51 53 52
rect 51 51 52 52
rect 50 51 51 52
rect 49 51 50 52
rect 48 51 49 52
rect 47 51 48 52
rect 46 51 47 52
rect 45 51 46 52
rect 44 51 45 52
rect 43 51 44 52
rect 42 51 43 52
rect 41 51 42 52
rect 40 51 41 52
rect 33 51 34 52
rect 32 51 33 52
rect 31 51 32 52
rect 30 51 31 52
rect 29 51 30 52
rect 28 51 29 52
rect 27 51 28 52
rect 26 51 27 52
rect 25 51 26 52
rect 24 51 25 52
rect 23 51 24 52
rect 181 52 182 53
rect 180 52 181 53
rect 179 52 180 53
rect 178 52 179 53
rect 177 52 178 53
rect 176 52 177 53
rect 175 52 176 53
rect 174 52 175 53
rect 173 52 174 53
rect 172 52 173 53
rect 171 52 172 53
rect 170 52 171 53
rect 169 52 170 53
rect 168 52 169 53
rect 167 52 168 53
rect 166 52 167 53
rect 165 52 166 53
rect 117 52 118 53
rect 116 52 117 53
rect 115 52 116 53
rect 114 52 115 53
rect 113 52 114 53
rect 112 52 113 53
rect 111 52 112 53
rect 110 52 111 53
rect 109 52 110 53
rect 108 52 109 53
rect 107 52 108 53
rect 106 52 107 53
rect 105 52 106 53
rect 104 52 105 53
rect 103 52 104 53
rect 102 52 103 53
rect 101 52 102 53
rect 100 52 101 53
rect 99 52 100 53
rect 98 52 99 53
rect 97 52 98 53
rect 96 52 97 53
rect 95 52 96 53
rect 94 52 95 53
rect 93 52 94 53
rect 92 52 93 53
rect 91 52 92 53
rect 90 52 91 53
rect 89 52 90 53
rect 88 52 89 53
rect 87 52 88 53
rect 86 52 87 53
rect 85 52 86 53
rect 84 52 85 53
rect 83 52 84 53
rect 82 52 83 53
rect 81 52 82 53
rect 80 52 81 53
rect 79 52 80 53
rect 78 52 79 53
rect 77 52 78 53
rect 76 52 77 53
rect 69 52 70 53
rect 68 52 69 53
rect 67 52 68 53
rect 66 52 67 53
rect 65 52 66 53
rect 64 52 65 53
rect 63 52 64 53
rect 62 52 63 53
rect 61 52 62 53
rect 60 52 61 53
rect 59 52 60 53
rect 58 52 59 53
rect 57 52 58 53
rect 56 52 57 53
rect 55 52 56 53
rect 54 52 55 53
rect 53 52 54 53
rect 52 52 53 53
rect 51 52 52 53
rect 50 52 51 53
rect 49 52 50 53
rect 48 52 49 53
rect 47 52 48 53
rect 46 52 47 53
rect 45 52 46 53
rect 44 52 45 53
rect 43 52 44 53
rect 42 52 43 53
rect 41 52 42 53
rect 40 52 41 53
rect 39 52 40 53
rect 32 52 33 53
rect 31 52 32 53
rect 30 52 31 53
rect 29 52 30 53
rect 28 52 29 53
rect 27 52 28 53
rect 26 52 27 53
rect 25 52 26 53
rect 24 52 25 53
rect 23 52 24 53
rect 22 52 23 53
rect 21 52 22 53
rect 199 53 200 54
rect 198 53 199 54
rect 197 53 198 54
rect 196 53 197 54
rect 195 53 196 54
rect 194 53 195 54
rect 193 53 194 54
rect 192 53 193 54
rect 191 53 192 54
rect 182 53 183 54
rect 181 53 182 54
rect 180 53 181 54
rect 179 53 180 54
rect 178 53 179 54
rect 177 53 178 54
rect 176 53 177 54
rect 175 53 176 54
rect 174 53 175 54
rect 173 53 174 54
rect 172 53 173 54
rect 171 53 172 54
rect 170 53 171 54
rect 169 53 170 54
rect 168 53 169 54
rect 167 53 168 54
rect 166 53 167 54
rect 165 53 166 54
rect 112 53 113 54
rect 111 53 112 54
rect 110 53 111 54
rect 109 53 110 54
rect 108 53 109 54
rect 107 53 108 54
rect 106 53 107 54
rect 105 53 106 54
rect 104 53 105 54
rect 103 53 104 54
rect 102 53 103 54
rect 101 53 102 54
rect 100 53 101 54
rect 99 53 100 54
rect 98 53 99 54
rect 97 53 98 54
rect 96 53 97 54
rect 95 53 96 54
rect 94 53 95 54
rect 93 53 94 54
rect 92 53 93 54
rect 91 53 92 54
rect 90 53 91 54
rect 89 53 90 54
rect 88 53 89 54
rect 87 53 88 54
rect 86 53 87 54
rect 85 53 86 54
rect 84 53 85 54
rect 83 53 84 54
rect 82 53 83 54
rect 81 53 82 54
rect 80 53 81 54
rect 79 53 80 54
rect 78 53 79 54
rect 77 53 78 54
rect 76 53 77 54
rect 68 53 69 54
rect 67 53 68 54
rect 66 53 67 54
rect 65 53 66 54
rect 64 53 65 54
rect 63 53 64 54
rect 62 53 63 54
rect 61 53 62 54
rect 60 53 61 54
rect 59 53 60 54
rect 58 53 59 54
rect 57 53 58 54
rect 56 53 57 54
rect 55 53 56 54
rect 54 53 55 54
rect 53 53 54 54
rect 52 53 53 54
rect 51 53 52 54
rect 50 53 51 54
rect 49 53 50 54
rect 48 53 49 54
rect 47 53 48 54
rect 46 53 47 54
rect 45 53 46 54
rect 44 53 45 54
rect 43 53 44 54
rect 42 53 43 54
rect 41 53 42 54
rect 40 53 41 54
rect 39 53 40 54
rect 38 53 39 54
rect 37 53 38 54
rect 32 53 33 54
rect 31 53 32 54
rect 30 53 31 54
rect 29 53 30 54
rect 28 53 29 54
rect 27 53 28 54
rect 26 53 27 54
rect 25 53 26 54
rect 24 53 25 54
rect 23 53 24 54
rect 22 53 23 54
rect 21 53 22 54
rect 20 53 21 54
rect 199 54 200 55
rect 198 54 199 55
rect 193 54 194 55
rect 192 54 193 55
rect 191 54 192 55
rect 182 54 183 55
rect 181 54 182 55
rect 180 54 181 55
rect 179 54 180 55
rect 178 54 179 55
rect 177 54 178 55
rect 176 54 177 55
rect 175 54 176 55
rect 174 54 175 55
rect 173 54 174 55
rect 172 54 173 55
rect 171 54 172 55
rect 170 54 171 55
rect 169 54 170 55
rect 168 54 169 55
rect 167 54 168 55
rect 166 54 167 55
rect 165 54 166 55
rect 106 54 107 55
rect 105 54 106 55
rect 104 54 105 55
rect 103 54 104 55
rect 102 54 103 55
rect 101 54 102 55
rect 100 54 101 55
rect 99 54 100 55
rect 98 54 99 55
rect 97 54 98 55
rect 96 54 97 55
rect 95 54 96 55
rect 94 54 95 55
rect 93 54 94 55
rect 92 54 93 55
rect 91 54 92 55
rect 90 54 91 55
rect 89 54 90 55
rect 88 54 89 55
rect 87 54 88 55
rect 86 54 87 55
rect 85 54 86 55
rect 84 54 85 55
rect 83 54 84 55
rect 82 54 83 55
rect 81 54 82 55
rect 80 54 81 55
rect 79 54 80 55
rect 78 54 79 55
rect 77 54 78 55
rect 76 54 77 55
rect 75 54 76 55
rect 68 54 69 55
rect 67 54 68 55
rect 66 54 67 55
rect 65 54 66 55
rect 64 54 65 55
rect 63 54 64 55
rect 62 54 63 55
rect 61 54 62 55
rect 60 54 61 55
rect 59 54 60 55
rect 58 54 59 55
rect 57 54 58 55
rect 56 54 57 55
rect 55 54 56 55
rect 54 54 55 55
rect 53 54 54 55
rect 52 54 53 55
rect 51 54 52 55
rect 50 54 51 55
rect 49 54 50 55
rect 48 54 49 55
rect 47 54 48 55
rect 46 54 47 55
rect 45 54 46 55
rect 44 54 45 55
rect 43 54 44 55
rect 42 54 43 55
rect 41 54 42 55
rect 40 54 41 55
rect 39 54 40 55
rect 38 54 39 55
rect 37 54 38 55
rect 36 54 37 55
rect 32 54 33 55
rect 31 54 32 55
rect 30 54 31 55
rect 29 54 30 55
rect 28 54 29 55
rect 27 54 28 55
rect 26 54 27 55
rect 25 54 26 55
rect 24 54 25 55
rect 23 54 24 55
rect 22 54 23 55
rect 21 54 22 55
rect 20 54 21 55
rect 194 55 195 56
rect 193 55 194 56
rect 192 55 193 56
rect 191 55 192 56
rect 182 55 183 56
rect 181 55 182 56
rect 180 55 181 56
rect 179 55 180 56
rect 166 55 167 56
rect 165 55 166 56
rect 104 55 105 56
rect 103 55 104 56
rect 102 55 103 56
rect 101 55 102 56
rect 100 55 101 56
rect 99 55 100 56
rect 98 55 99 56
rect 97 55 98 56
rect 96 55 97 56
rect 95 55 96 56
rect 94 55 95 56
rect 93 55 94 56
rect 92 55 93 56
rect 91 55 92 56
rect 90 55 91 56
rect 89 55 90 56
rect 88 55 89 56
rect 87 55 88 56
rect 86 55 87 56
rect 85 55 86 56
rect 84 55 85 56
rect 83 55 84 56
rect 82 55 83 56
rect 81 55 82 56
rect 80 55 81 56
rect 79 55 80 56
rect 78 55 79 56
rect 77 55 78 56
rect 76 55 77 56
rect 75 55 76 56
rect 68 55 69 56
rect 67 55 68 56
rect 66 55 67 56
rect 65 55 66 56
rect 64 55 65 56
rect 63 55 64 56
rect 62 55 63 56
rect 61 55 62 56
rect 60 55 61 56
rect 59 55 60 56
rect 58 55 59 56
rect 57 55 58 56
rect 56 55 57 56
rect 55 55 56 56
rect 54 55 55 56
rect 53 55 54 56
rect 52 55 53 56
rect 51 55 52 56
rect 50 55 51 56
rect 49 55 50 56
rect 48 55 49 56
rect 47 55 48 56
rect 46 55 47 56
rect 45 55 46 56
rect 44 55 45 56
rect 43 55 44 56
rect 42 55 43 56
rect 41 55 42 56
rect 40 55 41 56
rect 39 55 40 56
rect 38 55 39 56
rect 37 55 38 56
rect 36 55 37 56
rect 35 55 36 56
rect 31 55 32 56
rect 30 55 31 56
rect 29 55 30 56
rect 28 55 29 56
rect 27 55 28 56
rect 26 55 27 56
rect 25 55 26 56
rect 24 55 25 56
rect 23 55 24 56
rect 22 55 23 56
rect 21 55 22 56
rect 20 55 21 56
rect 19 55 20 56
rect 195 56 196 57
rect 194 56 195 57
rect 193 56 194 57
rect 183 56 184 57
rect 182 56 183 57
rect 181 56 182 57
rect 180 56 181 57
rect 165 56 166 57
rect 102 56 103 57
rect 101 56 102 57
rect 100 56 101 57
rect 99 56 100 57
rect 98 56 99 57
rect 97 56 98 57
rect 96 56 97 57
rect 95 56 96 57
rect 94 56 95 57
rect 93 56 94 57
rect 92 56 93 57
rect 91 56 92 57
rect 90 56 91 57
rect 89 56 90 57
rect 88 56 89 57
rect 87 56 88 57
rect 86 56 87 57
rect 85 56 86 57
rect 84 56 85 57
rect 83 56 84 57
rect 82 56 83 57
rect 81 56 82 57
rect 80 56 81 57
rect 79 56 80 57
rect 78 56 79 57
rect 77 56 78 57
rect 76 56 77 57
rect 75 56 76 57
rect 74 56 75 57
rect 67 56 68 57
rect 66 56 67 57
rect 65 56 66 57
rect 64 56 65 57
rect 63 56 64 57
rect 62 56 63 57
rect 61 56 62 57
rect 60 56 61 57
rect 59 56 60 57
rect 58 56 59 57
rect 57 56 58 57
rect 56 56 57 57
rect 55 56 56 57
rect 54 56 55 57
rect 53 56 54 57
rect 52 56 53 57
rect 51 56 52 57
rect 50 56 51 57
rect 49 56 50 57
rect 48 56 49 57
rect 47 56 48 57
rect 46 56 47 57
rect 45 56 46 57
rect 44 56 45 57
rect 43 56 44 57
rect 42 56 43 57
rect 41 56 42 57
rect 40 56 41 57
rect 39 56 40 57
rect 38 56 39 57
rect 37 56 38 57
rect 36 56 37 57
rect 35 56 36 57
rect 34 56 35 57
rect 31 56 32 57
rect 30 56 31 57
rect 29 56 30 57
rect 28 56 29 57
rect 27 56 28 57
rect 26 56 27 57
rect 25 56 26 57
rect 24 56 25 57
rect 23 56 24 57
rect 22 56 23 57
rect 21 56 22 57
rect 20 56 21 57
rect 19 56 20 57
rect 196 57 197 58
rect 195 57 196 58
rect 194 57 195 58
rect 183 57 184 58
rect 182 57 183 58
rect 181 57 182 58
rect 124 57 125 58
rect 123 57 124 58
rect 122 57 123 58
rect 121 57 122 58
rect 120 57 121 58
rect 119 57 120 58
rect 118 57 119 58
rect 117 57 118 58
rect 100 57 101 58
rect 99 57 100 58
rect 98 57 99 58
rect 97 57 98 58
rect 96 57 97 58
rect 95 57 96 58
rect 94 57 95 58
rect 93 57 94 58
rect 92 57 93 58
rect 91 57 92 58
rect 90 57 91 58
rect 89 57 90 58
rect 88 57 89 58
rect 87 57 88 58
rect 86 57 87 58
rect 85 57 86 58
rect 84 57 85 58
rect 83 57 84 58
rect 82 57 83 58
rect 81 57 82 58
rect 80 57 81 58
rect 79 57 80 58
rect 78 57 79 58
rect 77 57 78 58
rect 76 57 77 58
rect 75 57 76 58
rect 74 57 75 58
rect 67 57 68 58
rect 66 57 67 58
rect 65 57 66 58
rect 64 57 65 58
rect 63 57 64 58
rect 62 57 63 58
rect 61 57 62 58
rect 60 57 61 58
rect 59 57 60 58
rect 58 57 59 58
rect 57 57 58 58
rect 56 57 57 58
rect 55 57 56 58
rect 54 57 55 58
rect 53 57 54 58
rect 52 57 53 58
rect 51 57 52 58
rect 50 57 51 58
rect 49 57 50 58
rect 48 57 49 58
rect 47 57 48 58
rect 46 57 47 58
rect 45 57 46 58
rect 44 57 45 58
rect 43 57 44 58
rect 42 57 43 58
rect 41 57 42 58
rect 40 57 41 58
rect 39 57 40 58
rect 38 57 39 58
rect 37 57 38 58
rect 36 57 37 58
rect 35 57 36 58
rect 34 57 35 58
rect 31 57 32 58
rect 30 57 31 58
rect 29 57 30 58
rect 28 57 29 58
rect 27 57 28 58
rect 26 57 27 58
rect 25 57 26 58
rect 24 57 25 58
rect 23 57 24 58
rect 22 57 23 58
rect 21 57 22 58
rect 20 57 21 58
rect 19 57 20 58
rect 197 58 198 59
rect 196 58 197 59
rect 195 58 196 59
rect 183 58 184 59
rect 182 58 183 59
rect 181 58 182 59
rect 126 58 127 59
rect 125 58 126 59
rect 124 58 125 59
rect 123 58 124 59
rect 122 58 123 59
rect 121 58 122 59
rect 120 58 121 59
rect 119 58 120 59
rect 118 58 119 59
rect 117 58 118 59
rect 116 58 117 59
rect 115 58 116 59
rect 114 58 115 59
rect 99 58 100 59
rect 98 58 99 59
rect 97 58 98 59
rect 96 58 97 59
rect 95 58 96 59
rect 94 58 95 59
rect 93 58 94 59
rect 92 58 93 59
rect 91 58 92 59
rect 90 58 91 59
rect 89 58 90 59
rect 88 58 89 59
rect 87 58 88 59
rect 86 58 87 59
rect 85 58 86 59
rect 84 58 85 59
rect 83 58 84 59
rect 82 58 83 59
rect 81 58 82 59
rect 80 58 81 59
rect 79 58 80 59
rect 78 58 79 59
rect 77 58 78 59
rect 76 58 77 59
rect 75 58 76 59
rect 74 58 75 59
rect 66 58 67 59
rect 65 58 66 59
rect 64 58 65 59
rect 63 58 64 59
rect 62 58 63 59
rect 61 58 62 59
rect 60 58 61 59
rect 59 58 60 59
rect 58 58 59 59
rect 57 58 58 59
rect 56 58 57 59
rect 55 58 56 59
rect 54 58 55 59
rect 53 58 54 59
rect 52 58 53 59
rect 51 58 52 59
rect 50 58 51 59
rect 49 58 50 59
rect 48 58 49 59
rect 47 58 48 59
rect 46 58 47 59
rect 45 58 46 59
rect 44 58 45 59
rect 43 58 44 59
rect 42 58 43 59
rect 41 58 42 59
rect 40 58 41 59
rect 39 58 40 59
rect 38 58 39 59
rect 37 58 38 59
rect 36 58 37 59
rect 35 58 36 59
rect 34 58 35 59
rect 33 58 34 59
rect 31 58 32 59
rect 30 58 31 59
rect 29 58 30 59
rect 28 58 29 59
rect 27 58 28 59
rect 26 58 27 59
rect 25 58 26 59
rect 24 58 25 59
rect 23 58 24 59
rect 22 58 23 59
rect 21 58 22 59
rect 20 58 21 59
rect 19 58 20 59
rect 199 59 200 60
rect 198 59 199 60
rect 197 59 198 60
rect 196 59 197 60
rect 195 59 196 60
rect 193 59 194 60
rect 192 59 193 60
rect 191 59 192 60
rect 183 59 184 60
rect 182 59 183 60
rect 181 59 182 60
rect 127 59 128 60
rect 126 59 127 60
rect 125 59 126 60
rect 124 59 125 60
rect 123 59 124 60
rect 122 59 123 60
rect 121 59 122 60
rect 120 59 121 60
rect 119 59 120 60
rect 118 59 119 60
rect 117 59 118 60
rect 116 59 117 60
rect 115 59 116 60
rect 114 59 115 60
rect 113 59 114 60
rect 112 59 113 60
rect 99 59 100 60
rect 98 59 99 60
rect 97 59 98 60
rect 96 59 97 60
rect 95 59 96 60
rect 94 59 95 60
rect 93 59 94 60
rect 92 59 93 60
rect 91 59 92 60
rect 90 59 91 60
rect 89 59 90 60
rect 88 59 89 60
rect 87 59 88 60
rect 86 59 87 60
rect 85 59 86 60
rect 84 59 85 60
rect 83 59 84 60
rect 82 59 83 60
rect 81 59 82 60
rect 80 59 81 60
rect 79 59 80 60
rect 78 59 79 60
rect 77 59 78 60
rect 76 59 77 60
rect 75 59 76 60
rect 74 59 75 60
rect 73 59 74 60
rect 66 59 67 60
rect 65 59 66 60
rect 64 59 65 60
rect 63 59 64 60
rect 62 59 63 60
rect 61 59 62 60
rect 60 59 61 60
rect 59 59 60 60
rect 58 59 59 60
rect 57 59 58 60
rect 56 59 57 60
rect 55 59 56 60
rect 54 59 55 60
rect 53 59 54 60
rect 52 59 53 60
rect 51 59 52 60
rect 50 59 51 60
rect 49 59 50 60
rect 48 59 49 60
rect 47 59 48 60
rect 46 59 47 60
rect 45 59 46 60
rect 44 59 45 60
rect 43 59 44 60
rect 42 59 43 60
rect 41 59 42 60
rect 40 59 41 60
rect 39 59 40 60
rect 38 59 39 60
rect 37 59 38 60
rect 36 59 37 60
rect 35 59 36 60
rect 34 59 35 60
rect 33 59 34 60
rect 30 59 31 60
rect 29 59 30 60
rect 28 59 29 60
rect 27 59 28 60
rect 26 59 27 60
rect 25 59 26 60
rect 24 59 25 60
rect 23 59 24 60
rect 22 59 23 60
rect 21 59 22 60
rect 20 59 21 60
rect 19 59 20 60
rect 199 60 200 61
rect 198 60 199 61
rect 197 60 198 61
rect 196 60 197 61
rect 195 60 196 61
rect 194 60 195 61
rect 193 60 194 61
rect 192 60 193 61
rect 191 60 192 61
rect 183 60 184 61
rect 182 60 183 61
rect 181 60 182 61
rect 165 60 166 61
rect 129 60 130 61
rect 128 60 129 61
rect 127 60 128 61
rect 126 60 127 61
rect 125 60 126 61
rect 124 60 125 61
rect 123 60 124 61
rect 122 60 123 61
rect 121 60 122 61
rect 120 60 121 61
rect 119 60 120 61
rect 118 60 119 61
rect 117 60 118 61
rect 116 60 117 61
rect 115 60 116 61
rect 114 60 115 61
rect 113 60 114 61
rect 112 60 113 61
rect 111 60 112 61
rect 110 60 111 61
rect 98 60 99 61
rect 97 60 98 61
rect 96 60 97 61
rect 95 60 96 61
rect 94 60 95 61
rect 93 60 94 61
rect 92 60 93 61
rect 91 60 92 61
rect 90 60 91 61
rect 89 60 90 61
rect 88 60 89 61
rect 87 60 88 61
rect 86 60 87 61
rect 85 60 86 61
rect 84 60 85 61
rect 83 60 84 61
rect 82 60 83 61
rect 81 60 82 61
rect 80 60 81 61
rect 79 60 80 61
rect 78 60 79 61
rect 77 60 78 61
rect 76 60 77 61
rect 75 60 76 61
rect 74 60 75 61
rect 73 60 74 61
rect 65 60 66 61
rect 64 60 65 61
rect 63 60 64 61
rect 62 60 63 61
rect 61 60 62 61
rect 60 60 61 61
rect 59 60 60 61
rect 58 60 59 61
rect 57 60 58 61
rect 56 60 57 61
rect 55 60 56 61
rect 54 60 55 61
rect 53 60 54 61
rect 52 60 53 61
rect 51 60 52 61
rect 50 60 51 61
rect 49 60 50 61
rect 48 60 49 61
rect 47 60 48 61
rect 46 60 47 61
rect 45 60 46 61
rect 44 60 45 61
rect 43 60 44 61
rect 42 60 43 61
rect 41 60 42 61
rect 40 60 41 61
rect 39 60 40 61
rect 38 60 39 61
rect 37 60 38 61
rect 36 60 37 61
rect 35 60 36 61
rect 34 60 35 61
rect 33 60 34 61
rect 32 60 33 61
rect 30 60 31 61
rect 29 60 30 61
rect 28 60 29 61
rect 27 60 28 61
rect 26 60 27 61
rect 25 60 26 61
rect 24 60 25 61
rect 23 60 24 61
rect 22 60 23 61
rect 21 60 22 61
rect 20 60 21 61
rect 182 61 183 62
rect 181 61 182 62
rect 180 61 181 62
rect 165 61 166 62
rect 130 61 131 62
rect 129 61 130 62
rect 128 61 129 62
rect 127 61 128 62
rect 126 61 127 62
rect 125 61 126 62
rect 124 61 125 62
rect 123 61 124 62
rect 122 61 123 62
rect 121 61 122 62
rect 120 61 121 62
rect 119 61 120 62
rect 118 61 119 62
rect 117 61 118 62
rect 116 61 117 62
rect 115 61 116 62
rect 114 61 115 62
rect 113 61 114 62
rect 112 61 113 62
rect 111 61 112 62
rect 110 61 111 62
rect 109 61 110 62
rect 97 61 98 62
rect 96 61 97 62
rect 95 61 96 62
rect 94 61 95 62
rect 93 61 94 62
rect 92 61 93 62
rect 91 61 92 62
rect 90 61 91 62
rect 89 61 90 62
rect 88 61 89 62
rect 87 61 88 62
rect 86 61 87 62
rect 85 61 86 62
rect 84 61 85 62
rect 83 61 84 62
rect 82 61 83 62
rect 81 61 82 62
rect 80 61 81 62
rect 79 61 80 62
rect 78 61 79 62
rect 77 61 78 62
rect 76 61 77 62
rect 75 61 76 62
rect 74 61 75 62
rect 73 61 74 62
rect 72 61 73 62
rect 65 61 66 62
rect 64 61 65 62
rect 63 61 64 62
rect 62 61 63 62
rect 61 61 62 62
rect 60 61 61 62
rect 59 61 60 62
rect 58 61 59 62
rect 57 61 58 62
rect 56 61 57 62
rect 55 61 56 62
rect 54 61 55 62
rect 53 61 54 62
rect 52 61 53 62
rect 51 61 52 62
rect 50 61 51 62
rect 49 61 50 62
rect 48 61 49 62
rect 47 61 48 62
rect 46 61 47 62
rect 45 61 46 62
rect 44 61 45 62
rect 43 61 44 62
rect 42 61 43 62
rect 41 61 42 62
rect 40 61 41 62
rect 39 61 40 62
rect 38 61 39 62
rect 37 61 38 62
rect 36 61 37 62
rect 35 61 36 62
rect 34 61 35 62
rect 33 61 34 62
rect 32 61 33 62
rect 31 61 32 62
rect 30 61 31 62
rect 29 61 30 62
rect 28 61 29 62
rect 27 61 28 62
rect 26 61 27 62
rect 25 61 26 62
rect 24 61 25 62
rect 23 61 24 62
rect 22 61 23 62
rect 21 61 22 62
rect 20 61 21 62
rect 182 62 183 63
rect 181 62 182 63
rect 180 62 181 63
rect 179 62 180 63
rect 166 62 167 63
rect 165 62 166 63
rect 131 62 132 63
rect 130 62 131 63
rect 129 62 130 63
rect 128 62 129 63
rect 127 62 128 63
rect 126 62 127 63
rect 125 62 126 63
rect 124 62 125 63
rect 123 62 124 63
rect 122 62 123 63
rect 121 62 122 63
rect 120 62 121 63
rect 119 62 120 63
rect 118 62 119 63
rect 117 62 118 63
rect 116 62 117 63
rect 115 62 116 63
rect 114 62 115 63
rect 113 62 114 63
rect 112 62 113 63
rect 111 62 112 63
rect 110 62 111 63
rect 109 62 110 63
rect 108 62 109 63
rect 107 62 108 63
rect 97 62 98 63
rect 96 62 97 63
rect 95 62 96 63
rect 94 62 95 63
rect 93 62 94 63
rect 92 62 93 63
rect 91 62 92 63
rect 90 62 91 63
rect 89 62 90 63
rect 88 62 89 63
rect 87 62 88 63
rect 86 62 87 63
rect 85 62 86 63
rect 84 62 85 63
rect 83 62 84 63
rect 82 62 83 63
rect 81 62 82 63
rect 80 62 81 63
rect 79 62 80 63
rect 78 62 79 63
rect 77 62 78 63
rect 76 62 77 63
rect 75 62 76 63
rect 74 62 75 63
rect 73 62 74 63
rect 72 62 73 63
rect 64 62 65 63
rect 63 62 64 63
rect 62 62 63 63
rect 61 62 62 63
rect 60 62 61 63
rect 59 62 60 63
rect 58 62 59 63
rect 57 62 58 63
rect 56 62 57 63
rect 55 62 56 63
rect 54 62 55 63
rect 53 62 54 63
rect 52 62 53 63
rect 51 62 52 63
rect 50 62 51 63
rect 49 62 50 63
rect 48 62 49 63
rect 47 62 48 63
rect 46 62 47 63
rect 45 62 46 63
rect 44 62 45 63
rect 43 62 44 63
rect 42 62 43 63
rect 41 62 42 63
rect 40 62 41 63
rect 39 62 40 63
rect 38 62 39 63
rect 37 62 38 63
rect 36 62 37 63
rect 35 62 36 63
rect 34 62 35 63
rect 33 62 34 63
rect 32 62 33 63
rect 31 62 32 63
rect 30 62 31 63
rect 29 62 30 63
rect 28 62 29 63
rect 27 62 28 63
rect 26 62 27 63
rect 25 62 26 63
rect 24 62 25 63
rect 23 62 24 63
rect 22 62 23 63
rect 21 62 22 63
rect 181 63 182 64
rect 180 63 181 64
rect 179 63 180 64
rect 178 63 179 64
rect 177 63 178 64
rect 176 63 177 64
rect 175 63 176 64
rect 174 63 175 64
rect 173 63 174 64
rect 172 63 173 64
rect 171 63 172 64
rect 170 63 171 64
rect 169 63 170 64
rect 168 63 169 64
rect 167 63 168 64
rect 166 63 167 64
rect 165 63 166 64
rect 132 63 133 64
rect 131 63 132 64
rect 130 63 131 64
rect 129 63 130 64
rect 128 63 129 64
rect 127 63 128 64
rect 126 63 127 64
rect 125 63 126 64
rect 124 63 125 64
rect 123 63 124 64
rect 122 63 123 64
rect 121 63 122 64
rect 120 63 121 64
rect 119 63 120 64
rect 118 63 119 64
rect 117 63 118 64
rect 116 63 117 64
rect 115 63 116 64
rect 114 63 115 64
rect 113 63 114 64
rect 112 63 113 64
rect 111 63 112 64
rect 110 63 111 64
rect 109 63 110 64
rect 108 63 109 64
rect 107 63 108 64
rect 106 63 107 64
rect 96 63 97 64
rect 95 63 96 64
rect 94 63 95 64
rect 93 63 94 64
rect 92 63 93 64
rect 91 63 92 64
rect 90 63 91 64
rect 89 63 90 64
rect 88 63 89 64
rect 87 63 88 64
rect 86 63 87 64
rect 85 63 86 64
rect 84 63 85 64
rect 83 63 84 64
rect 82 63 83 64
rect 81 63 82 64
rect 80 63 81 64
rect 79 63 80 64
rect 78 63 79 64
rect 77 63 78 64
rect 76 63 77 64
rect 75 63 76 64
rect 74 63 75 64
rect 73 63 74 64
rect 72 63 73 64
rect 71 63 72 64
rect 63 63 64 64
rect 62 63 63 64
rect 61 63 62 64
rect 60 63 61 64
rect 59 63 60 64
rect 58 63 59 64
rect 57 63 58 64
rect 56 63 57 64
rect 55 63 56 64
rect 54 63 55 64
rect 53 63 54 64
rect 52 63 53 64
rect 51 63 52 64
rect 50 63 51 64
rect 49 63 50 64
rect 48 63 49 64
rect 47 63 48 64
rect 46 63 47 64
rect 45 63 46 64
rect 44 63 45 64
rect 43 63 44 64
rect 42 63 43 64
rect 41 63 42 64
rect 40 63 41 64
rect 39 63 40 64
rect 38 63 39 64
rect 37 63 38 64
rect 36 63 37 64
rect 35 63 36 64
rect 34 63 35 64
rect 33 63 34 64
rect 32 63 33 64
rect 31 63 32 64
rect 30 63 31 64
rect 29 63 30 64
rect 28 63 29 64
rect 27 63 28 64
rect 26 63 27 64
rect 25 63 26 64
rect 24 63 25 64
rect 23 63 24 64
rect 22 63 23 64
rect 180 64 181 65
rect 179 64 180 65
rect 178 64 179 65
rect 177 64 178 65
rect 176 64 177 65
rect 175 64 176 65
rect 174 64 175 65
rect 173 64 174 65
rect 172 64 173 65
rect 171 64 172 65
rect 170 64 171 65
rect 169 64 170 65
rect 168 64 169 65
rect 167 64 168 65
rect 166 64 167 65
rect 165 64 166 65
rect 132 64 133 65
rect 131 64 132 65
rect 130 64 131 65
rect 129 64 130 65
rect 128 64 129 65
rect 127 64 128 65
rect 126 64 127 65
rect 125 64 126 65
rect 124 64 125 65
rect 123 64 124 65
rect 122 64 123 65
rect 121 64 122 65
rect 120 64 121 65
rect 119 64 120 65
rect 118 64 119 65
rect 117 64 118 65
rect 116 64 117 65
rect 115 64 116 65
rect 114 64 115 65
rect 113 64 114 65
rect 112 64 113 65
rect 111 64 112 65
rect 110 64 111 65
rect 109 64 110 65
rect 108 64 109 65
rect 107 64 108 65
rect 106 64 107 65
rect 105 64 106 65
rect 96 64 97 65
rect 95 64 96 65
rect 94 64 95 65
rect 93 64 94 65
rect 92 64 93 65
rect 91 64 92 65
rect 90 64 91 65
rect 89 64 90 65
rect 88 64 89 65
rect 87 64 88 65
rect 86 64 87 65
rect 85 64 86 65
rect 84 64 85 65
rect 83 64 84 65
rect 82 64 83 65
rect 81 64 82 65
rect 80 64 81 65
rect 79 64 80 65
rect 78 64 79 65
rect 77 64 78 65
rect 76 64 77 65
rect 75 64 76 65
rect 74 64 75 65
rect 73 64 74 65
rect 72 64 73 65
rect 71 64 72 65
rect 62 64 63 65
rect 61 64 62 65
rect 60 64 61 65
rect 59 64 60 65
rect 58 64 59 65
rect 57 64 58 65
rect 56 64 57 65
rect 55 64 56 65
rect 54 64 55 65
rect 53 64 54 65
rect 52 64 53 65
rect 51 64 52 65
rect 50 64 51 65
rect 49 64 50 65
rect 48 64 49 65
rect 47 64 48 65
rect 46 64 47 65
rect 45 64 46 65
rect 44 64 45 65
rect 43 64 44 65
rect 42 64 43 65
rect 41 64 42 65
rect 40 64 41 65
rect 39 64 40 65
rect 38 64 39 65
rect 37 64 38 65
rect 36 64 37 65
rect 35 64 36 65
rect 34 64 35 65
rect 33 64 34 65
rect 32 64 33 65
rect 31 64 32 65
rect 30 64 31 65
rect 29 64 30 65
rect 28 64 29 65
rect 27 64 28 65
rect 26 64 27 65
rect 25 64 26 65
rect 24 64 25 65
rect 23 64 24 65
rect 16 64 17 65
rect 199 65 200 66
rect 198 65 199 66
rect 191 65 192 66
rect 177 65 178 66
rect 169 65 170 66
rect 168 65 169 66
rect 167 65 168 66
rect 166 65 167 66
rect 165 65 166 66
rect 133 65 134 66
rect 132 65 133 66
rect 131 65 132 66
rect 130 65 131 66
rect 129 65 130 66
rect 128 65 129 66
rect 127 65 128 66
rect 126 65 127 66
rect 125 65 126 66
rect 124 65 125 66
rect 123 65 124 66
rect 122 65 123 66
rect 121 65 122 66
rect 120 65 121 66
rect 119 65 120 66
rect 118 65 119 66
rect 117 65 118 66
rect 116 65 117 66
rect 115 65 116 66
rect 114 65 115 66
rect 113 65 114 66
rect 112 65 113 66
rect 111 65 112 66
rect 110 65 111 66
rect 109 65 110 66
rect 108 65 109 66
rect 107 65 108 66
rect 106 65 107 66
rect 105 65 106 66
rect 104 65 105 66
rect 95 65 96 66
rect 94 65 95 66
rect 93 65 94 66
rect 92 65 93 66
rect 91 65 92 66
rect 90 65 91 66
rect 89 65 90 66
rect 88 65 89 66
rect 87 65 88 66
rect 86 65 87 66
rect 85 65 86 66
rect 84 65 85 66
rect 83 65 84 66
rect 82 65 83 66
rect 81 65 82 66
rect 80 65 81 66
rect 79 65 80 66
rect 78 65 79 66
rect 77 65 78 66
rect 76 65 77 66
rect 75 65 76 66
rect 74 65 75 66
rect 73 65 74 66
rect 72 65 73 66
rect 71 65 72 66
rect 70 65 71 66
rect 61 65 62 66
rect 60 65 61 66
rect 59 65 60 66
rect 58 65 59 66
rect 57 65 58 66
rect 56 65 57 66
rect 55 65 56 66
rect 54 65 55 66
rect 53 65 54 66
rect 52 65 53 66
rect 51 65 52 66
rect 50 65 51 66
rect 49 65 50 66
rect 48 65 49 66
rect 47 65 48 66
rect 46 65 47 66
rect 45 65 46 66
rect 44 65 45 66
rect 43 65 44 66
rect 42 65 43 66
rect 41 65 42 66
rect 40 65 41 66
rect 39 65 40 66
rect 38 65 39 66
rect 37 65 38 66
rect 36 65 37 66
rect 35 65 36 66
rect 34 65 35 66
rect 33 65 34 66
rect 32 65 33 66
rect 31 65 32 66
rect 30 65 31 66
rect 29 65 30 66
rect 28 65 29 66
rect 27 65 28 66
rect 26 65 27 66
rect 25 65 26 66
rect 24 65 25 66
rect 23 65 24 66
rect 18 65 19 66
rect 17 65 18 66
rect 16 65 17 66
rect 15 65 16 66
rect 14 65 15 66
rect 198 66 199 67
rect 197 66 198 67
rect 196 66 197 67
rect 195 66 196 67
rect 194 66 195 67
rect 193 66 194 67
rect 192 66 193 67
rect 191 66 192 67
rect 166 66 167 67
rect 165 66 166 67
rect 134 66 135 67
rect 133 66 134 67
rect 132 66 133 67
rect 131 66 132 67
rect 130 66 131 67
rect 129 66 130 67
rect 128 66 129 67
rect 127 66 128 67
rect 126 66 127 67
rect 125 66 126 67
rect 124 66 125 67
rect 123 66 124 67
rect 122 66 123 67
rect 121 66 122 67
rect 120 66 121 67
rect 119 66 120 67
rect 118 66 119 67
rect 117 66 118 67
rect 116 66 117 67
rect 115 66 116 67
rect 114 66 115 67
rect 113 66 114 67
rect 112 66 113 67
rect 111 66 112 67
rect 110 66 111 67
rect 109 66 110 67
rect 108 66 109 67
rect 107 66 108 67
rect 106 66 107 67
rect 105 66 106 67
rect 104 66 105 67
rect 95 66 96 67
rect 94 66 95 67
rect 93 66 94 67
rect 92 66 93 67
rect 91 66 92 67
rect 90 66 91 67
rect 89 66 90 67
rect 88 66 89 67
rect 87 66 88 67
rect 86 66 87 67
rect 85 66 86 67
rect 84 66 85 67
rect 83 66 84 67
rect 82 66 83 67
rect 81 66 82 67
rect 80 66 81 67
rect 79 66 80 67
rect 78 66 79 67
rect 77 66 78 67
rect 76 66 77 67
rect 75 66 76 67
rect 74 66 75 67
rect 73 66 74 67
rect 72 66 73 67
rect 71 66 72 67
rect 70 66 71 67
rect 60 66 61 67
rect 59 66 60 67
rect 58 66 59 67
rect 57 66 58 67
rect 56 66 57 67
rect 55 66 56 67
rect 54 66 55 67
rect 53 66 54 67
rect 52 66 53 67
rect 51 66 52 67
rect 50 66 51 67
rect 49 66 50 67
rect 48 66 49 67
rect 47 66 48 67
rect 46 66 47 67
rect 45 66 46 67
rect 44 66 45 67
rect 43 66 44 67
rect 42 66 43 67
rect 41 66 42 67
rect 40 66 41 67
rect 39 66 40 67
rect 38 66 39 67
rect 37 66 38 67
rect 36 66 37 67
rect 35 66 36 67
rect 34 66 35 67
rect 33 66 34 67
rect 32 66 33 67
rect 31 66 32 67
rect 30 66 31 67
rect 29 66 30 67
rect 28 66 29 67
rect 27 66 28 67
rect 26 66 27 67
rect 25 66 26 67
rect 24 66 25 67
rect 23 66 24 67
rect 18 66 19 67
rect 17 66 18 67
rect 16 66 17 67
rect 15 66 16 67
rect 14 66 15 67
rect 13 66 14 67
rect 12 66 13 67
rect 198 67 199 68
rect 197 67 198 68
rect 196 67 197 68
rect 195 67 196 68
rect 194 67 195 68
rect 193 67 194 68
rect 192 67 193 68
rect 191 67 192 68
rect 165 67 166 68
rect 134 67 135 68
rect 133 67 134 68
rect 132 67 133 68
rect 131 67 132 68
rect 130 67 131 68
rect 129 67 130 68
rect 128 67 129 68
rect 127 67 128 68
rect 126 67 127 68
rect 125 67 126 68
rect 124 67 125 68
rect 123 67 124 68
rect 122 67 123 68
rect 121 67 122 68
rect 120 67 121 68
rect 119 67 120 68
rect 118 67 119 68
rect 117 67 118 68
rect 116 67 117 68
rect 115 67 116 68
rect 114 67 115 68
rect 113 67 114 68
rect 112 67 113 68
rect 111 67 112 68
rect 110 67 111 68
rect 109 67 110 68
rect 108 67 109 68
rect 107 67 108 68
rect 106 67 107 68
rect 105 67 106 68
rect 104 67 105 68
rect 103 67 104 68
rect 94 67 95 68
rect 93 67 94 68
rect 92 67 93 68
rect 91 67 92 68
rect 90 67 91 68
rect 89 67 90 68
rect 88 67 89 68
rect 87 67 88 68
rect 86 67 87 68
rect 85 67 86 68
rect 84 67 85 68
rect 83 67 84 68
rect 82 67 83 68
rect 81 67 82 68
rect 80 67 81 68
rect 79 67 80 68
rect 78 67 79 68
rect 77 67 78 68
rect 76 67 77 68
rect 75 67 76 68
rect 74 67 75 68
rect 73 67 74 68
rect 72 67 73 68
rect 71 67 72 68
rect 70 67 71 68
rect 69 67 70 68
rect 59 67 60 68
rect 58 67 59 68
rect 57 67 58 68
rect 56 67 57 68
rect 55 67 56 68
rect 54 67 55 68
rect 53 67 54 68
rect 52 67 53 68
rect 51 67 52 68
rect 50 67 51 68
rect 49 67 50 68
rect 48 67 49 68
rect 47 67 48 68
rect 46 67 47 68
rect 45 67 46 68
rect 44 67 45 68
rect 43 67 44 68
rect 42 67 43 68
rect 41 67 42 68
rect 40 67 41 68
rect 39 67 40 68
rect 38 67 39 68
rect 37 67 38 68
rect 36 67 37 68
rect 35 67 36 68
rect 34 67 35 68
rect 33 67 34 68
rect 32 67 33 68
rect 31 67 32 68
rect 30 67 31 68
rect 29 67 30 68
rect 28 67 29 68
rect 27 67 28 68
rect 26 67 27 68
rect 25 67 26 68
rect 24 67 25 68
rect 23 67 24 68
rect 19 67 20 68
rect 18 67 19 68
rect 17 67 18 68
rect 16 67 17 68
rect 15 67 16 68
rect 14 67 15 68
rect 13 67 14 68
rect 12 67 13 68
rect 135 68 136 69
rect 134 68 135 69
rect 133 68 134 69
rect 132 68 133 69
rect 131 68 132 69
rect 130 68 131 69
rect 129 68 130 69
rect 128 68 129 69
rect 127 68 128 69
rect 126 68 127 69
rect 125 68 126 69
rect 124 68 125 69
rect 123 68 124 69
rect 122 68 123 69
rect 121 68 122 69
rect 120 68 121 69
rect 119 68 120 69
rect 118 68 119 69
rect 117 68 118 69
rect 116 68 117 69
rect 115 68 116 69
rect 114 68 115 69
rect 113 68 114 69
rect 112 68 113 69
rect 111 68 112 69
rect 110 68 111 69
rect 109 68 110 69
rect 108 68 109 69
rect 107 68 108 69
rect 106 68 107 69
rect 105 68 106 69
rect 104 68 105 69
rect 103 68 104 69
rect 102 68 103 69
rect 94 68 95 69
rect 93 68 94 69
rect 92 68 93 69
rect 91 68 92 69
rect 90 68 91 69
rect 89 68 90 69
rect 88 68 89 69
rect 87 68 88 69
rect 86 68 87 69
rect 85 68 86 69
rect 84 68 85 69
rect 83 68 84 69
rect 82 68 83 69
rect 81 68 82 69
rect 80 68 81 69
rect 79 68 80 69
rect 78 68 79 69
rect 77 68 78 69
rect 76 68 77 69
rect 75 68 76 69
rect 74 68 75 69
rect 73 68 74 69
rect 72 68 73 69
rect 71 68 72 69
rect 70 68 71 69
rect 69 68 70 69
rect 68 68 69 69
rect 57 68 58 69
rect 56 68 57 69
rect 55 68 56 69
rect 54 68 55 69
rect 53 68 54 69
rect 52 68 53 69
rect 51 68 52 69
rect 50 68 51 69
rect 49 68 50 69
rect 48 68 49 69
rect 47 68 48 69
rect 46 68 47 69
rect 45 68 46 69
rect 44 68 45 69
rect 43 68 44 69
rect 42 68 43 69
rect 41 68 42 69
rect 40 68 41 69
rect 39 68 40 69
rect 38 68 39 69
rect 37 68 38 69
rect 36 68 37 69
rect 35 68 36 69
rect 34 68 35 69
rect 33 68 34 69
rect 32 68 33 69
rect 31 68 32 69
rect 30 68 31 69
rect 29 68 30 69
rect 28 68 29 69
rect 27 68 28 69
rect 26 68 27 69
rect 25 68 26 69
rect 24 68 25 69
rect 23 68 24 69
rect 22 68 23 69
rect 18 68 19 69
rect 17 68 18 69
rect 16 68 17 69
rect 15 68 16 69
rect 14 68 15 69
rect 13 68 14 69
rect 12 68 13 69
rect 11 68 12 69
rect 165 69 166 70
rect 136 69 137 70
rect 135 69 136 70
rect 134 69 135 70
rect 133 69 134 70
rect 132 69 133 70
rect 131 69 132 70
rect 130 69 131 70
rect 129 69 130 70
rect 128 69 129 70
rect 127 69 128 70
rect 126 69 127 70
rect 125 69 126 70
rect 124 69 125 70
rect 123 69 124 70
rect 122 69 123 70
rect 121 69 122 70
rect 120 69 121 70
rect 119 69 120 70
rect 118 69 119 70
rect 117 69 118 70
rect 116 69 117 70
rect 115 69 116 70
rect 114 69 115 70
rect 113 69 114 70
rect 112 69 113 70
rect 111 69 112 70
rect 110 69 111 70
rect 109 69 110 70
rect 108 69 109 70
rect 107 69 108 70
rect 106 69 107 70
rect 105 69 106 70
rect 104 69 105 70
rect 103 69 104 70
rect 102 69 103 70
rect 94 69 95 70
rect 93 69 94 70
rect 92 69 93 70
rect 91 69 92 70
rect 90 69 91 70
rect 89 69 90 70
rect 88 69 89 70
rect 87 69 88 70
rect 86 69 87 70
rect 85 69 86 70
rect 84 69 85 70
rect 83 69 84 70
rect 82 69 83 70
rect 81 69 82 70
rect 80 69 81 70
rect 79 69 80 70
rect 78 69 79 70
rect 77 69 78 70
rect 76 69 77 70
rect 75 69 76 70
rect 74 69 75 70
rect 73 69 74 70
rect 72 69 73 70
rect 71 69 72 70
rect 70 69 71 70
rect 69 69 70 70
rect 68 69 69 70
rect 67 69 68 70
rect 56 69 57 70
rect 55 69 56 70
rect 54 69 55 70
rect 53 69 54 70
rect 52 69 53 70
rect 51 69 52 70
rect 50 69 51 70
rect 49 69 50 70
rect 48 69 49 70
rect 47 69 48 70
rect 46 69 47 70
rect 45 69 46 70
rect 44 69 45 70
rect 43 69 44 70
rect 42 69 43 70
rect 41 69 42 70
rect 40 69 41 70
rect 39 69 40 70
rect 38 69 39 70
rect 37 69 38 70
rect 36 69 37 70
rect 35 69 36 70
rect 34 69 35 70
rect 33 69 34 70
rect 32 69 33 70
rect 31 69 32 70
rect 30 69 31 70
rect 29 69 30 70
rect 28 69 29 70
rect 27 69 28 70
rect 26 69 27 70
rect 25 69 26 70
rect 24 69 25 70
rect 23 69 24 70
rect 22 69 23 70
rect 18 69 19 70
rect 17 69 18 70
rect 16 69 17 70
rect 15 69 16 70
rect 14 69 15 70
rect 13 69 14 70
rect 12 69 13 70
rect 11 69 12 70
rect 10 69 11 70
rect 182 70 183 71
rect 165 70 166 71
rect 137 70 138 71
rect 136 70 137 71
rect 135 70 136 71
rect 134 70 135 71
rect 133 70 134 71
rect 132 70 133 71
rect 131 70 132 71
rect 130 70 131 71
rect 129 70 130 71
rect 128 70 129 71
rect 127 70 128 71
rect 126 70 127 71
rect 125 70 126 71
rect 124 70 125 71
rect 123 70 124 71
rect 122 70 123 71
rect 121 70 122 71
rect 120 70 121 71
rect 119 70 120 71
rect 118 70 119 71
rect 117 70 118 71
rect 116 70 117 71
rect 115 70 116 71
rect 114 70 115 71
rect 113 70 114 71
rect 112 70 113 71
rect 111 70 112 71
rect 110 70 111 71
rect 109 70 110 71
rect 108 70 109 71
rect 107 70 108 71
rect 106 70 107 71
rect 105 70 106 71
rect 104 70 105 71
rect 103 70 104 71
rect 102 70 103 71
rect 101 70 102 71
rect 93 70 94 71
rect 92 70 93 71
rect 91 70 92 71
rect 90 70 91 71
rect 89 70 90 71
rect 88 70 89 71
rect 87 70 88 71
rect 86 70 87 71
rect 85 70 86 71
rect 84 70 85 71
rect 83 70 84 71
rect 82 70 83 71
rect 81 70 82 71
rect 80 70 81 71
rect 79 70 80 71
rect 78 70 79 71
rect 77 70 78 71
rect 76 70 77 71
rect 75 70 76 71
rect 74 70 75 71
rect 73 70 74 71
rect 72 70 73 71
rect 71 70 72 71
rect 70 70 71 71
rect 69 70 70 71
rect 68 70 69 71
rect 67 70 68 71
rect 66 70 67 71
rect 54 70 55 71
rect 53 70 54 71
rect 52 70 53 71
rect 51 70 52 71
rect 50 70 51 71
rect 49 70 50 71
rect 48 70 49 71
rect 47 70 48 71
rect 46 70 47 71
rect 45 70 46 71
rect 44 70 45 71
rect 43 70 44 71
rect 42 70 43 71
rect 41 70 42 71
rect 40 70 41 71
rect 39 70 40 71
rect 38 70 39 71
rect 37 70 38 71
rect 36 70 37 71
rect 35 70 36 71
rect 34 70 35 71
rect 33 70 34 71
rect 32 70 33 71
rect 31 70 32 71
rect 30 70 31 71
rect 29 70 30 71
rect 28 70 29 71
rect 27 70 28 71
rect 26 70 27 71
rect 25 70 26 71
rect 24 70 25 71
rect 23 70 24 71
rect 22 70 23 71
rect 21 70 22 71
rect 18 70 19 71
rect 17 70 18 71
rect 16 70 17 71
rect 15 70 16 71
rect 14 70 15 71
rect 13 70 14 71
rect 12 70 13 71
rect 11 70 12 71
rect 10 70 11 71
rect 182 71 183 72
rect 181 71 182 72
rect 166 71 167 72
rect 165 71 166 72
rect 138 71 139 72
rect 137 71 138 72
rect 136 71 137 72
rect 135 71 136 72
rect 124 71 125 72
rect 123 71 124 72
rect 122 71 123 72
rect 121 71 122 72
rect 120 71 121 72
rect 119 71 120 72
rect 118 71 119 72
rect 117 71 118 72
rect 116 71 117 72
rect 115 71 116 72
rect 114 71 115 72
rect 113 71 114 72
rect 112 71 113 72
rect 111 71 112 72
rect 110 71 111 72
rect 109 71 110 72
rect 108 71 109 72
rect 107 71 108 72
rect 106 71 107 72
rect 105 71 106 72
rect 104 71 105 72
rect 103 71 104 72
rect 102 71 103 72
rect 101 71 102 72
rect 100 71 101 72
rect 93 71 94 72
rect 92 71 93 72
rect 91 71 92 72
rect 90 71 91 72
rect 89 71 90 72
rect 88 71 89 72
rect 87 71 88 72
rect 86 71 87 72
rect 85 71 86 72
rect 84 71 85 72
rect 83 71 84 72
rect 82 71 83 72
rect 81 71 82 72
rect 80 71 81 72
rect 79 71 80 72
rect 78 71 79 72
rect 77 71 78 72
rect 76 71 77 72
rect 75 71 76 72
rect 74 71 75 72
rect 73 71 74 72
rect 72 71 73 72
rect 71 71 72 72
rect 70 71 71 72
rect 69 71 70 72
rect 68 71 69 72
rect 67 71 68 72
rect 66 71 67 72
rect 53 71 54 72
rect 52 71 53 72
rect 51 71 52 72
rect 50 71 51 72
rect 49 71 50 72
rect 48 71 49 72
rect 47 71 48 72
rect 46 71 47 72
rect 45 71 46 72
rect 44 71 45 72
rect 43 71 44 72
rect 42 71 43 72
rect 41 71 42 72
rect 40 71 41 72
rect 39 71 40 72
rect 38 71 39 72
rect 37 71 38 72
rect 36 71 37 72
rect 35 71 36 72
rect 34 71 35 72
rect 33 71 34 72
rect 32 71 33 72
rect 31 71 32 72
rect 30 71 31 72
rect 29 71 30 72
rect 28 71 29 72
rect 27 71 28 72
rect 26 71 27 72
rect 25 71 26 72
rect 24 71 25 72
rect 23 71 24 72
rect 22 71 23 72
rect 21 71 22 72
rect 17 71 18 72
rect 16 71 17 72
rect 15 71 16 72
rect 14 71 15 72
rect 13 71 14 72
rect 12 71 13 72
rect 11 71 12 72
rect 10 71 11 72
rect 191 72 192 73
rect 182 72 183 73
rect 181 72 182 73
rect 180 72 181 73
rect 179 72 180 73
rect 178 72 179 73
rect 177 72 178 73
rect 176 72 177 73
rect 175 72 176 73
rect 174 72 175 73
rect 173 72 174 73
rect 172 72 173 73
rect 171 72 172 73
rect 170 72 171 73
rect 169 72 170 73
rect 168 72 169 73
rect 167 72 168 73
rect 166 72 167 73
rect 165 72 166 73
rect 121 72 122 73
rect 120 72 121 73
rect 119 72 120 73
rect 118 72 119 73
rect 117 72 118 73
rect 116 72 117 73
rect 115 72 116 73
rect 114 72 115 73
rect 113 72 114 73
rect 112 72 113 73
rect 111 72 112 73
rect 110 72 111 73
rect 109 72 110 73
rect 108 72 109 73
rect 107 72 108 73
rect 106 72 107 73
rect 105 72 106 73
rect 104 72 105 73
rect 103 72 104 73
rect 102 72 103 73
rect 101 72 102 73
rect 100 72 101 73
rect 92 72 93 73
rect 91 72 92 73
rect 90 72 91 73
rect 89 72 90 73
rect 88 72 89 73
rect 87 72 88 73
rect 86 72 87 73
rect 85 72 86 73
rect 84 72 85 73
rect 83 72 84 73
rect 82 72 83 73
rect 81 72 82 73
rect 80 72 81 73
rect 79 72 80 73
rect 78 72 79 73
rect 77 72 78 73
rect 76 72 77 73
rect 75 72 76 73
rect 74 72 75 73
rect 73 72 74 73
rect 72 72 73 73
rect 71 72 72 73
rect 70 72 71 73
rect 69 72 70 73
rect 68 72 69 73
rect 67 72 68 73
rect 66 72 67 73
rect 65 72 66 73
rect 51 72 52 73
rect 50 72 51 73
rect 49 72 50 73
rect 48 72 49 73
rect 47 72 48 73
rect 46 72 47 73
rect 45 72 46 73
rect 44 72 45 73
rect 43 72 44 73
rect 42 72 43 73
rect 41 72 42 73
rect 40 72 41 73
rect 39 72 40 73
rect 38 72 39 73
rect 37 72 38 73
rect 36 72 37 73
rect 35 72 36 73
rect 34 72 35 73
rect 33 72 34 73
rect 32 72 33 73
rect 31 72 32 73
rect 30 72 31 73
rect 29 72 30 73
rect 28 72 29 73
rect 27 72 28 73
rect 26 72 27 73
rect 25 72 26 73
rect 24 72 25 73
rect 23 72 24 73
rect 22 72 23 73
rect 21 72 22 73
rect 17 72 18 73
rect 16 72 17 73
rect 15 72 16 73
rect 14 72 15 73
rect 13 72 14 73
rect 12 72 13 73
rect 11 72 12 73
rect 10 72 11 73
rect 193 73 194 74
rect 192 73 193 74
rect 191 73 192 74
rect 182 73 183 74
rect 181 73 182 74
rect 180 73 181 74
rect 179 73 180 74
rect 178 73 179 74
rect 177 73 178 74
rect 176 73 177 74
rect 175 73 176 74
rect 174 73 175 74
rect 173 73 174 74
rect 172 73 173 74
rect 171 73 172 74
rect 170 73 171 74
rect 169 73 170 74
rect 168 73 169 74
rect 167 73 168 74
rect 166 73 167 74
rect 165 73 166 74
rect 119 73 120 74
rect 118 73 119 74
rect 117 73 118 74
rect 116 73 117 74
rect 115 73 116 74
rect 114 73 115 74
rect 113 73 114 74
rect 112 73 113 74
rect 111 73 112 74
rect 110 73 111 74
rect 109 73 110 74
rect 108 73 109 74
rect 107 73 108 74
rect 106 73 107 74
rect 105 73 106 74
rect 104 73 105 74
rect 103 73 104 74
rect 102 73 103 74
rect 101 73 102 74
rect 100 73 101 74
rect 99 73 100 74
rect 92 73 93 74
rect 91 73 92 74
rect 90 73 91 74
rect 89 73 90 74
rect 88 73 89 74
rect 87 73 88 74
rect 86 73 87 74
rect 85 73 86 74
rect 84 73 85 74
rect 83 73 84 74
rect 82 73 83 74
rect 81 73 82 74
rect 80 73 81 74
rect 79 73 80 74
rect 78 73 79 74
rect 77 73 78 74
rect 76 73 77 74
rect 75 73 76 74
rect 74 73 75 74
rect 73 73 74 74
rect 72 73 73 74
rect 71 73 72 74
rect 70 73 71 74
rect 69 73 70 74
rect 68 73 69 74
rect 67 73 68 74
rect 66 73 67 74
rect 65 73 66 74
rect 64 73 65 74
rect 63 73 64 74
rect 50 73 51 74
rect 49 73 50 74
rect 48 73 49 74
rect 47 73 48 74
rect 46 73 47 74
rect 45 73 46 74
rect 44 73 45 74
rect 43 73 44 74
rect 42 73 43 74
rect 41 73 42 74
rect 40 73 41 74
rect 39 73 40 74
rect 38 73 39 74
rect 37 73 38 74
rect 36 73 37 74
rect 34 73 35 74
rect 33 73 34 74
rect 32 73 33 74
rect 31 73 32 74
rect 30 73 31 74
rect 29 73 30 74
rect 28 73 29 74
rect 27 73 28 74
rect 26 73 27 74
rect 25 73 26 74
rect 24 73 25 74
rect 23 73 24 74
rect 22 73 23 74
rect 21 73 22 74
rect 20 73 21 74
rect 16 73 17 74
rect 15 73 16 74
rect 14 73 15 74
rect 13 73 14 74
rect 12 73 13 74
rect 11 73 12 74
rect 10 73 11 74
rect 195 74 196 75
rect 194 74 195 75
rect 193 74 194 75
rect 192 74 193 75
rect 191 74 192 75
rect 182 74 183 75
rect 181 74 182 75
rect 170 74 171 75
rect 169 74 170 75
rect 168 74 169 75
rect 167 74 168 75
rect 166 74 167 75
rect 165 74 166 75
rect 117 74 118 75
rect 116 74 117 75
rect 115 74 116 75
rect 114 74 115 75
rect 113 74 114 75
rect 112 74 113 75
rect 111 74 112 75
rect 110 74 111 75
rect 109 74 110 75
rect 108 74 109 75
rect 107 74 108 75
rect 106 74 107 75
rect 105 74 106 75
rect 104 74 105 75
rect 103 74 104 75
rect 102 74 103 75
rect 101 74 102 75
rect 100 74 101 75
rect 99 74 100 75
rect 91 74 92 75
rect 90 74 91 75
rect 89 74 90 75
rect 88 74 89 75
rect 87 74 88 75
rect 86 74 87 75
rect 85 74 86 75
rect 84 74 85 75
rect 83 74 84 75
rect 82 74 83 75
rect 81 74 82 75
rect 80 74 81 75
rect 79 74 80 75
rect 78 74 79 75
rect 77 74 78 75
rect 76 74 77 75
rect 75 74 76 75
rect 74 74 75 75
rect 73 74 74 75
rect 72 74 73 75
rect 71 74 72 75
rect 70 74 71 75
rect 69 74 70 75
rect 68 74 69 75
rect 67 74 68 75
rect 66 74 67 75
rect 65 74 66 75
rect 64 74 65 75
rect 63 74 64 75
rect 62 74 63 75
rect 47 74 48 75
rect 46 74 47 75
rect 45 74 46 75
rect 44 74 45 75
rect 43 74 44 75
rect 42 74 43 75
rect 41 74 42 75
rect 40 74 41 75
rect 32 74 33 75
rect 31 74 32 75
rect 30 74 31 75
rect 29 74 30 75
rect 28 74 29 75
rect 27 74 28 75
rect 26 74 27 75
rect 25 74 26 75
rect 24 74 25 75
rect 23 74 24 75
rect 22 74 23 75
rect 21 74 22 75
rect 20 74 21 75
rect 16 74 17 75
rect 15 74 16 75
rect 14 74 15 75
rect 13 74 14 75
rect 12 74 13 75
rect 11 74 12 75
rect 198 75 199 76
rect 197 75 198 76
rect 196 75 197 76
rect 195 75 196 76
rect 194 75 195 76
rect 193 75 194 76
rect 191 75 192 76
rect 182 75 183 76
rect 171 75 172 76
rect 170 75 171 76
rect 169 75 170 76
rect 168 75 169 76
rect 167 75 168 76
rect 166 75 167 76
rect 116 75 117 76
rect 115 75 116 76
rect 114 75 115 76
rect 113 75 114 76
rect 112 75 113 76
rect 111 75 112 76
rect 110 75 111 76
rect 109 75 110 76
rect 108 75 109 76
rect 107 75 108 76
rect 106 75 107 76
rect 105 75 106 76
rect 104 75 105 76
rect 103 75 104 76
rect 102 75 103 76
rect 101 75 102 76
rect 100 75 101 76
rect 99 75 100 76
rect 98 75 99 76
rect 91 75 92 76
rect 90 75 91 76
rect 89 75 90 76
rect 88 75 89 76
rect 87 75 88 76
rect 86 75 87 76
rect 85 75 86 76
rect 84 75 85 76
rect 83 75 84 76
rect 82 75 83 76
rect 81 75 82 76
rect 80 75 81 76
rect 79 75 80 76
rect 78 75 79 76
rect 77 75 78 76
rect 76 75 77 76
rect 75 75 76 76
rect 74 75 75 76
rect 73 75 74 76
rect 72 75 73 76
rect 71 75 72 76
rect 70 75 71 76
rect 69 75 70 76
rect 68 75 69 76
rect 67 75 68 76
rect 66 75 67 76
rect 65 75 66 76
rect 64 75 65 76
rect 63 75 64 76
rect 62 75 63 76
rect 61 75 62 76
rect 31 75 32 76
rect 30 75 31 76
rect 29 75 30 76
rect 28 75 29 76
rect 27 75 28 76
rect 26 75 27 76
rect 25 75 26 76
rect 24 75 25 76
rect 23 75 24 76
rect 22 75 23 76
rect 21 75 22 76
rect 20 75 21 76
rect 16 75 17 76
rect 15 75 16 76
rect 14 75 15 76
rect 13 75 14 76
rect 12 75 13 76
rect 11 75 12 76
rect 199 76 200 77
rect 198 76 199 77
rect 197 76 198 77
rect 196 76 197 77
rect 182 76 183 77
rect 172 76 173 77
rect 171 76 172 77
rect 170 76 171 77
rect 169 76 170 77
rect 168 76 169 77
rect 167 76 168 77
rect 115 76 116 77
rect 114 76 115 77
rect 113 76 114 77
rect 112 76 113 77
rect 111 76 112 77
rect 110 76 111 77
rect 109 76 110 77
rect 108 76 109 77
rect 107 76 108 77
rect 106 76 107 77
rect 105 76 106 77
rect 104 76 105 77
rect 103 76 104 77
rect 102 76 103 77
rect 101 76 102 77
rect 100 76 101 77
rect 99 76 100 77
rect 98 76 99 77
rect 90 76 91 77
rect 89 76 90 77
rect 88 76 89 77
rect 87 76 88 77
rect 86 76 87 77
rect 85 76 86 77
rect 84 76 85 77
rect 83 76 84 77
rect 82 76 83 77
rect 81 76 82 77
rect 80 76 81 77
rect 79 76 80 77
rect 78 76 79 77
rect 77 76 78 77
rect 76 76 77 77
rect 75 76 76 77
rect 74 76 75 77
rect 73 76 74 77
rect 72 76 73 77
rect 71 76 72 77
rect 70 76 71 77
rect 69 76 70 77
rect 68 76 69 77
rect 67 76 68 77
rect 66 76 67 77
rect 65 76 66 77
rect 64 76 65 77
rect 63 76 64 77
rect 62 76 63 77
rect 61 76 62 77
rect 60 76 61 77
rect 59 76 60 77
rect 30 76 31 77
rect 29 76 30 77
rect 28 76 29 77
rect 27 76 28 77
rect 26 76 27 77
rect 25 76 26 77
rect 24 76 25 77
rect 23 76 24 77
rect 22 76 23 77
rect 21 76 22 77
rect 16 76 17 77
rect 15 76 16 77
rect 14 76 15 77
rect 13 76 14 77
rect 12 76 13 77
rect 11 76 12 77
rect 197 77 198 78
rect 196 77 197 78
rect 195 77 196 78
rect 173 77 174 78
rect 172 77 173 78
rect 171 77 172 78
rect 170 77 171 78
rect 169 77 170 78
rect 168 77 169 78
rect 114 77 115 78
rect 113 77 114 78
rect 112 77 113 78
rect 111 77 112 78
rect 110 77 111 78
rect 109 77 110 78
rect 108 77 109 78
rect 107 77 108 78
rect 106 77 107 78
rect 105 77 106 78
rect 104 77 105 78
rect 103 77 104 78
rect 102 77 103 78
rect 101 77 102 78
rect 100 77 101 78
rect 99 77 100 78
rect 98 77 99 78
rect 97 77 98 78
rect 89 77 90 78
rect 88 77 89 78
rect 87 77 88 78
rect 86 77 87 78
rect 85 77 86 78
rect 84 77 85 78
rect 83 77 84 78
rect 82 77 83 78
rect 81 77 82 78
rect 80 77 81 78
rect 79 77 80 78
rect 78 77 79 78
rect 77 77 78 78
rect 76 77 77 78
rect 75 77 76 78
rect 74 77 75 78
rect 73 77 74 78
rect 72 77 73 78
rect 71 77 72 78
rect 70 77 71 78
rect 69 77 70 78
rect 68 77 69 78
rect 67 77 68 78
rect 66 77 67 78
rect 65 77 66 78
rect 64 77 65 78
rect 63 77 64 78
rect 62 77 63 78
rect 61 77 62 78
rect 60 77 61 78
rect 59 77 60 78
rect 58 77 59 78
rect 30 77 31 78
rect 29 77 30 78
rect 28 77 29 78
rect 27 77 28 78
rect 26 77 27 78
rect 25 77 26 78
rect 24 77 25 78
rect 23 77 24 78
rect 22 77 23 78
rect 21 77 22 78
rect 16 77 17 78
rect 15 77 16 78
rect 14 77 15 78
rect 13 77 14 78
rect 12 77 13 78
rect 195 78 196 79
rect 194 78 195 79
rect 193 78 194 79
rect 192 78 193 79
rect 191 78 192 79
rect 174 78 175 79
rect 173 78 174 79
rect 172 78 173 79
rect 171 78 172 79
rect 170 78 171 79
rect 169 78 170 79
rect 113 78 114 79
rect 112 78 113 79
rect 111 78 112 79
rect 110 78 111 79
rect 109 78 110 79
rect 108 78 109 79
rect 107 78 108 79
rect 106 78 107 79
rect 105 78 106 79
rect 104 78 105 79
rect 103 78 104 79
rect 102 78 103 79
rect 101 78 102 79
rect 100 78 101 79
rect 99 78 100 79
rect 98 78 99 79
rect 97 78 98 79
rect 89 78 90 79
rect 88 78 89 79
rect 87 78 88 79
rect 86 78 87 79
rect 85 78 86 79
rect 84 78 85 79
rect 83 78 84 79
rect 82 78 83 79
rect 81 78 82 79
rect 80 78 81 79
rect 79 78 80 79
rect 78 78 79 79
rect 77 78 78 79
rect 76 78 77 79
rect 75 78 76 79
rect 74 78 75 79
rect 73 78 74 79
rect 72 78 73 79
rect 71 78 72 79
rect 70 78 71 79
rect 69 78 70 79
rect 68 78 69 79
rect 67 78 68 79
rect 66 78 67 79
rect 65 78 66 79
rect 64 78 65 79
rect 63 78 64 79
rect 62 78 63 79
rect 61 78 62 79
rect 60 78 61 79
rect 59 78 60 79
rect 58 78 59 79
rect 57 78 58 79
rect 56 78 57 79
rect 29 78 30 79
rect 28 78 29 79
rect 27 78 28 79
rect 26 78 27 79
rect 25 78 26 79
rect 24 78 25 79
rect 23 78 24 79
rect 22 78 23 79
rect 16 78 17 79
rect 15 78 16 79
rect 14 78 15 79
rect 13 78 14 79
rect 12 78 13 79
rect 192 79 193 80
rect 191 79 192 80
rect 176 79 177 80
rect 175 79 176 80
rect 174 79 175 80
rect 173 79 174 80
rect 172 79 173 80
rect 171 79 172 80
rect 170 79 171 80
rect 133 79 134 80
rect 132 79 133 80
rect 131 79 132 80
rect 130 79 131 80
rect 129 79 130 80
rect 128 79 129 80
rect 112 79 113 80
rect 111 79 112 80
rect 110 79 111 80
rect 109 79 110 80
rect 108 79 109 80
rect 107 79 108 80
rect 106 79 107 80
rect 105 79 106 80
rect 104 79 105 80
rect 103 79 104 80
rect 102 79 103 80
rect 101 79 102 80
rect 100 79 101 80
rect 99 79 100 80
rect 98 79 99 80
rect 97 79 98 80
rect 96 79 97 80
rect 88 79 89 80
rect 87 79 88 80
rect 86 79 87 80
rect 85 79 86 80
rect 84 79 85 80
rect 83 79 84 80
rect 82 79 83 80
rect 81 79 82 80
rect 80 79 81 80
rect 79 79 80 80
rect 78 79 79 80
rect 77 79 78 80
rect 76 79 77 80
rect 75 79 76 80
rect 74 79 75 80
rect 73 79 74 80
rect 72 79 73 80
rect 71 79 72 80
rect 70 79 71 80
rect 69 79 70 80
rect 68 79 69 80
rect 67 79 68 80
rect 66 79 67 80
rect 65 79 66 80
rect 64 79 65 80
rect 63 79 64 80
rect 62 79 63 80
rect 61 79 62 80
rect 60 79 61 80
rect 59 79 60 80
rect 58 79 59 80
rect 57 79 58 80
rect 56 79 57 80
rect 55 79 56 80
rect 54 79 55 80
rect 53 79 54 80
rect 28 79 29 80
rect 27 79 28 80
rect 26 79 27 80
rect 25 79 26 80
rect 24 79 25 80
rect 23 79 24 80
rect 22 79 23 80
rect 16 79 17 80
rect 15 79 16 80
rect 14 79 15 80
rect 13 79 14 80
rect 12 79 13 80
rect 177 80 178 81
rect 176 80 177 81
rect 175 80 176 81
rect 174 80 175 81
rect 173 80 174 81
rect 172 80 173 81
rect 137 80 138 81
rect 136 80 137 81
rect 135 80 136 81
rect 134 80 135 81
rect 133 80 134 81
rect 132 80 133 81
rect 131 80 132 81
rect 130 80 131 81
rect 129 80 130 81
rect 128 80 129 81
rect 127 80 128 81
rect 126 80 127 81
rect 125 80 126 81
rect 124 80 125 81
rect 111 80 112 81
rect 110 80 111 81
rect 109 80 110 81
rect 108 80 109 81
rect 107 80 108 81
rect 106 80 107 81
rect 105 80 106 81
rect 104 80 105 81
rect 103 80 104 81
rect 102 80 103 81
rect 101 80 102 81
rect 100 80 101 81
rect 99 80 100 81
rect 98 80 99 81
rect 97 80 98 81
rect 96 80 97 81
rect 87 80 88 81
rect 86 80 87 81
rect 85 80 86 81
rect 84 80 85 81
rect 83 80 84 81
rect 82 80 83 81
rect 81 80 82 81
rect 80 80 81 81
rect 79 80 80 81
rect 78 80 79 81
rect 77 80 78 81
rect 76 80 77 81
rect 75 80 76 81
rect 74 80 75 81
rect 73 80 74 81
rect 72 80 73 81
rect 71 80 72 81
rect 70 80 71 81
rect 69 80 70 81
rect 68 80 69 81
rect 67 80 68 81
rect 66 80 67 81
rect 65 80 66 81
rect 64 80 65 81
rect 63 80 64 81
rect 62 80 63 81
rect 61 80 62 81
rect 60 80 61 81
rect 59 80 60 81
rect 58 80 59 81
rect 57 80 58 81
rect 56 80 57 81
rect 55 80 56 81
rect 54 80 55 81
rect 53 80 54 81
rect 52 80 53 81
rect 51 80 52 81
rect 50 80 51 81
rect 37 80 38 81
rect 36 80 37 81
rect 35 80 36 81
rect 26 80 27 81
rect 25 80 26 81
rect 24 80 25 81
rect 16 80 17 81
rect 15 80 16 81
rect 14 80 15 81
rect 13 80 14 81
rect 12 80 13 81
rect 178 81 179 82
rect 177 81 178 82
rect 176 81 177 82
rect 175 81 176 82
rect 174 81 175 82
rect 173 81 174 82
rect 139 81 140 82
rect 138 81 139 82
rect 137 81 138 82
rect 136 81 137 82
rect 135 81 136 82
rect 134 81 135 82
rect 133 81 134 82
rect 132 81 133 82
rect 131 81 132 82
rect 130 81 131 82
rect 129 81 130 82
rect 128 81 129 82
rect 127 81 128 82
rect 126 81 127 82
rect 125 81 126 82
rect 124 81 125 82
rect 123 81 124 82
rect 122 81 123 82
rect 121 81 122 82
rect 111 81 112 82
rect 110 81 111 82
rect 109 81 110 82
rect 108 81 109 82
rect 107 81 108 82
rect 106 81 107 82
rect 105 81 106 82
rect 104 81 105 82
rect 103 81 104 82
rect 102 81 103 82
rect 101 81 102 82
rect 100 81 101 82
rect 99 81 100 82
rect 98 81 99 82
rect 97 81 98 82
rect 96 81 97 82
rect 95 81 96 82
rect 86 81 87 82
rect 85 81 86 82
rect 84 81 85 82
rect 83 81 84 82
rect 82 81 83 82
rect 81 81 82 82
rect 80 81 81 82
rect 79 81 80 82
rect 78 81 79 82
rect 77 81 78 82
rect 76 81 77 82
rect 75 81 76 82
rect 74 81 75 82
rect 73 81 74 82
rect 72 81 73 82
rect 71 81 72 82
rect 70 81 71 82
rect 69 81 70 82
rect 68 81 69 82
rect 67 81 68 82
rect 66 81 67 82
rect 65 81 66 82
rect 64 81 65 82
rect 63 81 64 82
rect 62 81 63 82
rect 61 81 62 82
rect 60 81 61 82
rect 59 81 60 82
rect 58 81 59 82
rect 57 81 58 82
rect 56 81 57 82
rect 55 81 56 82
rect 54 81 55 82
rect 53 81 54 82
rect 52 81 53 82
rect 51 81 52 82
rect 50 81 51 82
rect 49 81 50 82
rect 48 81 49 82
rect 47 81 48 82
rect 46 81 47 82
rect 45 81 46 82
rect 44 81 45 82
rect 43 81 44 82
rect 42 81 43 82
rect 40 81 41 82
rect 39 81 40 82
rect 38 81 39 82
rect 37 81 38 82
rect 36 81 37 82
rect 35 81 36 82
rect 17 81 18 82
rect 16 81 17 82
rect 15 81 16 82
rect 14 81 15 82
rect 13 81 14 82
rect 12 81 13 82
rect 179 82 180 83
rect 178 82 179 83
rect 177 82 178 83
rect 176 82 177 83
rect 175 82 176 83
rect 174 82 175 83
rect 165 82 166 83
rect 140 82 141 83
rect 139 82 140 83
rect 138 82 139 83
rect 137 82 138 83
rect 136 82 137 83
rect 135 82 136 83
rect 134 82 135 83
rect 133 82 134 83
rect 132 82 133 83
rect 131 82 132 83
rect 130 82 131 83
rect 129 82 130 83
rect 128 82 129 83
rect 127 82 128 83
rect 126 82 127 83
rect 125 82 126 83
rect 124 82 125 83
rect 123 82 124 83
rect 122 82 123 83
rect 121 82 122 83
rect 120 82 121 83
rect 119 82 120 83
rect 110 82 111 83
rect 109 82 110 83
rect 108 82 109 83
rect 107 82 108 83
rect 106 82 107 83
rect 105 82 106 83
rect 104 82 105 83
rect 103 82 104 83
rect 102 82 103 83
rect 101 82 102 83
rect 100 82 101 83
rect 99 82 100 83
rect 98 82 99 83
rect 97 82 98 83
rect 96 82 97 83
rect 95 82 96 83
rect 94 82 95 83
rect 85 82 86 83
rect 84 82 85 83
rect 83 82 84 83
rect 82 82 83 83
rect 81 82 82 83
rect 80 82 81 83
rect 79 82 80 83
rect 78 82 79 83
rect 77 82 78 83
rect 76 82 77 83
rect 75 82 76 83
rect 74 82 75 83
rect 73 82 74 83
rect 72 82 73 83
rect 71 82 72 83
rect 70 82 71 83
rect 69 82 70 83
rect 68 82 69 83
rect 67 82 68 83
rect 66 82 67 83
rect 65 82 66 83
rect 64 82 65 83
rect 63 82 64 83
rect 62 82 63 83
rect 61 82 62 83
rect 60 82 61 83
rect 59 82 60 83
rect 58 82 59 83
rect 57 82 58 83
rect 56 82 57 83
rect 55 82 56 83
rect 54 82 55 83
rect 53 82 54 83
rect 52 82 53 83
rect 51 82 52 83
rect 50 82 51 83
rect 49 82 50 83
rect 48 82 49 83
rect 47 82 48 83
rect 46 82 47 83
rect 45 82 46 83
rect 44 82 45 83
rect 43 82 44 83
rect 42 82 43 83
rect 41 82 42 83
rect 40 82 41 83
rect 39 82 40 83
rect 38 82 39 83
rect 37 82 38 83
rect 36 82 37 83
rect 35 82 36 83
rect 17 82 18 83
rect 16 82 17 83
rect 15 82 16 83
rect 14 82 15 83
rect 13 82 14 83
rect 12 82 13 83
rect 181 83 182 84
rect 180 83 181 84
rect 179 83 180 84
rect 178 83 179 84
rect 177 83 178 84
rect 176 83 177 84
rect 175 83 176 84
rect 165 83 166 84
rect 142 83 143 84
rect 141 83 142 84
rect 140 83 141 84
rect 139 83 140 84
rect 138 83 139 84
rect 137 83 138 84
rect 136 83 137 84
rect 135 83 136 84
rect 134 83 135 84
rect 133 83 134 84
rect 132 83 133 84
rect 131 83 132 84
rect 130 83 131 84
rect 129 83 130 84
rect 128 83 129 84
rect 127 83 128 84
rect 126 83 127 84
rect 125 83 126 84
rect 124 83 125 84
rect 123 83 124 84
rect 122 83 123 84
rect 121 83 122 84
rect 120 83 121 84
rect 119 83 120 84
rect 118 83 119 84
rect 117 83 118 84
rect 109 83 110 84
rect 108 83 109 84
rect 107 83 108 84
rect 106 83 107 84
rect 105 83 106 84
rect 104 83 105 84
rect 103 83 104 84
rect 102 83 103 84
rect 101 83 102 84
rect 100 83 101 84
rect 99 83 100 84
rect 98 83 99 84
rect 97 83 98 84
rect 96 83 97 84
rect 95 83 96 84
rect 94 83 95 84
rect 84 83 85 84
rect 83 83 84 84
rect 82 83 83 84
rect 81 83 82 84
rect 80 83 81 84
rect 79 83 80 84
rect 78 83 79 84
rect 77 83 78 84
rect 76 83 77 84
rect 75 83 76 84
rect 74 83 75 84
rect 73 83 74 84
rect 72 83 73 84
rect 71 83 72 84
rect 70 83 71 84
rect 69 83 70 84
rect 68 83 69 84
rect 67 83 68 84
rect 66 83 67 84
rect 65 83 66 84
rect 64 83 65 84
rect 63 83 64 84
rect 62 83 63 84
rect 61 83 62 84
rect 60 83 61 84
rect 59 83 60 84
rect 58 83 59 84
rect 57 83 58 84
rect 56 83 57 84
rect 55 83 56 84
rect 54 83 55 84
rect 53 83 54 84
rect 52 83 53 84
rect 51 83 52 84
rect 50 83 51 84
rect 49 83 50 84
rect 48 83 49 84
rect 47 83 48 84
rect 46 83 47 84
rect 45 83 46 84
rect 44 83 45 84
rect 43 83 44 84
rect 42 83 43 84
rect 41 83 42 84
rect 40 83 41 84
rect 39 83 40 84
rect 38 83 39 84
rect 37 83 38 84
rect 36 83 37 84
rect 35 83 36 84
rect 18 83 19 84
rect 17 83 18 84
rect 16 83 17 84
rect 15 83 16 84
rect 14 83 15 84
rect 13 83 14 84
rect 12 83 13 84
rect 199 84 200 85
rect 198 84 199 85
rect 191 84 192 85
rect 182 84 183 85
rect 181 84 182 85
rect 180 84 181 85
rect 179 84 180 85
rect 178 84 179 85
rect 177 84 178 85
rect 176 84 177 85
rect 166 84 167 85
rect 165 84 166 85
rect 143 84 144 85
rect 142 84 143 85
rect 141 84 142 85
rect 140 84 141 85
rect 139 84 140 85
rect 138 84 139 85
rect 137 84 138 85
rect 136 84 137 85
rect 135 84 136 85
rect 134 84 135 85
rect 133 84 134 85
rect 132 84 133 85
rect 131 84 132 85
rect 130 84 131 85
rect 129 84 130 85
rect 128 84 129 85
rect 127 84 128 85
rect 126 84 127 85
rect 125 84 126 85
rect 124 84 125 85
rect 123 84 124 85
rect 122 84 123 85
rect 121 84 122 85
rect 120 84 121 85
rect 119 84 120 85
rect 118 84 119 85
rect 117 84 118 85
rect 116 84 117 85
rect 109 84 110 85
rect 108 84 109 85
rect 107 84 108 85
rect 106 84 107 85
rect 105 84 106 85
rect 104 84 105 85
rect 103 84 104 85
rect 102 84 103 85
rect 101 84 102 85
rect 100 84 101 85
rect 99 84 100 85
rect 98 84 99 85
rect 97 84 98 85
rect 96 84 97 85
rect 95 84 96 85
rect 94 84 95 85
rect 93 84 94 85
rect 83 84 84 85
rect 82 84 83 85
rect 81 84 82 85
rect 80 84 81 85
rect 79 84 80 85
rect 78 84 79 85
rect 77 84 78 85
rect 76 84 77 85
rect 75 84 76 85
rect 74 84 75 85
rect 73 84 74 85
rect 72 84 73 85
rect 71 84 72 85
rect 70 84 71 85
rect 69 84 70 85
rect 68 84 69 85
rect 67 84 68 85
rect 66 84 67 85
rect 65 84 66 85
rect 64 84 65 85
rect 63 84 64 85
rect 62 84 63 85
rect 61 84 62 85
rect 60 84 61 85
rect 59 84 60 85
rect 58 84 59 85
rect 57 84 58 85
rect 56 84 57 85
rect 55 84 56 85
rect 54 84 55 85
rect 53 84 54 85
rect 52 84 53 85
rect 51 84 52 85
rect 50 84 51 85
rect 49 84 50 85
rect 48 84 49 85
rect 47 84 48 85
rect 46 84 47 85
rect 45 84 46 85
rect 44 84 45 85
rect 43 84 44 85
rect 42 84 43 85
rect 41 84 42 85
rect 40 84 41 85
rect 39 84 40 85
rect 38 84 39 85
rect 37 84 38 85
rect 36 84 37 85
rect 35 84 36 85
rect 18 84 19 85
rect 17 84 18 85
rect 16 84 17 85
rect 15 84 16 85
rect 14 84 15 85
rect 13 84 14 85
rect 12 84 13 85
rect 198 85 199 86
rect 197 85 198 86
rect 196 85 197 86
rect 195 85 196 86
rect 194 85 195 86
rect 193 85 194 86
rect 192 85 193 86
rect 191 85 192 86
rect 183 85 184 86
rect 182 85 183 86
rect 181 85 182 86
rect 180 85 181 86
rect 179 85 180 86
rect 178 85 179 86
rect 177 85 178 86
rect 176 85 177 86
rect 175 85 176 86
rect 174 85 175 86
rect 173 85 174 86
rect 172 85 173 86
rect 171 85 172 86
rect 170 85 171 86
rect 169 85 170 86
rect 168 85 169 86
rect 167 85 168 86
rect 166 85 167 86
rect 165 85 166 86
rect 144 85 145 86
rect 143 85 144 86
rect 142 85 143 86
rect 141 85 142 86
rect 140 85 141 86
rect 139 85 140 86
rect 138 85 139 86
rect 137 85 138 86
rect 136 85 137 86
rect 135 85 136 86
rect 134 85 135 86
rect 133 85 134 86
rect 132 85 133 86
rect 131 85 132 86
rect 130 85 131 86
rect 129 85 130 86
rect 128 85 129 86
rect 127 85 128 86
rect 126 85 127 86
rect 125 85 126 86
rect 124 85 125 86
rect 123 85 124 86
rect 122 85 123 86
rect 121 85 122 86
rect 120 85 121 86
rect 119 85 120 86
rect 118 85 119 86
rect 117 85 118 86
rect 116 85 117 86
rect 115 85 116 86
rect 108 85 109 86
rect 107 85 108 86
rect 106 85 107 86
rect 105 85 106 86
rect 104 85 105 86
rect 103 85 104 86
rect 102 85 103 86
rect 101 85 102 86
rect 100 85 101 86
rect 99 85 100 86
rect 98 85 99 86
rect 97 85 98 86
rect 96 85 97 86
rect 95 85 96 86
rect 94 85 95 86
rect 93 85 94 86
rect 92 85 93 86
rect 82 85 83 86
rect 81 85 82 86
rect 80 85 81 86
rect 79 85 80 86
rect 78 85 79 86
rect 77 85 78 86
rect 76 85 77 86
rect 75 85 76 86
rect 74 85 75 86
rect 73 85 74 86
rect 72 85 73 86
rect 71 85 72 86
rect 70 85 71 86
rect 69 85 70 86
rect 68 85 69 86
rect 67 85 68 86
rect 66 85 67 86
rect 65 85 66 86
rect 64 85 65 86
rect 63 85 64 86
rect 62 85 63 86
rect 61 85 62 86
rect 60 85 61 86
rect 59 85 60 86
rect 58 85 59 86
rect 57 85 58 86
rect 56 85 57 86
rect 55 85 56 86
rect 54 85 55 86
rect 53 85 54 86
rect 52 85 53 86
rect 51 85 52 86
rect 50 85 51 86
rect 49 85 50 86
rect 48 85 49 86
rect 47 85 48 86
rect 46 85 47 86
rect 45 85 46 86
rect 44 85 45 86
rect 43 85 44 86
rect 42 85 43 86
rect 41 85 42 86
rect 40 85 41 86
rect 39 85 40 86
rect 38 85 39 86
rect 37 85 38 86
rect 36 85 37 86
rect 35 85 36 86
rect 27 85 28 86
rect 26 85 27 86
rect 25 85 26 86
rect 19 85 20 86
rect 18 85 19 86
rect 17 85 18 86
rect 16 85 17 86
rect 15 85 16 86
rect 14 85 15 86
rect 13 85 14 86
rect 12 85 13 86
rect 199 86 200 87
rect 198 86 199 87
rect 197 86 198 87
rect 196 86 197 87
rect 195 86 196 87
rect 194 86 195 87
rect 193 86 194 87
rect 192 86 193 87
rect 191 86 192 87
rect 182 86 183 87
rect 181 86 182 87
rect 180 86 181 87
rect 179 86 180 87
rect 178 86 179 87
rect 177 86 178 87
rect 176 86 177 87
rect 175 86 176 87
rect 174 86 175 87
rect 173 86 174 87
rect 172 86 173 87
rect 171 86 172 87
rect 170 86 171 87
rect 169 86 170 87
rect 168 86 169 87
rect 167 86 168 87
rect 166 86 167 87
rect 165 86 166 87
rect 145 86 146 87
rect 144 86 145 87
rect 143 86 144 87
rect 142 86 143 87
rect 141 86 142 87
rect 140 86 141 87
rect 139 86 140 87
rect 138 86 139 87
rect 137 86 138 87
rect 136 86 137 87
rect 135 86 136 87
rect 134 86 135 87
rect 133 86 134 87
rect 132 86 133 87
rect 131 86 132 87
rect 130 86 131 87
rect 129 86 130 87
rect 128 86 129 87
rect 127 86 128 87
rect 126 86 127 87
rect 125 86 126 87
rect 124 86 125 87
rect 123 86 124 87
rect 122 86 123 87
rect 121 86 122 87
rect 120 86 121 87
rect 119 86 120 87
rect 118 86 119 87
rect 117 86 118 87
rect 116 86 117 87
rect 115 86 116 87
rect 114 86 115 87
rect 113 86 114 87
rect 108 86 109 87
rect 107 86 108 87
rect 106 86 107 87
rect 105 86 106 87
rect 104 86 105 87
rect 103 86 104 87
rect 102 86 103 87
rect 101 86 102 87
rect 100 86 101 87
rect 99 86 100 87
rect 98 86 99 87
rect 97 86 98 87
rect 96 86 97 87
rect 95 86 96 87
rect 94 86 95 87
rect 93 86 94 87
rect 92 86 93 87
rect 81 86 82 87
rect 80 86 81 87
rect 79 86 80 87
rect 78 86 79 87
rect 77 86 78 87
rect 76 86 77 87
rect 75 86 76 87
rect 74 86 75 87
rect 73 86 74 87
rect 72 86 73 87
rect 71 86 72 87
rect 70 86 71 87
rect 69 86 70 87
rect 68 86 69 87
rect 67 86 68 87
rect 66 86 67 87
rect 65 86 66 87
rect 64 86 65 87
rect 63 86 64 87
rect 62 86 63 87
rect 61 86 62 87
rect 60 86 61 87
rect 59 86 60 87
rect 58 86 59 87
rect 57 86 58 87
rect 56 86 57 87
rect 55 86 56 87
rect 54 86 55 87
rect 53 86 54 87
rect 52 86 53 87
rect 51 86 52 87
rect 50 86 51 87
rect 49 86 50 87
rect 48 86 49 87
rect 47 86 48 87
rect 46 86 47 87
rect 45 86 46 87
rect 44 86 45 87
rect 43 86 44 87
rect 42 86 43 87
rect 41 86 42 87
rect 40 86 41 87
rect 39 86 40 87
rect 38 86 39 87
rect 37 86 38 87
rect 36 86 37 87
rect 35 86 36 87
rect 28 86 29 87
rect 27 86 28 87
rect 26 86 27 87
rect 25 86 26 87
rect 24 86 25 87
rect 23 86 24 87
rect 22 86 23 87
rect 21 86 22 87
rect 20 86 21 87
rect 19 86 20 87
rect 18 86 19 87
rect 17 86 18 87
rect 16 86 17 87
rect 15 86 16 87
rect 14 86 15 87
rect 13 86 14 87
rect 12 86 13 87
rect 199 87 200 88
rect 195 87 196 88
rect 194 87 195 88
rect 166 87 167 88
rect 165 87 166 88
rect 146 87 147 88
rect 145 87 146 88
rect 144 87 145 88
rect 143 87 144 88
rect 142 87 143 88
rect 141 87 142 88
rect 140 87 141 88
rect 139 87 140 88
rect 138 87 139 88
rect 137 87 138 88
rect 136 87 137 88
rect 135 87 136 88
rect 134 87 135 88
rect 133 87 134 88
rect 132 87 133 88
rect 131 87 132 88
rect 130 87 131 88
rect 129 87 130 88
rect 128 87 129 88
rect 127 87 128 88
rect 126 87 127 88
rect 125 87 126 88
rect 124 87 125 88
rect 123 87 124 88
rect 122 87 123 88
rect 121 87 122 88
rect 120 87 121 88
rect 119 87 120 88
rect 118 87 119 88
rect 117 87 118 88
rect 116 87 117 88
rect 115 87 116 88
rect 114 87 115 88
rect 113 87 114 88
rect 112 87 113 88
rect 107 87 108 88
rect 106 87 107 88
rect 105 87 106 88
rect 104 87 105 88
rect 103 87 104 88
rect 102 87 103 88
rect 101 87 102 88
rect 100 87 101 88
rect 99 87 100 88
rect 98 87 99 88
rect 97 87 98 88
rect 96 87 97 88
rect 95 87 96 88
rect 94 87 95 88
rect 93 87 94 88
rect 92 87 93 88
rect 91 87 92 88
rect 80 87 81 88
rect 79 87 80 88
rect 78 87 79 88
rect 77 87 78 88
rect 76 87 77 88
rect 75 87 76 88
rect 74 87 75 88
rect 73 87 74 88
rect 72 87 73 88
rect 71 87 72 88
rect 70 87 71 88
rect 69 87 70 88
rect 68 87 69 88
rect 67 87 68 88
rect 66 87 67 88
rect 65 87 66 88
rect 64 87 65 88
rect 63 87 64 88
rect 62 87 63 88
rect 61 87 62 88
rect 60 87 61 88
rect 59 87 60 88
rect 58 87 59 88
rect 57 87 58 88
rect 56 87 57 88
rect 55 87 56 88
rect 54 87 55 88
rect 53 87 54 88
rect 52 87 53 88
rect 51 87 52 88
rect 50 87 51 88
rect 49 87 50 88
rect 48 87 49 88
rect 47 87 48 88
rect 46 87 47 88
rect 45 87 46 88
rect 44 87 45 88
rect 43 87 44 88
rect 42 87 43 88
rect 41 87 42 88
rect 40 87 41 88
rect 39 87 40 88
rect 38 87 39 88
rect 37 87 38 88
rect 36 87 37 88
rect 29 87 30 88
rect 28 87 29 88
rect 27 87 28 88
rect 26 87 27 88
rect 25 87 26 88
rect 24 87 25 88
rect 23 87 24 88
rect 22 87 23 88
rect 21 87 22 88
rect 20 87 21 88
rect 19 87 20 88
rect 18 87 19 88
rect 17 87 18 88
rect 16 87 17 88
rect 15 87 16 88
rect 14 87 15 88
rect 13 87 14 88
rect 12 87 13 88
rect 195 88 196 89
rect 194 88 195 89
rect 191 88 192 89
rect 165 88 166 89
rect 147 88 148 89
rect 146 88 147 89
rect 145 88 146 89
rect 144 88 145 89
rect 143 88 144 89
rect 142 88 143 89
rect 141 88 142 89
rect 140 88 141 89
rect 139 88 140 89
rect 138 88 139 89
rect 137 88 138 89
rect 136 88 137 89
rect 135 88 136 89
rect 134 88 135 89
rect 133 88 134 89
rect 132 88 133 89
rect 131 88 132 89
rect 130 88 131 89
rect 129 88 130 89
rect 128 88 129 89
rect 127 88 128 89
rect 126 88 127 89
rect 125 88 126 89
rect 124 88 125 89
rect 123 88 124 89
rect 122 88 123 89
rect 121 88 122 89
rect 120 88 121 89
rect 119 88 120 89
rect 118 88 119 89
rect 117 88 118 89
rect 116 88 117 89
rect 115 88 116 89
rect 114 88 115 89
rect 113 88 114 89
rect 112 88 113 89
rect 111 88 112 89
rect 110 88 111 89
rect 106 88 107 89
rect 105 88 106 89
rect 104 88 105 89
rect 103 88 104 89
rect 102 88 103 89
rect 101 88 102 89
rect 100 88 101 89
rect 99 88 100 89
rect 98 88 99 89
rect 97 88 98 89
rect 96 88 97 89
rect 95 88 96 89
rect 94 88 95 89
rect 93 88 94 89
rect 92 88 93 89
rect 91 88 92 89
rect 90 88 91 89
rect 79 88 80 89
rect 78 88 79 89
rect 77 88 78 89
rect 76 88 77 89
rect 75 88 76 89
rect 74 88 75 89
rect 73 88 74 89
rect 72 88 73 89
rect 71 88 72 89
rect 70 88 71 89
rect 69 88 70 89
rect 68 88 69 89
rect 67 88 68 89
rect 66 88 67 89
rect 65 88 66 89
rect 64 88 65 89
rect 63 88 64 89
rect 62 88 63 89
rect 61 88 62 89
rect 60 88 61 89
rect 59 88 60 89
rect 58 88 59 89
rect 57 88 58 89
rect 56 88 57 89
rect 55 88 56 89
rect 54 88 55 89
rect 53 88 54 89
rect 52 88 53 89
rect 51 88 52 89
rect 50 88 51 89
rect 49 88 50 89
rect 48 88 49 89
rect 47 88 48 89
rect 46 88 47 89
rect 45 88 46 89
rect 44 88 45 89
rect 43 88 44 89
rect 42 88 43 89
rect 41 88 42 89
rect 40 88 41 89
rect 39 88 40 89
rect 38 88 39 89
rect 37 88 38 89
rect 36 88 37 89
rect 29 88 30 89
rect 28 88 29 89
rect 27 88 28 89
rect 26 88 27 89
rect 25 88 26 89
rect 24 88 25 89
rect 23 88 24 89
rect 22 88 23 89
rect 21 88 22 89
rect 20 88 21 89
rect 19 88 20 89
rect 18 88 19 89
rect 17 88 18 89
rect 16 88 17 89
rect 15 88 16 89
rect 14 88 15 89
rect 13 88 14 89
rect 12 88 13 89
rect 199 89 200 90
rect 198 89 199 90
rect 195 89 196 90
rect 194 89 195 90
rect 192 89 193 90
rect 191 89 192 90
rect 148 89 149 90
rect 147 89 148 90
rect 146 89 147 90
rect 145 89 146 90
rect 144 89 145 90
rect 143 89 144 90
rect 142 89 143 90
rect 141 89 142 90
rect 140 89 141 90
rect 139 89 140 90
rect 138 89 139 90
rect 137 89 138 90
rect 136 89 137 90
rect 135 89 136 90
rect 134 89 135 90
rect 133 89 134 90
rect 132 89 133 90
rect 131 89 132 90
rect 130 89 131 90
rect 129 89 130 90
rect 128 89 129 90
rect 127 89 128 90
rect 126 89 127 90
rect 125 89 126 90
rect 124 89 125 90
rect 123 89 124 90
rect 122 89 123 90
rect 121 89 122 90
rect 120 89 121 90
rect 119 89 120 90
rect 118 89 119 90
rect 117 89 118 90
rect 116 89 117 90
rect 115 89 116 90
rect 114 89 115 90
rect 113 89 114 90
rect 112 89 113 90
rect 111 89 112 90
rect 110 89 111 90
rect 109 89 110 90
rect 106 89 107 90
rect 105 89 106 90
rect 104 89 105 90
rect 103 89 104 90
rect 102 89 103 90
rect 101 89 102 90
rect 100 89 101 90
rect 99 89 100 90
rect 98 89 99 90
rect 97 89 98 90
rect 96 89 97 90
rect 95 89 96 90
rect 94 89 95 90
rect 93 89 94 90
rect 92 89 93 90
rect 91 89 92 90
rect 90 89 91 90
rect 89 89 90 90
rect 77 89 78 90
rect 76 89 77 90
rect 75 89 76 90
rect 74 89 75 90
rect 73 89 74 90
rect 72 89 73 90
rect 71 89 72 90
rect 70 89 71 90
rect 69 89 70 90
rect 68 89 69 90
rect 67 89 68 90
rect 66 89 67 90
rect 65 89 66 90
rect 64 89 65 90
rect 63 89 64 90
rect 62 89 63 90
rect 61 89 62 90
rect 60 89 61 90
rect 59 89 60 90
rect 58 89 59 90
rect 57 89 58 90
rect 56 89 57 90
rect 55 89 56 90
rect 54 89 55 90
rect 53 89 54 90
rect 52 89 53 90
rect 51 89 52 90
rect 50 89 51 90
rect 49 89 50 90
rect 48 89 49 90
rect 47 89 48 90
rect 46 89 47 90
rect 45 89 46 90
rect 44 89 45 90
rect 43 89 44 90
rect 42 89 43 90
rect 41 89 42 90
rect 40 89 41 90
rect 39 89 40 90
rect 38 89 39 90
rect 37 89 38 90
rect 30 89 31 90
rect 29 89 30 90
rect 28 89 29 90
rect 27 89 28 90
rect 26 89 27 90
rect 25 89 26 90
rect 24 89 25 90
rect 23 89 24 90
rect 22 89 23 90
rect 21 89 22 90
rect 20 89 21 90
rect 19 89 20 90
rect 18 89 19 90
rect 17 89 18 90
rect 16 89 17 90
rect 15 89 16 90
rect 14 89 15 90
rect 13 89 14 90
rect 12 89 13 90
rect 11 89 12 90
rect 198 90 199 91
rect 197 90 198 91
rect 192 90 193 91
rect 175 90 176 91
rect 174 90 175 91
rect 173 90 174 91
rect 172 90 173 91
rect 148 90 149 91
rect 147 90 148 91
rect 146 90 147 91
rect 145 90 146 91
rect 144 90 145 91
rect 143 90 144 91
rect 142 90 143 91
rect 141 90 142 91
rect 140 90 141 91
rect 139 90 140 91
rect 138 90 139 91
rect 137 90 138 91
rect 136 90 137 91
rect 135 90 136 91
rect 134 90 135 91
rect 133 90 134 91
rect 132 90 133 91
rect 131 90 132 91
rect 130 90 131 91
rect 129 90 130 91
rect 128 90 129 91
rect 127 90 128 91
rect 126 90 127 91
rect 125 90 126 91
rect 124 90 125 91
rect 123 90 124 91
rect 122 90 123 91
rect 121 90 122 91
rect 120 90 121 91
rect 119 90 120 91
rect 118 90 119 91
rect 117 90 118 91
rect 116 90 117 91
rect 115 90 116 91
rect 114 90 115 91
rect 113 90 114 91
rect 112 90 113 91
rect 111 90 112 91
rect 110 90 111 91
rect 109 90 110 91
rect 108 90 109 91
rect 107 90 108 91
rect 106 90 107 91
rect 105 90 106 91
rect 104 90 105 91
rect 103 90 104 91
rect 102 90 103 91
rect 101 90 102 91
rect 100 90 101 91
rect 99 90 100 91
rect 98 90 99 91
rect 97 90 98 91
rect 96 90 97 91
rect 95 90 96 91
rect 94 90 95 91
rect 93 90 94 91
rect 92 90 93 91
rect 91 90 92 91
rect 90 90 91 91
rect 89 90 90 91
rect 88 90 89 91
rect 75 90 76 91
rect 74 90 75 91
rect 73 90 74 91
rect 72 90 73 91
rect 71 90 72 91
rect 70 90 71 91
rect 69 90 70 91
rect 68 90 69 91
rect 67 90 68 91
rect 66 90 67 91
rect 65 90 66 91
rect 64 90 65 91
rect 63 90 64 91
rect 62 90 63 91
rect 61 90 62 91
rect 60 90 61 91
rect 59 90 60 91
rect 58 90 59 91
rect 57 90 58 91
rect 56 90 57 91
rect 55 90 56 91
rect 54 90 55 91
rect 53 90 54 91
rect 52 90 53 91
rect 51 90 52 91
rect 50 90 51 91
rect 49 90 50 91
rect 48 90 49 91
rect 47 90 48 91
rect 46 90 47 91
rect 45 90 46 91
rect 44 90 45 91
rect 43 90 44 91
rect 42 90 43 91
rect 41 90 42 91
rect 40 90 41 91
rect 39 90 40 91
rect 38 90 39 91
rect 31 90 32 91
rect 30 90 31 91
rect 29 90 30 91
rect 28 90 29 91
rect 27 90 28 91
rect 26 90 27 91
rect 25 90 26 91
rect 24 90 25 91
rect 23 90 24 91
rect 22 90 23 91
rect 21 90 22 91
rect 20 90 21 91
rect 19 90 20 91
rect 18 90 19 91
rect 17 90 18 91
rect 16 90 17 91
rect 15 90 16 91
rect 14 90 15 91
rect 13 90 14 91
rect 12 90 13 91
rect 11 90 12 91
rect 178 91 179 92
rect 177 91 178 92
rect 176 91 177 92
rect 175 91 176 92
rect 174 91 175 92
rect 173 91 174 92
rect 172 91 173 92
rect 171 91 172 92
rect 170 91 171 92
rect 169 91 170 92
rect 149 91 150 92
rect 148 91 149 92
rect 147 91 148 92
rect 146 91 147 92
rect 145 91 146 92
rect 144 91 145 92
rect 143 91 144 92
rect 142 91 143 92
rect 141 91 142 92
rect 140 91 141 92
rect 139 91 140 92
rect 138 91 139 92
rect 137 91 138 92
rect 136 91 137 92
rect 135 91 136 92
rect 134 91 135 92
rect 133 91 134 92
rect 132 91 133 92
rect 131 91 132 92
rect 130 91 131 92
rect 129 91 130 92
rect 128 91 129 92
rect 127 91 128 92
rect 126 91 127 92
rect 125 91 126 92
rect 124 91 125 92
rect 123 91 124 92
rect 122 91 123 92
rect 121 91 122 92
rect 120 91 121 92
rect 119 91 120 92
rect 118 91 119 92
rect 117 91 118 92
rect 116 91 117 92
rect 115 91 116 92
rect 114 91 115 92
rect 113 91 114 92
rect 112 91 113 92
rect 111 91 112 92
rect 110 91 111 92
rect 109 91 110 92
rect 108 91 109 92
rect 107 91 108 92
rect 106 91 107 92
rect 105 91 106 92
rect 104 91 105 92
rect 103 91 104 92
rect 102 91 103 92
rect 101 91 102 92
rect 100 91 101 92
rect 99 91 100 92
rect 98 91 99 92
rect 97 91 98 92
rect 96 91 97 92
rect 95 91 96 92
rect 94 91 95 92
rect 93 91 94 92
rect 92 91 93 92
rect 91 91 92 92
rect 90 91 91 92
rect 89 91 90 92
rect 88 91 89 92
rect 87 91 88 92
rect 73 91 74 92
rect 72 91 73 92
rect 71 91 72 92
rect 70 91 71 92
rect 69 91 70 92
rect 68 91 69 92
rect 67 91 68 92
rect 66 91 67 92
rect 65 91 66 92
rect 64 91 65 92
rect 63 91 64 92
rect 62 91 63 92
rect 61 91 62 92
rect 60 91 61 92
rect 59 91 60 92
rect 58 91 59 92
rect 57 91 58 92
rect 56 91 57 92
rect 55 91 56 92
rect 54 91 55 92
rect 53 91 54 92
rect 52 91 53 92
rect 51 91 52 92
rect 50 91 51 92
rect 49 91 50 92
rect 48 91 49 92
rect 47 91 48 92
rect 46 91 47 92
rect 45 91 46 92
rect 44 91 45 92
rect 43 91 44 92
rect 42 91 43 92
rect 41 91 42 92
rect 40 91 41 92
rect 31 91 32 92
rect 30 91 31 92
rect 29 91 30 92
rect 28 91 29 92
rect 27 91 28 92
rect 26 91 27 92
rect 25 91 26 92
rect 24 91 25 92
rect 23 91 24 92
rect 22 91 23 92
rect 21 91 22 92
rect 20 91 21 92
rect 19 91 20 92
rect 18 91 19 92
rect 17 91 18 92
rect 16 91 17 92
rect 15 91 16 92
rect 14 91 15 92
rect 13 91 14 92
rect 12 91 13 92
rect 11 91 12 92
rect 179 92 180 93
rect 178 92 179 93
rect 177 92 178 93
rect 176 92 177 93
rect 175 92 176 93
rect 174 92 175 93
rect 173 92 174 93
rect 172 92 173 93
rect 171 92 172 93
rect 170 92 171 93
rect 169 92 170 93
rect 168 92 169 93
rect 149 92 150 93
rect 148 92 149 93
rect 147 92 148 93
rect 146 92 147 93
rect 145 92 146 93
rect 144 92 145 93
rect 143 92 144 93
rect 142 92 143 93
rect 141 92 142 93
rect 140 92 141 93
rect 139 92 140 93
rect 138 92 139 93
rect 137 92 138 93
rect 136 92 137 93
rect 135 92 136 93
rect 134 92 135 93
rect 133 92 134 93
rect 132 92 133 93
rect 131 92 132 93
rect 130 92 131 93
rect 129 92 130 93
rect 128 92 129 93
rect 127 92 128 93
rect 126 92 127 93
rect 125 92 126 93
rect 124 92 125 93
rect 123 92 124 93
rect 122 92 123 93
rect 121 92 122 93
rect 120 92 121 93
rect 119 92 120 93
rect 118 92 119 93
rect 117 92 118 93
rect 116 92 117 93
rect 115 92 116 93
rect 114 92 115 93
rect 113 92 114 93
rect 112 92 113 93
rect 111 92 112 93
rect 110 92 111 93
rect 109 92 110 93
rect 108 92 109 93
rect 107 92 108 93
rect 106 92 107 93
rect 105 92 106 93
rect 104 92 105 93
rect 103 92 104 93
rect 102 92 103 93
rect 101 92 102 93
rect 100 92 101 93
rect 99 92 100 93
rect 98 92 99 93
rect 97 92 98 93
rect 96 92 97 93
rect 95 92 96 93
rect 94 92 95 93
rect 93 92 94 93
rect 92 92 93 93
rect 91 92 92 93
rect 90 92 91 93
rect 89 92 90 93
rect 88 92 89 93
rect 87 92 88 93
rect 86 92 87 93
rect 85 92 86 93
rect 70 92 71 93
rect 69 92 70 93
rect 68 92 69 93
rect 67 92 68 93
rect 66 92 67 93
rect 65 92 66 93
rect 64 92 65 93
rect 63 92 64 93
rect 62 92 63 93
rect 61 92 62 93
rect 60 92 61 93
rect 59 92 60 93
rect 58 92 59 93
rect 57 92 58 93
rect 56 92 57 93
rect 55 92 56 93
rect 54 92 55 93
rect 53 92 54 93
rect 52 92 53 93
rect 51 92 52 93
rect 50 92 51 93
rect 49 92 50 93
rect 48 92 49 93
rect 47 92 48 93
rect 46 92 47 93
rect 45 92 46 93
rect 44 92 45 93
rect 43 92 44 93
rect 42 92 43 93
rect 41 92 42 93
rect 32 92 33 93
rect 31 92 32 93
rect 30 92 31 93
rect 29 92 30 93
rect 28 92 29 93
rect 27 92 28 93
rect 26 92 27 93
rect 25 92 26 93
rect 24 92 25 93
rect 23 92 24 93
rect 22 92 23 93
rect 21 92 22 93
rect 20 92 21 93
rect 19 92 20 93
rect 18 92 19 93
rect 17 92 18 93
rect 16 92 17 93
rect 15 92 16 93
rect 14 92 15 93
rect 13 92 14 93
rect 12 92 13 93
rect 11 92 12 93
rect 180 93 181 94
rect 179 93 180 94
rect 178 93 179 94
rect 177 93 178 94
rect 176 93 177 94
rect 175 93 176 94
rect 174 93 175 94
rect 173 93 174 94
rect 172 93 173 94
rect 171 93 172 94
rect 170 93 171 94
rect 169 93 170 94
rect 168 93 169 94
rect 167 93 168 94
rect 150 93 151 94
rect 149 93 150 94
rect 148 93 149 94
rect 147 93 148 94
rect 146 93 147 94
rect 145 93 146 94
rect 144 93 145 94
rect 143 93 144 94
rect 142 93 143 94
rect 141 93 142 94
rect 140 93 141 94
rect 139 93 140 94
rect 138 93 139 94
rect 137 93 138 94
rect 136 93 137 94
rect 135 93 136 94
rect 134 93 135 94
rect 133 93 134 94
rect 132 93 133 94
rect 131 93 132 94
rect 130 93 131 94
rect 129 93 130 94
rect 128 93 129 94
rect 127 93 128 94
rect 126 93 127 94
rect 125 93 126 94
rect 124 93 125 94
rect 123 93 124 94
rect 122 93 123 94
rect 121 93 122 94
rect 120 93 121 94
rect 119 93 120 94
rect 118 93 119 94
rect 117 93 118 94
rect 116 93 117 94
rect 115 93 116 94
rect 114 93 115 94
rect 113 93 114 94
rect 112 93 113 94
rect 111 93 112 94
rect 110 93 111 94
rect 109 93 110 94
rect 108 93 109 94
rect 107 93 108 94
rect 106 93 107 94
rect 105 93 106 94
rect 104 93 105 94
rect 103 93 104 94
rect 102 93 103 94
rect 101 93 102 94
rect 100 93 101 94
rect 99 93 100 94
rect 98 93 99 94
rect 97 93 98 94
rect 96 93 97 94
rect 95 93 96 94
rect 94 93 95 94
rect 93 93 94 94
rect 92 93 93 94
rect 91 93 92 94
rect 90 93 91 94
rect 89 93 90 94
rect 88 93 89 94
rect 87 93 88 94
rect 86 93 87 94
rect 85 93 86 94
rect 84 93 85 94
rect 67 93 68 94
rect 66 93 67 94
rect 65 93 66 94
rect 64 93 65 94
rect 63 93 64 94
rect 62 93 63 94
rect 61 93 62 94
rect 60 93 61 94
rect 59 93 60 94
rect 58 93 59 94
rect 57 93 58 94
rect 56 93 57 94
rect 55 93 56 94
rect 54 93 55 94
rect 53 93 54 94
rect 52 93 53 94
rect 51 93 52 94
rect 50 93 51 94
rect 49 93 50 94
rect 48 93 49 94
rect 47 93 48 94
rect 46 93 47 94
rect 45 93 46 94
rect 44 93 45 94
rect 43 93 44 94
rect 33 93 34 94
rect 32 93 33 94
rect 31 93 32 94
rect 30 93 31 94
rect 29 93 30 94
rect 28 93 29 94
rect 27 93 28 94
rect 26 93 27 94
rect 25 93 26 94
rect 24 93 25 94
rect 23 93 24 94
rect 22 93 23 94
rect 21 93 22 94
rect 20 93 21 94
rect 19 93 20 94
rect 18 93 19 94
rect 17 93 18 94
rect 16 93 17 94
rect 15 93 16 94
rect 14 93 15 94
rect 13 93 14 94
rect 12 93 13 94
rect 11 93 12 94
rect 10 93 11 94
rect 191 94 192 95
rect 181 94 182 95
rect 180 94 181 95
rect 179 94 180 95
rect 178 94 179 95
rect 177 94 178 95
rect 176 94 177 95
rect 175 94 176 95
rect 174 94 175 95
rect 173 94 174 95
rect 172 94 173 95
rect 171 94 172 95
rect 170 94 171 95
rect 169 94 170 95
rect 168 94 169 95
rect 167 94 168 95
rect 166 94 167 95
rect 150 94 151 95
rect 149 94 150 95
rect 148 94 149 95
rect 147 94 148 95
rect 146 94 147 95
rect 145 94 146 95
rect 144 94 145 95
rect 143 94 144 95
rect 142 94 143 95
rect 128 94 129 95
rect 127 94 128 95
rect 126 94 127 95
rect 125 94 126 95
rect 124 94 125 95
rect 123 94 124 95
rect 122 94 123 95
rect 121 94 122 95
rect 120 94 121 95
rect 119 94 120 95
rect 118 94 119 95
rect 117 94 118 95
rect 116 94 117 95
rect 115 94 116 95
rect 114 94 115 95
rect 113 94 114 95
rect 112 94 113 95
rect 111 94 112 95
rect 110 94 111 95
rect 109 94 110 95
rect 108 94 109 95
rect 107 94 108 95
rect 106 94 107 95
rect 105 94 106 95
rect 104 94 105 95
rect 103 94 104 95
rect 102 94 103 95
rect 101 94 102 95
rect 100 94 101 95
rect 99 94 100 95
rect 98 94 99 95
rect 97 94 98 95
rect 96 94 97 95
rect 95 94 96 95
rect 94 94 95 95
rect 93 94 94 95
rect 92 94 93 95
rect 91 94 92 95
rect 90 94 91 95
rect 89 94 90 95
rect 88 94 89 95
rect 87 94 88 95
rect 86 94 87 95
rect 85 94 86 95
rect 84 94 85 95
rect 83 94 84 95
rect 82 94 83 95
rect 66 94 67 95
rect 65 94 66 95
rect 64 94 65 95
rect 63 94 64 95
rect 62 94 63 95
rect 61 94 62 95
rect 60 94 61 95
rect 59 94 60 95
rect 58 94 59 95
rect 57 94 58 95
rect 56 94 57 95
rect 55 94 56 95
rect 54 94 55 95
rect 53 94 54 95
rect 52 94 53 95
rect 51 94 52 95
rect 50 94 51 95
rect 49 94 50 95
rect 48 94 49 95
rect 47 94 48 95
rect 46 94 47 95
rect 34 94 35 95
rect 33 94 34 95
rect 32 94 33 95
rect 31 94 32 95
rect 30 94 31 95
rect 29 94 30 95
rect 28 94 29 95
rect 27 94 28 95
rect 26 94 27 95
rect 25 94 26 95
rect 24 94 25 95
rect 23 94 24 95
rect 22 94 23 95
rect 21 94 22 95
rect 20 94 21 95
rect 19 94 20 95
rect 18 94 19 95
rect 17 94 18 95
rect 16 94 17 95
rect 15 94 16 95
rect 14 94 15 95
rect 13 94 14 95
rect 12 94 13 95
rect 11 94 12 95
rect 10 94 11 95
rect 199 95 200 96
rect 198 95 199 96
rect 197 95 198 96
rect 196 95 197 96
rect 195 95 196 96
rect 194 95 195 96
rect 193 95 194 96
rect 192 95 193 96
rect 191 95 192 96
rect 182 95 183 96
rect 181 95 182 96
rect 180 95 181 96
rect 179 95 180 96
rect 178 95 179 96
rect 177 95 178 96
rect 169 95 170 96
rect 168 95 169 96
rect 167 95 168 96
rect 166 95 167 96
rect 151 95 152 96
rect 150 95 151 96
rect 149 95 150 96
rect 148 95 149 96
rect 147 95 148 96
rect 146 95 147 96
rect 125 95 126 96
rect 124 95 125 96
rect 123 95 124 96
rect 122 95 123 96
rect 121 95 122 96
rect 120 95 121 96
rect 119 95 120 96
rect 118 95 119 96
rect 117 95 118 96
rect 116 95 117 96
rect 115 95 116 96
rect 114 95 115 96
rect 113 95 114 96
rect 112 95 113 96
rect 111 95 112 96
rect 110 95 111 96
rect 109 95 110 96
rect 108 95 109 96
rect 107 95 108 96
rect 106 95 107 96
rect 105 95 106 96
rect 104 95 105 96
rect 103 95 104 96
rect 102 95 103 96
rect 101 95 102 96
rect 100 95 101 96
rect 99 95 100 96
rect 98 95 99 96
rect 97 95 98 96
rect 96 95 97 96
rect 95 95 96 96
rect 94 95 95 96
rect 93 95 94 96
rect 92 95 93 96
rect 91 95 92 96
rect 90 95 91 96
rect 89 95 90 96
rect 88 95 89 96
rect 87 95 88 96
rect 86 95 87 96
rect 85 95 86 96
rect 84 95 85 96
rect 83 95 84 96
rect 82 95 83 96
rect 81 95 82 96
rect 80 95 81 96
rect 79 95 80 96
rect 65 95 66 96
rect 64 95 65 96
rect 63 95 64 96
rect 62 95 63 96
rect 61 95 62 96
rect 60 95 61 96
rect 59 95 60 96
rect 58 95 59 96
rect 57 95 58 96
rect 56 95 57 96
rect 55 95 56 96
rect 54 95 55 96
rect 53 95 54 96
rect 52 95 53 96
rect 51 95 52 96
rect 50 95 51 96
rect 49 95 50 96
rect 48 95 49 96
rect 35 95 36 96
rect 34 95 35 96
rect 33 95 34 96
rect 32 95 33 96
rect 31 95 32 96
rect 30 95 31 96
rect 29 95 30 96
rect 28 95 29 96
rect 27 95 28 96
rect 26 95 27 96
rect 25 95 26 96
rect 24 95 25 96
rect 23 95 24 96
rect 22 95 23 96
rect 21 95 22 96
rect 20 95 21 96
rect 19 95 20 96
rect 18 95 19 96
rect 17 95 18 96
rect 16 95 17 96
rect 15 95 16 96
rect 14 95 15 96
rect 13 95 14 96
rect 12 95 13 96
rect 11 95 12 96
rect 10 95 11 96
rect 199 96 200 97
rect 198 96 199 97
rect 197 96 198 97
rect 196 96 197 97
rect 195 96 196 97
rect 194 96 195 97
rect 193 96 194 97
rect 192 96 193 97
rect 191 96 192 97
rect 182 96 183 97
rect 181 96 182 97
rect 180 96 181 97
rect 179 96 180 97
rect 167 96 168 97
rect 166 96 167 97
rect 165 96 166 97
rect 151 96 152 97
rect 150 96 151 97
rect 149 96 150 97
rect 123 96 124 97
rect 122 96 123 97
rect 121 96 122 97
rect 120 96 121 97
rect 119 96 120 97
rect 118 96 119 97
rect 117 96 118 97
rect 116 96 117 97
rect 115 96 116 97
rect 114 96 115 97
rect 113 96 114 97
rect 112 96 113 97
rect 111 96 112 97
rect 110 96 111 97
rect 109 96 110 97
rect 108 96 109 97
rect 107 96 108 97
rect 106 96 107 97
rect 105 96 106 97
rect 104 96 105 97
rect 103 96 104 97
rect 102 96 103 97
rect 101 96 102 97
rect 100 96 101 97
rect 99 96 100 97
rect 98 96 99 97
rect 97 96 98 97
rect 96 96 97 97
rect 95 96 96 97
rect 94 96 95 97
rect 93 96 94 97
rect 92 96 93 97
rect 91 96 92 97
rect 90 96 91 97
rect 89 96 90 97
rect 88 96 89 97
rect 87 96 88 97
rect 86 96 87 97
rect 85 96 86 97
rect 84 96 85 97
rect 83 96 84 97
rect 82 96 83 97
rect 81 96 82 97
rect 80 96 81 97
rect 79 96 80 97
rect 78 96 79 97
rect 77 96 78 97
rect 65 96 66 97
rect 64 96 65 97
rect 63 96 64 97
rect 62 96 63 97
rect 61 96 62 97
rect 60 96 61 97
rect 59 96 60 97
rect 58 96 59 97
rect 57 96 58 97
rect 56 96 57 97
rect 55 96 56 97
rect 54 96 55 97
rect 53 96 54 97
rect 52 96 53 97
rect 51 96 52 97
rect 50 96 51 97
rect 49 96 50 97
rect 36 96 37 97
rect 35 96 36 97
rect 34 96 35 97
rect 33 96 34 97
rect 32 96 33 97
rect 31 96 32 97
rect 30 96 31 97
rect 29 96 30 97
rect 28 96 29 97
rect 27 96 28 97
rect 26 96 27 97
rect 25 96 26 97
rect 24 96 25 97
rect 23 96 24 97
rect 22 96 23 97
rect 21 96 22 97
rect 20 96 21 97
rect 19 96 20 97
rect 18 96 19 97
rect 17 96 18 97
rect 16 96 17 97
rect 15 96 16 97
rect 14 96 15 97
rect 13 96 14 97
rect 12 96 13 97
rect 11 96 12 97
rect 10 96 11 97
rect 199 97 200 98
rect 195 97 196 98
rect 191 97 192 98
rect 182 97 183 98
rect 181 97 182 98
rect 166 97 167 98
rect 165 97 166 98
rect 151 97 152 98
rect 121 97 122 98
rect 120 97 121 98
rect 119 97 120 98
rect 118 97 119 98
rect 117 97 118 98
rect 116 97 117 98
rect 115 97 116 98
rect 114 97 115 98
rect 113 97 114 98
rect 112 97 113 98
rect 111 97 112 98
rect 110 97 111 98
rect 109 97 110 98
rect 108 97 109 98
rect 107 97 108 98
rect 106 97 107 98
rect 105 97 106 98
rect 104 97 105 98
rect 103 97 104 98
rect 102 97 103 98
rect 101 97 102 98
rect 100 97 101 98
rect 99 97 100 98
rect 98 97 99 98
rect 97 97 98 98
rect 96 97 97 98
rect 95 97 96 98
rect 94 97 95 98
rect 93 97 94 98
rect 92 97 93 98
rect 91 97 92 98
rect 90 97 91 98
rect 89 97 90 98
rect 88 97 89 98
rect 87 97 88 98
rect 86 97 87 98
rect 85 97 86 98
rect 84 97 85 98
rect 83 97 84 98
rect 82 97 83 98
rect 81 97 82 98
rect 80 97 81 98
rect 79 97 80 98
rect 78 97 79 98
rect 77 97 78 98
rect 76 97 77 98
rect 75 97 76 98
rect 65 97 66 98
rect 64 97 65 98
rect 63 97 64 98
rect 62 97 63 98
rect 61 97 62 98
rect 60 97 61 98
rect 59 97 60 98
rect 58 97 59 98
rect 57 97 58 98
rect 56 97 57 98
rect 55 97 56 98
rect 54 97 55 98
rect 53 97 54 98
rect 52 97 53 98
rect 51 97 52 98
rect 38 97 39 98
rect 37 97 38 98
rect 36 97 37 98
rect 35 97 36 98
rect 34 97 35 98
rect 33 97 34 98
rect 32 97 33 98
rect 31 97 32 98
rect 30 97 31 98
rect 29 97 30 98
rect 28 97 29 98
rect 27 97 28 98
rect 26 97 27 98
rect 25 97 26 98
rect 24 97 25 98
rect 23 97 24 98
rect 22 97 23 98
rect 21 97 22 98
rect 20 97 21 98
rect 19 97 20 98
rect 18 97 19 98
rect 17 97 18 98
rect 16 97 17 98
rect 15 97 16 98
rect 14 97 15 98
rect 13 97 14 98
rect 12 97 13 98
rect 11 97 12 98
rect 10 97 11 98
rect 197 98 198 99
rect 196 98 197 99
rect 195 98 196 99
rect 194 98 195 99
rect 191 98 192 99
rect 183 98 184 99
rect 182 98 183 99
rect 181 98 182 99
rect 166 98 167 99
rect 165 98 166 99
rect 119 98 120 99
rect 118 98 119 99
rect 117 98 118 99
rect 116 98 117 99
rect 115 98 116 99
rect 114 98 115 99
rect 113 98 114 99
rect 112 98 113 99
rect 111 98 112 99
rect 110 98 111 99
rect 109 98 110 99
rect 108 98 109 99
rect 107 98 108 99
rect 106 98 107 99
rect 105 98 106 99
rect 104 98 105 99
rect 103 98 104 99
rect 102 98 103 99
rect 101 98 102 99
rect 100 98 101 99
rect 99 98 100 99
rect 98 98 99 99
rect 97 98 98 99
rect 96 98 97 99
rect 95 98 96 99
rect 94 98 95 99
rect 93 98 94 99
rect 92 98 93 99
rect 91 98 92 99
rect 90 98 91 99
rect 89 98 90 99
rect 88 98 89 99
rect 87 98 88 99
rect 86 98 87 99
rect 85 98 86 99
rect 84 98 85 99
rect 83 98 84 99
rect 82 98 83 99
rect 81 98 82 99
rect 80 98 81 99
rect 79 98 80 99
rect 78 98 79 99
rect 77 98 78 99
rect 76 98 77 99
rect 75 98 76 99
rect 74 98 75 99
rect 73 98 74 99
rect 65 98 66 99
rect 64 98 65 99
rect 63 98 64 99
rect 62 98 63 99
rect 61 98 62 99
rect 60 98 61 99
rect 59 98 60 99
rect 58 98 59 99
rect 57 98 58 99
rect 56 98 57 99
rect 55 98 56 99
rect 54 98 55 99
rect 53 98 54 99
rect 52 98 53 99
rect 39 98 40 99
rect 38 98 39 99
rect 37 98 38 99
rect 36 98 37 99
rect 35 98 36 99
rect 34 98 35 99
rect 33 98 34 99
rect 32 98 33 99
rect 31 98 32 99
rect 30 98 31 99
rect 29 98 30 99
rect 28 98 29 99
rect 27 98 28 99
rect 26 98 27 99
rect 25 98 26 99
rect 24 98 25 99
rect 23 98 24 99
rect 22 98 23 99
rect 21 98 22 99
rect 20 98 21 99
rect 19 98 20 99
rect 18 98 19 99
rect 17 98 18 99
rect 16 98 17 99
rect 15 98 16 99
rect 14 98 15 99
rect 13 98 14 99
rect 12 98 13 99
rect 11 98 12 99
rect 10 98 11 99
rect 9 98 10 99
rect 198 99 199 100
rect 197 99 198 100
rect 196 99 197 100
rect 195 99 196 100
rect 194 99 195 100
rect 193 99 194 100
rect 192 99 193 100
rect 191 99 192 100
rect 183 99 184 100
rect 182 99 183 100
rect 165 99 166 100
rect 164 99 165 100
rect 118 99 119 100
rect 117 99 118 100
rect 116 99 117 100
rect 115 99 116 100
rect 114 99 115 100
rect 113 99 114 100
rect 112 99 113 100
rect 111 99 112 100
rect 110 99 111 100
rect 109 99 110 100
rect 108 99 109 100
rect 107 99 108 100
rect 106 99 107 100
rect 105 99 106 100
rect 104 99 105 100
rect 103 99 104 100
rect 102 99 103 100
rect 101 99 102 100
rect 100 99 101 100
rect 99 99 100 100
rect 98 99 99 100
rect 97 99 98 100
rect 96 99 97 100
rect 95 99 96 100
rect 94 99 95 100
rect 93 99 94 100
rect 92 99 93 100
rect 91 99 92 100
rect 90 99 91 100
rect 89 99 90 100
rect 88 99 89 100
rect 87 99 88 100
rect 86 99 87 100
rect 85 99 86 100
rect 84 99 85 100
rect 83 99 84 100
rect 82 99 83 100
rect 81 99 82 100
rect 80 99 81 100
rect 79 99 80 100
rect 78 99 79 100
rect 77 99 78 100
rect 76 99 77 100
rect 75 99 76 100
rect 74 99 75 100
rect 73 99 74 100
rect 72 99 73 100
rect 65 99 66 100
rect 64 99 65 100
rect 63 99 64 100
rect 62 99 63 100
rect 61 99 62 100
rect 60 99 61 100
rect 59 99 60 100
rect 58 99 59 100
rect 57 99 58 100
rect 56 99 57 100
rect 55 99 56 100
rect 54 99 55 100
rect 53 99 54 100
rect 52 99 53 100
rect 41 99 42 100
rect 40 99 41 100
rect 39 99 40 100
rect 38 99 39 100
rect 37 99 38 100
rect 36 99 37 100
rect 35 99 36 100
rect 34 99 35 100
rect 33 99 34 100
rect 32 99 33 100
rect 31 99 32 100
rect 30 99 31 100
rect 29 99 30 100
rect 28 99 29 100
rect 27 99 28 100
rect 26 99 27 100
rect 25 99 26 100
rect 24 99 25 100
rect 23 99 24 100
rect 22 99 23 100
rect 21 99 22 100
rect 20 99 21 100
rect 19 99 20 100
rect 18 99 19 100
rect 17 99 18 100
rect 16 99 17 100
rect 15 99 16 100
rect 14 99 15 100
rect 13 99 14 100
rect 12 99 13 100
rect 11 99 12 100
rect 10 99 11 100
rect 9 99 10 100
rect 199 100 200 101
rect 198 100 199 101
rect 197 100 198 101
rect 194 100 195 101
rect 193 100 194 101
rect 192 100 193 101
rect 191 100 192 101
rect 183 100 184 101
rect 182 100 183 101
rect 174 100 175 101
rect 165 100 166 101
rect 164 100 165 101
rect 117 100 118 101
rect 116 100 117 101
rect 115 100 116 101
rect 114 100 115 101
rect 113 100 114 101
rect 112 100 113 101
rect 111 100 112 101
rect 110 100 111 101
rect 109 100 110 101
rect 108 100 109 101
rect 107 100 108 101
rect 106 100 107 101
rect 105 100 106 101
rect 104 100 105 101
rect 103 100 104 101
rect 102 100 103 101
rect 101 100 102 101
rect 100 100 101 101
rect 99 100 100 101
rect 98 100 99 101
rect 97 100 98 101
rect 96 100 97 101
rect 95 100 96 101
rect 94 100 95 101
rect 93 100 94 101
rect 92 100 93 101
rect 91 100 92 101
rect 90 100 91 101
rect 89 100 90 101
rect 88 100 89 101
rect 87 100 88 101
rect 86 100 87 101
rect 85 100 86 101
rect 84 100 85 101
rect 83 100 84 101
rect 82 100 83 101
rect 81 100 82 101
rect 80 100 81 101
rect 79 100 80 101
rect 78 100 79 101
rect 77 100 78 101
rect 76 100 77 101
rect 75 100 76 101
rect 74 100 75 101
rect 73 100 74 101
rect 65 100 66 101
rect 64 100 65 101
rect 63 100 64 101
rect 62 100 63 101
rect 61 100 62 101
rect 60 100 61 101
rect 59 100 60 101
rect 58 100 59 101
rect 57 100 58 101
rect 56 100 57 101
rect 55 100 56 101
rect 54 100 55 101
rect 53 100 54 101
rect 43 100 44 101
rect 42 100 43 101
rect 41 100 42 101
rect 40 100 41 101
rect 39 100 40 101
rect 38 100 39 101
rect 37 100 38 101
rect 36 100 37 101
rect 35 100 36 101
rect 34 100 35 101
rect 33 100 34 101
rect 32 100 33 101
rect 31 100 32 101
rect 30 100 31 101
rect 29 100 30 101
rect 28 100 29 101
rect 27 100 28 101
rect 26 100 27 101
rect 25 100 26 101
rect 24 100 25 101
rect 23 100 24 101
rect 22 100 23 101
rect 21 100 22 101
rect 20 100 21 101
rect 19 100 20 101
rect 18 100 19 101
rect 17 100 18 101
rect 16 100 17 101
rect 15 100 16 101
rect 14 100 15 101
rect 13 100 14 101
rect 12 100 13 101
rect 11 100 12 101
rect 10 100 11 101
rect 9 100 10 101
rect 199 101 200 102
rect 198 101 199 102
rect 183 101 184 102
rect 182 101 183 102
rect 175 101 176 102
rect 174 101 175 102
rect 165 101 166 102
rect 164 101 165 102
rect 116 101 117 102
rect 115 101 116 102
rect 114 101 115 102
rect 113 101 114 102
rect 112 101 113 102
rect 111 101 112 102
rect 110 101 111 102
rect 109 101 110 102
rect 108 101 109 102
rect 107 101 108 102
rect 106 101 107 102
rect 105 101 106 102
rect 104 101 105 102
rect 103 101 104 102
rect 102 101 103 102
rect 101 101 102 102
rect 100 101 101 102
rect 99 101 100 102
rect 98 101 99 102
rect 97 101 98 102
rect 96 101 97 102
rect 95 101 96 102
rect 94 101 95 102
rect 93 101 94 102
rect 92 101 93 102
rect 91 101 92 102
rect 90 101 91 102
rect 89 101 90 102
rect 88 101 89 102
rect 87 101 88 102
rect 86 101 87 102
rect 85 101 86 102
rect 84 101 85 102
rect 83 101 84 102
rect 82 101 83 102
rect 81 101 82 102
rect 80 101 81 102
rect 79 101 80 102
rect 78 101 79 102
rect 77 101 78 102
rect 76 101 77 102
rect 75 101 76 102
rect 74 101 75 102
rect 65 101 66 102
rect 64 101 65 102
rect 63 101 64 102
rect 62 101 63 102
rect 61 101 62 102
rect 60 101 61 102
rect 59 101 60 102
rect 58 101 59 102
rect 57 101 58 102
rect 56 101 57 102
rect 55 101 56 102
rect 54 101 55 102
rect 45 101 46 102
rect 44 101 45 102
rect 43 101 44 102
rect 42 101 43 102
rect 41 101 42 102
rect 40 101 41 102
rect 39 101 40 102
rect 38 101 39 102
rect 37 101 38 102
rect 36 101 37 102
rect 35 101 36 102
rect 34 101 35 102
rect 33 101 34 102
rect 32 101 33 102
rect 31 101 32 102
rect 30 101 31 102
rect 29 101 30 102
rect 28 101 29 102
rect 27 101 28 102
rect 26 101 27 102
rect 25 101 26 102
rect 24 101 25 102
rect 23 101 24 102
rect 22 101 23 102
rect 21 101 22 102
rect 20 101 21 102
rect 19 101 20 102
rect 18 101 19 102
rect 16 101 17 102
rect 15 101 16 102
rect 14 101 15 102
rect 13 101 14 102
rect 12 101 13 102
rect 11 101 12 102
rect 10 101 11 102
rect 9 101 10 102
rect 183 102 184 103
rect 182 102 183 103
rect 175 102 176 103
rect 174 102 175 103
rect 165 102 166 103
rect 164 102 165 103
rect 115 102 116 103
rect 114 102 115 103
rect 113 102 114 103
rect 112 102 113 103
rect 111 102 112 103
rect 110 102 111 103
rect 109 102 110 103
rect 108 102 109 103
rect 107 102 108 103
rect 106 102 107 103
rect 105 102 106 103
rect 104 102 105 103
rect 103 102 104 103
rect 102 102 103 103
rect 101 102 102 103
rect 100 102 101 103
rect 99 102 100 103
rect 98 102 99 103
rect 97 102 98 103
rect 96 102 97 103
rect 95 102 96 103
rect 94 102 95 103
rect 93 102 94 103
rect 92 102 93 103
rect 91 102 92 103
rect 90 102 91 103
rect 89 102 90 103
rect 88 102 89 103
rect 87 102 88 103
rect 86 102 87 103
rect 85 102 86 103
rect 84 102 85 103
rect 83 102 84 103
rect 82 102 83 103
rect 81 102 82 103
rect 80 102 81 103
rect 79 102 80 103
rect 78 102 79 103
rect 77 102 78 103
rect 76 102 77 103
rect 66 102 67 103
rect 65 102 66 103
rect 64 102 65 103
rect 63 102 64 103
rect 62 102 63 103
rect 61 102 62 103
rect 60 102 61 103
rect 59 102 60 103
rect 58 102 59 103
rect 57 102 58 103
rect 56 102 57 103
rect 55 102 56 103
rect 54 102 55 103
rect 46 102 47 103
rect 45 102 46 103
rect 44 102 45 103
rect 43 102 44 103
rect 42 102 43 103
rect 41 102 42 103
rect 40 102 41 103
rect 39 102 40 103
rect 38 102 39 103
rect 37 102 38 103
rect 36 102 37 103
rect 35 102 36 103
rect 34 102 35 103
rect 33 102 34 103
rect 32 102 33 103
rect 31 102 32 103
rect 30 102 31 103
rect 29 102 30 103
rect 28 102 29 103
rect 27 102 28 103
rect 26 102 27 103
rect 25 102 26 103
rect 24 102 25 103
rect 23 102 24 103
rect 22 102 23 103
rect 21 102 22 103
rect 20 102 21 103
rect 19 102 20 103
rect 18 102 19 103
rect 15 102 16 103
rect 14 102 15 103
rect 13 102 14 103
rect 12 102 13 103
rect 11 102 12 103
rect 10 102 11 103
rect 9 102 10 103
rect 183 103 184 104
rect 182 103 183 104
rect 181 103 182 104
rect 180 103 181 104
rect 179 103 180 104
rect 178 103 179 104
rect 177 103 178 104
rect 176 103 177 104
rect 175 103 176 104
rect 174 103 175 104
rect 166 103 167 104
rect 165 103 166 104
rect 164 103 165 104
rect 133 103 134 104
rect 132 103 133 104
rect 131 103 132 104
rect 130 103 131 104
rect 129 103 130 104
rect 128 103 129 104
rect 127 103 128 104
rect 126 103 127 104
rect 125 103 126 104
rect 124 103 125 104
rect 123 103 124 104
rect 122 103 123 104
rect 121 103 122 104
rect 114 103 115 104
rect 113 103 114 104
rect 112 103 113 104
rect 111 103 112 104
rect 110 103 111 104
rect 109 103 110 104
rect 108 103 109 104
rect 107 103 108 104
rect 106 103 107 104
rect 105 103 106 104
rect 104 103 105 104
rect 103 103 104 104
rect 102 103 103 104
rect 101 103 102 104
rect 100 103 101 104
rect 99 103 100 104
rect 98 103 99 104
rect 97 103 98 104
rect 96 103 97 104
rect 95 103 96 104
rect 94 103 95 104
rect 93 103 94 104
rect 92 103 93 104
rect 91 103 92 104
rect 90 103 91 104
rect 89 103 90 104
rect 88 103 89 104
rect 87 103 88 104
rect 86 103 87 104
rect 85 103 86 104
rect 84 103 85 104
rect 83 103 84 104
rect 82 103 83 104
rect 81 103 82 104
rect 80 103 81 104
rect 79 103 80 104
rect 78 103 79 104
rect 66 103 67 104
rect 65 103 66 104
rect 64 103 65 104
rect 63 103 64 104
rect 62 103 63 104
rect 61 103 62 104
rect 60 103 61 104
rect 59 103 60 104
rect 58 103 59 104
rect 57 103 58 104
rect 56 103 57 104
rect 55 103 56 104
rect 54 103 55 104
rect 47 103 48 104
rect 46 103 47 104
rect 45 103 46 104
rect 44 103 45 104
rect 43 103 44 104
rect 42 103 43 104
rect 41 103 42 104
rect 40 103 41 104
rect 39 103 40 104
rect 38 103 39 104
rect 37 103 38 104
rect 36 103 37 104
rect 35 103 36 104
rect 34 103 35 104
rect 33 103 34 104
rect 32 103 33 104
rect 31 103 32 104
rect 30 103 31 104
rect 29 103 30 104
rect 28 103 29 104
rect 27 103 28 104
rect 26 103 27 104
rect 25 103 26 104
rect 24 103 25 104
rect 23 103 24 104
rect 22 103 23 104
rect 21 103 22 104
rect 20 103 21 104
rect 19 103 20 104
rect 18 103 19 104
rect 15 103 16 104
rect 14 103 15 104
rect 13 103 14 104
rect 12 103 13 104
rect 11 103 12 104
rect 10 103 11 104
rect 9 103 10 104
rect 182 104 183 105
rect 181 104 182 105
rect 180 104 181 105
rect 179 104 180 105
rect 178 104 179 105
rect 177 104 178 105
rect 176 104 177 105
rect 175 104 176 105
rect 174 104 175 105
rect 167 104 168 105
rect 166 104 167 105
rect 165 104 166 105
rect 137 104 138 105
rect 136 104 137 105
rect 135 104 136 105
rect 134 104 135 105
rect 133 104 134 105
rect 132 104 133 105
rect 131 104 132 105
rect 130 104 131 105
rect 129 104 130 105
rect 128 104 129 105
rect 127 104 128 105
rect 126 104 127 105
rect 125 104 126 105
rect 124 104 125 105
rect 123 104 124 105
rect 122 104 123 105
rect 121 104 122 105
rect 120 104 121 105
rect 119 104 120 105
rect 118 104 119 105
rect 117 104 118 105
rect 114 104 115 105
rect 113 104 114 105
rect 112 104 113 105
rect 111 104 112 105
rect 110 104 111 105
rect 109 104 110 105
rect 108 104 109 105
rect 107 104 108 105
rect 106 104 107 105
rect 105 104 106 105
rect 104 104 105 105
rect 103 104 104 105
rect 102 104 103 105
rect 101 104 102 105
rect 100 104 101 105
rect 99 104 100 105
rect 98 104 99 105
rect 97 104 98 105
rect 96 104 97 105
rect 95 104 96 105
rect 94 104 95 105
rect 93 104 94 105
rect 92 104 93 105
rect 91 104 92 105
rect 90 104 91 105
rect 89 104 90 105
rect 88 104 89 105
rect 87 104 88 105
rect 86 104 87 105
rect 85 104 86 105
rect 84 104 85 105
rect 83 104 84 105
rect 82 104 83 105
rect 81 104 82 105
rect 80 104 81 105
rect 67 104 68 105
rect 66 104 67 105
rect 65 104 66 105
rect 64 104 65 105
rect 63 104 64 105
rect 62 104 63 105
rect 61 104 62 105
rect 60 104 61 105
rect 59 104 60 105
rect 58 104 59 105
rect 57 104 58 105
rect 56 104 57 105
rect 55 104 56 105
rect 48 104 49 105
rect 47 104 48 105
rect 46 104 47 105
rect 45 104 46 105
rect 44 104 45 105
rect 43 104 44 105
rect 42 104 43 105
rect 41 104 42 105
rect 40 104 41 105
rect 39 104 40 105
rect 38 104 39 105
rect 37 104 38 105
rect 36 104 37 105
rect 35 104 36 105
rect 34 104 35 105
rect 33 104 34 105
rect 32 104 33 105
rect 31 104 32 105
rect 30 104 31 105
rect 29 104 30 105
rect 28 104 29 105
rect 27 104 28 105
rect 26 104 27 105
rect 25 104 26 105
rect 24 104 25 105
rect 23 104 24 105
rect 22 104 23 105
rect 21 104 22 105
rect 20 104 21 105
rect 19 104 20 105
rect 15 104 16 105
rect 14 104 15 105
rect 13 104 14 105
rect 12 104 13 105
rect 11 104 12 105
rect 10 104 11 105
rect 9 104 10 105
rect 8 104 9 105
rect 198 105 199 106
rect 197 105 198 106
rect 193 105 194 106
rect 192 105 193 106
rect 182 105 183 106
rect 181 105 182 106
rect 180 105 181 106
rect 179 105 180 106
rect 178 105 179 106
rect 177 105 178 106
rect 176 105 177 106
rect 175 105 176 106
rect 174 105 175 106
rect 168 105 169 106
rect 167 105 168 106
rect 166 105 167 106
rect 165 105 166 106
rect 137 105 138 106
rect 136 105 137 106
rect 135 105 136 106
rect 134 105 135 106
rect 133 105 134 106
rect 132 105 133 106
rect 131 105 132 106
rect 130 105 131 106
rect 129 105 130 106
rect 128 105 129 106
rect 127 105 128 106
rect 126 105 127 106
rect 125 105 126 106
rect 124 105 125 106
rect 123 105 124 106
rect 122 105 123 106
rect 121 105 122 106
rect 120 105 121 106
rect 119 105 120 106
rect 118 105 119 106
rect 117 105 118 106
rect 116 105 117 106
rect 115 105 116 106
rect 113 105 114 106
rect 112 105 113 106
rect 111 105 112 106
rect 110 105 111 106
rect 109 105 110 106
rect 108 105 109 106
rect 107 105 108 106
rect 106 105 107 106
rect 105 105 106 106
rect 104 105 105 106
rect 103 105 104 106
rect 102 105 103 106
rect 101 105 102 106
rect 100 105 101 106
rect 95 105 96 106
rect 94 105 95 106
rect 93 105 94 106
rect 92 105 93 106
rect 91 105 92 106
rect 90 105 91 106
rect 89 105 90 106
rect 88 105 89 106
rect 87 105 88 106
rect 86 105 87 106
rect 85 105 86 106
rect 84 105 85 106
rect 83 105 84 106
rect 68 105 69 106
rect 67 105 68 106
rect 66 105 67 106
rect 65 105 66 106
rect 64 105 65 106
rect 63 105 64 106
rect 62 105 63 106
rect 61 105 62 106
rect 60 105 61 106
rect 59 105 60 106
rect 58 105 59 106
rect 57 105 58 106
rect 56 105 57 106
rect 55 105 56 106
rect 49 105 50 106
rect 48 105 49 106
rect 47 105 48 106
rect 46 105 47 106
rect 45 105 46 106
rect 44 105 45 106
rect 43 105 44 106
rect 42 105 43 106
rect 41 105 42 106
rect 40 105 41 106
rect 39 105 40 106
rect 38 105 39 106
rect 37 105 38 106
rect 36 105 37 106
rect 35 105 36 106
rect 34 105 35 106
rect 33 105 34 106
rect 32 105 33 106
rect 31 105 32 106
rect 30 105 31 106
rect 29 105 30 106
rect 28 105 29 106
rect 27 105 28 106
rect 26 105 27 106
rect 25 105 26 106
rect 24 105 25 106
rect 23 105 24 106
rect 22 105 23 106
rect 21 105 22 106
rect 20 105 21 106
rect 19 105 20 106
rect 15 105 16 106
rect 14 105 15 106
rect 13 105 14 106
rect 12 105 13 106
rect 11 105 12 106
rect 10 105 11 106
rect 9 105 10 106
rect 199 106 200 107
rect 198 106 199 107
rect 194 106 195 107
rect 193 106 194 107
rect 192 106 193 107
rect 191 106 192 107
rect 182 106 183 107
rect 181 106 182 107
rect 180 106 181 107
rect 179 106 180 107
rect 178 106 179 107
rect 177 106 178 107
rect 176 106 177 107
rect 175 106 176 107
rect 174 106 175 107
rect 169 106 170 107
rect 168 106 169 107
rect 167 106 168 107
rect 166 106 167 107
rect 165 106 166 107
rect 135 106 136 107
rect 134 106 135 107
rect 133 106 134 107
rect 132 106 133 107
rect 131 106 132 107
rect 130 106 131 107
rect 129 106 130 107
rect 128 106 129 107
rect 127 106 128 107
rect 126 106 127 107
rect 125 106 126 107
rect 124 106 125 107
rect 123 106 124 107
rect 122 106 123 107
rect 121 106 122 107
rect 120 106 121 107
rect 119 106 120 107
rect 118 106 119 107
rect 117 106 118 107
rect 116 106 117 107
rect 115 106 116 107
rect 114 106 115 107
rect 113 106 114 107
rect 112 106 113 107
rect 111 106 112 107
rect 110 106 111 107
rect 109 106 110 107
rect 108 106 109 107
rect 107 106 108 107
rect 106 106 107 107
rect 105 106 106 107
rect 104 106 105 107
rect 103 106 104 107
rect 102 106 103 107
rect 101 106 102 107
rect 100 106 101 107
rect 69 106 70 107
rect 68 106 69 107
rect 67 106 68 107
rect 66 106 67 107
rect 65 106 66 107
rect 64 106 65 107
rect 63 106 64 107
rect 62 106 63 107
rect 61 106 62 107
rect 60 106 61 107
rect 59 106 60 107
rect 58 106 59 107
rect 57 106 58 107
rect 56 106 57 107
rect 55 106 56 107
rect 49 106 50 107
rect 48 106 49 107
rect 47 106 48 107
rect 46 106 47 107
rect 45 106 46 107
rect 44 106 45 107
rect 43 106 44 107
rect 42 106 43 107
rect 41 106 42 107
rect 40 106 41 107
rect 39 106 40 107
rect 38 106 39 107
rect 37 106 38 107
rect 36 106 37 107
rect 35 106 36 107
rect 34 106 35 107
rect 33 106 34 107
rect 32 106 33 107
rect 31 106 32 107
rect 30 106 31 107
rect 29 106 30 107
rect 28 106 29 107
rect 27 106 28 107
rect 26 106 27 107
rect 25 106 26 107
rect 24 106 25 107
rect 23 106 24 107
rect 22 106 23 107
rect 21 106 22 107
rect 20 106 21 107
rect 19 106 20 107
rect 15 106 16 107
rect 14 106 15 107
rect 13 106 14 107
rect 12 106 13 107
rect 11 106 12 107
rect 10 106 11 107
rect 9 106 10 107
rect 8 106 9 107
rect 199 107 200 108
rect 195 107 196 108
rect 194 107 195 108
rect 193 107 194 108
rect 191 107 192 108
rect 190 107 191 108
rect 175 107 176 108
rect 174 107 175 108
rect 134 107 135 108
rect 133 107 134 108
rect 132 107 133 108
rect 131 107 132 108
rect 130 107 131 108
rect 129 107 130 108
rect 128 107 129 108
rect 127 107 128 108
rect 126 107 127 108
rect 125 107 126 108
rect 124 107 125 108
rect 123 107 124 108
rect 122 107 123 108
rect 121 107 122 108
rect 120 107 121 108
rect 119 107 120 108
rect 118 107 119 108
rect 117 107 118 108
rect 116 107 117 108
rect 115 107 116 108
rect 114 107 115 108
rect 113 107 114 108
rect 112 107 113 108
rect 111 107 112 108
rect 110 107 111 108
rect 109 107 110 108
rect 108 107 109 108
rect 107 107 108 108
rect 106 107 107 108
rect 105 107 106 108
rect 104 107 105 108
rect 103 107 104 108
rect 102 107 103 108
rect 101 107 102 108
rect 100 107 101 108
rect 99 107 100 108
rect 70 107 71 108
rect 69 107 70 108
rect 68 107 69 108
rect 67 107 68 108
rect 66 107 67 108
rect 65 107 66 108
rect 64 107 65 108
rect 63 107 64 108
rect 62 107 63 108
rect 61 107 62 108
rect 60 107 61 108
rect 59 107 60 108
rect 58 107 59 108
rect 57 107 58 108
rect 56 107 57 108
rect 55 107 56 108
rect 50 107 51 108
rect 49 107 50 108
rect 48 107 49 108
rect 47 107 48 108
rect 46 107 47 108
rect 45 107 46 108
rect 44 107 45 108
rect 43 107 44 108
rect 42 107 43 108
rect 41 107 42 108
rect 40 107 41 108
rect 39 107 40 108
rect 38 107 39 108
rect 37 107 38 108
rect 36 107 37 108
rect 35 107 36 108
rect 34 107 35 108
rect 33 107 34 108
rect 32 107 33 108
rect 31 107 32 108
rect 30 107 31 108
rect 29 107 30 108
rect 28 107 29 108
rect 27 107 28 108
rect 26 107 27 108
rect 25 107 26 108
rect 24 107 25 108
rect 23 107 24 108
rect 22 107 23 108
rect 21 107 22 108
rect 20 107 21 108
rect 15 107 16 108
rect 14 107 15 108
rect 13 107 14 108
rect 12 107 13 108
rect 11 107 12 108
rect 10 107 11 108
rect 9 107 10 108
rect 8 107 9 108
rect 199 108 200 109
rect 196 108 197 109
rect 195 108 196 109
rect 194 108 195 109
rect 191 108 192 109
rect 190 108 191 109
rect 175 108 176 109
rect 174 108 175 109
rect 132 108 133 109
rect 131 108 132 109
rect 130 108 131 109
rect 129 108 130 109
rect 128 108 129 109
rect 127 108 128 109
rect 126 108 127 109
rect 125 108 126 109
rect 124 108 125 109
rect 123 108 124 109
rect 122 108 123 109
rect 121 108 122 109
rect 120 108 121 109
rect 119 108 120 109
rect 118 108 119 109
rect 117 108 118 109
rect 116 108 117 109
rect 115 108 116 109
rect 114 108 115 109
rect 113 108 114 109
rect 112 108 113 109
rect 111 108 112 109
rect 110 108 111 109
rect 109 108 110 109
rect 108 108 109 109
rect 107 108 108 109
rect 106 108 107 109
rect 105 108 106 109
rect 104 108 105 109
rect 103 108 104 109
rect 102 108 103 109
rect 101 108 102 109
rect 100 108 101 109
rect 99 108 100 109
rect 71 108 72 109
rect 70 108 71 109
rect 69 108 70 109
rect 68 108 69 109
rect 67 108 68 109
rect 66 108 67 109
rect 65 108 66 109
rect 64 108 65 109
rect 63 108 64 109
rect 62 108 63 109
rect 61 108 62 109
rect 60 108 61 109
rect 59 108 60 109
rect 58 108 59 109
rect 57 108 58 109
rect 56 108 57 109
rect 50 108 51 109
rect 49 108 50 109
rect 48 108 49 109
rect 47 108 48 109
rect 46 108 47 109
rect 45 108 46 109
rect 44 108 45 109
rect 43 108 44 109
rect 42 108 43 109
rect 41 108 42 109
rect 40 108 41 109
rect 39 108 40 109
rect 38 108 39 109
rect 37 108 38 109
rect 36 108 37 109
rect 35 108 36 109
rect 34 108 35 109
rect 33 108 34 109
rect 32 108 33 109
rect 31 108 32 109
rect 30 108 31 109
rect 29 108 30 109
rect 28 108 29 109
rect 27 108 28 109
rect 26 108 27 109
rect 25 108 26 109
rect 24 108 25 109
rect 23 108 24 109
rect 22 108 23 109
rect 21 108 22 109
rect 20 108 21 109
rect 15 108 16 109
rect 14 108 15 109
rect 13 108 14 109
rect 12 108 13 109
rect 11 108 12 109
rect 10 108 11 109
rect 9 108 10 109
rect 8 108 9 109
rect 198 109 199 110
rect 197 109 198 110
rect 196 109 197 110
rect 195 109 196 110
rect 194 109 195 110
rect 191 109 192 110
rect 190 109 191 110
rect 131 109 132 110
rect 130 109 131 110
rect 129 109 130 110
rect 128 109 129 110
rect 127 109 128 110
rect 126 109 127 110
rect 125 109 126 110
rect 124 109 125 110
rect 123 109 124 110
rect 122 109 123 110
rect 121 109 122 110
rect 120 109 121 110
rect 119 109 120 110
rect 118 109 119 110
rect 117 109 118 110
rect 116 109 117 110
rect 115 109 116 110
rect 114 109 115 110
rect 113 109 114 110
rect 112 109 113 110
rect 111 109 112 110
rect 110 109 111 110
rect 109 109 110 110
rect 108 109 109 110
rect 107 109 108 110
rect 106 109 107 110
rect 105 109 106 110
rect 104 109 105 110
rect 103 109 104 110
rect 102 109 103 110
rect 101 109 102 110
rect 100 109 101 110
rect 99 109 100 110
rect 73 109 74 110
rect 72 109 73 110
rect 71 109 72 110
rect 70 109 71 110
rect 69 109 70 110
rect 68 109 69 110
rect 67 109 68 110
rect 66 109 67 110
rect 65 109 66 110
rect 64 109 65 110
rect 63 109 64 110
rect 62 109 63 110
rect 61 109 62 110
rect 60 109 61 110
rect 59 109 60 110
rect 58 109 59 110
rect 57 109 58 110
rect 56 109 57 110
rect 50 109 51 110
rect 49 109 50 110
rect 48 109 49 110
rect 47 109 48 110
rect 46 109 47 110
rect 45 109 46 110
rect 44 109 45 110
rect 43 109 44 110
rect 42 109 43 110
rect 41 109 42 110
rect 40 109 41 110
rect 39 109 40 110
rect 38 109 39 110
rect 37 109 38 110
rect 36 109 37 110
rect 35 109 36 110
rect 34 109 35 110
rect 33 109 34 110
rect 32 109 33 110
rect 31 109 32 110
rect 29 109 30 110
rect 28 109 29 110
rect 27 109 28 110
rect 26 109 27 110
rect 25 109 26 110
rect 24 109 25 110
rect 23 109 24 110
rect 22 109 23 110
rect 21 109 22 110
rect 20 109 21 110
rect 16 109 17 110
rect 15 109 16 110
rect 14 109 15 110
rect 13 109 14 110
rect 12 109 13 110
rect 11 109 12 110
rect 10 109 11 110
rect 9 109 10 110
rect 8 109 9 110
rect 197 110 198 111
rect 196 110 197 111
rect 195 110 196 111
rect 192 110 193 111
rect 191 110 192 111
rect 130 110 131 111
rect 129 110 130 111
rect 128 110 129 111
rect 127 110 128 111
rect 126 110 127 111
rect 125 110 126 111
rect 124 110 125 111
rect 123 110 124 111
rect 122 110 123 111
rect 121 110 122 111
rect 120 110 121 111
rect 119 110 120 111
rect 118 110 119 111
rect 117 110 118 111
rect 116 110 117 111
rect 115 110 116 111
rect 114 110 115 111
rect 113 110 114 111
rect 112 110 113 111
rect 111 110 112 111
rect 110 110 111 111
rect 109 110 110 111
rect 108 110 109 111
rect 107 110 108 111
rect 106 110 107 111
rect 105 110 106 111
rect 104 110 105 111
rect 103 110 104 111
rect 102 110 103 111
rect 101 110 102 111
rect 100 110 101 111
rect 99 110 100 111
rect 75 110 76 111
rect 74 110 75 111
rect 73 110 74 111
rect 72 110 73 111
rect 71 110 72 111
rect 70 110 71 111
rect 69 110 70 111
rect 68 110 69 111
rect 67 110 68 111
rect 66 110 67 111
rect 65 110 66 111
rect 64 110 65 111
rect 63 110 64 111
rect 62 110 63 111
rect 61 110 62 111
rect 60 110 61 111
rect 59 110 60 111
rect 58 110 59 111
rect 57 110 58 111
rect 56 110 57 111
rect 51 110 52 111
rect 50 110 51 111
rect 49 110 50 111
rect 48 110 49 111
rect 47 110 48 111
rect 46 110 47 111
rect 45 110 46 111
rect 44 110 45 111
rect 43 110 44 111
rect 42 110 43 111
rect 41 110 42 111
rect 40 110 41 111
rect 39 110 40 111
rect 38 110 39 111
rect 37 110 38 111
rect 36 110 37 111
rect 35 110 36 111
rect 34 110 35 111
rect 29 110 30 111
rect 28 110 29 111
rect 27 110 28 111
rect 26 110 27 111
rect 25 110 26 111
rect 24 110 25 111
rect 23 110 24 111
rect 22 110 23 111
rect 21 110 22 111
rect 16 110 17 111
rect 15 110 16 111
rect 14 110 15 111
rect 13 110 14 111
rect 12 110 13 111
rect 11 110 12 111
rect 10 110 11 111
rect 9 110 10 111
rect 8 110 9 111
rect 129 111 130 112
rect 128 111 129 112
rect 127 111 128 112
rect 126 111 127 112
rect 125 111 126 112
rect 124 111 125 112
rect 123 111 124 112
rect 122 111 123 112
rect 121 111 122 112
rect 120 111 121 112
rect 119 111 120 112
rect 118 111 119 112
rect 117 111 118 112
rect 116 111 117 112
rect 115 111 116 112
rect 114 111 115 112
rect 113 111 114 112
rect 112 111 113 112
rect 111 111 112 112
rect 110 111 111 112
rect 109 111 110 112
rect 108 111 109 112
rect 107 111 108 112
rect 106 111 107 112
rect 105 111 106 112
rect 104 111 105 112
rect 103 111 104 112
rect 102 111 103 112
rect 101 111 102 112
rect 100 111 101 112
rect 99 111 100 112
rect 98 111 99 112
rect 79 111 80 112
rect 78 111 79 112
rect 77 111 78 112
rect 76 111 77 112
rect 75 111 76 112
rect 74 111 75 112
rect 73 111 74 112
rect 72 111 73 112
rect 71 111 72 112
rect 70 111 71 112
rect 69 111 70 112
rect 68 111 69 112
rect 67 111 68 112
rect 66 111 67 112
rect 65 111 66 112
rect 64 111 65 112
rect 63 111 64 112
rect 62 111 63 112
rect 61 111 62 112
rect 60 111 61 112
rect 59 111 60 112
rect 58 111 59 112
rect 57 111 58 112
rect 56 111 57 112
rect 51 111 52 112
rect 50 111 51 112
rect 49 111 50 112
rect 48 111 49 112
rect 47 111 48 112
rect 46 111 47 112
rect 45 111 46 112
rect 44 111 45 112
rect 43 111 44 112
rect 42 111 43 112
rect 41 111 42 112
rect 40 111 41 112
rect 39 111 40 112
rect 38 111 39 112
rect 37 111 38 112
rect 36 111 37 112
rect 35 111 36 112
rect 29 111 30 112
rect 28 111 29 112
rect 27 111 28 112
rect 26 111 27 112
rect 25 111 26 112
rect 24 111 25 112
rect 23 111 24 112
rect 22 111 23 112
rect 21 111 22 112
rect 16 111 17 112
rect 15 111 16 112
rect 14 111 15 112
rect 13 111 14 112
rect 12 111 13 112
rect 11 111 12 112
rect 10 111 11 112
rect 9 111 10 112
rect 8 111 9 112
rect 128 112 129 113
rect 127 112 128 113
rect 126 112 127 113
rect 125 112 126 113
rect 124 112 125 113
rect 123 112 124 113
rect 122 112 123 113
rect 121 112 122 113
rect 120 112 121 113
rect 119 112 120 113
rect 118 112 119 113
rect 117 112 118 113
rect 116 112 117 113
rect 115 112 116 113
rect 114 112 115 113
rect 113 112 114 113
rect 112 112 113 113
rect 111 112 112 113
rect 110 112 111 113
rect 109 112 110 113
rect 108 112 109 113
rect 107 112 108 113
rect 106 112 107 113
rect 105 112 106 113
rect 104 112 105 113
rect 103 112 104 113
rect 102 112 103 113
rect 101 112 102 113
rect 100 112 101 113
rect 99 112 100 113
rect 98 112 99 113
rect 89 112 90 113
rect 88 112 89 113
rect 84 112 85 113
rect 83 112 84 113
rect 82 112 83 113
rect 81 112 82 113
rect 80 112 81 113
rect 79 112 80 113
rect 78 112 79 113
rect 77 112 78 113
rect 76 112 77 113
rect 75 112 76 113
rect 74 112 75 113
rect 73 112 74 113
rect 72 112 73 113
rect 71 112 72 113
rect 70 112 71 113
rect 69 112 70 113
rect 68 112 69 113
rect 67 112 68 113
rect 66 112 67 113
rect 65 112 66 113
rect 64 112 65 113
rect 63 112 64 113
rect 62 112 63 113
rect 61 112 62 113
rect 60 112 61 113
rect 59 112 60 113
rect 58 112 59 113
rect 57 112 58 113
rect 56 112 57 113
rect 51 112 52 113
rect 50 112 51 113
rect 49 112 50 113
rect 48 112 49 113
rect 47 112 48 113
rect 46 112 47 113
rect 45 112 46 113
rect 44 112 45 113
rect 43 112 44 113
rect 42 112 43 113
rect 41 112 42 113
rect 40 112 41 113
rect 39 112 40 113
rect 38 112 39 113
rect 37 112 38 113
rect 36 112 37 113
rect 29 112 30 113
rect 28 112 29 113
rect 27 112 28 113
rect 26 112 27 113
rect 25 112 26 113
rect 24 112 25 113
rect 23 112 24 113
rect 22 112 23 113
rect 21 112 22 113
rect 17 112 18 113
rect 16 112 17 113
rect 15 112 16 113
rect 14 112 15 113
rect 13 112 14 113
rect 12 112 13 113
rect 11 112 12 113
rect 10 112 11 113
rect 9 112 10 113
rect 8 112 9 113
rect 127 113 128 114
rect 126 113 127 114
rect 125 113 126 114
rect 124 113 125 114
rect 123 113 124 114
rect 122 113 123 114
rect 121 113 122 114
rect 120 113 121 114
rect 119 113 120 114
rect 118 113 119 114
rect 117 113 118 114
rect 116 113 117 114
rect 115 113 116 114
rect 114 113 115 114
rect 113 113 114 114
rect 112 113 113 114
rect 111 113 112 114
rect 110 113 111 114
rect 109 113 110 114
rect 108 113 109 114
rect 107 113 108 114
rect 106 113 107 114
rect 105 113 106 114
rect 104 113 105 114
rect 103 113 104 114
rect 102 113 103 114
rect 101 113 102 114
rect 100 113 101 114
rect 99 113 100 114
rect 98 113 99 114
rect 89 113 90 114
rect 88 113 89 114
rect 87 113 88 114
rect 86 113 87 114
rect 85 113 86 114
rect 84 113 85 114
rect 83 113 84 114
rect 82 113 83 114
rect 81 113 82 114
rect 80 113 81 114
rect 79 113 80 114
rect 78 113 79 114
rect 77 113 78 114
rect 76 113 77 114
rect 75 113 76 114
rect 74 113 75 114
rect 73 113 74 114
rect 72 113 73 114
rect 71 113 72 114
rect 70 113 71 114
rect 69 113 70 114
rect 68 113 69 114
rect 67 113 68 114
rect 66 113 67 114
rect 65 113 66 114
rect 64 113 65 114
rect 63 113 64 114
rect 62 113 63 114
rect 61 113 62 114
rect 60 113 61 114
rect 59 113 60 114
rect 58 113 59 114
rect 57 113 58 114
rect 51 113 52 114
rect 50 113 51 114
rect 49 113 50 114
rect 48 113 49 114
rect 47 113 48 114
rect 46 113 47 114
rect 45 113 46 114
rect 44 113 45 114
rect 43 113 44 114
rect 42 113 43 114
rect 41 113 42 114
rect 40 113 41 114
rect 39 113 40 114
rect 38 113 39 114
rect 37 113 38 114
rect 36 113 37 114
rect 30 113 31 114
rect 29 113 30 114
rect 28 113 29 114
rect 27 113 28 114
rect 26 113 27 114
rect 25 113 26 114
rect 24 113 25 114
rect 23 113 24 114
rect 22 113 23 114
rect 21 113 22 114
rect 17 113 18 114
rect 16 113 17 114
rect 15 113 16 114
rect 14 113 15 114
rect 13 113 14 114
rect 12 113 13 114
rect 11 113 12 114
rect 10 113 11 114
rect 9 113 10 114
rect 8 113 9 114
rect 191 114 192 115
rect 126 114 127 115
rect 125 114 126 115
rect 124 114 125 115
rect 123 114 124 115
rect 122 114 123 115
rect 121 114 122 115
rect 120 114 121 115
rect 119 114 120 115
rect 118 114 119 115
rect 117 114 118 115
rect 116 114 117 115
rect 115 114 116 115
rect 114 114 115 115
rect 113 114 114 115
rect 112 114 113 115
rect 111 114 112 115
rect 110 114 111 115
rect 109 114 110 115
rect 108 114 109 115
rect 107 114 108 115
rect 106 114 107 115
rect 105 114 106 115
rect 104 114 105 115
rect 103 114 104 115
rect 102 114 103 115
rect 101 114 102 115
rect 100 114 101 115
rect 99 114 100 115
rect 98 114 99 115
rect 97 114 98 115
rect 89 114 90 115
rect 88 114 89 115
rect 87 114 88 115
rect 86 114 87 115
rect 85 114 86 115
rect 84 114 85 115
rect 83 114 84 115
rect 82 114 83 115
rect 81 114 82 115
rect 80 114 81 115
rect 79 114 80 115
rect 78 114 79 115
rect 77 114 78 115
rect 76 114 77 115
rect 75 114 76 115
rect 74 114 75 115
rect 73 114 74 115
rect 72 114 73 115
rect 71 114 72 115
rect 70 114 71 115
rect 69 114 70 115
rect 68 114 69 115
rect 67 114 68 115
rect 66 114 67 115
rect 65 114 66 115
rect 64 114 65 115
rect 63 114 64 115
rect 62 114 63 115
rect 61 114 62 115
rect 60 114 61 115
rect 59 114 60 115
rect 58 114 59 115
rect 57 114 58 115
rect 51 114 52 115
rect 50 114 51 115
rect 49 114 50 115
rect 48 114 49 115
rect 47 114 48 115
rect 46 114 47 115
rect 45 114 46 115
rect 44 114 45 115
rect 43 114 44 115
rect 42 114 43 115
rect 41 114 42 115
rect 40 114 41 115
rect 39 114 40 115
rect 38 114 39 115
rect 37 114 38 115
rect 30 114 31 115
rect 29 114 30 115
rect 28 114 29 115
rect 27 114 28 115
rect 26 114 27 115
rect 25 114 26 115
rect 24 114 25 115
rect 23 114 24 115
rect 22 114 23 115
rect 17 114 18 115
rect 16 114 17 115
rect 15 114 16 115
rect 14 114 15 115
rect 13 114 14 115
rect 12 114 13 115
rect 11 114 12 115
rect 10 114 11 115
rect 9 114 10 115
rect 8 114 9 115
rect 199 115 200 116
rect 198 115 199 116
rect 197 115 198 116
rect 196 115 197 116
rect 195 115 196 116
rect 194 115 195 116
rect 193 115 194 116
rect 192 115 193 116
rect 191 115 192 116
rect 126 115 127 116
rect 125 115 126 116
rect 124 115 125 116
rect 123 115 124 116
rect 122 115 123 116
rect 121 115 122 116
rect 120 115 121 116
rect 119 115 120 116
rect 118 115 119 116
rect 117 115 118 116
rect 116 115 117 116
rect 115 115 116 116
rect 114 115 115 116
rect 113 115 114 116
rect 112 115 113 116
rect 111 115 112 116
rect 110 115 111 116
rect 109 115 110 116
rect 108 115 109 116
rect 107 115 108 116
rect 106 115 107 116
rect 105 115 106 116
rect 104 115 105 116
rect 103 115 104 116
rect 102 115 103 116
rect 101 115 102 116
rect 100 115 101 116
rect 99 115 100 116
rect 98 115 99 116
rect 97 115 98 116
rect 88 115 89 116
rect 87 115 88 116
rect 86 115 87 116
rect 85 115 86 116
rect 84 115 85 116
rect 83 115 84 116
rect 82 115 83 116
rect 81 115 82 116
rect 80 115 81 116
rect 79 115 80 116
rect 78 115 79 116
rect 77 115 78 116
rect 76 115 77 116
rect 75 115 76 116
rect 74 115 75 116
rect 73 115 74 116
rect 72 115 73 116
rect 71 115 72 116
rect 70 115 71 116
rect 69 115 70 116
rect 68 115 69 116
rect 67 115 68 116
rect 66 115 67 116
rect 65 115 66 116
rect 64 115 65 116
rect 63 115 64 116
rect 62 115 63 116
rect 61 115 62 116
rect 60 115 61 116
rect 59 115 60 116
rect 58 115 59 116
rect 57 115 58 116
rect 51 115 52 116
rect 50 115 51 116
rect 49 115 50 116
rect 48 115 49 116
rect 47 115 48 116
rect 46 115 47 116
rect 45 115 46 116
rect 44 115 45 116
rect 43 115 44 116
rect 42 115 43 116
rect 41 115 42 116
rect 40 115 41 116
rect 39 115 40 116
rect 38 115 39 116
rect 31 115 32 116
rect 30 115 31 116
rect 29 115 30 116
rect 28 115 29 116
rect 27 115 28 116
rect 26 115 27 116
rect 25 115 26 116
rect 24 115 25 116
rect 23 115 24 116
rect 22 115 23 116
rect 17 115 18 116
rect 16 115 17 116
rect 15 115 16 116
rect 14 115 15 116
rect 13 115 14 116
rect 12 115 13 116
rect 11 115 12 116
rect 10 115 11 116
rect 9 115 10 116
rect 8 115 9 116
rect 199 116 200 117
rect 198 116 199 117
rect 197 116 198 117
rect 196 116 197 117
rect 195 116 196 117
rect 194 116 195 117
rect 193 116 194 117
rect 192 116 193 117
rect 191 116 192 117
rect 125 116 126 117
rect 124 116 125 117
rect 123 116 124 117
rect 122 116 123 117
rect 121 116 122 117
rect 120 116 121 117
rect 119 116 120 117
rect 118 116 119 117
rect 117 116 118 117
rect 116 116 117 117
rect 115 116 116 117
rect 114 116 115 117
rect 113 116 114 117
rect 112 116 113 117
rect 111 116 112 117
rect 110 116 111 117
rect 109 116 110 117
rect 108 116 109 117
rect 107 116 108 117
rect 106 116 107 117
rect 105 116 106 117
rect 104 116 105 117
rect 103 116 104 117
rect 102 116 103 117
rect 101 116 102 117
rect 100 116 101 117
rect 99 116 100 117
rect 98 116 99 117
rect 97 116 98 117
rect 88 116 89 117
rect 87 116 88 117
rect 86 116 87 117
rect 85 116 86 117
rect 84 116 85 117
rect 83 116 84 117
rect 82 116 83 117
rect 81 116 82 117
rect 80 116 81 117
rect 79 116 80 117
rect 78 116 79 117
rect 77 116 78 117
rect 76 116 77 117
rect 75 116 76 117
rect 74 116 75 117
rect 73 116 74 117
rect 72 116 73 117
rect 71 116 72 117
rect 70 116 71 117
rect 69 116 70 117
rect 68 116 69 117
rect 67 116 68 117
rect 66 116 67 117
rect 65 116 66 117
rect 64 116 65 117
rect 63 116 64 117
rect 62 116 63 117
rect 61 116 62 117
rect 60 116 61 117
rect 59 116 60 117
rect 58 116 59 117
rect 52 116 53 117
rect 51 116 52 117
rect 50 116 51 117
rect 49 116 50 117
rect 48 116 49 117
rect 47 116 48 117
rect 46 116 47 117
rect 45 116 46 117
rect 44 116 45 117
rect 43 116 44 117
rect 42 116 43 117
rect 41 116 42 117
rect 40 116 41 117
rect 39 116 40 117
rect 38 116 39 117
rect 31 116 32 117
rect 30 116 31 117
rect 29 116 30 117
rect 28 116 29 117
rect 27 116 28 117
rect 26 116 27 117
rect 25 116 26 117
rect 24 116 25 117
rect 23 116 24 117
rect 22 116 23 117
rect 17 116 18 117
rect 16 116 17 117
rect 15 116 16 117
rect 14 116 15 117
rect 13 116 14 117
rect 12 116 13 117
rect 11 116 12 117
rect 10 116 11 117
rect 9 116 10 117
rect 8 116 9 117
rect 198 117 199 118
rect 191 117 192 118
rect 182 117 183 118
rect 165 117 166 118
rect 124 117 125 118
rect 123 117 124 118
rect 122 117 123 118
rect 121 117 122 118
rect 120 117 121 118
rect 119 117 120 118
rect 118 117 119 118
rect 117 117 118 118
rect 116 117 117 118
rect 115 117 116 118
rect 114 117 115 118
rect 113 117 114 118
rect 112 117 113 118
rect 111 117 112 118
rect 110 117 111 118
rect 109 117 110 118
rect 108 117 109 118
rect 107 117 108 118
rect 106 117 107 118
rect 105 117 106 118
rect 104 117 105 118
rect 103 117 104 118
rect 102 117 103 118
rect 101 117 102 118
rect 100 117 101 118
rect 99 117 100 118
rect 98 117 99 118
rect 97 117 98 118
rect 96 117 97 118
rect 87 117 88 118
rect 86 117 87 118
rect 85 117 86 118
rect 84 117 85 118
rect 83 117 84 118
rect 82 117 83 118
rect 81 117 82 118
rect 80 117 81 118
rect 79 117 80 118
rect 78 117 79 118
rect 77 117 78 118
rect 76 117 77 118
rect 75 117 76 118
rect 74 117 75 118
rect 73 117 74 118
rect 72 117 73 118
rect 71 117 72 118
rect 70 117 71 118
rect 69 117 70 118
rect 68 117 69 118
rect 67 117 68 118
rect 66 117 67 118
rect 65 117 66 118
rect 64 117 65 118
rect 63 117 64 118
rect 62 117 63 118
rect 61 117 62 118
rect 60 117 61 118
rect 59 117 60 118
rect 58 117 59 118
rect 52 117 53 118
rect 51 117 52 118
rect 50 117 51 118
rect 49 117 50 118
rect 48 117 49 118
rect 47 117 48 118
rect 46 117 47 118
rect 45 117 46 118
rect 44 117 45 118
rect 43 117 44 118
rect 42 117 43 118
rect 41 117 42 118
rect 40 117 41 118
rect 39 117 40 118
rect 32 117 33 118
rect 31 117 32 118
rect 30 117 31 118
rect 29 117 30 118
rect 28 117 29 118
rect 27 117 28 118
rect 26 117 27 118
rect 25 117 26 118
rect 24 117 25 118
rect 23 117 24 118
rect 22 117 23 118
rect 18 117 19 118
rect 17 117 18 118
rect 16 117 17 118
rect 15 117 16 118
rect 14 117 15 118
rect 13 117 14 118
rect 12 117 13 118
rect 11 117 12 118
rect 10 117 11 118
rect 9 117 10 118
rect 8 117 9 118
rect 182 118 183 119
rect 166 118 167 119
rect 165 118 166 119
rect 123 118 124 119
rect 122 118 123 119
rect 121 118 122 119
rect 120 118 121 119
rect 119 118 120 119
rect 118 118 119 119
rect 117 118 118 119
rect 116 118 117 119
rect 115 118 116 119
rect 114 118 115 119
rect 113 118 114 119
rect 112 118 113 119
rect 111 118 112 119
rect 110 118 111 119
rect 109 118 110 119
rect 108 118 109 119
rect 107 118 108 119
rect 106 118 107 119
rect 105 118 106 119
rect 104 118 105 119
rect 103 118 104 119
rect 102 118 103 119
rect 101 118 102 119
rect 100 118 101 119
rect 99 118 100 119
rect 98 118 99 119
rect 97 118 98 119
rect 96 118 97 119
rect 87 118 88 119
rect 86 118 87 119
rect 85 118 86 119
rect 84 118 85 119
rect 83 118 84 119
rect 82 118 83 119
rect 81 118 82 119
rect 80 118 81 119
rect 79 118 80 119
rect 78 118 79 119
rect 77 118 78 119
rect 76 118 77 119
rect 75 118 76 119
rect 74 118 75 119
rect 73 118 74 119
rect 72 118 73 119
rect 71 118 72 119
rect 70 118 71 119
rect 69 118 70 119
rect 68 118 69 119
rect 67 118 68 119
rect 66 118 67 119
rect 65 118 66 119
rect 64 118 65 119
rect 63 118 64 119
rect 62 118 63 119
rect 61 118 62 119
rect 60 118 61 119
rect 59 118 60 119
rect 58 118 59 119
rect 52 118 53 119
rect 51 118 52 119
rect 50 118 51 119
rect 49 118 50 119
rect 48 118 49 119
rect 47 118 48 119
rect 46 118 47 119
rect 45 118 46 119
rect 44 118 45 119
rect 43 118 44 119
rect 42 118 43 119
rect 41 118 42 119
rect 40 118 41 119
rect 39 118 40 119
rect 32 118 33 119
rect 31 118 32 119
rect 30 118 31 119
rect 29 118 30 119
rect 28 118 29 119
rect 27 118 28 119
rect 26 118 27 119
rect 25 118 26 119
rect 24 118 25 119
rect 23 118 24 119
rect 22 118 23 119
rect 18 118 19 119
rect 17 118 18 119
rect 16 118 17 119
rect 15 118 16 119
rect 14 118 15 119
rect 13 118 14 119
rect 12 118 13 119
rect 11 118 12 119
rect 10 118 11 119
rect 9 118 10 119
rect 8 118 9 119
rect 182 119 183 120
rect 181 119 182 120
rect 180 119 181 120
rect 179 119 180 120
rect 178 119 179 120
rect 177 119 178 120
rect 176 119 177 120
rect 175 119 176 120
rect 174 119 175 120
rect 173 119 174 120
rect 172 119 173 120
rect 171 119 172 120
rect 170 119 171 120
rect 169 119 170 120
rect 168 119 169 120
rect 167 119 168 120
rect 166 119 167 120
rect 165 119 166 120
rect 123 119 124 120
rect 122 119 123 120
rect 121 119 122 120
rect 120 119 121 120
rect 119 119 120 120
rect 118 119 119 120
rect 117 119 118 120
rect 116 119 117 120
rect 115 119 116 120
rect 114 119 115 120
rect 113 119 114 120
rect 112 119 113 120
rect 111 119 112 120
rect 110 119 111 120
rect 109 119 110 120
rect 108 119 109 120
rect 107 119 108 120
rect 106 119 107 120
rect 105 119 106 120
rect 104 119 105 120
rect 103 119 104 120
rect 102 119 103 120
rect 101 119 102 120
rect 100 119 101 120
rect 99 119 100 120
rect 98 119 99 120
rect 97 119 98 120
rect 96 119 97 120
rect 95 119 96 120
rect 86 119 87 120
rect 85 119 86 120
rect 84 119 85 120
rect 83 119 84 120
rect 82 119 83 120
rect 81 119 82 120
rect 80 119 81 120
rect 79 119 80 120
rect 78 119 79 120
rect 77 119 78 120
rect 76 119 77 120
rect 75 119 76 120
rect 74 119 75 120
rect 73 119 74 120
rect 72 119 73 120
rect 71 119 72 120
rect 70 119 71 120
rect 69 119 70 120
rect 68 119 69 120
rect 67 119 68 120
rect 66 119 67 120
rect 65 119 66 120
rect 64 119 65 120
rect 63 119 64 120
rect 62 119 63 120
rect 61 119 62 120
rect 60 119 61 120
rect 59 119 60 120
rect 52 119 53 120
rect 51 119 52 120
rect 50 119 51 120
rect 49 119 50 120
rect 48 119 49 120
rect 47 119 48 120
rect 46 119 47 120
rect 45 119 46 120
rect 44 119 45 120
rect 43 119 44 120
rect 42 119 43 120
rect 41 119 42 120
rect 40 119 41 120
rect 39 119 40 120
rect 32 119 33 120
rect 31 119 32 120
rect 30 119 31 120
rect 29 119 30 120
rect 28 119 29 120
rect 27 119 28 120
rect 26 119 27 120
rect 25 119 26 120
rect 24 119 25 120
rect 23 119 24 120
rect 22 119 23 120
rect 18 119 19 120
rect 17 119 18 120
rect 16 119 17 120
rect 15 119 16 120
rect 14 119 15 120
rect 13 119 14 120
rect 12 119 13 120
rect 11 119 12 120
rect 10 119 11 120
rect 9 119 10 120
rect 8 119 9 120
rect 182 120 183 121
rect 181 120 182 121
rect 180 120 181 121
rect 179 120 180 121
rect 178 120 179 121
rect 177 120 178 121
rect 176 120 177 121
rect 175 120 176 121
rect 174 120 175 121
rect 173 120 174 121
rect 172 120 173 121
rect 171 120 172 121
rect 170 120 171 121
rect 169 120 170 121
rect 168 120 169 121
rect 167 120 168 121
rect 166 120 167 121
rect 165 120 166 121
rect 122 120 123 121
rect 121 120 122 121
rect 120 120 121 121
rect 119 120 120 121
rect 118 120 119 121
rect 117 120 118 121
rect 116 120 117 121
rect 115 120 116 121
rect 114 120 115 121
rect 113 120 114 121
rect 112 120 113 121
rect 111 120 112 121
rect 110 120 111 121
rect 109 120 110 121
rect 108 120 109 121
rect 107 120 108 121
rect 106 120 107 121
rect 105 120 106 121
rect 104 120 105 121
rect 103 120 104 121
rect 102 120 103 121
rect 101 120 102 121
rect 100 120 101 121
rect 99 120 100 121
rect 98 120 99 121
rect 97 120 98 121
rect 96 120 97 121
rect 95 120 96 121
rect 86 120 87 121
rect 85 120 86 121
rect 84 120 85 121
rect 83 120 84 121
rect 82 120 83 121
rect 81 120 82 121
rect 80 120 81 121
rect 79 120 80 121
rect 78 120 79 121
rect 77 120 78 121
rect 76 120 77 121
rect 75 120 76 121
rect 74 120 75 121
rect 73 120 74 121
rect 72 120 73 121
rect 71 120 72 121
rect 70 120 71 121
rect 69 120 70 121
rect 68 120 69 121
rect 67 120 68 121
rect 66 120 67 121
rect 65 120 66 121
rect 64 120 65 121
rect 63 120 64 121
rect 62 120 63 121
rect 61 120 62 121
rect 60 120 61 121
rect 59 120 60 121
rect 53 120 54 121
rect 52 120 53 121
rect 51 120 52 121
rect 50 120 51 121
rect 49 120 50 121
rect 48 120 49 121
rect 47 120 48 121
rect 46 120 47 121
rect 45 120 46 121
rect 44 120 45 121
rect 43 120 44 121
rect 42 120 43 121
rect 41 120 42 121
rect 40 120 41 121
rect 39 120 40 121
rect 33 120 34 121
rect 32 120 33 121
rect 31 120 32 121
rect 30 120 31 121
rect 29 120 30 121
rect 28 120 29 121
rect 27 120 28 121
rect 26 120 27 121
rect 25 120 26 121
rect 24 120 25 121
rect 23 120 24 121
rect 22 120 23 121
rect 18 120 19 121
rect 17 120 18 121
rect 16 120 17 121
rect 15 120 16 121
rect 14 120 15 121
rect 13 120 14 121
rect 12 120 13 121
rect 11 120 12 121
rect 10 120 11 121
rect 9 120 10 121
rect 8 120 9 121
rect 192 121 193 122
rect 191 121 192 122
rect 182 121 183 122
rect 181 121 182 122
rect 180 121 181 122
rect 179 121 180 122
rect 178 121 179 122
rect 177 121 178 122
rect 176 121 177 122
rect 175 121 176 122
rect 174 121 175 122
rect 173 121 174 122
rect 172 121 173 122
rect 171 121 172 122
rect 170 121 171 122
rect 169 121 170 122
rect 168 121 169 122
rect 167 121 168 122
rect 166 121 167 122
rect 165 121 166 122
rect 121 121 122 122
rect 120 121 121 122
rect 119 121 120 122
rect 118 121 119 122
rect 117 121 118 122
rect 116 121 117 122
rect 115 121 116 122
rect 114 121 115 122
rect 113 121 114 122
rect 112 121 113 122
rect 111 121 112 122
rect 110 121 111 122
rect 109 121 110 122
rect 108 121 109 122
rect 107 121 108 122
rect 106 121 107 122
rect 105 121 106 122
rect 104 121 105 122
rect 103 121 104 122
rect 102 121 103 122
rect 101 121 102 122
rect 100 121 101 122
rect 99 121 100 122
rect 98 121 99 122
rect 97 121 98 122
rect 96 121 97 122
rect 95 121 96 122
rect 94 121 95 122
rect 85 121 86 122
rect 84 121 85 122
rect 83 121 84 122
rect 82 121 83 122
rect 81 121 82 122
rect 80 121 81 122
rect 79 121 80 122
rect 78 121 79 122
rect 77 121 78 122
rect 76 121 77 122
rect 75 121 76 122
rect 74 121 75 122
rect 73 121 74 122
rect 72 121 73 122
rect 71 121 72 122
rect 70 121 71 122
rect 69 121 70 122
rect 68 121 69 122
rect 67 121 68 122
rect 66 121 67 122
rect 65 121 66 122
rect 64 121 65 122
rect 63 121 64 122
rect 62 121 63 122
rect 61 121 62 122
rect 60 121 61 122
rect 53 121 54 122
rect 52 121 53 122
rect 51 121 52 122
rect 50 121 51 122
rect 49 121 50 122
rect 48 121 49 122
rect 47 121 48 122
rect 46 121 47 122
rect 45 121 46 122
rect 44 121 45 122
rect 43 121 44 122
rect 42 121 43 122
rect 41 121 42 122
rect 40 121 41 122
rect 33 121 34 122
rect 32 121 33 122
rect 31 121 32 122
rect 30 121 31 122
rect 29 121 30 122
rect 28 121 29 122
rect 27 121 28 122
rect 26 121 27 122
rect 25 121 26 122
rect 24 121 25 122
rect 23 121 24 122
rect 22 121 23 122
rect 18 121 19 122
rect 17 121 18 122
rect 16 121 17 122
rect 15 121 16 122
rect 14 121 15 122
rect 13 121 14 122
rect 12 121 13 122
rect 11 121 12 122
rect 10 121 11 122
rect 9 121 10 122
rect 8 121 9 122
rect 191 122 192 123
rect 182 122 183 123
rect 181 122 182 123
rect 180 122 181 123
rect 179 122 180 123
rect 178 122 179 123
rect 177 122 178 123
rect 176 122 177 123
rect 175 122 176 123
rect 174 122 175 123
rect 173 122 174 123
rect 172 122 173 123
rect 171 122 172 123
rect 170 122 171 123
rect 169 122 170 123
rect 168 122 169 123
rect 167 122 168 123
rect 166 122 167 123
rect 165 122 166 123
rect 120 122 121 123
rect 119 122 120 123
rect 118 122 119 123
rect 117 122 118 123
rect 116 122 117 123
rect 115 122 116 123
rect 114 122 115 123
rect 113 122 114 123
rect 112 122 113 123
rect 111 122 112 123
rect 110 122 111 123
rect 109 122 110 123
rect 108 122 109 123
rect 107 122 108 123
rect 106 122 107 123
rect 105 122 106 123
rect 104 122 105 123
rect 103 122 104 123
rect 102 122 103 123
rect 101 122 102 123
rect 100 122 101 123
rect 99 122 100 123
rect 98 122 99 123
rect 97 122 98 123
rect 96 122 97 123
rect 95 122 96 123
rect 94 122 95 123
rect 84 122 85 123
rect 83 122 84 123
rect 82 122 83 123
rect 81 122 82 123
rect 80 122 81 123
rect 79 122 80 123
rect 78 122 79 123
rect 77 122 78 123
rect 76 122 77 123
rect 75 122 76 123
rect 74 122 75 123
rect 73 122 74 123
rect 72 122 73 123
rect 71 122 72 123
rect 70 122 71 123
rect 69 122 70 123
rect 68 122 69 123
rect 67 122 68 123
rect 66 122 67 123
rect 65 122 66 123
rect 64 122 65 123
rect 63 122 64 123
rect 62 122 63 123
rect 61 122 62 123
rect 60 122 61 123
rect 53 122 54 123
rect 52 122 53 123
rect 51 122 52 123
rect 50 122 51 123
rect 49 122 50 123
rect 48 122 49 123
rect 47 122 48 123
rect 46 122 47 123
rect 45 122 46 123
rect 44 122 45 123
rect 43 122 44 123
rect 42 122 43 123
rect 41 122 42 123
rect 40 122 41 123
rect 33 122 34 123
rect 32 122 33 123
rect 31 122 32 123
rect 30 122 31 123
rect 29 122 30 123
rect 28 122 29 123
rect 27 122 28 123
rect 26 122 27 123
rect 25 122 26 123
rect 24 122 25 123
rect 23 122 24 123
rect 22 122 23 123
rect 19 122 20 123
rect 18 122 19 123
rect 17 122 18 123
rect 16 122 17 123
rect 15 122 16 123
rect 14 122 15 123
rect 13 122 14 123
rect 12 122 13 123
rect 11 122 12 123
rect 10 122 11 123
rect 9 122 10 123
rect 8 122 9 123
rect 182 123 183 124
rect 181 123 182 124
rect 174 123 175 124
rect 173 123 174 124
rect 172 123 173 124
rect 167 123 168 124
rect 166 123 167 124
rect 165 123 166 124
rect 119 123 120 124
rect 118 123 119 124
rect 117 123 118 124
rect 116 123 117 124
rect 115 123 116 124
rect 114 123 115 124
rect 113 123 114 124
rect 112 123 113 124
rect 111 123 112 124
rect 110 123 111 124
rect 109 123 110 124
rect 108 123 109 124
rect 107 123 108 124
rect 106 123 107 124
rect 105 123 106 124
rect 104 123 105 124
rect 103 123 104 124
rect 102 123 103 124
rect 101 123 102 124
rect 100 123 101 124
rect 99 123 100 124
rect 98 123 99 124
rect 97 123 98 124
rect 96 123 97 124
rect 95 123 96 124
rect 94 123 95 124
rect 93 123 94 124
rect 84 123 85 124
rect 83 123 84 124
rect 82 123 83 124
rect 81 123 82 124
rect 80 123 81 124
rect 79 123 80 124
rect 78 123 79 124
rect 77 123 78 124
rect 76 123 77 124
rect 75 123 76 124
rect 74 123 75 124
rect 73 123 74 124
rect 72 123 73 124
rect 71 123 72 124
rect 70 123 71 124
rect 69 123 70 124
rect 68 123 69 124
rect 67 123 68 124
rect 66 123 67 124
rect 65 123 66 124
rect 64 123 65 124
rect 63 123 64 124
rect 62 123 63 124
rect 61 123 62 124
rect 54 123 55 124
rect 53 123 54 124
rect 52 123 53 124
rect 51 123 52 124
rect 50 123 51 124
rect 49 123 50 124
rect 48 123 49 124
rect 47 123 48 124
rect 46 123 47 124
rect 45 123 46 124
rect 44 123 45 124
rect 43 123 44 124
rect 42 123 43 124
rect 41 123 42 124
rect 40 123 41 124
rect 34 123 35 124
rect 33 123 34 124
rect 32 123 33 124
rect 31 123 32 124
rect 30 123 31 124
rect 29 123 30 124
rect 28 123 29 124
rect 27 123 28 124
rect 26 123 27 124
rect 25 123 26 124
rect 24 123 25 124
rect 23 123 24 124
rect 22 123 23 124
rect 19 123 20 124
rect 18 123 19 124
rect 17 123 18 124
rect 16 123 17 124
rect 15 123 16 124
rect 14 123 15 124
rect 13 123 14 124
rect 12 123 13 124
rect 11 123 12 124
rect 10 123 11 124
rect 9 123 10 124
rect 8 123 9 124
rect 199 124 200 125
rect 198 124 199 125
rect 197 124 198 125
rect 196 124 197 125
rect 195 124 196 125
rect 194 124 195 125
rect 193 124 194 125
rect 192 124 193 125
rect 191 124 192 125
rect 182 124 183 125
rect 173 124 174 125
rect 172 124 173 125
rect 165 124 166 125
rect 118 124 119 125
rect 117 124 118 125
rect 116 124 117 125
rect 115 124 116 125
rect 114 124 115 125
rect 113 124 114 125
rect 112 124 113 125
rect 111 124 112 125
rect 110 124 111 125
rect 109 124 110 125
rect 108 124 109 125
rect 107 124 108 125
rect 106 124 107 125
rect 105 124 106 125
rect 104 124 105 125
rect 103 124 104 125
rect 102 124 103 125
rect 101 124 102 125
rect 100 124 101 125
rect 99 124 100 125
rect 98 124 99 125
rect 97 124 98 125
rect 96 124 97 125
rect 95 124 96 125
rect 94 124 95 125
rect 93 124 94 125
rect 92 124 93 125
rect 83 124 84 125
rect 82 124 83 125
rect 81 124 82 125
rect 80 124 81 125
rect 79 124 80 125
rect 78 124 79 125
rect 77 124 78 125
rect 76 124 77 125
rect 75 124 76 125
rect 74 124 75 125
rect 73 124 74 125
rect 72 124 73 125
rect 71 124 72 125
rect 70 124 71 125
rect 69 124 70 125
rect 68 124 69 125
rect 67 124 68 125
rect 66 124 67 125
rect 65 124 66 125
rect 64 124 65 125
rect 63 124 64 125
rect 62 124 63 125
rect 61 124 62 125
rect 54 124 55 125
rect 53 124 54 125
rect 52 124 53 125
rect 51 124 52 125
rect 50 124 51 125
rect 49 124 50 125
rect 48 124 49 125
rect 47 124 48 125
rect 46 124 47 125
rect 45 124 46 125
rect 44 124 45 125
rect 43 124 44 125
rect 42 124 43 125
rect 41 124 42 125
rect 40 124 41 125
rect 34 124 35 125
rect 33 124 34 125
rect 32 124 33 125
rect 31 124 32 125
rect 30 124 31 125
rect 29 124 30 125
rect 28 124 29 125
rect 27 124 28 125
rect 26 124 27 125
rect 25 124 26 125
rect 24 124 25 125
rect 23 124 24 125
rect 19 124 20 125
rect 18 124 19 125
rect 17 124 18 125
rect 16 124 17 125
rect 15 124 16 125
rect 14 124 15 125
rect 13 124 14 125
rect 12 124 13 125
rect 11 124 12 125
rect 10 124 11 125
rect 9 124 10 125
rect 8 124 9 125
rect 198 125 199 126
rect 197 125 198 126
rect 196 125 197 126
rect 195 125 196 126
rect 194 125 195 126
rect 193 125 194 126
rect 192 125 193 126
rect 191 125 192 126
rect 182 125 183 126
rect 173 125 174 126
rect 172 125 173 126
rect 165 125 166 126
rect 117 125 118 126
rect 116 125 117 126
rect 115 125 116 126
rect 114 125 115 126
rect 113 125 114 126
rect 112 125 113 126
rect 111 125 112 126
rect 110 125 111 126
rect 109 125 110 126
rect 108 125 109 126
rect 107 125 108 126
rect 106 125 107 126
rect 105 125 106 126
rect 104 125 105 126
rect 103 125 104 126
rect 102 125 103 126
rect 101 125 102 126
rect 100 125 101 126
rect 99 125 100 126
rect 98 125 99 126
rect 97 125 98 126
rect 96 125 97 126
rect 95 125 96 126
rect 94 125 95 126
rect 93 125 94 126
rect 92 125 93 126
rect 82 125 83 126
rect 81 125 82 126
rect 80 125 81 126
rect 79 125 80 126
rect 78 125 79 126
rect 77 125 78 126
rect 76 125 77 126
rect 75 125 76 126
rect 74 125 75 126
rect 73 125 74 126
rect 72 125 73 126
rect 71 125 72 126
rect 70 125 71 126
rect 69 125 70 126
rect 68 125 69 126
rect 67 125 68 126
rect 66 125 67 126
rect 65 125 66 126
rect 64 125 65 126
rect 63 125 64 126
rect 62 125 63 126
rect 55 125 56 126
rect 54 125 55 126
rect 53 125 54 126
rect 52 125 53 126
rect 51 125 52 126
rect 50 125 51 126
rect 49 125 50 126
rect 48 125 49 126
rect 47 125 48 126
rect 46 125 47 126
rect 45 125 46 126
rect 44 125 45 126
rect 43 125 44 126
rect 42 125 43 126
rect 41 125 42 126
rect 34 125 35 126
rect 33 125 34 126
rect 32 125 33 126
rect 31 125 32 126
rect 30 125 31 126
rect 29 125 30 126
rect 28 125 29 126
rect 27 125 28 126
rect 26 125 27 126
rect 25 125 26 126
rect 24 125 25 126
rect 23 125 24 126
rect 19 125 20 126
rect 18 125 19 126
rect 17 125 18 126
rect 16 125 17 126
rect 15 125 16 126
rect 14 125 15 126
rect 13 125 14 126
rect 12 125 13 126
rect 11 125 12 126
rect 10 125 11 126
rect 9 125 10 126
rect 198 126 199 127
rect 196 126 197 127
rect 195 126 196 127
rect 194 126 195 127
rect 193 126 194 127
rect 191 126 192 127
rect 173 126 174 127
rect 172 126 173 127
rect 116 126 117 127
rect 115 126 116 127
rect 114 126 115 127
rect 113 126 114 127
rect 112 126 113 127
rect 111 126 112 127
rect 110 126 111 127
rect 109 126 110 127
rect 108 126 109 127
rect 107 126 108 127
rect 106 126 107 127
rect 105 126 106 127
rect 104 126 105 127
rect 103 126 104 127
rect 102 126 103 127
rect 101 126 102 127
rect 100 126 101 127
rect 99 126 100 127
rect 98 126 99 127
rect 97 126 98 127
rect 96 126 97 127
rect 95 126 96 127
rect 94 126 95 127
rect 93 126 94 127
rect 92 126 93 127
rect 91 126 92 127
rect 81 126 82 127
rect 80 126 81 127
rect 79 126 80 127
rect 78 126 79 127
rect 77 126 78 127
rect 76 126 77 127
rect 75 126 76 127
rect 74 126 75 127
rect 73 126 74 127
rect 72 126 73 127
rect 71 126 72 127
rect 70 126 71 127
rect 69 126 70 127
rect 68 126 69 127
rect 67 126 68 127
rect 66 126 67 127
rect 65 126 66 127
rect 64 126 65 127
rect 63 126 64 127
rect 55 126 56 127
rect 54 126 55 127
rect 53 126 54 127
rect 52 126 53 127
rect 51 126 52 127
rect 50 126 51 127
rect 49 126 50 127
rect 48 126 49 127
rect 47 126 48 127
rect 46 126 47 127
rect 45 126 46 127
rect 44 126 45 127
rect 43 126 44 127
rect 42 126 43 127
rect 41 126 42 127
rect 34 126 35 127
rect 33 126 34 127
rect 32 126 33 127
rect 31 126 32 127
rect 30 126 31 127
rect 29 126 30 127
rect 28 126 29 127
rect 27 126 28 127
rect 26 126 27 127
rect 25 126 26 127
rect 24 126 25 127
rect 23 126 24 127
rect 19 126 20 127
rect 18 126 19 127
rect 17 126 18 127
rect 16 126 17 127
rect 15 126 16 127
rect 14 126 15 127
rect 13 126 14 127
rect 12 126 13 127
rect 11 126 12 127
rect 10 126 11 127
rect 9 126 10 127
rect 191 127 192 128
rect 173 127 174 128
rect 172 127 173 128
rect 115 127 116 128
rect 114 127 115 128
rect 113 127 114 128
rect 112 127 113 128
rect 111 127 112 128
rect 110 127 111 128
rect 109 127 110 128
rect 108 127 109 128
rect 107 127 108 128
rect 106 127 107 128
rect 105 127 106 128
rect 104 127 105 128
rect 103 127 104 128
rect 102 127 103 128
rect 101 127 102 128
rect 100 127 101 128
rect 99 127 100 128
rect 98 127 99 128
rect 97 127 98 128
rect 96 127 97 128
rect 95 127 96 128
rect 94 127 95 128
rect 93 127 94 128
rect 92 127 93 128
rect 91 127 92 128
rect 90 127 91 128
rect 80 127 81 128
rect 79 127 80 128
rect 78 127 79 128
rect 77 127 78 128
rect 76 127 77 128
rect 75 127 76 128
rect 74 127 75 128
rect 73 127 74 128
rect 72 127 73 128
rect 71 127 72 128
rect 70 127 71 128
rect 69 127 70 128
rect 68 127 69 128
rect 67 127 68 128
rect 66 127 67 128
rect 65 127 66 128
rect 64 127 65 128
rect 55 127 56 128
rect 54 127 55 128
rect 53 127 54 128
rect 52 127 53 128
rect 51 127 52 128
rect 50 127 51 128
rect 49 127 50 128
rect 48 127 49 128
rect 47 127 48 128
rect 46 127 47 128
rect 45 127 46 128
rect 44 127 45 128
rect 43 127 44 128
rect 42 127 43 128
rect 41 127 42 128
rect 35 127 36 128
rect 34 127 35 128
rect 33 127 34 128
rect 32 127 33 128
rect 31 127 32 128
rect 30 127 31 128
rect 29 127 30 128
rect 28 127 29 128
rect 27 127 28 128
rect 26 127 27 128
rect 25 127 26 128
rect 24 127 25 128
rect 23 127 24 128
rect 19 127 20 128
rect 18 127 19 128
rect 17 127 18 128
rect 16 127 17 128
rect 15 127 16 128
rect 14 127 15 128
rect 13 127 14 128
rect 12 127 13 128
rect 11 127 12 128
rect 10 127 11 128
rect 9 127 10 128
rect 192 128 193 129
rect 191 128 192 129
rect 190 128 191 129
rect 182 128 183 129
rect 173 128 174 129
rect 172 128 173 129
rect 165 128 166 129
rect 113 128 114 129
rect 112 128 113 129
rect 111 128 112 129
rect 110 128 111 129
rect 109 128 110 129
rect 108 128 109 129
rect 107 128 108 129
rect 106 128 107 129
rect 105 128 106 129
rect 104 128 105 129
rect 103 128 104 129
rect 102 128 103 129
rect 101 128 102 129
rect 100 128 101 129
rect 99 128 100 129
rect 98 128 99 129
rect 97 128 98 129
rect 96 128 97 129
rect 95 128 96 129
rect 94 128 95 129
rect 93 128 94 129
rect 92 128 93 129
rect 91 128 92 129
rect 90 128 91 129
rect 78 128 79 129
rect 77 128 78 129
rect 76 128 77 129
rect 75 128 76 129
rect 74 128 75 129
rect 73 128 74 129
rect 72 128 73 129
rect 71 128 72 129
rect 70 128 71 129
rect 69 128 70 129
rect 68 128 69 129
rect 67 128 68 129
rect 66 128 67 129
rect 56 128 57 129
rect 55 128 56 129
rect 54 128 55 129
rect 53 128 54 129
rect 52 128 53 129
rect 51 128 52 129
rect 50 128 51 129
rect 49 128 50 129
rect 48 128 49 129
rect 47 128 48 129
rect 46 128 47 129
rect 45 128 46 129
rect 44 128 45 129
rect 43 128 44 129
rect 42 128 43 129
rect 41 128 42 129
rect 35 128 36 129
rect 34 128 35 129
rect 33 128 34 129
rect 32 128 33 129
rect 31 128 32 129
rect 30 128 31 129
rect 29 128 30 129
rect 28 128 29 129
rect 27 128 28 129
rect 26 128 27 129
rect 25 128 26 129
rect 24 128 25 129
rect 19 128 20 129
rect 18 128 19 129
rect 17 128 18 129
rect 16 128 17 129
rect 15 128 16 129
rect 14 128 15 129
rect 13 128 14 129
rect 12 128 13 129
rect 11 128 12 129
rect 10 128 11 129
rect 182 129 183 130
rect 173 129 174 130
rect 172 129 173 130
rect 165 129 166 130
rect 112 129 113 130
rect 111 129 112 130
rect 110 129 111 130
rect 109 129 110 130
rect 108 129 109 130
rect 107 129 108 130
rect 106 129 107 130
rect 105 129 106 130
rect 104 129 105 130
rect 103 129 104 130
rect 102 129 103 130
rect 101 129 102 130
rect 100 129 101 130
rect 99 129 100 130
rect 98 129 99 130
rect 97 129 98 130
rect 96 129 97 130
rect 95 129 96 130
rect 94 129 95 130
rect 93 129 94 130
rect 92 129 93 130
rect 91 129 92 130
rect 90 129 91 130
rect 89 129 90 130
rect 77 129 78 130
rect 76 129 77 130
rect 75 129 76 130
rect 74 129 75 130
rect 73 129 74 130
rect 72 129 73 130
rect 71 129 72 130
rect 70 129 71 130
rect 69 129 70 130
rect 68 129 69 130
rect 56 129 57 130
rect 55 129 56 130
rect 54 129 55 130
rect 53 129 54 130
rect 52 129 53 130
rect 51 129 52 130
rect 50 129 51 130
rect 49 129 50 130
rect 48 129 49 130
rect 47 129 48 130
rect 46 129 47 130
rect 45 129 46 130
rect 44 129 45 130
rect 43 129 44 130
rect 42 129 43 130
rect 35 129 36 130
rect 34 129 35 130
rect 33 129 34 130
rect 32 129 33 130
rect 31 129 32 130
rect 30 129 31 130
rect 29 129 30 130
rect 28 129 29 130
rect 27 129 28 130
rect 26 129 27 130
rect 25 129 26 130
rect 24 129 25 130
rect 19 129 20 130
rect 18 129 19 130
rect 17 129 18 130
rect 16 129 17 130
rect 15 129 16 130
rect 14 129 15 130
rect 13 129 14 130
rect 12 129 13 130
rect 11 129 12 130
rect 10 129 11 130
rect 182 130 183 131
rect 181 130 182 131
rect 174 130 175 131
rect 173 130 174 131
rect 172 130 173 131
rect 166 130 167 131
rect 165 130 166 131
rect 111 130 112 131
rect 110 130 111 131
rect 109 130 110 131
rect 108 130 109 131
rect 107 130 108 131
rect 106 130 107 131
rect 105 130 106 131
rect 104 130 105 131
rect 103 130 104 131
rect 102 130 103 131
rect 101 130 102 131
rect 100 130 101 131
rect 99 130 100 131
rect 98 130 99 131
rect 97 130 98 131
rect 96 130 97 131
rect 95 130 96 131
rect 94 130 95 131
rect 93 130 94 131
rect 92 130 93 131
rect 91 130 92 131
rect 90 130 91 131
rect 89 130 90 131
rect 88 130 89 131
rect 74 130 75 131
rect 73 130 74 131
rect 72 130 73 131
rect 71 130 72 131
rect 70 130 71 131
rect 57 130 58 131
rect 56 130 57 131
rect 55 130 56 131
rect 54 130 55 131
rect 53 130 54 131
rect 52 130 53 131
rect 51 130 52 131
rect 50 130 51 131
rect 49 130 50 131
rect 48 130 49 131
rect 47 130 48 131
rect 46 130 47 131
rect 45 130 46 131
rect 44 130 45 131
rect 43 130 44 131
rect 42 130 43 131
rect 36 130 37 131
rect 35 130 36 131
rect 34 130 35 131
rect 33 130 34 131
rect 32 130 33 131
rect 31 130 32 131
rect 30 130 31 131
rect 29 130 30 131
rect 28 130 29 131
rect 27 130 28 131
rect 26 130 27 131
rect 25 130 26 131
rect 24 130 25 131
rect 20 130 21 131
rect 19 130 20 131
rect 18 130 19 131
rect 17 130 18 131
rect 16 130 17 131
rect 15 130 16 131
rect 14 130 15 131
rect 13 130 14 131
rect 12 130 13 131
rect 11 130 12 131
rect 182 131 183 132
rect 181 131 182 132
rect 180 131 181 132
rect 179 131 180 132
rect 178 131 179 132
rect 177 131 178 132
rect 176 131 177 132
rect 175 131 176 132
rect 174 131 175 132
rect 173 131 174 132
rect 172 131 173 132
rect 171 131 172 132
rect 170 131 171 132
rect 169 131 170 132
rect 168 131 169 132
rect 167 131 168 132
rect 166 131 167 132
rect 165 131 166 132
rect 109 131 110 132
rect 108 131 109 132
rect 107 131 108 132
rect 106 131 107 132
rect 105 131 106 132
rect 104 131 105 132
rect 103 131 104 132
rect 102 131 103 132
rect 101 131 102 132
rect 100 131 101 132
rect 99 131 100 132
rect 98 131 99 132
rect 97 131 98 132
rect 96 131 97 132
rect 95 131 96 132
rect 94 131 95 132
rect 93 131 94 132
rect 92 131 93 132
rect 91 131 92 132
rect 90 131 91 132
rect 89 131 90 132
rect 88 131 89 132
rect 87 131 88 132
rect 58 131 59 132
rect 57 131 58 132
rect 56 131 57 132
rect 55 131 56 132
rect 54 131 55 132
rect 53 131 54 132
rect 52 131 53 132
rect 51 131 52 132
rect 50 131 51 132
rect 49 131 50 132
rect 48 131 49 132
rect 47 131 48 132
rect 46 131 47 132
rect 45 131 46 132
rect 44 131 45 132
rect 43 131 44 132
rect 36 131 37 132
rect 35 131 36 132
rect 34 131 35 132
rect 33 131 34 132
rect 32 131 33 132
rect 31 131 32 132
rect 30 131 31 132
rect 29 131 30 132
rect 28 131 29 132
rect 27 131 28 132
rect 26 131 27 132
rect 25 131 26 132
rect 20 131 21 132
rect 19 131 20 132
rect 18 131 19 132
rect 17 131 18 132
rect 16 131 17 132
rect 15 131 16 132
rect 14 131 15 132
rect 13 131 14 132
rect 12 131 13 132
rect 11 131 12 132
rect 182 132 183 133
rect 181 132 182 133
rect 180 132 181 133
rect 179 132 180 133
rect 178 132 179 133
rect 177 132 178 133
rect 176 132 177 133
rect 175 132 176 133
rect 174 132 175 133
rect 173 132 174 133
rect 172 132 173 133
rect 171 132 172 133
rect 170 132 171 133
rect 169 132 170 133
rect 168 132 169 133
rect 167 132 168 133
rect 166 132 167 133
rect 165 132 166 133
rect 107 132 108 133
rect 106 132 107 133
rect 105 132 106 133
rect 104 132 105 133
rect 103 132 104 133
rect 102 132 103 133
rect 101 132 102 133
rect 100 132 101 133
rect 99 132 100 133
rect 98 132 99 133
rect 97 132 98 133
rect 96 132 97 133
rect 95 132 96 133
rect 94 132 95 133
rect 93 132 94 133
rect 92 132 93 133
rect 91 132 92 133
rect 90 132 91 133
rect 89 132 90 133
rect 88 132 89 133
rect 87 132 88 133
rect 86 132 87 133
rect 59 132 60 133
rect 58 132 59 133
rect 57 132 58 133
rect 56 132 57 133
rect 55 132 56 133
rect 54 132 55 133
rect 53 132 54 133
rect 52 132 53 133
rect 51 132 52 133
rect 50 132 51 133
rect 49 132 50 133
rect 48 132 49 133
rect 47 132 48 133
rect 46 132 47 133
rect 45 132 46 133
rect 44 132 45 133
rect 43 132 44 133
rect 36 132 37 133
rect 35 132 36 133
rect 34 132 35 133
rect 33 132 34 133
rect 32 132 33 133
rect 31 132 32 133
rect 30 132 31 133
rect 29 132 30 133
rect 28 132 29 133
rect 27 132 28 133
rect 26 132 27 133
rect 25 132 26 133
rect 20 132 21 133
rect 19 132 20 133
rect 18 132 19 133
rect 17 132 18 133
rect 16 132 17 133
rect 15 132 16 133
rect 14 132 15 133
rect 13 132 14 133
rect 12 132 13 133
rect 191 133 192 134
rect 182 133 183 134
rect 181 133 182 134
rect 180 133 181 134
rect 179 133 180 134
rect 178 133 179 134
rect 177 133 178 134
rect 176 133 177 134
rect 175 133 176 134
rect 174 133 175 134
rect 173 133 174 134
rect 172 133 173 134
rect 171 133 172 134
rect 170 133 171 134
rect 169 133 170 134
rect 168 133 169 134
rect 167 133 168 134
rect 166 133 167 134
rect 165 133 166 134
rect 105 133 106 134
rect 104 133 105 134
rect 103 133 104 134
rect 102 133 103 134
rect 101 133 102 134
rect 100 133 101 134
rect 99 133 100 134
rect 98 133 99 134
rect 97 133 98 134
rect 96 133 97 134
rect 95 133 96 134
rect 94 133 95 134
rect 93 133 94 134
rect 92 133 93 134
rect 91 133 92 134
rect 90 133 91 134
rect 89 133 90 134
rect 88 133 89 134
rect 87 133 88 134
rect 86 133 87 134
rect 85 133 86 134
rect 60 133 61 134
rect 59 133 60 134
rect 58 133 59 134
rect 57 133 58 134
rect 56 133 57 134
rect 55 133 56 134
rect 54 133 55 134
rect 53 133 54 134
rect 52 133 53 134
rect 51 133 52 134
rect 50 133 51 134
rect 49 133 50 134
rect 48 133 49 134
rect 47 133 48 134
rect 46 133 47 134
rect 45 133 46 134
rect 44 133 45 134
rect 37 133 38 134
rect 36 133 37 134
rect 35 133 36 134
rect 34 133 35 134
rect 33 133 34 134
rect 32 133 33 134
rect 31 133 32 134
rect 30 133 31 134
rect 29 133 30 134
rect 28 133 29 134
rect 27 133 28 134
rect 26 133 27 134
rect 25 133 26 134
rect 20 133 21 134
rect 19 133 20 134
rect 18 133 19 134
rect 17 133 18 134
rect 16 133 17 134
rect 15 133 16 134
rect 14 133 15 134
rect 13 133 14 134
rect 12 133 13 134
rect 193 134 194 135
rect 192 134 193 135
rect 191 134 192 135
rect 182 134 183 135
rect 181 134 182 135
rect 180 134 181 135
rect 179 134 180 135
rect 178 134 179 135
rect 177 134 178 135
rect 176 134 177 135
rect 175 134 176 135
rect 174 134 175 135
rect 173 134 174 135
rect 172 134 173 135
rect 171 134 172 135
rect 170 134 171 135
rect 169 134 170 135
rect 168 134 169 135
rect 167 134 168 135
rect 166 134 167 135
rect 165 134 166 135
rect 103 134 104 135
rect 102 134 103 135
rect 101 134 102 135
rect 100 134 101 135
rect 99 134 100 135
rect 98 134 99 135
rect 97 134 98 135
rect 96 134 97 135
rect 95 134 96 135
rect 94 134 95 135
rect 93 134 94 135
rect 92 134 93 135
rect 91 134 92 135
rect 90 134 91 135
rect 89 134 90 135
rect 88 134 89 135
rect 87 134 88 135
rect 86 134 87 135
rect 85 134 86 135
rect 84 134 85 135
rect 61 134 62 135
rect 60 134 61 135
rect 59 134 60 135
rect 58 134 59 135
rect 57 134 58 135
rect 56 134 57 135
rect 55 134 56 135
rect 54 134 55 135
rect 53 134 54 135
rect 52 134 53 135
rect 51 134 52 135
rect 50 134 51 135
rect 49 134 50 135
rect 48 134 49 135
rect 47 134 48 135
rect 46 134 47 135
rect 45 134 46 135
rect 37 134 38 135
rect 36 134 37 135
rect 35 134 36 135
rect 34 134 35 135
rect 33 134 34 135
rect 32 134 33 135
rect 31 134 32 135
rect 30 134 31 135
rect 29 134 30 135
rect 28 134 29 135
rect 27 134 28 135
rect 26 134 27 135
rect 21 134 22 135
rect 20 134 21 135
rect 19 134 20 135
rect 18 134 19 135
rect 17 134 18 135
rect 16 134 17 135
rect 15 134 16 135
rect 14 134 15 135
rect 13 134 14 135
rect 199 135 200 136
rect 198 135 199 136
rect 197 135 198 136
rect 196 135 197 136
rect 195 135 196 136
rect 194 135 195 136
rect 193 135 194 136
rect 192 135 193 136
rect 191 135 192 136
rect 182 135 183 136
rect 181 135 182 136
rect 165 135 166 136
rect 100 135 101 136
rect 99 135 100 136
rect 98 135 99 136
rect 97 135 98 136
rect 96 135 97 136
rect 95 135 96 136
rect 94 135 95 136
rect 93 135 94 136
rect 92 135 93 136
rect 91 135 92 136
rect 90 135 91 136
rect 89 135 90 136
rect 88 135 89 136
rect 87 135 88 136
rect 86 135 87 136
rect 85 135 86 136
rect 84 135 85 136
rect 83 135 84 136
rect 63 135 64 136
rect 62 135 63 136
rect 61 135 62 136
rect 60 135 61 136
rect 59 135 60 136
rect 58 135 59 136
rect 57 135 58 136
rect 56 135 57 136
rect 55 135 56 136
rect 54 135 55 136
rect 53 135 54 136
rect 52 135 53 136
rect 51 135 52 136
rect 50 135 51 136
rect 49 135 50 136
rect 48 135 49 136
rect 47 135 48 136
rect 46 135 47 136
rect 45 135 46 136
rect 38 135 39 136
rect 37 135 38 136
rect 36 135 37 136
rect 35 135 36 136
rect 34 135 35 136
rect 33 135 34 136
rect 32 135 33 136
rect 31 135 32 136
rect 30 135 31 136
rect 29 135 30 136
rect 28 135 29 136
rect 27 135 28 136
rect 26 135 27 136
rect 21 135 22 136
rect 20 135 21 136
rect 19 135 20 136
rect 18 135 19 136
rect 17 135 18 136
rect 16 135 17 136
rect 15 135 16 136
rect 14 135 15 136
rect 198 136 199 137
rect 197 136 198 137
rect 196 136 197 137
rect 195 136 196 137
rect 194 136 195 137
rect 182 136 183 137
rect 165 136 166 137
rect 95 136 96 137
rect 94 136 95 137
rect 93 136 94 137
rect 92 136 93 137
rect 91 136 92 137
rect 90 136 91 137
rect 89 136 90 137
rect 88 136 89 137
rect 87 136 88 137
rect 85 136 86 137
rect 64 136 65 137
rect 63 136 64 137
rect 62 136 63 137
rect 61 136 62 137
rect 60 136 61 137
rect 59 136 60 137
rect 58 136 59 137
rect 57 136 58 137
rect 56 136 57 137
rect 55 136 56 137
rect 54 136 55 137
rect 53 136 54 137
rect 52 136 53 137
rect 51 136 52 137
rect 50 136 51 137
rect 49 136 50 137
rect 48 136 49 137
rect 47 136 48 137
rect 46 136 47 137
rect 38 136 39 137
rect 37 136 38 137
rect 36 136 37 137
rect 35 136 36 137
rect 34 136 35 137
rect 33 136 34 137
rect 32 136 33 137
rect 31 136 32 137
rect 30 136 31 137
rect 29 136 30 137
rect 28 136 29 137
rect 27 136 28 137
rect 26 136 27 137
rect 21 136 22 137
rect 20 136 21 137
rect 19 136 20 137
rect 18 136 19 137
rect 17 136 18 137
rect 16 136 17 137
rect 15 136 16 137
rect 198 137 199 138
rect 197 137 198 138
rect 196 137 197 138
rect 195 137 196 138
rect 194 137 195 138
rect 193 137 194 138
rect 66 137 67 138
rect 65 137 66 138
rect 64 137 65 138
rect 63 137 64 138
rect 62 137 63 138
rect 61 137 62 138
rect 60 137 61 138
rect 59 137 60 138
rect 58 137 59 138
rect 57 137 58 138
rect 56 137 57 138
rect 55 137 56 138
rect 54 137 55 138
rect 53 137 54 138
rect 52 137 53 138
rect 51 137 52 138
rect 50 137 51 138
rect 49 137 50 138
rect 48 137 49 138
rect 47 137 48 138
rect 39 137 40 138
rect 38 137 39 138
rect 37 137 38 138
rect 36 137 37 138
rect 35 137 36 138
rect 34 137 35 138
rect 33 137 34 138
rect 32 137 33 138
rect 31 137 32 138
rect 30 137 31 138
rect 29 137 30 138
rect 28 137 29 138
rect 27 137 28 138
rect 22 137 23 138
rect 21 137 22 138
rect 20 137 21 138
rect 19 137 20 138
rect 18 137 19 138
rect 17 137 18 138
rect 16 137 17 138
rect 15 137 16 138
rect 193 138 194 139
rect 192 138 193 139
rect 191 138 192 139
rect 68 138 69 139
rect 67 138 68 139
rect 66 138 67 139
rect 65 138 66 139
rect 64 138 65 139
rect 63 138 64 139
rect 62 138 63 139
rect 61 138 62 139
rect 60 138 61 139
rect 59 138 60 139
rect 58 138 59 139
rect 57 138 58 139
rect 56 138 57 139
rect 55 138 56 139
rect 54 138 55 139
rect 53 138 54 139
rect 52 138 53 139
rect 51 138 52 139
rect 50 138 51 139
rect 49 138 50 139
rect 48 138 49 139
rect 40 138 41 139
rect 39 138 40 139
rect 38 138 39 139
rect 37 138 38 139
rect 36 138 37 139
rect 35 138 36 139
rect 34 138 35 139
rect 33 138 34 139
rect 32 138 33 139
rect 31 138 32 139
rect 30 138 31 139
rect 29 138 30 139
rect 28 138 29 139
rect 27 138 28 139
rect 22 138 23 139
rect 21 138 22 139
rect 20 138 21 139
rect 19 138 20 139
rect 18 138 19 139
rect 17 138 18 139
rect 16 138 17 139
rect 191 139 192 140
rect 71 139 72 140
rect 70 139 71 140
rect 69 139 70 140
rect 68 139 69 140
rect 67 139 68 140
rect 66 139 67 140
rect 65 139 66 140
rect 64 139 65 140
rect 63 139 64 140
rect 62 139 63 140
rect 61 139 62 140
rect 60 139 61 140
rect 59 139 60 140
rect 58 139 59 140
rect 57 139 58 140
rect 56 139 57 140
rect 55 139 56 140
rect 54 139 55 140
rect 53 139 54 140
rect 52 139 53 140
rect 51 139 52 140
rect 50 139 51 140
rect 49 139 50 140
rect 40 139 41 140
rect 39 139 40 140
rect 38 139 39 140
rect 37 139 38 140
rect 36 139 37 140
rect 35 139 36 140
rect 34 139 35 140
rect 33 139 34 140
rect 32 139 33 140
rect 31 139 32 140
rect 30 139 31 140
rect 29 139 30 140
rect 28 139 29 140
rect 27 139 28 140
rect 22 139 23 140
rect 21 139 22 140
rect 20 139 21 140
rect 19 139 20 140
rect 18 139 19 140
rect 17 139 18 140
rect 182 140 183 141
rect 165 140 166 141
rect 74 140 75 141
rect 73 140 74 141
rect 72 140 73 141
rect 71 140 72 141
rect 70 140 71 141
rect 69 140 70 141
rect 68 140 69 141
rect 67 140 68 141
rect 66 140 67 141
rect 65 140 66 141
rect 64 140 65 141
rect 63 140 64 141
rect 62 140 63 141
rect 61 140 62 141
rect 60 140 61 141
rect 59 140 60 141
rect 58 140 59 141
rect 57 140 58 141
rect 56 140 57 141
rect 55 140 56 141
rect 54 140 55 141
rect 53 140 54 141
rect 52 140 53 141
rect 51 140 52 141
rect 50 140 51 141
rect 49 140 50 141
rect 41 140 42 141
rect 40 140 41 141
rect 39 140 40 141
rect 38 140 39 141
rect 37 140 38 141
rect 36 140 37 141
rect 35 140 36 141
rect 34 140 35 141
rect 33 140 34 141
rect 32 140 33 141
rect 31 140 32 141
rect 30 140 31 141
rect 29 140 30 141
rect 28 140 29 141
rect 23 140 24 141
rect 22 140 23 141
rect 21 140 22 141
rect 20 140 21 141
rect 19 140 20 141
rect 18 140 19 141
rect 182 141 183 142
rect 165 141 166 142
rect 78 141 79 142
rect 77 141 78 142
rect 76 141 77 142
rect 75 141 76 142
rect 74 141 75 142
rect 73 141 74 142
rect 72 141 73 142
rect 71 141 72 142
rect 70 141 71 142
rect 69 141 70 142
rect 68 141 69 142
rect 67 141 68 142
rect 66 141 67 142
rect 65 141 66 142
rect 64 141 65 142
rect 63 141 64 142
rect 62 141 63 142
rect 61 141 62 142
rect 60 141 61 142
rect 59 141 60 142
rect 58 141 59 142
rect 57 141 58 142
rect 56 141 57 142
rect 55 141 56 142
rect 54 141 55 142
rect 53 141 54 142
rect 52 141 53 142
rect 51 141 52 142
rect 50 141 51 142
rect 42 141 43 142
rect 41 141 42 142
rect 40 141 41 142
rect 39 141 40 142
rect 38 141 39 142
rect 37 141 38 142
rect 36 141 37 142
rect 35 141 36 142
rect 34 141 35 142
rect 33 141 34 142
rect 32 141 33 142
rect 31 141 32 142
rect 30 141 31 142
rect 29 141 30 142
rect 28 141 29 142
rect 23 141 24 142
rect 22 141 23 142
rect 21 141 22 142
rect 20 141 21 142
rect 19 141 20 142
rect 182 142 183 143
rect 181 142 182 143
rect 180 142 181 143
rect 179 142 180 143
rect 178 142 179 143
rect 177 142 178 143
rect 176 142 177 143
rect 175 142 176 143
rect 174 142 175 143
rect 173 142 174 143
rect 172 142 173 143
rect 171 142 172 143
rect 170 142 171 143
rect 169 142 170 143
rect 168 142 169 143
rect 167 142 168 143
rect 166 142 167 143
rect 165 142 166 143
rect 77 142 78 143
rect 76 142 77 143
rect 75 142 76 143
rect 74 142 75 143
rect 73 142 74 143
rect 72 142 73 143
rect 71 142 72 143
rect 70 142 71 143
rect 69 142 70 143
rect 68 142 69 143
rect 67 142 68 143
rect 66 142 67 143
rect 65 142 66 143
rect 64 142 65 143
rect 63 142 64 143
rect 62 142 63 143
rect 61 142 62 143
rect 60 142 61 143
rect 59 142 60 143
rect 58 142 59 143
rect 57 142 58 143
rect 56 142 57 143
rect 55 142 56 143
rect 54 142 55 143
rect 53 142 54 143
rect 52 142 53 143
rect 51 142 52 143
rect 43 142 44 143
rect 42 142 43 143
rect 41 142 42 143
rect 40 142 41 143
rect 39 142 40 143
rect 38 142 39 143
rect 37 142 38 143
rect 36 142 37 143
rect 35 142 36 143
rect 34 142 35 143
rect 33 142 34 143
rect 32 142 33 143
rect 31 142 32 143
rect 30 142 31 143
rect 29 142 30 143
rect 24 142 25 143
rect 23 142 24 143
rect 22 142 23 143
rect 21 142 22 143
rect 20 142 21 143
rect 182 143 183 144
rect 181 143 182 144
rect 180 143 181 144
rect 179 143 180 144
rect 178 143 179 144
rect 177 143 178 144
rect 176 143 177 144
rect 175 143 176 144
rect 174 143 175 144
rect 173 143 174 144
rect 172 143 173 144
rect 171 143 172 144
rect 170 143 171 144
rect 169 143 170 144
rect 168 143 169 144
rect 167 143 168 144
rect 166 143 167 144
rect 165 143 166 144
rect 76 143 77 144
rect 75 143 76 144
rect 74 143 75 144
rect 73 143 74 144
rect 72 143 73 144
rect 71 143 72 144
rect 70 143 71 144
rect 69 143 70 144
rect 68 143 69 144
rect 67 143 68 144
rect 66 143 67 144
rect 65 143 66 144
rect 64 143 65 144
rect 63 143 64 144
rect 62 143 63 144
rect 61 143 62 144
rect 60 143 61 144
rect 59 143 60 144
rect 58 143 59 144
rect 57 143 58 144
rect 56 143 57 144
rect 55 143 56 144
rect 54 143 55 144
rect 53 143 54 144
rect 52 143 53 144
rect 43 143 44 144
rect 42 143 43 144
rect 41 143 42 144
rect 40 143 41 144
rect 39 143 40 144
rect 38 143 39 144
rect 37 143 38 144
rect 36 143 37 144
rect 35 143 36 144
rect 34 143 35 144
rect 33 143 34 144
rect 32 143 33 144
rect 31 143 32 144
rect 30 143 31 144
rect 29 143 30 144
rect 24 143 25 144
rect 23 143 24 144
rect 22 143 23 144
rect 21 143 22 144
rect 182 144 183 145
rect 181 144 182 145
rect 180 144 181 145
rect 179 144 180 145
rect 178 144 179 145
rect 177 144 178 145
rect 176 144 177 145
rect 175 144 176 145
rect 174 144 175 145
rect 173 144 174 145
rect 172 144 173 145
rect 171 144 172 145
rect 170 144 171 145
rect 169 144 170 145
rect 168 144 169 145
rect 167 144 168 145
rect 166 144 167 145
rect 165 144 166 145
rect 74 144 75 145
rect 73 144 74 145
rect 72 144 73 145
rect 71 144 72 145
rect 70 144 71 145
rect 69 144 70 145
rect 68 144 69 145
rect 67 144 68 145
rect 66 144 67 145
rect 65 144 66 145
rect 64 144 65 145
rect 63 144 64 145
rect 62 144 63 145
rect 61 144 62 145
rect 60 144 61 145
rect 59 144 60 145
rect 58 144 59 145
rect 57 144 58 145
rect 56 144 57 145
rect 55 144 56 145
rect 54 144 55 145
rect 53 144 54 145
rect 44 144 45 145
rect 43 144 44 145
rect 42 144 43 145
rect 41 144 42 145
rect 40 144 41 145
rect 39 144 40 145
rect 38 144 39 145
rect 37 144 38 145
rect 36 144 37 145
rect 35 144 36 145
rect 34 144 35 145
rect 33 144 34 145
rect 32 144 33 145
rect 31 144 32 145
rect 30 144 31 145
rect 29 144 30 145
rect 25 144 26 145
rect 24 144 25 145
rect 23 144 24 145
rect 22 144 23 145
rect 182 145 183 146
rect 181 145 182 146
rect 180 145 181 146
rect 179 145 180 146
rect 178 145 179 146
rect 177 145 178 146
rect 176 145 177 146
rect 175 145 176 146
rect 174 145 175 146
rect 173 145 174 146
rect 172 145 173 146
rect 171 145 172 146
rect 170 145 171 146
rect 169 145 170 146
rect 168 145 169 146
rect 167 145 168 146
rect 166 145 167 146
rect 165 145 166 146
rect 72 145 73 146
rect 71 145 72 146
rect 70 145 71 146
rect 69 145 70 146
rect 68 145 69 146
rect 67 145 68 146
rect 66 145 67 146
rect 65 145 66 146
rect 64 145 65 146
rect 63 145 64 146
rect 62 145 63 146
rect 61 145 62 146
rect 60 145 61 146
rect 59 145 60 146
rect 58 145 59 146
rect 57 145 58 146
rect 56 145 57 146
rect 55 145 56 146
rect 45 145 46 146
rect 44 145 45 146
rect 43 145 44 146
rect 42 145 43 146
rect 41 145 42 146
rect 40 145 41 146
rect 39 145 40 146
rect 38 145 39 146
rect 37 145 38 146
rect 36 145 37 146
rect 35 145 36 146
rect 34 145 35 146
rect 33 145 34 146
rect 32 145 33 146
rect 31 145 32 146
rect 30 145 31 146
rect 25 145 26 146
rect 182 146 183 147
rect 181 146 182 147
rect 174 146 175 147
rect 173 146 174 147
rect 172 146 173 147
rect 166 146 167 147
rect 165 146 166 147
rect 67 146 68 147
rect 66 146 67 147
rect 65 146 66 147
rect 64 146 65 147
rect 63 146 64 147
rect 62 146 63 147
rect 61 146 62 147
rect 60 146 61 147
rect 59 146 60 147
rect 58 146 59 147
rect 46 146 47 147
rect 45 146 46 147
rect 44 146 45 147
rect 43 146 44 147
rect 42 146 43 147
rect 41 146 42 147
rect 40 146 41 147
rect 39 146 40 147
rect 38 146 39 147
rect 37 146 38 147
rect 36 146 37 147
rect 35 146 36 147
rect 34 146 35 147
rect 33 146 34 147
rect 32 146 33 147
rect 31 146 32 147
rect 30 146 31 147
rect 182 147 183 148
rect 174 147 175 148
rect 173 147 174 148
rect 165 147 166 148
rect 47 147 48 148
rect 46 147 47 148
rect 45 147 46 148
rect 44 147 45 148
rect 43 147 44 148
rect 42 147 43 148
rect 41 147 42 148
rect 40 147 41 148
rect 39 147 40 148
rect 38 147 39 148
rect 37 147 38 148
rect 36 147 37 148
rect 35 147 36 148
rect 34 147 35 148
rect 33 147 34 148
rect 32 147 33 148
rect 31 147 32 148
rect 182 148 183 149
rect 174 148 175 149
rect 173 148 174 149
rect 165 148 166 149
rect 49 148 50 149
rect 48 148 49 149
rect 47 148 48 149
rect 46 148 47 149
rect 45 148 46 149
rect 44 148 45 149
rect 43 148 44 149
rect 42 148 43 149
rect 41 148 42 149
rect 40 148 41 149
rect 39 148 40 149
rect 38 148 39 149
rect 37 148 38 149
rect 36 148 37 149
rect 35 148 36 149
rect 34 148 35 149
rect 33 148 34 149
rect 32 148 33 149
rect 182 149 183 150
rect 174 149 175 150
rect 173 149 174 150
rect 165 149 166 150
rect 50 149 51 150
rect 49 149 50 150
rect 48 149 49 150
rect 47 149 48 150
rect 46 149 47 150
rect 45 149 46 150
rect 44 149 45 150
rect 43 149 44 150
rect 42 149 43 150
rect 41 149 42 150
rect 40 149 41 150
rect 39 149 40 150
rect 38 149 39 150
rect 37 149 38 150
rect 36 149 37 150
rect 35 149 36 150
rect 34 149 35 150
rect 33 149 34 150
rect 182 150 183 151
rect 175 150 176 151
rect 174 150 175 151
rect 173 150 174 151
rect 172 150 173 151
rect 166 150 167 151
rect 165 150 166 151
rect 52 150 53 151
rect 51 150 52 151
rect 50 150 51 151
rect 49 150 50 151
rect 48 150 49 151
rect 47 150 48 151
rect 46 150 47 151
rect 45 150 46 151
rect 44 150 45 151
rect 43 150 44 151
rect 42 150 43 151
rect 41 150 42 151
rect 40 150 41 151
rect 39 150 40 151
rect 38 150 39 151
rect 37 150 38 151
rect 36 150 37 151
rect 35 150 36 151
rect 34 150 35 151
rect 182 151 183 152
rect 181 151 182 152
rect 176 151 177 152
rect 175 151 176 152
rect 174 151 175 152
rect 173 151 174 152
rect 172 151 173 152
rect 171 151 172 152
rect 166 151 167 152
rect 165 151 166 152
rect 53 151 54 152
rect 52 151 53 152
rect 51 151 52 152
rect 50 151 51 152
rect 49 151 50 152
rect 48 151 49 152
rect 47 151 48 152
rect 46 151 47 152
rect 45 151 46 152
rect 44 151 45 152
rect 43 151 44 152
rect 42 151 43 152
rect 41 151 42 152
rect 40 151 41 152
rect 39 151 40 152
rect 38 151 39 152
rect 37 151 38 152
rect 36 151 37 152
rect 182 152 183 153
rect 181 152 182 153
rect 180 152 181 153
rect 169 152 170 153
rect 168 152 169 153
rect 167 152 168 153
rect 166 152 167 153
rect 165 152 166 153
rect 53 152 54 153
rect 52 152 53 153
rect 51 152 52 153
rect 50 152 51 153
rect 49 152 50 153
rect 48 152 49 153
rect 47 152 48 153
rect 46 152 47 153
rect 45 152 46 153
rect 44 152 45 153
rect 43 152 44 153
rect 42 152 43 153
rect 41 152 42 153
rect 40 152 41 153
rect 39 152 40 153
rect 182 153 183 154
rect 181 153 182 154
rect 180 153 181 154
rect 179 153 180 154
rect 178 153 179 154
rect 168 153 169 154
rect 167 153 168 154
rect 166 153 167 154
rect 49 153 50 154
rect 48 153 49 154
rect 47 153 48 154
rect 46 153 47 154
rect 45 153 46 154
rect 44 153 45 154
rect 180 154 181 155
rect 179 154 180 155
rect 178 154 179 155
rect 182 157 183 158
rect 165 157 166 158
rect 182 158 183 159
rect 165 158 166 159
rect 182 159 183 160
rect 181 159 182 160
rect 180 159 181 160
rect 179 159 180 160
rect 178 159 179 160
rect 177 159 178 160
rect 176 159 177 160
rect 175 159 176 160
rect 174 159 175 160
rect 173 159 174 160
rect 172 159 173 160
rect 171 159 172 160
rect 170 159 171 160
rect 169 159 170 160
rect 168 159 169 160
rect 167 159 168 160
rect 166 159 167 160
rect 165 159 166 160
rect 182 160 183 161
rect 181 160 182 161
rect 180 160 181 161
rect 179 160 180 161
rect 178 160 179 161
rect 177 160 178 161
rect 176 160 177 161
rect 175 160 176 161
rect 174 160 175 161
rect 173 160 174 161
rect 172 160 173 161
rect 171 160 172 161
rect 170 160 171 161
rect 169 160 170 161
rect 168 160 169 161
rect 167 160 168 161
rect 166 160 167 161
rect 165 160 166 161
rect 182 161 183 162
rect 181 161 182 162
rect 180 161 181 162
rect 179 161 180 162
rect 178 161 179 162
rect 177 161 178 162
rect 176 161 177 162
rect 175 161 176 162
rect 174 161 175 162
rect 173 161 174 162
rect 172 161 173 162
rect 171 161 172 162
rect 170 161 171 162
rect 169 161 170 162
rect 168 161 169 162
rect 167 161 168 162
rect 166 161 167 162
rect 165 161 166 162
rect 182 162 183 163
rect 181 162 182 163
rect 180 162 181 163
rect 179 162 180 163
rect 178 162 179 163
rect 177 162 178 163
rect 176 162 177 163
rect 175 162 176 163
rect 174 162 175 163
rect 173 162 174 163
rect 172 162 173 163
rect 171 162 172 163
rect 170 162 171 163
rect 169 162 170 163
rect 168 162 169 163
rect 167 162 168 163
rect 166 162 167 163
rect 165 162 166 163
rect 182 163 183 164
rect 181 163 182 164
rect 180 163 181 164
rect 179 163 180 164
rect 178 163 179 164
rect 177 163 178 164
rect 176 163 177 164
rect 175 163 176 164
rect 174 163 175 164
rect 173 163 174 164
rect 172 163 173 164
rect 171 163 172 164
rect 170 163 171 164
rect 169 163 170 164
rect 168 163 169 164
rect 167 163 168 164
rect 166 163 167 164
rect 165 163 166 164
rect 182 164 183 165
rect 181 164 182 165
rect 174 164 175 165
rect 173 164 174 165
rect 165 164 166 165
rect 182 165 183 166
rect 174 165 175 166
rect 173 165 174 166
rect 165 165 166 166
rect 182 166 183 167
rect 174 166 175 167
rect 173 166 174 167
rect 165 166 166 167
rect 182 167 183 168
rect 174 167 175 168
rect 173 167 174 168
rect 172 167 173 168
rect 166 167 167 168
rect 165 167 166 168
rect 182 168 183 169
rect 181 168 182 169
rect 176 168 177 169
rect 175 168 176 169
rect 174 168 175 169
rect 173 168 174 169
rect 172 168 173 169
rect 171 168 172 169
rect 166 168 167 169
rect 165 168 166 169
rect 182 169 183 170
rect 181 169 182 170
rect 180 169 181 170
rect 175 169 176 170
rect 174 169 175 170
rect 173 169 174 170
rect 172 169 173 170
rect 171 169 172 170
rect 168 169 169 170
rect 167 169 168 170
rect 166 169 167 170
rect 165 169 166 170
rect 182 170 183 171
rect 181 170 182 171
rect 180 170 181 171
rect 179 170 180 171
rect 168 170 169 171
rect 167 170 168 171
rect 166 170 167 171
rect 165 170 166 171
rect 181 171 182 172
rect 180 171 181 172
rect 179 171 180 172
rect 178 171 179 172
rect 145 178 146 179
rect 144 178 145 179
rect 143 178 144 179
rect 142 178 143 179
rect 141 178 142 179
rect 140 178 141 179
rect 139 178 140 179
rect 138 178 139 179
rect 137 178 138 179
rect 136 178 137 179
rect 135 178 136 179
rect 134 178 135 179
rect 133 178 134 179
rect 132 178 133 179
rect 131 178 132 179
rect 130 178 131 179
rect 129 178 130 179
rect 128 178 129 179
rect 127 178 128 179
rect 126 178 127 179
rect 125 178 126 179
rect 124 178 125 179
rect 123 178 124 179
rect 122 178 123 179
rect 121 178 122 179
rect 120 178 121 179
rect 119 178 120 179
rect 118 178 119 179
rect 117 178 118 179
rect 116 178 117 179
rect 115 178 116 179
rect 114 178 115 179
rect 113 178 114 179
rect 112 178 113 179
rect 111 178 112 179
rect 110 178 111 179
rect 109 178 110 179
rect 108 178 109 179
rect 107 178 108 179
rect 106 178 107 179
rect 105 178 106 179
rect 104 178 105 179
rect 147 179 148 180
rect 146 179 147 180
rect 145 179 146 180
rect 144 179 145 180
rect 143 179 144 180
rect 142 179 143 180
rect 141 179 142 180
rect 140 179 141 180
rect 139 179 140 180
rect 138 179 139 180
rect 137 179 138 180
rect 136 179 137 180
rect 135 179 136 180
rect 134 179 135 180
rect 133 179 134 180
rect 132 179 133 180
rect 131 179 132 180
rect 130 179 131 180
rect 129 179 130 180
rect 128 179 129 180
rect 127 179 128 180
rect 126 179 127 180
rect 125 179 126 180
rect 124 179 125 180
rect 123 179 124 180
rect 122 179 123 180
rect 121 179 122 180
rect 120 179 121 180
rect 119 179 120 180
rect 118 179 119 180
rect 117 179 118 180
rect 116 179 117 180
rect 115 179 116 180
rect 114 179 115 180
rect 113 179 114 180
rect 112 179 113 180
rect 111 179 112 180
rect 110 179 111 180
rect 109 179 110 180
rect 108 179 109 180
rect 107 179 108 180
rect 106 179 107 180
rect 105 179 106 180
rect 104 179 105 180
rect 198 180 199 181
rect 197 180 198 181
rect 196 180 197 181
rect 195 180 196 181
rect 194 180 195 181
rect 193 180 194 181
rect 192 180 193 181
rect 191 180 192 181
rect 174 180 175 181
rect 169 180 170 181
rect 168 180 169 181
rect 167 180 168 181
rect 148 180 149 181
rect 147 180 148 181
rect 146 180 147 181
rect 145 180 146 181
rect 144 180 145 181
rect 143 180 144 181
rect 142 180 143 181
rect 141 180 142 181
rect 140 180 141 181
rect 139 180 140 181
rect 138 180 139 181
rect 137 180 138 181
rect 136 180 137 181
rect 135 180 136 181
rect 134 180 135 181
rect 133 180 134 181
rect 132 180 133 181
rect 131 180 132 181
rect 130 180 131 181
rect 129 180 130 181
rect 128 180 129 181
rect 127 180 128 181
rect 126 180 127 181
rect 125 180 126 181
rect 124 180 125 181
rect 123 180 124 181
rect 122 180 123 181
rect 121 180 122 181
rect 120 180 121 181
rect 119 180 120 181
rect 118 180 119 181
rect 117 180 118 181
rect 116 180 117 181
rect 115 180 116 181
rect 114 180 115 181
rect 113 180 114 181
rect 112 180 113 181
rect 111 180 112 181
rect 110 180 111 181
rect 109 180 110 181
rect 108 180 109 181
rect 107 180 108 181
rect 106 180 107 181
rect 105 180 106 181
rect 104 180 105 181
rect 199 181 200 182
rect 198 181 199 182
rect 197 181 198 182
rect 196 181 197 182
rect 195 181 196 182
rect 194 181 195 182
rect 193 181 194 182
rect 192 181 193 182
rect 191 181 192 182
rect 176 181 177 182
rect 175 181 176 182
rect 174 181 175 182
rect 173 181 174 182
rect 172 181 173 182
rect 169 181 170 182
rect 168 181 169 182
rect 167 181 168 182
rect 149 181 150 182
rect 148 181 149 182
rect 147 181 148 182
rect 146 181 147 182
rect 145 181 146 182
rect 144 181 145 182
rect 143 181 144 182
rect 142 181 143 182
rect 141 181 142 182
rect 140 181 141 182
rect 139 181 140 182
rect 138 181 139 182
rect 137 181 138 182
rect 136 181 137 182
rect 135 181 136 182
rect 134 181 135 182
rect 133 181 134 182
rect 132 181 133 182
rect 131 181 132 182
rect 130 181 131 182
rect 129 181 130 182
rect 128 181 129 182
rect 127 181 128 182
rect 126 181 127 182
rect 125 181 126 182
rect 124 181 125 182
rect 123 181 124 182
rect 122 181 123 182
rect 121 181 122 182
rect 120 181 121 182
rect 119 181 120 182
rect 118 181 119 182
rect 117 181 118 182
rect 116 181 117 182
rect 115 181 116 182
rect 114 181 115 182
rect 113 181 114 182
rect 112 181 113 182
rect 111 181 112 182
rect 110 181 111 182
rect 109 181 110 182
rect 108 181 109 182
rect 107 181 108 182
rect 106 181 107 182
rect 105 181 106 182
rect 104 181 105 182
rect 198 182 199 183
rect 197 182 198 183
rect 196 182 197 183
rect 195 182 196 183
rect 194 182 195 183
rect 193 182 194 183
rect 192 182 193 183
rect 191 182 192 183
rect 176 182 177 183
rect 175 182 176 183
rect 174 182 175 183
rect 173 182 174 183
rect 172 182 173 183
rect 171 182 172 183
rect 169 182 170 183
rect 168 182 169 183
rect 167 182 168 183
rect 150 182 151 183
rect 149 182 150 183
rect 148 182 149 183
rect 147 182 148 183
rect 146 182 147 183
rect 145 182 146 183
rect 144 182 145 183
rect 143 182 144 183
rect 142 182 143 183
rect 141 182 142 183
rect 140 182 141 183
rect 139 182 140 183
rect 138 182 139 183
rect 137 182 138 183
rect 136 182 137 183
rect 135 182 136 183
rect 134 182 135 183
rect 133 182 134 183
rect 132 182 133 183
rect 131 182 132 183
rect 130 182 131 183
rect 129 182 130 183
rect 128 182 129 183
rect 127 182 128 183
rect 126 182 127 183
rect 125 182 126 183
rect 124 182 125 183
rect 123 182 124 183
rect 122 182 123 183
rect 121 182 122 183
rect 120 182 121 183
rect 119 182 120 183
rect 118 182 119 183
rect 117 182 118 183
rect 116 182 117 183
rect 115 182 116 183
rect 114 182 115 183
rect 113 182 114 183
rect 112 182 113 183
rect 111 182 112 183
rect 110 182 111 183
rect 109 182 110 183
rect 108 182 109 183
rect 107 182 108 183
rect 106 182 107 183
rect 105 182 106 183
rect 104 182 105 183
rect 198 183 199 184
rect 195 183 196 184
rect 194 183 195 184
rect 191 183 192 184
rect 184 183 185 184
rect 183 183 184 184
rect 182 183 183 184
rect 181 183 182 184
rect 180 183 181 184
rect 177 183 178 184
rect 176 183 177 184
rect 175 183 176 184
rect 174 183 175 184
rect 173 183 174 184
rect 172 183 173 184
rect 171 183 172 184
rect 169 183 170 184
rect 168 183 169 184
rect 167 183 168 184
rect 165 183 166 184
rect 164 183 165 184
rect 150 183 151 184
rect 149 183 150 184
rect 148 183 149 184
rect 147 183 148 184
rect 146 183 147 184
rect 145 183 146 184
rect 144 183 145 184
rect 143 183 144 184
rect 142 183 143 184
rect 141 183 142 184
rect 140 183 141 184
rect 139 183 140 184
rect 138 183 139 184
rect 137 183 138 184
rect 136 183 137 184
rect 135 183 136 184
rect 134 183 135 184
rect 133 183 134 184
rect 132 183 133 184
rect 131 183 132 184
rect 130 183 131 184
rect 129 183 130 184
rect 128 183 129 184
rect 127 183 128 184
rect 126 183 127 184
rect 125 183 126 184
rect 124 183 125 184
rect 123 183 124 184
rect 122 183 123 184
rect 121 183 122 184
rect 120 183 121 184
rect 119 183 120 184
rect 118 183 119 184
rect 117 183 118 184
rect 116 183 117 184
rect 115 183 116 184
rect 114 183 115 184
rect 113 183 114 184
rect 112 183 113 184
rect 111 183 112 184
rect 110 183 111 184
rect 109 183 110 184
rect 108 183 109 184
rect 107 183 108 184
rect 106 183 107 184
rect 105 183 106 184
rect 104 183 105 184
rect 198 184 199 185
rect 195 184 196 185
rect 194 184 195 185
rect 191 184 192 185
rect 185 184 186 185
rect 184 184 185 185
rect 183 184 184 185
rect 182 184 183 185
rect 181 184 182 185
rect 180 184 181 185
rect 179 184 180 185
rect 177 184 178 185
rect 176 184 177 185
rect 175 184 176 185
rect 174 184 175 185
rect 173 184 174 185
rect 172 184 173 185
rect 171 184 172 185
rect 169 184 170 185
rect 168 184 169 185
rect 167 184 168 185
rect 165 184 166 185
rect 164 184 165 185
rect 151 184 152 185
rect 150 184 151 185
rect 149 184 150 185
rect 148 184 149 185
rect 147 184 148 185
rect 146 184 147 185
rect 145 184 146 185
rect 144 184 145 185
rect 143 184 144 185
rect 142 184 143 185
rect 141 184 142 185
rect 140 184 141 185
rect 139 184 140 185
rect 138 184 139 185
rect 137 184 138 185
rect 136 184 137 185
rect 135 184 136 185
rect 134 184 135 185
rect 133 184 134 185
rect 132 184 133 185
rect 131 184 132 185
rect 130 184 131 185
rect 129 184 130 185
rect 128 184 129 185
rect 127 184 128 185
rect 126 184 127 185
rect 125 184 126 185
rect 124 184 125 185
rect 123 184 124 185
rect 122 184 123 185
rect 121 184 122 185
rect 120 184 121 185
rect 119 184 120 185
rect 118 184 119 185
rect 117 184 118 185
rect 116 184 117 185
rect 115 184 116 185
rect 114 184 115 185
rect 113 184 114 185
rect 112 184 113 185
rect 111 184 112 185
rect 110 184 111 185
rect 109 184 110 185
rect 108 184 109 185
rect 107 184 108 185
rect 106 184 107 185
rect 105 184 106 185
rect 104 184 105 185
rect 64 184 65 185
rect 63 184 64 185
rect 62 184 63 185
rect 61 184 62 185
rect 199 185 200 186
rect 198 185 199 186
rect 195 185 196 186
rect 194 185 195 186
rect 191 185 192 186
rect 185 185 186 186
rect 184 185 185 186
rect 183 185 184 186
rect 182 185 183 186
rect 181 185 182 186
rect 180 185 181 186
rect 179 185 180 186
rect 177 185 178 186
rect 176 185 177 186
rect 175 185 176 186
rect 173 185 174 186
rect 172 185 173 186
rect 171 185 172 186
rect 170 185 171 186
rect 169 185 170 186
rect 168 185 169 186
rect 167 185 168 186
rect 165 185 166 186
rect 164 185 165 186
rect 151 185 152 186
rect 150 185 151 186
rect 149 185 150 186
rect 148 185 149 186
rect 147 185 148 186
rect 146 185 147 186
rect 145 185 146 186
rect 144 185 145 186
rect 143 185 144 186
rect 142 185 143 186
rect 141 185 142 186
rect 140 185 141 186
rect 139 185 140 186
rect 138 185 139 186
rect 137 185 138 186
rect 136 185 137 186
rect 135 185 136 186
rect 134 185 135 186
rect 133 185 134 186
rect 132 185 133 186
rect 131 185 132 186
rect 130 185 131 186
rect 129 185 130 186
rect 128 185 129 186
rect 127 185 128 186
rect 126 185 127 186
rect 125 185 126 186
rect 124 185 125 186
rect 123 185 124 186
rect 122 185 123 186
rect 121 185 122 186
rect 120 185 121 186
rect 119 185 120 186
rect 118 185 119 186
rect 117 185 118 186
rect 116 185 117 186
rect 115 185 116 186
rect 114 185 115 186
rect 113 185 114 186
rect 112 185 113 186
rect 111 185 112 186
rect 110 185 111 186
rect 109 185 110 186
rect 108 185 109 186
rect 107 185 108 186
rect 106 185 107 186
rect 105 185 106 186
rect 104 185 105 186
rect 64 185 65 186
rect 63 185 64 186
rect 62 185 63 186
rect 61 185 62 186
rect 31 185 32 186
rect 30 185 31 186
rect 185 186 186 187
rect 184 186 185 187
rect 183 186 184 187
rect 182 186 183 187
rect 181 186 182 187
rect 180 186 181 187
rect 179 186 180 187
rect 177 186 178 187
rect 176 186 177 187
rect 172 186 173 187
rect 171 186 172 187
rect 170 186 171 187
rect 169 186 170 187
rect 168 186 169 187
rect 167 186 168 187
rect 165 186 166 187
rect 164 186 165 187
rect 151 186 152 187
rect 150 186 151 187
rect 149 186 150 187
rect 148 186 149 187
rect 147 186 148 187
rect 146 186 147 187
rect 145 186 146 187
rect 144 186 145 187
rect 143 186 144 187
rect 142 186 143 187
rect 141 186 142 187
rect 140 186 141 187
rect 139 186 140 187
rect 138 186 139 187
rect 137 186 138 187
rect 136 186 137 187
rect 135 186 136 187
rect 134 186 135 187
rect 133 186 134 187
rect 132 186 133 187
rect 131 186 132 187
rect 130 186 131 187
rect 129 186 130 187
rect 128 186 129 187
rect 127 186 128 187
rect 126 186 127 187
rect 125 186 126 187
rect 124 186 125 187
rect 123 186 124 187
rect 122 186 123 187
rect 121 186 122 187
rect 120 186 121 187
rect 119 186 120 187
rect 118 186 119 187
rect 117 186 118 187
rect 116 186 117 187
rect 115 186 116 187
rect 114 186 115 187
rect 113 186 114 187
rect 112 186 113 187
rect 111 186 112 187
rect 110 186 111 187
rect 109 186 110 187
rect 108 186 109 187
rect 107 186 108 187
rect 106 186 107 187
rect 105 186 106 187
rect 104 186 105 187
rect 64 186 65 187
rect 63 186 64 187
rect 62 186 63 187
rect 61 186 62 187
rect 31 186 32 187
rect 30 186 31 187
rect 29 186 30 187
rect 28 186 29 187
rect 20 186 21 187
rect 198 187 199 188
rect 197 187 198 188
rect 196 187 197 188
rect 195 187 196 188
rect 194 187 195 188
rect 193 187 194 188
rect 192 187 193 188
rect 191 187 192 188
rect 190 187 191 188
rect 185 187 186 188
rect 184 187 185 188
rect 183 187 184 188
rect 182 187 183 188
rect 181 187 182 188
rect 180 187 181 188
rect 177 187 178 188
rect 176 187 177 188
rect 172 187 173 188
rect 171 187 172 188
rect 170 187 171 188
rect 169 187 170 188
rect 168 187 169 188
rect 167 187 168 188
rect 165 187 166 188
rect 164 187 165 188
rect 151 187 152 188
rect 150 187 151 188
rect 149 187 150 188
rect 148 187 149 188
rect 147 187 148 188
rect 146 187 147 188
rect 145 187 146 188
rect 144 187 145 188
rect 143 187 144 188
rect 142 187 143 188
rect 141 187 142 188
rect 140 187 141 188
rect 139 187 140 188
rect 138 187 139 188
rect 137 187 138 188
rect 136 187 137 188
rect 135 187 136 188
rect 134 187 135 188
rect 133 187 134 188
rect 132 187 133 188
rect 131 187 132 188
rect 130 187 131 188
rect 129 187 130 188
rect 128 187 129 188
rect 127 187 128 188
rect 126 187 127 188
rect 125 187 126 188
rect 124 187 125 188
rect 123 187 124 188
rect 122 187 123 188
rect 121 187 122 188
rect 120 187 121 188
rect 119 187 120 188
rect 118 187 119 188
rect 117 187 118 188
rect 116 187 117 188
rect 115 187 116 188
rect 114 187 115 188
rect 113 187 114 188
rect 112 187 113 188
rect 111 187 112 188
rect 110 187 111 188
rect 109 187 110 188
rect 108 187 109 188
rect 107 187 108 188
rect 106 187 107 188
rect 105 187 106 188
rect 104 187 105 188
rect 80 187 81 188
rect 79 187 80 188
rect 78 187 79 188
rect 77 187 78 188
rect 76 187 77 188
rect 75 187 76 188
rect 74 187 75 188
rect 73 187 74 188
rect 72 187 73 188
rect 71 187 72 188
rect 70 187 71 188
rect 69 187 70 188
rect 68 187 69 188
rect 67 187 68 188
rect 66 187 67 188
rect 65 187 66 188
rect 64 187 65 188
rect 63 187 64 188
rect 62 187 63 188
rect 61 187 62 188
rect 60 187 61 188
rect 59 187 60 188
rect 58 187 59 188
rect 57 187 58 188
rect 56 187 57 188
rect 31 187 32 188
rect 30 187 31 188
rect 29 187 30 188
rect 28 187 29 188
rect 27 187 28 188
rect 21 187 22 188
rect 20 187 21 188
rect 19 187 20 188
rect 198 188 199 189
rect 197 188 198 189
rect 196 188 197 189
rect 195 188 196 189
rect 194 188 195 189
rect 193 188 194 189
rect 192 188 193 189
rect 191 188 192 189
rect 190 188 191 189
rect 185 188 186 189
rect 184 188 185 189
rect 183 188 184 189
rect 182 188 183 189
rect 177 188 178 189
rect 176 188 177 189
rect 172 188 173 189
rect 171 188 172 189
rect 170 188 171 189
rect 169 188 170 189
rect 168 188 169 189
rect 167 188 168 189
rect 165 188 166 189
rect 164 188 165 189
rect 151 188 152 189
rect 150 188 151 189
rect 149 188 150 189
rect 148 188 149 189
rect 147 188 148 189
rect 146 188 147 189
rect 145 188 146 189
rect 144 188 145 189
rect 143 188 144 189
rect 142 188 143 189
rect 141 188 142 189
rect 140 188 141 189
rect 139 188 140 189
rect 138 188 139 189
rect 137 188 138 189
rect 136 188 137 189
rect 135 188 136 189
rect 134 188 135 189
rect 133 188 134 189
rect 132 188 133 189
rect 131 188 132 189
rect 130 188 131 189
rect 129 188 130 189
rect 128 188 129 189
rect 127 188 128 189
rect 126 188 127 189
rect 125 188 126 189
rect 124 188 125 189
rect 123 188 124 189
rect 122 188 123 189
rect 121 188 122 189
rect 120 188 121 189
rect 119 188 120 189
rect 118 188 119 189
rect 117 188 118 189
rect 116 188 117 189
rect 115 188 116 189
rect 114 188 115 189
rect 113 188 114 189
rect 112 188 113 189
rect 111 188 112 189
rect 110 188 111 189
rect 109 188 110 189
rect 108 188 109 189
rect 107 188 108 189
rect 106 188 107 189
rect 105 188 106 189
rect 104 188 105 189
rect 80 188 81 189
rect 79 188 80 189
rect 78 188 79 189
rect 77 188 78 189
rect 76 188 77 189
rect 75 188 76 189
rect 74 188 75 189
rect 73 188 74 189
rect 72 188 73 189
rect 71 188 72 189
rect 70 188 71 189
rect 69 188 70 189
rect 68 188 69 189
rect 67 188 68 189
rect 66 188 67 189
rect 65 188 66 189
rect 64 188 65 189
rect 63 188 64 189
rect 62 188 63 189
rect 61 188 62 189
rect 60 188 61 189
rect 59 188 60 189
rect 58 188 59 189
rect 57 188 58 189
rect 56 188 57 189
rect 55 188 56 189
rect 54 188 55 189
rect 31 188 32 189
rect 30 188 31 189
rect 29 188 30 189
rect 28 188 29 189
rect 27 188 28 189
rect 26 188 27 189
rect 21 188 22 189
rect 20 188 21 189
rect 19 188 20 189
rect 18 188 19 189
rect 185 189 186 190
rect 184 189 185 190
rect 183 189 184 190
rect 182 189 183 190
rect 177 189 178 190
rect 176 189 177 190
rect 175 189 176 190
rect 173 189 174 190
rect 172 189 173 190
rect 171 189 172 190
rect 170 189 171 190
rect 169 189 170 190
rect 168 189 169 190
rect 167 189 168 190
rect 165 189 166 190
rect 164 189 165 190
rect 151 189 152 190
rect 150 189 151 190
rect 149 189 150 190
rect 148 189 149 190
rect 147 189 148 190
rect 146 189 147 190
rect 145 189 146 190
rect 144 189 145 190
rect 143 189 144 190
rect 142 189 143 190
rect 141 189 142 190
rect 140 189 141 190
rect 139 189 140 190
rect 138 189 139 190
rect 137 189 138 190
rect 136 189 137 190
rect 135 189 136 190
rect 134 189 135 190
rect 133 189 134 190
rect 132 189 133 190
rect 131 189 132 190
rect 130 189 131 190
rect 129 189 130 190
rect 128 189 129 190
rect 127 189 128 190
rect 126 189 127 190
rect 125 189 126 190
rect 124 189 125 190
rect 123 189 124 190
rect 122 189 123 190
rect 121 189 122 190
rect 120 189 121 190
rect 119 189 120 190
rect 118 189 119 190
rect 117 189 118 190
rect 116 189 117 190
rect 115 189 116 190
rect 114 189 115 190
rect 113 189 114 190
rect 112 189 113 190
rect 111 189 112 190
rect 110 189 111 190
rect 109 189 110 190
rect 108 189 109 190
rect 107 189 108 190
rect 106 189 107 190
rect 105 189 106 190
rect 104 189 105 190
rect 80 189 81 190
rect 79 189 80 190
rect 78 189 79 190
rect 77 189 78 190
rect 76 189 77 190
rect 75 189 76 190
rect 74 189 75 190
rect 73 189 74 190
rect 72 189 73 190
rect 71 189 72 190
rect 70 189 71 190
rect 69 189 70 190
rect 68 189 69 190
rect 67 189 68 190
rect 66 189 67 190
rect 65 189 66 190
rect 64 189 65 190
rect 63 189 64 190
rect 62 189 63 190
rect 61 189 62 190
rect 60 189 61 190
rect 59 189 60 190
rect 58 189 59 190
rect 57 189 58 190
rect 56 189 57 190
rect 55 189 56 190
rect 54 189 55 190
rect 31 189 32 190
rect 30 189 31 190
rect 29 189 30 190
rect 28 189 29 190
rect 27 189 28 190
rect 26 189 27 190
rect 25 189 26 190
rect 21 189 22 190
rect 20 189 21 190
rect 19 189 20 190
rect 18 189 19 190
rect 17 189 18 190
rect 198 190 199 191
rect 197 190 198 191
rect 196 190 197 191
rect 195 190 196 191
rect 194 190 195 191
rect 185 190 186 191
rect 184 190 185 191
rect 183 190 184 191
rect 182 190 183 191
rect 177 190 178 191
rect 176 190 177 191
rect 175 190 176 191
rect 173 190 174 191
rect 172 190 173 191
rect 171 190 172 191
rect 170 190 171 191
rect 169 190 170 191
rect 168 190 169 191
rect 167 190 168 191
rect 165 190 166 191
rect 164 190 165 191
rect 151 190 152 191
rect 150 190 151 191
rect 149 190 150 191
rect 148 190 149 191
rect 147 190 148 191
rect 146 190 147 191
rect 145 190 146 191
rect 144 190 145 191
rect 143 190 144 191
rect 142 190 143 191
rect 141 190 142 191
rect 140 190 141 191
rect 139 190 140 191
rect 138 190 139 191
rect 137 190 138 191
rect 136 190 137 191
rect 135 190 136 191
rect 134 190 135 191
rect 133 190 134 191
rect 132 190 133 191
rect 131 190 132 191
rect 130 190 131 191
rect 129 190 130 191
rect 128 190 129 191
rect 127 190 128 191
rect 126 190 127 191
rect 125 190 126 191
rect 124 190 125 191
rect 123 190 124 191
rect 122 190 123 191
rect 121 190 122 191
rect 120 190 121 191
rect 119 190 120 191
rect 118 190 119 191
rect 117 190 118 191
rect 116 190 117 191
rect 115 190 116 191
rect 114 190 115 191
rect 113 190 114 191
rect 112 190 113 191
rect 111 190 112 191
rect 110 190 111 191
rect 109 190 110 191
rect 108 190 109 191
rect 107 190 108 191
rect 106 190 107 191
rect 105 190 106 191
rect 104 190 105 191
rect 80 190 81 191
rect 79 190 80 191
rect 78 190 79 191
rect 77 190 78 191
rect 76 190 77 191
rect 75 190 76 191
rect 74 190 75 191
rect 73 190 74 191
rect 72 190 73 191
rect 71 190 72 191
rect 70 190 71 191
rect 69 190 70 191
rect 68 190 69 191
rect 67 190 68 191
rect 66 190 67 191
rect 65 190 66 191
rect 64 190 65 191
rect 63 190 64 191
rect 62 190 63 191
rect 61 190 62 191
rect 60 190 61 191
rect 59 190 60 191
rect 58 190 59 191
rect 57 190 58 191
rect 56 190 57 191
rect 55 190 56 191
rect 54 190 55 191
rect 53 190 54 191
rect 31 190 32 191
rect 30 190 31 191
rect 29 190 30 191
rect 27 190 28 191
rect 26 190 27 191
rect 25 190 26 191
rect 24 190 25 191
rect 19 190 20 191
rect 18 190 19 191
rect 17 190 18 191
rect 198 191 199 192
rect 197 191 198 192
rect 196 191 197 192
rect 195 191 196 192
rect 194 191 195 192
rect 193 191 194 192
rect 185 191 186 192
rect 184 191 185 192
rect 183 191 184 192
rect 182 191 183 192
rect 177 191 178 192
rect 176 191 177 192
rect 175 191 176 192
rect 174 191 175 192
rect 173 191 174 192
rect 172 191 173 192
rect 171 191 172 192
rect 169 191 170 192
rect 168 191 169 192
rect 167 191 168 192
rect 165 191 166 192
rect 164 191 165 192
rect 151 191 152 192
rect 150 191 151 192
rect 149 191 150 192
rect 148 191 149 192
rect 147 191 148 192
rect 146 191 147 192
rect 145 191 146 192
rect 144 191 145 192
rect 143 191 144 192
rect 142 191 143 192
rect 141 191 142 192
rect 140 191 141 192
rect 139 191 140 192
rect 138 191 139 192
rect 137 191 138 192
rect 136 191 137 192
rect 135 191 136 192
rect 134 191 135 192
rect 133 191 134 192
rect 132 191 133 192
rect 131 191 132 192
rect 130 191 131 192
rect 129 191 130 192
rect 128 191 129 192
rect 127 191 128 192
rect 126 191 127 192
rect 125 191 126 192
rect 124 191 125 192
rect 123 191 124 192
rect 122 191 123 192
rect 121 191 122 192
rect 120 191 121 192
rect 119 191 120 192
rect 118 191 119 192
rect 117 191 118 192
rect 116 191 117 192
rect 115 191 116 192
rect 114 191 115 192
rect 113 191 114 192
rect 112 191 113 192
rect 111 191 112 192
rect 110 191 111 192
rect 109 191 110 192
rect 108 191 109 192
rect 107 191 108 192
rect 106 191 107 192
rect 105 191 106 192
rect 104 191 105 192
rect 80 191 81 192
rect 79 191 80 192
rect 78 191 79 192
rect 77 191 78 192
rect 76 191 77 192
rect 75 191 76 192
rect 74 191 75 192
rect 73 191 74 192
rect 72 191 73 192
rect 71 191 72 192
rect 70 191 71 192
rect 69 191 70 192
rect 68 191 69 192
rect 67 191 68 192
rect 66 191 67 192
rect 65 191 66 192
rect 64 191 65 192
rect 63 191 64 192
rect 62 191 63 192
rect 61 191 62 192
rect 60 191 61 192
rect 59 191 60 192
rect 58 191 59 192
rect 57 191 58 192
rect 56 191 57 192
rect 55 191 56 192
rect 54 191 55 192
rect 53 191 54 192
rect 31 191 32 192
rect 30 191 31 192
rect 29 191 30 192
rect 26 191 27 192
rect 25 191 26 192
rect 24 191 25 192
rect 23 191 24 192
rect 19 191 20 192
rect 18 191 19 192
rect 17 191 18 192
rect 199 192 200 193
rect 198 192 199 193
rect 196 192 197 193
rect 194 192 195 193
rect 193 192 194 193
rect 185 192 186 193
rect 184 192 185 193
rect 183 192 184 193
rect 182 192 183 193
rect 177 192 178 193
rect 176 192 177 193
rect 175 192 176 193
rect 174 192 175 193
rect 173 192 174 193
rect 172 192 173 193
rect 171 192 172 193
rect 169 192 170 193
rect 168 192 169 193
rect 167 192 168 193
rect 151 192 152 193
rect 150 192 151 193
rect 149 192 150 193
rect 148 192 149 193
rect 147 192 148 193
rect 146 192 147 193
rect 145 192 146 193
rect 144 192 145 193
rect 143 192 144 193
rect 142 192 143 193
rect 141 192 142 193
rect 140 192 141 193
rect 139 192 140 193
rect 138 192 139 193
rect 137 192 138 193
rect 136 192 137 193
rect 135 192 136 193
rect 134 192 135 193
rect 133 192 134 193
rect 132 192 133 193
rect 131 192 132 193
rect 130 192 131 193
rect 129 192 130 193
rect 128 192 129 193
rect 127 192 128 193
rect 126 192 127 193
rect 125 192 126 193
rect 124 192 125 193
rect 123 192 124 193
rect 122 192 123 193
rect 121 192 122 193
rect 120 192 121 193
rect 119 192 120 193
rect 118 192 119 193
rect 117 192 118 193
rect 116 192 117 193
rect 115 192 116 193
rect 114 192 115 193
rect 113 192 114 193
rect 112 192 113 193
rect 111 192 112 193
rect 110 192 111 193
rect 109 192 110 193
rect 108 192 109 193
rect 107 192 108 193
rect 106 192 107 193
rect 105 192 106 193
rect 104 192 105 193
rect 80 192 81 193
rect 79 192 80 193
rect 78 192 79 193
rect 77 192 78 193
rect 76 192 77 193
rect 75 192 76 193
rect 74 192 75 193
rect 73 192 74 193
rect 72 192 73 193
rect 71 192 72 193
rect 70 192 71 193
rect 69 192 70 193
rect 68 192 69 193
rect 67 192 68 193
rect 66 192 67 193
rect 65 192 66 193
rect 64 192 65 193
rect 63 192 64 193
rect 62 192 63 193
rect 61 192 62 193
rect 60 192 61 193
rect 59 192 60 193
rect 58 192 59 193
rect 57 192 58 193
rect 56 192 57 193
rect 55 192 56 193
rect 54 192 55 193
rect 53 192 54 193
rect 31 192 32 193
rect 30 192 31 193
rect 29 192 30 193
rect 25 192 26 193
rect 24 192 25 193
rect 23 192 24 193
rect 22 192 23 193
rect 19 192 20 193
rect 18 192 19 193
rect 17 192 18 193
rect 199 193 200 194
rect 198 193 199 194
rect 196 193 197 194
rect 195 193 196 194
rect 194 193 195 194
rect 193 193 194 194
rect 185 193 186 194
rect 184 193 185 194
rect 183 193 184 194
rect 182 193 183 194
rect 176 193 177 194
rect 175 193 176 194
rect 174 193 175 194
rect 173 193 174 194
rect 172 193 173 194
rect 169 193 170 194
rect 168 193 169 194
rect 167 193 168 194
rect 151 193 152 194
rect 150 193 151 194
rect 149 193 150 194
rect 148 193 149 194
rect 147 193 148 194
rect 146 193 147 194
rect 145 193 146 194
rect 144 193 145 194
rect 143 193 144 194
rect 142 193 143 194
rect 141 193 142 194
rect 140 193 141 194
rect 139 193 140 194
rect 138 193 139 194
rect 137 193 138 194
rect 136 193 137 194
rect 135 193 136 194
rect 134 193 135 194
rect 133 193 134 194
rect 132 193 133 194
rect 131 193 132 194
rect 130 193 131 194
rect 129 193 130 194
rect 128 193 129 194
rect 127 193 128 194
rect 126 193 127 194
rect 125 193 126 194
rect 124 193 125 194
rect 123 193 124 194
rect 122 193 123 194
rect 121 193 122 194
rect 120 193 121 194
rect 119 193 120 194
rect 118 193 119 194
rect 117 193 118 194
rect 116 193 117 194
rect 115 193 116 194
rect 114 193 115 194
rect 113 193 114 194
rect 112 193 113 194
rect 111 193 112 194
rect 110 193 111 194
rect 109 193 110 194
rect 108 193 109 194
rect 107 193 108 194
rect 106 193 107 194
rect 105 193 106 194
rect 104 193 105 194
rect 64 193 65 194
rect 63 193 64 194
rect 62 193 63 194
rect 61 193 62 194
rect 56 193 57 194
rect 55 193 56 194
rect 54 193 55 194
rect 53 193 54 194
rect 31 193 32 194
rect 30 193 31 194
rect 29 193 30 194
rect 24 193 25 194
rect 23 193 24 194
rect 22 193 23 194
rect 21 193 22 194
rect 20 193 21 194
rect 19 193 20 194
rect 18 193 19 194
rect 17 193 18 194
rect 198 194 199 195
rect 196 194 197 195
rect 195 194 196 195
rect 194 194 195 195
rect 193 194 194 195
rect 185 194 186 195
rect 184 194 185 195
rect 183 194 184 195
rect 182 194 183 195
rect 175 194 176 195
rect 174 194 175 195
rect 173 194 174 195
rect 169 194 170 195
rect 168 194 169 195
rect 167 194 168 195
rect 151 194 152 195
rect 150 194 151 195
rect 149 194 150 195
rect 148 194 149 195
rect 147 194 148 195
rect 146 194 147 195
rect 145 194 146 195
rect 144 194 145 195
rect 143 194 144 195
rect 142 194 143 195
rect 141 194 142 195
rect 140 194 141 195
rect 139 194 140 195
rect 138 194 139 195
rect 137 194 138 195
rect 136 194 137 195
rect 135 194 136 195
rect 134 194 135 195
rect 133 194 134 195
rect 132 194 133 195
rect 131 194 132 195
rect 130 194 131 195
rect 129 194 130 195
rect 128 194 129 195
rect 127 194 128 195
rect 126 194 127 195
rect 125 194 126 195
rect 124 194 125 195
rect 123 194 124 195
rect 122 194 123 195
rect 121 194 122 195
rect 120 194 121 195
rect 119 194 120 195
rect 118 194 119 195
rect 117 194 118 195
rect 116 194 117 195
rect 115 194 116 195
rect 114 194 115 195
rect 113 194 114 195
rect 112 194 113 195
rect 111 194 112 195
rect 110 194 111 195
rect 109 194 110 195
rect 108 194 109 195
rect 107 194 108 195
rect 106 194 107 195
rect 105 194 106 195
rect 104 194 105 195
rect 64 194 65 195
rect 63 194 64 195
rect 62 194 63 195
rect 61 194 62 195
rect 56 194 57 195
rect 55 194 56 195
rect 54 194 55 195
rect 53 194 54 195
rect 30 194 31 195
rect 29 194 30 195
rect 23 194 24 195
rect 22 194 23 195
rect 21 194 22 195
rect 20 194 21 195
rect 19 194 20 195
rect 18 194 19 195
rect 198 195 199 196
rect 196 195 197 196
rect 195 195 196 196
rect 185 195 186 196
rect 184 195 185 196
rect 183 195 184 196
rect 182 195 183 196
rect 168 195 169 196
rect 167 195 168 196
rect 151 195 152 196
rect 150 195 151 196
rect 149 195 150 196
rect 148 195 149 196
rect 147 195 148 196
rect 146 195 147 196
rect 145 195 146 196
rect 144 195 145 196
rect 143 195 144 196
rect 142 195 143 196
rect 141 195 142 196
rect 140 195 141 196
rect 139 195 140 196
rect 138 195 139 196
rect 137 195 138 196
rect 136 195 137 196
rect 135 195 136 196
rect 134 195 135 196
rect 133 195 134 196
rect 132 195 133 196
rect 131 195 132 196
rect 130 195 131 196
rect 129 195 130 196
rect 128 195 129 196
rect 127 195 128 196
rect 126 195 127 196
rect 125 195 126 196
rect 124 195 125 196
rect 123 195 124 196
rect 122 195 123 196
rect 121 195 122 196
rect 120 195 121 196
rect 119 195 120 196
rect 118 195 119 196
rect 117 195 118 196
rect 116 195 117 196
rect 115 195 116 196
rect 114 195 115 196
rect 113 195 114 196
rect 112 195 113 196
rect 111 195 112 196
rect 110 195 111 196
rect 109 195 110 196
rect 108 195 109 196
rect 107 195 108 196
rect 106 195 107 196
rect 105 195 106 196
rect 104 195 105 196
rect 64 195 65 196
rect 63 195 64 196
rect 62 195 63 196
rect 61 195 62 196
rect 56 195 57 196
rect 55 195 56 196
rect 54 195 55 196
rect 53 195 54 196
rect 22 195 23 196
rect 21 195 22 196
rect 20 195 21 196
rect 19 195 20 196
rect 197 196 198 197
rect 196 196 197 197
rect 195 196 196 197
rect 185 196 186 197
rect 184 196 185 197
rect 183 196 184 197
rect 182 196 183 197
rect 151 196 152 197
rect 150 196 151 197
rect 149 196 150 197
rect 148 196 149 197
rect 147 196 148 197
rect 146 196 147 197
rect 145 196 146 197
rect 144 196 145 197
rect 143 196 144 197
rect 142 196 143 197
rect 141 196 142 197
rect 140 196 141 197
rect 139 196 140 197
rect 138 196 139 197
rect 137 196 138 197
rect 136 196 137 197
rect 135 196 136 197
rect 134 196 135 197
rect 133 196 134 197
rect 132 196 133 197
rect 131 196 132 197
rect 130 196 131 197
rect 129 196 130 197
rect 128 196 129 197
rect 127 196 128 197
rect 126 196 127 197
rect 125 196 126 197
rect 124 196 125 197
rect 123 196 124 197
rect 122 196 123 197
rect 121 196 122 197
rect 120 196 121 197
rect 119 196 120 197
rect 118 196 119 197
rect 117 196 118 197
rect 116 196 117 197
rect 115 196 116 197
rect 114 196 115 197
rect 113 196 114 197
rect 112 196 113 197
rect 111 196 112 197
rect 110 196 111 197
rect 109 196 110 197
rect 108 196 109 197
rect 107 196 108 197
rect 106 196 107 197
rect 105 196 106 197
rect 104 196 105 197
rect 64 196 65 197
rect 63 196 64 197
rect 62 196 63 197
rect 61 196 62 197
rect 56 196 57 197
rect 55 196 56 197
rect 54 196 55 197
rect 53 196 54 197
rect 198 197 199 198
rect 197 197 198 198
rect 196 197 197 198
rect 195 197 196 198
rect 194 197 195 198
rect 193 197 194 198
rect 185 197 186 198
rect 184 197 185 198
rect 183 197 184 198
rect 182 197 183 198
rect 151 197 152 198
rect 150 197 151 198
rect 149 197 150 198
rect 148 197 149 198
rect 147 197 148 198
rect 146 197 147 198
rect 145 197 146 198
rect 144 197 145 198
rect 143 197 144 198
rect 142 197 143 198
rect 141 197 142 198
rect 140 197 141 198
rect 139 197 140 198
rect 138 197 139 198
rect 137 197 138 198
rect 136 197 137 198
rect 135 197 136 198
rect 134 197 135 198
rect 133 197 134 198
rect 132 197 133 198
rect 131 197 132 198
rect 130 197 131 198
rect 129 197 130 198
rect 128 197 129 198
rect 127 197 128 198
rect 126 197 127 198
rect 125 197 126 198
rect 124 197 125 198
rect 123 197 124 198
rect 122 197 123 198
rect 121 197 122 198
rect 120 197 121 198
rect 119 197 120 198
rect 118 197 119 198
rect 117 197 118 198
rect 116 197 117 198
rect 115 197 116 198
rect 114 197 115 198
rect 113 197 114 198
rect 112 197 113 198
rect 111 197 112 198
rect 110 197 111 198
rect 109 197 110 198
rect 108 197 109 198
rect 107 197 108 198
rect 106 197 107 198
rect 105 197 106 198
rect 104 197 105 198
rect 55 197 56 198
rect 54 197 55 198
rect 53 197 54 198
rect 29 197 30 198
rect 28 197 29 198
rect 27 197 28 198
rect 26 197 27 198
rect 25 197 26 198
rect 24 197 25 198
rect 23 197 24 198
rect 198 198 199 199
rect 197 198 198 199
rect 194 198 195 199
rect 193 198 194 199
rect 185 198 186 199
rect 184 198 185 199
rect 183 198 184 199
rect 182 198 183 199
rect 179 198 180 199
rect 178 198 179 199
rect 177 198 178 199
rect 176 198 177 199
rect 175 198 176 199
rect 174 198 175 199
rect 173 198 174 199
rect 172 198 173 199
rect 171 198 172 199
rect 170 198 171 199
rect 169 198 170 199
rect 168 198 169 199
rect 167 198 168 199
rect 166 198 167 199
rect 165 198 166 199
rect 164 198 165 199
rect 151 198 152 199
rect 150 198 151 199
rect 149 198 150 199
rect 148 198 149 199
rect 147 198 148 199
rect 146 198 147 199
rect 145 198 146 199
rect 144 198 145 199
rect 143 198 144 199
rect 142 198 143 199
rect 141 198 142 199
rect 140 198 141 199
rect 139 198 140 199
rect 138 198 139 199
rect 137 198 138 199
rect 136 198 137 199
rect 135 198 136 199
rect 134 198 135 199
rect 133 198 134 199
rect 132 198 133 199
rect 131 198 132 199
rect 130 198 131 199
rect 129 198 130 199
rect 128 198 129 199
rect 127 198 128 199
rect 126 198 127 199
rect 125 198 126 199
rect 124 198 125 199
rect 123 198 124 199
rect 122 198 123 199
rect 121 198 122 199
rect 120 198 121 199
rect 119 198 120 199
rect 118 198 119 199
rect 117 198 118 199
rect 116 198 117 199
rect 115 198 116 199
rect 114 198 115 199
rect 113 198 114 199
rect 112 198 113 199
rect 111 198 112 199
rect 110 198 111 199
rect 109 198 110 199
rect 108 198 109 199
rect 107 198 108 199
rect 106 198 107 199
rect 105 198 106 199
rect 104 198 105 199
rect 30 198 31 199
rect 29 198 30 199
rect 28 198 29 199
rect 27 198 28 199
rect 26 198 27 199
rect 25 198 26 199
rect 24 198 25 199
rect 23 198 24 199
rect 22 198 23 199
rect 21 198 22 199
rect 20 198 21 199
rect 199 199 200 200
rect 198 199 199 200
rect 194 199 195 200
rect 193 199 194 200
rect 185 199 186 200
rect 184 199 185 200
rect 183 199 184 200
rect 182 199 183 200
rect 179 199 180 200
rect 178 199 179 200
rect 177 199 178 200
rect 176 199 177 200
rect 175 199 176 200
rect 174 199 175 200
rect 173 199 174 200
rect 172 199 173 200
rect 171 199 172 200
rect 170 199 171 200
rect 169 199 170 200
rect 168 199 169 200
rect 167 199 168 200
rect 166 199 167 200
rect 165 199 166 200
rect 164 199 165 200
rect 151 199 152 200
rect 150 199 151 200
rect 149 199 150 200
rect 148 199 149 200
rect 147 199 148 200
rect 146 199 147 200
rect 145 199 146 200
rect 144 199 145 200
rect 143 199 144 200
rect 142 199 143 200
rect 141 199 142 200
rect 140 199 141 200
rect 139 199 140 200
rect 138 199 139 200
rect 137 199 138 200
rect 136 199 137 200
rect 135 199 136 200
rect 134 199 135 200
rect 133 199 134 200
rect 132 199 133 200
rect 131 199 132 200
rect 130 199 131 200
rect 129 199 130 200
rect 128 199 129 200
rect 127 199 128 200
rect 126 199 127 200
rect 125 199 126 200
rect 124 199 125 200
rect 123 199 124 200
rect 122 199 123 200
rect 121 199 122 200
rect 120 199 121 200
rect 119 199 120 200
rect 118 199 119 200
rect 117 199 118 200
rect 116 199 117 200
rect 115 199 116 200
rect 114 199 115 200
rect 113 199 114 200
rect 112 199 113 200
rect 111 199 112 200
rect 110 199 111 200
rect 109 199 110 200
rect 108 199 109 200
rect 107 199 108 200
rect 106 199 107 200
rect 105 199 106 200
rect 104 199 105 200
rect 80 199 81 200
rect 79 199 80 200
rect 78 199 79 200
rect 77 199 78 200
rect 76 199 77 200
rect 75 199 76 200
rect 74 199 75 200
rect 73 199 74 200
rect 72 199 73 200
rect 71 199 72 200
rect 70 199 71 200
rect 69 199 70 200
rect 68 199 69 200
rect 67 199 68 200
rect 66 199 67 200
rect 65 199 66 200
rect 64 199 65 200
rect 63 199 64 200
rect 62 199 63 200
rect 61 199 62 200
rect 57 199 58 200
rect 56 199 57 200
rect 55 199 56 200
rect 54 199 55 200
rect 53 199 54 200
rect 31 199 32 200
rect 30 199 31 200
rect 29 199 30 200
rect 28 199 29 200
rect 27 199 28 200
rect 26 199 27 200
rect 25 199 26 200
rect 24 199 25 200
rect 23 199 24 200
rect 22 199 23 200
rect 21 199 22 200
rect 20 199 21 200
rect 19 199 20 200
rect 199 200 200 201
rect 198 200 199 201
rect 194 200 195 201
rect 193 200 194 201
rect 185 200 186 201
rect 184 200 185 201
rect 183 200 184 201
rect 182 200 183 201
rect 179 200 180 201
rect 178 200 179 201
rect 177 200 178 201
rect 176 200 177 201
rect 175 200 176 201
rect 174 200 175 201
rect 173 200 174 201
rect 172 200 173 201
rect 171 200 172 201
rect 170 200 171 201
rect 169 200 170 201
rect 168 200 169 201
rect 167 200 168 201
rect 166 200 167 201
rect 165 200 166 201
rect 164 200 165 201
rect 151 200 152 201
rect 150 200 151 201
rect 149 200 150 201
rect 148 200 149 201
rect 147 200 148 201
rect 146 200 147 201
rect 145 200 146 201
rect 144 200 145 201
rect 143 200 144 201
rect 142 200 143 201
rect 141 200 142 201
rect 140 200 141 201
rect 139 200 140 201
rect 138 200 139 201
rect 137 200 138 201
rect 136 200 137 201
rect 135 200 136 201
rect 134 200 135 201
rect 133 200 134 201
rect 132 200 133 201
rect 131 200 132 201
rect 130 200 131 201
rect 129 200 130 201
rect 128 200 129 201
rect 127 200 128 201
rect 126 200 127 201
rect 125 200 126 201
rect 124 200 125 201
rect 123 200 124 201
rect 122 200 123 201
rect 121 200 122 201
rect 120 200 121 201
rect 119 200 120 201
rect 118 200 119 201
rect 117 200 118 201
rect 116 200 117 201
rect 115 200 116 201
rect 114 200 115 201
rect 113 200 114 201
rect 112 200 113 201
rect 111 200 112 201
rect 110 200 111 201
rect 109 200 110 201
rect 108 200 109 201
rect 107 200 108 201
rect 106 200 107 201
rect 105 200 106 201
rect 104 200 105 201
rect 80 200 81 201
rect 79 200 80 201
rect 78 200 79 201
rect 77 200 78 201
rect 76 200 77 201
rect 75 200 76 201
rect 74 200 75 201
rect 73 200 74 201
rect 72 200 73 201
rect 71 200 72 201
rect 70 200 71 201
rect 69 200 70 201
rect 68 200 69 201
rect 67 200 68 201
rect 66 200 67 201
rect 65 200 66 201
rect 64 200 65 201
rect 63 200 64 201
rect 62 200 63 201
rect 61 200 62 201
rect 57 200 58 201
rect 56 200 57 201
rect 55 200 56 201
rect 54 200 55 201
rect 53 200 54 201
rect 31 200 32 201
rect 30 200 31 201
rect 29 200 30 201
rect 23 200 24 201
rect 22 200 23 201
rect 21 200 22 201
rect 20 200 21 201
rect 19 200 20 201
rect 18 200 19 201
rect 193 201 194 202
rect 184 201 185 202
rect 183 201 184 202
rect 172 201 173 202
rect 171 201 172 202
rect 170 201 171 202
rect 151 201 152 202
rect 150 201 151 202
rect 149 201 150 202
rect 148 201 149 202
rect 147 201 148 202
rect 146 201 147 202
rect 145 201 146 202
rect 144 201 145 202
rect 143 201 144 202
rect 142 201 143 202
rect 141 201 142 202
rect 139 201 140 202
rect 138 201 139 202
rect 137 201 138 202
rect 136 201 137 202
rect 135 201 136 202
rect 134 201 135 202
rect 133 201 134 202
rect 132 201 133 202
rect 131 201 132 202
rect 130 201 131 202
rect 129 201 130 202
rect 128 201 129 202
rect 127 201 128 202
rect 126 201 127 202
rect 125 201 126 202
rect 124 201 125 202
rect 123 201 124 202
rect 122 201 123 202
rect 120 201 121 202
rect 119 201 120 202
rect 118 201 119 202
rect 117 201 118 202
rect 116 201 117 202
rect 114 201 115 202
rect 113 201 114 202
rect 112 201 113 202
rect 111 201 112 202
rect 110 201 111 202
rect 109 201 110 202
rect 108 201 109 202
rect 107 201 108 202
rect 106 201 107 202
rect 105 201 106 202
rect 104 201 105 202
rect 80 201 81 202
rect 79 201 80 202
rect 78 201 79 202
rect 77 201 78 202
rect 76 201 77 202
rect 75 201 76 202
rect 74 201 75 202
rect 73 201 74 202
rect 72 201 73 202
rect 71 201 72 202
rect 70 201 71 202
rect 69 201 70 202
rect 68 201 69 202
rect 67 201 68 202
rect 66 201 67 202
rect 65 201 66 202
rect 64 201 65 202
rect 63 201 64 202
rect 62 201 63 202
rect 61 201 62 202
rect 57 201 58 202
rect 56 201 57 202
rect 55 201 56 202
rect 54 201 55 202
rect 53 201 54 202
rect 31 201 32 202
rect 30 201 31 202
rect 29 201 30 202
rect 20 201 21 202
rect 19 201 20 202
rect 18 201 19 202
rect 17 201 18 202
rect 197 202 198 203
rect 196 202 197 203
rect 195 202 196 203
rect 194 202 195 203
rect 193 202 194 203
rect 192 202 193 203
rect 172 202 173 203
rect 171 202 172 203
rect 170 202 171 203
rect 151 202 152 203
rect 150 202 151 203
rect 149 202 150 203
rect 148 202 149 203
rect 147 202 148 203
rect 146 202 147 203
rect 145 202 146 203
rect 144 202 145 203
rect 143 202 144 203
rect 142 202 143 203
rect 133 202 134 203
rect 132 202 133 203
rect 131 202 132 203
rect 130 202 131 203
rect 129 202 130 203
rect 128 202 129 203
rect 127 202 128 203
rect 126 202 127 203
rect 125 202 126 203
rect 124 202 125 203
rect 123 202 124 203
rect 114 202 115 203
rect 113 202 114 203
rect 112 202 113 203
rect 111 202 112 203
rect 110 202 111 203
rect 109 202 110 203
rect 108 202 109 203
rect 107 202 108 203
rect 106 202 107 203
rect 105 202 106 203
rect 104 202 105 203
rect 80 202 81 203
rect 79 202 80 203
rect 78 202 79 203
rect 77 202 78 203
rect 76 202 77 203
rect 75 202 76 203
rect 74 202 75 203
rect 73 202 74 203
rect 72 202 73 203
rect 71 202 72 203
rect 70 202 71 203
rect 69 202 70 203
rect 68 202 69 203
rect 67 202 68 203
rect 66 202 67 203
rect 65 202 66 203
rect 64 202 65 203
rect 63 202 64 203
rect 62 202 63 203
rect 61 202 62 203
rect 57 202 58 203
rect 56 202 57 203
rect 55 202 56 203
rect 54 202 55 203
rect 53 202 54 203
rect 31 202 32 203
rect 30 202 31 203
rect 29 202 30 203
rect 19 202 20 203
rect 18 202 19 203
rect 17 202 18 203
rect 198 203 199 204
rect 197 203 198 204
rect 196 203 197 204
rect 195 203 196 204
rect 194 203 195 204
rect 193 203 194 204
rect 192 203 193 204
rect 191 203 192 204
rect 172 203 173 204
rect 171 203 172 204
rect 170 203 171 204
rect 151 203 152 204
rect 150 203 151 204
rect 149 203 150 204
rect 148 203 149 204
rect 147 203 148 204
rect 146 203 147 204
rect 145 203 146 204
rect 144 203 145 204
rect 143 203 144 204
rect 142 203 143 204
rect 132 203 133 204
rect 131 203 132 204
rect 130 203 131 204
rect 129 203 130 204
rect 128 203 129 204
rect 127 203 128 204
rect 126 203 127 204
rect 125 203 126 204
rect 124 203 125 204
rect 123 203 124 204
rect 114 203 115 204
rect 113 203 114 204
rect 112 203 113 204
rect 111 203 112 204
rect 110 203 111 204
rect 109 203 110 204
rect 108 203 109 204
rect 107 203 108 204
rect 106 203 107 204
rect 105 203 106 204
rect 104 203 105 204
rect 80 203 81 204
rect 79 203 80 204
rect 78 203 79 204
rect 77 203 78 204
rect 76 203 77 204
rect 75 203 76 204
rect 74 203 75 204
rect 73 203 74 204
rect 72 203 73 204
rect 71 203 72 204
rect 70 203 71 204
rect 69 203 70 204
rect 68 203 69 204
rect 67 203 68 204
rect 66 203 67 204
rect 65 203 66 204
rect 64 203 65 204
rect 63 203 64 204
rect 62 203 63 204
rect 61 203 62 204
rect 57 203 58 204
rect 56 203 57 204
rect 55 203 56 204
rect 54 203 55 204
rect 53 203 54 204
rect 30 203 31 204
rect 29 203 30 204
rect 28 203 29 204
rect 27 203 28 204
rect 19 203 20 204
rect 18 203 19 204
rect 17 203 18 204
rect 198 204 199 205
rect 197 204 198 205
rect 196 204 197 205
rect 195 204 196 205
rect 194 204 195 205
rect 193 204 194 205
rect 192 204 193 205
rect 191 204 192 205
rect 151 204 152 205
rect 150 204 151 205
rect 149 204 150 205
rect 148 204 149 205
rect 147 204 148 205
rect 146 204 147 205
rect 145 204 146 205
rect 144 204 145 205
rect 143 204 144 205
rect 142 204 143 205
rect 132 204 133 205
rect 131 204 132 205
rect 130 204 131 205
rect 129 204 130 205
rect 128 204 129 205
rect 127 204 128 205
rect 126 204 127 205
rect 125 204 126 205
rect 124 204 125 205
rect 123 204 124 205
rect 114 204 115 205
rect 113 204 114 205
rect 112 204 113 205
rect 111 204 112 205
rect 110 204 111 205
rect 109 204 110 205
rect 108 204 109 205
rect 107 204 108 205
rect 106 204 107 205
rect 105 204 106 205
rect 104 204 105 205
rect 80 204 81 205
rect 79 204 80 205
rect 78 204 79 205
rect 77 204 78 205
rect 76 204 77 205
rect 75 204 76 205
rect 74 204 75 205
rect 73 204 74 205
rect 72 204 73 205
rect 71 204 72 205
rect 70 204 71 205
rect 69 204 70 205
rect 68 204 69 205
rect 67 204 68 205
rect 66 204 67 205
rect 65 204 66 205
rect 64 204 65 205
rect 63 204 64 205
rect 62 204 63 205
rect 61 204 62 205
rect 57 204 58 205
rect 56 204 57 205
rect 55 204 56 205
rect 54 204 55 205
rect 53 204 54 205
rect 30 204 31 205
rect 29 204 30 205
rect 28 204 29 205
rect 27 204 28 205
rect 26 204 27 205
rect 25 204 26 205
rect 24 204 25 205
rect 23 204 24 205
rect 19 204 20 205
rect 18 204 19 205
rect 17 204 18 205
rect 198 205 199 206
rect 193 205 194 206
rect 151 205 152 206
rect 150 205 151 206
rect 149 205 150 206
rect 148 205 149 206
rect 147 205 148 206
rect 146 205 147 206
rect 145 205 146 206
rect 144 205 145 206
rect 143 205 144 206
rect 142 205 143 206
rect 132 205 133 206
rect 131 205 132 206
rect 130 205 131 206
rect 129 205 130 206
rect 128 205 129 206
rect 127 205 128 206
rect 126 205 127 206
rect 125 205 126 206
rect 124 205 125 206
rect 123 205 124 206
rect 114 205 115 206
rect 113 205 114 206
rect 112 205 113 206
rect 111 205 112 206
rect 110 205 111 206
rect 109 205 110 206
rect 108 205 109 206
rect 107 205 108 206
rect 106 205 107 206
rect 105 205 106 206
rect 104 205 105 206
rect 29 205 30 206
rect 28 205 29 206
rect 27 205 28 206
rect 26 205 27 206
rect 25 205 26 206
rect 24 205 25 206
rect 23 205 24 206
rect 22 205 23 206
rect 21 205 22 206
rect 20 205 21 206
rect 19 205 20 206
rect 18 205 19 206
rect 17 205 18 206
rect 198 206 199 207
rect 197 206 198 207
rect 196 206 197 207
rect 195 206 196 207
rect 194 206 195 207
rect 193 206 194 207
rect 151 206 152 207
rect 150 206 151 207
rect 149 206 150 207
rect 148 206 149 207
rect 147 206 148 207
rect 146 206 147 207
rect 145 206 146 207
rect 144 206 145 207
rect 143 206 144 207
rect 142 206 143 207
rect 132 206 133 207
rect 131 206 132 207
rect 130 206 131 207
rect 129 206 130 207
rect 128 206 129 207
rect 127 206 128 207
rect 126 206 127 207
rect 125 206 126 207
rect 124 206 125 207
rect 123 206 124 207
rect 114 206 115 207
rect 113 206 114 207
rect 112 206 113 207
rect 111 206 112 207
rect 110 206 111 207
rect 109 206 110 207
rect 108 206 109 207
rect 107 206 108 207
rect 106 206 107 207
rect 105 206 106 207
rect 104 206 105 207
rect 27 206 28 207
rect 26 206 27 207
rect 25 206 26 207
rect 24 206 25 207
rect 23 206 24 207
rect 22 206 23 207
rect 21 206 22 207
rect 20 206 21 207
rect 19 206 20 207
rect 18 206 19 207
rect 199 207 200 208
rect 198 207 199 208
rect 197 207 198 208
rect 196 207 197 208
rect 195 207 196 208
rect 194 207 195 208
rect 193 207 194 208
rect 151 207 152 208
rect 150 207 151 208
rect 149 207 150 208
rect 148 207 149 208
rect 147 207 148 208
rect 146 207 147 208
rect 145 207 146 208
rect 144 207 145 208
rect 143 207 144 208
rect 142 207 143 208
rect 132 207 133 208
rect 131 207 132 208
rect 130 207 131 208
rect 129 207 130 208
rect 128 207 129 208
rect 127 207 128 208
rect 126 207 127 208
rect 125 207 126 208
rect 124 207 125 208
rect 123 207 124 208
rect 114 207 115 208
rect 113 207 114 208
rect 112 207 113 208
rect 111 207 112 208
rect 110 207 111 208
rect 109 207 110 208
rect 108 207 109 208
rect 107 207 108 208
rect 106 207 107 208
rect 105 207 106 208
rect 104 207 105 208
rect 24 207 25 208
rect 23 207 24 208
rect 22 207 23 208
rect 21 207 22 208
rect 20 207 21 208
rect 198 208 199 209
rect 197 208 198 209
rect 196 208 197 209
rect 195 208 196 209
rect 194 208 195 209
rect 193 208 194 209
rect 151 208 152 209
rect 150 208 151 209
rect 149 208 150 209
rect 148 208 149 209
rect 147 208 148 209
rect 146 208 147 209
rect 145 208 146 209
rect 144 208 145 209
rect 143 208 144 209
rect 142 208 143 209
rect 132 208 133 209
rect 131 208 132 209
rect 130 208 131 209
rect 129 208 130 209
rect 128 208 129 209
rect 127 208 128 209
rect 126 208 127 209
rect 125 208 126 209
rect 124 208 125 209
rect 123 208 124 209
rect 114 208 115 209
rect 113 208 114 209
rect 112 208 113 209
rect 111 208 112 209
rect 110 208 111 209
rect 109 208 110 209
rect 108 208 109 209
rect 107 208 108 209
rect 106 208 107 209
rect 105 208 106 209
rect 104 208 105 209
rect 194 209 195 210
rect 193 209 194 210
rect 151 209 152 210
rect 150 209 151 210
rect 149 209 150 210
rect 148 209 149 210
rect 147 209 148 210
rect 146 209 147 210
rect 145 209 146 210
rect 144 209 145 210
rect 143 209 144 210
rect 142 209 143 210
rect 132 209 133 210
rect 131 209 132 210
rect 130 209 131 210
rect 129 209 130 210
rect 128 209 129 210
rect 127 209 128 210
rect 126 209 127 210
rect 125 209 126 210
rect 124 209 125 210
rect 123 209 124 210
rect 114 209 115 210
rect 113 209 114 210
rect 112 209 113 210
rect 111 209 112 210
rect 110 209 111 210
rect 109 209 110 210
rect 108 209 109 210
rect 107 209 108 210
rect 106 209 107 210
rect 105 209 106 210
rect 104 209 105 210
rect 31 209 32 210
rect 30 209 31 210
rect 29 209 30 210
rect 197 210 198 211
rect 196 210 197 211
rect 195 210 196 211
rect 194 210 195 211
rect 193 210 194 211
rect 151 210 152 211
rect 150 210 151 211
rect 149 210 150 211
rect 148 210 149 211
rect 147 210 148 211
rect 146 210 147 211
rect 145 210 146 211
rect 144 210 145 211
rect 143 210 144 211
rect 142 210 143 211
rect 132 210 133 211
rect 131 210 132 211
rect 130 210 131 211
rect 129 210 130 211
rect 128 210 129 211
rect 127 210 128 211
rect 126 210 127 211
rect 125 210 126 211
rect 124 210 125 211
rect 123 210 124 211
rect 114 210 115 211
rect 113 210 114 211
rect 112 210 113 211
rect 111 210 112 211
rect 110 210 111 211
rect 109 210 110 211
rect 108 210 109 211
rect 107 210 108 211
rect 106 210 107 211
rect 105 210 106 211
rect 104 210 105 211
rect 80 210 81 211
rect 79 210 80 211
rect 78 210 79 211
rect 77 210 78 211
rect 76 210 77 211
rect 75 210 76 211
rect 74 210 75 211
rect 73 210 74 211
rect 72 210 73 211
rect 71 210 72 211
rect 70 210 71 211
rect 69 210 70 211
rect 68 210 69 211
rect 67 210 68 211
rect 66 210 67 211
rect 65 210 66 211
rect 64 210 65 211
rect 63 210 64 211
rect 62 210 63 211
rect 61 210 62 211
rect 31 210 32 211
rect 30 210 31 211
rect 29 210 30 211
rect 28 210 29 211
rect 21 210 22 211
rect 20 210 21 211
rect 198 211 199 212
rect 197 211 198 212
rect 196 211 197 212
rect 195 211 196 212
rect 194 211 195 212
rect 151 211 152 212
rect 150 211 151 212
rect 149 211 150 212
rect 148 211 149 212
rect 147 211 148 212
rect 146 211 147 212
rect 145 211 146 212
rect 144 211 145 212
rect 143 211 144 212
rect 142 211 143 212
rect 132 211 133 212
rect 131 211 132 212
rect 130 211 131 212
rect 129 211 130 212
rect 128 211 129 212
rect 127 211 128 212
rect 126 211 127 212
rect 125 211 126 212
rect 124 211 125 212
rect 123 211 124 212
rect 114 211 115 212
rect 113 211 114 212
rect 112 211 113 212
rect 111 211 112 212
rect 110 211 111 212
rect 109 211 110 212
rect 108 211 109 212
rect 107 211 108 212
rect 106 211 107 212
rect 105 211 106 212
rect 104 211 105 212
rect 80 211 81 212
rect 79 211 80 212
rect 78 211 79 212
rect 77 211 78 212
rect 76 211 77 212
rect 75 211 76 212
rect 74 211 75 212
rect 73 211 74 212
rect 72 211 73 212
rect 71 211 72 212
rect 70 211 71 212
rect 69 211 70 212
rect 68 211 69 212
rect 67 211 68 212
rect 66 211 67 212
rect 65 211 66 212
rect 64 211 65 212
rect 63 211 64 212
rect 62 211 63 212
rect 61 211 62 212
rect 31 211 32 212
rect 30 211 31 212
rect 29 211 30 212
rect 28 211 29 212
rect 27 211 28 212
rect 21 211 22 212
rect 20 211 21 212
rect 19 211 20 212
rect 18 211 19 212
rect 198 212 199 213
rect 197 212 198 213
rect 196 212 197 213
rect 195 212 196 213
rect 194 212 195 213
rect 193 212 194 213
rect 151 212 152 213
rect 150 212 151 213
rect 149 212 150 213
rect 148 212 149 213
rect 147 212 148 213
rect 146 212 147 213
rect 145 212 146 213
rect 144 212 145 213
rect 143 212 144 213
rect 142 212 143 213
rect 132 212 133 213
rect 131 212 132 213
rect 130 212 131 213
rect 129 212 130 213
rect 128 212 129 213
rect 127 212 128 213
rect 126 212 127 213
rect 125 212 126 213
rect 124 212 125 213
rect 123 212 124 213
rect 114 212 115 213
rect 113 212 114 213
rect 112 212 113 213
rect 111 212 112 213
rect 110 212 111 213
rect 109 212 110 213
rect 108 212 109 213
rect 107 212 108 213
rect 106 212 107 213
rect 105 212 106 213
rect 104 212 105 213
rect 80 212 81 213
rect 79 212 80 213
rect 78 212 79 213
rect 77 212 78 213
rect 76 212 77 213
rect 75 212 76 213
rect 74 212 75 213
rect 73 212 74 213
rect 72 212 73 213
rect 71 212 72 213
rect 70 212 71 213
rect 69 212 70 213
rect 68 212 69 213
rect 67 212 68 213
rect 66 212 67 213
rect 65 212 66 213
rect 64 212 65 213
rect 63 212 64 213
rect 62 212 63 213
rect 61 212 62 213
rect 31 212 32 213
rect 30 212 31 213
rect 29 212 30 213
rect 28 212 29 213
rect 27 212 28 213
rect 26 212 27 213
rect 21 212 22 213
rect 20 212 21 213
rect 19 212 20 213
rect 18 212 19 213
rect 17 212 18 213
rect 199 213 200 214
rect 198 213 199 214
rect 194 213 195 214
rect 193 213 194 214
rect 173 213 174 214
rect 151 213 152 214
rect 150 213 151 214
rect 149 213 150 214
rect 148 213 149 214
rect 147 213 148 214
rect 146 213 147 214
rect 145 213 146 214
rect 144 213 145 214
rect 143 213 144 214
rect 142 213 143 214
rect 132 213 133 214
rect 131 213 132 214
rect 130 213 131 214
rect 129 213 130 214
rect 128 213 129 214
rect 127 213 128 214
rect 126 213 127 214
rect 125 213 126 214
rect 124 213 125 214
rect 123 213 124 214
rect 114 213 115 214
rect 113 213 114 214
rect 112 213 113 214
rect 111 213 112 214
rect 110 213 111 214
rect 109 213 110 214
rect 108 213 109 214
rect 107 213 108 214
rect 106 213 107 214
rect 105 213 106 214
rect 104 213 105 214
rect 80 213 81 214
rect 79 213 80 214
rect 78 213 79 214
rect 77 213 78 214
rect 76 213 77 214
rect 75 213 76 214
rect 74 213 75 214
rect 73 213 74 214
rect 72 213 73 214
rect 71 213 72 214
rect 70 213 71 214
rect 69 213 70 214
rect 68 213 69 214
rect 67 213 68 214
rect 66 213 67 214
rect 65 213 66 214
rect 64 213 65 214
rect 63 213 64 214
rect 62 213 63 214
rect 61 213 62 214
rect 31 213 32 214
rect 30 213 31 214
rect 29 213 30 214
rect 28 213 29 214
rect 27 213 28 214
rect 26 213 27 214
rect 25 213 26 214
rect 20 213 21 214
rect 19 213 20 214
rect 18 213 19 214
rect 17 213 18 214
rect 199 214 200 215
rect 198 214 199 215
rect 194 214 195 215
rect 193 214 194 215
rect 175 214 176 215
rect 174 214 175 215
rect 173 214 174 215
rect 172 214 173 215
rect 151 214 152 215
rect 150 214 151 215
rect 149 214 150 215
rect 148 214 149 215
rect 147 214 148 215
rect 146 214 147 215
rect 145 214 146 215
rect 144 214 145 215
rect 143 214 144 215
rect 142 214 143 215
rect 132 214 133 215
rect 131 214 132 215
rect 130 214 131 215
rect 129 214 130 215
rect 128 214 129 215
rect 127 214 128 215
rect 126 214 127 215
rect 125 214 126 215
rect 124 214 125 215
rect 123 214 124 215
rect 114 214 115 215
rect 113 214 114 215
rect 112 214 113 215
rect 111 214 112 215
rect 110 214 111 215
rect 109 214 110 215
rect 108 214 109 215
rect 107 214 108 215
rect 106 214 107 215
rect 105 214 106 215
rect 104 214 105 215
rect 80 214 81 215
rect 79 214 80 215
rect 78 214 79 215
rect 77 214 78 215
rect 76 214 77 215
rect 75 214 76 215
rect 74 214 75 215
rect 73 214 74 215
rect 72 214 73 215
rect 71 214 72 215
rect 70 214 71 215
rect 69 214 70 215
rect 68 214 69 215
rect 67 214 68 215
rect 66 214 67 215
rect 65 214 66 215
rect 64 214 65 215
rect 63 214 64 215
rect 62 214 63 215
rect 61 214 62 215
rect 31 214 32 215
rect 30 214 31 215
rect 29 214 30 215
rect 27 214 28 215
rect 26 214 27 215
rect 25 214 26 215
rect 24 214 25 215
rect 19 214 20 215
rect 18 214 19 215
rect 17 214 18 215
rect 198 215 199 216
rect 197 215 198 216
rect 196 215 197 216
rect 195 215 196 216
rect 194 215 195 216
rect 193 215 194 216
rect 175 215 176 216
rect 174 215 175 216
rect 173 215 174 216
rect 172 215 173 216
rect 151 215 152 216
rect 150 215 151 216
rect 149 215 150 216
rect 148 215 149 216
rect 147 215 148 216
rect 146 215 147 216
rect 145 215 146 216
rect 144 215 145 216
rect 143 215 144 216
rect 142 215 143 216
rect 132 215 133 216
rect 131 215 132 216
rect 130 215 131 216
rect 129 215 130 216
rect 128 215 129 216
rect 127 215 128 216
rect 126 215 127 216
rect 125 215 126 216
rect 124 215 125 216
rect 123 215 124 216
rect 114 215 115 216
rect 113 215 114 216
rect 112 215 113 216
rect 111 215 112 216
rect 110 215 111 216
rect 109 215 110 216
rect 108 215 109 216
rect 107 215 108 216
rect 106 215 107 216
rect 105 215 106 216
rect 104 215 105 216
rect 68 215 69 216
rect 67 215 68 216
rect 66 215 67 216
rect 65 215 66 216
rect 64 215 65 216
rect 63 215 64 216
rect 62 215 63 216
rect 31 215 32 216
rect 30 215 31 216
rect 29 215 30 216
rect 26 215 27 216
rect 25 215 26 216
rect 24 215 25 216
rect 23 215 24 216
rect 19 215 20 216
rect 18 215 19 216
rect 17 215 18 216
rect 198 216 199 217
rect 197 216 198 217
rect 196 216 197 217
rect 195 216 196 217
rect 194 216 195 217
rect 180 216 181 217
rect 179 216 180 217
rect 175 216 176 217
rect 174 216 175 217
rect 173 216 174 217
rect 172 216 173 217
rect 166 216 167 217
rect 165 216 166 217
rect 151 216 152 217
rect 150 216 151 217
rect 149 216 150 217
rect 148 216 149 217
rect 147 216 148 217
rect 146 216 147 217
rect 145 216 146 217
rect 144 216 145 217
rect 143 216 144 217
rect 142 216 143 217
rect 132 216 133 217
rect 131 216 132 217
rect 130 216 131 217
rect 129 216 130 217
rect 128 216 129 217
rect 127 216 128 217
rect 126 216 127 217
rect 125 216 126 217
rect 124 216 125 217
rect 123 216 124 217
rect 114 216 115 217
rect 113 216 114 217
rect 112 216 113 217
rect 111 216 112 217
rect 110 216 111 217
rect 109 216 110 217
rect 108 216 109 217
rect 107 216 108 217
rect 106 216 107 217
rect 105 216 106 217
rect 104 216 105 217
rect 66 216 67 217
rect 65 216 66 217
rect 64 216 65 217
rect 63 216 64 217
rect 62 216 63 217
rect 61 216 62 217
rect 31 216 32 217
rect 30 216 31 217
rect 29 216 30 217
rect 25 216 26 217
rect 24 216 25 217
rect 23 216 24 217
rect 22 216 23 217
rect 21 216 22 217
rect 20 216 21 217
rect 19 216 20 217
rect 18 216 19 217
rect 17 216 18 217
rect 181 217 182 218
rect 180 217 181 218
rect 179 217 180 218
rect 178 217 179 218
rect 175 217 176 218
rect 174 217 175 218
rect 173 217 174 218
rect 172 217 173 218
rect 167 217 168 218
rect 166 217 167 218
rect 165 217 166 218
rect 164 217 165 218
rect 151 217 152 218
rect 150 217 151 218
rect 149 217 150 218
rect 148 217 149 218
rect 147 217 148 218
rect 146 217 147 218
rect 145 217 146 218
rect 144 217 145 218
rect 143 217 144 218
rect 142 217 143 218
rect 132 217 133 218
rect 131 217 132 218
rect 130 217 131 218
rect 129 217 130 218
rect 128 217 129 218
rect 127 217 128 218
rect 126 217 127 218
rect 125 217 126 218
rect 124 217 125 218
rect 123 217 124 218
rect 114 217 115 218
rect 113 217 114 218
rect 112 217 113 218
rect 111 217 112 218
rect 110 217 111 218
rect 109 217 110 218
rect 108 217 109 218
rect 107 217 108 218
rect 106 217 107 218
rect 105 217 106 218
rect 104 217 105 218
rect 65 217 66 218
rect 64 217 65 218
rect 63 217 64 218
rect 62 217 63 218
rect 61 217 62 218
rect 31 217 32 218
rect 30 217 31 218
rect 29 217 30 218
rect 24 217 25 218
rect 23 217 24 218
rect 22 217 23 218
rect 21 217 22 218
rect 20 217 21 218
rect 19 217 20 218
rect 18 217 19 218
rect 17 217 18 218
rect 198 218 199 219
rect 197 218 198 219
rect 196 218 197 219
rect 195 218 196 219
rect 194 218 195 219
rect 193 218 194 219
rect 181 218 182 219
rect 180 218 181 219
rect 179 218 180 219
rect 178 218 179 219
rect 175 218 176 219
rect 174 218 175 219
rect 173 218 174 219
rect 172 218 173 219
rect 167 218 168 219
rect 166 218 167 219
rect 165 218 166 219
rect 164 218 165 219
rect 151 218 152 219
rect 150 218 151 219
rect 149 218 150 219
rect 148 218 149 219
rect 147 218 148 219
rect 146 218 147 219
rect 145 218 146 219
rect 144 218 145 219
rect 143 218 144 219
rect 142 218 143 219
rect 132 218 133 219
rect 131 218 132 219
rect 130 218 131 219
rect 129 218 130 219
rect 128 218 129 219
rect 127 218 128 219
rect 126 218 127 219
rect 125 218 126 219
rect 124 218 125 219
rect 123 218 124 219
rect 114 218 115 219
rect 113 218 114 219
rect 112 218 113 219
rect 111 218 112 219
rect 110 218 111 219
rect 109 218 110 219
rect 108 218 109 219
rect 107 218 108 219
rect 106 218 107 219
rect 105 218 106 219
rect 104 218 105 219
rect 65 218 66 219
rect 64 218 65 219
rect 63 218 64 219
rect 62 218 63 219
rect 61 218 62 219
rect 60 218 61 219
rect 23 218 24 219
rect 22 218 23 219
rect 21 218 22 219
rect 20 218 21 219
rect 19 218 20 219
rect 18 218 19 219
rect 199 219 200 220
rect 198 219 199 220
rect 197 219 198 220
rect 196 219 197 220
rect 195 219 196 220
rect 194 219 195 220
rect 193 219 194 220
rect 181 219 182 220
rect 180 219 181 220
rect 179 219 180 220
rect 178 219 179 220
rect 175 219 176 220
rect 174 219 175 220
rect 173 219 174 220
rect 172 219 173 220
rect 167 219 168 220
rect 166 219 167 220
rect 165 219 166 220
rect 164 219 165 220
rect 151 219 152 220
rect 150 219 151 220
rect 149 219 150 220
rect 148 219 149 220
rect 147 219 148 220
rect 146 219 147 220
rect 145 219 146 220
rect 144 219 145 220
rect 143 219 144 220
rect 142 219 143 220
rect 132 219 133 220
rect 131 219 132 220
rect 130 219 131 220
rect 129 219 130 220
rect 128 219 129 220
rect 127 219 128 220
rect 126 219 127 220
rect 125 219 126 220
rect 124 219 125 220
rect 123 219 124 220
rect 114 219 115 220
rect 113 219 114 220
rect 112 219 113 220
rect 111 219 112 220
rect 110 219 111 220
rect 109 219 110 220
rect 108 219 109 220
rect 107 219 108 220
rect 106 219 107 220
rect 105 219 106 220
rect 104 219 105 220
rect 65 219 66 220
rect 64 219 65 220
rect 63 219 64 220
rect 62 219 63 220
rect 61 219 62 220
rect 60 219 61 220
rect 21 219 22 220
rect 20 219 21 220
rect 194 220 195 221
rect 193 220 194 221
rect 181 220 182 221
rect 180 220 181 221
rect 179 220 180 221
rect 178 220 179 221
rect 175 220 176 221
rect 174 220 175 221
rect 173 220 174 221
rect 172 220 173 221
rect 167 220 168 221
rect 166 220 167 221
rect 165 220 166 221
rect 164 220 165 221
rect 151 220 152 221
rect 150 220 151 221
rect 149 220 150 221
rect 148 220 149 221
rect 147 220 148 221
rect 146 220 147 221
rect 145 220 146 221
rect 144 220 145 221
rect 143 220 144 221
rect 142 220 143 221
rect 132 220 133 221
rect 131 220 132 221
rect 130 220 131 221
rect 129 220 130 221
rect 128 220 129 221
rect 127 220 128 221
rect 126 220 127 221
rect 125 220 126 221
rect 124 220 125 221
rect 123 220 124 221
rect 114 220 115 221
rect 113 220 114 221
rect 112 220 113 221
rect 111 220 112 221
rect 110 220 111 221
rect 109 220 110 221
rect 108 220 109 221
rect 107 220 108 221
rect 106 220 107 221
rect 105 220 106 221
rect 104 220 105 221
rect 65 220 66 221
rect 64 220 65 221
rect 63 220 64 221
rect 62 220 63 221
rect 61 220 62 221
rect 28 220 29 221
rect 27 220 28 221
rect 26 220 27 221
rect 194 221 195 222
rect 193 221 194 222
rect 181 221 182 222
rect 180 221 181 222
rect 179 221 180 222
rect 178 221 179 222
rect 175 221 176 222
rect 174 221 175 222
rect 173 221 174 222
rect 172 221 173 222
rect 167 221 168 222
rect 166 221 167 222
rect 165 221 166 222
rect 164 221 165 222
rect 151 221 152 222
rect 150 221 151 222
rect 149 221 150 222
rect 148 221 149 222
rect 147 221 148 222
rect 146 221 147 222
rect 145 221 146 222
rect 144 221 145 222
rect 143 221 144 222
rect 142 221 143 222
rect 132 221 133 222
rect 131 221 132 222
rect 130 221 131 222
rect 129 221 130 222
rect 128 221 129 222
rect 127 221 128 222
rect 126 221 127 222
rect 125 221 126 222
rect 124 221 125 222
rect 123 221 124 222
rect 114 221 115 222
rect 113 221 114 222
rect 112 221 113 222
rect 111 221 112 222
rect 110 221 111 222
rect 109 221 110 222
rect 108 221 109 222
rect 107 221 108 222
rect 106 221 107 222
rect 105 221 106 222
rect 104 221 105 222
rect 87 221 88 222
rect 86 221 87 222
rect 85 221 86 222
rect 65 221 66 222
rect 64 221 65 222
rect 63 221 64 222
rect 62 221 63 222
rect 61 221 62 222
rect 28 221 29 222
rect 27 221 28 222
rect 26 221 27 222
rect 25 221 26 222
rect 198 222 199 223
rect 197 222 198 223
rect 196 222 197 223
rect 195 222 196 223
rect 194 222 195 223
rect 193 222 194 223
rect 181 222 182 223
rect 180 222 181 223
rect 179 222 180 223
rect 178 222 179 223
rect 175 222 176 223
rect 174 222 175 223
rect 173 222 174 223
rect 172 222 173 223
rect 167 222 168 223
rect 166 222 167 223
rect 165 222 166 223
rect 164 222 165 223
rect 151 222 152 223
rect 150 222 151 223
rect 149 222 150 223
rect 148 222 149 223
rect 147 222 148 223
rect 146 222 147 223
rect 145 222 146 223
rect 144 222 145 223
rect 143 222 144 223
rect 142 222 143 223
rect 132 222 133 223
rect 131 222 132 223
rect 130 222 131 223
rect 129 222 130 223
rect 128 222 129 223
rect 127 222 128 223
rect 126 222 127 223
rect 125 222 126 223
rect 124 222 125 223
rect 123 222 124 223
rect 114 222 115 223
rect 113 222 114 223
rect 112 222 113 223
rect 111 222 112 223
rect 110 222 111 223
rect 109 222 110 223
rect 108 222 109 223
rect 107 222 108 223
rect 106 222 107 223
rect 105 222 106 223
rect 104 222 105 223
rect 88 222 89 223
rect 87 222 88 223
rect 86 222 87 223
rect 85 222 86 223
rect 62 222 63 223
rect 61 222 62 223
rect 28 222 29 223
rect 27 222 28 223
rect 26 222 27 223
rect 25 222 26 223
rect 24 222 25 223
rect 199 223 200 224
rect 198 223 199 224
rect 197 223 198 224
rect 196 223 197 224
rect 195 223 196 224
rect 194 223 195 224
rect 193 223 194 224
rect 181 223 182 224
rect 180 223 181 224
rect 179 223 180 224
rect 178 223 179 224
rect 175 223 176 224
rect 174 223 175 224
rect 173 223 174 224
rect 172 223 173 224
rect 167 223 168 224
rect 166 223 167 224
rect 165 223 166 224
rect 164 223 165 224
rect 151 223 152 224
rect 150 223 151 224
rect 149 223 150 224
rect 148 223 149 224
rect 147 223 148 224
rect 146 223 147 224
rect 145 223 146 224
rect 144 223 145 224
rect 143 223 144 224
rect 142 223 143 224
rect 132 223 133 224
rect 131 223 132 224
rect 130 223 131 224
rect 129 223 130 224
rect 128 223 129 224
rect 127 223 128 224
rect 126 223 127 224
rect 125 223 126 224
rect 124 223 125 224
rect 123 223 124 224
rect 114 223 115 224
rect 113 223 114 224
rect 112 223 113 224
rect 111 223 112 224
rect 110 223 111 224
rect 109 223 110 224
rect 108 223 109 224
rect 107 223 108 224
rect 106 223 107 224
rect 105 223 106 224
rect 104 223 105 224
rect 88 223 89 224
rect 87 223 88 224
rect 86 223 87 224
rect 85 223 86 224
rect 28 223 29 224
rect 27 223 28 224
rect 26 223 27 224
rect 25 223 26 224
rect 24 223 25 224
rect 23 223 24 224
rect 181 224 182 225
rect 180 224 181 225
rect 179 224 180 225
rect 178 224 179 225
rect 177 224 178 225
rect 176 224 177 225
rect 175 224 176 225
rect 174 224 175 225
rect 173 224 174 225
rect 172 224 173 225
rect 167 224 168 225
rect 166 224 167 225
rect 165 224 166 225
rect 164 224 165 225
rect 151 224 152 225
rect 150 224 151 225
rect 149 224 150 225
rect 148 224 149 225
rect 147 224 148 225
rect 146 224 147 225
rect 145 224 146 225
rect 144 224 145 225
rect 143 224 144 225
rect 142 224 143 225
rect 132 224 133 225
rect 131 224 132 225
rect 130 224 131 225
rect 129 224 130 225
rect 128 224 129 225
rect 127 224 128 225
rect 126 224 127 225
rect 125 224 126 225
rect 124 224 125 225
rect 123 224 124 225
rect 114 224 115 225
rect 113 224 114 225
rect 112 224 113 225
rect 111 224 112 225
rect 110 224 111 225
rect 109 224 110 225
rect 108 224 109 225
rect 107 224 108 225
rect 106 224 107 225
rect 105 224 106 225
rect 104 224 105 225
rect 88 224 89 225
rect 87 224 88 225
rect 86 224 87 225
rect 85 224 86 225
rect 28 224 29 225
rect 27 224 28 225
rect 26 224 27 225
rect 24 224 25 225
rect 23 224 24 225
rect 22 224 23 225
rect 198 225 199 226
rect 197 225 198 226
rect 196 225 197 226
rect 195 225 196 226
rect 194 225 195 226
rect 193 225 194 226
rect 191 225 192 226
rect 190 225 191 226
rect 181 225 182 226
rect 180 225 181 226
rect 179 225 180 226
rect 178 225 179 226
rect 177 225 178 226
rect 176 225 177 226
rect 175 225 176 226
rect 174 225 175 226
rect 173 225 174 226
rect 172 225 173 226
rect 167 225 168 226
rect 166 225 167 226
rect 165 225 166 226
rect 164 225 165 226
rect 151 225 152 226
rect 150 225 151 226
rect 149 225 150 226
rect 148 225 149 226
rect 147 225 148 226
rect 146 225 147 226
rect 145 225 146 226
rect 144 225 145 226
rect 143 225 144 226
rect 142 225 143 226
rect 132 225 133 226
rect 131 225 132 226
rect 130 225 131 226
rect 129 225 130 226
rect 128 225 129 226
rect 127 225 128 226
rect 126 225 127 226
rect 125 225 126 226
rect 124 225 125 226
rect 123 225 124 226
rect 114 225 115 226
rect 113 225 114 226
rect 112 225 113 226
rect 111 225 112 226
rect 110 225 111 226
rect 109 225 110 226
rect 108 225 109 226
rect 107 225 108 226
rect 106 225 107 226
rect 105 225 106 226
rect 104 225 105 226
rect 88 225 89 226
rect 87 225 88 226
rect 86 225 87 226
rect 85 225 86 226
rect 31 225 32 226
rect 30 225 31 226
rect 28 225 29 226
rect 27 225 28 226
rect 26 225 27 226
rect 23 225 24 226
rect 22 225 23 226
rect 21 225 22 226
rect 20 225 21 226
rect 198 226 199 227
rect 197 226 198 227
rect 196 226 197 227
rect 195 226 196 227
rect 194 226 195 227
rect 193 226 194 227
rect 191 226 192 227
rect 190 226 191 227
rect 181 226 182 227
rect 180 226 181 227
rect 179 226 180 227
rect 178 226 179 227
rect 177 226 178 227
rect 176 226 177 227
rect 175 226 176 227
rect 174 226 175 227
rect 173 226 174 227
rect 172 226 173 227
rect 167 226 168 227
rect 166 226 167 227
rect 165 226 166 227
rect 164 226 165 227
rect 151 226 152 227
rect 150 226 151 227
rect 149 226 150 227
rect 148 226 149 227
rect 147 226 148 227
rect 146 226 147 227
rect 145 226 146 227
rect 144 226 145 227
rect 143 226 144 227
rect 142 226 143 227
rect 132 226 133 227
rect 131 226 132 227
rect 130 226 131 227
rect 129 226 130 227
rect 128 226 129 227
rect 127 226 128 227
rect 126 226 127 227
rect 125 226 126 227
rect 124 226 125 227
rect 123 226 124 227
rect 114 226 115 227
rect 113 226 114 227
rect 112 226 113 227
rect 111 226 112 227
rect 110 226 111 227
rect 109 226 110 227
rect 108 226 109 227
rect 107 226 108 227
rect 106 226 107 227
rect 105 226 106 227
rect 104 226 105 227
rect 88 226 89 227
rect 87 226 88 227
rect 86 226 87 227
rect 85 226 86 227
rect 31 226 32 227
rect 30 226 31 227
rect 29 226 30 227
rect 28 226 29 227
rect 27 226 28 227
rect 26 226 27 227
rect 25 226 26 227
rect 22 226 23 227
rect 21 226 22 227
rect 20 226 21 227
rect 19 226 20 227
rect 181 227 182 228
rect 180 227 181 228
rect 179 227 180 228
rect 178 227 179 228
rect 175 227 176 228
rect 174 227 175 228
rect 173 227 174 228
rect 172 227 173 228
rect 167 227 168 228
rect 166 227 167 228
rect 165 227 166 228
rect 164 227 165 228
rect 151 227 152 228
rect 150 227 151 228
rect 149 227 150 228
rect 148 227 149 228
rect 147 227 148 228
rect 146 227 147 228
rect 145 227 146 228
rect 144 227 145 228
rect 143 227 144 228
rect 142 227 143 228
rect 132 227 133 228
rect 131 227 132 228
rect 130 227 131 228
rect 129 227 130 228
rect 128 227 129 228
rect 127 227 128 228
rect 126 227 127 228
rect 125 227 126 228
rect 124 227 125 228
rect 123 227 124 228
rect 114 227 115 228
rect 113 227 114 228
rect 112 227 113 228
rect 111 227 112 228
rect 110 227 111 228
rect 109 227 110 228
rect 108 227 109 228
rect 107 227 108 228
rect 106 227 107 228
rect 105 227 106 228
rect 104 227 105 228
rect 88 227 89 228
rect 87 227 88 228
rect 86 227 87 228
rect 85 227 86 228
rect 31 227 32 228
rect 30 227 31 228
rect 29 227 30 228
rect 28 227 29 228
rect 27 227 28 228
rect 26 227 27 228
rect 25 227 26 228
rect 24 227 25 228
rect 23 227 24 228
rect 22 227 23 228
rect 21 227 22 228
rect 20 227 21 228
rect 19 227 20 228
rect 18 227 19 228
rect 197 228 198 229
rect 196 228 197 229
rect 195 228 196 229
rect 194 228 195 229
rect 181 228 182 229
rect 180 228 181 229
rect 179 228 180 229
rect 178 228 179 229
rect 175 228 176 229
rect 174 228 175 229
rect 173 228 174 229
rect 172 228 173 229
rect 167 228 168 229
rect 166 228 167 229
rect 165 228 166 229
rect 164 228 165 229
rect 151 228 152 229
rect 150 228 151 229
rect 149 228 150 229
rect 148 228 149 229
rect 147 228 148 229
rect 146 228 147 229
rect 145 228 146 229
rect 144 228 145 229
rect 143 228 144 229
rect 142 228 143 229
rect 132 228 133 229
rect 131 228 132 229
rect 130 228 131 229
rect 129 228 130 229
rect 128 228 129 229
rect 127 228 128 229
rect 126 228 127 229
rect 125 228 126 229
rect 124 228 125 229
rect 123 228 124 229
rect 114 228 115 229
rect 113 228 114 229
rect 112 228 113 229
rect 111 228 112 229
rect 110 228 111 229
rect 109 228 110 229
rect 108 228 109 229
rect 107 228 108 229
rect 106 228 107 229
rect 105 228 106 229
rect 104 228 105 229
rect 88 228 89 229
rect 87 228 88 229
rect 86 228 87 229
rect 85 228 86 229
rect 29 228 30 229
rect 28 228 29 229
rect 27 228 28 229
rect 26 228 27 229
rect 25 228 26 229
rect 24 228 25 229
rect 23 228 24 229
rect 22 228 23 229
rect 21 228 22 229
rect 20 228 21 229
rect 19 228 20 229
rect 18 228 19 229
rect 17 228 18 229
rect 198 229 199 230
rect 197 229 198 230
rect 196 229 197 230
rect 195 229 196 230
rect 194 229 195 230
rect 193 229 194 230
rect 181 229 182 230
rect 180 229 181 230
rect 179 229 180 230
rect 178 229 179 230
rect 175 229 176 230
rect 174 229 175 230
rect 173 229 174 230
rect 172 229 173 230
rect 167 229 168 230
rect 166 229 167 230
rect 165 229 166 230
rect 164 229 165 230
rect 151 229 152 230
rect 150 229 151 230
rect 149 229 150 230
rect 148 229 149 230
rect 147 229 148 230
rect 146 229 147 230
rect 145 229 146 230
rect 144 229 145 230
rect 143 229 144 230
rect 142 229 143 230
rect 132 229 133 230
rect 131 229 132 230
rect 130 229 131 230
rect 129 229 130 230
rect 128 229 129 230
rect 127 229 128 230
rect 126 229 127 230
rect 125 229 126 230
rect 124 229 125 230
rect 123 229 124 230
rect 114 229 115 230
rect 113 229 114 230
rect 112 229 113 230
rect 111 229 112 230
rect 110 229 111 230
rect 109 229 110 230
rect 108 229 109 230
rect 107 229 108 230
rect 106 229 107 230
rect 105 229 106 230
rect 104 229 105 230
rect 88 229 89 230
rect 87 229 88 230
rect 86 229 87 230
rect 85 229 86 230
rect 28 229 29 230
rect 27 229 28 230
rect 26 229 27 230
rect 24 229 25 230
rect 23 229 24 230
rect 22 229 23 230
rect 21 229 22 230
rect 20 229 21 230
rect 19 229 20 230
rect 18 229 19 230
rect 17 229 18 230
rect 198 230 199 231
rect 197 230 198 231
rect 194 230 195 231
rect 193 230 194 231
rect 181 230 182 231
rect 180 230 181 231
rect 179 230 180 231
rect 178 230 179 231
rect 175 230 176 231
rect 174 230 175 231
rect 173 230 174 231
rect 172 230 173 231
rect 167 230 168 231
rect 166 230 167 231
rect 165 230 166 231
rect 164 230 165 231
rect 151 230 152 231
rect 150 230 151 231
rect 149 230 150 231
rect 148 230 149 231
rect 147 230 148 231
rect 146 230 147 231
rect 145 230 146 231
rect 144 230 145 231
rect 143 230 144 231
rect 142 230 143 231
rect 132 230 133 231
rect 131 230 132 231
rect 130 230 131 231
rect 129 230 130 231
rect 128 230 129 231
rect 127 230 128 231
rect 126 230 127 231
rect 125 230 126 231
rect 124 230 125 231
rect 123 230 124 231
rect 114 230 115 231
rect 113 230 114 231
rect 112 230 113 231
rect 111 230 112 231
rect 110 230 111 231
rect 109 230 110 231
rect 108 230 109 231
rect 107 230 108 231
rect 106 230 107 231
rect 105 230 106 231
rect 104 230 105 231
rect 88 230 89 231
rect 87 230 88 231
rect 86 230 87 231
rect 85 230 86 231
rect 27 230 28 231
rect 26 230 27 231
rect 20 230 21 231
rect 19 230 20 231
rect 18 230 19 231
rect 17 230 18 231
rect 199 231 200 232
rect 198 231 199 232
rect 194 231 195 232
rect 193 231 194 232
rect 185 231 186 232
rect 184 231 185 232
rect 183 231 184 232
rect 182 231 183 232
rect 181 231 182 232
rect 180 231 181 232
rect 179 231 180 232
rect 178 231 179 232
rect 175 231 176 232
rect 174 231 175 232
rect 173 231 174 232
rect 172 231 173 232
rect 171 231 172 232
rect 170 231 171 232
rect 169 231 170 232
rect 168 231 169 232
rect 167 231 168 232
rect 166 231 167 232
rect 165 231 166 232
rect 164 231 165 232
rect 151 231 152 232
rect 150 231 151 232
rect 149 231 150 232
rect 148 231 149 232
rect 147 231 148 232
rect 146 231 147 232
rect 145 231 146 232
rect 144 231 145 232
rect 143 231 144 232
rect 142 231 143 232
rect 132 231 133 232
rect 131 231 132 232
rect 130 231 131 232
rect 129 231 130 232
rect 128 231 129 232
rect 127 231 128 232
rect 126 231 127 232
rect 125 231 126 232
rect 124 231 125 232
rect 123 231 124 232
rect 114 231 115 232
rect 113 231 114 232
rect 112 231 113 232
rect 111 231 112 232
rect 110 231 111 232
rect 109 231 110 232
rect 108 231 109 232
rect 107 231 108 232
rect 106 231 107 232
rect 105 231 106 232
rect 104 231 105 232
rect 88 231 89 232
rect 87 231 88 232
rect 86 231 87 232
rect 85 231 86 232
rect 198 232 199 233
rect 193 232 194 233
rect 185 232 186 233
rect 184 232 185 233
rect 183 232 184 233
rect 182 232 183 233
rect 181 232 182 233
rect 180 232 181 233
rect 179 232 180 233
rect 178 232 179 233
rect 175 232 176 233
rect 174 232 175 233
rect 173 232 174 233
rect 172 232 173 233
rect 171 232 172 233
rect 170 232 171 233
rect 169 232 170 233
rect 168 232 169 233
rect 167 232 168 233
rect 166 232 167 233
rect 165 232 166 233
rect 164 232 165 233
rect 151 232 152 233
rect 150 232 151 233
rect 149 232 150 233
rect 148 232 149 233
rect 147 232 148 233
rect 146 232 147 233
rect 145 232 146 233
rect 144 232 145 233
rect 143 232 144 233
rect 142 232 143 233
rect 132 232 133 233
rect 131 232 132 233
rect 130 232 131 233
rect 129 232 130 233
rect 128 232 129 233
rect 127 232 128 233
rect 126 232 127 233
rect 125 232 126 233
rect 124 232 125 233
rect 123 232 124 233
rect 114 232 115 233
rect 113 232 114 233
rect 112 232 113 233
rect 111 232 112 233
rect 110 232 111 233
rect 109 232 110 233
rect 108 232 109 233
rect 107 232 108 233
rect 106 232 107 233
rect 105 232 106 233
rect 104 232 105 233
rect 88 232 89 233
rect 87 232 88 233
rect 86 232 87 233
rect 85 232 86 233
rect 27 232 28 233
rect 26 232 27 233
rect 25 232 26 233
rect 198 233 199 234
rect 195 233 196 234
rect 194 233 195 234
rect 185 233 186 234
rect 184 233 185 234
rect 183 233 184 234
rect 182 233 183 234
rect 181 233 182 234
rect 180 233 181 234
rect 179 233 180 234
rect 178 233 179 234
rect 175 233 176 234
rect 174 233 175 234
rect 173 233 174 234
rect 172 233 173 234
rect 171 233 172 234
rect 170 233 171 234
rect 169 233 170 234
rect 168 233 169 234
rect 167 233 168 234
rect 166 233 167 234
rect 165 233 166 234
rect 164 233 165 234
rect 151 233 152 234
rect 150 233 151 234
rect 149 233 150 234
rect 148 233 149 234
rect 147 233 148 234
rect 146 233 147 234
rect 145 233 146 234
rect 144 233 145 234
rect 143 233 144 234
rect 142 233 143 234
rect 132 233 133 234
rect 131 233 132 234
rect 130 233 131 234
rect 129 233 130 234
rect 128 233 129 234
rect 127 233 128 234
rect 126 233 127 234
rect 125 233 126 234
rect 124 233 125 234
rect 123 233 124 234
rect 114 233 115 234
rect 113 233 114 234
rect 112 233 113 234
rect 111 233 112 234
rect 110 233 111 234
rect 109 233 110 234
rect 108 233 109 234
rect 107 233 108 234
rect 106 233 107 234
rect 105 233 106 234
rect 104 233 105 234
rect 88 233 89 234
rect 87 233 88 234
rect 86 233 87 234
rect 85 233 86 234
rect 27 233 28 234
rect 26 233 27 234
rect 25 233 26 234
rect 199 234 200 235
rect 198 234 199 235
rect 196 234 197 235
rect 195 234 196 235
rect 194 234 195 235
rect 193 234 194 235
rect 185 234 186 235
rect 184 234 185 235
rect 183 234 184 235
rect 182 234 183 235
rect 181 234 182 235
rect 180 234 181 235
rect 179 234 180 235
rect 178 234 179 235
rect 175 234 176 235
rect 174 234 175 235
rect 173 234 174 235
rect 172 234 173 235
rect 171 234 172 235
rect 170 234 171 235
rect 169 234 170 235
rect 168 234 169 235
rect 167 234 168 235
rect 166 234 167 235
rect 165 234 166 235
rect 164 234 165 235
rect 151 234 152 235
rect 150 234 151 235
rect 149 234 150 235
rect 148 234 149 235
rect 147 234 148 235
rect 146 234 147 235
rect 145 234 146 235
rect 144 234 145 235
rect 143 234 144 235
rect 142 234 143 235
rect 132 234 133 235
rect 131 234 132 235
rect 130 234 131 235
rect 129 234 130 235
rect 128 234 129 235
rect 127 234 128 235
rect 126 234 127 235
rect 125 234 126 235
rect 124 234 125 235
rect 123 234 124 235
rect 114 234 115 235
rect 113 234 114 235
rect 112 234 113 235
rect 111 234 112 235
rect 110 234 111 235
rect 109 234 110 235
rect 108 234 109 235
rect 107 234 108 235
rect 106 234 107 235
rect 105 234 106 235
rect 104 234 105 235
rect 88 234 89 235
rect 87 234 88 235
rect 86 234 87 235
rect 85 234 86 235
rect 27 234 28 235
rect 26 234 27 235
rect 25 234 26 235
rect 199 235 200 236
rect 198 235 199 236
rect 196 235 197 236
rect 195 235 196 236
rect 194 235 195 236
rect 193 235 194 236
rect 175 235 176 236
rect 174 235 175 236
rect 173 235 174 236
rect 172 235 173 236
rect 166 235 167 236
rect 165 235 166 236
rect 151 235 152 236
rect 150 235 151 236
rect 149 235 150 236
rect 148 235 149 236
rect 147 235 148 236
rect 146 235 147 236
rect 145 235 146 236
rect 144 235 145 236
rect 143 235 144 236
rect 142 235 143 236
rect 132 235 133 236
rect 131 235 132 236
rect 130 235 131 236
rect 129 235 130 236
rect 128 235 129 236
rect 127 235 128 236
rect 126 235 127 236
rect 125 235 126 236
rect 124 235 125 236
rect 123 235 124 236
rect 114 235 115 236
rect 113 235 114 236
rect 112 235 113 236
rect 111 235 112 236
rect 110 235 111 236
rect 109 235 110 236
rect 108 235 109 236
rect 107 235 108 236
rect 106 235 107 236
rect 105 235 106 236
rect 104 235 105 236
rect 88 235 89 236
rect 87 235 88 236
rect 86 235 87 236
rect 85 235 86 236
rect 27 235 28 236
rect 26 235 27 236
rect 25 235 26 236
rect 199 236 200 237
rect 198 236 199 237
rect 197 236 198 237
rect 196 236 197 237
rect 194 236 195 237
rect 193 236 194 237
rect 175 236 176 237
rect 174 236 175 237
rect 173 236 174 237
rect 172 236 173 237
rect 151 236 152 237
rect 150 236 151 237
rect 149 236 150 237
rect 148 236 149 237
rect 147 236 148 237
rect 146 236 147 237
rect 145 236 146 237
rect 144 236 145 237
rect 143 236 144 237
rect 142 236 143 237
rect 132 236 133 237
rect 131 236 132 237
rect 130 236 131 237
rect 129 236 130 237
rect 128 236 129 237
rect 127 236 128 237
rect 126 236 127 237
rect 125 236 126 237
rect 124 236 125 237
rect 123 236 124 237
rect 114 236 115 237
rect 113 236 114 237
rect 112 236 113 237
rect 111 236 112 237
rect 110 236 111 237
rect 109 236 110 237
rect 108 236 109 237
rect 107 236 108 237
rect 106 236 107 237
rect 105 236 106 237
rect 104 236 105 237
rect 88 236 89 237
rect 87 236 88 237
rect 86 236 87 237
rect 85 236 86 237
rect 27 236 28 237
rect 26 236 27 237
rect 25 236 26 237
rect 198 237 199 238
rect 197 237 198 238
rect 196 237 197 238
rect 194 237 195 238
rect 193 237 194 238
rect 175 237 176 238
rect 174 237 175 238
rect 173 237 174 238
rect 172 237 173 238
rect 151 237 152 238
rect 150 237 151 238
rect 149 237 150 238
rect 148 237 149 238
rect 147 237 148 238
rect 146 237 147 238
rect 145 237 146 238
rect 144 237 145 238
rect 143 237 144 238
rect 142 237 143 238
rect 132 237 133 238
rect 131 237 132 238
rect 130 237 131 238
rect 129 237 130 238
rect 128 237 129 238
rect 127 237 128 238
rect 126 237 127 238
rect 125 237 126 238
rect 124 237 125 238
rect 123 237 124 238
rect 114 237 115 238
rect 113 237 114 238
rect 112 237 113 238
rect 111 237 112 238
rect 110 237 111 238
rect 109 237 110 238
rect 108 237 109 238
rect 107 237 108 238
rect 106 237 107 238
rect 105 237 106 238
rect 104 237 105 238
rect 88 237 89 238
rect 87 237 88 238
rect 86 237 87 238
rect 85 237 86 238
rect 27 237 28 238
rect 26 237 27 238
rect 25 237 26 238
rect 174 238 175 239
rect 173 238 174 239
rect 151 238 152 239
rect 150 238 151 239
rect 149 238 150 239
rect 148 238 149 239
rect 147 238 148 239
rect 146 238 147 239
rect 145 238 146 239
rect 144 238 145 239
rect 143 238 144 239
rect 142 238 143 239
rect 132 238 133 239
rect 131 238 132 239
rect 130 238 131 239
rect 129 238 130 239
rect 128 238 129 239
rect 127 238 128 239
rect 126 238 127 239
rect 125 238 126 239
rect 124 238 125 239
rect 123 238 124 239
rect 114 238 115 239
rect 113 238 114 239
rect 112 238 113 239
rect 111 238 112 239
rect 110 238 111 239
rect 109 238 110 239
rect 108 238 109 239
rect 107 238 108 239
rect 106 238 107 239
rect 105 238 106 239
rect 104 238 105 239
rect 88 238 89 239
rect 87 238 88 239
rect 86 238 87 239
rect 85 238 86 239
rect 151 239 152 240
rect 150 239 151 240
rect 149 239 150 240
rect 148 239 149 240
rect 147 239 148 240
rect 146 239 147 240
rect 145 239 146 240
rect 144 239 145 240
rect 143 239 144 240
rect 142 239 143 240
rect 132 239 133 240
rect 131 239 132 240
rect 130 239 131 240
rect 129 239 130 240
rect 128 239 129 240
rect 127 239 128 240
rect 126 239 127 240
rect 125 239 126 240
rect 124 239 125 240
rect 123 239 124 240
rect 114 239 115 240
rect 113 239 114 240
rect 112 239 113 240
rect 111 239 112 240
rect 110 239 111 240
rect 109 239 110 240
rect 108 239 109 240
rect 107 239 108 240
rect 106 239 107 240
rect 105 239 106 240
rect 104 239 105 240
rect 88 239 89 240
rect 87 239 88 240
rect 86 239 87 240
rect 85 239 86 240
rect 28 239 29 240
rect 27 239 28 240
rect 151 240 152 241
rect 150 240 151 241
rect 149 240 150 241
rect 148 240 149 241
rect 147 240 148 241
rect 146 240 147 241
rect 145 240 146 241
rect 144 240 145 241
rect 143 240 144 241
rect 142 240 143 241
rect 132 240 133 241
rect 131 240 132 241
rect 130 240 131 241
rect 129 240 130 241
rect 128 240 129 241
rect 127 240 128 241
rect 126 240 127 241
rect 125 240 126 241
rect 124 240 125 241
rect 123 240 124 241
rect 114 240 115 241
rect 113 240 114 241
rect 112 240 113 241
rect 111 240 112 241
rect 110 240 111 241
rect 109 240 110 241
rect 108 240 109 241
rect 107 240 108 241
rect 106 240 107 241
rect 105 240 106 241
rect 104 240 105 241
rect 88 240 89 241
rect 87 240 88 241
rect 86 240 87 241
rect 85 240 86 241
rect 30 240 31 241
rect 29 240 30 241
rect 28 240 29 241
rect 27 240 28 241
rect 151 241 152 242
rect 150 241 151 242
rect 149 241 150 242
rect 148 241 149 242
rect 147 241 148 242
rect 146 241 147 242
rect 145 241 146 242
rect 144 241 145 242
rect 143 241 144 242
rect 142 241 143 242
rect 132 241 133 242
rect 131 241 132 242
rect 130 241 131 242
rect 129 241 130 242
rect 128 241 129 242
rect 127 241 128 242
rect 126 241 127 242
rect 125 241 126 242
rect 124 241 125 242
rect 123 241 124 242
rect 114 241 115 242
rect 113 241 114 242
rect 112 241 113 242
rect 111 241 112 242
rect 110 241 111 242
rect 109 241 110 242
rect 108 241 109 242
rect 107 241 108 242
rect 106 241 107 242
rect 105 241 106 242
rect 104 241 105 242
rect 88 241 89 242
rect 87 241 88 242
rect 86 241 87 242
rect 85 241 86 242
rect 30 241 31 242
rect 29 241 30 242
rect 28 241 29 242
rect 27 241 28 242
rect 21 241 22 242
rect 20 241 21 242
rect 19 241 20 242
rect 198 242 199 243
rect 197 242 198 243
rect 196 242 197 243
rect 194 242 195 243
rect 193 242 194 243
rect 151 242 152 243
rect 150 242 151 243
rect 149 242 150 243
rect 148 242 149 243
rect 147 242 148 243
rect 146 242 147 243
rect 145 242 146 243
rect 144 242 145 243
rect 143 242 144 243
rect 142 242 143 243
rect 132 242 133 243
rect 131 242 132 243
rect 130 242 131 243
rect 129 242 130 243
rect 128 242 129 243
rect 127 242 128 243
rect 126 242 127 243
rect 125 242 126 243
rect 124 242 125 243
rect 123 242 124 243
rect 114 242 115 243
rect 113 242 114 243
rect 112 242 113 243
rect 111 242 112 243
rect 110 242 111 243
rect 109 242 110 243
rect 108 242 109 243
rect 107 242 108 243
rect 106 242 107 243
rect 105 242 106 243
rect 104 242 105 243
rect 88 242 89 243
rect 87 242 88 243
rect 86 242 87 243
rect 85 242 86 243
rect 31 242 32 243
rect 30 242 31 243
rect 29 242 30 243
rect 28 242 29 243
rect 21 242 22 243
rect 20 242 21 243
rect 19 242 20 243
rect 18 242 19 243
rect 198 243 199 244
rect 197 243 198 244
rect 196 243 197 244
rect 195 243 196 244
rect 194 243 195 244
rect 193 243 194 244
rect 151 243 152 244
rect 150 243 151 244
rect 149 243 150 244
rect 148 243 149 244
rect 147 243 148 244
rect 146 243 147 244
rect 145 243 146 244
rect 144 243 145 244
rect 143 243 144 244
rect 142 243 143 244
rect 132 243 133 244
rect 131 243 132 244
rect 130 243 131 244
rect 129 243 130 244
rect 128 243 129 244
rect 127 243 128 244
rect 126 243 127 244
rect 125 243 126 244
rect 124 243 125 244
rect 123 243 124 244
rect 114 243 115 244
rect 113 243 114 244
rect 112 243 113 244
rect 111 243 112 244
rect 110 243 111 244
rect 109 243 110 244
rect 108 243 109 244
rect 107 243 108 244
rect 106 243 107 244
rect 105 243 106 244
rect 104 243 105 244
rect 87 243 88 244
rect 86 243 87 244
rect 85 243 86 244
rect 31 243 32 244
rect 30 243 31 244
rect 29 243 30 244
rect 21 243 22 244
rect 20 243 21 244
rect 19 243 20 244
rect 18 243 19 244
rect 17 243 18 244
rect 199 244 200 245
rect 198 244 199 245
rect 196 244 197 245
rect 195 244 196 245
rect 194 244 195 245
rect 193 244 194 245
rect 151 244 152 245
rect 150 244 151 245
rect 149 244 150 245
rect 148 244 149 245
rect 147 244 148 245
rect 146 244 147 245
rect 145 244 146 245
rect 144 244 145 245
rect 143 244 144 245
rect 142 244 143 245
rect 132 244 133 245
rect 131 244 132 245
rect 130 244 131 245
rect 129 244 130 245
rect 128 244 129 245
rect 127 244 128 245
rect 126 244 127 245
rect 125 244 126 245
rect 124 244 125 245
rect 123 244 124 245
rect 114 244 115 245
rect 113 244 114 245
rect 112 244 113 245
rect 111 244 112 245
rect 110 244 111 245
rect 109 244 110 245
rect 108 244 109 245
rect 107 244 108 245
rect 106 244 107 245
rect 105 244 106 245
rect 104 244 105 245
rect 31 244 32 245
rect 30 244 31 245
rect 29 244 30 245
rect 24 244 25 245
rect 23 244 24 245
rect 19 244 20 245
rect 18 244 19 245
rect 17 244 18 245
rect 198 245 199 246
rect 197 245 198 246
rect 196 245 197 246
rect 195 245 196 246
rect 194 245 195 246
rect 193 245 194 246
rect 151 245 152 246
rect 150 245 151 246
rect 149 245 150 246
rect 148 245 149 246
rect 147 245 148 246
rect 146 245 147 246
rect 145 245 146 246
rect 144 245 145 246
rect 143 245 144 246
rect 142 245 143 246
rect 132 245 133 246
rect 131 245 132 246
rect 130 245 131 246
rect 129 245 130 246
rect 128 245 129 246
rect 127 245 128 246
rect 126 245 127 246
rect 125 245 126 246
rect 124 245 125 246
rect 123 245 124 246
rect 114 245 115 246
rect 113 245 114 246
rect 112 245 113 246
rect 111 245 112 246
rect 110 245 111 246
rect 109 245 110 246
rect 108 245 109 246
rect 107 245 108 246
rect 106 245 107 246
rect 105 245 106 246
rect 104 245 105 246
rect 31 245 32 246
rect 30 245 31 246
rect 29 245 30 246
rect 25 245 26 246
rect 24 245 25 246
rect 23 245 24 246
rect 22 245 23 246
rect 19 245 20 246
rect 18 245 19 246
rect 17 245 18 246
rect 199 246 200 247
rect 198 246 199 247
rect 197 246 198 247
rect 196 246 197 247
rect 195 246 196 247
rect 194 246 195 247
rect 193 246 194 247
rect 151 246 152 247
rect 150 246 151 247
rect 149 246 150 247
rect 148 246 149 247
rect 147 246 148 247
rect 146 246 147 247
rect 145 246 146 247
rect 144 246 145 247
rect 143 246 144 247
rect 142 246 143 247
rect 132 246 133 247
rect 131 246 132 247
rect 130 246 131 247
rect 129 246 130 247
rect 128 246 129 247
rect 127 246 128 247
rect 126 246 127 247
rect 125 246 126 247
rect 124 246 125 247
rect 123 246 124 247
rect 114 246 115 247
rect 113 246 114 247
rect 112 246 113 247
rect 111 246 112 247
rect 110 246 111 247
rect 109 246 110 247
rect 108 246 109 247
rect 107 246 108 247
rect 106 246 107 247
rect 105 246 106 247
rect 104 246 105 247
rect 88 246 89 247
rect 87 246 88 247
rect 86 246 87 247
rect 85 246 86 247
rect 84 246 85 247
rect 83 246 84 247
rect 82 246 83 247
rect 81 246 82 247
rect 80 246 81 247
rect 79 246 80 247
rect 78 246 79 247
rect 77 246 78 247
rect 76 246 77 247
rect 75 246 76 247
rect 74 246 75 247
rect 73 246 74 247
rect 72 246 73 247
rect 71 246 72 247
rect 70 246 71 247
rect 69 246 70 247
rect 68 246 69 247
rect 67 246 68 247
rect 66 246 67 247
rect 65 246 66 247
rect 64 246 65 247
rect 63 246 64 247
rect 62 246 63 247
rect 61 246 62 247
rect 30 246 31 247
rect 29 246 30 247
rect 28 246 29 247
rect 27 246 28 247
rect 26 246 27 247
rect 25 246 26 247
rect 24 246 25 247
rect 23 246 24 247
rect 22 246 23 247
rect 19 246 20 247
rect 18 246 19 247
rect 17 246 18 247
rect 198 247 199 248
rect 197 247 198 248
rect 196 247 197 248
rect 195 247 196 248
rect 194 247 195 248
rect 151 247 152 248
rect 150 247 151 248
rect 149 247 150 248
rect 148 247 149 248
rect 147 247 148 248
rect 146 247 147 248
rect 145 247 146 248
rect 144 247 145 248
rect 143 247 144 248
rect 142 247 143 248
rect 132 247 133 248
rect 131 247 132 248
rect 130 247 131 248
rect 129 247 130 248
rect 128 247 129 248
rect 127 247 128 248
rect 126 247 127 248
rect 125 247 126 248
rect 124 247 125 248
rect 123 247 124 248
rect 114 247 115 248
rect 113 247 114 248
rect 112 247 113 248
rect 111 247 112 248
rect 110 247 111 248
rect 109 247 110 248
rect 108 247 109 248
rect 107 247 108 248
rect 106 247 107 248
rect 105 247 106 248
rect 104 247 105 248
rect 88 247 89 248
rect 87 247 88 248
rect 86 247 87 248
rect 85 247 86 248
rect 84 247 85 248
rect 83 247 84 248
rect 82 247 83 248
rect 81 247 82 248
rect 80 247 81 248
rect 79 247 80 248
rect 78 247 79 248
rect 77 247 78 248
rect 76 247 77 248
rect 75 247 76 248
rect 74 247 75 248
rect 73 247 74 248
rect 72 247 73 248
rect 71 247 72 248
rect 70 247 71 248
rect 69 247 70 248
rect 68 247 69 248
rect 67 247 68 248
rect 66 247 67 248
rect 65 247 66 248
rect 64 247 65 248
rect 63 247 64 248
rect 62 247 63 248
rect 61 247 62 248
rect 30 247 31 248
rect 29 247 30 248
rect 28 247 29 248
rect 27 247 28 248
rect 26 247 27 248
rect 25 247 26 248
rect 24 247 25 248
rect 23 247 24 248
rect 22 247 23 248
rect 21 247 22 248
rect 20 247 21 248
rect 19 247 20 248
rect 18 247 19 248
rect 17 247 18 248
rect 151 248 152 249
rect 150 248 151 249
rect 149 248 150 249
rect 148 248 149 249
rect 147 248 148 249
rect 146 248 147 249
rect 145 248 146 249
rect 144 248 145 249
rect 143 248 144 249
rect 142 248 143 249
rect 132 248 133 249
rect 131 248 132 249
rect 130 248 131 249
rect 129 248 130 249
rect 128 248 129 249
rect 127 248 128 249
rect 126 248 127 249
rect 125 248 126 249
rect 124 248 125 249
rect 123 248 124 249
rect 114 248 115 249
rect 113 248 114 249
rect 112 248 113 249
rect 111 248 112 249
rect 110 248 111 249
rect 109 248 110 249
rect 108 248 109 249
rect 107 248 108 249
rect 106 248 107 249
rect 105 248 106 249
rect 104 248 105 249
rect 88 248 89 249
rect 87 248 88 249
rect 86 248 87 249
rect 85 248 86 249
rect 84 248 85 249
rect 83 248 84 249
rect 82 248 83 249
rect 81 248 82 249
rect 80 248 81 249
rect 79 248 80 249
rect 78 248 79 249
rect 77 248 78 249
rect 76 248 77 249
rect 75 248 76 249
rect 74 248 75 249
rect 73 248 74 249
rect 72 248 73 249
rect 71 248 72 249
rect 70 248 71 249
rect 69 248 70 249
rect 68 248 69 249
rect 67 248 68 249
rect 66 248 67 249
rect 65 248 66 249
rect 64 248 65 249
rect 63 248 64 249
rect 62 248 63 249
rect 61 248 62 249
rect 29 248 30 249
rect 28 248 29 249
rect 27 248 28 249
rect 26 248 27 249
rect 25 248 26 249
rect 23 248 24 249
rect 22 248 23 249
rect 21 248 22 249
rect 20 248 21 249
rect 19 248 20 249
rect 18 248 19 249
rect 199 249 200 250
rect 198 249 199 250
rect 197 249 198 250
rect 196 249 197 250
rect 195 249 196 250
rect 194 249 195 250
rect 193 249 194 250
rect 175 249 176 250
rect 174 249 175 250
rect 151 249 152 250
rect 150 249 151 250
rect 149 249 150 250
rect 148 249 149 250
rect 147 249 148 250
rect 146 249 147 250
rect 145 249 146 250
rect 144 249 145 250
rect 143 249 144 250
rect 142 249 143 250
rect 132 249 133 250
rect 131 249 132 250
rect 130 249 131 250
rect 129 249 130 250
rect 128 249 129 250
rect 127 249 128 250
rect 126 249 127 250
rect 125 249 126 250
rect 124 249 125 250
rect 123 249 124 250
rect 114 249 115 250
rect 113 249 114 250
rect 112 249 113 250
rect 111 249 112 250
rect 110 249 111 250
rect 109 249 110 250
rect 108 249 109 250
rect 107 249 108 250
rect 106 249 107 250
rect 105 249 106 250
rect 104 249 105 250
rect 88 249 89 250
rect 87 249 88 250
rect 86 249 87 250
rect 85 249 86 250
rect 84 249 85 250
rect 83 249 84 250
rect 82 249 83 250
rect 81 249 82 250
rect 80 249 81 250
rect 79 249 80 250
rect 78 249 79 250
rect 77 249 78 250
rect 76 249 77 250
rect 75 249 76 250
rect 74 249 75 250
rect 73 249 74 250
rect 72 249 73 250
rect 71 249 72 250
rect 70 249 71 250
rect 69 249 70 250
rect 68 249 69 250
rect 67 249 68 250
rect 66 249 67 250
rect 65 249 66 250
rect 64 249 65 250
rect 63 249 64 250
rect 62 249 63 250
rect 61 249 62 250
rect 27 249 28 250
rect 26 249 27 250
rect 22 249 23 250
rect 21 249 22 250
rect 20 249 21 250
rect 19 249 20 250
rect 198 250 199 251
rect 197 250 198 251
rect 196 250 197 251
rect 195 250 196 251
rect 194 250 195 251
rect 193 250 194 251
rect 176 250 177 251
rect 175 250 176 251
rect 174 250 175 251
rect 167 250 168 251
rect 166 250 167 251
rect 165 250 166 251
rect 151 250 152 251
rect 150 250 151 251
rect 149 250 150 251
rect 148 250 149 251
rect 147 250 148 251
rect 146 250 147 251
rect 145 250 146 251
rect 144 250 145 251
rect 143 250 144 251
rect 142 250 143 251
rect 132 250 133 251
rect 131 250 132 251
rect 130 250 131 251
rect 129 250 130 251
rect 128 250 129 251
rect 127 250 128 251
rect 126 250 127 251
rect 125 250 126 251
rect 124 250 125 251
rect 123 250 124 251
rect 114 250 115 251
rect 113 250 114 251
rect 112 250 113 251
rect 111 250 112 251
rect 110 250 111 251
rect 109 250 110 251
rect 108 250 109 251
rect 107 250 108 251
rect 106 250 107 251
rect 105 250 106 251
rect 104 250 105 251
rect 88 250 89 251
rect 87 250 88 251
rect 86 250 87 251
rect 85 250 86 251
rect 84 250 85 251
rect 83 250 84 251
rect 82 250 83 251
rect 81 250 82 251
rect 80 250 81 251
rect 79 250 80 251
rect 78 250 79 251
rect 77 250 78 251
rect 76 250 77 251
rect 75 250 76 251
rect 74 250 75 251
rect 73 250 74 251
rect 72 250 73 251
rect 71 250 72 251
rect 70 250 71 251
rect 69 250 70 251
rect 68 250 69 251
rect 67 250 68 251
rect 66 250 67 251
rect 65 250 66 251
rect 64 250 65 251
rect 63 250 64 251
rect 62 250 63 251
rect 61 250 62 251
rect 194 251 195 252
rect 193 251 194 252
rect 176 251 177 252
rect 175 251 176 252
rect 174 251 175 252
rect 173 251 174 252
rect 167 251 168 252
rect 166 251 167 252
rect 165 251 166 252
rect 151 251 152 252
rect 150 251 151 252
rect 149 251 150 252
rect 148 251 149 252
rect 147 251 148 252
rect 146 251 147 252
rect 145 251 146 252
rect 144 251 145 252
rect 143 251 144 252
rect 142 251 143 252
rect 132 251 133 252
rect 131 251 132 252
rect 130 251 131 252
rect 129 251 130 252
rect 128 251 129 252
rect 127 251 128 252
rect 126 251 127 252
rect 125 251 126 252
rect 124 251 125 252
rect 123 251 124 252
rect 114 251 115 252
rect 113 251 114 252
rect 112 251 113 252
rect 111 251 112 252
rect 110 251 111 252
rect 109 251 110 252
rect 108 251 109 252
rect 107 251 108 252
rect 106 251 107 252
rect 105 251 106 252
rect 104 251 105 252
rect 78 251 79 252
rect 77 251 78 252
rect 76 251 77 252
rect 75 251 76 252
rect 74 251 75 252
rect 73 251 74 252
rect 72 251 73 252
rect 68 251 69 252
rect 67 251 68 252
rect 66 251 67 252
rect 65 251 66 252
rect 64 251 65 252
rect 63 251 64 252
rect 198 252 199 253
rect 197 252 198 253
rect 196 252 197 253
rect 195 252 196 253
rect 194 252 195 253
rect 193 252 194 253
rect 176 252 177 253
rect 175 252 176 253
rect 174 252 175 253
rect 173 252 174 253
rect 172 252 173 253
rect 167 252 168 253
rect 166 252 167 253
rect 165 252 166 253
rect 151 252 152 253
rect 150 252 151 253
rect 149 252 150 253
rect 148 252 149 253
rect 147 252 148 253
rect 146 252 147 253
rect 145 252 146 253
rect 144 252 145 253
rect 143 252 144 253
rect 142 252 143 253
rect 132 252 133 253
rect 131 252 132 253
rect 130 252 131 253
rect 129 252 130 253
rect 128 252 129 253
rect 127 252 128 253
rect 126 252 127 253
rect 125 252 126 253
rect 124 252 125 253
rect 123 252 124 253
rect 114 252 115 253
rect 113 252 114 253
rect 112 252 113 253
rect 111 252 112 253
rect 110 252 111 253
rect 109 252 110 253
rect 108 252 109 253
rect 107 252 108 253
rect 106 252 107 253
rect 105 252 106 253
rect 104 252 105 253
rect 79 252 80 253
rect 78 252 79 253
rect 77 252 78 253
rect 76 252 77 253
rect 75 252 76 253
rect 65 252 66 253
rect 64 252 65 253
rect 63 252 64 253
rect 62 252 63 253
rect 199 253 200 254
rect 198 253 199 254
rect 197 253 198 254
rect 196 253 197 254
rect 195 253 196 254
rect 194 253 195 254
rect 193 253 194 254
rect 184 253 185 254
rect 183 253 184 254
rect 182 253 183 254
rect 181 253 182 254
rect 180 253 181 254
rect 179 253 180 254
rect 178 253 179 254
rect 175 253 176 254
rect 174 253 175 254
rect 173 253 174 254
rect 172 253 173 254
rect 171 253 172 254
rect 167 253 168 254
rect 166 253 167 254
rect 165 253 166 254
rect 151 253 152 254
rect 150 253 151 254
rect 149 253 150 254
rect 148 253 149 254
rect 147 253 148 254
rect 146 253 147 254
rect 145 253 146 254
rect 144 253 145 254
rect 143 253 144 254
rect 142 253 143 254
rect 132 253 133 254
rect 131 253 132 254
rect 130 253 131 254
rect 129 253 130 254
rect 128 253 129 254
rect 127 253 128 254
rect 126 253 127 254
rect 125 253 126 254
rect 124 253 125 254
rect 123 253 124 254
rect 114 253 115 254
rect 113 253 114 254
rect 112 253 113 254
rect 111 253 112 254
rect 110 253 111 254
rect 109 253 110 254
rect 108 253 109 254
rect 107 253 108 254
rect 106 253 107 254
rect 105 253 106 254
rect 104 253 105 254
rect 79 253 80 254
rect 78 253 79 254
rect 77 253 78 254
rect 76 253 77 254
rect 64 253 65 254
rect 63 253 64 254
rect 62 253 63 254
rect 61 253 62 254
rect 198 254 199 255
rect 197 254 198 255
rect 196 254 197 255
rect 195 254 196 255
rect 194 254 195 255
rect 185 254 186 255
rect 184 254 185 255
rect 183 254 184 255
rect 182 254 183 255
rect 181 254 182 255
rect 180 254 181 255
rect 179 254 180 255
rect 178 254 179 255
rect 175 254 176 255
rect 174 254 175 255
rect 173 254 174 255
rect 172 254 173 255
rect 171 254 172 255
rect 170 254 171 255
rect 167 254 168 255
rect 166 254 167 255
rect 165 254 166 255
rect 80 254 81 255
rect 79 254 80 255
rect 78 254 79 255
rect 77 254 78 255
rect 64 254 65 255
rect 63 254 64 255
rect 62 254 63 255
rect 61 254 62 255
rect 197 255 198 256
rect 196 255 197 256
rect 195 255 196 256
rect 185 255 186 256
rect 184 255 185 256
rect 183 255 184 256
rect 182 255 183 256
rect 181 255 182 256
rect 180 255 181 256
rect 179 255 180 256
rect 178 255 179 256
rect 174 255 175 256
rect 173 255 174 256
rect 172 255 173 256
rect 171 255 172 256
rect 170 255 171 256
rect 169 255 170 256
rect 168 255 169 256
rect 167 255 168 256
rect 166 255 167 256
rect 165 255 166 256
rect 80 255 81 256
rect 79 255 80 256
rect 78 255 79 256
rect 77 255 78 256
rect 64 255 65 256
rect 63 255 64 256
rect 62 255 63 256
rect 61 255 62 256
rect 198 256 199 257
rect 197 256 198 257
rect 196 256 197 257
rect 195 256 196 257
rect 194 256 195 257
rect 193 256 194 257
rect 185 256 186 257
rect 184 256 185 257
rect 183 256 184 257
rect 182 256 183 257
rect 181 256 182 257
rect 180 256 181 257
rect 179 256 180 257
rect 178 256 179 257
rect 173 256 174 257
rect 172 256 173 257
rect 171 256 172 257
rect 170 256 171 257
rect 169 256 170 257
rect 168 256 169 257
rect 167 256 168 257
rect 166 256 167 257
rect 165 256 166 257
rect 80 256 81 257
rect 79 256 80 257
rect 78 256 79 257
rect 77 256 78 257
rect 64 256 65 257
rect 63 256 64 257
rect 62 256 63 257
rect 61 256 62 257
rect 60 256 61 257
rect 198 257 199 258
rect 197 257 198 258
rect 196 257 197 258
rect 195 257 196 258
rect 194 257 195 258
rect 193 257 194 258
rect 185 257 186 258
rect 184 257 185 258
rect 183 257 184 258
rect 182 257 183 258
rect 173 257 174 258
rect 172 257 173 258
rect 171 257 172 258
rect 170 257 171 258
rect 169 257 170 258
rect 168 257 169 258
rect 167 257 168 258
rect 166 257 167 258
rect 165 257 166 258
rect 80 257 81 258
rect 79 257 80 258
rect 78 257 79 258
rect 77 257 78 258
rect 64 257 65 258
rect 63 257 64 258
rect 62 257 63 258
rect 61 257 62 258
rect 60 257 61 258
rect 31 257 32 258
rect 30 257 31 258
rect 29 257 30 258
rect 28 257 29 258
rect 199 258 200 259
rect 198 258 199 259
rect 194 258 195 259
rect 193 258 194 259
rect 185 258 186 259
rect 184 258 185 259
rect 183 258 184 259
rect 182 258 183 259
rect 174 258 175 259
rect 173 258 174 259
rect 172 258 173 259
rect 171 258 172 259
rect 170 258 171 259
rect 169 258 170 259
rect 168 258 169 259
rect 167 258 168 259
rect 166 258 167 259
rect 165 258 166 259
rect 80 258 81 259
rect 79 258 80 259
rect 78 258 79 259
rect 77 258 78 259
rect 76 258 77 259
rect 65 258 66 259
rect 64 258 65 259
rect 63 258 64 259
rect 62 258 63 259
rect 61 258 62 259
rect 60 258 61 259
rect 31 258 32 259
rect 30 258 31 259
rect 29 258 30 259
rect 28 258 29 259
rect 27 258 28 259
rect 26 258 27 259
rect 25 258 26 259
rect 24 258 25 259
rect 23 258 24 259
rect 199 259 200 260
rect 198 259 199 260
rect 197 259 198 260
rect 196 259 197 260
rect 195 259 196 260
rect 194 259 195 260
rect 193 259 194 260
rect 192 259 193 260
rect 191 259 192 260
rect 190 259 191 260
rect 185 259 186 260
rect 184 259 185 260
rect 183 259 184 260
rect 182 259 183 260
rect 174 259 175 260
rect 173 259 174 260
rect 172 259 173 260
rect 171 259 172 260
rect 170 259 171 260
rect 167 259 168 260
rect 166 259 167 260
rect 165 259 166 260
rect 80 259 81 260
rect 79 259 80 260
rect 78 259 79 260
rect 77 259 78 260
rect 76 259 77 260
rect 75 259 76 260
rect 74 259 75 260
rect 67 259 68 260
rect 66 259 67 260
rect 65 259 66 260
rect 64 259 65 260
rect 63 259 64 260
rect 62 259 63 260
rect 61 259 62 260
rect 31 259 32 260
rect 30 259 31 260
rect 29 259 30 260
rect 28 259 29 260
rect 27 259 28 260
rect 26 259 27 260
rect 25 259 26 260
rect 24 259 25 260
rect 23 259 24 260
rect 22 259 23 260
rect 21 259 22 260
rect 20 259 21 260
rect 19 259 20 260
rect 18 259 19 260
rect 199 260 200 261
rect 198 260 199 261
rect 197 260 198 261
rect 196 260 197 261
rect 195 260 196 261
rect 194 260 195 261
rect 193 260 194 261
rect 192 260 193 261
rect 191 260 192 261
rect 190 260 191 261
rect 185 260 186 261
rect 184 260 185 261
rect 183 260 184 261
rect 182 260 183 261
rect 175 260 176 261
rect 174 260 175 261
rect 173 260 174 261
rect 172 260 173 261
rect 167 260 168 261
rect 166 260 167 261
rect 165 260 166 261
rect 80 260 81 261
rect 79 260 80 261
rect 78 260 79 261
rect 77 260 78 261
rect 76 260 77 261
rect 75 260 76 261
rect 74 260 75 261
rect 73 260 74 261
rect 72 260 73 261
rect 71 260 72 261
rect 70 260 71 261
rect 69 260 70 261
rect 68 260 69 261
rect 67 260 68 261
rect 66 260 67 261
rect 65 260 66 261
rect 64 260 65 261
rect 63 260 64 261
rect 62 260 63 261
rect 61 260 62 261
rect 28 260 29 261
rect 27 260 28 261
rect 26 260 27 261
rect 25 260 26 261
rect 24 260 25 261
rect 23 260 24 261
rect 22 260 23 261
rect 21 260 22 261
rect 20 260 21 261
rect 19 260 20 261
rect 18 260 19 261
rect 17 260 18 261
rect 16 260 17 261
rect 198 261 199 262
rect 197 261 198 262
rect 196 261 197 262
rect 195 261 196 262
rect 194 261 195 262
rect 193 261 194 262
rect 192 261 193 262
rect 191 261 192 262
rect 190 261 191 262
rect 185 261 186 262
rect 184 261 185 262
rect 183 261 184 262
rect 182 261 183 262
rect 175 261 176 262
rect 174 261 175 262
rect 173 261 174 262
rect 172 261 173 262
rect 167 261 168 262
rect 166 261 167 262
rect 165 261 166 262
rect 79 261 80 262
rect 78 261 79 262
rect 77 261 78 262
rect 76 261 77 262
rect 75 261 76 262
rect 74 261 75 262
rect 73 261 74 262
rect 72 261 73 262
rect 71 261 72 262
rect 70 261 71 262
rect 69 261 70 262
rect 68 261 69 262
rect 67 261 68 262
rect 66 261 67 262
rect 65 261 66 262
rect 64 261 65 262
rect 63 261 64 262
rect 62 261 63 262
rect 22 261 23 262
rect 21 261 22 262
rect 20 261 21 262
rect 19 261 20 262
rect 18 261 19 262
rect 17 261 18 262
rect 16 261 17 262
rect 185 262 186 263
rect 184 262 185 263
rect 183 262 184 263
rect 182 262 183 263
rect 176 262 177 263
rect 175 262 176 263
rect 174 262 175 263
rect 173 262 174 263
rect 167 262 168 263
rect 166 262 167 263
rect 165 262 166 263
rect 78 262 79 263
rect 77 262 78 263
rect 76 262 77 263
rect 75 262 76 263
rect 74 262 75 263
rect 73 262 74 263
rect 72 262 73 263
rect 71 262 72 263
rect 70 262 71 263
rect 69 262 70 263
rect 68 262 69 263
rect 67 262 68 263
rect 66 262 67 263
rect 65 262 66 263
rect 64 262 65 263
rect 63 262 64 263
rect 31 262 32 263
rect 30 262 31 263
rect 29 262 30 263
rect 28 262 29 263
rect 27 262 28 263
rect 26 262 27 263
rect 25 262 26 263
rect 24 262 25 263
rect 23 262 24 263
rect 22 262 23 263
rect 21 262 22 263
rect 20 262 21 263
rect 19 262 20 263
rect 18 262 19 263
rect 17 262 18 263
rect 16 262 17 263
rect 185 263 186 264
rect 184 263 185 264
rect 183 263 184 264
rect 182 263 183 264
rect 175 263 176 264
rect 174 263 175 264
rect 171 263 172 264
rect 170 263 171 264
rect 169 263 170 264
rect 168 263 169 264
rect 167 263 168 264
rect 166 263 167 264
rect 165 263 166 264
rect 77 263 78 264
rect 76 263 77 264
rect 75 263 76 264
rect 74 263 75 264
rect 73 263 74 264
rect 72 263 73 264
rect 71 263 72 264
rect 70 263 71 264
rect 69 263 70 264
rect 68 263 69 264
rect 67 263 68 264
rect 66 263 67 264
rect 65 263 66 264
rect 64 263 65 264
rect 31 263 32 264
rect 30 263 31 264
rect 29 263 30 264
rect 28 263 29 264
rect 27 263 28 264
rect 26 263 27 264
rect 25 263 26 264
rect 24 263 25 264
rect 23 263 24 264
rect 22 263 23 264
rect 21 263 22 264
rect 20 263 21 264
rect 19 263 20 264
rect 18 263 19 264
rect 17 263 18 264
rect 16 263 17 264
rect 185 264 186 265
rect 184 264 185 265
rect 183 264 184 265
rect 182 264 183 265
rect 174 264 175 265
rect 171 264 172 265
rect 170 264 171 265
rect 169 264 170 265
rect 168 264 169 265
rect 75 264 76 265
rect 74 264 75 265
rect 73 264 74 265
rect 72 264 73 265
rect 71 264 72 265
rect 70 264 71 265
rect 69 264 70 265
rect 68 264 69 265
rect 67 264 68 265
rect 66 264 67 265
rect 65 264 66 265
rect 31 264 32 265
rect 30 264 31 265
rect 29 264 30 265
rect 28 264 29 265
rect 27 264 28 265
rect 26 264 27 265
rect 25 264 26 265
rect 24 264 25 265
rect 23 264 24 265
rect 22 264 23 265
rect 21 264 22 265
rect 20 264 21 265
rect 19 264 20 265
rect 18 264 19 265
rect 17 264 18 265
rect 191 265 192 266
rect 185 265 186 266
rect 184 265 185 266
rect 183 265 184 266
rect 182 265 183 266
rect 171 265 172 266
rect 170 265 171 266
rect 169 265 170 266
rect 168 265 169 266
rect 71 265 72 266
rect 70 265 71 266
rect 69 265 70 266
rect 31 265 32 266
rect 30 265 31 266
rect 29 265 30 266
rect 28 265 29 266
rect 27 265 28 266
rect 26 265 27 266
rect 25 265 26 266
rect 191 266 192 267
rect 185 266 186 267
rect 184 266 185 267
rect 183 266 184 267
rect 182 266 183 267
rect 171 266 172 267
rect 170 266 171 267
rect 169 266 170 267
rect 168 266 169 267
rect 29 266 30 267
rect 28 266 29 267
rect 27 266 28 267
rect 26 266 27 267
rect 25 266 26 267
rect 24 266 25 267
rect 23 266 24 267
rect 192 267 193 268
rect 191 267 192 268
rect 185 267 186 268
rect 184 267 185 268
rect 183 267 184 268
rect 182 267 183 268
rect 179 267 180 268
rect 178 267 179 268
rect 177 267 178 268
rect 176 267 177 268
rect 175 267 176 268
rect 174 267 175 268
rect 173 267 174 268
rect 172 267 173 268
rect 171 267 172 268
rect 170 267 171 268
rect 169 267 170 268
rect 168 267 169 268
rect 167 267 168 268
rect 166 267 167 268
rect 165 267 166 268
rect 164 267 165 268
rect 114 267 115 268
rect 113 267 114 268
rect 112 267 113 268
rect 111 267 112 268
rect 110 267 111 268
rect 109 267 110 268
rect 108 267 109 268
rect 107 267 108 268
rect 106 267 107 268
rect 105 267 106 268
rect 104 267 105 268
rect 27 267 28 268
rect 26 267 27 268
rect 25 267 26 268
rect 24 267 25 268
rect 23 267 24 268
rect 22 267 23 268
rect 21 267 22 268
rect 199 268 200 269
rect 198 268 199 269
rect 197 268 198 269
rect 196 268 197 269
rect 195 268 196 269
rect 194 268 195 269
rect 193 268 194 269
rect 192 268 193 269
rect 191 268 192 269
rect 185 268 186 269
rect 184 268 185 269
rect 183 268 184 269
rect 182 268 183 269
rect 179 268 180 269
rect 178 268 179 269
rect 177 268 178 269
rect 176 268 177 269
rect 175 268 176 269
rect 174 268 175 269
rect 173 268 174 269
rect 172 268 173 269
rect 171 268 172 269
rect 170 268 171 269
rect 169 268 170 269
rect 168 268 169 269
rect 167 268 168 269
rect 166 268 167 269
rect 165 268 166 269
rect 164 268 165 269
rect 114 268 115 269
rect 113 268 114 269
rect 112 268 113 269
rect 111 268 112 269
rect 110 268 111 269
rect 109 268 110 269
rect 108 268 109 269
rect 107 268 108 269
rect 106 268 107 269
rect 105 268 106 269
rect 104 268 105 269
rect 75 268 76 269
rect 74 268 75 269
rect 73 268 74 269
rect 72 268 73 269
rect 71 268 72 269
rect 70 268 71 269
rect 69 268 70 269
rect 68 268 69 269
rect 67 268 68 269
rect 66 268 67 269
rect 31 268 32 269
rect 24 268 25 269
rect 23 268 24 269
rect 22 268 23 269
rect 21 268 22 269
rect 20 268 21 269
rect 19 268 20 269
rect 198 269 199 270
rect 197 269 198 270
rect 196 269 197 270
rect 195 269 196 270
rect 194 269 195 270
rect 193 269 194 270
rect 192 269 193 270
rect 191 269 192 270
rect 185 269 186 270
rect 184 269 185 270
rect 183 269 184 270
rect 182 269 183 270
rect 179 269 180 270
rect 178 269 179 270
rect 177 269 178 270
rect 176 269 177 270
rect 175 269 176 270
rect 174 269 175 270
rect 173 269 174 270
rect 172 269 173 270
rect 171 269 172 270
rect 170 269 171 270
rect 169 269 170 270
rect 168 269 169 270
rect 167 269 168 270
rect 166 269 167 270
rect 165 269 166 270
rect 164 269 165 270
rect 114 269 115 270
rect 113 269 114 270
rect 112 269 113 270
rect 111 269 112 270
rect 110 269 111 270
rect 109 269 110 270
rect 108 269 109 270
rect 107 269 108 270
rect 106 269 107 270
rect 105 269 106 270
rect 104 269 105 270
rect 77 269 78 270
rect 76 269 77 270
rect 75 269 76 270
rect 74 269 75 270
rect 73 269 74 270
rect 72 269 73 270
rect 71 269 72 270
rect 70 269 71 270
rect 69 269 70 270
rect 68 269 69 270
rect 67 269 68 270
rect 66 269 67 270
rect 65 269 66 270
rect 64 269 65 270
rect 31 269 32 270
rect 30 269 31 270
rect 29 269 30 270
rect 28 269 29 270
rect 27 269 28 270
rect 26 269 27 270
rect 22 269 23 270
rect 21 269 22 270
rect 20 269 21 270
rect 19 269 20 270
rect 18 269 19 270
rect 17 269 18 270
rect 191 270 192 271
rect 185 270 186 271
rect 184 270 185 271
rect 183 270 184 271
rect 182 270 183 271
rect 179 270 180 271
rect 178 270 179 271
rect 177 270 178 271
rect 176 270 177 271
rect 175 270 176 271
rect 174 270 175 271
rect 173 270 174 271
rect 172 270 173 271
rect 171 270 172 271
rect 170 270 171 271
rect 169 270 170 271
rect 168 270 169 271
rect 167 270 168 271
rect 166 270 167 271
rect 165 270 166 271
rect 164 270 165 271
rect 114 270 115 271
rect 113 270 114 271
rect 112 270 113 271
rect 111 270 112 271
rect 110 270 111 271
rect 109 270 110 271
rect 108 270 109 271
rect 107 270 108 271
rect 106 270 107 271
rect 105 270 106 271
rect 104 270 105 271
rect 78 270 79 271
rect 77 270 78 271
rect 76 270 77 271
rect 75 270 76 271
rect 74 270 75 271
rect 73 270 74 271
rect 72 270 73 271
rect 71 270 72 271
rect 70 270 71 271
rect 69 270 70 271
rect 68 270 69 271
rect 67 270 68 271
rect 66 270 67 271
rect 65 270 66 271
rect 64 270 65 271
rect 63 270 64 271
rect 31 270 32 271
rect 30 270 31 271
rect 29 270 30 271
rect 28 270 29 271
rect 27 270 28 271
rect 26 270 27 271
rect 25 270 26 271
rect 24 270 25 271
rect 23 270 24 271
rect 22 270 23 271
rect 21 270 22 271
rect 20 270 21 271
rect 19 270 20 271
rect 18 270 19 271
rect 17 270 18 271
rect 16 270 17 271
rect 197 271 198 272
rect 196 271 197 272
rect 195 271 196 272
rect 194 271 195 272
rect 191 271 192 272
rect 184 271 185 272
rect 183 271 184 272
rect 114 271 115 272
rect 113 271 114 272
rect 112 271 113 272
rect 111 271 112 272
rect 110 271 111 272
rect 109 271 110 272
rect 108 271 109 272
rect 107 271 108 272
rect 106 271 107 272
rect 105 271 106 272
rect 104 271 105 272
rect 79 271 80 272
rect 78 271 79 272
rect 77 271 78 272
rect 76 271 77 272
rect 75 271 76 272
rect 74 271 75 272
rect 73 271 74 272
rect 72 271 73 272
rect 71 271 72 272
rect 70 271 71 272
rect 69 271 70 272
rect 68 271 69 272
rect 67 271 68 272
rect 66 271 67 272
rect 65 271 66 272
rect 64 271 65 272
rect 63 271 64 272
rect 62 271 63 272
rect 30 271 31 272
rect 29 271 30 272
rect 28 271 29 272
rect 27 271 28 272
rect 26 271 27 272
rect 25 271 26 272
rect 24 271 25 272
rect 23 271 24 272
rect 22 271 23 272
rect 21 271 22 272
rect 20 271 21 272
rect 19 271 20 272
rect 18 271 19 272
rect 17 271 18 272
rect 16 271 17 272
rect 198 272 199 273
rect 197 272 198 273
rect 196 272 197 273
rect 195 272 196 273
rect 194 272 195 273
rect 193 272 194 273
rect 114 272 115 273
rect 113 272 114 273
rect 112 272 113 273
rect 111 272 112 273
rect 110 272 111 273
rect 109 272 110 273
rect 108 272 109 273
rect 107 272 108 273
rect 106 272 107 273
rect 105 272 106 273
rect 104 272 105 273
rect 79 272 80 273
rect 78 272 79 273
rect 77 272 78 273
rect 76 272 77 273
rect 75 272 76 273
rect 74 272 75 273
rect 73 272 74 273
rect 72 272 73 273
rect 71 272 72 273
rect 70 272 71 273
rect 69 272 70 273
rect 68 272 69 273
rect 67 272 68 273
rect 66 272 67 273
rect 65 272 66 273
rect 64 272 65 273
rect 63 272 64 273
rect 62 272 63 273
rect 25 272 26 273
rect 24 272 25 273
rect 23 272 24 273
rect 22 272 23 273
rect 21 272 22 273
rect 20 272 21 273
rect 19 272 20 273
rect 18 272 19 273
rect 17 272 18 273
rect 16 272 17 273
rect 199 273 200 274
rect 198 273 199 274
rect 197 273 198 274
rect 196 273 197 274
rect 195 273 196 274
rect 194 273 195 274
rect 193 273 194 274
rect 114 273 115 274
rect 113 273 114 274
rect 112 273 113 274
rect 111 273 112 274
rect 110 273 111 274
rect 109 273 110 274
rect 108 273 109 274
rect 107 273 108 274
rect 106 273 107 274
rect 105 273 106 274
rect 104 273 105 274
rect 80 273 81 274
rect 79 273 80 274
rect 78 273 79 274
rect 77 273 78 274
rect 76 273 77 274
rect 75 273 76 274
rect 74 273 75 274
rect 73 273 74 274
rect 72 273 73 274
rect 71 273 72 274
rect 70 273 71 274
rect 69 273 70 274
rect 68 273 69 274
rect 67 273 68 274
rect 66 273 67 274
rect 65 273 66 274
rect 64 273 65 274
rect 63 273 64 274
rect 62 273 63 274
rect 61 273 62 274
rect 20 273 21 274
rect 19 273 20 274
rect 18 273 19 274
rect 17 273 18 274
rect 16 273 17 274
rect 199 274 200 275
rect 198 274 199 275
rect 196 274 197 275
rect 194 274 195 275
rect 193 274 194 275
rect 114 274 115 275
rect 113 274 114 275
rect 112 274 113 275
rect 111 274 112 275
rect 110 274 111 275
rect 109 274 110 275
rect 108 274 109 275
rect 107 274 108 275
rect 106 274 107 275
rect 105 274 106 275
rect 104 274 105 275
rect 80 274 81 275
rect 79 274 80 275
rect 78 274 79 275
rect 77 274 78 275
rect 76 274 77 275
rect 72 274 73 275
rect 71 274 72 275
rect 70 274 71 275
rect 69 274 70 275
rect 65 274 66 275
rect 64 274 65 275
rect 63 274 64 275
rect 62 274 63 275
rect 61 274 62 275
rect 35 274 36 275
rect 34 274 35 275
rect 199 275 200 276
rect 198 275 199 276
rect 196 275 197 276
rect 195 275 196 276
rect 194 275 195 276
rect 193 275 194 276
rect 114 275 115 276
rect 113 275 114 276
rect 112 275 113 276
rect 111 275 112 276
rect 110 275 111 276
rect 109 275 110 276
rect 108 275 109 276
rect 107 275 108 276
rect 106 275 107 276
rect 105 275 106 276
rect 104 275 105 276
rect 80 275 81 276
rect 79 275 80 276
rect 78 275 79 276
rect 77 275 78 276
rect 76 275 77 276
rect 72 275 73 276
rect 71 275 72 276
rect 70 275 71 276
rect 69 275 70 276
rect 64 275 65 276
rect 63 275 64 276
rect 62 275 63 276
rect 61 275 62 276
rect 60 275 61 276
rect 35 275 36 276
rect 34 275 35 276
rect 21 275 22 276
rect 198 276 199 277
rect 196 276 197 277
rect 195 276 196 277
rect 194 276 195 277
rect 114 276 115 277
rect 113 276 114 277
rect 112 276 113 277
rect 111 276 112 277
rect 110 276 111 277
rect 109 276 110 277
rect 108 276 109 277
rect 107 276 108 277
rect 106 276 107 277
rect 105 276 106 277
rect 104 276 105 277
rect 80 276 81 277
rect 79 276 80 277
rect 78 276 79 277
rect 77 276 78 277
rect 72 276 73 277
rect 71 276 72 277
rect 70 276 71 277
rect 69 276 70 277
rect 64 276 65 277
rect 63 276 64 277
rect 62 276 63 277
rect 61 276 62 277
rect 60 276 61 277
rect 35 276 36 277
rect 34 276 35 277
rect 33 276 34 277
rect 27 276 28 277
rect 26 276 27 277
rect 25 276 26 277
rect 24 276 25 277
rect 23 276 24 277
rect 22 276 23 277
rect 21 276 22 277
rect 20 276 21 277
rect 114 277 115 278
rect 113 277 114 278
rect 112 277 113 278
rect 111 277 112 278
rect 110 277 111 278
rect 109 277 110 278
rect 108 277 109 278
rect 107 277 108 278
rect 106 277 107 278
rect 105 277 106 278
rect 104 277 105 278
rect 80 277 81 278
rect 79 277 80 278
rect 78 277 79 278
rect 77 277 78 278
rect 72 277 73 278
rect 71 277 72 278
rect 70 277 71 278
rect 69 277 70 278
rect 64 277 65 278
rect 63 277 64 278
rect 62 277 63 278
rect 61 277 62 278
rect 60 277 61 278
rect 35 277 36 278
rect 34 277 35 278
rect 33 277 34 278
rect 32 277 33 278
rect 31 277 32 278
rect 30 277 31 278
rect 29 277 30 278
rect 28 277 29 278
rect 27 277 28 278
rect 26 277 27 278
rect 25 277 26 278
rect 24 277 25 278
rect 23 277 24 278
rect 22 277 23 278
rect 21 277 22 278
rect 20 277 21 278
rect 198 278 199 279
rect 197 278 198 279
rect 196 278 197 279
rect 195 278 196 279
rect 194 278 195 279
rect 193 278 194 279
rect 192 278 193 279
rect 191 278 192 279
rect 190 278 191 279
rect 114 278 115 279
rect 113 278 114 279
rect 112 278 113 279
rect 111 278 112 279
rect 110 278 111 279
rect 109 278 110 279
rect 108 278 109 279
rect 107 278 108 279
rect 106 278 107 279
rect 105 278 106 279
rect 104 278 105 279
rect 80 278 81 279
rect 79 278 80 279
rect 78 278 79 279
rect 77 278 78 279
rect 72 278 73 279
rect 71 278 72 279
rect 70 278 71 279
rect 69 278 70 279
rect 64 278 65 279
rect 63 278 64 279
rect 62 278 63 279
rect 61 278 62 279
rect 60 278 61 279
rect 34 278 35 279
rect 33 278 34 279
rect 32 278 33 279
rect 31 278 32 279
rect 30 278 31 279
rect 29 278 30 279
rect 28 278 29 279
rect 27 278 28 279
rect 26 278 27 279
rect 25 278 26 279
rect 24 278 25 279
rect 23 278 24 279
rect 22 278 23 279
rect 21 278 22 279
rect 198 279 199 280
rect 197 279 198 280
rect 196 279 197 280
rect 195 279 196 280
rect 194 279 195 280
rect 193 279 194 280
rect 192 279 193 280
rect 191 279 192 280
rect 190 279 191 280
rect 114 279 115 280
rect 113 279 114 280
rect 112 279 113 280
rect 111 279 112 280
rect 110 279 111 280
rect 109 279 110 280
rect 108 279 109 280
rect 107 279 108 280
rect 106 279 107 280
rect 105 279 106 280
rect 104 279 105 280
rect 80 279 81 280
rect 79 279 80 280
rect 78 279 79 280
rect 77 279 78 280
rect 72 279 73 280
rect 71 279 72 280
rect 70 279 71 280
rect 69 279 70 280
rect 64 279 65 280
rect 63 279 64 280
rect 62 279 63 280
rect 61 279 62 280
rect 33 279 34 280
rect 32 279 33 280
rect 31 279 32 280
rect 30 279 31 280
rect 29 279 30 280
rect 28 279 29 280
rect 27 279 28 280
rect 114 280 115 281
rect 113 280 114 281
rect 112 280 113 281
rect 111 280 112 281
rect 110 280 111 281
rect 109 280 110 281
rect 108 280 109 281
rect 107 280 108 281
rect 106 280 107 281
rect 105 280 106 281
rect 104 280 105 281
rect 80 280 81 281
rect 79 280 80 281
rect 78 280 79 281
rect 77 280 78 281
rect 76 280 77 281
rect 75 280 76 281
rect 72 280 73 281
rect 71 280 72 281
rect 70 280 71 281
rect 69 280 70 281
rect 66 280 67 281
rect 65 280 66 281
rect 64 280 65 281
rect 63 280 64 281
rect 62 280 63 281
rect 61 280 62 281
rect 31 280 32 281
rect 30 280 31 281
rect 29 280 30 281
rect 28 280 29 281
rect 27 280 28 281
rect 26 280 27 281
rect 198 281 199 282
rect 197 281 198 282
rect 196 281 197 282
rect 195 281 196 282
rect 194 281 195 282
rect 114 281 115 282
rect 113 281 114 282
rect 112 281 113 282
rect 111 281 112 282
rect 110 281 111 282
rect 109 281 110 282
rect 108 281 109 282
rect 107 281 108 282
rect 106 281 107 282
rect 105 281 106 282
rect 104 281 105 282
rect 80 281 81 282
rect 79 281 80 282
rect 78 281 79 282
rect 77 281 78 282
rect 76 281 77 282
rect 75 281 76 282
rect 74 281 75 282
rect 72 281 73 282
rect 71 281 72 282
rect 70 281 71 282
rect 69 281 70 282
rect 68 281 69 282
rect 67 281 68 282
rect 66 281 67 282
rect 65 281 66 282
rect 64 281 65 282
rect 63 281 64 282
rect 62 281 63 282
rect 61 281 62 282
rect 30 281 31 282
rect 29 281 30 282
rect 28 281 29 282
rect 27 281 28 282
rect 26 281 27 282
rect 25 281 26 282
rect 24 281 25 282
rect 198 282 199 283
rect 197 282 198 283
rect 196 282 197 283
rect 195 282 196 283
rect 194 282 195 283
rect 193 282 194 283
rect 180 282 181 283
rect 114 282 115 283
rect 113 282 114 283
rect 112 282 113 283
rect 111 282 112 283
rect 110 282 111 283
rect 109 282 110 283
rect 108 282 109 283
rect 107 282 108 283
rect 106 282 107 283
rect 105 282 106 283
rect 104 282 105 283
rect 79 282 80 283
rect 78 282 79 283
rect 77 282 78 283
rect 76 282 77 283
rect 75 282 76 283
rect 72 282 73 283
rect 71 282 72 283
rect 70 282 71 283
rect 69 282 70 283
rect 68 282 69 283
rect 67 282 68 283
rect 66 282 67 283
rect 65 282 66 283
rect 64 282 65 283
rect 63 282 64 283
rect 62 282 63 283
rect 28 282 29 283
rect 27 282 28 283
rect 26 282 27 283
rect 25 282 26 283
rect 24 282 25 283
rect 23 282 24 283
rect 22 282 23 283
rect 199 283 200 284
rect 198 283 199 284
rect 196 283 197 284
rect 195 283 196 284
rect 194 283 195 284
rect 193 283 194 284
rect 181 283 182 284
rect 180 283 181 284
rect 179 283 180 284
rect 168 283 169 284
rect 114 283 115 284
rect 113 283 114 284
rect 112 283 113 284
rect 111 283 112 284
rect 110 283 111 284
rect 109 283 110 284
rect 108 283 109 284
rect 107 283 108 284
rect 106 283 107 284
rect 105 283 106 284
rect 104 283 105 284
rect 79 283 80 284
rect 78 283 79 284
rect 77 283 78 284
rect 76 283 77 284
rect 75 283 76 284
rect 72 283 73 284
rect 71 283 72 284
rect 70 283 71 284
rect 69 283 70 284
rect 68 283 69 284
rect 67 283 68 284
rect 66 283 67 284
rect 65 283 66 284
rect 64 283 65 284
rect 63 283 64 284
rect 26 283 27 284
rect 25 283 26 284
rect 24 283 25 284
rect 23 283 24 284
rect 22 283 23 284
rect 21 283 22 284
rect 199 284 200 285
rect 198 284 199 285
rect 196 284 197 285
rect 194 284 195 285
rect 193 284 194 285
rect 181 284 182 285
rect 180 284 181 285
rect 179 284 180 285
rect 178 284 179 285
rect 168 284 169 285
rect 167 284 168 285
rect 166 284 167 285
rect 114 284 115 285
rect 113 284 114 285
rect 112 284 113 285
rect 111 284 112 285
rect 110 284 111 285
rect 109 284 110 285
rect 108 284 109 285
rect 107 284 108 285
rect 106 284 107 285
rect 105 284 106 285
rect 104 284 105 285
rect 78 284 79 285
rect 77 284 78 285
rect 76 284 77 285
rect 75 284 76 285
rect 72 284 73 285
rect 71 284 72 285
rect 70 284 71 285
rect 69 284 70 285
rect 68 284 69 285
rect 67 284 68 285
rect 66 284 67 285
rect 65 284 66 285
rect 64 284 65 285
rect 24 284 25 285
rect 23 284 24 285
rect 22 284 23 285
rect 21 284 22 285
rect 20 284 21 285
rect 198 285 199 286
rect 196 285 197 286
rect 195 285 196 286
rect 194 285 195 286
rect 193 285 194 286
rect 181 285 182 286
rect 180 285 181 286
rect 179 285 180 286
rect 178 285 179 286
rect 177 285 178 286
rect 168 285 169 286
rect 167 285 168 286
rect 166 285 167 286
rect 114 285 115 286
rect 113 285 114 286
rect 112 285 113 286
rect 111 285 112 286
rect 110 285 111 286
rect 109 285 110 286
rect 108 285 109 286
rect 107 285 108 286
rect 106 285 107 286
rect 105 285 106 286
rect 104 285 105 286
rect 76 285 77 286
rect 75 285 76 286
rect 72 285 73 286
rect 71 285 72 286
rect 70 285 71 286
rect 69 285 70 286
rect 68 285 69 286
rect 67 285 68 286
rect 66 285 67 286
rect 65 285 66 286
rect 22 285 23 286
rect 21 285 22 286
rect 20 285 21 286
rect 198 286 199 287
rect 196 286 197 287
rect 195 286 196 287
rect 194 286 195 287
rect 181 286 182 287
rect 180 286 181 287
rect 179 286 180 287
rect 178 286 179 287
rect 177 286 178 287
rect 176 286 177 287
rect 168 286 169 287
rect 167 286 168 287
rect 166 286 167 287
rect 114 286 115 287
rect 113 286 114 287
rect 112 286 113 287
rect 111 286 112 287
rect 110 286 111 287
rect 109 286 110 287
rect 108 286 109 287
rect 107 286 108 287
rect 106 286 107 287
rect 105 286 106 287
rect 104 286 105 287
rect 71 286 72 287
rect 70 286 71 287
rect 69 286 70 287
rect 197 287 198 288
rect 196 287 197 288
rect 195 287 196 288
rect 180 287 181 288
rect 179 287 180 288
rect 178 287 179 288
rect 177 287 178 288
rect 176 287 177 288
rect 175 287 176 288
rect 168 287 169 288
rect 167 287 168 288
rect 166 287 167 288
rect 114 287 115 288
rect 113 287 114 288
rect 112 287 113 288
rect 111 287 112 288
rect 110 287 111 288
rect 109 287 110 288
rect 108 287 109 288
rect 107 287 108 288
rect 106 287 107 288
rect 105 287 106 288
rect 104 287 105 288
rect 198 288 199 289
rect 197 288 198 289
rect 196 288 197 289
rect 195 288 196 289
rect 194 288 195 289
rect 193 288 194 289
rect 179 288 180 289
rect 178 288 179 289
rect 177 288 178 289
rect 176 288 177 289
rect 175 288 176 289
rect 174 288 175 289
rect 173 288 174 289
rect 172 288 173 289
rect 171 288 172 289
rect 168 288 169 289
rect 167 288 168 289
rect 166 288 167 289
rect 114 288 115 289
rect 113 288 114 289
rect 112 288 113 289
rect 111 288 112 289
rect 110 288 111 289
rect 109 288 110 289
rect 108 288 109 289
rect 107 288 108 289
rect 106 288 107 289
rect 105 288 106 289
rect 104 288 105 289
rect 198 289 199 290
rect 197 289 198 290
rect 196 289 197 290
rect 195 289 196 290
rect 194 289 195 290
rect 193 289 194 290
rect 178 289 179 290
rect 177 289 178 290
rect 176 289 177 290
rect 175 289 176 290
rect 174 289 175 290
rect 173 289 174 290
rect 172 289 173 290
rect 171 289 172 290
rect 170 289 171 290
rect 169 289 170 290
rect 168 289 169 290
rect 167 289 168 290
rect 166 289 167 290
rect 114 289 115 290
rect 113 289 114 290
rect 112 289 113 290
rect 111 289 112 290
rect 110 289 111 290
rect 109 289 110 290
rect 108 289 109 290
rect 107 289 108 290
rect 106 289 107 290
rect 105 289 106 290
rect 104 289 105 290
rect 199 290 200 291
rect 198 290 199 291
rect 194 290 195 291
rect 193 290 194 291
rect 176 290 177 291
rect 175 290 176 291
rect 174 290 175 291
rect 173 290 174 291
rect 172 290 173 291
rect 171 290 172 291
rect 170 290 171 291
rect 169 290 170 291
rect 168 290 169 291
rect 167 290 168 291
rect 166 290 167 291
rect 114 290 115 291
rect 113 290 114 291
rect 112 290 113 291
rect 111 290 112 291
rect 110 290 111 291
rect 109 290 110 291
rect 108 290 109 291
rect 107 290 108 291
rect 106 290 107 291
rect 105 290 106 291
rect 104 290 105 291
rect 199 291 200 292
rect 198 291 199 292
rect 194 291 195 292
rect 193 291 194 292
rect 176 291 177 292
rect 175 291 176 292
rect 174 291 175 292
rect 173 291 174 292
rect 172 291 173 292
rect 171 291 172 292
rect 170 291 171 292
rect 169 291 170 292
rect 168 291 169 292
rect 167 291 168 292
rect 166 291 167 292
rect 114 291 115 292
rect 113 291 114 292
rect 112 291 113 292
rect 111 291 112 292
rect 110 291 111 292
rect 109 291 110 292
rect 108 291 109 292
rect 107 291 108 292
rect 106 291 107 292
rect 105 291 106 292
rect 104 291 105 292
rect 198 292 199 293
rect 197 292 198 293
rect 195 292 196 293
rect 178 292 179 293
rect 177 292 178 293
rect 176 292 177 293
rect 175 292 176 293
rect 174 292 175 293
rect 173 292 174 293
rect 172 292 173 293
rect 171 292 172 293
rect 170 292 171 293
rect 169 292 170 293
rect 168 292 169 293
rect 167 292 168 293
rect 166 292 167 293
rect 114 292 115 293
rect 113 292 114 293
rect 112 292 113 293
rect 111 292 112 293
rect 110 292 111 293
rect 109 292 110 293
rect 108 292 109 293
rect 107 292 108 293
rect 106 292 107 293
rect 105 292 106 293
rect 104 292 105 293
rect 198 293 199 294
rect 197 293 198 294
rect 196 293 197 294
rect 195 293 196 294
rect 194 293 195 294
rect 179 293 180 294
rect 178 293 179 294
rect 177 293 178 294
rect 176 293 177 294
rect 175 293 176 294
rect 174 293 175 294
rect 173 293 174 294
rect 168 293 169 294
rect 167 293 168 294
rect 166 293 167 294
rect 114 293 115 294
rect 113 293 114 294
rect 112 293 113 294
rect 111 293 112 294
rect 110 293 111 294
rect 109 293 110 294
rect 108 293 109 294
rect 107 293 108 294
rect 106 293 107 294
rect 105 293 106 294
rect 104 293 105 294
rect 27 293 28 294
rect 26 293 27 294
rect 25 293 26 294
rect 24 293 25 294
rect 23 293 24 294
rect 198 294 199 295
rect 197 294 198 295
rect 196 294 197 295
rect 195 294 196 295
rect 194 294 195 295
rect 193 294 194 295
rect 179 294 180 295
rect 178 294 179 295
rect 177 294 178 295
rect 176 294 177 295
rect 175 294 176 295
rect 168 294 169 295
rect 167 294 168 295
rect 166 294 167 295
rect 151 294 152 295
rect 150 294 151 295
rect 149 294 150 295
rect 148 294 149 295
rect 147 294 148 295
rect 146 294 147 295
rect 145 294 146 295
rect 144 294 145 295
rect 143 294 144 295
rect 142 294 143 295
rect 141 294 142 295
rect 140 294 141 295
rect 139 294 140 295
rect 138 294 139 295
rect 137 294 138 295
rect 136 294 137 295
rect 135 294 136 295
rect 134 294 135 295
rect 133 294 134 295
rect 132 294 133 295
rect 131 294 132 295
rect 130 294 131 295
rect 129 294 130 295
rect 128 294 129 295
rect 127 294 128 295
rect 126 294 127 295
rect 125 294 126 295
rect 124 294 125 295
rect 123 294 124 295
rect 122 294 123 295
rect 121 294 122 295
rect 120 294 121 295
rect 119 294 120 295
rect 118 294 119 295
rect 117 294 118 295
rect 116 294 117 295
rect 115 294 116 295
rect 114 294 115 295
rect 113 294 114 295
rect 112 294 113 295
rect 111 294 112 295
rect 110 294 111 295
rect 109 294 110 295
rect 108 294 109 295
rect 107 294 108 295
rect 106 294 107 295
rect 105 294 106 295
rect 104 294 105 295
rect 29 294 30 295
rect 28 294 29 295
rect 27 294 28 295
rect 26 294 27 295
rect 25 294 26 295
rect 24 294 25 295
rect 23 294 24 295
rect 22 294 23 295
rect 21 294 22 295
rect 20 294 21 295
rect 199 295 200 296
rect 198 295 199 296
rect 194 295 195 296
rect 193 295 194 296
rect 180 295 181 296
rect 179 295 180 296
rect 178 295 179 296
rect 177 295 178 296
rect 168 295 169 296
rect 167 295 168 296
rect 166 295 167 296
rect 151 295 152 296
rect 150 295 151 296
rect 149 295 150 296
rect 148 295 149 296
rect 147 295 148 296
rect 146 295 147 296
rect 145 295 146 296
rect 144 295 145 296
rect 143 295 144 296
rect 142 295 143 296
rect 141 295 142 296
rect 140 295 141 296
rect 139 295 140 296
rect 138 295 139 296
rect 137 295 138 296
rect 136 295 137 296
rect 135 295 136 296
rect 134 295 135 296
rect 133 295 134 296
rect 132 295 133 296
rect 131 295 132 296
rect 130 295 131 296
rect 129 295 130 296
rect 128 295 129 296
rect 127 295 128 296
rect 126 295 127 296
rect 125 295 126 296
rect 124 295 125 296
rect 123 295 124 296
rect 122 295 123 296
rect 121 295 122 296
rect 120 295 121 296
rect 119 295 120 296
rect 118 295 119 296
rect 117 295 118 296
rect 116 295 117 296
rect 115 295 116 296
rect 114 295 115 296
rect 113 295 114 296
rect 112 295 113 296
rect 111 295 112 296
rect 110 295 111 296
rect 109 295 110 296
rect 108 295 109 296
rect 107 295 108 296
rect 106 295 107 296
rect 105 295 106 296
rect 104 295 105 296
rect 30 295 31 296
rect 29 295 30 296
rect 28 295 29 296
rect 27 295 28 296
rect 26 295 27 296
rect 25 295 26 296
rect 24 295 25 296
rect 23 295 24 296
rect 22 295 23 296
rect 21 295 22 296
rect 20 295 21 296
rect 19 295 20 296
rect 199 296 200 297
rect 198 296 199 297
rect 194 296 195 297
rect 193 296 194 297
rect 181 296 182 297
rect 180 296 181 297
rect 179 296 180 297
rect 178 296 179 297
rect 177 296 178 297
rect 168 296 169 297
rect 167 296 168 297
rect 166 296 167 297
rect 151 296 152 297
rect 150 296 151 297
rect 149 296 150 297
rect 148 296 149 297
rect 147 296 148 297
rect 146 296 147 297
rect 145 296 146 297
rect 144 296 145 297
rect 143 296 144 297
rect 142 296 143 297
rect 141 296 142 297
rect 140 296 141 297
rect 139 296 140 297
rect 138 296 139 297
rect 137 296 138 297
rect 136 296 137 297
rect 135 296 136 297
rect 134 296 135 297
rect 133 296 134 297
rect 132 296 133 297
rect 131 296 132 297
rect 130 296 131 297
rect 129 296 130 297
rect 128 296 129 297
rect 127 296 128 297
rect 126 296 127 297
rect 125 296 126 297
rect 124 296 125 297
rect 123 296 124 297
rect 122 296 123 297
rect 121 296 122 297
rect 120 296 121 297
rect 119 296 120 297
rect 118 296 119 297
rect 117 296 118 297
rect 116 296 117 297
rect 115 296 116 297
rect 114 296 115 297
rect 113 296 114 297
rect 112 296 113 297
rect 111 296 112 297
rect 110 296 111 297
rect 109 296 110 297
rect 108 296 109 297
rect 107 296 108 297
rect 106 296 107 297
rect 105 296 106 297
rect 104 296 105 297
rect 31 296 32 297
rect 30 296 31 297
rect 29 296 30 297
rect 28 296 29 297
rect 27 296 28 297
rect 26 296 27 297
rect 25 296 26 297
rect 24 296 25 297
rect 23 296 24 297
rect 22 296 23 297
rect 21 296 22 297
rect 20 296 21 297
rect 19 296 20 297
rect 18 296 19 297
rect 198 297 199 298
rect 197 297 198 298
rect 196 297 197 298
rect 195 297 196 298
rect 194 297 195 298
rect 193 297 194 298
rect 180 297 181 298
rect 179 297 180 298
rect 178 297 179 298
rect 168 297 169 298
rect 167 297 168 298
rect 166 297 167 298
rect 151 297 152 298
rect 150 297 151 298
rect 149 297 150 298
rect 148 297 149 298
rect 147 297 148 298
rect 146 297 147 298
rect 145 297 146 298
rect 144 297 145 298
rect 143 297 144 298
rect 142 297 143 298
rect 141 297 142 298
rect 140 297 141 298
rect 139 297 140 298
rect 138 297 139 298
rect 137 297 138 298
rect 136 297 137 298
rect 135 297 136 298
rect 134 297 135 298
rect 133 297 134 298
rect 132 297 133 298
rect 131 297 132 298
rect 130 297 131 298
rect 129 297 130 298
rect 128 297 129 298
rect 127 297 128 298
rect 126 297 127 298
rect 125 297 126 298
rect 124 297 125 298
rect 123 297 124 298
rect 122 297 123 298
rect 121 297 122 298
rect 120 297 121 298
rect 119 297 120 298
rect 118 297 119 298
rect 117 297 118 298
rect 116 297 117 298
rect 115 297 116 298
rect 114 297 115 298
rect 113 297 114 298
rect 112 297 113 298
rect 111 297 112 298
rect 110 297 111 298
rect 109 297 110 298
rect 108 297 109 298
rect 107 297 108 298
rect 106 297 107 298
rect 105 297 106 298
rect 104 297 105 298
rect 31 297 32 298
rect 30 297 31 298
rect 29 297 30 298
rect 28 297 29 298
rect 21 297 22 298
rect 20 297 21 298
rect 19 297 20 298
rect 18 297 19 298
rect 17 297 18 298
rect 198 298 199 299
rect 197 298 198 299
rect 196 298 197 299
rect 195 298 196 299
rect 194 298 195 299
rect 179 298 180 299
rect 151 298 152 299
rect 150 298 151 299
rect 149 298 150 299
rect 148 298 149 299
rect 147 298 148 299
rect 146 298 147 299
rect 145 298 146 299
rect 144 298 145 299
rect 143 298 144 299
rect 142 298 143 299
rect 141 298 142 299
rect 140 298 141 299
rect 139 298 140 299
rect 138 298 139 299
rect 137 298 138 299
rect 136 298 137 299
rect 135 298 136 299
rect 134 298 135 299
rect 133 298 134 299
rect 132 298 133 299
rect 131 298 132 299
rect 130 298 131 299
rect 129 298 130 299
rect 128 298 129 299
rect 127 298 128 299
rect 126 298 127 299
rect 125 298 126 299
rect 124 298 125 299
rect 123 298 124 299
rect 122 298 123 299
rect 121 298 122 299
rect 120 298 121 299
rect 119 298 120 299
rect 118 298 119 299
rect 117 298 118 299
rect 116 298 117 299
rect 115 298 116 299
rect 114 298 115 299
rect 113 298 114 299
rect 112 298 113 299
rect 111 298 112 299
rect 110 298 111 299
rect 109 298 110 299
rect 108 298 109 299
rect 107 298 108 299
rect 106 298 107 299
rect 105 298 106 299
rect 104 298 105 299
rect 31 298 32 299
rect 30 298 31 299
rect 29 298 30 299
rect 19 298 20 299
rect 18 298 19 299
rect 17 298 18 299
rect 196 299 197 300
rect 151 299 152 300
rect 150 299 151 300
rect 149 299 150 300
rect 148 299 149 300
rect 147 299 148 300
rect 146 299 147 300
rect 145 299 146 300
rect 144 299 145 300
rect 143 299 144 300
rect 142 299 143 300
rect 141 299 142 300
rect 140 299 141 300
rect 139 299 140 300
rect 138 299 139 300
rect 137 299 138 300
rect 136 299 137 300
rect 135 299 136 300
rect 134 299 135 300
rect 133 299 134 300
rect 132 299 133 300
rect 131 299 132 300
rect 130 299 131 300
rect 129 299 130 300
rect 128 299 129 300
rect 127 299 128 300
rect 126 299 127 300
rect 125 299 126 300
rect 124 299 125 300
rect 123 299 124 300
rect 122 299 123 300
rect 121 299 122 300
rect 120 299 121 300
rect 119 299 120 300
rect 118 299 119 300
rect 117 299 118 300
rect 116 299 117 300
rect 115 299 116 300
rect 114 299 115 300
rect 113 299 114 300
rect 112 299 113 300
rect 111 299 112 300
rect 110 299 111 300
rect 109 299 110 300
rect 108 299 109 300
rect 107 299 108 300
rect 106 299 107 300
rect 105 299 106 300
rect 104 299 105 300
rect 31 299 32 300
rect 30 299 31 300
rect 29 299 30 300
rect 19 299 20 300
rect 18 299 19 300
rect 17 299 18 300
rect 16 299 17 300
rect 198 300 199 301
rect 197 300 198 301
rect 196 300 197 301
rect 195 300 196 301
rect 194 300 195 301
rect 193 300 194 301
rect 184 300 185 301
rect 183 300 184 301
rect 182 300 183 301
rect 181 300 182 301
rect 180 300 181 301
rect 179 300 180 301
rect 178 300 179 301
rect 177 300 178 301
rect 176 300 177 301
rect 175 300 176 301
rect 174 300 175 301
rect 173 300 174 301
rect 172 300 173 301
rect 171 300 172 301
rect 170 300 171 301
rect 169 300 170 301
rect 168 300 169 301
rect 167 300 168 301
rect 166 300 167 301
rect 165 300 166 301
rect 151 300 152 301
rect 150 300 151 301
rect 149 300 150 301
rect 148 300 149 301
rect 147 300 148 301
rect 146 300 147 301
rect 145 300 146 301
rect 144 300 145 301
rect 143 300 144 301
rect 142 300 143 301
rect 141 300 142 301
rect 140 300 141 301
rect 139 300 140 301
rect 138 300 139 301
rect 137 300 138 301
rect 136 300 137 301
rect 135 300 136 301
rect 134 300 135 301
rect 133 300 134 301
rect 132 300 133 301
rect 131 300 132 301
rect 130 300 131 301
rect 129 300 130 301
rect 128 300 129 301
rect 127 300 128 301
rect 126 300 127 301
rect 125 300 126 301
rect 124 300 125 301
rect 123 300 124 301
rect 122 300 123 301
rect 121 300 122 301
rect 120 300 121 301
rect 119 300 120 301
rect 118 300 119 301
rect 117 300 118 301
rect 116 300 117 301
rect 115 300 116 301
rect 114 300 115 301
rect 113 300 114 301
rect 112 300 113 301
rect 111 300 112 301
rect 110 300 111 301
rect 109 300 110 301
rect 108 300 109 301
rect 107 300 108 301
rect 106 300 107 301
rect 105 300 106 301
rect 104 300 105 301
rect 71 300 72 301
rect 70 300 71 301
rect 69 300 70 301
rect 31 300 32 301
rect 30 300 31 301
rect 29 300 30 301
rect 18 300 19 301
rect 17 300 18 301
rect 16 300 17 301
rect 199 301 200 302
rect 198 301 199 302
rect 197 301 198 302
rect 196 301 197 302
rect 195 301 196 302
rect 194 301 195 302
rect 193 301 194 302
rect 185 301 186 302
rect 184 301 185 302
rect 183 301 184 302
rect 182 301 183 302
rect 181 301 182 302
rect 180 301 181 302
rect 179 301 180 302
rect 178 301 179 302
rect 177 301 178 302
rect 176 301 177 302
rect 175 301 176 302
rect 174 301 175 302
rect 173 301 174 302
rect 172 301 173 302
rect 171 301 172 302
rect 170 301 171 302
rect 169 301 170 302
rect 168 301 169 302
rect 167 301 168 302
rect 166 301 167 302
rect 165 301 166 302
rect 164 301 165 302
rect 151 301 152 302
rect 150 301 151 302
rect 149 301 150 302
rect 148 301 149 302
rect 147 301 148 302
rect 146 301 147 302
rect 145 301 146 302
rect 144 301 145 302
rect 143 301 144 302
rect 142 301 143 302
rect 141 301 142 302
rect 140 301 141 302
rect 139 301 140 302
rect 138 301 139 302
rect 137 301 138 302
rect 136 301 137 302
rect 135 301 136 302
rect 134 301 135 302
rect 133 301 134 302
rect 132 301 133 302
rect 131 301 132 302
rect 130 301 131 302
rect 129 301 130 302
rect 128 301 129 302
rect 127 301 128 302
rect 126 301 127 302
rect 125 301 126 302
rect 124 301 125 302
rect 123 301 124 302
rect 122 301 123 302
rect 121 301 122 302
rect 120 301 121 302
rect 119 301 120 302
rect 118 301 119 302
rect 117 301 118 302
rect 116 301 117 302
rect 115 301 116 302
rect 114 301 115 302
rect 113 301 114 302
rect 112 301 113 302
rect 111 301 112 302
rect 110 301 111 302
rect 109 301 110 302
rect 108 301 109 302
rect 107 301 108 302
rect 106 301 107 302
rect 105 301 106 302
rect 104 301 105 302
rect 77 301 78 302
rect 76 301 77 302
rect 75 301 76 302
rect 74 301 75 302
rect 73 301 74 302
rect 72 301 73 302
rect 71 301 72 302
rect 70 301 71 302
rect 69 301 70 302
rect 68 301 69 302
rect 67 301 68 302
rect 66 301 67 302
rect 65 301 66 302
rect 64 301 65 302
rect 63 301 64 302
rect 31 301 32 302
rect 30 301 31 302
rect 29 301 30 302
rect 18 301 19 302
rect 17 301 18 302
rect 16 301 17 302
rect 194 302 195 303
rect 193 302 194 303
rect 185 302 186 303
rect 184 302 185 303
rect 183 302 184 303
rect 182 302 183 303
rect 181 302 182 303
rect 180 302 181 303
rect 179 302 180 303
rect 178 302 179 303
rect 177 302 178 303
rect 176 302 177 303
rect 175 302 176 303
rect 174 302 175 303
rect 173 302 174 303
rect 172 302 173 303
rect 171 302 172 303
rect 170 302 171 303
rect 169 302 170 303
rect 168 302 169 303
rect 167 302 168 303
rect 166 302 167 303
rect 165 302 166 303
rect 164 302 165 303
rect 151 302 152 303
rect 150 302 151 303
rect 149 302 150 303
rect 148 302 149 303
rect 147 302 148 303
rect 146 302 147 303
rect 145 302 146 303
rect 144 302 145 303
rect 143 302 144 303
rect 142 302 143 303
rect 141 302 142 303
rect 140 302 141 303
rect 139 302 140 303
rect 138 302 139 303
rect 137 302 138 303
rect 136 302 137 303
rect 135 302 136 303
rect 134 302 135 303
rect 133 302 134 303
rect 132 302 133 303
rect 131 302 132 303
rect 130 302 131 303
rect 129 302 130 303
rect 128 302 129 303
rect 127 302 128 303
rect 126 302 127 303
rect 125 302 126 303
rect 124 302 125 303
rect 123 302 124 303
rect 122 302 123 303
rect 121 302 122 303
rect 120 302 121 303
rect 119 302 120 303
rect 118 302 119 303
rect 117 302 118 303
rect 116 302 117 303
rect 115 302 116 303
rect 114 302 115 303
rect 113 302 114 303
rect 112 302 113 303
rect 111 302 112 303
rect 110 302 111 303
rect 109 302 110 303
rect 108 302 109 303
rect 107 302 108 303
rect 106 302 107 303
rect 105 302 106 303
rect 104 302 105 303
rect 80 302 81 303
rect 79 302 80 303
rect 78 302 79 303
rect 77 302 78 303
rect 76 302 77 303
rect 75 302 76 303
rect 74 302 75 303
rect 73 302 74 303
rect 72 302 73 303
rect 71 302 72 303
rect 70 302 71 303
rect 69 302 70 303
rect 68 302 69 303
rect 67 302 68 303
rect 66 302 67 303
rect 65 302 66 303
rect 64 302 65 303
rect 63 302 64 303
rect 62 302 63 303
rect 61 302 62 303
rect 60 302 61 303
rect 31 302 32 303
rect 30 302 31 303
rect 29 302 30 303
rect 28 302 29 303
rect 18 302 19 303
rect 17 302 18 303
rect 16 302 17 303
rect 194 303 195 304
rect 193 303 194 304
rect 185 303 186 304
rect 184 303 185 304
rect 183 303 184 304
rect 182 303 183 304
rect 181 303 182 304
rect 180 303 181 304
rect 179 303 180 304
rect 178 303 179 304
rect 177 303 178 304
rect 176 303 177 304
rect 175 303 176 304
rect 174 303 175 304
rect 173 303 174 304
rect 172 303 173 304
rect 171 303 172 304
rect 170 303 171 304
rect 169 303 170 304
rect 168 303 169 304
rect 167 303 168 304
rect 166 303 167 304
rect 165 303 166 304
rect 164 303 165 304
rect 151 303 152 304
rect 150 303 151 304
rect 149 303 150 304
rect 148 303 149 304
rect 147 303 148 304
rect 146 303 147 304
rect 145 303 146 304
rect 144 303 145 304
rect 143 303 144 304
rect 142 303 143 304
rect 141 303 142 304
rect 140 303 141 304
rect 139 303 140 304
rect 138 303 139 304
rect 137 303 138 304
rect 136 303 137 304
rect 135 303 136 304
rect 134 303 135 304
rect 133 303 134 304
rect 132 303 133 304
rect 131 303 132 304
rect 130 303 131 304
rect 129 303 130 304
rect 128 303 129 304
rect 127 303 128 304
rect 126 303 127 304
rect 125 303 126 304
rect 124 303 125 304
rect 123 303 124 304
rect 122 303 123 304
rect 121 303 122 304
rect 120 303 121 304
rect 119 303 120 304
rect 118 303 119 304
rect 117 303 118 304
rect 116 303 117 304
rect 115 303 116 304
rect 114 303 115 304
rect 113 303 114 304
rect 112 303 113 304
rect 111 303 112 304
rect 110 303 111 304
rect 109 303 110 304
rect 108 303 109 304
rect 107 303 108 304
rect 106 303 107 304
rect 105 303 106 304
rect 104 303 105 304
rect 83 303 84 304
rect 82 303 83 304
rect 81 303 82 304
rect 80 303 81 304
rect 79 303 80 304
rect 78 303 79 304
rect 77 303 78 304
rect 76 303 77 304
rect 75 303 76 304
rect 74 303 75 304
rect 73 303 74 304
rect 72 303 73 304
rect 71 303 72 304
rect 70 303 71 304
rect 69 303 70 304
rect 68 303 69 304
rect 67 303 68 304
rect 66 303 67 304
rect 65 303 66 304
rect 64 303 65 304
rect 63 303 64 304
rect 62 303 63 304
rect 61 303 62 304
rect 60 303 61 304
rect 59 303 60 304
rect 58 303 59 304
rect 30 303 31 304
rect 29 303 30 304
rect 28 303 29 304
rect 27 303 28 304
rect 19 303 20 304
rect 18 303 19 304
rect 17 303 18 304
rect 16 303 17 304
rect 199 304 200 305
rect 198 304 199 305
rect 197 304 198 305
rect 196 304 197 305
rect 195 304 196 305
rect 194 304 195 305
rect 193 304 194 305
rect 175 304 176 305
rect 174 304 175 305
rect 173 304 174 305
rect 172 304 173 305
rect 151 304 152 305
rect 150 304 151 305
rect 149 304 150 305
rect 148 304 149 305
rect 147 304 148 305
rect 146 304 147 305
rect 145 304 146 305
rect 144 304 145 305
rect 143 304 144 305
rect 142 304 143 305
rect 141 304 142 305
rect 140 304 141 305
rect 139 304 140 305
rect 138 304 139 305
rect 137 304 138 305
rect 136 304 137 305
rect 135 304 136 305
rect 134 304 135 305
rect 133 304 134 305
rect 132 304 133 305
rect 131 304 132 305
rect 130 304 131 305
rect 129 304 130 305
rect 128 304 129 305
rect 127 304 128 305
rect 126 304 127 305
rect 125 304 126 305
rect 124 304 125 305
rect 123 304 124 305
rect 122 304 123 305
rect 121 304 122 305
rect 120 304 121 305
rect 119 304 120 305
rect 118 304 119 305
rect 117 304 118 305
rect 116 304 117 305
rect 115 304 116 305
rect 114 304 115 305
rect 113 304 114 305
rect 112 304 113 305
rect 111 304 112 305
rect 110 304 111 305
rect 109 304 110 305
rect 108 304 109 305
rect 107 304 108 305
rect 106 304 107 305
rect 105 304 106 305
rect 104 304 105 305
rect 84 304 85 305
rect 83 304 84 305
rect 82 304 83 305
rect 81 304 82 305
rect 80 304 81 305
rect 79 304 80 305
rect 78 304 79 305
rect 77 304 78 305
rect 76 304 77 305
rect 75 304 76 305
rect 74 304 75 305
rect 73 304 74 305
rect 72 304 73 305
rect 71 304 72 305
rect 70 304 71 305
rect 69 304 70 305
rect 68 304 69 305
rect 67 304 68 305
rect 66 304 67 305
rect 65 304 66 305
rect 64 304 65 305
rect 63 304 64 305
rect 62 304 63 305
rect 61 304 62 305
rect 60 304 61 305
rect 59 304 60 305
rect 58 304 59 305
rect 57 304 58 305
rect 56 304 57 305
rect 29 304 30 305
rect 28 304 29 305
rect 27 304 28 305
rect 21 304 22 305
rect 20 304 21 305
rect 19 304 20 305
rect 18 304 19 305
rect 17 304 18 305
rect 198 305 199 306
rect 197 305 198 306
rect 196 305 197 306
rect 195 305 196 306
rect 194 305 195 306
rect 193 305 194 306
rect 175 305 176 306
rect 174 305 175 306
rect 173 305 174 306
rect 172 305 173 306
rect 151 305 152 306
rect 150 305 151 306
rect 149 305 150 306
rect 148 305 149 306
rect 147 305 148 306
rect 146 305 147 306
rect 145 305 146 306
rect 144 305 145 306
rect 143 305 144 306
rect 142 305 143 306
rect 141 305 142 306
rect 140 305 141 306
rect 139 305 140 306
rect 138 305 139 306
rect 137 305 138 306
rect 136 305 137 306
rect 135 305 136 306
rect 134 305 135 306
rect 133 305 134 306
rect 132 305 133 306
rect 131 305 132 306
rect 130 305 131 306
rect 129 305 130 306
rect 128 305 129 306
rect 127 305 128 306
rect 126 305 127 306
rect 125 305 126 306
rect 124 305 125 306
rect 123 305 124 306
rect 122 305 123 306
rect 121 305 122 306
rect 120 305 121 306
rect 119 305 120 306
rect 118 305 119 306
rect 117 305 118 306
rect 116 305 117 306
rect 115 305 116 306
rect 114 305 115 306
rect 113 305 114 306
rect 112 305 113 306
rect 111 305 112 306
rect 110 305 111 306
rect 109 305 110 306
rect 108 305 109 306
rect 107 305 108 306
rect 106 305 107 306
rect 105 305 106 306
rect 104 305 105 306
rect 86 305 87 306
rect 85 305 86 306
rect 84 305 85 306
rect 83 305 84 306
rect 82 305 83 306
rect 81 305 82 306
rect 80 305 81 306
rect 79 305 80 306
rect 78 305 79 306
rect 77 305 78 306
rect 76 305 77 306
rect 75 305 76 306
rect 74 305 75 306
rect 73 305 74 306
rect 72 305 73 306
rect 71 305 72 306
rect 70 305 71 306
rect 69 305 70 306
rect 68 305 69 306
rect 67 305 68 306
rect 66 305 67 306
rect 65 305 66 306
rect 64 305 65 306
rect 63 305 64 306
rect 62 305 63 306
rect 61 305 62 306
rect 60 305 61 306
rect 59 305 60 306
rect 58 305 59 306
rect 57 305 58 306
rect 56 305 57 306
rect 55 305 56 306
rect 28 305 29 306
rect 27 305 28 306
rect 21 305 22 306
rect 20 305 21 306
rect 19 305 20 306
rect 18 305 19 306
rect 194 306 195 307
rect 193 306 194 307
rect 175 306 176 307
rect 174 306 175 307
rect 173 306 174 307
rect 172 306 173 307
rect 151 306 152 307
rect 150 306 151 307
rect 149 306 150 307
rect 148 306 149 307
rect 147 306 148 307
rect 146 306 147 307
rect 145 306 146 307
rect 144 306 145 307
rect 143 306 144 307
rect 142 306 143 307
rect 141 306 142 307
rect 140 306 141 307
rect 139 306 140 307
rect 138 306 139 307
rect 137 306 138 307
rect 136 306 137 307
rect 135 306 136 307
rect 134 306 135 307
rect 133 306 134 307
rect 132 306 133 307
rect 131 306 132 307
rect 130 306 131 307
rect 129 306 130 307
rect 128 306 129 307
rect 127 306 128 307
rect 126 306 127 307
rect 125 306 126 307
rect 124 306 125 307
rect 123 306 124 307
rect 122 306 123 307
rect 121 306 122 307
rect 120 306 121 307
rect 119 306 120 307
rect 118 306 119 307
rect 117 306 118 307
rect 116 306 117 307
rect 115 306 116 307
rect 114 306 115 307
rect 113 306 114 307
rect 112 306 113 307
rect 111 306 112 307
rect 110 306 111 307
rect 109 306 110 307
rect 108 306 109 307
rect 107 306 108 307
rect 106 306 107 307
rect 105 306 106 307
rect 104 306 105 307
rect 87 306 88 307
rect 86 306 87 307
rect 85 306 86 307
rect 84 306 85 307
rect 83 306 84 307
rect 82 306 83 307
rect 81 306 82 307
rect 80 306 81 307
rect 79 306 80 307
rect 78 306 79 307
rect 77 306 78 307
rect 63 306 64 307
rect 62 306 63 307
rect 61 306 62 307
rect 60 306 61 307
rect 59 306 60 307
rect 58 306 59 307
rect 57 306 58 307
rect 56 306 57 307
rect 55 306 56 307
rect 54 306 55 307
rect 53 306 54 307
rect 20 306 21 307
rect 19 306 20 307
rect 198 307 199 308
rect 197 307 198 308
rect 196 307 197 308
rect 195 307 196 308
rect 194 307 195 308
rect 193 307 194 308
rect 174 307 175 308
rect 173 307 174 308
rect 151 307 152 308
rect 150 307 151 308
rect 149 307 150 308
rect 148 307 149 308
rect 147 307 148 308
rect 146 307 147 308
rect 145 307 146 308
rect 144 307 145 308
rect 143 307 144 308
rect 142 307 143 308
rect 141 307 142 308
rect 140 307 141 308
rect 139 307 140 308
rect 138 307 139 308
rect 137 307 138 308
rect 136 307 137 308
rect 135 307 136 308
rect 134 307 135 308
rect 133 307 134 308
rect 132 307 133 308
rect 131 307 132 308
rect 130 307 131 308
rect 129 307 130 308
rect 128 307 129 308
rect 127 307 128 308
rect 126 307 127 308
rect 125 307 126 308
rect 124 307 125 308
rect 123 307 124 308
rect 122 307 123 308
rect 121 307 122 308
rect 120 307 121 308
rect 119 307 120 308
rect 118 307 119 308
rect 117 307 118 308
rect 116 307 117 308
rect 115 307 116 308
rect 114 307 115 308
rect 113 307 114 308
rect 112 307 113 308
rect 111 307 112 308
rect 110 307 111 308
rect 109 307 110 308
rect 108 307 109 308
rect 107 307 108 308
rect 106 307 107 308
rect 105 307 106 308
rect 104 307 105 308
rect 88 307 89 308
rect 87 307 88 308
rect 86 307 87 308
rect 85 307 86 308
rect 84 307 85 308
rect 83 307 84 308
rect 82 307 83 308
rect 59 307 60 308
rect 58 307 59 308
rect 57 307 58 308
rect 56 307 57 308
rect 55 307 56 308
rect 54 307 55 308
rect 53 307 54 308
rect 199 308 200 309
rect 198 308 199 309
rect 197 308 198 309
rect 196 308 197 309
rect 195 308 196 309
rect 194 308 195 309
rect 193 308 194 309
rect 151 308 152 309
rect 150 308 151 309
rect 149 308 150 309
rect 148 308 149 309
rect 147 308 148 309
rect 146 308 147 309
rect 145 308 146 309
rect 144 308 145 309
rect 143 308 144 309
rect 142 308 143 309
rect 141 308 142 309
rect 140 308 141 309
rect 139 308 140 309
rect 138 308 139 309
rect 137 308 138 309
rect 136 308 137 309
rect 135 308 136 309
rect 134 308 135 309
rect 133 308 134 309
rect 132 308 133 309
rect 131 308 132 309
rect 130 308 131 309
rect 129 308 130 309
rect 128 308 129 309
rect 127 308 128 309
rect 126 308 127 309
rect 125 308 126 309
rect 124 308 125 309
rect 123 308 124 309
rect 122 308 123 309
rect 121 308 122 309
rect 120 308 121 309
rect 119 308 120 309
rect 118 308 119 309
rect 117 308 118 309
rect 116 308 117 309
rect 115 308 116 309
rect 114 308 115 309
rect 113 308 114 309
rect 112 308 113 309
rect 111 308 112 309
rect 110 308 111 309
rect 109 308 110 309
rect 108 308 109 309
rect 107 308 108 309
rect 106 308 107 309
rect 105 308 106 309
rect 104 308 105 309
rect 88 308 89 309
rect 87 308 88 309
rect 86 308 87 309
rect 85 308 86 309
rect 84 308 85 309
rect 57 308 58 309
rect 56 308 57 309
rect 55 308 56 309
rect 54 308 55 309
rect 53 308 54 309
rect 31 308 32 309
rect 30 308 31 309
rect 29 308 30 309
rect 28 308 29 309
rect 27 308 28 309
rect 198 309 199 310
rect 197 309 198 310
rect 196 309 197 310
rect 195 309 196 310
rect 194 309 195 310
rect 151 309 152 310
rect 150 309 151 310
rect 149 309 150 310
rect 148 309 149 310
rect 147 309 148 310
rect 146 309 147 310
rect 145 309 146 310
rect 144 309 145 310
rect 143 309 144 310
rect 142 309 143 310
rect 141 309 142 310
rect 140 309 141 310
rect 139 309 140 310
rect 138 309 139 310
rect 137 309 138 310
rect 136 309 137 310
rect 135 309 136 310
rect 134 309 135 310
rect 133 309 134 310
rect 132 309 133 310
rect 131 309 132 310
rect 130 309 131 310
rect 129 309 130 310
rect 128 309 129 310
rect 127 309 128 310
rect 126 309 127 310
rect 125 309 126 310
rect 124 309 125 310
rect 123 309 124 310
rect 122 309 123 310
rect 121 309 122 310
rect 120 309 121 310
rect 119 309 120 310
rect 118 309 119 310
rect 117 309 118 310
rect 116 309 117 310
rect 115 309 116 310
rect 114 309 115 310
rect 113 309 114 310
rect 112 309 113 310
rect 111 309 112 310
rect 110 309 111 310
rect 109 309 110 310
rect 108 309 109 310
rect 107 309 108 310
rect 106 309 107 310
rect 105 309 106 310
rect 104 309 105 310
rect 88 309 89 310
rect 87 309 88 310
rect 54 309 55 310
rect 53 309 54 310
rect 31 309 32 310
rect 30 309 31 310
rect 29 309 30 310
rect 28 309 29 310
rect 27 309 28 310
rect 26 309 27 310
rect 25 309 26 310
rect 24 309 25 310
rect 23 309 24 310
rect 22 309 23 310
rect 198 310 199 311
rect 194 310 195 311
rect 151 310 152 311
rect 150 310 151 311
rect 149 310 150 311
rect 148 310 149 311
rect 147 310 148 311
rect 146 310 147 311
rect 145 310 146 311
rect 144 310 145 311
rect 143 310 144 311
rect 142 310 143 311
rect 141 310 142 311
rect 140 310 141 311
rect 139 310 140 311
rect 138 310 139 311
rect 137 310 138 311
rect 136 310 137 311
rect 135 310 136 311
rect 134 310 135 311
rect 133 310 134 311
rect 132 310 133 311
rect 131 310 132 311
rect 130 310 131 311
rect 129 310 130 311
rect 128 310 129 311
rect 127 310 128 311
rect 126 310 127 311
rect 125 310 126 311
rect 124 310 125 311
rect 123 310 124 311
rect 122 310 123 311
rect 121 310 122 311
rect 120 310 121 311
rect 119 310 120 311
rect 118 310 119 311
rect 117 310 118 311
rect 116 310 117 311
rect 115 310 116 311
rect 114 310 115 311
rect 113 310 114 311
rect 112 310 113 311
rect 111 310 112 311
rect 110 310 111 311
rect 109 310 110 311
rect 108 310 109 311
rect 107 310 108 311
rect 106 310 107 311
rect 105 310 106 311
rect 104 310 105 311
rect 31 310 32 311
rect 30 310 31 311
rect 29 310 30 311
rect 28 310 29 311
rect 27 310 28 311
rect 26 310 27 311
rect 25 310 26 311
rect 24 310 25 311
rect 23 310 24 311
rect 22 310 23 311
rect 21 310 22 311
rect 20 310 21 311
rect 19 310 20 311
rect 18 310 19 311
rect 17 310 18 311
rect 199 311 200 312
rect 198 311 199 312
rect 197 311 198 312
rect 196 311 197 312
rect 195 311 196 312
rect 194 311 195 312
rect 193 311 194 312
rect 151 311 152 312
rect 150 311 151 312
rect 149 311 150 312
rect 148 311 149 312
rect 147 311 148 312
rect 146 311 147 312
rect 145 311 146 312
rect 144 311 145 312
rect 143 311 144 312
rect 142 311 143 312
rect 141 311 142 312
rect 140 311 141 312
rect 139 311 140 312
rect 138 311 139 312
rect 137 311 138 312
rect 136 311 137 312
rect 135 311 136 312
rect 134 311 135 312
rect 133 311 134 312
rect 132 311 133 312
rect 131 311 132 312
rect 130 311 131 312
rect 129 311 130 312
rect 128 311 129 312
rect 127 311 128 312
rect 126 311 127 312
rect 125 311 126 312
rect 124 311 125 312
rect 123 311 124 312
rect 122 311 123 312
rect 121 311 122 312
rect 120 311 121 312
rect 119 311 120 312
rect 118 311 119 312
rect 117 311 118 312
rect 116 311 117 312
rect 115 311 116 312
rect 114 311 115 312
rect 113 311 114 312
rect 112 311 113 312
rect 111 311 112 312
rect 110 311 111 312
rect 109 311 110 312
rect 108 311 109 312
rect 107 311 108 312
rect 106 311 107 312
rect 105 311 106 312
rect 104 311 105 312
rect 27 311 28 312
rect 26 311 27 312
rect 25 311 26 312
rect 24 311 25 312
rect 23 311 24 312
rect 22 311 23 312
rect 21 311 22 312
rect 20 311 21 312
rect 19 311 20 312
rect 18 311 19 312
rect 17 311 18 312
rect 16 311 17 312
rect 198 312 199 313
rect 197 312 198 313
rect 196 312 197 313
rect 195 312 196 313
rect 194 312 195 313
rect 193 312 194 313
rect 151 312 152 313
rect 150 312 151 313
rect 149 312 150 313
rect 148 312 149 313
rect 147 312 148 313
rect 146 312 147 313
rect 145 312 146 313
rect 144 312 145 313
rect 143 312 144 313
rect 142 312 143 313
rect 141 312 142 313
rect 140 312 141 313
rect 139 312 140 313
rect 138 312 139 313
rect 137 312 138 313
rect 136 312 137 313
rect 135 312 136 313
rect 134 312 135 313
rect 133 312 134 313
rect 132 312 133 313
rect 131 312 132 313
rect 130 312 131 313
rect 129 312 130 313
rect 128 312 129 313
rect 127 312 128 313
rect 126 312 127 313
rect 125 312 126 313
rect 124 312 125 313
rect 123 312 124 313
rect 122 312 123 313
rect 121 312 122 313
rect 120 312 121 313
rect 119 312 120 313
rect 118 312 119 313
rect 117 312 118 313
rect 116 312 117 313
rect 115 312 116 313
rect 114 312 115 313
rect 113 312 114 313
rect 112 312 113 313
rect 111 312 112 313
rect 110 312 111 313
rect 109 312 110 313
rect 108 312 109 313
rect 107 312 108 313
rect 106 312 107 313
rect 105 312 106 313
rect 104 312 105 313
rect 23 312 24 313
rect 22 312 23 313
rect 21 312 22 313
rect 20 312 21 313
rect 19 312 20 313
rect 18 312 19 313
rect 17 312 18 313
rect 16 312 17 313
rect 194 313 195 314
rect 193 313 194 314
rect 151 313 152 314
rect 150 313 151 314
rect 149 313 150 314
rect 148 313 149 314
rect 147 313 148 314
rect 146 313 147 314
rect 145 313 146 314
rect 144 313 145 314
rect 143 313 144 314
rect 142 313 143 314
rect 141 313 142 314
rect 140 313 141 314
rect 139 313 140 314
rect 138 313 139 314
rect 137 313 138 314
rect 136 313 137 314
rect 135 313 136 314
rect 134 313 135 314
rect 133 313 134 314
rect 132 313 133 314
rect 131 313 132 314
rect 130 313 131 314
rect 129 313 130 314
rect 128 313 129 314
rect 127 313 128 314
rect 126 313 127 314
rect 125 313 126 314
rect 124 313 125 314
rect 123 313 124 314
rect 122 313 123 314
rect 121 313 122 314
rect 120 313 121 314
rect 119 313 120 314
rect 118 313 119 314
rect 117 313 118 314
rect 116 313 117 314
rect 115 313 116 314
rect 114 313 115 314
rect 113 313 114 314
rect 112 313 113 314
rect 111 313 112 314
rect 110 313 111 314
rect 109 313 110 314
rect 108 313 109 314
rect 107 313 108 314
rect 106 313 107 314
rect 105 313 106 314
rect 104 313 105 314
rect 22 313 23 314
rect 21 313 22 314
rect 18 313 19 314
rect 17 313 18 314
rect 198 314 199 315
rect 197 314 198 315
rect 196 314 197 315
rect 195 314 196 315
rect 194 314 195 315
rect 193 314 194 315
rect 151 314 152 315
rect 150 314 151 315
rect 149 314 150 315
rect 148 314 149 315
rect 147 314 148 315
rect 146 314 147 315
rect 145 314 146 315
rect 144 314 145 315
rect 143 314 144 315
rect 142 314 143 315
rect 141 314 142 315
rect 140 314 141 315
rect 139 314 140 315
rect 138 314 139 315
rect 137 314 138 315
rect 136 314 137 315
rect 135 314 136 315
rect 134 314 135 315
rect 133 314 134 315
rect 132 314 133 315
rect 131 314 132 315
rect 130 314 131 315
rect 129 314 130 315
rect 128 314 129 315
rect 127 314 128 315
rect 126 314 127 315
rect 125 314 126 315
rect 124 314 125 315
rect 123 314 124 315
rect 122 314 123 315
rect 121 314 122 315
rect 120 314 121 315
rect 119 314 120 315
rect 118 314 119 315
rect 117 314 118 315
rect 116 314 117 315
rect 115 314 116 315
rect 114 314 115 315
rect 113 314 114 315
rect 112 314 113 315
rect 111 314 112 315
rect 110 314 111 315
rect 109 314 110 315
rect 108 314 109 315
rect 107 314 108 315
rect 106 314 107 315
rect 105 314 106 315
rect 104 314 105 315
rect 80 314 81 315
rect 79 314 80 315
rect 78 314 79 315
rect 77 314 78 315
rect 76 314 77 315
rect 75 314 76 315
rect 74 314 75 315
rect 73 314 74 315
rect 72 314 73 315
rect 71 314 72 315
rect 70 314 71 315
rect 69 314 70 315
rect 68 314 69 315
rect 67 314 68 315
rect 66 314 67 315
rect 65 314 66 315
rect 64 314 65 315
rect 63 314 64 315
rect 62 314 63 315
rect 61 314 62 315
rect 60 314 61 315
rect 59 314 60 315
rect 58 314 59 315
rect 57 314 58 315
rect 56 314 57 315
rect 55 314 56 315
rect 54 314 55 315
rect 53 314 54 315
rect 22 314 23 315
rect 21 314 22 315
rect 199 315 200 316
rect 198 315 199 316
rect 197 315 198 316
rect 196 315 197 316
rect 195 315 196 316
rect 194 315 195 316
rect 193 315 194 316
rect 151 315 152 316
rect 150 315 151 316
rect 149 315 150 316
rect 148 315 149 316
rect 147 315 148 316
rect 146 315 147 316
rect 145 315 146 316
rect 144 315 145 316
rect 143 315 144 316
rect 142 315 143 316
rect 141 315 142 316
rect 140 315 141 316
rect 139 315 140 316
rect 138 315 139 316
rect 137 315 138 316
rect 136 315 137 316
rect 135 315 136 316
rect 134 315 135 316
rect 133 315 134 316
rect 132 315 133 316
rect 131 315 132 316
rect 130 315 131 316
rect 129 315 130 316
rect 128 315 129 316
rect 127 315 128 316
rect 126 315 127 316
rect 125 315 126 316
rect 124 315 125 316
rect 123 315 124 316
rect 122 315 123 316
rect 121 315 122 316
rect 120 315 121 316
rect 119 315 120 316
rect 118 315 119 316
rect 117 315 118 316
rect 116 315 117 316
rect 115 315 116 316
rect 114 315 115 316
rect 113 315 114 316
rect 112 315 113 316
rect 111 315 112 316
rect 110 315 111 316
rect 109 315 110 316
rect 108 315 109 316
rect 107 315 108 316
rect 106 315 107 316
rect 105 315 106 316
rect 104 315 105 316
rect 80 315 81 316
rect 79 315 80 316
rect 78 315 79 316
rect 77 315 78 316
rect 76 315 77 316
rect 75 315 76 316
rect 74 315 75 316
rect 73 315 74 316
rect 72 315 73 316
rect 71 315 72 316
rect 70 315 71 316
rect 69 315 70 316
rect 68 315 69 316
rect 67 315 68 316
rect 66 315 67 316
rect 65 315 66 316
rect 64 315 65 316
rect 63 315 64 316
rect 62 315 63 316
rect 61 315 62 316
rect 60 315 61 316
rect 59 315 60 316
rect 58 315 59 316
rect 57 315 58 316
rect 56 315 57 316
rect 55 315 56 316
rect 54 315 55 316
rect 53 315 54 316
rect 31 315 32 316
rect 30 315 31 316
rect 29 315 30 316
rect 28 315 29 316
rect 27 315 28 316
rect 22 315 23 316
rect 21 315 22 316
rect 20 315 21 316
rect 194 316 195 317
rect 193 316 194 317
rect 176 316 177 317
rect 151 316 152 317
rect 150 316 151 317
rect 149 316 150 317
rect 148 316 149 317
rect 147 316 148 317
rect 146 316 147 317
rect 145 316 146 317
rect 144 316 145 317
rect 143 316 144 317
rect 142 316 143 317
rect 141 316 142 317
rect 140 316 141 317
rect 139 316 140 317
rect 138 316 139 317
rect 137 316 138 317
rect 136 316 137 317
rect 135 316 136 317
rect 134 316 135 317
rect 133 316 134 317
rect 132 316 133 317
rect 131 316 132 317
rect 130 316 131 317
rect 129 316 130 317
rect 128 316 129 317
rect 127 316 128 317
rect 126 316 127 317
rect 125 316 126 317
rect 124 316 125 317
rect 123 316 124 317
rect 122 316 123 317
rect 121 316 122 317
rect 120 316 121 317
rect 119 316 120 317
rect 118 316 119 317
rect 117 316 118 317
rect 116 316 117 317
rect 115 316 116 317
rect 114 316 115 317
rect 113 316 114 317
rect 112 316 113 317
rect 111 316 112 317
rect 110 316 111 317
rect 109 316 110 317
rect 108 316 109 317
rect 107 316 108 317
rect 106 316 107 317
rect 105 316 106 317
rect 104 316 105 317
rect 80 316 81 317
rect 79 316 80 317
rect 78 316 79 317
rect 77 316 78 317
rect 76 316 77 317
rect 75 316 76 317
rect 74 316 75 317
rect 73 316 74 317
rect 72 316 73 317
rect 71 316 72 317
rect 70 316 71 317
rect 69 316 70 317
rect 68 316 69 317
rect 67 316 68 317
rect 66 316 67 317
rect 65 316 66 317
rect 64 316 65 317
rect 63 316 64 317
rect 62 316 63 317
rect 61 316 62 317
rect 60 316 61 317
rect 59 316 60 317
rect 58 316 59 317
rect 57 316 58 317
rect 56 316 57 317
rect 55 316 56 317
rect 54 316 55 317
rect 53 316 54 317
rect 31 316 32 317
rect 30 316 31 317
rect 29 316 30 317
rect 28 316 29 317
rect 27 316 28 317
rect 26 316 27 317
rect 25 316 26 317
rect 24 316 25 317
rect 23 316 24 317
rect 22 316 23 317
rect 21 316 22 317
rect 20 316 21 317
rect 194 317 195 318
rect 193 317 194 318
rect 177 317 178 318
rect 176 317 177 318
rect 175 317 176 318
rect 151 317 152 318
rect 150 317 151 318
rect 149 317 150 318
rect 148 317 149 318
rect 147 317 148 318
rect 146 317 147 318
rect 145 317 146 318
rect 144 317 145 318
rect 143 317 144 318
rect 142 317 143 318
rect 141 317 142 318
rect 140 317 141 318
rect 139 317 140 318
rect 138 317 139 318
rect 137 317 138 318
rect 136 317 137 318
rect 135 317 136 318
rect 134 317 135 318
rect 133 317 134 318
rect 132 317 133 318
rect 131 317 132 318
rect 130 317 131 318
rect 129 317 130 318
rect 128 317 129 318
rect 127 317 128 318
rect 126 317 127 318
rect 125 317 126 318
rect 124 317 125 318
rect 123 317 124 318
rect 122 317 123 318
rect 121 317 122 318
rect 120 317 121 318
rect 119 317 120 318
rect 118 317 119 318
rect 117 317 118 318
rect 116 317 117 318
rect 115 317 116 318
rect 114 317 115 318
rect 113 317 114 318
rect 112 317 113 318
rect 111 317 112 318
rect 110 317 111 318
rect 109 317 110 318
rect 108 317 109 318
rect 107 317 108 318
rect 106 317 107 318
rect 105 317 106 318
rect 104 317 105 318
rect 80 317 81 318
rect 79 317 80 318
rect 78 317 79 318
rect 77 317 78 318
rect 76 317 77 318
rect 75 317 76 318
rect 74 317 75 318
rect 73 317 74 318
rect 72 317 73 318
rect 71 317 72 318
rect 70 317 71 318
rect 69 317 70 318
rect 68 317 69 318
rect 67 317 68 318
rect 66 317 67 318
rect 65 317 66 318
rect 64 317 65 318
rect 63 317 64 318
rect 62 317 63 318
rect 61 317 62 318
rect 60 317 61 318
rect 59 317 60 318
rect 58 317 59 318
rect 57 317 58 318
rect 56 317 57 318
rect 55 317 56 318
rect 54 317 55 318
rect 53 317 54 318
rect 31 317 32 318
rect 30 317 31 318
rect 29 317 30 318
rect 28 317 29 318
rect 27 317 28 318
rect 26 317 27 318
rect 25 317 26 318
rect 24 317 25 318
rect 23 317 24 318
rect 22 317 23 318
rect 21 317 22 318
rect 20 317 21 318
rect 198 318 199 319
rect 197 318 198 319
rect 196 318 197 319
rect 195 318 196 319
rect 194 318 195 319
rect 193 318 194 319
rect 177 318 178 319
rect 176 318 177 319
rect 175 318 176 319
rect 114 318 115 319
rect 113 318 114 319
rect 112 318 113 319
rect 111 318 112 319
rect 110 318 111 319
rect 109 318 110 319
rect 108 318 109 319
rect 107 318 108 319
rect 106 318 107 319
rect 105 318 106 319
rect 104 318 105 319
rect 80 318 81 319
rect 79 318 80 319
rect 78 318 79 319
rect 77 318 78 319
rect 76 318 77 319
rect 75 318 76 319
rect 74 318 75 319
rect 73 318 74 319
rect 72 318 73 319
rect 71 318 72 319
rect 70 318 71 319
rect 69 318 70 319
rect 68 318 69 319
rect 67 318 68 319
rect 66 318 67 319
rect 65 318 66 319
rect 64 318 65 319
rect 63 318 64 319
rect 62 318 63 319
rect 61 318 62 319
rect 60 318 61 319
rect 59 318 60 319
rect 58 318 59 319
rect 57 318 58 319
rect 56 318 57 319
rect 55 318 56 319
rect 54 318 55 319
rect 53 318 54 319
rect 28 318 29 319
rect 27 318 28 319
rect 26 318 27 319
rect 25 318 26 319
rect 24 318 25 319
rect 23 318 24 319
rect 22 318 23 319
rect 21 318 22 319
rect 198 319 199 320
rect 197 319 198 320
rect 196 319 197 320
rect 195 319 196 320
rect 194 319 195 320
rect 183 319 184 320
rect 182 319 183 320
rect 181 319 182 320
rect 177 319 178 320
rect 176 319 177 320
rect 175 319 176 320
rect 114 319 115 320
rect 113 319 114 320
rect 112 319 113 320
rect 111 319 112 320
rect 110 319 111 320
rect 109 319 110 320
rect 108 319 109 320
rect 107 319 108 320
rect 106 319 107 320
rect 105 319 106 320
rect 104 319 105 320
rect 80 319 81 320
rect 79 319 80 320
rect 78 319 79 320
rect 77 319 78 320
rect 76 319 77 320
rect 75 319 76 320
rect 74 319 75 320
rect 73 319 74 320
rect 72 319 73 320
rect 71 319 72 320
rect 70 319 71 320
rect 69 319 70 320
rect 68 319 69 320
rect 67 319 68 320
rect 66 319 67 320
rect 65 319 66 320
rect 64 319 65 320
rect 63 319 64 320
rect 62 319 63 320
rect 61 319 62 320
rect 60 319 61 320
rect 59 319 60 320
rect 58 319 59 320
rect 57 319 58 320
rect 56 319 57 320
rect 55 319 56 320
rect 54 319 55 320
rect 53 319 54 320
rect 23 319 24 320
rect 184 320 185 321
rect 183 320 184 321
rect 182 320 183 321
rect 181 320 182 321
rect 180 320 181 321
rect 177 320 178 321
rect 176 320 177 321
rect 175 320 176 321
rect 173 320 174 321
rect 172 320 173 321
rect 171 320 172 321
rect 170 320 171 321
rect 169 320 170 321
rect 168 320 169 321
rect 167 320 168 321
rect 166 320 167 321
rect 165 320 166 321
rect 164 320 165 321
rect 114 320 115 321
rect 113 320 114 321
rect 112 320 113 321
rect 111 320 112 321
rect 110 320 111 321
rect 109 320 110 321
rect 108 320 109 321
rect 107 320 108 321
rect 106 320 107 321
rect 105 320 106 321
rect 104 320 105 321
rect 68 320 69 321
rect 67 320 68 321
rect 66 320 67 321
rect 65 320 66 321
rect 64 320 65 321
rect 57 320 58 321
rect 56 320 57 321
rect 55 320 56 321
rect 54 320 55 321
rect 53 320 54 321
rect 198 321 199 322
rect 197 321 198 322
rect 196 321 197 322
rect 195 321 196 322
rect 194 321 195 322
rect 193 321 194 322
rect 184 321 185 322
rect 183 321 184 322
rect 182 321 183 322
rect 181 321 182 322
rect 180 321 181 322
rect 179 321 180 322
rect 177 321 178 322
rect 176 321 177 322
rect 175 321 176 322
rect 173 321 174 322
rect 172 321 173 322
rect 171 321 172 322
rect 170 321 171 322
rect 169 321 170 322
rect 168 321 169 322
rect 167 321 168 322
rect 166 321 167 322
rect 165 321 166 322
rect 164 321 165 322
rect 114 321 115 322
rect 113 321 114 322
rect 112 321 113 322
rect 111 321 112 322
rect 110 321 111 322
rect 109 321 110 322
rect 108 321 109 322
rect 107 321 108 322
rect 106 321 107 322
rect 105 321 106 322
rect 104 321 105 322
rect 68 321 69 322
rect 67 321 68 322
rect 66 321 67 322
rect 65 321 66 322
rect 64 321 65 322
rect 57 321 58 322
rect 56 321 57 322
rect 55 321 56 322
rect 54 321 55 322
rect 53 321 54 322
rect 31 321 32 322
rect 30 321 31 322
rect 29 321 30 322
rect 28 321 29 322
rect 27 321 28 322
rect 199 322 200 323
rect 198 322 199 323
rect 197 322 198 323
rect 196 322 197 323
rect 195 322 196 323
rect 194 322 195 323
rect 193 322 194 323
rect 185 322 186 323
rect 184 322 185 323
rect 183 322 184 323
rect 182 322 183 323
rect 181 322 182 323
rect 180 322 181 323
rect 179 322 180 323
rect 177 322 178 323
rect 176 322 177 323
rect 175 322 176 323
rect 173 322 174 323
rect 172 322 173 323
rect 171 322 172 323
rect 170 322 171 323
rect 169 322 170 323
rect 168 322 169 323
rect 167 322 168 323
rect 166 322 167 323
rect 165 322 166 323
rect 164 322 165 323
rect 114 322 115 323
rect 113 322 114 323
rect 112 322 113 323
rect 111 322 112 323
rect 110 322 111 323
rect 109 322 110 323
rect 108 322 109 323
rect 107 322 108 323
rect 106 322 107 323
rect 105 322 106 323
rect 104 322 105 323
rect 68 322 69 323
rect 67 322 68 323
rect 66 322 67 323
rect 65 322 66 323
rect 64 322 65 323
rect 57 322 58 323
rect 56 322 57 323
rect 55 322 56 323
rect 54 322 55 323
rect 53 322 54 323
rect 31 322 32 323
rect 30 322 31 323
rect 29 322 30 323
rect 28 322 29 323
rect 27 322 28 323
rect 26 322 27 323
rect 25 322 26 323
rect 24 322 25 323
rect 23 322 24 323
rect 22 322 23 323
rect 198 323 199 324
rect 185 323 186 324
rect 184 323 185 324
rect 183 323 184 324
rect 182 323 183 324
rect 181 323 182 324
rect 180 323 181 324
rect 179 323 180 324
rect 177 323 178 324
rect 176 323 177 324
rect 175 323 176 324
rect 173 323 174 324
rect 172 323 173 324
rect 171 323 172 324
rect 170 323 171 324
rect 169 323 170 324
rect 168 323 169 324
rect 167 323 168 324
rect 166 323 167 324
rect 165 323 166 324
rect 164 323 165 324
rect 114 323 115 324
rect 113 323 114 324
rect 112 323 113 324
rect 111 323 112 324
rect 110 323 111 324
rect 109 323 110 324
rect 108 323 109 324
rect 107 323 108 324
rect 106 323 107 324
rect 105 323 106 324
rect 104 323 105 324
rect 68 323 69 324
rect 67 323 68 324
rect 66 323 67 324
rect 65 323 66 324
rect 64 323 65 324
rect 57 323 58 324
rect 56 323 57 324
rect 55 323 56 324
rect 54 323 55 324
rect 53 323 54 324
rect 31 323 32 324
rect 30 323 31 324
rect 29 323 30 324
rect 28 323 29 324
rect 27 323 28 324
rect 26 323 27 324
rect 25 323 26 324
rect 24 323 25 324
rect 23 323 24 324
rect 22 323 23 324
rect 21 323 22 324
rect 18 323 19 324
rect 17 323 18 324
rect 198 324 199 325
rect 185 324 186 325
rect 184 324 185 325
rect 183 324 184 325
rect 181 324 182 325
rect 180 324 181 325
rect 179 324 180 325
rect 177 324 178 325
rect 176 324 177 325
rect 175 324 176 325
rect 173 324 174 325
rect 172 324 173 325
rect 171 324 172 325
rect 169 324 170 325
rect 168 324 169 325
rect 166 324 167 325
rect 165 324 166 325
rect 164 324 165 325
rect 114 324 115 325
rect 113 324 114 325
rect 112 324 113 325
rect 111 324 112 325
rect 110 324 111 325
rect 109 324 110 325
rect 108 324 109 325
rect 107 324 108 325
rect 106 324 107 325
rect 105 324 106 325
rect 104 324 105 325
rect 68 324 69 325
rect 67 324 68 325
rect 66 324 67 325
rect 65 324 66 325
rect 64 324 65 325
rect 57 324 58 325
rect 56 324 57 325
rect 55 324 56 325
rect 54 324 55 325
rect 53 324 54 325
rect 27 324 28 325
rect 26 324 27 325
rect 25 324 26 325
rect 24 324 25 325
rect 23 324 24 325
rect 22 324 23 325
rect 21 324 22 325
rect 20 324 21 325
rect 18 324 19 325
rect 17 324 18 325
rect 16 324 17 325
rect 199 325 200 326
rect 198 325 199 326
rect 197 325 198 326
rect 196 325 197 326
rect 195 325 196 326
rect 194 325 195 326
rect 193 325 194 326
rect 185 325 186 326
rect 184 325 185 326
rect 180 325 181 326
rect 179 325 180 326
rect 177 325 178 326
rect 176 325 177 326
rect 175 325 176 326
rect 173 325 174 326
rect 172 325 173 326
rect 171 325 172 326
rect 169 325 170 326
rect 168 325 169 326
rect 166 325 167 326
rect 165 325 166 326
rect 164 325 165 326
rect 114 325 115 326
rect 113 325 114 326
rect 112 325 113 326
rect 111 325 112 326
rect 110 325 111 326
rect 109 325 110 326
rect 108 325 109 326
rect 107 325 108 326
rect 106 325 107 326
rect 105 325 106 326
rect 104 325 105 326
rect 68 325 69 326
rect 67 325 68 326
rect 66 325 67 326
rect 65 325 66 326
rect 64 325 65 326
rect 57 325 58 326
rect 56 325 57 326
rect 55 325 56 326
rect 54 325 55 326
rect 53 325 54 326
rect 23 325 24 326
rect 22 325 23 326
rect 21 325 22 326
rect 18 325 19 326
rect 17 325 18 326
rect 16 325 17 326
rect 198 326 199 327
rect 197 326 198 327
rect 196 326 197 327
rect 195 326 196 327
rect 194 326 195 327
rect 193 326 194 327
rect 186 326 187 327
rect 185 326 186 327
rect 184 326 185 327
rect 180 326 181 327
rect 179 326 180 327
rect 178 326 179 327
rect 177 326 178 327
rect 176 326 177 327
rect 175 326 176 327
rect 173 326 174 327
rect 172 326 173 327
rect 171 326 172 327
rect 169 326 170 327
rect 168 326 169 327
rect 166 326 167 327
rect 165 326 166 327
rect 164 326 165 327
rect 114 326 115 327
rect 113 326 114 327
rect 112 326 113 327
rect 111 326 112 327
rect 110 326 111 327
rect 109 326 110 327
rect 108 326 109 327
rect 107 326 108 327
rect 106 326 107 327
rect 105 326 106 327
rect 104 326 105 327
rect 68 326 69 327
rect 67 326 68 327
rect 66 326 67 327
rect 65 326 66 327
rect 64 326 65 327
rect 57 326 58 327
rect 56 326 57 327
rect 55 326 56 327
rect 54 326 55 327
rect 53 326 54 327
rect 35 326 36 327
rect 34 326 35 327
rect 33 326 34 327
rect 32 326 33 327
rect 31 326 32 327
rect 30 326 31 327
rect 18 326 19 327
rect 17 326 18 327
rect 186 327 187 328
rect 185 327 186 328
rect 184 327 185 328
rect 180 327 181 328
rect 179 327 180 328
rect 178 327 179 328
rect 177 327 178 328
rect 176 327 177 328
rect 175 327 176 328
rect 174 327 175 328
rect 173 327 174 328
rect 172 327 173 328
rect 171 327 172 328
rect 169 327 170 328
rect 168 327 169 328
rect 166 327 167 328
rect 165 327 166 328
rect 164 327 165 328
rect 114 327 115 328
rect 113 327 114 328
rect 112 327 113 328
rect 111 327 112 328
rect 110 327 111 328
rect 109 327 110 328
rect 108 327 109 328
rect 107 327 108 328
rect 106 327 107 328
rect 105 327 106 328
rect 104 327 105 328
rect 68 327 69 328
rect 67 327 68 328
rect 66 327 67 328
rect 65 327 66 328
rect 64 327 65 328
rect 57 327 58 328
rect 56 327 57 328
rect 55 327 56 328
rect 54 327 55 328
rect 53 327 54 328
rect 35 327 36 328
rect 34 327 35 328
rect 33 327 34 328
rect 32 327 33 328
rect 31 327 32 328
rect 30 327 31 328
rect 29 327 30 328
rect 28 327 29 328
rect 27 327 28 328
rect 26 327 27 328
rect 198 328 199 329
rect 197 328 198 329
rect 196 328 197 329
rect 195 328 196 329
rect 194 328 195 329
rect 193 328 194 329
rect 186 328 187 329
rect 185 328 186 329
rect 184 328 185 329
rect 180 328 181 329
rect 179 328 180 329
rect 178 328 179 329
rect 177 328 178 329
rect 176 328 177 329
rect 175 328 176 329
rect 174 328 175 329
rect 173 328 174 329
rect 172 328 173 329
rect 171 328 172 329
rect 169 328 170 329
rect 168 328 169 329
rect 166 328 167 329
rect 165 328 166 329
rect 164 328 165 329
rect 114 328 115 329
rect 113 328 114 329
rect 112 328 113 329
rect 111 328 112 329
rect 110 328 111 329
rect 109 328 110 329
rect 108 328 109 329
rect 107 328 108 329
rect 106 328 107 329
rect 105 328 106 329
rect 104 328 105 329
rect 68 328 69 329
rect 67 328 68 329
rect 66 328 67 329
rect 65 328 66 329
rect 64 328 65 329
rect 57 328 58 329
rect 56 328 57 329
rect 55 328 56 329
rect 54 328 55 329
rect 53 328 54 329
rect 35 328 36 329
rect 34 328 35 329
rect 33 328 34 329
rect 32 328 33 329
rect 31 328 32 329
rect 30 328 31 329
rect 29 328 30 329
rect 28 328 29 329
rect 27 328 28 329
rect 26 328 27 329
rect 25 328 26 329
rect 24 328 25 329
rect 23 328 24 329
rect 22 328 23 329
rect 21 328 22 329
rect 199 329 200 330
rect 198 329 199 330
rect 197 329 198 330
rect 196 329 197 330
rect 195 329 196 330
rect 194 329 195 330
rect 193 329 194 330
rect 186 329 187 330
rect 185 329 186 330
rect 184 329 185 330
rect 180 329 181 330
rect 179 329 180 330
rect 178 329 179 330
rect 177 329 178 330
rect 176 329 177 330
rect 175 329 176 330
rect 174 329 175 330
rect 173 329 174 330
rect 172 329 173 330
rect 171 329 172 330
rect 169 329 170 330
rect 168 329 169 330
rect 166 329 167 330
rect 165 329 166 330
rect 164 329 165 330
rect 114 329 115 330
rect 113 329 114 330
rect 112 329 113 330
rect 111 329 112 330
rect 110 329 111 330
rect 109 329 110 330
rect 108 329 109 330
rect 107 329 108 330
rect 106 329 107 330
rect 105 329 106 330
rect 104 329 105 330
rect 68 329 69 330
rect 67 329 68 330
rect 66 329 67 330
rect 65 329 66 330
rect 64 329 65 330
rect 57 329 58 330
rect 56 329 57 330
rect 55 329 56 330
rect 54 329 55 330
rect 53 329 54 330
rect 31 329 32 330
rect 30 329 31 330
rect 29 329 30 330
rect 28 329 29 330
rect 27 329 28 330
rect 26 329 27 330
rect 25 329 26 330
rect 24 329 25 330
rect 23 329 24 330
rect 22 329 23 330
rect 21 329 22 330
rect 20 329 21 330
rect 198 330 199 331
rect 195 330 196 331
rect 194 330 195 331
rect 193 330 194 331
rect 186 330 187 331
rect 185 330 186 331
rect 184 330 185 331
rect 180 330 181 331
rect 179 330 180 331
rect 178 330 179 331
rect 177 330 178 331
rect 176 330 177 331
rect 175 330 176 331
rect 174 330 175 331
rect 173 330 174 331
rect 172 330 173 331
rect 171 330 172 331
rect 169 330 170 331
rect 168 330 169 331
rect 166 330 167 331
rect 165 330 166 331
rect 164 330 165 331
rect 114 330 115 331
rect 113 330 114 331
rect 112 330 113 331
rect 111 330 112 331
rect 110 330 111 331
rect 109 330 110 331
rect 108 330 109 331
rect 107 330 108 331
rect 106 330 107 331
rect 105 330 106 331
rect 104 330 105 331
rect 68 330 69 331
rect 67 330 68 331
rect 66 330 67 331
rect 65 330 66 331
rect 64 330 65 331
rect 57 330 58 331
rect 56 330 57 331
rect 55 330 56 331
rect 54 330 55 331
rect 53 330 54 331
rect 30 330 31 331
rect 29 330 30 331
rect 28 330 29 331
rect 27 330 28 331
rect 26 330 27 331
rect 25 330 26 331
rect 24 330 25 331
rect 23 330 24 331
rect 22 330 23 331
rect 21 330 22 331
rect 20 330 21 331
rect 194 331 195 332
rect 193 331 194 332
rect 186 331 187 332
rect 185 331 186 332
rect 184 331 185 332
rect 180 331 181 332
rect 179 331 180 332
rect 178 331 179 332
rect 177 331 178 332
rect 176 331 177 332
rect 175 331 176 332
rect 173 331 174 332
rect 172 331 173 332
rect 171 331 172 332
rect 169 331 170 332
rect 168 331 169 332
rect 166 331 167 332
rect 165 331 166 332
rect 164 331 165 332
rect 114 331 115 332
rect 113 331 114 332
rect 112 331 113 332
rect 111 331 112 332
rect 110 331 111 332
rect 109 331 110 332
rect 108 331 109 332
rect 107 331 108 332
rect 106 331 107 332
rect 105 331 106 332
rect 104 331 105 332
rect 57 331 58 332
rect 56 331 57 332
rect 55 331 56 332
rect 54 331 55 332
rect 53 331 54 332
rect 31 331 32 332
rect 30 331 31 332
rect 29 331 30 332
rect 23 331 24 332
rect 22 331 23 332
rect 21 331 22 332
rect 198 332 199 333
rect 197 332 198 333
rect 196 332 197 333
rect 195 332 196 333
rect 194 332 195 333
rect 193 332 194 333
rect 186 332 187 333
rect 185 332 186 333
rect 184 332 185 333
rect 181 332 182 333
rect 180 332 181 333
rect 179 332 180 333
rect 177 332 178 333
rect 176 332 177 333
rect 175 332 176 333
rect 173 332 174 333
rect 172 332 173 333
rect 171 332 172 333
rect 169 332 170 333
rect 168 332 169 333
rect 166 332 167 333
rect 165 332 166 333
rect 164 332 165 333
rect 114 332 115 333
rect 113 332 114 333
rect 112 332 113 333
rect 111 332 112 333
rect 110 332 111 333
rect 109 332 110 333
rect 108 332 109 333
rect 107 332 108 333
rect 106 332 107 333
rect 105 332 106 333
rect 104 332 105 333
rect 57 332 58 333
rect 56 332 57 333
rect 55 332 56 333
rect 54 332 55 333
rect 53 332 54 333
rect 31 332 32 333
rect 30 332 31 333
rect 22 332 23 333
rect 21 332 22 333
rect 199 333 200 334
rect 198 333 199 334
rect 197 333 198 334
rect 196 333 197 334
rect 195 333 196 334
rect 194 333 195 334
rect 193 333 194 334
rect 185 333 186 334
rect 184 333 185 334
rect 183 333 184 334
rect 181 333 182 334
rect 180 333 181 334
rect 179 333 180 334
rect 177 333 178 334
rect 176 333 177 334
rect 175 333 176 334
rect 173 333 174 334
rect 172 333 173 334
rect 171 333 172 334
rect 169 333 170 334
rect 168 333 169 334
rect 166 333 167 334
rect 165 333 166 334
rect 164 333 165 334
rect 114 333 115 334
rect 113 333 114 334
rect 112 333 113 334
rect 111 333 112 334
rect 110 333 111 334
rect 109 333 110 334
rect 108 333 109 334
rect 107 333 108 334
rect 106 333 107 334
rect 105 333 106 334
rect 104 333 105 334
rect 31 333 32 334
rect 30 333 31 334
rect 29 333 30 334
rect 21 333 22 334
rect 20 333 21 334
rect 185 334 186 335
rect 184 334 185 335
rect 183 334 184 335
rect 181 334 182 335
rect 180 334 181 335
rect 179 334 180 335
rect 177 334 178 335
rect 176 334 177 335
rect 175 334 176 335
rect 173 334 174 335
rect 172 334 173 335
rect 171 334 172 335
rect 169 334 170 335
rect 168 334 169 335
rect 166 334 167 335
rect 165 334 166 335
rect 164 334 165 335
rect 114 334 115 335
rect 113 334 114 335
rect 112 334 113 335
rect 111 334 112 335
rect 110 334 111 335
rect 109 334 110 335
rect 108 334 109 335
rect 107 334 108 335
rect 106 334 107 335
rect 105 334 106 335
rect 104 334 105 335
rect 31 334 32 335
rect 30 334 31 335
rect 29 334 30 335
rect 28 334 29 335
rect 22 334 23 335
rect 21 334 22 335
rect 20 334 21 335
rect 198 335 199 336
rect 197 335 198 336
rect 196 335 197 336
rect 195 335 196 336
rect 194 335 195 336
rect 193 335 194 336
rect 191 335 192 336
rect 190 335 191 336
rect 185 335 186 336
rect 184 335 185 336
rect 183 335 184 336
rect 182 335 183 336
rect 181 335 182 336
rect 180 335 181 336
rect 179 335 180 336
rect 177 335 178 336
rect 176 335 177 336
rect 175 335 176 336
rect 173 335 174 336
rect 172 335 173 336
rect 171 335 172 336
rect 169 335 170 336
rect 168 335 169 336
rect 166 335 167 336
rect 165 335 166 336
rect 164 335 165 336
rect 114 335 115 336
rect 113 335 114 336
rect 112 335 113 336
rect 111 335 112 336
rect 110 335 111 336
rect 109 335 110 336
rect 108 335 109 336
rect 107 335 108 336
rect 106 335 107 336
rect 105 335 106 336
rect 104 335 105 336
rect 30 335 31 336
rect 29 335 30 336
rect 28 335 29 336
rect 27 335 28 336
rect 26 335 27 336
rect 25 335 26 336
rect 24 335 25 336
rect 23 335 24 336
rect 22 335 23 336
rect 21 335 22 336
rect 20 335 21 336
rect 199 336 200 337
rect 198 336 199 337
rect 197 336 198 337
rect 196 336 197 337
rect 195 336 196 337
rect 194 336 195 337
rect 193 336 194 337
rect 191 336 192 337
rect 190 336 191 337
rect 185 336 186 337
rect 184 336 185 337
rect 183 336 184 337
rect 182 336 183 337
rect 181 336 182 337
rect 180 336 181 337
rect 177 336 178 337
rect 176 336 177 337
rect 175 336 176 337
rect 173 336 174 337
rect 172 336 173 337
rect 171 336 172 337
rect 169 336 170 337
rect 168 336 169 337
rect 166 336 167 337
rect 165 336 166 337
rect 164 336 165 337
rect 114 336 115 337
rect 113 336 114 337
rect 112 336 113 337
rect 111 336 112 337
rect 110 336 111 337
rect 109 336 110 337
rect 108 336 109 337
rect 107 336 108 337
rect 106 336 107 337
rect 105 336 106 337
rect 104 336 105 337
rect 29 336 30 337
rect 28 336 29 337
rect 27 336 28 337
rect 26 336 27 337
rect 25 336 26 337
rect 24 336 25 337
rect 23 336 24 337
rect 22 336 23 337
rect 21 336 22 337
rect 198 337 199 338
rect 196 337 197 338
rect 191 337 192 338
rect 184 337 185 338
rect 183 337 184 338
rect 182 337 183 338
rect 181 337 182 338
rect 180 337 181 338
rect 177 337 178 338
rect 176 337 177 338
rect 175 337 176 338
rect 173 337 174 338
rect 172 337 173 338
rect 171 337 172 338
rect 169 337 170 338
rect 168 337 169 338
rect 166 337 167 338
rect 165 337 166 338
rect 164 337 165 338
rect 114 337 115 338
rect 113 337 114 338
rect 112 337 113 338
rect 111 337 112 338
rect 110 337 111 338
rect 109 337 110 338
rect 108 337 109 338
rect 107 337 108 338
rect 106 337 107 338
rect 105 337 106 338
rect 104 337 105 338
rect 80 337 81 338
rect 79 337 80 338
rect 78 337 79 338
rect 77 337 78 338
rect 76 337 77 338
rect 75 337 76 338
rect 74 337 75 338
rect 73 337 74 338
rect 72 337 73 338
rect 71 337 72 338
rect 70 337 71 338
rect 69 337 70 338
rect 68 337 69 338
rect 67 337 68 338
rect 66 337 67 338
rect 65 337 66 338
rect 64 337 65 338
rect 63 337 64 338
rect 62 337 63 338
rect 61 337 62 338
rect 60 337 61 338
rect 59 337 60 338
rect 58 337 59 338
rect 57 337 58 338
rect 56 337 57 338
rect 55 337 56 338
rect 54 337 55 338
rect 53 337 54 338
rect 28 337 29 338
rect 27 337 28 338
rect 26 337 27 338
rect 25 337 26 338
rect 24 337 25 338
rect 23 337 24 338
rect 22 337 23 338
rect 21 337 22 338
rect 197 338 198 339
rect 196 338 197 339
rect 195 338 196 339
rect 194 338 195 339
rect 183 338 184 339
rect 182 338 183 339
rect 181 338 182 339
rect 177 338 178 339
rect 176 338 177 339
rect 175 338 176 339
rect 172 338 173 339
rect 171 338 172 339
rect 114 338 115 339
rect 113 338 114 339
rect 112 338 113 339
rect 111 338 112 339
rect 110 338 111 339
rect 109 338 110 339
rect 108 338 109 339
rect 107 338 108 339
rect 106 338 107 339
rect 105 338 106 339
rect 104 338 105 339
rect 80 338 81 339
rect 79 338 80 339
rect 78 338 79 339
rect 77 338 78 339
rect 76 338 77 339
rect 75 338 76 339
rect 74 338 75 339
rect 73 338 74 339
rect 72 338 73 339
rect 71 338 72 339
rect 70 338 71 339
rect 69 338 70 339
rect 68 338 69 339
rect 67 338 68 339
rect 66 338 67 339
rect 65 338 66 339
rect 64 338 65 339
rect 63 338 64 339
rect 62 338 63 339
rect 61 338 62 339
rect 60 338 61 339
rect 59 338 60 339
rect 58 338 59 339
rect 57 338 58 339
rect 56 338 57 339
rect 55 338 56 339
rect 54 338 55 339
rect 53 338 54 339
rect 26 338 27 339
rect 25 338 26 339
rect 24 338 25 339
rect 23 338 24 339
rect 198 339 199 340
rect 197 339 198 340
rect 196 339 197 340
rect 195 339 196 340
rect 194 339 195 340
rect 193 339 194 340
rect 177 339 178 340
rect 176 339 177 340
rect 175 339 176 340
rect 114 339 115 340
rect 113 339 114 340
rect 112 339 113 340
rect 111 339 112 340
rect 110 339 111 340
rect 109 339 110 340
rect 108 339 109 340
rect 107 339 108 340
rect 106 339 107 340
rect 105 339 106 340
rect 104 339 105 340
rect 80 339 81 340
rect 79 339 80 340
rect 78 339 79 340
rect 77 339 78 340
rect 76 339 77 340
rect 75 339 76 340
rect 74 339 75 340
rect 73 339 74 340
rect 72 339 73 340
rect 71 339 72 340
rect 70 339 71 340
rect 69 339 70 340
rect 68 339 69 340
rect 67 339 68 340
rect 66 339 67 340
rect 65 339 66 340
rect 64 339 65 340
rect 63 339 64 340
rect 62 339 63 340
rect 61 339 62 340
rect 60 339 61 340
rect 59 339 60 340
rect 58 339 59 340
rect 57 339 58 340
rect 56 339 57 340
rect 55 339 56 340
rect 54 339 55 340
rect 53 339 54 340
rect 198 340 199 341
rect 197 340 198 341
rect 194 340 195 341
rect 193 340 194 341
rect 177 340 178 341
rect 176 340 177 341
rect 175 340 176 341
rect 114 340 115 341
rect 113 340 114 341
rect 112 340 113 341
rect 111 340 112 341
rect 110 340 111 341
rect 109 340 110 341
rect 108 340 109 341
rect 107 340 108 341
rect 106 340 107 341
rect 105 340 106 341
rect 104 340 105 341
rect 80 340 81 341
rect 79 340 80 341
rect 78 340 79 341
rect 77 340 78 341
rect 76 340 77 341
rect 75 340 76 341
rect 74 340 75 341
rect 73 340 74 341
rect 72 340 73 341
rect 71 340 72 341
rect 70 340 71 341
rect 69 340 70 341
rect 68 340 69 341
rect 67 340 68 341
rect 66 340 67 341
rect 65 340 66 341
rect 64 340 65 341
rect 63 340 64 341
rect 62 340 63 341
rect 61 340 62 341
rect 60 340 61 341
rect 59 340 60 341
rect 58 340 59 341
rect 57 340 58 341
rect 56 340 57 341
rect 55 340 56 341
rect 54 340 55 341
rect 53 340 54 341
rect 199 341 200 342
rect 198 341 199 342
rect 194 341 195 342
rect 193 341 194 342
rect 176 341 177 342
rect 114 341 115 342
rect 113 341 114 342
rect 112 341 113 342
rect 111 341 112 342
rect 110 341 111 342
rect 109 341 110 342
rect 108 341 109 342
rect 107 341 108 342
rect 106 341 107 342
rect 105 341 106 342
rect 104 341 105 342
rect 80 341 81 342
rect 79 341 80 342
rect 78 341 79 342
rect 77 341 78 342
rect 76 341 77 342
rect 75 341 76 342
rect 74 341 75 342
rect 73 341 74 342
rect 72 341 73 342
rect 71 341 72 342
rect 70 341 71 342
rect 69 341 70 342
rect 68 341 69 342
rect 67 341 68 342
rect 66 341 67 342
rect 65 341 66 342
rect 64 341 65 342
rect 63 341 64 342
rect 62 341 63 342
rect 61 341 62 342
rect 60 341 61 342
rect 59 341 60 342
rect 58 341 59 342
rect 57 341 58 342
rect 56 341 57 342
rect 55 341 56 342
rect 54 341 55 342
rect 53 341 54 342
rect 198 342 199 343
rect 194 342 195 343
rect 193 342 194 343
rect 114 342 115 343
rect 113 342 114 343
rect 112 342 113 343
rect 111 342 112 343
rect 110 342 111 343
rect 109 342 110 343
rect 108 342 109 343
rect 107 342 108 343
rect 106 342 107 343
rect 105 342 106 343
rect 104 342 105 343
rect 80 342 81 343
rect 79 342 80 343
rect 78 342 79 343
rect 77 342 78 343
rect 76 342 77 343
rect 75 342 76 343
rect 74 342 75 343
rect 73 342 74 343
rect 72 342 73 343
rect 71 342 72 343
rect 70 342 71 343
rect 69 342 70 343
rect 68 342 69 343
rect 67 342 68 343
rect 66 342 67 343
rect 65 342 66 343
rect 64 342 65 343
rect 63 342 64 343
rect 62 342 63 343
rect 61 342 62 343
rect 60 342 61 343
rect 59 342 60 343
rect 58 342 59 343
rect 57 342 58 343
rect 56 342 57 343
rect 55 342 56 343
rect 54 342 55 343
rect 53 342 54 343
rect 197 343 198 344
rect 114 343 115 344
rect 113 343 114 344
rect 112 343 113 344
rect 111 343 112 344
rect 110 343 111 344
rect 109 343 110 344
rect 108 343 109 344
rect 107 343 108 344
rect 106 343 107 344
rect 105 343 106 344
rect 104 343 105 344
rect 198 344 199 345
rect 197 344 198 345
rect 196 344 197 345
rect 194 344 195 345
rect 193 344 194 345
rect 114 344 115 345
rect 113 344 114 345
rect 112 344 113 345
rect 111 344 112 345
rect 110 344 111 345
rect 109 344 110 345
rect 108 344 109 345
rect 107 344 108 345
rect 106 344 107 345
rect 105 344 106 345
rect 104 344 105 345
rect 199 345 200 346
rect 198 345 199 346
rect 197 345 198 346
rect 196 345 197 346
rect 195 345 196 346
rect 194 345 195 346
rect 193 345 194 346
rect 31 345 32 346
rect 30 345 31 346
rect 199 346 200 347
rect 198 346 199 347
rect 196 346 197 347
rect 195 346 196 347
rect 194 346 195 347
rect 193 346 194 347
rect 31 346 32 347
rect 30 346 31 347
rect 29 346 30 347
rect 28 346 29 347
rect 27 346 28 347
rect 26 346 27 347
rect 198 347 199 348
rect 197 347 198 348
rect 196 347 197 348
rect 195 347 196 348
rect 194 347 195 348
rect 193 347 194 348
rect 31 347 32 348
rect 30 347 31 348
rect 29 347 30 348
rect 28 347 29 348
rect 27 347 28 348
rect 26 347 27 348
rect 25 347 26 348
rect 24 347 25 348
rect 23 347 24 348
rect 22 347 23 348
rect 21 347 22 348
rect 199 348 200 349
rect 198 348 199 349
rect 197 348 198 349
rect 196 348 197 349
rect 195 348 196 349
rect 194 348 195 349
rect 193 348 194 349
rect 80 348 81 349
rect 79 348 80 349
rect 78 348 79 349
rect 77 348 78 349
rect 76 348 77 349
rect 75 348 76 349
rect 74 348 75 349
rect 73 348 74 349
rect 72 348 73 349
rect 71 348 72 349
rect 70 348 71 349
rect 69 348 70 349
rect 68 348 69 349
rect 67 348 68 349
rect 66 348 67 349
rect 65 348 66 349
rect 64 348 65 349
rect 63 348 64 349
rect 62 348 63 349
rect 61 348 62 349
rect 60 348 61 349
rect 59 348 60 349
rect 58 348 59 349
rect 57 348 58 349
rect 56 348 57 349
rect 55 348 56 349
rect 54 348 55 349
rect 53 348 54 349
rect 30 348 31 349
rect 29 348 30 349
rect 28 348 29 349
rect 27 348 28 349
rect 26 348 27 349
rect 25 348 26 349
rect 24 348 25 349
rect 23 348 24 349
rect 22 348 23 349
rect 21 348 22 349
rect 20 348 21 349
rect 19 348 20 349
rect 18 348 19 349
rect 17 348 18 349
rect 198 349 199 350
rect 80 349 81 350
rect 79 349 80 350
rect 78 349 79 350
rect 77 349 78 350
rect 76 349 77 350
rect 75 349 76 350
rect 74 349 75 350
rect 73 349 74 350
rect 72 349 73 350
rect 71 349 72 350
rect 70 349 71 350
rect 69 349 70 350
rect 68 349 69 350
rect 67 349 68 350
rect 66 349 67 350
rect 65 349 66 350
rect 64 349 65 350
rect 63 349 64 350
rect 62 349 63 350
rect 61 349 62 350
rect 60 349 61 350
rect 59 349 60 350
rect 58 349 59 350
rect 57 349 58 350
rect 56 349 57 350
rect 55 349 56 350
rect 54 349 55 350
rect 53 349 54 350
rect 25 349 26 350
rect 24 349 25 350
rect 23 349 24 350
rect 22 349 23 350
rect 21 349 22 350
rect 20 349 21 350
rect 19 349 20 350
rect 18 349 19 350
rect 17 349 18 350
rect 16 349 17 350
rect 194 350 195 351
rect 193 350 194 351
rect 80 350 81 351
rect 79 350 80 351
rect 78 350 79 351
rect 77 350 78 351
rect 76 350 77 351
rect 75 350 76 351
rect 74 350 75 351
rect 73 350 74 351
rect 72 350 73 351
rect 71 350 72 351
rect 70 350 71 351
rect 69 350 70 351
rect 68 350 69 351
rect 67 350 68 351
rect 66 350 67 351
rect 65 350 66 351
rect 64 350 65 351
rect 63 350 64 351
rect 62 350 63 351
rect 61 350 62 351
rect 60 350 61 351
rect 59 350 60 351
rect 58 350 59 351
rect 57 350 58 351
rect 56 350 57 351
rect 55 350 56 351
rect 54 350 55 351
rect 53 350 54 351
rect 22 350 23 351
rect 21 350 22 351
rect 20 350 21 351
rect 19 350 20 351
rect 18 350 19 351
rect 17 350 18 351
rect 16 350 17 351
rect 198 351 199 352
rect 197 351 198 352
rect 196 351 197 352
rect 195 351 196 352
rect 194 351 195 352
rect 193 351 194 352
rect 192 351 193 352
rect 191 351 192 352
rect 175 351 176 352
rect 80 351 81 352
rect 79 351 80 352
rect 78 351 79 352
rect 77 351 78 352
rect 76 351 77 352
rect 75 351 76 352
rect 74 351 75 352
rect 73 351 74 352
rect 72 351 73 352
rect 71 351 72 352
rect 70 351 71 352
rect 69 351 70 352
rect 68 351 69 352
rect 67 351 68 352
rect 66 351 67 352
rect 65 351 66 352
rect 64 351 65 352
rect 63 351 64 352
rect 62 351 63 352
rect 61 351 62 352
rect 60 351 61 352
rect 59 351 60 352
rect 58 351 59 352
rect 57 351 58 352
rect 56 351 57 352
rect 55 351 56 352
rect 54 351 55 352
rect 53 351 54 352
rect 31 351 32 352
rect 30 351 31 352
rect 29 351 30 352
rect 28 351 29 352
rect 27 351 28 352
rect 26 351 27 352
rect 25 351 26 352
rect 24 351 25 352
rect 23 351 24 352
rect 22 351 23 352
rect 21 351 22 352
rect 20 351 21 352
rect 19 351 20 352
rect 18 351 19 352
rect 17 351 18 352
rect 16 351 17 352
rect 198 352 199 353
rect 197 352 198 353
rect 196 352 197 353
rect 195 352 196 353
rect 194 352 195 353
rect 193 352 194 353
rect 192 352 193 353
rect 191 352 192 353
rect 176 352 177 353
rect 175 352 176 353
rect 174 352 175 353
rect 80 352 81 353
rect 79 352 80 353
rect 78 352 79 353
rect 77 352 78 353
rect 76 352 77 353
rect 75 352 76 353
rect 74 352 75 353
rect 73 352 74 353
rect 72 352 73 353
rect 71 352 72 353
rect 70 352 71 353
rect 69 352 70 353
rect 68 352 69 353
rect 67 352 68 353
rect 66 352 67 353
rect 65 352 66 353
rect 64 352 65 353
rect 63 352 64 353
rect 62 352 63 353
rect 61 352 62 353
rect 60 352 61 353
rect 59 352 60 353
rect 58 352 59 353
rect 57 352 58 353
rect 56 352 57 353
rect 55 352 56 353
rect 54 352 55 353
rect 53 352 54 353
rect 31 352 32 353
rect 30 352 31 353
rect 29 352 30 353
rect 28 352 29 353
rect 27 352 28 353
rect 26 352 27 353
rect 25 352 26 353
rect 24 352 25 353
rect 23 352 24 353
rect 22 352 23 353
rect 21 352 22 353
rect 20 352 21 353
rect 19 352 20 353
rect 18 352 19 353
rect 17 352 18 353
rect 199 353 200 354
rect 198 353 199 354
rect 194 353 195 354
rect 193 353 194 354
rect 176 353 177 354
rect 175 353 176 354
rect 174 353 175 354
rect 80 353 81 354
rect 79 353 80 354
rect 78 353 79 354
rect 77 353 78 354
rect 76 353 77 354
rect 75 353 76 354
rect 74 353 75 354
rect 73 353 74 354
rect 72 353 73 354
rect 71 353 72 354
rect 70 353 71 354
rect 69 353 70 354
rect 68 353 69 354
rect 67 353 68 354
rect 66 353 67 354
rect 65 353 66 354
rect 64 353 65 354
rect 63 353 64 354
rect 62 353 63 354
rect 61 353 62 354
rect 60 353 61 354
rect 59 353 60 354
rect 58 353 59 354
rect 57 353 58 354
rect 56 353 57 354
rect 55 353 56 354
rect 54 353 55 354
rect 53 353 54 354
rect 31 353 32 354
rect 30 353 31 354
rect 29 353 30 354
rect 28 353 29 354
rect 27 353 28 354
rect 26 353 27 354
rect 198 354 199 355
rect 193 354 194 355
rect 176 354 177 355
rect 175 354 176 355
rect 174 354 175 355
rect 173 354 174 355
rect 69 354 70 355
rect 68 354 69 355
rect 67 354 68 355
rect 66 354 67 355
rect 65 354 66 355
rect 64 354 65 355
rect 57 354 58 355
rect 56 354 57 355
rect 55 354 56 355
rect 54 354 55 355
rect 53 354 54 355
rect 30 354 31 355
rect 29 354 30 355
rect 28 354 29 355
rect 27 354 28 355
rect 26 354 27 355
rect 25 354 26 355
rect 24 354 25 355
rect 198 355 199 356
rect 197 355 198 356
rect 196 355 197 356
rect 195 355 196 356
rect 194 355 195 356
rect 193 355 194 356
rect 191 355 192 356
rect 190 355 191 356
rect 175 355 176 356
rect 174 355 175 356
rect 173 355 174 356
rect 172 355 173 356
rect 68 355 69 356
rect 67 355 68 356
rect 66 355 67 356
rect 65 355 66 356
rect 64 355 65 356
rect 57 355 58 356
rect 56 355 57 356
rect 55 355 56 356
rect 54 355 55 356
rect 53 355 54 356
rect 28 355 29 356
rect 27 355 28 356
rect 26 355 27 356
rect 25 355 26 356
rect 24 355 25 356
rect 23 355 24 356
rect 22 355 23 356
rect 198 356 199 357
rect 197 356 198 357
rect 196 356 197 357
rect 195 356 196 357
rect 194 356 195 357
rect 193 356 194 357
rect 191 356 192 357
rect 190 356 191 357
rect 184 356 185 357
rect 183 356 184 357
rect 182 356 183 357
rect 181 356 182 357
rect 180 356 181 357
rect 179 356 180 357
rect 178 356 179 357
rect 175 356 176 357
rect 174 356 175 357
rect 173 356 174 357
rect 172 356 173 357
rect 171 356 172 357
rect 151 356 152 357
rect 150 356 151 357
rect 149 356 150 357
rect 148 356 149 357
rect 147 356 148 357
rect 146 356 147 357
rect 145 356 146 357
rect 144 356 145 357
rect 143 356 144 357
rect 142 356 143 357
rect 141 356 142 357
rect 140 356 141 357
rect 139 356 140 357
rect 138 356 139 357
rect 137 356 138 357
rect 136 356 137 357
rect 135 356 136 357
rect 134 356 135 357
rect 133 356 134 357
rect 132 356 133 357
rect 131 356 132 357
rect 130 356 131 357
rect 129 356 130 357
rect 128 356 129 357
rect 127 356 128 357
rect 126 356 127 357
rect 125 356 126 357
rect 124 356 125 357
rect 123 356 124 357
rect 122 356 123 357
rect 121 356 122 357
rect 120 356 121 357
rect 119 356 120 357
rect 118 356 119 357
rect 117 356 118 357
rect 116 356 117 357
rect 115 356 116 357
rect 114 356 115 357
rect 113 356 114 357
rect 112 356 113 357
rect 111 356 112 357
rect 110 356 111 357
rect 109 356 110 357
rect 108 356 109 357
rect 107 356 108 357
rect 106 356 107 357
rect 105 356 106 357
rect 104 356 105 357
rect 69 356 70 357
rect 68 356 69 357
rect 67 356 68 357
rect 66 356 67 357
rect 65 356 66 357
rect 64 356 65 357
rect 57 356 58 357
rect 56 356 57 357
rect 55 356 56 357
rect 54 356 55 357
rect 53 356 54 357
rect 26 356 27 357
rect 25 356 26 357
rect 24 356 25 357
rect 23 356 24 357
rect 22 356 23 357
rect 21 356 22 357
rect 20 356 21 357
rect 185 357 186 358
rect 184 357 185 358
rect 183 357 184 358
rect 182 357 183 358
rect 181 357 182 358
rect 180 357 181 358
rect 179 357 180 358
rect 178 357 179 358
rect 174 357 175 358
rect 173 357 174 358
rect 172 357 173 358
rect 171 357 172 358
rect 170 357 171 358
rect 169 357 170 358
rect 168 357 169 358
rect 151 357 152 358
rect 150 357 151 358
rect 149 357 150 358
rect 148 357 149 358
rect 147 357 148 358
rect 146 357 147 358
rect 145 357 146 358
rect 144 357 145 358
rect 143 357 144 358
rect 142 357 143 358
rect 141 357 142 358
rect 140 357 141 358
rect 139 357 140 358
rect 138 357 139 358
rect 137 357 138 358
rect 136 357 137 358
rect 135 357 136 358
rect 134 357 135 358
rect 133 357 134 358
rect 132 357 133 358
rect 131 357 132 358
rect 130 357 131 358
rect 129 357 130 358
rect 128 357 129 358
rect 127 357 128 358
rect 126 357 127 358
rect 125 357 126 358
rect 124 357 125 358
rect 123 357 124 358
rect 122 357 123 358
rect 121 357 122 358
rect 120 357 121 358
rect 119 357 120 358
rect 118 357 119 358
rect 117 357 118 358
rect 116 357 117 358
rect 115 357 116 358
rect 114 357 115 358
rect 113 357 114 358
rect 112 357 113 358
rect 111 357 112 358
rect 110 357 111 358
rect 109 357 110 358
rect 108 357 109 358
rect 107 357 108 358
rect 106 357 107 358
rect 105 357 106 358
rect 104 357 105 358
rect 69 357 70 358
rect 68 357 69 358
rect 67 357 68 358
rect 66 357 67 358
rect 65 357 66 358
rect 64 357 65 358
rect 57 357 58 358
rect 56 357 57 358
rect 55 357 56 358
rect 54 357 55 358
rect 53 357 54 358
rect 31 357 32 358
rect 30 357 31 358
rect 29 357 30 358
rect 23 357 24 358
rect 22 357 23 358
rect 21 357 22 358
rect 20 357 21 358
rect 19 357 20 358
rect 18 357 19 358
rect 198 358 199 359
rect 197 358 198 359
rect 196 358 197 359
rect 195 358 196 359
rect 194 358 195 359
rect 185 358 186 359
rect 184 358 185 359
rect 183 358 184 359
rect 182 358 183 359
rect 181 358 182 359
rect 180 358 181 359
rect 179 358 180 359
rect 178 358 179 359
rect 173 358 174 359
rect 172 358 173 359
rect 171 358 172 359
rect 170 358 171 359
rect 169 358 170 359
rect 168 358 169 359
rect 167 358 168 359
rect 166 358 167 359
rect 165 358 166 359
rect 164 358 165 359
rect 151 358 152 359
rect 150 358 151 359
rect 149 358 150 359
rect 148 358 149 359
rect 147 358 148 359
rect 146 358 147 359
rect 145 358 146 359
rect 144 358 145 359
rect 143 358 144 359
rect 142 358 143 359
rect 141 358 142 359
rect 140 358 141 359
rect 139 358 140 359
rect 138 358 139 359
rect 137 358 138 359
rect 136 358 137 359
rect 135 358 136 359
rect 134 358 135 359
rect 133 358 134 359
rect 132 358 133 359
rect 131 358 132 359
rect 130 358 131 359
rect 129 358 130 359
rect 128 358 129 359
rect 127 358 128 359
rect 126 358 127 359
rect 125 358 126 359
rect 124 358 125 359
rect 123 358 124 359
rect 122 358 123 359
rect 121 358 122 359
rect 120 358 121 359
rect 119 358 120 359
rect 118 358 119 359
rect 117 358 118 359
rect 116 358 117 359
rect 115 358 116 359
rect 114 358 115 359
rect 113 358 114 359
rect 112 358 113 359
rect 111 358 112 359
rect 110 358 111 359
rect 109 358 110 359
rect 108 358 109 359
rect 107 358 108 359
rect 106 358 107 359
rect 105 358 106 359
rect 104 358 105 359
rect 69 358 70 359
rect 68 358 69 359
rect 67 358 68 359
rect 66 358 67 359
rect 65 358 66 359
rect 64 358 65 359
rect 57 358 58 359
rect 56 358 57 359
rect 55 358 56 359
rect 54 358 55 359
rect 53 358 54 359
rect 31 358 32 359
rect 30 358 31 359
rect 29 358 30 359
rect 28 358 29 359
rect 27 358 28 359
rect 26 358 27 359
rect 25 358 26 359
rect 24 358 25 359
rect 22 358 23 359
rect 21 358 22 359
rect 20 358 21 359
rect 19 358 20 359
rect 18 358 19 359
rect 17 358 18 359
rect 198 359 199 360
rect 197 359 198 360
rect 196 359 197 360
rect 195 359 196 360
rect 194 359 195 360
rect 193 359 194 360
rect 185 359 186 360
rect 184 359 185 360
rect 183 359 184 360
rect 182 359 183 360
rect 172 359 173 360
rect 171 359 172 360
rect 170 359 171 360
rect 169 359 170 360
rect 168 359 169 360
rect 167 359 168 360
rect 166 359 167 360
rect 165 359 166 360
rect 164 359 165 360
rect 151 359 152 360
rect 150 359 151 360
rect 149 359 150 360
rect 148 359 149 360
rect 147 359 148 360
rect 146 359 147 360
rect 145 359 146 360
rect 144 359 145 360
rect 143 359 144 360
rect 142 359 143 360
rect 141 359 142 360
rect 140 359 141 360
rect 139 359 140 360
rect 138 359 139 360
rect 137 359 138 360
rect 136 359 137 360
rect 135 359 136 360
rect 134 359 135 360
rect 133 359 134 360
rect 132 359 133 360
rect 131 359 132 360
rect 130 359 131 360
rect 129 359 130 360
rect 128 359 129 360
rect 127 359 128 360
rect 126 359 127 360
rect 125 359 126 360
rect 124 359 125 360
rect 123 359 124 360
rect 122 359 123 360
rect 121 359 122 360
rect 120 359 121 360
rect 119 359 120 360
rect 118 359 119 360
rect 117 359 118 360
rect 116 359 117 360
rect 115 359 116 360
rect 114 359 115 360
rect 113 359 114 360
rect 112 359 113 360
rect 111 359 112 360
rect 110 359 111 360
rect 109 359 110 360
rect 108 359 109 360
rect 107 359 108 360
rect 106 359 107 360
rect 105 359 106 360
rect 104 359 105 360
rect 70 359 71 360
rect 69 359 70 360
rect 68 359 69 360
rect 67 359 68 360
rect 66 359 67 360
rect 65 359 66 360
rect 64 359 65 360
rect 57 359 58 360
rect 56 359 57 360
rect 55 359 56 360
rect 54 359 55 360
rect 53 359 54 360
rect 31 359 32 360
rect 30 359 31 360
rect 29 359 30 360
rect 28 359 29 360
rect 27 359 28 360
rect 26 359 27 360
rect 25 359 26 360
rect 24 359 25 360
rect 23 359 24 360
rect 22 359 23 360
rect 21 359 22 360
rect 20 359 21 360
rect 19 359 20 360
rect 18 359 19 360
rect 17 359 18 360
rect 16 359 17 360
rect 198 360 199 361
rect 194 360 195 361
rect 193 360 194 361
rect 185 360 186 361
rect 184 360 185 361
rect 183 360 184 361
rect 182 360 183 361
rect 173 360 174 361
rect 172 360 173 361
rect 171 360 172 361
rect 170 360 171 361
rect 169 360 170 361
rect 168 360 169 361
rect 167 360 168 361
rect 166 360 167 361
rect 165 360 166 361
rect 164 360 165 361
rect 151 360 152 361
rect 150 360 151 361
rect 149 360 150 361
rect 148 360 149 361
rect 147 360 148 361
rect 146 360 147 361
rect 145 360 146 361
rect 144 360 145 361
rect 143 360 144 361
rect 142 360 143 361
rect 141 360 142 361
rect 140 360 141 361
rect 139 360 140 361
rect 138 360 139 361
rect 137 360 138 361
rect 136 360 137 361
rect 135 360 136 361
rect 134 360 135 361
rect 133 360 134 361
rect 132 360 133 361
rect 131 360 132 361
rect 130 360 131 361
rect 129 360 130 361
rect 128 360 129 361
rect 127 360 128 361
rect 126 360 127 361
rect 125 360 126 361
rect 124 360 125 361
rect 123 360 124 361
rect 122 360 123 361
rect 121 360 122 361
rect 120 360 121 361
rect 119 360 120 361
rect 118 360 119 361
rect 117 360 118 361
rect 116 360 117 361
rect 115 360 116 361
rect 114 360 115 361
rect 113 360 114 361
rect 112 360 113 361
rect 111 360 112 361
rect 110 360 111 361
rect 109 360 110 361
rect 108 360 109 361
rect 107 360 108 361
rect 106 360 107 361
rect 105 360 106 361
rect 104 360 105 361
rect 72 360 73 361
rect 71 360 72 361
rect 70 360 71 361
rect 69 360 70 361
rect 68 360 69 361
rect 67 360 68 361
rect 66 360 67 361
rect 65 360 66 361
rect 64 360 65 361
rect 57 360 58 361
rect 56 360 57 361
rect 55 360 56 361
rect 54 360 55 361
rect 53 360 54 361
rect 28 360 29 361
rect 27 360 28 361
rect 26 360 27 361
rect 25 360 26 361
rect 24 360 25 361
rect 23 360 24 361
rect 22 360 23 361
rect 21 360 22 361
rect 20 360 21 361
rect 19 360 20 361
rect 18 360 19 361
rect 17 360 18 361
rect 16 360 17 361
rect 199 361 200 362
rect 198 361 199 362
rect 194 361 195 362
rect 193 361 194 362
rect 185 361 186 362
rect 184 361 185 362
rect 183 361 184 362
rect 182 361 183 362
rect 173 361 174 362
rect 172 361 173 362
rect 171 361 172 362
rect 170 361 171 362
rect 169 361 170 362
rect 168 361 169 362
rect 167 361 168 362
rect 166 361 167 362
rect 165 361 166 362
rect 164 361 165 362
rect 151 361 152 362
rect 150 361 151 362
rect 149 361 150 362
rect 148 361 149 362
rect 147 361 148 362
rect 146 361 147 362
rect 145 361 146 362
rect 144 361 145 362
rect 143 361 144 362
rect 142 361 143 362
rect 141 361 142 362
rect 140 361 141 362
rect 139 361 140 362
rect 138 361 139 362
rect 137 361 138 362
rect 136 361 137 362
rect 135 361 136 362
rect 134 361 135 362
rect 133 361 134 362
rect 132 361 133 362
rect 131 361 132 362
rect 130 361 131 362
rect 129 361 130 362
rect 128 361 129 362
rect 127 361 128 362
rect 126 361 127 362
rect 125 361 126 362
rect 124 361 125 362
rect 123 361 124 362
rect 122 361 123 362
rect 121 361 122 362
rect 120 361 121 362
rect 119 361 120 362
rect 118 361 119 362
rect 117 361 118 362
rect 116 361 117 362
rect 115 361 116 362
rect 114 361 115 362
rect 113 361 114 362
rect 112 361 113 362
rect 111 361 112 362
rect 110 361 111 362
rect 109 361 110 362
rect 108 361 109 362
rect 107 361 108 362
rect 106 361 107 362
rect 105 361 106 362
rect 104 361 105 362
rect 73 361 74 362
rect 72 361 73 362
rect 71 361 72 362
rect 70 361 71 362
rect 69 361 70 362
rect 68 361 69 362
rect 67 361 68 362
rect 66 361 67 362
rect 65 361 66 362
rect 64 361 65 362
rect 57 361 58 362
rect 56 361 57 362
rect 55 361 56 362
rect 54 361 55 362
rect 53 361 54 362
rect 23 361 24 362
rect 22 361 23 362
rect 21 361 22 362
rect 20 361 21 362
rect 19 361 20 362
rect 18 361 19 362
rect 17 361 18 362
rect 16 361 17 362
rect 198 362 199 363
rect 197 362 198 363
rect 196 362 197 363
rect 195 362 196 363
rect 194 362 195 363
rect 193 362 194 363
rect 185 362 186 363
rect 184 362 185 363
rect 183 362 184 363
rect 182 362 183 363
rect 174 362 175 363
rect 173 362 174 363
rect 172 362 173 363
rect 171 362 172 363
rect 170 362 171 363
rect 151 362 152 363
rect 150 362 151 363
rect 149 362 150 363
rect 148 362 149 363
rect 147 362 148 363
rect 146 362 147 363
rect 145 362 146 363
rect 144 362 145 363
rect 143 362 144 363
rect 142 362 143 363
rect 141 362 142 363
rect 140 362 141 363
rect 139 362 140 363
rect 138 362 139 363
rect 137 362 138 363
rect 136 362 137 363
rect 135 362 136 363
rect 134 362 135 363
rect 133 362 134 363
rect 132 362 133 363
rect 131 362 132 363
rect 130 362 131 363
rect 129 362 130 363
rect 128 362 129 363
rect 127 362 128 363
rect 126 362 127 363
rect 125 362 126 363
rect 124 362 125 363
rect 123 362 124 363
rect 122 362 123 363
rect 121 362 122 363
rect 120 362 121 363
rect 119 362 120 363
rect 118 362 119 363
rect 117 362 118 363
rect 116 362 117 363
rect 115 362 116 363
rect 114 362 115 363
rect 113 362 114 363
rect 112 362 113 363
rect 111 362 112 363
rect 110 362 111 363
rect 109 362 110 363
rect 108 362 109 363
rect 107 362 108 363
rect 106 362 107 363
rect 105 362 106 363
rect 104 362 105 363
rect 75 362 76 363
rect 74 362 75 363
rect 73 362 74 363
rect 72 362 73 363
rect 71 362 72 363
rect 70 362 71 363
rect 69 362 70 363
rect 68 362 69 363
rect 67 362 68 363
rect 66 362 67 363
rect 65 362 66 363
rect 64 362 65 363
rect 58 362 59 363
rect 57 362 58 363
rect 56 362 57 363
rect 55 362 56 363
rect 54 362 55 363
rect 53 362 54 363
rect 17 362 18 363
rect 198 363 199 364
rect 197 363 198 364
rect 196 363 197 364
rect 195 363 196 364
rect 194 363 195 364
rect 193 363 194 364
rect 185 363 186 364
rect 184 363 185 364
rect 183 363 184 364
rect 182 363 183 364
rect 175 363 176 364
rect 174 363 175 364
rect 173 363 174 364
rect 172 363 173 364
rect 171 363 172 364
rect 151 363 152 364
rect 150 363 151 364
rect 149 363 150 364
rect 148 363 149 364
rect 147 363 148 364
rect 146 363 147 364
rect 145 363 146 364
rect 144 363 145 364
rect 143 363 144 364
rect 142 363 143 364
rect 141 363 142 364
rect 140 363 141 364
rect 139 363 140 364
rect 138 363 139 364
rect 137 363 138 364
rect 136 363 137 364
rect 135 363 136 364
rect 134 363 135 364
rect 133 363 134 364
rect 132 363 133 364
rect 131 363 132 364
rect 130 363 131 364
rect 129 363 130 364
rect 128 363 129 364
rect 127 363 128 364
rect 126 363 127 364
rect 125 363 126 364
rect 124 363 125 364
rect 123 363 124 364
rect 122 363 123 364
rect 121 363 122 364
rect 120 363 121 364
rect 119 363 120 364
rect 118 363 119 364
rect 117 363 118 364
rect 116 363 117 364
rect 115 363 116 364
rect 114 363 115 364
rect 113 363 114 364
rect 112 363 113 364
rect 111 363 112 364
rect 110 363 111 364
rect 109 363 110 364
rect 108 363 109 364
rect 107 363 108 364
rect 106 363 107 364
rect 105 363 106 364
rect 104 363 105 364
rect 76 363 77 364
rect 75 363 76 364
rect 74 363 75 364
rect 73 363 74 364
rect 72 363 73 364
rect 71 363 72 364
rect 70 363 71 364
rect 69 363 70 364
rect 68 363 69 364
rect 67 363 68 364
rect 66 363 67 364
rect 65 363 66 364
rect 64 363 65 364
rect 58 363 59 364
rect 57 363 58 364
rect 56 363 57 364
rect 55 363 56 364
rect 54 363 55 364
rect 53 363 54 364
rect 31 363 32 364
rect 30 363 31 364
rect 29 363 30 364
rect 196 364 197 365
rect 185 364 186 365
rect 184 364 185 365
rect 183 364 184 365
rect 182 364 183 365
rect 175 364 176 365
rect 174 364 175 365
rect 173 364 174 365
rect 172 364 173 365
rect 151 364 152 365
rect 150 364 151 365
rect 149 364 150 365
rect 148 364 149 365
rect 147 364 148 365
rect 146 364 147 365
rect 145 364 146 365
rect 144 364 145 365
rect 143 364 144 365
rect 142 364 143 365
rect 141 364 142 365
rect 140 364 141 365
rect 139 364 140 365
rect 138 364 139 365
rect 137 364 138 365
rect 136 364 137 365
rect 135 364 136 365
rect 134 364 135 365
rect 133 364 134 365
rect 132 364 133 365
rect 131 364 132 365
rect 130 364 131 365
rect 129 364 130 365
rect 128 364 129 365
rect 127 364 128 365
rect 126 364 127 365
rect 125 364 126 365
rect 124 364 125 365
rect 123 364 124 365
rect 122 364 123 365
rect 121 364 122 365
rect 120 364 121 365
rect 119 364 120 365
rect 118 364 119 365
rect 117 364 118 365
rect 116 364 117 365
rect 115 364 116 365
rect 114 364 115 365
rect 113 364 114 365
rect 112 364 113 365
rect 111 364 112 365
rect 110 364 111 365
rect 109 364 110 365
rect 108 364 109 365
rect 107 364 108 365
rect 106 364 107 365
rect 105 364 106 365
rect 104 364 105 365
rect 77 364 78 365
rect 76 364 77 365
rect 75 364 76 365
rect 74 364 75 365
rect 73 364 74 365
rect 72 364 73 365
rect 71 364 72 365
rect 70 364 71 365
rect 69 364 70 365
rect 68 364 69 365
rect 67 364 68 365
rect 66 364 67 365
rect 65 364 66 365
rect 64 364 65 365
rect 63 364 64 365
rect 59 364 60 365
rect 58 364 59 365
rect 57 364 58 365
rect 56 364 57 365
rect 55 364 56 365
rect 54 364 55 365
rect 53 364 54 365
rect 31 364 32 365
rect 30 364 31 365
rect 29 364 30 365
rect 28 364 29 365
rect 27 364 28 365
rect 26 364 27 365
rect 25 364 26 365
rect 198 365 199 366
rect 197 365 198 366
rect 195 365 196 366
rect 194 365 195 366
rect 193 365 194 366
rect 185 365 186 366
rect 184 365 185 366
rect 183 365 184 366
rect 182 365 183 366
rect 176 365 177 366
rect 175 365 176 366
rect 174 365 175 366
rect 173 365 174 366
rect 151 365 152 366
rect 150 365 151 366
rect 149 365 150 366
rect 148 365 149 366
rect 147 365 148 366
rect 146 365 147 366
rect 145 365 146 366
rect 144 365 145 366
rect 143 365 144 366
rect 142 365 143 366
rect 141 365 142 366
rect 140 365 141 366
rect 139 365 140 366
rect 138 365 139 366
rect 137 365 138 366
rect 136 365 137 366
rect 135 365 136 366
rect 134 365 135 366
rect 133 365 134 366
rect 132 365 133 366
rect 131 365 132 366
rect 130 365 131 366
rect 129 365 130 366
rect 128 365 129 366
rect 127 365 128 366
rect 126 365 127 366
rect 125 365 126 366
rect 124 365 125 366
rect 123 365 124 366
rect 122 365 123 366
rect 121 365 122 366
rect 120 365 121 366
rect 119 365 120 366
rect 118 365 119 366
rect 117 365 118 366
rect 116 365 117 366
rect 115 365 116 366
rect 114 365 115 366
rect 113 365 114 366
rect 112 365 113 366
rect 111 365 112 366
rect 110 365 111 366
rect 109 365 110 366
rect 108 365 109 366
rect 107 365 108 366
rect 106 365 107 366
rect 105 365 106 366
rect 104 365 105 366
rect 79 365 80 366
rect 78 365 79 366
rect 77 365 78 366
rect 76 365 77 366
rect 75 365 76 366
rect 74 365 75 366
rect 73 365 74 366
rect 72 365 73 366
rect 71 365 72 366
rect 70 365 71 366
rect 67 365 68 366
rect 66 365 67 366
rect 65 365 66 366
rect 64 365 65 366
rect 63 365 64 366
rect 62 365 63 366
rect 61 365 62 366
rect 60 365 61 366
rect 59 365 60 366
rect 58 365 59 366
rect 57 365 58 366
rect 56 365 57 366
rect 55 365 56 366
rect 54 365 55 366
rect 31 365 32 366
rect 30 365 31 366
rect 29 365 30 366
rect 28 365 29 366
rect 27 365 28 366
rect 26 365 27 366
rect 25 365 26 366
rect 24 365 25 366
rect 23 365 24 366
rect 22 365 23 366
rect 21 365 22 366
rect 20 365 21 366
rect 199 366 200 367
rect 198 366 199 367
rect 197 366 198 367
rect 196 366 197 367
rect 195 366 196 367
rect 194 366 195 367
rect 193 366 194 367
rect 185 366 186 367
rect 184 366 185 367
rect 183 366 184 367
rect 182 366 183 367
rect 176 366 177 367
rect 175 366 176 367
rect 174 366 175 367
rect 173 366 174 367
rect 151 366 152 367
rect 150 366 151 367
rect 149 366 150 367
rect 148 366 149 367
rect 147 366 148 367
rect 146 366 147 367
rect 145 366 146 367
rect 144 366 145 367
rect 143 366 144 367
rect 142 366 143 367
rect 141 366 142 367
rect 140 366 141 367
rect 139 366 140 367
rect 138 366 139 367
rect 137 366 138 367
rect 136 366 137 367
rect 135 366 136 367
rect 134 366 135 367
rect 133 366 134 367
rect 132 366 133 367
rect 131 366 132 367
rect 130 366 131 367
rect 129 366 130 367
rect 128 366 129 367
rect 127 366 128 367
rect 126 366 127 367
rect 125 366 126 367
rect 124 366 125 367
rect 123 366 124 367
rect 122 366 123 367
rect 121 366 122 367
rect 120 366 121 367
rect 119 366 120 367
rect 118 366 119 367
rect 117 366 118 367
rect 116 366 117 367
rect 115 366 116 367
rect 114 366 115 367
rect 113 366 114 367
rect 112 366 113 367
rect 111 366 112 367
rect 110 366 111 367
rect 109 366 110 367
rect 108 366 109 367
rect 107 366 108 367
rect 106 366 107 367
rect 105 366 106 367
rect 104 366 105 367
rect 80 366 81 367
rect 79 366 80 367
rect 78 366 79 367
rect 77 366 78 367
rect 76 366 77 367
rect 75 366 76 367
rect 74 366 75 367
rect 73 366 74 367
rect 72 366 73 367
rect 71 366 72 367
rect 67 366 68 367
rect 66 366 67 367
rect 65 366 66 367
rect 64 366 65 367
rect 63 366 64 367
rect 62 366 63 367
rect 61 366 62 367
rect 60 366 61 367
rect 59 366 60 367
rect 58 366 59 367
rect 57 366 58 367
rect 56 366 57 367
rect 55 366 56 367
rect 54 366 55 367
rect 30 366 31 367
rect 29 366 30 367
rect 28 366 29 367
rect 27 366 28 367
rect 26 366 27 367
rect 25 366 26 367
rect 24 366 25 367
rect 23 366 24 367
rect 22 366 23 367
rect 21 366 22 367
rect 20 366 21 367
rect 19 366 20 367
rect 18 366 19 367
rect 17 366 18 367
rect 198 367 199 368
rect 195 367 196 368
rect 194 367 195 368
rect 193 367 194 368
rect 185 367 186 368
rect 184 367 185 368
rect 183 367 184 368
rect 182 367 183 368
rect 174 367 175 368
rect 151 367 152 368
rect 150 367 151 368
rect 149 367 150 368
rect 148 367 149 368
rect 147 367 148 368
rect 146 367 147 368
rect 145 367 146 368
rect 144 367 145 368
rect 143 367 144 368
rect 142 367 143 368
rect 141 367 142 368
rect 140 367 141 368
rect 139 367 140 368
rect 138 367 139 368
rect 137 367 138 368
rect 136 367 137 368
rect 135 367 136 368
rect 134 367 135 368
rect 133 367 134 368
rect 132 367 133 368
rect 131 367 132 368
rect 130 367 131 368
rect 129 367 130 368
rect 128 367 129 368
rect 127 367 128 368
rect 126 367 127 368
rect 125 367 126 368
rect 124 367 125 368
rect 123 367 124 368
rect 122 367 123 368
rect 121 367 122 368
rect 120 367 121 368
rect 119 367 120 368
rect 118 367 119 368
rect 117 367 118 368
rect 116 367 117 368
rect 115 367 116 368
rect 114 367 115 368
rect 113 367 114 368
rect 112 367 113 368
rect 111 367 112 368
rect 110 367 111 368
rect 109 367 110 368
rect 108 367 109 368
rect 107 367 108 368
rect 106 367 107 368
rect 105 367 106 368
rect 104 367 105 368
rect 80 367 81 368
rect 79 367 80 368
rect 78 367 79 368
rect 77 367 78 368
rect 76 367 77 368
rect 75 367 76 368
rect 74 367 75 368
rect 73 367 74 368
rect 72 367 73 368
rect 66 367 67 368
rect 65 367 66 368
rect 64 367 65 368
rect 63 367 64 368
rect 62 367 63 368
rect 61 367 62 368
rect 60 367 61 368
rect 59 367 60 368
rect 58 367 59 368
rect 57 367 58 368
rect 56 367 57 368
rect 55 367 56 368
rect 26 367 27 368
rect 25 367 26 368
rect 24 367 25 368
rect 23 367 24 368
rect 22 367 23 368
rect 21 367 22 368
rect 20 367 21 368
rect 19 367 20 368
rect 18 367 19 368
rect 17 367 18 368
rect 16 367 17 368
rect 194 368 195 369
rect 193 368 194 369
rect 185 368 186 369
rect 184 368 185 369
rect 183 368 184 369
rect 182 368 183 369
rect 151 368 152 369
rect 150 368 151 369
rect 149 368 150 369
rect 148 368 149 369
rect 147 368 148 369
rect 146 368 147 369
rect 145 368 146 369
rect 144 368 145 369
rect 143 368 144 369
rect 142 368 143 369
rect 141 368 142 369
rect 140 368 141 369
rect 139 368 140 369
rect 138 368 139 369
rect 137 368 138 369
rect 136 368 137 369
rect 135 368 136 369
rect 134 368 135 369
rect 133 368 134 369
rect 132 368 133 369
rect 131 368 132 369
rect 130 368 131 369
rect 129 368 130 369
rect 128 368 129 369
rect 127 368 128 369
rect 126 368 127 369
rect 125 368 126 369
rect 124 368 125 369
rect 123 368 124 369
rect 122 368 123 369
rect 121 368 122 369
rect 120 368 121 369
rect 119 368 120 369
rect 118 368 119 369
rect 117 368 118 369
rect 116 368 117 369
rect 115 368 116 369
rect 114 368 115 369
rect 113 368 114 369
rect 112 368 113 369
rect 111 368 112 369
rect 110 368 111 369
rect 109 368 110 369
rect 108 368 109 369
rect 107 368 108 369
rect 106 368 107 369
rect 105 368 106 369
rect 104 368 105 369
rect 80 368 81 369
rect 79 368 80 369
rect 78 368 79 369
rect 77 368 78 369
rect 76 368 77 369
rect 75 368 76 369
rect 74 368 75 369
rect 73 368 74 369
rect 66 368 67 369
rect 65 368 66 369
rect 64 368 65 369
rect 63 368 64 369
rect 62 368 63 369
rect 61 368 62 369
rect 60 368 61 369
rect 59 368 60 369
rect 58 368 59 369
rect 57 368 58 369
rect 56 368 57 369
rect 55 368 56 369
rect 25 368 26 369
rect 24 368 25 369
rect 23 368 24 369
rect 21 368 22 369
rect 20 368 21 369
rect 19 368 20 369
rect 18 368 19 369
rect 17 368 18 369
rect 16 368 17 369
rect 198 369 199 370
rect 197 369 198 370
rect 196 369 197 370
rect 195 369 196 370
rect 194 369 195 370
rect 193 369 194 370
rect 185 369 186 370
rect 184 369 185 370
rect 183 369 184 370
rect 182 369 183 370
rect 151 369 152 370
rect 150 369 151 370
rect 149 369 150 370
rect 148 369 149 370
rect 147 369 148 370
rect 146 369 147 370
rect 145 369 146 370
rect 144 369 145 370
rect 143 369 144 370
rect 142 369 143 370
rect 141 369 142 370
rect 140 369 141 370
rect 139 369 140 370
rect 138 369 139 370
rect 137 369 138 370
rect 136 369 137 370
rect 135 369 136 370
rect 134 369 135 370
rect 133 369 134 370
rect 132 369 133 370
rect 131 369 132 370
rect 130 369 131 370
rect 129 369 130 370
rect 128 369 129 370
rect 127 369 128 370
rect 126 369 127 370
rect 125 369 126 370
rect 124 369 125 370
rect 123 369 124 370
rect 122 369 123 370
rect 121 369 122 370
rect 120 369 121 370
rect 119 369 120 370
rect 118 369 119 370
rect 117 369 118 370
rect 116 369 117 370
rect 115 369 116 370
rect 114 369 115 370
rect 113 369 114 370
rect 112 369 113 370
rect 111 369 112 370
rect 110 369 111 370
rect 109 369 110 370
rect 108 369 109 370
rect 107 369 108 370
rect 106 369 107 370
rect 105 369 106 370
rect 104 369 105 370
rect 80 369 81 370
rect 79 369 80 370
rect 78 369 79 370
rect 77 369 78 370
rect 76 369 77 370
rect 75 369 76 370
rect 65 369 66 370
rect 64 369 65 370
rect 63 369 64 370
rect 62 369 63 370
rect 61 369 62 370
rect 60 369 61 370
rect 59 369 60 370
rect 58 369 59 370
rect 57 369 58 370
rect 56 369 57 370
rect 25 369 26 370
rect 24 369 25 370
rect 23 369 24 370
rect 18 369 19 370
rect 17 369 18 370
rect 16 369 17 370
rect 199 370 200 371
rect 198 370 199 371
rect 197 370 198 371
rect 196 370 197 371
rect 195 370 196 371
rect 194 370 195 371
rect 193 370 194 371
rect 185 370 186 371
rect 184 370 185 371
rect 183 370 184 371
rect 182 370 183 371
rect 179 370 180 371
rect 178 370 179 371
rect 177 370 178 371
rect 176 370 177 371
rect 175 370 176 371
rect 174 370 175 371
rect 173 370 174 371
rect 172 370 173 371
rect 171 370 172 371
rect 170 370 171 371
rect 169 370 170 371
rect 168 370 169 371
rect 167 370 168 371
rect 166 370 167 371
rect 165 370 166 371
rect 164 370 165 371
rect 151 370 152 371
rect 150 370 151 371
rect 149 370 150 371
rect 148 370 149 371
rect 147 370 148 371
rect 146 370 147 371
rect 145 370 146 371
rect 144 370 145 371
rect 143 370 144 371
rect 142 370 143 371
rect 141 370 142 371
rect 140 370 141 371
rect 139 370 140 371
rect 138 370 139 371
rect 137 370 138 371
rect 136 370 137 371
rect 135 370 136 371
rect 134 370 135 371
rect 133 370 134 371
rect 132 370 133 371
rect 131 370 132 371
rect 130 370 131 371
rect 129 370 130 371
rect 128 370 129 371
rect 127 370 128 371
rect 126 370 127 371
rect 125 370 126 371
rect 124 370 125 371
rect 123 370 124 371
rect 122 370 123 371
rect 121 370 122 371
rect 120 370 121 371
rect 119 370 120 371
rect 118 370 119 371
rect 117 370 118 371
rect 116 370 117 371
rect 115 370 116 371
rect 114 370 115 371
rect 113 370 114 371
rect 112 370 113 371
rect 111 370 112 371
rect 110 370 111 371
rect 109 370 110 371
rect 108 370 109 371
rect 107 370 108 371
rect 106 370 107 371
rect 105 370 106 371
rect 104 370 105 371
rect 80 370 81 371
rect 79 370 80 371
rect 78 370 79 371
rect 77 370 78 371
rect 63 370 64 371
rect 62 370 63 371
rect 61 370 62 371
rect 60 370 61 371
rect 59 370 60 371
rect 58 370 59 371
rect 25 370 26 371
rect 24 370 25 371
rect 23 370 24 371
rect 18 370 19 371
rect 17 370 18 371
rect 16 370 17 371
rect 185 371 186 372
rect 184 371 185 372
rect 183 371 184 372
rect 182 371 183 372
rect 179 371 180 372
rect 178 371 179 372
rect 177 371 178 372
rect 176 371 177 372
rect 175 371 176 372
rect 174 371 175 372
rect 173 371 174 372
rect 172 371 173 372
rect 171 371 172 372
rect 170 371 171 372
rect 169 371 170 372
rect 168 371 169 372
rect 167 371 168 372
rect 166 371 167 372
rect 165 371 166 372
rect 164 371 165 372
rect 151 371 152 372
rect 150 371 151 372
rect 149 371 150 372
rect 148 371 149 372
rect 147 371 148 372
rect 146 371 147 372
rect 145 371 146 372
rect 144 371 145 372
rect 143 371 144 372
rect 142 371 143 372
rect 141 371 142 372
rect 140 371 141 372
rect 139 371 140 372
rect 138 371 139 372
rect 137 371 138 372
rect 136 371 137 372
rect 135 371 136 372
rect 134 371 135 372
rect 133 371 134 372
rect 132 371 133 372
rect 131 371 132 372
rect 130 371 131 372
rect 129 371 130 372
rect 128 371 129 372
rect 127 371 128 372
rect 126 371 127 372
rect 125 371 126 372
rect 124 371 125 372
rect 123 371 124 372
rect 122 371 123 372
rect 121 371 122 372
rect 120 371 121 372
rect 119 371 120 372
rect 118 371 119 372
rect 117 371 118 372
rect 116 371 117 372
rect 115 371 116 372
rect 114 371 115 372
rect 113 371 114 372
rect 112 371 113 372
rect 111 371 112 372
rect 110 371 111 372
rect 109 371 110 372
rect 108 371 109 372
rect 107 371 108 372
rect 106 371 107 372
rect 105 371 106 372
rect 104 371 105 372
rect 80 371 81 372
rect 79 371 80 372
rect 78 371 79 372
rect 25 371 26 372
rect 24 371 25 372
rect 23 371 24 372
rect 18 371 19 372
rect 17 371 18 372
rect 16 371 17 372
rect 198 372 199 373
rect 195 372 196 373
rect 194 372 195 373
rect 185 372 186 373
rect 184 372 185 373
rect 183 372 184 373
rect 182 372 183 373
rect 179 372 180 373
rect 178 372 179 373
rect 177 372 178 373
rect 176 372 177 373
rect 175 372 176 373
rect 174 372 175 373
rect 173 372 174 373
rect 172 372 173 373
rect 171 372 172 373
rect 170 372 171 373
rect 169 372 170 373
rect 168 372 169 373
rect 167 372 168 373
rect 166 372 167 373
rect 165 372 166 373
rect 164 372 165 373
rect 151 372 152 373
rect 150 372 151 373
rect 149 372 150 373
rect 148 372 149 373
rect 147 372 148 373
rect 146 372 147 373
rect 145 372 146 373
rect 144 372 145 373
rect 143 372 144 373
rect 142 372 143 373
rect 141 372 142 373
rect 140 372 141 373
rect 139 372 140 373
rect 138 372 139 373
rect 137 372 138 373
rect 136 372 137 373
rect 135 372 136 373
rect 134 372 135 373
rect 133 372 134 373
rect 132 372 133 373
rect 131 372 132 373
rect 130 372 131 373
rect 129 372 130 373
rect 128 372 129 373
rect 127 372 128 373
rect 126 372 127 373
rect 125 372 126 373
rect 124 372 125 373
rect 123 372 124 373
rect 122 372 123 373
rect 121 372 122 373
rect 120 372 121 373
rect 119 372 120 373
rect 118 372 119 373
rect 117 372 118 373
rect 116 372 117 373
rect 115 372 116 373
rect 114 372 115 373
rect 113 372 114 373
rect 112 372 113 373
rect 111 372 112 373
rect 110 372 111 373
rect 109 372 110 373
rect 108 372 109 373
rect 107 372 108 373
rect 106 372 107 373
rect 105 372 106 373
rect 104 372 105 373
rect 80 372 81 373
rect 25 372 26 373
rect 24 372 25 373
rect 23 372 24 373
rect 18 372 19 373
rect 17 372 18 373
rect 16 372 17 373
rect 199 373 200 374
rect 198 373 199 374
rect 196 373 197 374
rect 195 373 196 374
rect 194 373 195 374
rect 193 373 194 374
rect 185 373 186 374
rect 184 373 185 374
rect 183 373 184 374
rect 182 373 183 374
rect 179 373 180 374
rect 178 373 179 374
rect 177 373 178 374
rect 176 373 177 374
rect 175 373 176 374
rect 174 373 175 374
rect 173 373 174 374
rect 172 373 173 374
rect 171 373 172 374
rect 170 373 171 374
rect 169 373 170 374
rect 168 373 169 374
rect 167 373 168 374
rect 166 373 167 374
rect 165 373 166 374
rect 164 373 165 374
rect 151 373 152 374
rect 150 373 151 374
rect 149 373 150 374
rect 148 373 149 374
rect 147 373 148 374
rect 146 373 147 374
rect 145 373 146 374
rect 144 373 145 374
rect 143 373 144 374
rect 142 373 143 374
rect 141 373 142 374
rect 140 373 141 374
rect 139 373 140 374
rect 138 373 139 374
rect 137 373 138 374
rect 136 373 137 374
rect 135 373 136 374
rect 134 373 135 374
rect 133 373 134 374
rect 132 373 133 374
rect 131 373 132 374
rect 130 373 131 374
rect 129 373 130 374
rect 128 373 129 374
rect 127 373 128 374
rect 126 373 127 374
rect 125 373 126 374
rect 124 373 125 374
rect 123 373 124 374
rect 122 373 123 374
rect 121 373 122 374
rect 120 373 121 374
rect 119 373 120 374
rect 118 373 119 374
rect 117 373 118 374
rect 116 373 117 374
rect 115 373 116 374
rect 114 373 115 374
rect 113 373 114 374
rect 112 373 113 374
rect 111 373 112 374
rect 110 373 111 374
rect 109 373 110 374
rect 108 373 109 374
rect 107 373 108 374
rect 106 373 107 374
rect 105 373 106 374
rect 104 373 105 374
rect 25 373 26 374
rect 24 373 25 374
rect 23 373 24 374
rect 22 373 23 374
rect 19 373 20 374
rect 18 373 19 374
rect 17 373 18 374
rect 199 374 200 375
rect 198 374 199 375
rect 197 374 198 375
rect 196 374 197 375
rect 195 374 196 375
rect 194 374 195 375
rect 193 374 194 375
rect 184 374 185 375
rect 183 374 184 375
rect 151 374 152 375
rect 150 374 151 375
rect 149 374 150 375
rect 148 374 149 375
rect 147 374 148 375
rect 146 374 147 375
rect 145 374 146 375
rect 144 374 145 375
rect 143 374 144 375
rect 142 374 143 375
rect 141 374 142 375
rect 140 374 141 375
rect 139 374 140 375
rect 138 374 139 375
rect 137 374 138 375
rect 136 374 137 375
rect 135 374 136 375
rect 134 374 135 375
rect 133 374 134 375
rect 132 374 133 375
rect 131 374 132 375
rect 130 374 131 375
rect 129 374 130 375
rect 128 374 129 375
rect 127 374 128 375
rect 126 374 127 375
rect 125 374 126 375
rect 124 374 125 375
rect 123 374 124 375
rect 122 374 123 375
rect 121 374 122 375
rect 120 374 121 375
rect 119 374 120 375
rect 118 374 119 375
rect 117 374 118 375
rect 116 374 117 375
rect 115 374 116 375
rect 114 374 115 375
rect 113 374 114 375
rect 112 374 113 375
rect 111 374 112 375
rect 110 374 111 375
rect 109 374 110 375
rect 108 374 109 375
rect 107 374 108 375
rect 106 374 107 375
rect 105 374 106 375
rect 104 374 105 375
rect 24 374 25 375
rect 23 374 24 375
rect 22 374 23 375
rect 21 374 22 375
rect 20 374 21 375
rect 19 374 20 375
rect 18 374 19 375
rect 17 374 18 375
rect 198 375 199 376
rect 197 375 198 376
rect 196 375 197 376
rect 194 375 195 376
rect 193 375 194 376
rect 151 375 152 376
rect 150 375 151 376
rect 149 375 150 376
rect 148 375 149 376
rect 147 375 148 376
rect 146 375 147 376
rect 145 375 146 376
rect 144 375 145 376
rect 143 375 144 376
rect 142 375 143 376
rect 141 375 142 376
rect 140 375 141 376
rect 139 375 140 376
rect 138 375 139 376
rect 137 375 138 376
rect 136 375 137 376
rect 135 375 136 376
rect 134 375 135 376
rect 133 375 134 376
rect 132 375 133 376
rect 131 375 132 376
rect 130 375 131 376
rect 129 375 130 376
rect 128 375 129 376
rect 127 375 128 376
rect 126 375 127 376
rect 125 375 126 376
rect 124 375 125 376
rect 123 375 124 376
rect 122 375 123 376
rect 121 375 122 376
rect 120 375 121 376
rect 119 375 120 376
rect 118 375 119 376
rect 117 375 118 376
rect 116 375 117 376
rect 115 375 116 376
rect 114 375 115 376
rect 113 375 114 376
rect 112 375 113 376
rect 111 375 112 376
rect 110 375 111 376
rect 109 375 110 376
rect 108 375 109 376
rect 107 375 108 376
rect 106 375 107 376
rect 105 375 106 376
rect 104 375 105 376
rect 76 375 77 376
rect 75 375 76 376
rect 74 375 75 376
rect 73 375 74 376
rect 72 375 73 376
rect 71 375 72 376
rect 70 375 71 376
rect 69 375 70 376
rect 61 375 62 376
rect 60 375 61 376
rect 59 375 60 376
rect 58 375 59 376
rect 24 375 25 376
rect 23 375 24 376
rect 22 375 23 376
rect 21 375 22 376
rect 20 375 21 376
rect 19 375 20 376
rect 18 375 19 376
rect 17 375 18 376
rect 198 376 199 377
rect 197 376 198 377
rect 196 376 197 377
rect 193 376 194 377
rect 151 376 152 377
rect 150 376 151 377
rect 149 376 150 377
rect 148 376 149 377
rect 147 376 148 377
rect 146 376 147 377
rect 145 376 146 377
rect 144 376 145 377
rect 143 376 144 377
rect 142 376 143 377
rect 141 376 142 377
rect 140 376 141 377
rect 139 376 140 377
rect 138 376 139 377
rect 137 376 138 377
rect 136 376 137 377
rect 135 376 136 377
rect 134 376 135 377
rect 133 376 134 377
rect 132 376 133 377
rect 131 376 132 377
rect 130 376 131 377
rect 129 376 130 377
rect 128 376 129 377
rect 127 376 128 377
rect 126 376 127 377
rect 125 376 126 377
rect 124 376 125 377
rect 123 376 124 377
rect 122 376 123 377
rect 121 376 122 377
rect 120 376 121 377
rect 119 376 120 377
rect 118 376 119 377
rect 117 376 118 377
rect 116 376 117 377
rect 115 376 116 377
rect 114 376 115 377
rect 113 376 114 377
rect 112 376 113 377
rect 111 376 112 377
rect 110 376 111 377
rect 109 376 110 377
rect 108 376 109 377
rect 107 376 108 377
rect 106 376 107 377
rect 105 376 106 377
rect 104 376 105 377
rect 77 376 78 377
rect 76 376 77 377
rect 75 376 76 377
rect 74 376 75 377
rect 73 376 74 377
rect 72 376 73 377
rect 71 376 72 377
rect 70 376 71 377
rect 69 376 70 377
rect 68 376 69 377
rect 63 376 64 377
rect 62 376 63 377
rect 61 376 62 377
rect 60 376 61 377
rect 59 376 60 377
rect 58 376 59 377
rect 57 376 58 377
rect 56 376 57 377
rect 22 376 23 377
rect 21 376 22 377
rect 20 376 21 377
rect 19 376 20 377
rect 18 376 19 377
rect 151 377 152 378
rect 150 377 151 378
rect 149 377 150 378
rect 148 377 149 378
rect 147 377 148 378
rect 146 377 147 378
rect 145 377 146 378
rect 144 377 145 378
rect 143 377 144 378
rect 142 377 143 378
rect 141 377 142 378
rect 140 377 141 378
rect 139 377 140 378
rect 138 377 139 378
rect 137 377 138 378
rect 136 377 137 378
rect 135 377 136 378
rect 134 377 135 378
rect 133 377 134 378
rect 132 377 133 378
rect 131 377 132 378
rect 130 377 131 378
rect 129 377 130 378
rect 128 377 129 378
rect 127 377 128 378
rect 126 377 127 378
rect 125 377 126 378
rect 124 377 125 378
rect 123 377 124 378
rect 122 377 123 378
rect 121 377 122 378
rect 120 377 121 378
rect 119 377 120 378
rect 118 377 119 378
rect 117 377 118 378
rect 116 377 117 378
rect 115 377 116 378
rect 114 377 115 378
rect 113 377 114 378
rect 112 377 113 378
rect 111 377 112 378
rect 110 377 111 378
rect 109 377 110 378
rect 108 377 109 378
rect 107 377 108 378
rect 106 377 107 378
rect 105 377 106 378
rect 104 377 105 378
rect 78 377 79 378
rect 77 377 78 378
rect 76 377 77 378
rect 75 377 76 378
rect 74 377 75 378
rect 73 377 74 378
rect 72 377 73 378
rect 71 377 72 378
rect 70 377 71 378
rect 69 377 70 378
rect 68 377 69 378
rect 67 377 68 378
rect 64 377 65 378
rect 63 377 64 378
rect 62 377 63 378
rect 61 377 62 378
rect 60 377 61 378
rect 59 377 60 378
rect 58 377 59 378
rect 57 377 58 378
rect 56 377 57 378
rect 55 377 56 378
rect 151 378 152 379
rect 150 378 151 379
rect 149 378 150 379
rect 148 378 149 379
rect 147 378 148 379
rect 146 378 147 379
rect 145 378 146 379
rect 144 378 145 379
rect 143 378 144 379
rect 142 378 143 379
rect 141 378 142 379
rect 140 378 141 379
rect 139 378 140 379
rect 138 378 139 379
rect 137 378 138 379
rect 136 378 137 379
rect 135 378 136 379
rect 134 378 135 379
rect 133 378 134 379
rect 132 378 133 379
rect 131 378 132 379
rect 130 378 131 379
rect 129 378 130 379
rect 128 378 129 379
rect 127 378 128 379
rect 126 378 127 379
rect 125 378 126 379
rect 124 378 125 379
rect 123 378 124 379
rect 122 378 123 379
rect 121 378 122 379
rect 120 378 121 379
rect 119 378 120 379
rect 118 378 119 379
rect 117 378 118 379
rect 116 378 117 379
rect 115 378 116 379
rect 114 378 115 379
rect 113 378 114 379
rect 112 378 113 379
rect 111 378 112 379
rect 110 378 111 379
rect 109 378 110 379
rect 108 378 109 379
rect 107 378 108 379
rect 106 378 107 379
rect 105 378 106 379
rect 104 378 105 379
rect 79 378 80 379
rect 78 378 79 379
rect 77 378 78 379
rect 76 378 77 379
rect 75 378 76 379
rect 74 378 75 379
rect 73 378 74 379
rect 72 378 73 379
rect 71 378 72 379
rect 70 378 71 379
rect 69 378 70 379
rect 68 378 69 379
rect 67 378 68 379
rect 66 378 67 379
rect 65 378 66 379
rect 64 378 65 379
rect 63 378 64 379
rect 62 378 63 379
rect 61 378 62 379
rect 60 378 61 379
rect 59 378 60 379
rect 58 378 59 379
rect 57 378 58 379
rect 56 378 57 379
rect 55 378 56 379
rect 54 378 55 379
rect 151 379 152 380
rect 150 379 151 380
rect 149 379 150 380
rect 148 379 149 380
rect 147 379 148 380
rect 146 379 147 380
rect 145 379 146 380
rect 144 379 145 380
rect 143 379 144 380
rect 142 379 143 380
rect 141 379 142 380
rect 140 379 141 380
rect 139 379 140 380
rect 138 379 139 380
rect 137 379 138 380
rect 136 379 137 380
rect 135 379 136 380
rect 134 379 135 380
rect 133 379 134 380
rect 132 379 133 380
rect 131 379 132 380
rect 130 379 131 380
rect 129 379 130 380
rect 128 379 129 380
rect 127 379 128 380
rect 126 379 127 380
rect 125 379 126 380
rect 124 379 125 380
rect 123 379 124 380
rect 122 379 123 380
rect 121 379 122 380
rect 120 379 121 380
rect 119 379 120 380
rect 118 379 119 380
rect 117 379 118 380
rect 116 379 117 380
rect 115 379 116 380
rect 114 379 115 380
rect 113 379 114 380
rect 112 379 113 380
rect 111 379 112 380
rect 110 379 111 380
rect 109 379 110 380
rect 108 379 109 380
rect 107 379 108 380
rect 106 379 107 380
rect 105 379 106 380
rect 104 379 105 380
rect 80 379 81 380
rect 79 379 80 380
rect 78 379 79 380
rect 77 379 78 380
rect 76 379 77 380
rect 75 379 76 380
rect 74 379 75 380
rect 73 379 74 380
rect 72 379 73 380
rect 71 379 72 380
rect 70 379 71 380
rect 69 379 70 380
rect 68 379 69 380
rect 67 379 68 380
rect 66 379 67 380
rect 65 379 66 380
rect 64 379 65 380
rect 63 379 64 380
rect 62 379 63 380
rect 61 379 62 380
rect 60 379 61 380
rect 59 379 60 380
rect 58 379 59 380
rect 57 379 58 380
rect 56 379 57 380
rect 55 379 56 380
rect 54 379 55 380
rect 31 379 32 380
rect 30 379 31 380
rect 29 379 30 380
rect 28 379 29 380
rect 27 379 28 380
rect 26 379 27 380
rect 25 379 26 380
rect 24 379 25 380
rect 23 379 24 380
rect 22 379 23 380
rect 21 379 22 380
rect 20 379 21 380
rect 19 379 20 380
rect 18 379 19 380
rect 17 379 18 380
rect 16 379 17 380
rect 114 380 115 381
rect 113 380 114 381
rect 112 380 113 381
rect 111 380 112 381
rect 110 380 111 381
rect 109 380 110 381
rect 108 380 109 381
rect 107 380 108 381
rect 106 380 107 381
rect 105 380 106 381
rect 104 380 105 381
rect 80 380 81 381
rect 79 380 80 381
rect 78 380 79 381
rect 77 380 78 381
rect 76 380 77 381
rect 75 380 76 381
rect 69 380 70 381
rect 68 380 69 381
rect 67 380 68 381
rect 66 380 67 381
rect 65 380 66 381
rect 64 380 65 381
rect 63 380 64 381
rect 62 380 63 381
rect 61 380 62 381
rect 60 380 61 381
rect 59 380 60 381
rect 58 380 59 381
rect 57 380 58 381
rect 56 380 57 381
rect 55 380 56 381
rect 54 380 55 381
rect 31 380 32 381
rect 30 380 31 381
rect 29 380 30 381
rect 28 380 29 381
rect 27 380 28 381
rect 26 380 27 381
rect 25 380 26 381
rect 24 380 25 381
rect 23 380 24 381
rect 22 380 23 381
rect 21 380 22 381
rect 20 380 21 381
rect 19 380 20 381
rect 18 380 19 381
rect 17 380 18 381
rect 16 380 17 381
rect 199 381 200 382
rect 198 381 199 382
rect 197 381 198 382
rect 196 381 197 382
rect 195 381 196 382
rect 194 381 195 382
rect 193 381 194 382
rect 192 381 193 382
rect 191 381 192 382
rect 114 381 115 382
rect 113 381 114 382
rect 112 381 113 382
rect 111 381 112 382
rect 110 381 111 382
rect 109 381 110 382
rect 108 381 109 382
rect 107 381 108 382
rect 106 381 107 382
rect 105 381 106 382
rect 104 381 105 382
rect 80 381 81 382
rect 79 381 80 382
rect 78 381 79 382
rect 77 381 78 382
rect 76 381 77 382
rect 68 381 69 382
rect 67 381 68 382
rect 66 381 67 382
rect 65 381 66 382
rect 64 381 65 382
rect 63 381 64 382
rect 57 381 58 382
rect 56 381 57 382
rect 55 381 56 382
rect 54 381 55 382
rect 53 381 54 382
rect 31 381 32 382
rect 30 381 31 382
rect 29 381 30 382
rect 28 381 29 382
rect 27 381 28 382
rect 26 381 27 382
rect 25 381 26 382
rect 24 381 25 382
rect 23 381 24 382
rect 22 381 23 382
rect 21 381 22 382
rect 20 381 21 382
rect 19 381 20 382
rect 18 381 19 382
rect 17 381 18 382
rect 198 382 199 383
rect 197 382 198 383
rect 196 382 197 383
rect 195 382 196 383
rect 194 382 195 383
rect 193 382 194 383
rect 192 382 193 383
rect 191 382 192 383
rect 114 382 115 383
rect 113 382 114 383
rect 112 382 113 383
rect 111 382 112 383
rect 110 382 111 383
rect 109 382 110 383
rect 108 382 109 383
rect 107 382 108 383
rect 106 382 107 383
rect 105 382 106 383
rect 104 382 105 383
rect 80 382 81 383
rect 79 382 80 383
rect 78 382 79 383
rect 77 382 78 383
rect 67 382 68 383
rect 66 382 67 383
rect 65 382 66 383
rect 64 382 65 383
rect 57 382 58 383
rect 56 382 57 383
rect 55 382 56 383
rect 54 382 55 383
rect 53 382 54 383
rect 31 382 32 383
rect 30 382 31 383
rect 29 382 30 383
rect 28 382 29 383
rect 27 382 28 383
rect 26 382 27 383
rect 195 383 196 384
rect 194 383 195 384
rect 191 383 192 384
rect 114 383 115 384
rect 113 383 114 384
rect 112 383 113 384
rect 111 383 112 384
rect 110 383 111 384
rect 109 383 110 384
rect 108 383 109 384
rect 107 383 108 384
rect 106 383 107 384
rect 105 383 106 384
rect 104 383 105 384
rect 80 383 81 384
rect 79 383 80 384
rect 78 383 79 384
rect 77 383 78 384
rect 67 383 68 384
rect 66 383 67 384
rect 65 383 66 384
rect 64 383 65 384
rect 57 383 58 384
rect 56 383 57 384
rect 55 383 56 384
rect 54 383 55 384
rect 53 383 54 384
rect 30 383 31 384
rect 29 383 30 384
rect 28 383 29 384
rect 27 383 28 384
rect 26 383 27 384
rect 25 383 26 384
rect 24 383 25 384
rect 196 384 197 385
rect 195 384 196 385
rect 194 384 195 385
rect 192 384 193 385
rect 191 384 192 385
rect 114 384 115 385
rect 113 384 114 385
rect 112 384 113 385
rect 111 384 112 385
rect 110 384 111 385
rect 109 384 110 385
rect 108 384 109 385
rect 107 384 108 385
rect 106 384 107 385
rect 105 384 106 385
rect 104 384 105 385
rect 80 384 81 385
rect 79 384 80 385
rect 78 384 79 385
rect 77 384 78 385
rect 67 384 68 385
rect 66 384 67 385
rect 65 384 66 385
rect 64 384 65 385
rect 57 384 58 385
rect 56 384 57 385
rect 55 384 56 385
rect 54 384 55 385
rect 53 384 54 385
rect 28 384 29 385
rect 27 384 28 385
rect 26 384 27 385
rect 25 384 26 385
rect 24 384 25 385
rect 23 384 24 385
rect 22 384 23 385
rect 198 385 199 386
rect 197 385 198 386
rect 196 385 197 386
rect 195 385 196 386
rect 194 385 195 386
rect 193 385 194 386
rect 192 385 193 386
rect 191 385 192 386
rect 114 385 115 386
rect 113 385 114 386
rect 112 385 113 386
rect 111 385 112 386
rect 110 385 111 386
rect 109 385 110 386
rect 108 385 109 386
rect 107 385 108 386
rect 106 385 107 386
rect 105 385 106 386
rect 104 385 105 386
rect 80 385 81 386
rect 79 385 80 386
rect 78 385 79 386
rect 77 385 78 386
rect 68 385 69 386
rect 67 385 68 386
rect 66 385 67 386
rect 65 385 66 386
rect 64 385 65 386
rect 63 385 64 386
rect 57 385 58 386
rect 56 385 57 386
rect 55 385 56 386
rect 54 385 55 386
rect 53 385 54 386
rect 26 385 27 386
rect 25 385 26 386
rect 24 385 25 386
rect 23 385 24 386
rect 22 385 23 386
rect 21 385 22 386
rect 20 385 21 386
rect 198 386 199 387
rect 197 386 198 387
rect 196 386 197 387
rect 194 386 195 387
rect 193 386 194 387
rect 192 386 193 387
rect 191 386 192 387
rect 114 386 115 387
rect 113 386 114 387
rect 112 386 113 387
rect 111 386 112 387
rect 110 386 111 387
rect 109 386 110 387
rect 108 386 109 387
rect 107 386 108 387
rect 106 386 107 387
rect 105 386 106 387
rect 104 386 105 387
rect 80 386 81 387
rect 79 386 80 387
rect 78 386 79 387
rect 77 386 78 387
rect 76 386 77 387
rect 69 386 70 387
rect 68 386 69 387
rect 67 386 68 387
rect 66 386 67 387
rect 65 386 66 387
rect 64 386 65 387
rect 63 386 64 387
rect 62 386 63 387
rect 58 386 59 387
rect 57 386 58 387
rect 56 386 57 387
rect 55 386 56 387
rect 54 386 55 387
rect 53 386 54 387
rect 24 386 25 387
rect 23 386 24 387
rect 22 386 23 387
rect 21 386 22 387
rect 20 386 21 387
rect 19 386 20 387
rect 18 386 19 387
rect 198 387 199 388
rect 196 387 197 388
rect 172 387 173 388
rect 171 387 172 388
rect 170 387 171 388
rect 169 387 170 388
rect 168 387 169 388
rect 167 387 168 388
rect 114 387 115 388
rect 113 387 114 388
rect 112 387 113 388
rect 111 387 112 388
rect 110 387 111 388
rect 109 387 110 388
rect 108 387 109 388
rect 107 387 108 388
rect 106 387 107 388
rect 105 387 106 388
rect 104 387 105 388
rect 80 387 81 388
rect 79 387 80 388
rect 78 387 79 388
rect 77 387 78 388
rect 76 387 77 388
rect 75 387 76 388
rect 74 387 75 388
rect 73 387 74 388
rect 72 387 73 388
rect 71 387 72 388
rect 70 387 71 388
rect 69 387 70 388
rect 68 387 69 388
rect 67 387 68 388
rect 66 387 67 388
rect 65 387 66 388
rect 64 387 65 388
rect 63 387 64 388
rect 62 387 63 388
rect 61 387 62 388
rect 60 387 61 388
rect 59 387 60 388
rect 58 387 59 388
rect 57 387 58 388
rect 56 387 57 388
rect 55 387 56 388
rect 54 387 55 388
rect 21 387 22 388
rect 20 387 21 388
rect 19 387 20 388
rect 18 387 19 388
rect 17 387 18 388
rect 198 388 199 389
rect 197 388 198 389
rect 196 388 197 389
rect 195 388 196 389
rect 194 388 195 389
rect 173 388 174 389
rect 172 388 173 389
rect 171 388 172 389
rect 170 388 171 389
rect 169 388 170 389
rect 168 388 169 389
rect 167 388 168 389
rect 166 388 167 389
rect 130 388 131 389
rect 114 388 115 389
rect 113 388 114 389
rect 112 388 113 389
rect 111 388 112 389
rect 110 388 111 389
rect 109 388 110 389
rect 108 388 109 389
rect 107 388 108 389
rect 106 388 107 389
rect 105 388 106 389
rect 104 388 105 389
rect 79 388 80 389
rect 78 388 79 389
rect 77 388 78 389
rect 76 388 77 389
rect 75 388 76 389
rect 74 388 75 389
rect 73 388 74 389
rect 72 388 73 389
rect 71 388 72 389
rect 70 388 71 389
rect 69 388 70 389
rect 68 388 69 389
rect 67 388 68 389
rect 66 388 67 389
rect 65 388 66 389
rect 64 388 65 389
rect 63 388 64 389
rect 62 388 63 389
rect 61 388 62 389
rect 60 388 61 389
rect 59 388 60 389
rect 58 388 59 389
rect 57 388 58 389
rect 56 388 57 389
rect 55 388 56 389
rect 54 388 55 389
rect 31 388 32 389
rect 30 388 31 389
rect 29 388 30 389
rect 28 388 29 389
rect 27 388 28 389
rect 26 388 27 389
rect 25 388 26 389
rect 24 388 25 389
rect 23 388 24 389
rect 22 388 23 389
rect 21 388 22 389
rect 20 388 21 389
rect 19 388 20 389
rect 18 388 19 389
rect 17 388 18 389
rect 16 388 17 389
rect 198 389 199 390
rect 197 389 198 390
rect 196 389 197 390
rect 195 389 196 390
rect 194 389 195 390
rect 193 389 194 390
rect 174 389 175 390
rect 173 389 174 390
rect 172 389 173 390
rect 171 389 172 390
rect 170 389 171 390
rect 169 389 170 390
rect 168 389 169 390
rect 167 389 168 390
rect 166 389 167 390
rect 165 389 166 390
rect 131 389 132 390
rect 130 389 131 390
rect 129 389 130 390
rect 114 389 115 390
rect 113 389 114 390
rect 112 389 113 390
rect 111 389 112 390
rect 110 389 111 390
rect 109 389 110 390
rect 108 389 109 390
rect 107 389 108 390
rect 106 389 107 390
rect 105 389 106 390
rect 104 389 105 390
rect 79 389 80 390
rect 78 389 79 390
rect 77 389 78 390
rect 76 389 77 390
rect 75 389 76 390
rect 74 389 75 390
rect 73 389 74 390
rect 72 389 73 390
rect 71 389 72 390
rect 70 389 71 390
rect 69 389 70 390
rect 68 389 69 390
rect 67 389 68 390
rect 64 389 65 390
rect 63 389 64 390
rect 62 389 63 390
rect 61 389 62 390
rect 60 389 61 390
rect 59 389 60 390
rect 58 389 59 390
rect 57 389 58 390
rect 56 389 57 390
rect 55 389 56 390
rect 31 389 32 390
rect 30 389 31 390
rect 29 389 30 390
rect 28 389 29 390
rect 27 389 28 390
rect 26 389 27 390
rect 25 389 26 390
rect 24 389 25 390
rect 23 389 24 390
rect 22 389 23 390
rect 21 389 22 390
rect 20 389 21 390
rect 19 389 20 390
rect 18 389 19 390
rect 17 389 18 390
rect 16 389 17 390
rect 199 390 200 391
rect 198 390 199 391
rect 196 390 197 391
rect 194 390 195 391
rect 193 390 194 391
rect 185 390 186 391
rect 184 390 185 391
rect 183 390 184 391
rect 182 390 183 391
rect 181 390 182 391
rect 180 390 181 391
rect 179 390 180 391
rect 178 390 179 391
rect 175 390 176 391
rect 174 390 175 391
rect 173 390 174 391
rect 172 390 173 391
rect 171 390 172 391
rect 168 390 169 391
rect 167 390 168 391
rect 166 390 167 391
rect 165 390 166 391
rect 132 390 133 391
rect 131 390 132 391
rect 130 390 131 391
rect 129 390 130 391
rect 114 390 115 391
rect 113 390 114 391
rect 112 390 113 391
rect 111 390 112 391
rect 110 390 111 391
rect 109 390 110 391
rect 108 390 109 391
rect 107 390 108 391
rect 106 390 107 391
rect 105 390 106 391
rect 104 390 105 391
rect 78 390 79 391
rect 77 390 78 391
rect 76 390 77 391
rect 75 390 76 391
rect 74 390 75 391
rect 73 390 74 391
rect 72 390 73 391
rect 71 390 72 391
rect 70 390 71 391
rect 69 390 70 391
rect 68 390 69 391
rect 67 390 68 391
rect 63 390 64 391
rect 62 390 63 391
rect 61 390 62 391
rect 60 390 61 391
rect 59 390 60 391
rect 58 390 59 391
rect 57 390 58 391
rect 56 390 57 391
rect 31 390 32 391
rect 30 390 31 391
rect 29 390 30 391
rect 28 390 29 391
rect 27 390 28 391
rect 26 390 27 391
rect 25 390 26 391
rect 24 390 25 391
rect 23 390 24 391
rect 22 390 23 391
rect 21 390 22 391
rect 20 390 21 391
rect 19 390 20 391
rect 18 390 19 391
rect 17 390 18 391
rect 199 391 200 392
rect 198 391 199 392
rect 196 391 197 392
rect 194 391 195 392
rect 193 391 194 392
rect 185 391 186 392
rect 184 391 185 392
rect 183 391 184 392
rect 182 391 183 392
rect 181 391 182 392
rect 180 391 181 392
rect 179 391 180 392
rect 178 391 179 392
rect 175 391 176 392
rect 174 391 175 392
rect 173 391 174 392
rect 172 391 173 392
rect 167 391 168 392
rect 166 391 167 392
rect 165 391 166 392
rect 133 391 134 392
rect 132 391 133 392
rect 131 391 132 392
rect 130 391 131 392
rect 129 391 130 392
rect 114 391 115 392
rect 113 391 114 392
rect 112 391 113 392
rect 111 391 112 392
rect 110 391 111 392
rect 109 391 110 392
rect 108 391 109 392
rect 107 391 108 392
rect 106 391 107 392
rect 105 391 106 392
rect 104 391 105 392
rect 77 391 78 392
rect 76 391 77 392
rect 75 391 76 392
rect 74 391 75 392
rect 73 391 74 392
rect 72 391 73 392
rect 71 391 72 392
rect 70 391 71 392
rect 69 391 70 392
rect 68 391 69 392
rect 62 391 63 392
rect 61 391 62 392
rect 60 391 61 392
rect 59 391 60 392
rect 58 391 59 392
rect 31 391 32 392
rect 30 391 31 392
rect 29 391 30 392
rect 28 391 29 392
rect 27 391 28 392
rect 26 391 27 392
rect 199 392 200 393
rect 198 392 199 393
rect 196 392 197 393
rect 195 392 196 393
rect 194 392 195 393
rect 193 392 194 393
rect 185 392 186 393
rect 184 392 185 393
rect 183 392 184 393
rect 182 392 183 393
rect 181 392 182 393
rect 180 392 181 393
rect 179 392 180 393
rect 178 392 179 393
rect 175 392 176 393
rect 174 392 175 393
rect 173 392 174 393
rect 167 392 168 393
rect 166 392 167 393
rect 165 392 166 393
rect 164 392 165 393
rect 133 392 134 393
rect 132 392 133 393
rect 131 392 132 393
rect 130 392 131 393
rect 129 392 130 393
rect 114 392 115 393
rect 113 392 114 393
rect 112 392 113 393
rect 111 392 112 393
rect 110 392 111 393
rect 109 392 110 393
rect 108 392 109 393
rect 107 392 108 393
rect 106 392 107 393
rect 105 392 106 393
rect 104 392 105 393
rect 75 392 76 393
rect 74 392 75 393
rect 73 392 74 393
rect 72 392 73 393
rect 71 392 72 393
rect 70 392 71 393
rect 29 392 30 393
rect 28 392 29 393
rect 27 392 28 393
rect 26 392 27 393
rect 25 392 26 393
rect 24 392 25 393
rect 198 393 199 394
rect 196 393 197 394
rect 195 393 196 394
rect 194 393 195 394
rect 185 393 186 394
rect 184 393 185 394
rect 183 393 184 394
rect 182 393 183 394
rect 181 393 182 394
rect 180 393 181 394
rect 179 393 180 394
rect 178 393 179 394
rect 175 393 176 394
rect 174 393 175 394
rect 173 393 174 394
rect 166 393 167 394
rect 165 393 166 394
rect 164 393 165 394
rect 134 393 135 394
rect 133 393 134 394
rect 132 393 133 394
rect 131 393 132 394
rect 130 393 131 394
rect 129 393 130 394
rect 114 393 115 394
rect 113 393 114 394
rect 112 393 113 394
rect 111 393 112 394
rect 110 393 111 394
rect 109 393 110 394
rect 108 393 109 394
rect 107 393 108 394
rect 106 393 107 394
rect 105 393 106 394
rect 104 393 105 394
rect 27 393 28 394
rect 26 393 27 394
rect 25 393 26 394
rect 24 393 25 394
rect 23 393 24 394
rect 22 393 23 394
rect 198 394 199 395
rect 195 394 196 395
rect 185 394 186 395
rect 184 394 185 395
rect 183 394 184 395
rect 182 394 183 395
rect 175 394 176 395
rect 174 394 175 395
rect 173 394 174 395
rect 167 394 168 395
rect 166 394 167 395
rect 165 394 166 395
rect 164 394 165 395
rect 135 394 136 395
rect 134 394 135 395
rect 133 394 134 395
rect 132 394 133 395
rect 131 394 132 395
rect 130 394 131 395
rect 129 394 130 395
rect 114 394 115 395
rect 113 394 114 395
rect 112 394 113 395
rect 111 394 112 395
rect 110 394 111 395
rect 109 394 110 395
rect 108 394 109 395
rect 107 394 108 395
rect 106 394 107 395
rect 105 394 106 395
rect 104 394 105 395
rect 25 394 26 395
rect 24 394 25 395
rect 23 394 24 395
rect 22 394 23 395
rect 21 394 22 395
rect 20 394 21 395
rect 19 394 20 395
rect 199 395 200 396
rect 198 395 199 396
rect 196 395 197 396
rect 195 395 196 396
rect 194 395 195 396
rect 193 395 194 396
rect 185 395 186 396
rect 184 395 185 396
rect 183 395 184 396
rect 182 395 183 396
rect 175 395 176 396
rect 174 395 175 396
rect 173 395 174 396
rect 172 395 173 396
rect 167 395 168 396
rect 166 395 167 396
rect 165 395 166 396
rect 136 395 137 396
rect 135 395 136 396
rect 134 395 135 396
rect 133 395 134 396
rect 132 395 133 396
rect 131 395 132 396
rect 130 395 131 396
rect 129 395 130 396
rect 114 395 115 396
rect 113 395 114 396
rect 112 395 113 396
rect 111 395 112 396
rect 110 395 111 396
rect 109 395 110 396
rect 108 395 109 396
rect 107 395 108 396
rect 106 395 107 396
rect 105 395 106 396
rect 104 395 105 396
rect 23 395 24 396
rect 22 395 23 396
rect 21 395 22 396
rect 20 395 21 396
rect 19 395 20 396
rect 18 395 19 396
rect 17 395 18 396
rect 199 396 200 397
rect 198 396 199 397
rect 196 396 197 397
rect 195 396 196 397
rect 194 396 195 397
rect 193 396 194 397
rect 185 396 186 397
rect 184 396 185 397
rect 183 396 184 397
rect 182 396 183 397
rect 175 396 176 397
rect 174 396 175 397
rect 173 396 174 397
rect 172 396 173 397
rect 171 396 172 397
rect 168 396 169 397
rect 167 396 168 397
rect 166 396 167 397
rect 165 396 166 397
rect 137 396 138 397
rect 136 396 137 397
rect 135 396 136 397
rect 134 396 135 397
rect 133 396 134 397
rect 132 396 133 397
rect 131 396 132 397
rect 130 396 131 397
rect 129 396 130 397
rect 114 396 115 397
rect 113 396 114 397
rect 112 396 113 397
rect 111 396 112 397
rect 110 396 111 397
rect 109 396 110 397
rect 108 396 109 397
rect 107 396 108 397
rect 106 396 107 397
rect 105 396 106 397
rect 104 396 105 397
rect 88 396 89 397
rect 87 396 88 397
rect 86 396 87 397
rect 55 396 56 397
rect 54 396 55 397
rect 53 396 54 397
rect 21 396 22 397
rect 20 396 21 397
rect 19 396 20 397
rect 18 396 19 397
rect 17 396 18 397
rect 16 396 17 397
rect 199 397 200 398
rect 198 397 199 398
rect 197 397 198 398
rect 196 397 197 398
rect 194 397 195 398
rect 193 397 194 398
rect 185 397 186 398
rect 184 397 185 398
rect 183 397 184 398
rect 182 397 183 398
rect 174 397 175 398
rect 173 397 174 398
rect 172 397 173 398
rect 171 397 172 398
rect 170 397 171 398
rect 169 397 170 398
rect 168 397 169 398
rect 167 397 168 398
rect 166 397 167 398
rect 165 397 166 398
rect 138 397 139 398
rect 137 397 138 398
rect 136 397 137 398
rect 135 397 136 398
rect 134 397 135 398
rect 133 397 134 398
rect 132 397 133 398
rect 131 397 132 398
rect 130 397 131 398
rect 129 397 130 398
rect 114 397 115 398
rect 113 397 114 398
rect 112 397 113 398
rect 111 397 112 398
rect 110 397 111 398
rect 109 397 110 398
rect 108 397 109 398
rect 107 397 108 398
rect 106 397 107 398
rect 105 397 106 398
rect 104 397 105 398
rect 88 397 89 398
rect 87 397 88 398
rect 86 397 87 398
rect 85 397 86 398
rect 84 397 85 398
rect 57 397 58 398
rect 56 397 57 398
rect 55 397 56 398
rect 54 397 55 398
rect 53 397 54 398
rect 19 397 20 398
rect 18 397 19 398
rect 17 397 18 398
rect 16 397 17 398
rect 198 398 199 399
rect 197 398 198 399
rect 196 398 197 399
rect 193 398 194 399
rect 185 398 186 399
rect 184 398 185 399
rect 183 398 184 399
rect 182 398 183 399
rect 174 398 175 399
rect 173 398 174 399
rect 172 398 173 399
rect 171 398 172 399
rect 170 398 171 399
rect 169 398 170 399
rect 168 398 169 399
rect 167 398 168 399
rect 166 398 167 399
rect 138 398 139 399
rect 137 398 138 399
rect 136 398 137 399
rect 135 398 136 399
rect 134 398 135 399
rect 133 398 134 399
rect 132 398 133 399
rect 131 398 132 399
rect 130 398 131 399
rect 129 398 130 399
rect 114 398 115 399
rect 113 398 114 399
rect 112 398 113 399
rect 111 398 112 399
rect 110 398 111 399
rect 109 398 110 399
rect 108 398 109 399
rect 107 398 108 399
rect 106 398 107 399
rect 105 398 106 399
rect 104 398 105 399
rect 88 398 89 399
rect 87 398 88 399
rect 86 398 87 399
rect 85 398 86 399
rect 84 398 85 399
rect 83 398 84 399
rect 82 398 83 399
rect 81 398 82 399
rect 60 398 61 399
rect 59 398 60 399
rect 58 398 59 399
rect 57 398 58 399
rect 56 398 57 399
rect 55 398 56 399
rect 54 398 55 399
rect 53 398 54 399
rect 17 398 18 399
rect 197 399 198 400
rect 196 399 197 400
rect 195 399 196 400
rect 185 399 186 400
rect 184 399 185 400
rect 183 399 184 400
rect 182 399 183 400
rect 173 399 174 400
rect 172 399 173 400
rect 171 399 172 400
rect 170 399 171 400
rect 169 399 170 400
rect 168 399 169 400
rect 167 399 168 400
rect 166 399 167 400
rect 139 399 140 400
rect 138 399 139 400
rect 137 399 138 400
rect 136 399 137 400
rect 135 399 136 400
rect 134 399 135 400
rect 133 399 134 400
rect 132 399 133 400
rect 131 399 132 400
rect 130 399 131 400
rect 129 399 130 400
rect 114 399 115 400
rect 113 399 114 400
rect 112 399 113 400
rect 111 399 112 400
rect 110 399 111 400
rect 109 399 110 400
rect 108 399 109 400
rect 107 399 108 400
rect 106 399 107 400
rect 105 399 106 400
rect 104 399 105 400
rect 87 399 88 400
rect 86 399 87 400
rect 85 399 86 400
rect 84 399 85 400
rect 83 399 84 400
rect 82 399 83 400
rect 81 399 82 400
rect 80 399 81 400
rect 79 399 80 400
rect 78 399 79 400
rect 77 399 78 400
rect 76 399 77 400
rect 65 399 66 400
rect 64 399 65 400
rect 63 399 64 400
rect 62 399 63 400
rect 61 399 62 400
rect 60 399 61 400
rect 59 399 60 400
rect 58 399 59 400
rect 57 399 58 400
rect 56 399 57 400
rect 55 399 56 400
rect 54 399 55 400
rect 198 400 199 401
rect 197 400 198 401
rect 196 400 197 401
rect 195 400 196 401
rect 194 400 195 401
rect 193 400 194 401
rect 185 400 186 401
rect 184 400 185 401
rect 183 400 184 401
rect 182 400 183 401
rect 173 400 174 401
rect 172 400 173 401
rect 171 400 172 401
rect 170 400 171 401
rect 169 400 170 401
rect 168 400 169 401
rect 167 400 168 401
rect 166 400 167 401
rect 140 400 141 401
rect 139 400 140 401
rect 138 400 139 401
rect 137 400 138 401
rect 136 400 137 401
rect 135 400 136 401
rect 134 400 135 401
rect 133 400 134 401
rect 132 400 133 401
rect 131 400 132 401
rect 130 400 131 401
rect 129 400 130 401
rect 114 400 115 401
rect 113 400 114 401
rect 112 400 113 401
rect 111 400 112 401
rect 110 400 111 401
rect 109 400 110 401
rect 108 400 109 401
rect 107 400 108 401
rect 106 400 107 401
rect 105 400 106 401
rect 104 400 105 401
rect 86 400 87 401
rect 85 400 86 401
rect 84 400 85 401
rect 83 400 84 401
rect 82 400 83 401
rect 81 400 82 401
rect 80 400 81 401
rect 79 400 80 401
rect 78 400 79 401
rect 77 400 78 401
rect 76 400 77 401
rect 75 400 76 401
rect 74 400 75 401
rect 73 400 74 401
rect 72 400 73 401
rect 71 400 72 401
rect 70 400 71 401
rect 69 400 70 401
rect 68 400 69 401
rect 67 400 68 401
rect 66 400 67 401
rect 65 400 66 401
rect 64 400 65 401
rect 63 400 64 401
rect 62 400 63 401
rect 61 400 62 401
rect 60 400 61 401
rect 59 400 60 401
rect 58 400 59 401
rect 57 400 58 401
rect 56 400 57 401
rect 55 400 56 401
rect 199 401 200 402
rect 198 401 199 402
rect 197 401 198 402
rect 196 401 197 402
rect 195 401 196 402
rect 194 401 195 402
rect 193 401 194 402
rect 185 401 186 402
rect 184 401 185 402
rect 183 401 184 402
rect 182 401 183 402
rect 173 401 174 402
rect 172 401 173 402
rect 171 401 172 402
rect 169 401 170 402
rect 168 401 169 402
rect 167 401 168 402
rect 166 401 167 402
rect 141 401 142 402
rect 140 401 141 402
rect 139 401 140 402
rect 138 401 139 402
rect 137 401 138 402
rect 136 401 137 402
rect 135 401 136 402
rect 134 401 135 402
rect 133 401 134 402
rect 132 401 133 402
rect 131 401 132 402
rect 130 401 131 402
rect 129 401 130 402
rect 114 401 115 402
rect 113 401 114 402
rect 112 401 113 402
rect 111 401 112 402
rect 110 401 111 402
rect 109 401 110 402
rect 108 401 109 402
rect 107 401 108 402
rect 106 401 107 402
rect 105 401 106 402
rect 104 401 105 402
rect 84 401 85 402
rect 83 401 84 402
rect 82 401 83 402
rect 81 401 82 402
rect 80 401 81 402
rect 79 401 80 402
rect 78 401 79 402
rect 77 401 78 402
rect 76 401 77 402
rect 75 401 76 402
rect 74 401 75 402
rect 73 401 74 402
rect 72 401 73 402
rect 71 401 72 402
rect 70 401 71 402
rect 69 401 70 402
rect 68 401 69 402
rect 67 401 68 402
rect 66 401 67 402
rect 65 401 66 402
rect 64 401 65 402
rect 63 401 64 402
rect 62 401 63 402
rect 61 401 62 402
rect 60 401 61 402
rect 59 401 60 402
rect 58 401 59 402
rect 57 401 58 402
rect 199 402 200 403
rect 198 402 199 403
rect 196 402 197 403
rect 194 402 195 403
rect 193 402 194 403
rect 185 402 186 403
rect 184 402 185 403
rect 183 402 184 403
rect 182 402 183 403
rect 173 402 174 403
rect 172 402 173 403
rect 171 402 172 403
rect 169 402 170 403
rect 168 402 169 403
rect 167 402 168 403
rect 166 402 167 403
rect 142 402 143 403
rect 141 402 142 403
rect 140 402 141 403
rect 139 402 140 403
rect 138 402 139 403
rect 137 402 138 403
rect 136 402 137 403
rect 135 402 136 403
rect 134 402 135 403
rect 133 402 134 403
rect 132 402 133 403
rect 131 402 132 403
rect 130 402 131 403
rect 129 402 130 403
rect 114 402 115 403
rect 113 402 114 403
rect 112 402 113 403
rect 111 402 112 403
rect 110 402 111 403
rect 109 402 110 403
rect 108 402 109 403
rect 107 402 108 403
rect 106 402 107 403
rect 105 402 106 403
rect 104 402 105 403
rect 82 402 83 403
rect 81 402 82 403
rect 80 402 81 403
rect 79 402 80 403
rect 78 402 79 403
rect 77 402 78 403
rect 76 402 77 403
rect 75 402 76 403
rect 74 402 75 403
rect 73 402 74 403
rect 72 402 73 403
rect 71 402 72 403
rect 70 402 71 403
rect 69 402 70 403
rect 68 402 69 403
rect 67 402 68 403
rect 66 402 67 403
rect 65 402 66 403
rect 64 402 65 403
rect 63 402 64 403
rect 62 402 63 403
rect 61 402 62 403
rect 60 402 61 403
rect 59 402 60 403
rect 199 403 200 404
rect 198 403 199 404
rect 196 403 197 404
rect 195 403 196 404
rect 194 403 195 404
rect 193 403 194 404
rect 185 403 186 404
rect 184 403 185 404
rect 183 403 184 404
rect 182 403 183 404
rect 173 403 174 404
rect 172 403 173 404
rect 171 403 172 404
rect 169 403 170 404
rect 168 403 169 404
rect 167 403 168 404
rect 166 403 167 404
rect 142 403 143 404
rect 141 403 142 404
rect 140 403 141 404
rect 139 403 140 404
rect 138 403 139 404
rect 137 403 138 404
rect 136 403 137 404
rect 135 403 136 404
rect 134 403 135 404
rect 133 403 134 404
rect 132 403 133 404
rect 131 403 132 404
rect 130 403 131 404
rect 129 403 130 404
rect 114 403 115 404
rect 113 403 114 404
rect 112 403 113 404
rect 111 403 112 404
rect 110 403 111 404
rect 109 403 110 404
rect 108 403 109 404
rect 107 403 108 404
rect 106 403 107 404
rect 105 403 106 404
rect 104 403 105 404
rect 80 403 81 404
rect 79 403 80 404
rect 78 403 79 404
rect 77 403 78 404
rect 76 403 77 404
rect 75 403 76 404
rect 74 403 75 404
rect 73 403 74 404
rect 72 403 73 404
rect 71 403 72 404
rect 70 403 71 404
rect 69 403 70 404
rect 68 403 69 404
rect 67 403 68 404
rect 66 403 67 404
rect 65 403 66 404
rect 64 403 65 404
rect 63 403 64 404
rect 62 403 63 404
rect 61 403 62 404
rect 198 404 199 405
rect 196 404 197 405
rect 195 404 196 405
rect 194 404 195 405
rect 193 404 194 405
rect 185 404 186 405
rect 184 404 185 405
rect 183 404 184 405
rect 182 404 183 405
rect 179 404 180 405
rect 178 404 179 405
rect 177 404 178 405
rect 176 404 177 405
rect 175 404 176 405
rect 174 404 175 405
rect 173 404 174 405
rect 172 404 173 405
rect 171 404 172 405
rect 170 404 171 405
rect 169 404 170 405
rect 168 404 169 405
rect 167 404 168 405
rect 166 404 167 405
rect 165 404 166 405
rect 164 404 165 405
rect 143 404 144 405
rect 142 404 143 405
rect 141 404 142 405
rect 140 404 141 405
rect 139 404 140 405
rect 138 404 139 405
rect 137 404 138 405
rect 136 404 137 405
rect 135 404 136 405
rect 134 404 135 405
rect 133 404 134 405
rect 132 404 133 405
rect 131 404 132 405
rect 130 404 131 405
rect 129 404 130 405
rect 114 404 115 405
rect 113 404 114 405
rect 112 404 113 405
rect 111 404 112 405
rect 110 404 111 405
rect 109 404 110 405
rect 108 404 109 405
rect 107 404 108 405
rect 106 404 107 405
rect 105 404 106 405
rect 104 404 105 405
rect 76 404 77 405
rect 75 404 76 405
rect 74 404 75 405
rect 73 404 74 405
rect 72 404 73 405
rect 71 404 72 405
rect 70 404 71 405
rect 69 404 70 405
rect 68 404 69 405
rect 67 404 68 405
rect 66 404 67 405
rect 65 404 66 405
rect 64 404 65 405
rect 196 405 197 406
rect 195 405 196 406
rect 185 405 186 406
rect 184 405 185 406
rect 183 405 184 406
rect 182 405 183 406
rect 179 405 180 406
rect 178 405 179 406
rect 177 405 178 406
rect 176 405 177 406
rect 175 405 176 406
rect 174 405 175 406
rect 173 405 174 406
rect 172 405 173 406
rect 171 405 172 406
rect 170 405 171 406
rect 169 405 170 406
rect 168 405 169 406
rect 167 405 168 406
rect 166 405 167 406
rect 165 405 166 406
rect 164 405 165 406
rect 144 405 145 406
rect 143 405 144 406
rect 142 405 143 406
rect 141 405 142 406
rect 140 405 141 406
rect 139 405 140 406
rect 138 405 139 406
rect 137 405 138 406
rect 136 405 137 406
rect 135 405 136 406
rect 134 405 135 406
rect 133 405 134 406
rect 132 405 133 406
rect 131 405 132 406
rect 130 405 131 406
rect 129 405 130 406
rect 114 405 115 406
rect 113 405 114 406
rect 112 405 113 406
rect 111 405 112 406
rect 110 405 111 406
rect 109 405 110 406
rect 108 405 109 406
rect 107 405 108 406
rect 106 405 107 406
rect 105 405 106 406
rect 104 405 105 406
rect 198 406 199 407
rect 197 406 198 407
rect 196 406 197 407
rect 185 406 186 407
rect 184 406 185 407
rect 183 406 184 407
rect 182 406 183 407
rect 179 406 180 407
rect 178 406 179 407
rect 177 406 178 407
rect 176 406 177 407
rect 175 406 176 407
rect 174 406 175 407
rect 173 406 174 407
rect 172 406 173 407
rect 171 406 172 407
rect 170 406 171 407
rect 169 406 170 407
rect 168 406 169 407
rect 167 406 168 407
rect 166 406 167 407
rect 165 406 166 407
rect 164 406 165 407
rect 145 406 146 407
rect 144 406 145 407
rect 143 406 144 407
rect 142 406 143 407
rect 141 406 142 407
rect 140 406 141 407
rect 139 406 140 407
rect 138 406 139 407
rect 137 406 138 407
rect 136 406 137 407
rect 135 406 136 407
rect 134 406 135 407
rect 133 406 134 407
rect 132 406 133 407
rect 131 406 132 407
rect 130 406 131 407
rect 129 406 130 407
rect 114 406 115 407
rect 113 406 114 407
rect 112 406 113 407
rect 111 406 112 407
rect 110 406 111 407
rect 109 406 110 407
rect 108 406 109 407
rect 107 406 108 407
rect 106 406 107 407
rect 105 406 106 407
rect 104 406 105 407
rect 199 407 200 408
rect 198 407 199 408
rect 197 407 198 408
rect 196 407 197 408
rect 194 407 195 408
rect 193 407 194 408
rect 185 407 186 408
rect 184 407 185 408
rect 183 407 184 408
rect 182 407 183 408
rect 179 407 180 408
rect 178 407 179 408
rect 177 407 178 408
rect 176 407 177 408
rect 175 407 176 408
rect 174 407 175 408
rect 173 407 174 408
rect 172 407 173 408
rect 171 407 172 408
rect 170 407 171 408
rect 169 407 170 408
rect 168 407 169 408
rect 167 407 168 408
rect 166 407 167 408
rect 165 407 166 408
rect 164 407 165 408
rect 146 407 147 408
rect 145 407 146 408
rect 144 407 145 408
rect 143 407 144 408
rect 142 407 143 408
rect 141 407 142 408
rect 140 407 141 408
rect 139 407 140 408
rect 138 407 139 408
rect 137 407 138 408
rect 136 407 137 408
rect 135 407 136 408
rect 134 407 135 408
rect 133 407 134 408
rect 132 407 133 408
rect 131 407 132 408
rect 130 407 131 408
rect 129 407 130 408
rect 114 407 115 408
rect 113 407 114 408
rect 112 407 113 408
rect 111 407 112 408
rect 110 407 111 408
rect 109 407 110 408
rect 108 407 109 408
rect 107 407 108 408
rect 106 407 107 408
rect 105 407 106 408
rect 104 407 105 408
rect 199 408 200 409
rect 198 408 199 409
rect 196 408 197 409
rect 195 408 196 409
rect 194 408 195 409
rect 193 408 194 409
rect 184 408 185 409
rect 183 408 184 409
rect 182 408 183 409
rect 178 408 179 409
rect 177 408 178 409
rect 176 408 177 409
rect 175 408 176 409
rect 174 408 175 409
rect 173 408 174 409
rect 172 408 173 409
rect 171 408 172 409
rect 170 408 171 409
rect 169 408 170 409
rect 168 408 169 409
rect 167 408 168 409
rect 166 408 167 409
rect 165 408 166 409
rect 146 408 147 409
rect 145 408 146 409
rect 144 408 145 409
rect 143 408 144 409
rect 142 408 143 409
rect 141 408 142 409
rect 140 408 141 409
rect 139 408 140 409
rect 138 408 139 409
rect 137 408 138 409
rect 136 408 137 409
rect 135 408 136 409
rect 134 408 135 409
rect 133 408 134 409
rect 132 408 133 409
rect 131 408 132 409
rect 130 408 131 409
rect 129 408 130 409
rect 114 408 115 409
rect 113 408 114 409
rect 112 408 113 409
rect 111 408 112 409
rect 110 408 111 409
rect 109 408 110 409
rect 108 408 109 409
rect 107 408 108 409
rect 106 408 107 409
rect 105 408 106 409
rect 104 408 105 409
rect 198 409 199 410
rect 196 409 197 410
rect 195 409 196 410
rect 194 409 195 410
rect 193 409 194 410
rect 147 409 148 410
rect 146 409 147 410
rect 145 409 146 410
rect 144 409 145 410
rect 143 409 144 410
rect 142 409 143 410
rect 141 409 142 410
rect 140 409 141 410
rect 139 409 140 410
rect 138 409 139 410
rect 137 409 138 410
rect 136 409 137 410
rect 135 409 136 410
rect 134 409 135 410
rect 133 409 134 410
rect 132 409 133 410
rect 131 409 132 410
rect 130 409 131 410
rect 129 409 130 410
rect 114 409 115 410
rect 113 409 114 410
rect 112 409 113 410
rect 111 409 112 410
rect 110 409 111 410
rect 109 409 110 410
rect 108 409 109 410
rect 107 409 108 410
rect 106 409 107 410
rect 105 409 106 410
rect 104 409 105 410
rect 199 410 200 411
rect 198 410 199 411
rect 197 410 198 411
rect 196 410 197 411
rect 195 410 196 411
rect 194 410 195 411
rect 193 410 194 411
rect 148 410 149 411
rect 147 410 148 411
rect 146 410 147 411
rect 145 410 146 411
rect 144 410 145 411
rect 143 410 144 411
rect 142 410 143 411
rect 141 410 142 411
rect 140 410 141 411
rect 139 410 140 411
rect 138 410 139 411
rect 137 410 138 411
rect 136 410 137 411
rect 135 410 136 411
rect 134 410 135 411
rect 133 410 134 411
rect 132 410 133 411
rect 131 410 132 411
rect 130 410 131 411
rect 129 410 130 411
rect 114 410 115 411
rect 113 410 114 411
rect 112 410 113 411
rect 111 410 112 411
rect 110 410 111 411
rect 109 410 110 411
rect 108 410 109 411
rect 107 410 108 411
rect 106 410 107 411
rect 105 410 106 411
rect 104 410 105 411
rect 198 411 199 412
rect 197 411 198 412
rect 196 411 197 412
rect 195 411 196 412
rect 194 411 195 412
rect 193 411 194 412
rect 149 411 150 412
rect 148 411 149 412
rect 147 411 148 412
rect 146 411 147 412
rect 145 411 146 412
rect 144 411 145 412
rect 143 411 144 412
rect 142 411 143 412
rect 141 411 142 412
rect 140 411 141 412
rect 139 411 140 412
rect 138 411 139 412
rect 137 411 138 412
rect 136 411 137 412
rect 135 411 136 412
rect 134 411 135 412
rect 133 411 134 412
rect 132 411 133 412
rect 131 411 132 412
rect 130 411 131 412
rect 129 411 130 412
rect 114 411 115 412
rect 113 411 114 412
rect 112 411 113 412
rect 111 411 112 412
rect 110 411 111 412
rect 109 411 110 412
rect 108 411 109 412
rect 107 411 108 412
rect 106 411 107 412
rect 105 411 106 412
rect 104 411 105 412
rect 150 412 151 413
rect 149 412 150 413
rect 148 412 149 413
rect 147 412 148 413
rect 146 412 147 413
rect 145 412 146 413
rect 144 412 145 413
rect 143 412 144 413
rect 142 412 143 413
rect 141 412 142 413
rect 140 412 141 413
rect 139 412 140 413
rect 138 412 139 413
rect 137 412 138 413
rect 136 412 137 413
rect 135 412 136 413
rect 134 412 135 413
rect 133 412 134 413
rect 132 412 133 413
rect 131 412 132 413
rect 130 412 131 413
rect 129 412 130 413
rect 114 412 115 413
rect 113 412 114 413
rect 112 412 113 413
rect 111 412 112 413
rect 110 412 111 413
rect 109 412 110 413
rect 108 412 109 413
rect 107 412 108 413
rect 106 412 107 413
rect 105 412 106 413
rect 104 412 105 413
rect 198 413 199 414
rect 197 413 198 414
rect 196 413 197 414
rect 195 413 196 414
rect 194 413 195 414
rect 193 413 194 414
rect 151 413 152 414
rect 150 413 151 414
rect 149 413 150 414
rect 148 413 149 414
rect 147 413 148 414
rect 146 413 147 414
rect 145 413 146 414
rect 144 413 145 414
rect 143 413 144 414
rect 142 413 143 414
rect 141 413 142 414
rect 140 413 141 414
rect 139 413 140 414
rect 138 413 139 414
rect 137 413 138 414
rect 136 413 137 414
rect 135 413 136 414
rect 134 413 135 414
rect 133 413 134 414
rect 132 413 133 414
rect 131 413 132 414
rect 130 413 131 414
rect 129 413 130 414
rect 114 413 115 414
rect 113 413 114 414
rect 112 413 113 414
rect 111 413 112 414
rect 110 413 111 414
rect 109 413 110 414
rect 108 413 109 414
rect 107 413 108 414
rect 106 413 107 414
rect 105 413 106 414
rect 104 413 105 414
rect 199 414 200 415
rect 198 414 199 415
rect 197 414 198 415
rect 196 414 197 415
rect 195 414 196 415
rect 194 414 195 415
rect 193 414 194 415
rect 151 414 152 415
rect 150 414 151 415
rect 149 414 150 415
rect 148 414 149 415
rect 147 414 148 415
rect 146 414 147 415
rect 145 414 146 415
rect 144 414 145 415
rect 143 414 144 415
rect 142 414 143 415
rect 141 414 142 415
rect 140 414 141 415
rect 139 414 140 415
rect 138 414 139 415
rect 137 414 138 415
rect 136 414 137 415
rect 135 414 136 415
rect 134 414 135 415
rect 133 414 134 415
rect 132 414 133 415
rect 131 414 132 415
rect 130 414 131 415
rect 129 414 130 415
rect 128 414 129 415
rect 127 414 128 415
rect 126 414 127 415
rect 125 414 126 415
rect 124 414 125 415
rect 123 414 124 415
rect 122 414 123 415
rect 121 414 122 415
rect 120 414 121 415
rect 119 414 120 415
rect 118 414 119 415
rect 117 414 118 415
rect 116 414 117 415
rect 115 414 116 415
rect 114 414 115 415
rect 113 414 114 415
rect 112 414 113 415
rect 111 414 112 415
rect 110 414 111 415
rect 109 414 110 415
rect 108 414 109 415
rect 107 414 108 415
rect 106 414 107 415
rect 105 414 106 415
rect 104 414 105 415
rect 194 415 195 416
rect 193 415 194 416
rect 152 415 153 416
rect 151 415 152 416
rect 150 415 151 416
rect 149 415 150 416
rect 148 415 149 416
rect 147 415 148 416
rect 146 415 147 416
rect 145 415 146 416
rect 144 415 145 416
rect 143 415 144 416
rect 142 415 143 416
rect 141 415 142 416
rect 140 415 141 416
rect 139 415 140 416
rect 138 415 139 416
rect 137 415 138 416
rect 136 415 137 416
rect 135 415 136 416
rect 134 415 135 416
rect 133 415 134 416
rect 132 415 133 416
rect 131 415 132 416
rect 130 415 131 416
rect 129 415 130 416
rect 128 415 129 416
rect 127 415 128 416
rect 126 415 127 416
rect 125 415 126 416
rect 124 415 125 416
rect 123 415 124 416
rect 122 415 123 416
rect 121 415 122 416
rect 120 415 121 416
rect 119 415 120 416
rect 118 415 119 416
rect 117 415 118 416
rect 116 415 117 416
rect 115 415 116 416
rect 114 415 115 416
rect 113 415 114 416
rect 112 415 113 416
rect 111 415 112 416
rect 110 415 111 416
rect 109 415 110 416
rect 108 415 109 416
rect 107 415 108 416
rect 106 415 107 416
rect 105 415 106 416
rect 104 415 105 416
rect 194 416 195 417
rect 193 416 194 417
rect 153 416 154 417
rect 152 416 153 417
rect 151 416 152 417
rect 150 416 151 417
rect 149 416 150 417
rect 148 416 149 417
rect 147 416 148 417
rect 146 416 147 417
rect 145 416 146 417
rect 144 416 145 417
rect 143 416 144 417
rect 142 416 143 417
rect 141 416 142 417
rect 140 416 141 417
rect 139 416 140 417
rect 138 416 139 417
rect 137 416 138 417
rect 136 416 137 417
rect 135 416 136 417
rect 134 416 135 417
rect 133 416 134 417
rect 132 416 133 417
rect 131 416 132 417
rect 129 416 130 417
rect 128 416 129 417
rect 127 416 128 417
rect 126 416 127 417
rect 125 416 126 417
rect 124 416 125 417
rect 123 416 124 417
rect 122 416 123 417
rect 121 416 122 417
rect 120 416 121 417
rect 119 416 120 417
rect 118 416 119 417
rect 117 416 118 417
rect 116 416 117 417
rect 115 416 116 417
rect 114 416 115 417
rect 113 416 114 417
rect 112 416 113 417
rect 111 416 112 417
rect 110 416 111 417
rect 109 416 110 417
rect 108 416 109 417
rect 107 416 108 417
rect 106 416 107 417
rect 105 416 106 417
rect 104 416 105 417
rect 198 417 199 418
rect 197 417 198 418
rect 196 417 197 418
rect 195 417 196 418
rect 194 417 195 418
rect 154 417 155 418
rect 153 417 154 418
rect 152 417 153 418
rect 151 417 152 418
rect 150 417 151 418
rect 149 417 150 418
rect 148 417 149 418
rect 147 417 148 418
rect 146 417 147 418
rect 145 417 146 418
rect 144 417 145 418
rect 143 417 144 418
rect 142 417 143 418
rect 141 417 142 418
rect 140 417 141 418
rect 139 417 140 418
rect 138 417 139 418
rect 137 417 138 418
rect 136 417 137 418
rect 135 417 136 418
rect 134 417 135 418
rect 133 417 134 418
rect 132 417 133 418
rect 129 417 130 418
rect 128 417 129 418
rect 127 417 128 418
rect 126 417 127 418
rect 125 417 126 418
rect 124 417 125 418
rect 123 417 124 418
rect 122 417 123 418
rect 121 417 122 418
rect 120 417 121 418
rect 119 417 120 418
rect 118 417 119 418
rect 117 417 118 418
rect 116 417 117 418
rect 115 417 116 418
rect 114 417 115 418
rect 113 417 114 418
rect 112 417 113 418
rect 111 417 112 418
rect 110 417 111 418
rect 109 417 110 418
rect 108 417 109 418
rect 107 417 108 418
rect 106 417 107 418
rect 105 417 106 418
rect 104 417 105 418
rect 198 418 199 419
rect 197 418 198 419
rect 196 418 197 419
rect 195 418 196 419
rect 194 418 195 419
rect 193 418 194 419
rect 155 418 156 419
rect 154 418 155 419
rect 153 418 154 419
rect 152 418 153 419
rect 151 418 152 419
rect 150 418 151 419
rect 149 418 150 419
rect 148 418 149 419
rect 147 418 148 419
rect 146 418 147 419
rect 145 418 146 419
rect 144 418 145 419
rect 143 418 144 419
rect 142 418 143 419
rect 141 418 142 419
rect 140 418 141 419
rect 139 418 140 419
rect 138 418 139 419
rect 137 418 138 419
rect 136 418 137 419
rect 135 418 136 419
rect 134 418 135 419
rect 133 418 134 419
rect 129 418 130 419
rect 128 418 129 419
rect 127 418 128 419
rect 126 418 127 419
rect 125 418 126 419
rect 124 418 125 419
rect 123 418 124 419
rect 122 418 123 419
rect 121 418 122 419
rect 120 418 121 419
rect 119 418 120 419
rect 118 418 119 419
rect 117 418 118 419
rect 116 418 117 419
rect 115 418 116 419
rect 114 418 115 419
rect 113 418 114 419
rect 112 418 113 419
rect 111 418 112 419
rect 110 418 111 419
rect 109 418 110 419
rect 108 418 109 419
rect 107 418 108 419
rect 106 418 107 419
rect 105 418 106 419
rect 104 418 105 419
rect 198 419 199 420
rect 197 419 198 420
rect 194 419 195 420
rect 193 419 194 420
rect 155 419 156 420
rect 154 419 155 420
rect 153 419 154 420
rect 152 419 153 420
rect 151 419 152 420
rect 150 419 151 420
rect 149 419 150 420
rect 148 419 149 420
rect 147 419 148 420
rect 146 419 147 420
rect 145 419 146 420
rect 144 419 145 420
rect 143 419 144 420
rect 142 419 143 420
rect 141 419 142 420
rect 140 419 141 420
rect 139 419 140 420
rect 138 419 139 420
rect 137 419 138 420
rect 136 419 137 420
rect 135 419 136 420
rect 134 419 135 420
rect 133 419 134 420
rect 129 419 130 420
rect 128 419 129 420
rect 127 419 128 420
rect 126 419 127 420
rect 125 419 126 420
rect 124 419 125 420
rect 123 419 124 420
rect 122 419 123 420
rect 121 419 122 420
rect 120 419 121 420
rect 119 419 120 420
rect 118 419 119 420
rect 117 419 118 420
rect 116 419 117 420
rect 115 419 116 420
rect 114 419 115 420
rect 113 419 114 420
rect 112 419 113 420
rect 111 419 112 420
rect 110 419 111 420
rect 109 419 110 420
rect 108 419 109 420
rect 107 419 108 420
rect 106 419 107 420
rect 105 419 106 420
rect 104 419 105 420
rect 199 420 200 421
rect 198 420 199 421
rect 194 420 195 421
rect 193 420 194 421
rect 176 420 177 421
rect 175 420 176 421
rect 174 420 175 421
rect 155 420 156 421
rect 154 420 155 421
rect 153 420 154 421
rect 152 420 153 421
rect 151 420 152 421
rect 150 420 151 421
rect 149 420 150 421
rect 148 420 149 421
rect 147 420 148 421
rect 146 420 147 421
rect 145 420 146 421
rect 144 420 145 421
rect 143 420 144 421
rect 142 420 143 421
rect 141 420 142 421
rect 140 420 141 421
rect 139 420 140 421
rect 138 420 139 421
rect 137 420 138 421
rect 136 420 137 421
rect 135 420 136 421
rect 134 420 135 421
rect 129 420 130 421
rect 128 420 129 421
rect 127 420 128 421
rect 126 420 127 421
rect 125 420 126 421
rect 124 420 125 421
rect 123 420 124 421
rect 122 420 123 421
rect 121 420 122 421
rect 120 420 121 421
rect 119 420 120 421
rect 118 420 119 421
rect 117 420 118 421
rect 116 420 117 421
rect 115 420 116 421
rect 114 420 115 421
rect 113 420 114 421
rect 112 420 113 421
rect 111 420 112 421
rect 110 420 111 421
rect 109 420 110 421
rect 108 420 109 421
rect 107 420 108 421
rect 106 420 107 421
rect 105 420 106 421
rect 104 420 105 421
rect 198 421 199 422
rect 193 421 194 422
rect 176 421 177 422
rect 175 421 176 422
rect 174 421 175 422
rect 155 421 156 422
rect 154 421 155 422
rect 153 421 154 422
rect 152 421 153 422
rect 151 421 152 422
rect 150 421 151 422
rect 149 421 150 422
rect 148 421 149 422
rect 147 421 148 422
rect 146 421 147 422
rect 145 421 146 422
rect 144 421 145 422
rect 143 421 144 422
rect 142 421 143 422
rect 141 421 142 422
rect 140 421 141 422
rect 139 421 140 422
rect 138 421 139 422
rect 137 421 138 422
rect 136 421 137 422
rect 135 421 136 422
rect 129 421 130 422
rect 128 421 129 422
rect 127 421 128 422
rect 126 421 127 422
rect 125 421 126 422
rect 124 421 125 422
rect 123 421 124 422
rect 122 421 123 422
rect 121 421 122 422
rect 120 421 121 422
rect 119 421 120 422
rect 118 421 119 422
rect 117 421 118 422
rect 116 421 117 422
rect 115 421 116 422
rect 114 421 115 422
rect 113 421 114 422
rect 112 421 113 422
rect 111 421 112 422
rect 110 421 111 422
rect 109 421 110 422
rect 108 421 109 422
rect 107 421 108 422
rect 106 421 107 422
rect 105 421 106 422
rect 104 421 105 422
rect 176 422 177 423
rect 175 422 176 423
rect 174 422 175 423
rect 166 422 167 423
rect 155 422 156 423
rect 154 422 155 423
rect 153 422 154 423
rect 152 422 153 423
rect 151 422 152 423
rect 150 422 151 423
rect 149 422 150 423
rect 148 422 149 423
rect 147 422 148 423
rect 146 422 147 423
rect 145 422 146 423
rect 144 422 145 423
rect 143 422 144 423
rect 142 422 143 423
rect 141 422 142 423
rect 140 422 141 423
rect 139 422 140 423
rect 138 422 139 423
rect 137 422 138 423
rect 136 422 137 423
rect 129 422 130 423
rect 128 422 129 423
rect 127 422 128 423
rect 126 422 127 423
rect 125 422 126 423
rect 124 422 125 423
rect 123 422 124 423
rect 122 422 123 423
rect 121 422 122 423
rect 120 422 121 423
rect 119 422 120 423
rect 118 422 119 423
rect 117 422 118 423
rect 116 422 117 423
rect 115 422 116 423
rect 114 422 115 423
rect 113 422 114 423
rect 112 422 113 423
rect 111 422 112 423
rect 110 422 111 423
rect 109 422 110 423
rect 108 422 109 423
rect 107 422 108 423
rect 106 422 107 423
rect 105 422 106 423
rect 104 422 105 423
rect 199 423 200 424
rect 198 423 199 424
rect 197 423 198 424
rect 196 423 197 424
rect 195 423 196 424
rect 194 423 195 424
rect 193 423 194 424
rect 192 423 193 424
rect 191 423 192 424
rect 190 423 191 424
rect 176 423 177 424
rect 175 423 176 424
rect 174 423 175 424
rect 167 423 168 424
rect 166 423 167 424
rect 165 423 166 424
rect 155 423 156 424
rect 154 423 155 424
rect 153 423 154 424
rect 152 423 153 424
rect 151 423 152 424
rect 150 423 151 424
rect 149 423 150 424
rect 148 423 149 424
rect 147 423 148 424
rect 146 423 147 424
rect 145 423 146 424
rect 144 423 145 424
rect 143 423 144 424
rect 142 423 143 424
rect 141 423 142 424
rect 140 423 141 424
rect 139 423 140 424
rect 138 423 139 424
rect 137 423 138 424
rect 129 423 130 424
rect 128 423 129 424
rect 127 423 128 424
rect 126 423 127 424
rect 125 423 126 424
rect 124 423 125 424
rect 123 423 124 424
rect 122 423 123 424
rect 121 423 122 424
rect 120 423 121 424
rect 119 423 120 424
rect 118 423 119 424
rect 117 423 118 424
rect 116 423 117 424
rect 115 423 116 424
rect 114 423 115 424
rect 113 423 114 424
rect 112 423 113 424
rect 111 423 112 424
rect 110 423 111 424
rect 109 423 110 424
rect 108 423 109 424
rect 107 423 108 424
rect 106 423 107 424
rect 105 423 106 424
rect 104 423 105 424
rect 198 424 199 425
rect 197 424 198 425
rect 196 424 197 425
rect 195 424 196 425
rect 194 424 195 425
rect 193 424 194 425
rect 192 424 193 425
rect 191 424 192 425
rect 190 424 191 425
rect 176 424 177 425
rect 175 424 176 425
rect 174 424 175 425
rect 167 424 168 425
rect 166 424 167 425
rect 165 424 166 425
rect 155 424 156 425
rect 154 424 155 425
rect 153 424 154 425
rect 152 424 153 425
rect 151 424 152 425
rect 150 424 151 425
rect 149 424 150 425
rect 148 424 149 425
rect 147 424 148 425
rect 146 424 147 425
rect 145 424 146 425
rect 144 424 145 425
rect 143 424 144 425
rect 142 424 143 425
rect 141 424 142 425
rect 140 424 141 425
rect 139 424 140 425
rect 138 424 139 425
rect 129 424 130 425
rect 128 424 129 425
rect 127 424 128 425
rect 126 424 127 425
rect 125 424 126 425
rect 124 424 125 425
rect 123 424 124 425
rect 122 424 123 425
rect 121 424 122 425
rect 120 424 121 425
rect 119 424 120 425
rect 118 424 119 425
rect 117 424 118 425
rect 116 424 117 425
rect 115 424 116 425
rect 114 424 115 425
rect 113 424 114 425
rect 112 424 113 425
rect 111 424 112 425
rect 110 424 111 425
rect 109 424 110 425
rect 108 424 109 425
rect 107 424 108 425
rect 106 424 107 425
rect 105 424 106 425
rect 104 424 105 425
rect 194 425 195 426
rect 193 425 194 426
rect 176 425 177 426
rect 175 425 176 426
rect 174 425 175 426
rect 167 425 168 426
rect 166 425 167 426
rect 165 425 166 426
rect 155 425 156 426
rect 154 425 155 426
rect 153 425 154 426
rect 152 425 153 426
rect 151 425 152 426
rect 150 425 151 426
rect 149 425 150 426
rect 148 425 149 426
rect 147 425 148 426
rect 146 425 147 426
rect 145 425 146 426
rect 144 425 145 426
rect 143 425 144 426
rect 142 425 143 426
rect 141 425 142 426
rect 140 425 141 426
rect 139 425 140 426
rect 138 425 139 426
rect 129 425 130 426
rect 128 425 129 426
rect 127 425 128 426
rect 126 425 127 426
rect 125 425 126 426
rect 124 425 125 426
rect 123 425 124 426
rect 122 425 123 426
rect 121 425 122 426
rect 120 425 121 426
rect 119 425 120 426
rect 118 425 119 426
rect 117 425 118 426
rect 116 425 117 426
rect 115 425 116 426
rect 114 425 115 426
rect 113 425 114 426
rect 112 425 113 426
rect 111 425 112 426
rect 110 425 111 426
rect 109 425 110 426
rect 108 425 109 426
rect 107 425 108 426
rect 106 425 107 426
rect 105 425 106 426
rect 104 425 105 426
rect 198 426 199 427
rect 197 426 198 427
rect 196 426 197 427
rect 194 426 195 427
rect 193 426 194 427
rect 176 426 177 427
rect 175 426 176 427
rect 174 426 175 427
rect 167 426 168 427
rect 166 426 167 427
rect 165 426 166 427
rect 155 426 156 427
rect 154 426 155 427
rect 153 426 154 427
rect 152 426 153 427
rect 151 426 152 427
rect 150 426 151 427
rect 149 426 150 427
rect 148 426 149 427
rect 147 426 148 427
rect 146 426 147 427
rect 145 426 146 427
rect 144 426 145 427
rect 143 426 144 427
rect 142 426 143 427
rect 141 426 142 427
rect 140 426 141 427
rect 139 426 140 427
rect 129 426 130 427
rect 128 426 129 427
rect 127 426 128 427
rect 126 426 127 427
rect 125 426 126 427
rect 124 426 125 427
rect 123 426 124 427
rect 122 426 123 427
rect 121 426 122 427
rect 120 426 121 427
rect 119 426 120 427
rect 118 426 119 427
rect 117 426 118 427
rect 116 426 117 427
rect 115 426 116 427
rect 114 426 115 427
rect 113 426 114 427
rect 112 426 113 427
rect 111 426 112 427
rect 110 426 111 427
rect 109 426 110 427
rect 108 426 109 427
rect 107 426 108 427
rect 106 426 107 427
rect 105 426 106 427
rect 104 426 105 427
rect 199 427 200 428
rect 198 427 199 428
rect 197 427 198 428
rect 196 427 197 428
rect 195 427 196 428
rect 194 427 195 428
rect 193 427 194 428
rect 176 427 177 428
rect 175 427 176 428
rect 174 427 175 428
rect 167 427 168 428
rect 166 427 167 428
rect 165 427 166 428
rect 155 427 156 428
rect 154 427 155 428
rect 153 427 154 428
rect 152 427 153 428
rect 151 427 152 428
rect 150 427 151 428
rect 149 427 150 428
rect 148 427 149 428
rect 147 427 148 428
rect 146 427 147 428
rect 145 427 146 428
rect 144 427 145 428
rect 143 427 144 428
rect 142 427 143 428
rect 141 427 142 428
rect 140 427 141 428
rect 129 427 130 428
rect 128 427 129 428
rect 127 427 128 428
rect 126 427 127 428
rect 125 427 126 428
rect 124 427 125 428
rect 123 427 124 428
rect 122 427 123 428
rect 121 427 122 428
rect 120 427 121 428
rect 119 427 120 428
rect 118 427 119 428
rect 117 427 118 428
rect 116 427 117 428
rect 115 427 116 428
rect 114 427 115 428
rect 113 427 114 428
rect 112 427 113 428
rect 111 427 112 428
rect 110 427 111 428
rect 109 427 110 428
rect 108 427 109 428
rect 107 427 108 428
rect 106 427 107 428
rect 105 427 106 428
rect 104 427 105 428
rect 176 428 177 429
rect 175 428 176 429
rect 174 428 175 429
rect 167 428 168 429
rect 166 428 167 429
rect 165 428 166 429
rect 155 428 156 429
rect 154 428 155 429
rect 153 428 154 429
rect 152 428 153 429
rect 151 428 152 429
rect 150 428 151 429
rect 149 428 150 429
rect 148 428 149 429
rect 147 428 148 429
rect 146 428 147 429
rect 145 428 146 429
rect 144 428 145 429
rect 143 428 144 429
rect 142 428 143 429
rect 141 428 142 429
rect 129 428 130 429
rect 128 428 129 429
rect 127 428 128 429
rect 126 428 127 429
rect 125 428 126 429
rect 124 428 125 429
rect 123 428 124 429
rect 122 428 123 429
rect 121 428 122 429
rect 120 428 121 429
rect 119 428 120 429
rect 118 428 119 429
rect 117 428 118 429
rect 116 428 117 429
rect 115 428 116 429
rect 114 428 115 429
rect 113 428 114 429
rect 112 428 113 429
rect 111 428 112 429
rect 110 428 111 429
rect 109 428 110 429
rect 108 428 109 429
rect 107 428 108 429
rect 106 428 107 429
rect 105 428 106 429
rect 104 428 105 429
rect 176 429 177 430
rect 175 429 176 430
rect 174 429 175 430
rect 167 429 168 430
rect 166 429 167 430
rect 165 429 166 430
rect 155 429 156 430
rect 154 429 155 430
rect 153 429 154 430
rect 152 429 153 430
rect 151 429 152 430
rect 150 429 151 430
rect 149 429 150 430
rect 148 429 149 430
rect 147 429 148 430
rect 146 429 147 430
rect 145 429 146 430
rect 144 429 145 430
rect 143 429 144 430
rect 142 429 143 430
rect 129 429 130 430
rect 128 429 129 430
rect 127 429 128 430
rect 126 429 127 430
rect 125 429 126 430
rect 124 429 125 430
rect 123 429 124 430
rect 122 429 123 430
rect 121 429 122 430
rect 120 429 121 430
rect 119 429 120 430
rect 118 429 119 430
rect 117 429 118 430
rect 116 429 117 430
rect 115 429 116 430
rect 114 429 115 430
rect 113 429 114 430
rect 112 429 113 430
rect 111 429 112 430
rect 110 429 111 430
rect 109 429 110 430
rect 108 429 109 430
rect 107 429 108 430
rect 106 429 107 430
rect 105 429 106 430
rect 104 429 105 430
rect 185 430 186 431
rect 184 430 185 431
rect 183 430 184 431
rect 182 430 183 431
rect 181 430 182 431
rect 180 430 181 431
rect 179 430 180 431
rect 178 430 179 431
rect 177 430 178 431
rect 176 430 177 431
rect 175 430 176 431
rect 174 430 175 431
rect 167 430 168 431
rect 166 430 167 431
rect 165 430 166 431
rect 155 430 156 431
rect 154 430 155 431
rect 153 430 154 431
rect 152 430 153 431
rect 151 430 152 431
rect 150 430 151 431
rect 149 430 150 431
rect 148 430 149 431
rect 147 430 148 431
rect 146 430 147 431
rect 145 430 146 431
rect 144 430 145 431
rect 143 430 144 431
rect 142 430 143 431
rect 129 430 130 431
rect 128 430 129 431
rect 127 430 128 431
rect 126 430 127 431
rect 125 430 126 431
rect 124 430 125 431
rect 123 430 124 431
rect 122 430 123 431
rect 121 430 122 431
rect 120 430 121 431
rect 119 430 120 431
rect 118 430 119 431
rect 117 430 118 431
rect 116 430 117 431
rect 115 430 116 431
rect 114 430 115 431
rect 113 430 114 431
rect 112 430 113 431
rect 111 430 112 431
rect 110 430 111 431
rect 109 430 110 431
rect 108 430 109 431
rect 107 430 108 431
rect 106 430 107 431
rect 105 430 106 431
rect 185 431 186 432
rect 184 431 185 432
rect 183 431 184 432
rect 182 431 183 432
rect 181 431 182 432
rect 180 431 181 432
rect 179 431 180 432
rect 178 431 179 432
rect 177 431 178 432
rect 176 431 177 432
rect 175 431 176 432
rect 174 431 175 432
rect 167 431 168 432
rect 166 431 167 432
rect 165 431 166 432
rect 155 431 156 432
rect 154 431 155 432
rect 153 431 154 432
rect 152 431 153 432
rect 151 431 152 432
rect 150 431 151 432
rect 149 431 150 432
rect 148 431 149 432
rect 147 431 148 432
rect 146 431 147 432
rect 145 431 146 432
rect 144 431 145 432
rect 143 431 144 432
rect 129 431 130 432
rect 128 431 129 432
rect 127 431 128 432
rect 126 431 127 432
rect 125 431 126 432
rect 124 431 125 432
rect 123 431 124 432
rect 122 431 123 432
rect 121 431 122 432
rect 120 431 121 432
rect 119 431 120 432
rect 118 431 119 432
rect 117 431 118 432
rect 116 431 117 432
rect 115 431 116 432
rect 114 431 115 432
rect 113 431 114 432
rect 112 431 113 432
rect 111 431 112 432
rect 110 431 111 432
rect 109 431 110 432
rect 108 431 109 432
rect 107 431 108 432
rect 106 431 107 432
rect 105 431 106 432
rect 198 432 199 433
rect 197 432 198 433
rect 196 432 197 433
rect 195 432 196 433
rect 194 432 195 433
rect 193 432 194 433
rect 192 432 193 433
rect 191 432 192 433
rect 185 432 186 433
rect 184 432 185 433
rect 183 432 184 433
rect 182 432 183 433
rect 181 432 182 433
rect 180 432 181 433
rect 179 432 180 433
rect 178 432 179 433
rect 177 432 178 433
rect 176 432 177 433
rect 175 432 176 433
rect 174 432 175 433
rect 167 432 168 433
rect 166 432 167 433
rect 165 432 166 433
rect 155 432 156 433
rect 154 432 155 433
rect 153 432 154 433
rect 152 432 153 433
rect 151 432 152 433
rect 150 432 151 433
rect 149 432 150 433
rect 148 432 149 433
rect 147 432 148 433
rect 146 432 147 433
rect 145 432 146 433
rect 144 432 145 433
rect 129 432 130 433
rect 128 432 129 433
rect 127 432 128 433
rect 126 432 127 433
rect 125 432 126 433
rect 124 432 125 433
rect 123 432 124 433
rect 122 432 123 433
rect 121 432 122 433
rect 120 432 121 433
rect 119 432 120 433
rect 118 432 119 433
rect 117 432 118 433
rect 116 432 117 433
rect 115 432 116 433
rect 114 432 115 433
rect 113 432 114 433
rect 112 432 113 433
rect 111 432 112 433
rect 110 432 111 433
rect 109 432 110 433
rect 108 432 109 433
rect 107 432 108 433
rect 106 432 107 433
rect 105 432 106 433
rect 199 433 200 434
rect 198 433 199 434
rect 197 433 198 434
rect 196 433 197 434
rect 195 433 196 434
rect 194 433 195 434
rect 193 433 194 434
rect 192 433 193 434
rect 191 433 192 434
rect 185 433 186 434
rect 184 433 185 434
rect 183 433 184 434
rect 182 433 183 434
rect 181 433 182 434
rect 180 433 181 434
rect 179 433 180 434
rect 178 433 179 434
rect 177 433 178 434
rect 176 433 177 434
rect 175 433 176 434
rect 174 433 175 434
rect 167 433 168 434
rect 166 433 167 434
rect 165 433 166 434
rect 155 433 156 434
rect 154 433 155 434
rect 153 433 154 434
rect 152 433 153 434
rect 151 433 152 434
rect 150 433 151 434
rect 149 433 150 434
rect 148 433 149 434
rect 147 433 148 434
rect 146 433 147 434
rect 145 433 146 434
rect 129 433 130 434
rect 128 433 129 434
rect 127 433 128 434
rect 126 433 127 434
rect 125 433 126 434
rect 124 433 125 434
rect 123 433 124 434
rect 122 433 123 434
rect 121 433 122 434
rect 120 433 121 434
rect 119 433 120 434
rect 118 433 119 434
rect 117 433 118 434
rect 116 433 117 434
rect 115 433 116 434
rect 114 433 115 434
rect 113 433 114 434
rect 112 433 113 434
rect 111 433 112 434
rect 110 433 111 434
rect 109 433 110 434
rect 108 433 109 434
rect 107 433 108 434
rect 106 433 107 434
rect 198 434 199 435
rect 197 434 198 435
rect 196 434 197 435
rect 195 434 196 435
rect 194 434 195 435
rect 193 434 194 435
rect 192 434 193 435
rect 191 434 192 435
rect 176 434 177 435
rect 175 434 176 435
rect 174 434 175 435
rect 167 434 168 435
rect 166 434 167 435
rect 165 434 166 435
rect 155 434 156 435
rect 154 434 155 435
rect 153 434 154 435
rect 152 434 153 435
rect 151 434 152 435
rect 150 434 151 435
rect 149 434 150 435
rect 148 434 149 435
rect 147 434 148 435
rect 146 434 147 435
rect 129 434 130 435
rect 128 434 129 435
rect 127 434 128 435
rect 126 434 127 435
rect 125 434 126 435
rect 124 434 125 435
rect 123 434 124 435
rect 122 434 123 435
rect 121 434 122 435
rect 120 434 121 435
rect 119 434 120 435
rect 118 434 119 435
rect 117 434 118 435
rect 116 434 117 435
rect 115 434 116 435
rect 114 434 115 435
rect 113 434 114 435
rect 112 434 113 435
rect 111 434 112 435
rect 110 434 111 435
rect 109 434 110 435
rect 108 434 109 435
rect 107 434 108 435
rect 176 435 177 436
rect 175 435 176 436
rect 174 435 175 436
rect 167 435 168 436
rect 166 435 167 436
rect 165 435 166 436
rect 155 435 156 436
rect 154 435 155 436
rect 153 435 154 436
rect 152 435 153 436
rect 151 435 152 436
rect 150 435 151 436
rect 149 435 150 436
rect 148 435 149 436
rect 147 435 148 436
rect 146 435 147 436
rect 129 435 130 436
rect 128 435 129 436
rect 127 435 128 436
rect 126 435 127 436
rect 125 435 126 436
rect 124 435 125 436
rect 123 435 124 436
rect 122 435 123 436
rect 121 435 122 436
rect 120 435 121 436
rect 119 435 120 436
rect 118 435 119 436
rect 117 435 118 436
rect 116 435 117 436
rect 115 435 116 436
rect 114 435 115 436
rect 113 435 114 436
rect 112 435 113 436
rect 111 435 112 436
rect 110 435 111 436
rect 109 435 110 436
rect 108 435 109 436
rect 198 436 199 437
rect 197 436 198 437
rect 196 436 197 437
rect 195 436 196 437
rect 194 436 195 437
rect 193 436 194 437
rect 176 436 177 437
rect 175 436 176 437
rect 174 436 175 437
rect 167 436 168 437
rect 166 436 167 437
rect 165 436 166 437
rect 155 436 156 437
rect 154 436 155 437
rect 153 436 154 437
rect 152 436 153 437
rect 151 436 152 437
rect 150 436 151 437
rect 149 436 150 437
rect 148 436 149 437
rect 147 436 148 437
rect 129 436 130 437
rect 128 436 129 437
rect 127 436 128 437
rect 126 436 127 437
rect 125 436 126 437
rect 124 436 125 437
rect 123 436 124 437
rect 122 436 123 437
rect 121 436 122 437
rect 120 436 121 437
rect 119 436 120 437
rect 118 436 119 437
rect 117 436 118 437
rect 116 436 117 437
rect 115 436 116 437
rect 114 436 115 437
rect 113 436 114 437
rect 112 436 113 437
rect 111 436 112 437
rect 110 436 111 437
rect 109 436 110 437
rect 199 437 200 438
rect 198 437 199 438
rect 197 437 198 438
rect 196 437 197 438
rect 195 437 196 438
rect 194 437 195 438
rect 193 437 194 438
rect 176 437 177 438
rect 175 437 176 438
rect 174 437 175 438
rect 173 437 174 438
rect 172 437 173 438
rect 171 437 172 438
rect 170 437 171 438
rect 169 437 170 438
rect 168 437 169 438
rect 167 437 168 438
rect 166 437 167 438
rect 165 437 166 438
rect 155 437 156 438
rect 154 437 155 438
rect 153 437 154 438
rect 152 437 153 438
rect 151 437 152 438
rect 150 437 151 438
rect 149 437 150 438
rect 148 437 149 438
rect 129 437 130 438
rect 128 437 129 438
rect 127 437 128 438
rect 126 437 127 438
rect 125 437 126 438
rect 124 437 125 438
rect 123 437 124 438
rect 122 437 123 438
rect 121 437 122 438
rect 120 437 121 438
rect 119 437 120 438
rect 118 437 119 438
rect 117 437 118 438
rect 116 437 117 438
rect 115 437 116 438
rect 114 437 115 438
rect 113 437 114 438
rect 112 437 113 438
rect 111 437 112 438
rect 110 437 111 438
rect 194 438 195 439
rect 193 438 194 439
rect 176 438 177 439
rect 175 438 176 439
rect 174 438 175 439
rect 173 438 174 439
rect 172 438 173 439
rect 171 438 172 439
rect 170 438 171 439
rect 169 438 170 439
rect 168 438 169 439
rect 167 438 168 439
rect 166 438 167 439
rect 165 438 166 439
rect 155 438 156 439
rect 154 438 155 439
rect 153 438 154 439
rect 152 438 153 439
rect 151 438 152 439
rect 150 438 151 439
rect 149 438 150 439
rect 194 439 195 440
rect 193 439 194 440
rect 176 439 177 440
rect 175 439 176 440
rect 174 439 175 440
rect 173 439 174 440
rect 172 439 173 440
rect 171 439 172 440
rect 170 439 171 440
rect 169 439 170 440
rect 168 439 169 440
rect 167 439 168 440
rect 166 439 167 440
rect 165 439 166 440
rect 155 439 156 440
rect 154 439 155 440
rect 153 439 154 440
rect 152 439 153 440
rect 151 439 152 440
rect 150 439 151 440
rect 198 440 199 441
rect 197 440 198 441
rect 196 440 197 441
rect 195 440 196 441
rect 194 440 195 441
rect 193 440 194 441
rect 176 440 177 441
rect 175 440 176 441
rect 174 440 175 441
rect 172 440 173 441
rect 171 440 172 441
rect 170 440 171 441
rect 169 440 170 441
rect 168 440 169 441
rect 167 440 168 441
rect 166 440 167 441
rect 165 440 166 441
rect 155 440 156 441
rect 154 440 155 441
rect 153 440 154 441
rect 152 440 153 441
rect 151 440 152 441
rect 199 441 200 442
rect 198 441 199 442
rect 197 441 198 442
rect 196 441 197 442
rect 195 441 196 442
rect 194 441 195 442
rect 193 441 194 442
rect 176 441 177 442
rect 175 441 176 442
rect 174 441 175 442
rect 169 441 170 442
rect 168 441 169 442
rect 167 441 168 442
rect 166 441 167 442
rect 165 441 166 442
rect 155 441 156 442
rect 154 441 155 442
rect 153 441 154 442
rect 152 441 153 442
rect 151 441 152 442
rect 194 442 195 443
rect 176 442 177 443
rect 175 442 176 443
rect 174 442 175 443
rect 155 442 156 443
rect 154 442 155 443
rect 153 442 154 443
rect 152 442 153 443
rect 198 443 199 444
rect 195 443 196 444
rect 194 443 195 444
rect 176 443 177 444
rect 175 443 176 444
rect 174 443 175 444
rect 155 443 156 444
rect 154 443 155 444
rect 153 443 154 444
rect 199 444 200 445
rect 198 444 199 445
rect 196 444 197 445
rect 195 444 196 445
rect 194 444 195 445
rect 193 444 194 445
rect 176 444 177 445
rect 175 444 176 445
rect 174 444 175 445
rect 155 444 156 445
rect 154 444 155 445
rect 199 445 200 446
rect 198 445 199 446
rect 197 445 198 446
rect 196 445 197 446
rect 195 445 196 446
rect 194 445 195 446
rect 193 445 194 446
rect 155 445 156 446
rect 154 445 155 446
rect 198 446 199 447
rect 197 446 198 447
rect 196 446 197 447
rect 194 446 195 447
rect 193 446 194 447
rect 198 447 199 448
rect 197 447 198 448
rect 196 447 197 448
rect 194 448 195 449
rect 193 448 194 449
rect 198 449 199 450
rect 197 449 198 450
rect 196 449 197 450
rect 195 449 196 450
rect 194 449 195 450
rect 193 449 194 450
rect 192 449 193 450
rect 199 450 200 451
rect 198 450 199 451
rect 197 450 198 451
rect 196 450 197 451
rect 195 450 196 451
rect 194 450 195 451
rect 193 450 194 451
rect 192 450 193 451
rect 191 450 192 451
rect 199 451 200 452
rect 198 451 199 452
rect 194 451 195 452
rect 193 451 194 452
rect 198 452 199 453
rect 198 453 199 454
rect 197 453 198 454
rect 196 453 197 454
rect 195 453 196 454
rect 194 453 195 454
rect 193 453 194 454
rect 191 453 192 454
rect 190 453 191 454
rect 199 454 200 455
rect 198 454 199 455
rect 197 454 198 455
rect 196 454 197 455
rect 195 454 196 455
rect 194 454 195 455
rect 193 454 194 455
rect 191 454 192 455
rect 190 454 191 455
rect 175 455 176 456
rect 174 455 175 456
rect 173 455 174 456
rect 151 455 152 456
rect 150 455 151 456
rect 149 455 150 456
rect 148 455 149 456
rect 147 455 148 456
rect 146 455 147 456
rect 145 455 146 456
rect 144 455 145 456
rect 143 455 144 456
rect 142 455 143 456
rect 141 455 142 456
rect 140 455 141 456
rect 139 455 140 456
rect 138 455 139 456
rect 137 455 138 456
rect 136 455 137 456
rect 135 455 136 456
rect 134 455 135 456
rect 133 455 134 456
rect 132 455 133 456
rect 131 455 132 456
rect 130 455 131 456
rect 129 455 130 456
rect 128 455 129 456
rect 127 455 128 456
rect 126 455 127 456
rect 125 455 126 456
rect 124 455 125 456
rect 123 455 124 456
rect 122 455 123 456
rect 121 455 122 456
rect 120 455 121 456
rect 119 455 120 456
rect 118 455 119 456
rect 117 455 118 456
rect 116 455 117 456
rect 115 455 116 456
rect 114 455 115 456
rect 113 455 114 456
rect 112 455 113 456
rect 111 455 112 456
rect 110 455 111 456
rect 109 455 110 456
rect 108 455 109 456
rect 107 455 108 456
rect 106 455 107 456
rect 105 455 106 456
rect 104 455 105 456
rect 194 456 195 457
rect 193 456 194 457
rect 175 456 176 457
rect 174 456 175 457
rect 173 456 174 457
rect 172 456 173 457
rect 151 456 152 457
rect 150 456 151 457
rect 149 456 150 457
rect 148 456 149 457
rect 147 456 148 457
rect 146 456 147 457
rect 145 456 146 457
rect 144 456 145 457
rect 143 456 144 457
rect 142 456 143 457
rect 141 456 142 457
rect 140 456 141 457
rect 139 456 140 457
rect 138 456 139 457
rect 137 456 138 457
rect 136 456 137 457
rect 135 456 136 457
rect 134 456 135 457
rect 133 456 134 457
rect 132 456 133 457
rect 131 456 132 457
rect 130 456 131 457
rect 129 456 130 457
rect 128 456 129 457
rect 127 456 128 457
rect 126 456 127 457
rect 125 456 126 457
rect 124 456 125 457
rect 123 456 124 457
rect 122 456 123 457
rect 121 456 122 457
rect 120 456 121 457
rect 119 456 120 457
rect 118 456 119 457
rect 117 456 118 457
rect 116 456 117 457
rect 115 456 116 457
rect 114 456 115 457
rect 113 456 114 457
rect 112 456 113 457
rect 111 456 112 457
rect 110 456 111 457
rect 109 456 110 457
rect 108 456 109 457
rect 107 456 108 457
rect 106 456 107 457
rect 105 456 106 457
rect 104 456 105 457
rect 198 457 199 458
rect 197 457 198 458
rect 196 457 197 458
rect 195 457 196 458
rect 194 457 195 458
rect 193 457 194 458
rect 192 457 193 458
rect 191 457 192 458
rect 175 457 176 458
rect 174 457 175 458
rect 173 457 174 458
rect 172 457 173 458
rect 169 457 170 458
rect 168 457 169 458
rect 167 457 168 458
rect 166 457 167 458
rect 151 457 152 458
rect 150 457 151 458
rect 149 457 150 458
rect 148 457 149 458
rect 147 457 148 458
rect 146 457 147 458
rect 145 457 146 458
rect 144 457 145 458
rect 143 457 144 458
rect 142 457 143 458
rect 141 457 142 458
rect 140 457 141 458
rect 139 457 140 458
rect 138 457 139 458
rect 137 457 138 458
rect 136 457 137 458
rect 135 457 136 458
rect 134 457 135 458
rect 133 457 134 458
rect 132 457 133 458
rect 131 457 132 458
rect 130 457 131 458
rect 129 457 130 458
rect 128 457 129 458
rect 127 457 128 458
rect 126 457 127 458
rect 125 457 126 458
rect 124 457 125 458
rect 123 457 124 458
rect 122 457 123 458
rect 121 457 122 458
rect 120 457 121 458
rect 119 457 120 458
rect 118 457 119 458
rect 117 457 118 458
rect 116 457 117 458
rect 115 457 116 458
rect 114 457 115 458
rect 113 457 114 458
rect 112 457 113 458
rect 111 457 112 458
rect 110 457 111 458
rect 109 457 110 458
rect 108 457 109 458
rect 107 457 108 458
rect 106 457 107 458
rect 105 457 106 458
rect 104 457 105 458
rect 199 458 200 459
rect 198 458 199 459
rect 197 458 198 459
rect 196 458 197 459
rect 195 458 196 459
rect 194 458 195 459
rect 193 458 194 459
rect 192 458 193 459
rect 191 458 192 459
rect 175 458 176 459
rect 174 458 175 459
rect 173 458 174 459
rect 172 458 173 459
rect 170 458 171 459
rect 169 458 170 459
rect 168 458 169 459
rect 167 458 168 459
rect 166 458 167 459
rect 165 458 166 459
rect 151 458 152 459
rect 150 458 151 459
rect 149 458 150 459
rect 148 458 149 459
rect 147 458 148 459
rect 146 458 147 459
rect 145 458 146 459
rect 144 458 145 459
rect 143 458 144 459
rect 142 458 143 459
rect 141 458 142 459
rect 140 458 141 459
rect 139 458 140 459
rect 138 458 139 459
rect 137 458 138 459
rect 136 458 137 459
rect 135 458 136 459
rect 134 458 135 459
rect 133 458 134 459
rect 132 458 133 459
rect 131 458 132 459
rect 130 458 131 459
rect 129 458 130 459
rect 128 458 129 459
rect 127 458 128 459
rect 126 458 127 459
rect 125 458 126 459
rect 124 458 125 459
rect 123 458 124 459
rect 122 458 123 459
rect 121 458 122 459
rect 120 458 121 459
rect 119 458 120 459
rect 118 458 119 459
rect 117 458 118 459
rect 116 458 117 459
rect 115 458 116 459
rect 114 458 115 459
rect 113 458 114 459
rect 112 458 113 459
rect 111 458 112 459
rect 110 458 111 459
rect 109 458 110 459
rect 108 458 109 459
rect 107 458 108 459
rect 106 458 107 459
rect 105 458 106 459
rect 104 458 105 459
rect 199 459 200 460
rect 198 459 199 460
rect 194 459 195 460
rect 193 459 194 460
rect 185 459 186 460
rect 184 459 185 460
rect 183 459 184 460
rect 182 459 183 460
rect 181 459 182 460
rect 180 459 181 460
rect 175 459 176 460
rect 174 459 175 460
rect 173 459 174 460
rect 172 459 173 460
rect 170 459 171 460
rect 169 459 170 460
rect 168 459 169 460
rect 167 459 168 460
rect 166 459 167 460
rect 165 459 166 460
rect 164 459 165 460
rect 151 459 152 460
rect 150 459 151 460
rect 149 459 150 460
rect 148 459 149 460
rect 147 459 148 460
rect 146 459 147 460
rect 145 459 146 460
rect 144 459 145 460
rect 143 459 144 460
rect 142 459 143 460
rect 141 459 142 460
rect 140 459 141 460
rect 139 459 140 460
rect 138 459 139 460
rect 137 459 138 460
rect 136 459 137 460
rect 135 459 136 460
rect 134 459 135 460
rect 133 459 134 460
rect 132 459 133 460
rect 131 459 132 460
rect 130 459 131 460
rect 129 459 130 460
rect 128 459 129 460
rect 127 459 128 460
rect 126 459 127 460
rect 125 459 126 460
rect 124 459 125 460
rect 123 459 124 460
rect 122 459 123 460
rect 121 459 122 460
rect 120 459 121 460
rect 119 459 120 460
rect 118 459 119 460
rect 117 459 118 460
rect 116 459 117 460
rect 115 459 116 460
rect 114 459 115 460
rect 113 459 114 460
rect 112 459 113 460
rect 111 459 112 460
rect 110 459 111 460
rect 109 459 110 460
rect 108 459 109 460
rect 107 459 108 460
rect 106 459 107 460
rect 105 459 106 460
rect 104 459 105 460
rect 198 460 199 461
rect 185 460 186 461
rect 184 460 185 461
rect 183 460 184 461
rect 182 460 183 461
rect 181 460 182 461
rect 180 460 181 461
rect 175 460 176 461
rect 174 460 175 461
rect 173 460 174 461
rect 172 460 173 461
rect 171 460 172 461
rect 170 460 171 461
rect 169 460 170 461
rect 168 460 169 461
rect 167 460 168 461
rect 166 460 167 461
rect 165 460 166 461
rect 164 460 165 461
rect 151 460 152 461
rect 150 460 151 461
rect 149 460 150 461
rect 148 460 149 461
rect 147 460 148 461
rect 146 460 147 461
rect 145 460 146 461
rect 144 460 145 461
rect 143 460 144 461
rect 142 460 143 461
rect 141 460 142 461
rect 140 460 141 461
rect 139 460 140 461
rect 138 460 139 461
rect 137 460 138 461
rect 136 460 137 461
rect 135 460 136 461
rect 134 460 135 461
rect 133 460 134 461
rect 132 460 133 461
rect 131 460 132 461
rect 130 460 131 461
rect 129 460 130 461
rect 128 460 129 461
rect 127 460 128 461
rect 126 460 127 461
rect 125 460 126 461
rect 124 460 125 461
rect 123 460 124 461
rect 122 460 123 461
rect 121 460 122 461
rect 120 460 121 461
rect 119 460 120 461
rect 118 460 119 461
rect 117 460 118 461
rect 116 460 117 461
rect 115 460 116 461
rect 114 460 115 461
rect 113 460 114 461
rect 112 460 113 461
rect 111 460 112 461
rect 110 460 111 461
rect 109 460 110 461
rect 108 460 109 461
rect 107 460 108 461
rect 106 460 107 461
rect 105 460 106 461
rect 104 460 105 461
rect 198 461 199 462
rect 197 461 198 462
rect 196 461 197 462
rect 195 461 196 462
rect 194 461 195 462
rect 193 461 194 462
rect 185 461 186 462
rect 184 461 185 462
rect 183 461 184 462
rect 182 461 183 462
rect 181 461 182 462
rect 180 461 181 462
rect 179 461 180 462
rect 178 461 179 462
rect 177 461 178 462
rect 176 461 177 462
rect 175 461 176 462
rect 174 461 175 462
rect 173 461 174 462
rect 172 461 173 462
rect 171 461 172 462
rect 170 461 171 462
rect 169 461 170 462
rect 168 461 169 462
rect 166 461 167 462
rect 165 461 166 462
rect 164 461 165 462
rect 163 461 164 462
rect 151 461 152 462
rect 150 461 151 462
rect 149 461 150 462
rect 148 461 149 462
rect 147 461 148 462
rect 146 461 147 462
rect 145 461 146 462
rect 144 461 145 462
rect 143 461 144 462
rect 142 461 143 462
rect 141 461 142 462
rect 140 461 141 462
rect 139 461 140 462
rect 138 461 139 462
rect 137 461 138 462
rect 136 461 137 462
rect 135 461 136 462
rect 134 461 135 462
rect 133 461 134 462
rect 132 461 133 462
rect 131 461 132 462
rect 130 461 131 462
rect 129 461 130 462
rect 128 461 129 462
rect 127 461 128 462
rect 126 461 127 462
rect 125 461 126 462
rect 124 461 125 462
rect 123 461 124 462
rect 122 461 123 462
rect 121 461 122 462
rect 120 461 121 462
rect 119 461 120 462
rect 118 461 119 462
rect 117 461 118 462
rect 116 461 117 462
rect 115 461 116 462
rect 114 461 115 462
rect 113 461 114 462
rect 112 461 113 462
rect 111 461 112 462
rect 110 461 111 462
rect 109 461 110 462
rect 108 461 109 462
rect 107 461 108 462
rect 106 461 107 462
rect 105 461 106 462
rect 104 461 105 462
rect 199 462 200 463
rect 198 462 199 463
rect 197 462 198 463
rect 196 462 197 463
rect 195 462 196 463
rect 194 462 195 463
rect 193 462 194 463
rect 185 462 186 463
rect 184 462 185 463
rect 183 462 184 463
rect 182 462 183 463
rect 181 462 182 463
rect 180 462 181 463
rect 179 462 180 463
rect 178 462 179 463
rect 177 462 178 463
rect 176 462 177 463
rect 175 462 176 463
rect 174 462 175 463
rect 173 462 174 463
rect 172 462 173 463
rect 171 462 172 463
rect 170 462 171 463
rect 169 462 170 463
rect 165 462 166 463
rect 164 462 165 463
rect 163 462 164 463
rect 151 462 152 463
rect 150 462 151 463
rect 149 462 150 463
rect 148 462 149 463
rect 147 462 148 463
rect 146 462 147 463
rect 145 462 146 463
rect 144 462 145 463
rect 143 462 144 463
rect 142 462 143 463
rect 141 462 142 463
rect 140 462 141 463
rect 139 462 140 463
rect 138 462 139 463
rect 137 462 138 463
rect 136 462 137 463
rect 135 462 136 463
rect 134 462 135 463
rect 133 462 134 463
rect 132 462 133 463
rect 131 462 132 463
rect 130 462 131 463
rect 129 462 130 463
rect 128 462 129 463
rect 127 462 128 463
rect 126 462 127 463
rect 125 462 126 463
rect 124 462 125 463
rect 123 462 124 463
rect 122 462 123 463
rect 121 462 122 463
rect 120 462 121 463
rect 119 462 120 463
rect 118 462 119 463
rect 117 462 118 463
rect 116 462 117 463
rect 115 462 116 463
rect 114 462 115 463
rect 113 462 114 463
rect 112 462 113 463
rect 111 462 112 463
rect 110 462 111 463
rect 109 462 110 463
rect 108 462 109 463
rect 107 462 108 463
rect 106 462 107 463
rect 105 462 106 463
rect 104 462 105 463
rect 199 463 200 464
rect 198 463 199 464
rect 185 463 186 464
rect 184 463 185 464
rect 183 463 184 464
rect 182 463 183 464
rect 178 463 179 464
rect 177 463 178 464
rect 176 463 177 464
rect 175 463 176 464
rect 174 463 175 464
rect 173 463 174 464
rect 172 463 173 464
rect 171 463 172 464
rect 170 463 171 464
rect 169 463 170 464
rect 165 463 166 464
rect 164 463 165 464
rect 163 463 164 464
rect 151 463 152 464
rect 150 463 151 464
rect 149 463 150 464
rect 148 463 149 464
rect 147 463 148 464
rect 146 463 147 464
rect 145 463 146 464
rect 144 463 145 464
rect 143 463 144 464
rect 142 463 143 464
rect 141 463 142 464
rect 140 463 141 464
rect 139 463 140 464
rect 138 463 139 464
rect 137 463 138 464
rect 136 463 137 464
rect 135 463 136 464
rect 134 463 135 464
rect 133 463 134 464
rect 132 463 133 464
rect 131 463 132 464
rect 130 463 131 464
rect 129 463 130 464
rect 128 463 129 464
rect 127 463 128 464
rect 126 463 127 464
rect 125 463 126 464
rect 124 463 125 464
rect 123 463 124 464
rect 122 463 123 464
rect 121 463 122 464
rect 120 463 121 464
rect 119 463 120 464
rect 118 463 119 464
rect 117 463 118 464
rect 116 463 117 464
rect 115 463 116 464
rect 114 463 115 464
rect 113 463 114 464
rect 112 463 113 464
rect 111 463 112 464
rect 110 463 111 464
rect 109 463 110 464
rect 108 463 109 464
rect 107 463 108 464
rect 106 463 107 464
rect 105 463 106 464
rect 104 463 105 464
rect 198 464 199 465
rect 185 464 186 465
rect 184 464 185 465
rect 183 464 184 465
rect 182 464 183 465
rect 175 464 176 465
rect 174 464 175 465
rect 173 464 174 465
rect 172 464 173 465
rect 171 464 172 465
rect 170 464 171 465
rect 169 464 170 465
rect 165 464 166 465
rect 164 464 165 465
rect 163 464 164 465
rect 151 464 152 465
rect 150 464 151 465
rect 149 464 150 465
rect 148 464 149 465
rect 147 464 148 465
rect 146 464 147 465
rect 145 464 146 465
rect 144 464 145 465
rect 143 464 144 465
rect 142 464 143 465
rect 141 464 142 465
rect 140 464 141 465
rect 139 464 140 465
rect 138 464 139 465
rect 137 464 138 465
rect 136 464 137 465
rect 135 464 136 465
rect 134 464 135 465
rect 133 464 134 465
rect 132 464 133 465
rect 131 464 132 465
rect 130 464 131 465
rect 129 464 130 465
rect 128 464 129 465
rect 127 464 128 465
rect 126 464 127 465
rect 125 464 126 465
rect 124 464 125 465
rect 123 464 124 465
rect 122 464 123 465
rect 121 464 122 465
rect 120 464 121 465
rect 119 464 120 465
rect 118 464 119 465
rect 117 464 118 465
rect 116 464 117 465
rect 115 464 116 465
rect 114 464 115 465
rect 113 464 114 465
rect 112 464 113 465
rect 111 464 112 465
rect 110 464 111 465
rect 109 464 110 465
rect 108 464 109 465
rect 107 464 108 465
rect 106 464 107 465
rect 105 464 106 465
rect 104 464 105 465
rect 199 465 200 466
rect 198 465 199 466
rect 197 465 198 466
rect 196 465 197 466
rect 195 465 196 466
rect 194 465 195 466
rect 193 465 194 466
rect 185 465 186 466
rect 184 465 185 466
rect 183 465 184 466
rect 182 465 183 466
rect 175 465 176 466
rect 174 465 175 466
rect 173 465 174 466
rect 172 465 173 466
rect 171 465 172 466
rect 170 465 171 466
rect 169 465 170 466
rect 165 465 166 466
rect 164 465 165 466
rect 163 465 164 466
rect 151 465 152 466
rect 150 465 151 466
rect 149 465 150 466
rect 148 465 149 466
rect 147 465 148 466
rect 146 465 147 466
rect 145 465 146 466
rect 144 465 145 466
rect 143 465 144 466
rect 142 465 143 466
rect 141 465 142 466
rect 140 465 141 466
rect 139 465 140 466
rect 138 465 139 466
rect 137 465 138 466
rect 136 465 137 466
rect 135 465 136 466
rect 134 465 135 466
rect 133 465 134 466
rect 132 465 133 466
rect 131 465 132 466
rect 130 465 131 466
rect 129 465 130 466
rect 128 465 129 466
rect 127 465 128 466
rect 126 465 127 466
rect 125 465 126 466
rect 124 465 125 466
rect 123 465 124 466
rect 122 465 123 466
rect 121 465 122 466
rect 120 465 121 466
rect 119 465 120 466
rect 118 465 119 466
rect 117 465 118 466
rect 116 465 117 466
rect 115 465 116 466
rect 114 465 115 466
rect 113 465 114 466
rect 112 465 113 466
rect 111 465 112 466
rect 110 465 111 466
rect 109 465 110 466
rect 108 465 109 466
rect 107 465 108 466
rect 106 465 107 466
rect 105 465 106 466
rect 104 465 105 466
rect 198 466 199 467
rect 197 466 198 467
rect 196 466 197 467
rect 195 466 196 467
rect 194 466 195 467
rect 193 466 194 467
rect 185 466 186 467
rect 184 466 185 467
rect 183 466 184 467
rect 182 466 183 467
rect 175 466 176 467
rect 174 466 175 467
rect 173 466 174 467
rect 172 466 173 467
rect 171 466 172 467
rect 170 466 171 467
rect 169 466 170 467
rect 168 466 169 467
rect 166 466 167 467
rect 165 466 166 467
rect 164 466 165 467
rect 151 466 152 467
rect 150 466 151 467
rect 149 466 150 467
rect 148 466 149 467
rect 147 466 148 467
rect 146 466 147 467
rect 145 466 146 467
rect 144 466 145 467
rect 143 466 144 467
rect 142 466 143 467
rect 141 466 142 467
rect 140 466 141 467
rect 139 466 140 467
rect 138 466 139 467
rect 137 466 138 467
rect 136 466 137 467
rect 135 466 136 467
rect 134 466 135 467
rect 133 466 134 467
rect 132 466 133 467
rect 131 466 132 467
rect 130 466 131 467
rect 129 466 130 467
rect 128 466 129 467
rect 127 466 128 467
rect 126 466 127 467
rect 125 466 126 467
rect 124 466 125 467
rect 123 466 124 467
rect 122 466 123 467
rect 121 466 122 467
rect 120 466 121 467
rect 119 466 120 467
rect 118 466 119 467
rect 117 466 118 467
rect 116 466 117 467
rect 115 466 116 467
rect 114 466 115 467
rect 113 466 114 467
rect 112 466 113 467
rect 111 466 112 467
rect 110 466 111 467
rect 109 466 110 467
rect 108 466 109 467
rect 107 466 108 467
rect 106 466 107 467
rect 105 466 106 467
rect 104 466 105 467
rect 185 467 186 468
rect 184 467 185 468
rect 183 467 184 468
rect 182 467 183 468
rect 175 467 176 468
rect 174 467 175 468
rect 173 467 174 468
rect 172 467 173 468
rect 170 467 171 468
rect 169 467 170 468
rect 168 467 169 468
rect 167 467 168 468
rect 166 467 167 468
rect 165 467 166 468
rect 164 467 165 468
rect 151 467 152 468
rect 150 467 151 468
rect 149 467 150 468
rect 148 467 149 468
rect 147 467 148 468
rect 146 467 147 468
rect 145 467 146 468
rect 144 467 145 468
rect 143 467 144 468
rect 142 467 143 468
rect 141 467 142 468
rect 140 467 141 468
rect 139 467 140 468
rect 138 467 139 468
rect 137 467 138 468
rect 136 467 137 468
rect 135 467 136 468
rect 134 467 135 468
rect 133 467 134 468
rect 132 467 133 468
rect 131 467 132 468
rect 130 467 131 468
rect 129 467 130 468
rect 128 467 129 468
rect 127 467 128 468
rect 126 467 127 468
rect 125 467 126 468
rect 124 467 125 468
rect 123 467 124 468
rect 122 467 123 468
rect 121 467 122 468
rect 120 467 121 468
rect 119 467 120 468
rect 118 467 119 468
rect 117 467 118 468
rect 116 467 117 468
rect 115 467 116 468
rect 114 467 115 468
rect 113 467 114 468
rect 112 467 113 468
rect 111 467 112 468
rect 110 467 111 468
rect 109 467 110 468
rect 108 467 109 468
rect 107 467 108 468
rect 106 467 107 468
rect 105 467 106 468
rect 104 467 105 468
rect 197 468 198 469
rect 196 468 197 469
rect 195 468 196 469
rect 194 468 195 469
rect 193 468 194 469
rect 192 468 193 469
rect 185 468 186 469
rect 184 468 185 469
rect 183 468 184 469
rect 182 468 183 469
rect 178 468 179 469
rect 177 468 178 469
rect 176 468 177 469
rect 175 468 176 469
rect 174 468 175 469
rect 173 468 174 469
rect 172 468 173 469
rect 170 468 171 469
rect 169 468 170 469
rect 168 468 169 469
rect 167 468 168 469
rect 166 468 167 469
rect 165 468 166 469
rect 151 468 152 469
rect 150 468 151 469
rect 149 468 150 469
rect 148 468 149 469
rect 147 468 148 469
rect 146 468 147 469
rect 145 468 146 469
rect 144 468 145 469
rect 143 468 144 469
rect 142 468 143 469
rect 141 468 142 469
rect 140 468 141 469
rect 139 468 140 469
rect 138 468 139 469
rect 137 468 138 469
rect 136 468 137 469
rect 135 468 136 469
rect 134 468 135 469
rect 133 468 134 469
rect 132 468 133 469
rect 131 468 132 469
rect 130 468 131 469
rect 129 468 130 469
rect 128 468 129 469
rect 127 468 128 469
rect 126 468 127 469
rect 125 468 126 469
rect 124 468 125 469
rect 123 468 124 469
rect 122 468 123 469
rect 121 468 122 469
rect 120 468 121 469
rect 119 468 120 469
rect 118 468 119 469
rect 117 468 118 469
rect 116 468 117 469
rect 115 468 116 469
rect 114 468 115 469
rect 113 468 114 469
rect 112 468 113 469
rect 111 468 112 469
rect 110 468 111 469
rect 109 468 110 469
rect 108 468 109 469
rect 107 468 108 469
rect 106 468 107 469
rect 105 468 106 469
rect 104 468 105 469
rect 198 469 199 470
rect 197 469 198 470
rect 196 469 197 470
rect 195 469 196 470
rect 194 469 195 470
rect 193 469 194 470
rect 192 469 193 470
rect 191 469 192 470
rect 185 469 186 470
rect 184 469 185 470
rect 183 469 184 470
rect 182 469 183 470
rect 178 469 179 470
rect 177 469 178 470
rect 176 469 177 470
rect 175 469 176 470
rect 174 469 175 470
rect 173 469 174 470
rect 172 469 173 470
rect 169 469 170 470
rect 168 469 169 470
rect 167 469 168 470
rect 166 469 167 470
rect 165 469 166 470
rect 151 469 152 470
rect 150 469 151 470
rect 149 469 150 470
rect 148 469 149 470
rect 147 469 148 470
rect 146 469 147 470
rect 145 469 146 470
rect 144 469 145 470
rect 143 469 144 470
rect 142 469 143 470
rect 141 469 142 470
rect 140 469 141 470
rect 139 469 140 470
rect 138 469 139 470
rect 137 469 138 470
rect 136 469 137 470
rect 135 469 136 470
rect 134 469 135 470
rect 133 469 134 470
rect 132 469 133 470
rect 131 469 132 470
rect 130 469 131 470
rect 129 469 130 470
rect 128 469 129 470
rect 127 469 128 470
rect 126 469 127 470
rect 125 469 126 470
rect 124 469 125 470
rect 123 469 124 470
rect 122 469 123 470
rect 121 469 122 470
rect 120 469 121 470
rect 119 469 120 470
rect 118 469 119 470
rect 117 469 118 470
rect 116 469 117 470
rect 115 469 116 470
rect 114 469 115 470
rect 113 469 114 470
rect 112 469 113 470
rect 111 469 112 470
rect 110 469 111 470
rect 109 469 110 470
rect 108 469 109 470
rect 107 469 108 470
rect 106 469 107 470
rect 105 469 106 470
rect 104 469 105 470
rect 198 470 199 471
rect 197 470 198 471
rect 196 470 197 471
rect 195 470 196 471
rect 194 470 195 471
rect 193 470 194 471
rect 192 470 193 471
rect 191 470 192 471
rect 185 470 186 471
rect 184 470 185 471
rect 183 470 184 471
rect 182 470 183 471
rect 178 470 179 471
rect 177 470 178 471
rect 176 470 177 471
rect 175 470 176 471
rect 174 470 175 471
rect 173 470 174 471
rect 172 470 173 471
rect 168 470 169 471
rect 167 470 168 471
rect 166 470 167 471
rect 151 470 152 471
rect 150 470 151 471
rect 149 470 150 471
rect 148 470 149 471
rect 147 470 148 471
rect 146 470 147 471
rect 145 470 146 471
rect 144 470 145 471
rect 143 470 144 471
rect 142 470 143 471
rect 141 470 142 471
rect 140 470 141 471
rect 139 470 140 471
rect 138 470 139 471
rect 137 470 138 471
rect 136 470 137 471
rect 135 470 136 471
rect 134 470 135 471
rect 133 470 134 471
rect 132 470 133 471
rect 131 470 132 471
rect 130 470 131 471
rect 129 470 130 471
rect 128 470 129 471
rect 127 470 128 471
rect 126 470 127 471
rect 125 470 126 471
rect 124 470 125 471
rect 123 470 124 471
rect 122 470 123 471
rect 121 470 122 471
rect 120 470 121 471
rect 119 470 120 471
rect 118 470 119 471
rect 117 470 118 471
rect 116 470 117 471
rect 115 470 116 471
rect 114 470 115 471
rect 113 470 114 471
rect 112 470 113 471
rect 111 470 112 471
rect 110 470 111 471
rect 109 470 110 471
rect 108 470 109 471
rect 107 470 108 471
rect 106 470 107 471
rect 105 470 106 471
rect 104 470 105 471
rect 199 471 200 472
rect 198 471 199 472
rect 194 471 195 472
rect 193 471 194 472
rect 185 471 186 472
rect 184 471 185 472
rect 183 471 184 472
rect 182 471 183 472
rect 178 471 179 472
rect 177 471 178 472
rect 176 471 177 472
rect 174 471 175 472
rect 173 471 174 472
rect 172 471 173 472
rect 151 471 152 472
rect 150 471 151 472
rect 149 471 150 472
rect 148 471 149 472
rect 147 471 148 472
rect 146 471 147 472
rect 145 471 146 472
rect 144 471 145 472
rect 143 471 144 472
rect 142 471 143 472
rect 141 471 142 472
rect 140 471 141 472
rect 139 471 140 472
rect 138 471 139 472
rect 137 471 138 472
rect 136 471 137 472
rect 135 471 136 472
rect 134 471 135 472
rect 133 471 134 472
rect 132 471 133 472
rect 131 471 132 472
rect 130 471 131 472
rect 129 471 130 472
rect 128 471 129 472
rect 127 471 128 472
rect 126 471 127 472
rect 125 471 126 472
rect 124 471 125 472
rect 123 471 124 472
rect 122 471 123 472
rect 121 471 122 472
rect 120 471 121 472
rect 119 471 120 472
rect 118 471 119 472
rect 117 471 118 472
rect 116 471 117 472
rect 115 471 116 472
rect 114 471 115 472
rect 113 471 114 472
rect 112 471 113 472
rect 111 471 112 472
rect 110 471 111 472
rect 109 471 110 472
rect 108 471 109 472
rect 107 471 108 472
rect 106 471 107 472
rect 105 471 106 472
rect 104 471 105 472
rect 197 472 198 473
rect 196 472 197 473
rect 195 472 196 473
rect 185 472 186 473
rect 184 472 185 473
rect 183 472 184 473
rect 182 472 183 473
rect 178 472 179 473
rect 177 472 178 473
rect 176 472 177 473
rect 174 472 175 473
rect 173 472 174 473
rect 172 472 173 473
rect 151 472 152 473
rect 150 472 151 473
rect 149 472 150 473
rect 148 472 149 473
rect 147 472 148 473
rect 146 472 147 473
rect 145 472 146 473
rect 144 472 145 473
rect 143 472 144 473
rect 142 472 143 473
rect 141 472 142 473
rect 140 472 141 473
rect 139 472 140 473
rect 138 472 139 473
rect 137 472 138 473
rect 136 472 137 473
rect 135 472 136 473
rect 134 472 135 473
rect 133 472 134 473
rect 132 472 133 473
rect 131 472 132 473
rect 130 472 131 473
rect 129 472 130 473
rect 128 472 129 473
rect 127 472 128 473
rect 126 472 127 473
rect 125 472 126 473
rect 124 472 125 473
rect 123 472 124 473
rect 122 472 123 473
rect 121 472 122 473
rect 120 472 121 473
rect 119 472 120 473
rect 118 472 119 473
rect 117 472 118 473
rect 116 472 117 473
rect 115 472 116 473
rect 114 472 115 473
rect 113 472 114 473
rect 112 472 113 473
rect 111 472 112 473
rect 110 472 111 473
rect 109 472 110 473
rect 108 472 109 473
rect 107 472 108 473
rect 106 472 107 473
rect 105 472 106 473
rect 104 472 105 473
rect 198 473 199 474
rect 197 473 198 474
rect 196 473 197 474
rect 195 473 196 474
rect 194 473 195 474
rect 193 473 194 474
rect 185 473 186 474
rect 184 473 185 474
rect 183 473 184 474
rect 182 473 183 474
rect 178 473 179 474
rect 177 473 178 474
rect 176 473 177 474
rect 175 473 176 474
rect 151 473 152 474
rect 150 473 151 474
rect 149 473 150 474
rect 148 473 149 474
rect 147 473 148 474
rect 146 473 147 474
rect 145 473 146 474
rect 144 473 145 474
rect 143 473 144 474
rect 142 473 143 474
rect 141 473 142 474
rect 140 473 141 474
rect 139 473 140 474
rect 138 473 139 474
rect 137 473 138 474
rect 136 473 137 474
rect 135 473 136 474
rect 134 473 135 474
rect 133 473 134 474
rect 132 473 133 474
rect 131 473 132 474
rect 130 473 131 474
rect 129 473 130 474
rect 128 473 129 474
rect 127 473 128 474
rect 126 473 127 474
rect 125 473 126 474
rect 124 473 125 474
rect 123 473 124 474
rect 122 473 123 474
rect 121 473 122 474
rect 120 473 121 474
rect 119 473 120 474
rect 118 473 119 474
rect 117 473 118 474
rect 116 473 117 474
rect 115 473 116 474
rect 114 473 115 474
rect 113 473 114 474
rect 112 473 113 474
rect 111 473 112 474
rect 110 473 111 474
rect 109 473 110 474
rect 108 473 109 474
rect 107 473 108 474
rect 106 473 107 474
rect 105 473 106 474
rect 104 473 105 474
rect 198 474 199 475
rect 197 474 198 475
rect 196 474 197 475
rect 195 474 196 475
rect 194 474 195 475
rect 193 474 194 475
rect 185 474 186 475
rect 184 474 185 475
rect 183 474 184 475
rect 182 474 183 475
rect 180 474 181 475
rect 179 474 180 475
rect 178 474 179 475
rect 177 474 178 475
rect 176 474 177 475
rect 175 474 176 475
rect 174 474 175 475
rect 173 474 174 475
rect 172 474 173 475
rect 171 474 172 475
rect 170 474 171 475
rect 169 474 170 475
rect 168 474 169 475
rect 167 474 168 475
rect 166 474 167 475
rect 165 474 166 475
rect 164 474 165 475
rect 151 474 152 475
rect 150 474 151 475
rect 149 474 150 475
rect 148 474 149 475
rect 147 474 148 475
rect 146 474 147 475
rect 145 474 146 475
rect 144 474 145 475
rect 143 474 144 475
rect 142 474 143 475
rect 141 474 142 475
rect 140 474 141 475
rect 139 474 140 475
rect 138 474 139 475
rect 137 474 138 475
rect 136 474 137 475
rect 135 474 136 475
rect 134 474 135 475
rect 133 474 134 475
rect 132 474 133 475
rect 131 474 132 475
rect 130 474 131 475
rect 129 474 130 475
rect 128 474 129 475
rect 127 474 128 475
rect 126 474 127 475
rect 125 474 126 475
rect 124 474 125 475
rect 123 474 124 475
rect 122 474 123 475
rect 121 474 122 475
rect 120 474 121 475
rect 119 474 120 475
rect 118 474 119 475
rect 117 474 118 475
rect 116 474 117 475
rect 115 474 116 475
rect 114 474 115 475
rect 113 474 114 475
rect 112 474 113 475
rect 111 474 112 475
rect 110 474 111 475
rect 109 474 110 475
rect 108 474 109 475
rect 107 474 108 475
rect 106 474 107 475
rect 105 474 106 475
rect 104 474 105 475
rect 199 475 200 476
rect 198 475 199 476
rect 196 475 197 476
rect 194 475 195 476
rect 193 475 194 476
rect 185 475 186 476
rect 184 475 185 476
rect 183 475 184 476
rect 182 475 183 476
rect 180 475 181 476
rect 179 475 180 476
rect 178 475 179 476
rect 177 475 178 476
rect 176 475 177 476
rect 175 475 176 476
rect 174 475 175 476
rect 173 475 174 476
rect 172 475 173 476
rect 171 475 172 476
rect 170 475 171 476
rect 169 475 170 476
rect 168 475 169 476
rect 167 475 168 476
rect 166 475 167 476
rect 165 475 166 476
rect 164 475 165 476
rect 151 475 152 476
rect 150 475 151 476
rect 149 475 150 476
rect 148 475 149 476
rect 147 475 148 476
rect 146 475 147 476
rect 145 475 146 476
rect 144 475 145 476
rect 143 475 144 476
rect 142 475 143 476
rect 141 475 142 476
rect 140 475 141 476
rect 139 475 140 476
rect 138 475 139 476
rect 137 475 138 476
rect 136 475 137 476
rect 135 475 136 476
rect 134 475 135 476
rect 133 475 134 476
rect 132 475 133 476
rect 131 475 132 476
rect 130 475 131 476
rect 129 475 130 476
rect 128 475 129 476
rect 127 475 128 476
rect 126 475 127 476
rect 125 475 126 476
rect 124 475 125 476
rect 123 475 124 476
rect 122 475 123 476
rect 121 475 122 476
rect 120 475 121 476
rect 119 475 120 476
rect 118 475 119 476
rect 117 475 118 476
rect 116 475 117 476
rect 115 475 116 476
rect 114 475 115 476
rect 113 475 114 476
rect 112 475 113 476
rect 111 475 112 476
rect 110 475 111 476
rect 109 475 110 476
rect 108 475 109 476
rect 107 475 108 476
rect 106 475 107 476
rect 105 475 106 476
rect 104 475 105 476
rect 199 476 200 477
rect 198 476 199 477
rect 196 476 197 477
rect 195 476 196 477
rect 194 476 195 477
rect 193 476 194 477
rect 185 476 186 477
rect 184 476 185 477
rect 183 476 184 477
rect 182 476 183 477
rect 180 476 181 477
rect 179 476 180 477
rect 178 476 179 477
rect 177 476 178 477
rect 176 476 177 477
rect 175 476 176 477
rect 174 476 175 477
rect 173 476 174 477
rect 172 476 173 477
rect 171 476 172 477
rect 170 476 171 477
rect 169 476 170 477
rect 168 476 169 477
rect 167 476 168 477
rect 166 476 167 477
rect 165 476 166 477
rect 164 476 165 477
rect 151 476 152 477
rect 150 476 151 477
rect 149 476 150 477
rect 148 476 149 477
rect 147 476 148 477
rect 146 476 147 477
rect 145 476 146 477
rect 144 476 145 477
rect 143 476 144 477
rect 142 476 143 477
rect 141 476 142 477
rect 140 476 141 477
rect 139 476 140 477
rect 138 476 139 477
rect 137 476 138 477
rect 136 476 137 477
rect 135 476 136 477
rect 134 476 135 477
rect 133 476 134 477
rect 132 476 133 477
rect 131 476 132 477
rect 130 476 131 477
rect 129 476 130 477
rect 128 476 129 477
rect 127 476 128 477
rect 126 476 127 477
rect 125 476 126 477
rect 124 476 125 477
rect 123 476 124 477
rect 122 476 123 477
rect 121 476 122 477
rect 120 476 121 477
rect 119 476 120 477
rect 118 476 119 477
rect 117 476 118 477
rect 116 476 117 477
rect 115 476 116 477
rect 114 476 115 477
rect 113 476 114 477
rect 112 476 113 477
rect 111 476 112 477
rect 110 476 111 477
rect 109 476 110 477
rect 108 476 109 477
rect 107 476 108 477
rect 106 476 107 477
rect 105 476 106 477
rect 104 476 105 477
rect 198 477 199 478
rect 196 477 197 478
rect 195 477 196 478
rect 194 477 195 478
rect 193 477 194 478
rect 184 477 185 478
rect 183 477 184 478
rect 182 477 183 478
rect 179 477 180 478
rect 178 477 179 478
rect 177 477 178 478
rect 176 477 177 478
rect 175 477 176 478
rect 174 477 175 478
rect 173 477 174 478
rect 172 477 173 478
rect 171 477 172 478
rect 170 477 171 478
rect 169 477 170 478
rect 168 477 169 478
rect 167 477 168 478
rect 166 477 167 478
rect 165 477 166 478
rect 164 477 165 478
rect 151 477 152 478
rect 150 477 151 478
rect 149 477 150 478
rect 148 477 149 478
rect 147 477 148 478
rect 146 477 147 478
rect 145 477 146 478
rect 144 477 145 478
rect 143 477 144 478
rect 142 477 143 478
rect 141 477 142 478
rect 140 477 141 478
rect 139 477 140 478
rect 138 477 139 478
rect 137 477 138 478
rect 136 477 137 478
rect 135 477 136 478
rect 134 477 135 478
rect 133 477 134 478
rect 132 477 133 478
rect 131 477 132 478
rect 130 477 131 478
rect 129 477 130 478
rect 128 477 129 478
rect 127 477 128 478
rect 126 477 127 478
rect 125 477 126 478
rect 124 477 125 478
rect 123 477 124 478
rect 122 477 123 478
rect 121 477 122 478
rect 120 477 121 478
rect 119 477 120 478
rect 118 477 119 478
rect 117 477 118 478
rect 116 477 117 478
rect 115 477 116 478
rect 114 477 115 478
rect 113 477 114 478
rect 112 477 113 478
rect 111 477 112 478
rect 110 477 111 478
rect 109 477 110 478
rect 108 477 109 478
rect 107 477 108 478
rect 106 477 107 478
rect 105 477 106 478
rect 104 477 105 478
rect 196 478 197 479
rect 151 478 152 479
rect 150 478 151 479
rect 149 478 150 479
rect 148 478 149 479
rect 147 478 148 479
rect 146 478 147 479
rect 145 478 146 479
rect 144 478 145 479
rect 143 478 144 479
rect 142 478 143 479
rect 141 478 142 479
rect 140 478 141 479
rect 139 478 140 479
rect 138 478 139 479
rect 137 478 138 479
rect 136 478 137 479
rect 135 478 136 479
rect 134 478 135 479
rect 133 478 134 479
rect 132 478 133 479
rect 131 478 132 479
rect 130 478 131 479
rect 129 478 130 479
rect 128 478 129 479
rect 127 478 128 479
rect 126 478 127 479
rect 125 478 126 479
rect 124 478 125 479
rect 123 478 124 479
rect 122 478 123 479
rect 121 478 122 479
rect 120 478 121 479
rect 119 478 120 479
rect 118 478 119 479
rect 117 478 118 479
rect 116 478 117 479
rect 115 478 116 479
rect 114 478 115 479
rect 113 478 114 479
rect 112 478 113 479
rect 111 478 112 479
rect 110 478 111 479
rect 109 478 110 479
rect 108 478 109 479
rect 107 478 108 479
rect 106 478 107 479
rect 105 478 106 479
rect 104 478 105 479
<< end >>
