magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -56 -56 162 162
<< diffusion >>
rect 5 5 101 101
<< genericcontact >>
rect 22 78 28 84
rect 50 78 56 84
rect 78 78 84 84
rect 22 50 28 56
rect 50 50 56 56
rect 78 50 84 56
rect 22 22 28 28
rect 50 22 56 28
rect 78 22 84 28
<< metal1 >>
rect 4 4 102 102
<< end >>
