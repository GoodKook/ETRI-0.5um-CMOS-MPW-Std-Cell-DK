magic
tech scmos
magscale 1 2
timestamp 1738238709
<< nwell >>
rect -2 4224 4782 4436
rect 2169 4220 2205 4224
rect -2 3744 4782 3956
rect 655 3740 691 3744
rect -3 3264 4782 3476
rect -3 2784 4782 2996
rect -3 2304 4782 2516
rect 875 2036 911 2040
rect -2 1942 4782 2036
rect -3 1824 4782 1942
rect -2 1462 4782 1556
rect -3 1344 4782 1462
rect 515 1076 551 1080
rect 3229 1076 3265 1080
rect -2 982 4782 1076
rect -3 864 4782 982
rect 3229 860 3265 864
rect 1069 596 1105 600
rect 2535 596 2571 600
rect -3 384 4782 596
rect 595 116 631 120
rect 3115 116 3151 120
rect -3 -2 4782 116
<< ntransistor >>
rect 43 4516 47 4556
rect 65 4536 69 4556
rect 133 4516 137 4556
rect 143 4516 147 4556
rect 205 4516 209 4556
rect 225 4516 229 4556
rect 245 4516 249 4556
rect 291 4536 295 4556
rect 313 4516 317 4556
rect 385 4536 389 4556
rect 405 4536 409 4556
rect 465 4536 469 4556
rect 485 4536 489 4556
rect 531 4536 535 4556
rect 553 4516 557 4556
rect 625 4536 629 4556
rect 671 4536 675 4556
rect 691 4536 695 4556
rect 751 4536 755 4556
rect 811 4516 815 4556
rect 833 4536 837 4556
rect 843 4536 847 4556
rect 863 4536 867 4556
rect 871 4536 875 4556
rect 917 4536 921 4556
rect 939 4536 943 4556
rect 949 4536 953 4556
rect 971 4536 975 4556
rect 981 4536 985 4556
rect 1001 4516 1005 4556
rect 1051 4516 1055 4556
rect 1071 4516 1075 4556
rect 1091 4516 1095 4556
rect 1151 4516 1155 4556
rect 1173 4536 1177 4556
rect 1183 4536 1187 4556
rect 1203 4536 1207 4556
rect 1211 4536 1215 4556
rect 1257 4536 1261 4556
rect 1279 4536 1283 4556
rect 1289 4536 1293 4556
rect 1311 4536 1315 4556
rect 1321 4536 1325 4556
rect 1341 4516 1345 4556
rect 1391 4516 1395 4556
rect 1411 4516 1415 4556
rect 1431 4516 1435 4556
rect 1495 4516 1499 4556
rect 1515 4536 1519 4556
rect 1525 4536 1529 4556
rect 1547 4536 1551 4556
rect 1557 4536 1561 4556
rect 1579 4536 1583 4556
rect 1625 4536 1629 4556
rect 1633 4536 1637 4556
rect 1653 4536 1657 4556
rect 1663 4536 1667 4556
rect 1685 4516 1689 4556
rect 1733 4516 1737 4556
rect 1743 4516 1747 4556
rect 1811 4516 1815 4556
rect 1833 4536 1837 4556
rect 1843 4536 1847 4556
rect 1863 4536 1867 4556
rect 1871 4536 1875 4556
rect 1917 4536 1921 4556
rect 1939 4536 1943 4556
rect 1949 4536 1953 4556
rect 1971 4536 1975 4556
rect 1981 4536 1985 4556
rect 2001 4516 2005 4556
rect 2051 4516 2055 4556
rect 2071 4516 2075 4556
rect 2091 4516 2095 4556
rect 2111 4516 2115 4556
rect 2208 4496 2212 4556
rect 2216 4496 2220 4556
rect 2224 4496 2228 4556
rect 2285 4516 2289 4556
rect 2305 4516 2309 4556
rect 2325 4516 2329 4556
rect 2385 4536 2389 4556
rect 2431 4536 2435 4556
rect 2451 4536 2455 4556
rect 2525 4536 2529 4556
rect 2571 4516 2575 4556
rect 2591 4516 2595 4556
rect 2611 4516 2615 4556
rect 2671 4536 2675 4556
rect 2693 4516 2697 4556
rect 2751 4536 2755 4556
rect 2773 4516 2777 4556
rect 2843 4516 2847 4556
rect 2865 4536 2869 4556
rect 2948 4496 2952 4556
rect 2956 4496 2960 4556
rect 2964 4496 2968 4556
rect 3035 4516 3039 4556
rect 3055 4516 3059 4556
rect 3065 4516 3069 4556
rect 3123 4516 3127 4556
rect 3145 4536 3149 4556
rect 3228 4496 3232 4556
rect 3236 4496 3240 4556
rect 3244 4496 3248 4556
rect 3293 4516 3297 4556
rect 3303 4516 3307 4556
rect 3374 4516 3378 4556
rect 3382 4516 3386 4556
rect 3404 4536 3408 4556
rect 3471 4536 3475 4556
rect 3533 4516 3537 4556
rect 3543 4516 3547 4556
rect 3612 4496 3616 4556
rect 3620 4496 3624 4556
rect 3628 4496 3632 4556
rect 3714 4516 3718 4556
rect 3722 4516 3726 4556
rect 3744 4536 3748 4556
rect 3811 4516 3815 4556
rect 3831 4516 3835 4556
rect 3851 4516 3855 4556
rect 3925 4516 3929 4556
rect 3945 4516 3949 4556
rect 3965 4516 3969 4556
rect 4048 4496 4052 4556
rect 4056 4496 4060 4556
rect 4064 4496 4068 4556
rect 4148 4496 4152 4556
rect 4156 4496 4160 4556
rect 4164 4496 4168 4556
rect 4214 4516 4218 4556
rect 4222 4516 4226 4556
rect 4244 4536 4248 4556
rect 4313 4516 4317 4556
rect 4323 4516 4327 4556
rect 4412 4536 4416 4556
rect 4434 4516 4438 4556
rect 4442 4516 4446 4556
rect 4505 4536 4509 4556
rect 4552 4496 4556 4556
rect 4560 4496 4564 4556
rect 4568 4496 4572 4556
rect 4652 4496 4656 4556
rect 4660 4496 4664 4556
rect 4668 4496 4672 4556
rect 45 4104 49 4144
rect 65 4104 69 4144
rect 85 4104 89 4144
rect 155 4104 159 4144
rect 175 4104 179 4144
rect 185 4104 189 4144
rect 231 4104 235 4124
rect 251 4104 255 4124
rect 332 4104 336 4124
rect 354 4104 358 4144
rect 362 4104 366 4144
rect 411 4104 415 4144
rect 421 4104 425 4144
rect 441 4104 445 4144
rect 532 4104 536 4124
rect 554 4104 558 4144
rect 562 4104 566 4144
rect 612 4104 616 4164
rect 620 4104 624 4164
rect 628 4104 632 4164
rect 714 4104 718 4144
rect 722 4104 726 4144
rect 744 4104 748 4124
rect 811 4104 815 4144
rect 821 4104 825 4144
rect 841 4104 845 4144
rect 925 4104 929 4144
rect 945 4104 949 4144
rect 965 4104 969 4144
rect 1025 4104 1029 4124
rect 1071 4104 1075 4124
rect 1091 4104 1095 4124
rect 1151 4104 1155 4124
rect 1171 4104 1175 4124
rect 1231 4104 1235 4124
rect 1251 4104 1255 4124
rect 1311 4104 1315 4124
rect 1371 4104 1375 4144
rect 1393 4104 1397 4124
rect 1403 4104 1407 4124
rect 1423 4104 1427 4124
rect 1431 4104 1435 4124
rect 1477 4104 1481 4124
rect 1499 4104 1503 4124
rect 1509 4104 1513 4124
rect 1531 4104 1535 4124
rect 1541 4104 1545 4124
rect 1561 4104 1565 4144
rect 1611 4104 1615 4144
rect 1631 4104 1635 4144
rect 1651 4104 1655 4144
rect 1711 4104 1715 4124
rect 1731 4104 1735 4124
rect 1805 4104 1809 4124
rect 1851 4104 1855 4144
rect 1873 4104 1877 4124
rect 1883 4104 1887 4124
rect 1903 4104 1907 4124
rect 1911 4104 1915 4124
rect 1957 4104 1961 4124
rect 1979 4104 1983 4124
rect 1989 4104 1993 4124
rect 2011 4104 2015 4124
rect 2021 4104 2025 4124
rect 2041 4104 2045 4144
rect 2113 4104 2117 4144
rect 2123 4104 2127 4144
rect 2171 4104 2175 4124
rect 2191 4104 2195 4124
rect 2211 4104 2215 4144
rect 2306 4104 2310 4144
rect 2314 4104 2318 4144
rect 2334 4104 2338 4144
rect 2342 4104 2346 4144
rect 2393 4104 2397 4144
rect 2403 4104 2407 4144
rect 2485 4104 2489 4144
rect 2505 4104 2509 4144
rect 2525 4104 2529 4144
rect 2585 4104 2589 4124
rect 2605 4104 2609 4124
rect 2654 4104 2658 4144
rect 2662 4104 2666 4144
rect 2684 4104 2688 4124
rect 2772 4104 2776 4124
rect 2794 4104 2798 4144
rect 2802 4104 2806 4144
rect 2851 4104 2855 4124
rect 2873 4104 2877 4144
rect 2968 4104 2972 4164
rect 2976 4104 2980 4164
rect 2984 4104 2988 4164
rect 3068 4104 3072 4164
rect 3076 4104 3080 4164
rect 3084 4104 3088 4164
rect 3133 4104 3137 4144
rect 3143 4104 3147 4144
rect 3225 4104 3229 4124
rect 3308 4104 3312 4164
rect 3316 4104 3320 4164
rect 3324 4104 3328 4164
rect 3408 4104 3412 4164
rect 3416 4104 3420 4164
rect 3424 4104 3428 4164
rect 3508 4104 3512 4164
rect 3516 4104 3520 4164
rect 3524 4104 3528 4164
rect 3608 4104 3612 4164
rect 3616 4104 3620 4164
rect 3624 4104 3628 4164
rect 3672 4104 3676 4164
rect 3680 4104 3684 4164
rect 3688 4104 3692 4164
rect 3774 4104 3778 4144
rect 3782 4104 3786 4144
rect 3804 4104 3808 4124
rect 3871 4104 3875 4144
rect 3891 4104 3895 4144
rect 3911 4104 3915 4144
rect 3971 4104 3975 4124
rect 4034 4104 4038 4144
rect 4042 4104 4046 4144
rect 4064 4104 4068 4124
rect 4168 4104 4172 4164
rect 4176 4104 4180 4164
rect 4184 4104 4188 4164
rect 4232 4104 4236 4164
rect 4240 4104 4244 4164
rect 4248 4104 4252 4164
rect 4334 4104 4338 4144
rect 4342 4104 4346 4144
rect 4364 4104 4368 4124
rect 4431 4104 4435 4144
rect 4451 4104 4455 4144
rect 4471 4104 4475 4144
rect 4534 4104 4538 4144
rect 4542 4104 4546 4144
rect 4562 4104 4566 4144
rect 4570 4104 4574 4144
rect 4665 4104 4669 4124
rect 4685 4104 4689 4124
rect 53 4036 57 4076
rect 63 4036 67 4076
rect 133 4036 137 4076
rect 143 4036 147 4076
rect 205 4056 209 4076
rect 225 4056 229 4076
rect 271 4036 275 4076
rect 291 4036 295 4076
rect 311 4036 315 4076
rect 385 4056 389 4076
rect 445 4056 449 4076
rect 505 4056 509 4076
rect 525 4056 529 4076
rect 571 4036 575 4076
rect 581 4036 585 4076
rect 601 4036 605 4076
rect 671 4036 675 4076
rect 691 4036 695 4076
rect 711 4036 715 4076
rect 771 4056 775 4076
rect 831 4036 835 4076
rect 851 4036 855 4076
rect 871 4036 875 4076
rect 933 4036 937 4076
rect 943 4036 947 4076
rect 1025 4056 1029 4076
rect 1085 4056 1089 4076
rect 1105 4056 1109 4076
rect 1151 4056 1155 4076
rect 1211 4056 1215 4076
rect 1231 4056 1235 4076
rect 1291 4056 1295 4076
rect 1365 4056 1369 4076
rect 1385 4056 1389 4076
rect 1445 4056 1449 4076
rect 1491 4036 1495 4076
rect 1511 4036 1515 4076
rect 1531 4036 1535 4076
rect 1591 4036 1595 4076
rect 1611 4036 1615 4076
rect 1631 4036 1635 4076
rect 1651 4036 1655 4076
rect 1713 4036 1717 4076
rect 1723 4036 1727 4076
rect 1812 4056 1816 4076
rect 1834 4036 1838 4076
rect 1842 4036 1846 4076
rect 1892 4016 1896 4076
rect 1900 4016 1904 4076
rect 1908 4016 1912 4076
rect 2005 4036 2009 4076
rect 2025 4036 2029 4076
rect 2045 4036 2049 4076
rect 2105 4056 2109 4076
rect 2188 4016 2192 4076
rect 2196 4016 2200 4076
rect 2204 4016 2208 4076
rect 2288 4016 2292 4076
rect 2296 4016 2300 4076
rect 2304 4016 2308 4076
rect 2372 4056 2376 4076
rect 2394 4036 2398 4076
rect 2402 4036 2406 4076
rect 2465 4056 2469 4076
rect 2525 4036 2529 4076
rect 2545 4036 2549 4076
rect 2565 4036 2569 4076
rect 2648 4016 2652 4076
rect 2656 4016 2660 4076
rect 2664 4016 2668 4076
rect 2732 4056 2736 4076
rect 2754 4036 2758 4076
rect 2762 4036 2766 4076
rect 2825 4036 2829 4076
rect 2845 4036 2849 4076
rect 2865 4036 2869 4076
rect 2911 4036 2915 4076
rect 2931 4036 2935 4076
rect 2951 4036 2955 4076
rect 3048 4016 3052 4076
rect 3056 4016 3060 4076
rect 3064 4016 3068 4076
rect 3125 4056 3129 4076
rect 3171 4036 3175 4076
rect 3191 4036 3195 4076
rect 3211 4036 3215 4076
rect 3274 4036 3278 4076
rect 3282 4036 3286 4076
rect 3304 4056 3308 4076
rect 3371 4036 3375 4076
rect 3391 4036 3395 4076
rect 3411 4036 3415 4076
rect 3485 4036 3489 4076
rect 3505 4036 3509 4076
rect 3525 4036 3529 4076
rect 3585 4036 3589 4076
rect 3605 4036 3609 4076
rect 3625 4036 3629 4076
rect 3692 4056 3696 4076
rect 3714 4036 3718 4076
rect 3722 4036 3726 4076
rect 3808 4016 3812 4076
rect 3816 4016 3820 4076
rect 3824 4016 3828 4076
rect 3893 4036 3897 4076
rect 3903 4036 3907 4076
rect 3973 4036 3977 4076
rect 3983 4036 3987 4076
rect 4033 4036 4037 4076
rect 4043 4036 4047 4076
rect 4148 4016 4152 4076
rect 4156 4016 4160 4076
rect 4164 4016 4168 4076
rect 4225 4036 4229 4076
rect 4245 4036 4249 4076
rect 4265 4036 4269 4076
rect 4311 4036 4315 4076
rect 4331 4036 4335 4076
rect 4351 4036 4355 4076
rect 4425 4056 4429 4076
rect 4508 4016 4512 4076
rect 4516 4016 4520 4076
rect 4524 4016 4528 4076
rect 4608 4016 4612 4076
rect 4616 4016 4620 4076
rect 4624 4016 4628 4076
rect 4674 4036 4678 4076
rect 4682 4036 4686 4076
rect 4704 4056 4708 4076
rect 45 3624 49 3664
rect 65 3624 69 3664
rect 85 3624 89 3664
rect 145 3624 149 3644
rect 191 3624 195 3664
rect 213 3624 217 3644
rect 223 3624 227 3644
rect 243 3624 247 3644
rect 251 3624 255 3644
rect 297 3624 301 3644
rect 319 3624 323 3644
rect 329 3624 333 3644
rect 351 3624 355 3644
rect 361 3624 365 3644
rect 381 3624 385 3664
rect 445 3624 449 3664
rect 465 3624 469 3664
rect 485 3624 489 3664
rect 531 3624 535 3664
rect 541 3624 545 3664
rect 561 3624 565 3664
rect 645 3624 649 3664
rect 665 3624 669 3644
rect 685 3624 689 3644
rect 753 3624 757 3664
rect 763 3624 767 3664
rect 815 3624 819 3664
rect 835 3624 839 3644
rect 845 3624 849 3644
rect 867 3624 871 3644
rect 877 3624 881 3644
rect 899 3624 903 3644
rect 945 3624 949 3644
rect 953 3624 957 3644
rect 973 3624 977 3644
rect 983 3624 987 3644
rect 1005 3624 1009 3664
rect 1063 3624 1067 3664
rect 1085 3624 1089 3644
rect 1131 3624 1135 3664
rect 1153 3624 1157 3644
rect 1163 3624 1167 3644
rect 1183 3624 1187 3644
rect 1191 3624 1195 3644
rect 1237 3624 1241 3644
rect 1259 3624 1263 3644
rect 1269 3624 1273 3644
rect 1291 3624 1295 3644
rect 1301 3624 1305 3644
rect 1321 3624 1325 3664
rect 1371 3624 1375 3664
rect 1391 3624 1395 3664
rect 1411 3624 1415 3664
rect 1473 3624 1477 3664
rect 1483 3624 1487 3664
rect 1553 3624 1557 3664
rect 1563 3624 1567 3664
rect 1631 3624 1635 3644
rect 1653 3624 1657 3664
rect 1711 3624 1715 3664
rect 1733 3624 1737 3644
rect 1743 3624 1747 3644
rect 1763 3624 1767 3644
rect 1771 3624 1775 3644
rect 1817 3624 1821 3644
rect 1839 3624 1843 3644
rect 1849 3624 1853 3644
rect 1871 3624 1875 3644
rect 1881 3624 1885 3644
rect 1901 3624 1905 3664
rect 1965 3624 1969 3644
rect 2032 3624 2036 3644
rect 2054 3624 2058 3664
rect 2062 3624 2066 3664
rect 2125 3624 2129 3644
rect 2172 3624 2176 3684
rect 2180 3624 2184 3684
rect 2188 3624 2192 3684
rect 2285 3624 2289 3664
rect 2305 3624 2309 3664
rect 2325 3624 2329 3664
rect 2408 3624 2412 3684
rect 2416 3624 2420 3684
rect 2424 3624 2428 3684
rect 2492 3624 2496 3644
rect 2514 3624 2518 3664
rect 2522 3624 2526 3664
rect 2608 3624 2612 3684
rect 2616 3624 2620 3684
rect 2624 3624 2628 3684
rect 2674 3624 2678 3664
rect 2682 3624 2686 3664
rect 2704 3624 2708 3644
rect 2792 3624 2796 3644
rect 2814 3624 2818 3664
rect 2822 3624 2826 3664
rect 2885 3624 2889 3644
rect 2945 3624 2949 3644
rect 3028 3624 3032 3684
rect 3036 3624 3040 3684
rect 3044 3624 3048 3684
rect 3112 3624 3116 3644
rect 3134 3624 3138 3664
rect 3142 3624 3146 3664
rect 3228 3624 3232 3684
rect 3236 3624 3240 3684
rect 3244 3624 3248 3684
rect 3305 3624 3309 3644
rect 3365 3624 3369 3664
rect 3385 3624 3389 3664
rect 3405 3624 3409 3664
rect 3473 3624 3477 3664
rect 3483 3624 3487 3664
rect 3531 3624 3535 3664
rect 3541 3624 3545 3664
rect 3561 3624 3565 3664
rect 3652 3624 3656 3644
rect 3674 3624 3678 3664
rect 3682 3624 3686 3664
rect 3768 3624 3772 3684
rect 3776 3624 3780 3684
rect 3784 3624 3788 3684
rect 3845 3624 3849 3644
rect 3894 3624 3898 3664
rect 3902 3624 3906 3664
rect 3924 3624 3928 3644
rect 4005 3624 4009 3664
rect 4025 3624 4029 3664
rect 4045 3624 4049 3664
rect 4091 3624 4095 3664
rect 4111 3624 4115 3664
rect 4131 3624 4135 3664
rect 4194 3624 4198 3664
rect 4202 3624 4206 3664
rect 4224 3624 4228 3644
rect 4312 3624 4316 3644
rect 4334 3624 4338 3664
rect 4342 3624 4346 3664
rect 4392 3624 4396 3684
rect 4400 3624 4404 3684
rect 4408 3624 4412 3684
rect 4505 3624 4509 3644
rect 4588 3624 4592 3684
rect 4596 3624 4600 3684
rect 4604 3624 4608 3684
rect 4652 3624 4656 3684
rect 4660 3624 4664 3684
rect 4668 3624 4672 3684
rect 35 3556 39 3596
rect 55 3576 59 3596
rect 65 3576 69 3596
rect 87 3576 91 3596
rect 97 3576 101 3596
rect 119 3576 123 3596
rect 165 3576 169 3596
rect 173 3576 177 3596
rect 193 3576 197 3596
rect 203 3576 207 3596
rect 225 3556 229 3596
rect 293 3556 297 3596
rect 303 3556 307 3596
rect 365 3556 369 3596
rect 385 3556 389 3596
rect 405 3556 409 3596
rect 473 3556 477 3596
rect 483 3556 487 3596
rect 568 3536 572 3596
rect 576 3536 580 3596
rect 584 3536 588 3596
rect 645 3576 649 3596
rect 705 3556 709 3596
rect 725 3556 729 3596
rect 745 3556 749 3596
rect 805 3556 809 3596
rect 825 3556 829 3596
rect 845 3556 849 3596
rect 891 3576 895 3596
rect 965 3576 969 3596
rect 985 3576 989 3596
rect 1031 3556 1035 3596
rect 1053 3576 1057 3596
rect 1063 3576 1067 3596
rect 1083 3576 1087 3596
rect 1091 3576 1095 3596
rect 1137 3576 1141 3596
rect 1159 3576 1163 3596
rect 1169 3576 1173 3596
rect 1191 3576 1195 3596
rect 1201 3576 1205 3596
rect 1221 3556 1225 3596
rect 1271 3576 1275 3596
rect 1331 3576 1335 3596
rect 1351 3576 1355 3596
rect 1411 3556 1415 3596
rect 1431 3556 1435 3596
rect 1451 3556 1455 3596
rect 1513 3556 1517 3596
rect 1523 3556 1527 3596
rect 1603 3556 1607 3596
rect 1625 3576 1629 3596
rect 1685 3576 1689 3596
rect 1731 3556 1735 3596
rect 1753 3576 1757 3596
rect 1763 3576 1767 3596
rect 1783 3576 1787 3596
rect 1791 3576 1795 3596
rect 1837 3576 1841 3596
rect 1859 3576 1863 3596
rect 1869 3576 1873 3596
rect 1891 3576 1895 3596
rect 1901 3576 1905 3596
rect 1921 3556 1925 3596
rect 1971 3556 1975 3596
rect 1991 3556 1995 3596
rect 2011 3556 2015 3596
rect 2031 3556 2035 3596
rect 2093 3556 2097 3596
rect 2103 3556 2107 3596
rect 2192 3576 2196 3596
rect 2214 3556 2218 3596
rect 2222 3556 2226 3596
rect 2308 3536 2312 3596
rect 2316 3536 2320 3596
rect 2324 3536 2328 3596
rect 2385 3576 2389 3596
rect 2468 3536 2472 3596
rect 2476 3536 2480 3596
rect 2484 3536 2488 3596
rect 2568 3536 2572 3596
rect 2576 3536 2580 3596
rect 2584 3536 2588 3596
rect 2645 3556 2649 3596
rect 2665 3556 2669 3596
rect 2685 3556 2689 3596
rect 2731 3556 2735 3596
rect 2751 3556 2755 3596
rect 2771 3556 2775 3596
rect 2833 3556 2837 3596
rect 2843 3556 2847 3596
rect 2911 3556 2915 3596
rect 2931 3556 2935 3596
rect 2951 3556 2955 3596
rect 3011 3576 3015 3596
rect 3031 3576 3035 3596
rect 3105 3556 3109 3596
rect 3125 3556 3129 3596
rect 3145 3556 3149 3596
rect 3194 3556 3198 3596
rect 3202 3556 3206 3596
rect 3222 3556 3226 3596
rect 3230 3556 3234 3596
rect 3313 3556 3317 3596
rect 3323 3556 3327 3596
rect 3393 3556 3397 3596
rect 3403 3556 3407 3596
rect 3473 3556 3477 3596
rect 3483 3556 3487 3596
rect 3551 3576 3555 3596
rect 3571 3576 3575 3596
rect 3633 3556 3637 3596
rect 3643 3556 3647 3596
rect 3713 3556 3717 3596
rect 3723 3556 3727 3596
rect 3813 3556 3817 3596
rect 3823 3556 3827 3596
rect 3885 3576 3889 3596
rect 3905 3576 3909 3596
rect 3953 3556 3957 3596
rect 3963 3556 3967 3596
rect 4033 3556 4037 3596
rect 4043 3556 4047 3596
rect 4111 3556 4115 3596
rect 4131 3556 4135 3596
rect 4151 3556 4155 3596
rect 4248 3536 4252 3596
rect 4256 3536 4260 3596
rect 4264 3536 4268 3596
rect 4312 3536 4316 3596
rect 4320 3536 4324 3596
rect 4328 3536 4332 3596
rect 4414 3556 4418 3596
rect 4422 3556 4426 3596
rect 4444 3576 4448 3596
rect 4511 3576 4515 3596
rect 4608 3536 4612 3596
rect 4616 3536 4620 3596
rect 4624 3536 4628 3596
rect 4672 3536 4676 3596
rect 4680 3536 4684 3596
rect 4688 3536 4692 3596
rect 35 3144 39 3184
rect 55 3144 59 3164
rect 65 3144 69 3164
rect 87 3144 91 3164
rect 97 3144 101 3164
rect 119 3144 123 3164
rect 165 3144 169 3164
rect 173 3144 177 3164
rect 193 3144 197 3164
rect 203 3144 207 3164
rect 225 3144 229 3184
rect 306 3144 310 3184
rect 314 3144 318 3184
rect 334 3144 338 3184
rect 342 3144 346 3184
rect 393 3144 397 3184
rect 403 3144 407 3184
rect 471 3144 475 3184
rect 491 3144 495 3184
rect 511 3144 515 3184
rect 571 3144 575 3184
rect 591 3144 595 3184
rect 611 3144 615 3184
rect 693 3144 697 3184
rect 703 3144 707 3184
rect 751 3144 755 3164
rect 825 3144 829 3184
rect 845 3144 849 3184
rect 865 3144 869 3184
rect 885 3144 889 3184
rect 905 3144 909 3184
rect 925 3144 929 3184
rect 945 3144 949 3184
rect 965 3144 969 3184
rect 1011 3144 1015 3184
rect 1031 3144 1035 3184
rect 1051 3144 1055 3184
rect 1071 3144 1075 3184
rect 1091 3144 1095 3184
rect 1111 3144 1115 3184
rect 1131 3144 1135 3184
rect 1151 3144 1155 3184
rect 1225 3144 1229 3164
rect 1271 3144 1275 3184
rect 1293 3144 1297 3164
rect 1303 3144 1307 3164
rect 1323 3144 1327 3164
rect 1331 3144 1335 3164
rect 1377 3144 1381 3164
rect 1399 3144 1403 3164
rect 1409 3144 1413 3164
rect 1431 3144 1435 3164
rect 1441 3144 1445 3164
rect 1461 3144 1465 3184
rect 1511 3144 1515 3184
rect 1531 3144 1535 3184
rect 1551 3144 1555 3184
rect 1625 3144 1629 3184
rect 1645 3144 1649 3184
rect 1665 3144 1669 3184
rect 1725 3144 1729 3184
rect 1745 3144 1749 3184
rect 1765 3144 1769 3184
rect 1825 3144 1829 3164
rect 1885 3144 1889 3184
rect 1905 3144 1909 3184
rect 1925 3144 1929 3184
rect 1985 3144 1989 3184
rect 2005 3144 2009 3184
rect 2025 3144 2029 3184
rect 2071 3144 2075 3184
rect 2093 3144 2097 3164
rect 2103 3144 2107 3164
rect 2123 3144 2127 3164
rect 2131 3144 2135 3164
rect 2177 3144 2181 3164
rect 2199 3144 2203 3164
rect 2209 3144 2213 3164
rect 2231 3144 2235 3164
rect 2241 3144 2245 3164
rect 2261 3144 2265 3184
rect 2325 3144 2329 3164
rect 2385 3144 2389 3164
rect 2468 3144 2472 3204
rect 2476 3144 2480 3204
rect 2484 3144 2488 3204
rect 2534 3144 2538 3184
rect 2542 3144 2546 3184
rect 2564 3144 2568 3164
rect 2645 3144 2649 3164
rect 2705 3144 2709 3184
rect 2725 3144 2729 3184
rect 2745 3144 2749 3184
rect 2791 3144 2795 3164
rect 2811 3144 2815 3164
rect 2871 3144 2875 3184
rect 2891 3144 2895 3184
rect 2911 3144 2915 3184
rect 2973 3144 2977 3184
rect 2983 3144 2987 3184
rect 3053 3144 3057 3184
rect 3063 3144 3067 3184
rect 3152 3144 3156 3164
rect 3174 3144 3178 3184
rect 3182 3144 3186 3184
rect 3268 3144 3272 3204
rect 3276 3144 3280 3204
rect 3284 3144 3288 3204
rect 3345 3144 3349 3184
rect 3365 3144 3369 3184
rect 3385 3144 3389 3184
rect 3455 3144 3459 3184
rect 3475 3144 3479 3184
rect 3485 3144 3489 3184
rect 3533 3144 3537 3184
rect 3543 3144 3547 3184
rect 3635 3144 3639 3184
rect 3655 3144 3659 3184
rect 3665 3144 3669 3184
rect 3746 3144 3750 3184
rect 3754 3144 3758 3184
rect 3774 3144 3778 3184
rect 3782 3144 3786 3184
rect 3853 3144 3857 3184
rect 3863 3144 3867 3184
rect 3911 3144 3915 3184
rect 3931 3144 3935 3184
rect 3951 3144 3955 3184
rect 4013 3144 4017 3184
rect 4023 3144 4027 3184
rect 4115 3144 4119 3184
rect 4135 3144 4139 3184
rect 4145 3144 4149 3184
rect 4193 3144 4197 3184
rect 4203 3144 4207 3184
rect 4271 3144 4275 3184
rect 4281 3144 4285 3184
rect 4301 3144 4305 3184
rect 4374 3144 4378 3184
rect 4382 3144 4386 3184
rect 4404 3144 4408 3164
rect 4471 3144 4475 3184
rect 4491 3144 4495 3184
rect 4511 3144 4515 3184
rect 4571 3144 4575 3184
rect 4591 3144 4595 3184
rect 4611 3144 4615 3184
rect 4708 3144 4712 3204
rect 4716 3144 4720 3204
rect 4724 3144 4728 3204
rect 35 3076 39 3116
rect 55 3096 59 3116
rect 65 3096 69 3116
rect 87 3096 91 3116
rect 97 3096 101 3116
rect 119 3096 123 3116
rect 165 3096 169 3116
rect 173 3096 177 3116
rect 193 3096 197 3116
rect 203 3096 207 3116
rect 225 3076 229 3116
rect 285 3076 289 3116
rect 305 3076 309 3116
rect 325 3076 329 3116
rect 393 3076 397 3116
rect 403 3076 407 3116
rect 451 3076 455 3116
rect 473 3096 477 3116
rect 483 3096 487 3116
rect 503 3096 507 3116
rect 511 3096 515 3116
rect 557 3096 561 3116
rect 579 3096 583 3116
rect 589 3096 593 3116
rect 611 3096 615 3116
rect 621 3096 625 3116
rect 641 3076 645 3116
rect 695 3076 699 3116
rect 715 3096 719 3116
rect 725 3096 729 3116
rect 747 3096 751 3116
rect 757 3096 761 3116
rect 779 3096 783 3116
rect 825 3096 829 3116
rect 833 3096 837 3116
rect 853 3096 857 3116
rect 863 3096 867 3116
rect 885 3076 889 3116
rect 931 3096 935 3116
rect 1005 3096 1009 3116
rect 1025 3096 1029 3116
rect 1093 3076 1097 3116
rect 1103 3076 1107 3116
rect 1151 3076 1155 3116
rect 1171 3076 1175 3116
rect 1191 3076 1195 3116
rect 1254 3076 1258 3116
rect 1262 3076 1266 3116
rect 1284 3096 1288 3116
rect 1355 3076 1359 3116
rect 1375 3096 1379 3116
rect 1385 3096 1389 3116
rect 1407 3096 1411 3116
rect 1417 3096 1421 3116
rect 1439 3096 1443 3116
rect 1485 3096 1489 3116
rect 1493 3096 1497 3116
rect 1513 3096 1517 3116
rect 1523 3096 1527 3116
rect 1545 3076 1549 3116
rect 1605 3096 1609 3116
rect 1625 3096 1629 3116
rect 1693 3076 1697 3116
rect 1703 3076 1707 3116
rect 1751 3076 1755 3116
rect 1771 3076 1775 3116
rect 1791 3076 1795 3116
rect 1865 3076 1869 3116
rect 1885 3076 1889 3116
rect 1905 3076 1909 3116
rect 1951 3076 1955 3116
rect 1973 3096 1977 3116
rect 1983 3096 1987 3116
rect 2003 3096 2007 3116
rect 2011 3096 2015 3116
rect 2057 3096 2061 3116
rect 2079 3096 2083 3116
rect 2089 3096 2093 3116
rect 2111 3096 2115 3116
rect 2121 3096 2125 3116
rect 2141 3076 2145 3116
rect 2205 3096 2209 3116
rect 2225 3096 2229 3116
rect 2285 3096 2289 3116
rect 2368 3056 2372 3116
rect 2376 3056 2380 3116
rect 2384 3056 2388 3116
rect 2452 3096 2456 3116
rect 2474 3076 2478 3116
rect 2482 3076 2486 3116
rect 2568 3056 2572 3116
rect 2576 3056 2580 3116
rect 2584 3056 2588 3116
rect 2645 3076 2649 3116
rect 2665 3076 2669 3116
rect 2685 3076 2689 3116
rect 2745 3096 2749 3116
rect 2765 3096 2769 3116
rect 2813 3076 2817 3116
rect 2823 3076 2827 3116
rect 2893 3076 2897 3116
rect 2903 3076 2907 3116
rect 2974 3076 2978 3116
rect 2982 3076 2986 3116
rect 3002 3076 3006 3116
rect 3010 3076 3014 3116
rect 3093 3076 3097 3116
rect 3103 3076 3107 3116
rect 3171 3076 3175 3116
rect 3191 3076 3195 3116
rect 3211 3076 3215 3116
rect 3271 3076 3275 3116
rect 3331 3076 3335 3116
rect 3341 3076 3345 3116
rect 3361 3076 3365 3116
rect 3443 3076 3447 3116
rect 3465 3096 3469 3116
rect 3523 3076 3527 3116
rect 3545 3096 3549 3116
rect 3593 3076 3597 3116
rect 3603 3076 3607 3116
rect 3671 3076 3675 3116
rect 3691 3076 3695 3116
rect 3711 3076 3715 3116
rect 3783 3076 3787 3116
rect 3805 3096 3809 3116
rect 3851 3076 3855 3116
rect 3871 3076 3875 3116
rect 3891 3076 3895 3116
rect 3952 3056 3956 3116
rect 3960 3056 3964 3116
rect 3968 3056 3972 3116
rect 4051 3096 4055 3116
rect 4073 3076 4077 3116
rect 4152 3096 4156 3116
rect 4174 3076 4178 3116
rect 4182 3076 4186 3116
rect 4232 3056 4236 3116
rect 4240 3056 4244 3116
rect 4248 3056 4252 3116
rect 4352 3096 4356 3116
rect 4374 3076 4378 3116
rect 4382 3076 4386 3116
rect 4468 3056 4472 3116
rect 4476 3056 4480 3116
rect 4484 3056 4488 3116
rect 4545 3096 4549 3116
rect 4605 3076 4609 3116
rect 4625 3076 4629 3116
rect 4645 3076 4649 3116
rect 4691 3076 4695 3116
rect 4711 3076 4715 3116
rect 4731 3076 4735 3116
rect 35 2664 39 2704
rect 55 2664 59 2684
rect 65 2664 69 2684
rect 87 2664 91 2684
rect 97 2664 101 2684
rect 119 2664 123 2684
rect 165 2664 169 2684
rect 173 2664 177 2684
rect 193 2664 197 2684
rect 203 2664 207 2684
rect 225 2664 229 2704
rect 306 2664 310 2704
rect 314 2664 318 2704
rect 334 2664 338 2704
rect 342 2664 346 2704
rect 393 2664 397 2704
rect 403 2664 407 2704
rect 485 2664 489 2704
rect 505 2664 509 2704
rect 525 2664 529 2704
rect 583 2664 587 2704
rect 605 2664 609 2684
rect 653 2664 657 2704
rect 663 2664 667 2704
rect 745 2664 749 2704
rect 765 2664 769 2704
rect 785 2664 789 2704
rect 845 2664 849 2684
rect 865 2664 869 2684
rect 933 2664 937 2704
rect 943 2664 947 2704
rect 991 2664 995 2684
rect 1073 2664 1077 2704
rect 1083 2664 1087 2704
rect 1131 2664 1135 2684
rect 1151 2664 1155 2684
rect 1223 2664 1227 2704
rect 1245 2664 1249 2684
rect 1295 2664 1299 2704
rect 1315 2664 1319 2684
rect 1325 2664 1329 2684
rect 1347 2664 1351 2684
rect 1357 2664 1361 2684
rect 1379 2664 1383 2684
rect 1425 2664 1429 2684
rect 1433 2664 1437 2684
rect 1453 2664 1457 2684
rect 1463 2664 1467 2684
rect 1485 2664 1489 2704
rect 1533 2664 1537 2704
rect 1543 2664 1547 2704
rect 1625 2664 1629 2704
rect 1645 2664 1649 2704
rect 1665 2664 1669 2704
rect 1725 2664 1729 2704
rect 1745 2664 1749 2704
rect 1765 2664 1769 2704
rect 1825 2664 1829 2684
rect 1845 2664 1849 2684
rect 1912 2664 1916 2684
rect 1934 2664 1938 2704
rect 1942 2664 1946 2704
rect 2003 2664 2007 2704
rect 2025 2664 2029 2684
rect 2108 2664 2112 2724
rect 2116 2664 2120 2724
rect 2124 2664 2128 2724
rect 2171 2664 2175 2684
rect 2193 2664 2197 2704
rect 2255 2664 2259 2704
rect 2275 2664 2279 2684
rect 2285 2664 2289 2684
rect 2307 2664 2311 2684
rect 2317 2664 2321 2684
rect 2339 2664 2343 2684
rect 2385 2664 2389 2684
rect 2393 2664 2397 2684
rect 2413 2664 2417 2684
rect 2423 2664 2427 2684
rect 2445 2664 2449 2704
rect 2505 2664 2509 2704
rect 2525 2664 2529 2704
rect 2545 2664 2549 2704
rect 2605 2664 2609 2704
rect 2625 2664 2629 2704
rect 2645 2664 2649 2704
rect 2691 2664 2695 2704
rect 2711 2664 2715 2704
rect 2731 2664 2735 2704
rect 2793 2664 2797 2704
rect 2803 2664 2807 2704
rect 2873 2664 2877 2704
rect 2883 2664 2887 2704
rect 2951 2664 2955 2704
rect 2971 2664 2975 2704
rect 2991 2664 2995 2704
rect 3051 2664 3055 2704
rect 3071 2664 3075 2704
rect 3091 2664 3095 2704
rect 3153 2664 3157 2704
rect 3163 2664 3167 2704
rect 3245 2664 3249 2704
rect 3265 2664 3269 2704
rect 3285 2664 3289 2704
rect 3353 2664 3357 2704
rect 3363 2664 3367 2704
rect 3412 2664 3416 2724
rect 3420 2664 3424 2724
rect 3428 2664 3432 2724
rect 3525 2664 3529 2704
rect 3545 2664 3549 2704
rect 3565 2664 3569 2704
rect 3611 2664 3615 2704
rect 3631 2664 3635 2704
rect 3651 2664 3655 2704
rect 3733 2664 3737 2704
rect 3743 2664 3747 2704
rect 3805 2664 3809 2704
rect 3825 2664 3829 2704
rect 3845 2664 3849 2704
rect 3892 2664 3896 2724
rect 3900 2664 3904 2724
rect 3908 2664 3912 2724
rect 3991 2664 3995 2684
rect 4086 2664 4090 2704
rect 4094 2664 4098 2704
rect 4114 2664 4118 2704
rect 4122 2664 4126 2704
rect 4172 2664 4176 2724
rect 4180 2664 4184 2724
rect 4188 2664 4192 2724
rect 4271 2664 4275 2704
rect 4291 2664 4295 2704
rect 4311 2664 4315 2704
rect 4371 2664 4375 2704
rect 4381 2664 4385 2704
rect 4401 2664 4405 2704
rect 4474 2664 4478 2704
rect 4482 2664 4486 2704
rect 4502 2664 4506 2704
rect 4510 2664 4514 2704
rect 4591 2664 4595 2684
rect 4654 2664 4658 2704
rect 4662 2664 4666 2704
rect 4684 2664 4688 2684
rect 35 2596 39 2636
rect 55 2616 59 2636
rect 65 2616 69 2636
rect 87 2616 91 2636
rect 97 2616 101 2636
rect 119 2616 123 2636
rect 165 2616 169 2636
rect 173 2616 177 2636
rect 193 2616 197 2636
rect 203 2616 207 2636
rect 225 2596 229 2636
rect 285 2596 289 2636
rect 305 2596 309 2636
rect 325 2596 329 2636
rect 371 2616 375 2636
rect 393 2596 397 2636
rect 453 2596 457 2636
rect 463 2596 467 2636
rect 545 2596 549 2636
rect 565 2596 569 2636
rect 585 2596 589 2636
rect 631 2616 635 2636
rect 653 2596 657 2636
rect 725 2596 729 2636
rect 745 2596 749 2636
rect 765 2596 769 2636
rect 811 2616 815 2636
rect 831 2616 835 2636
rect 895 2596 899 2636
rect 915 2616 919 2636
rect 925 2616 929 2636
rect 947 2616 951 2636
rect 957 2616 961 2636
rect 979 2616 983 2636
rect 1025 2616 1029 2636
rect 1033 2616 1037 2636
rect 1053 2616 1057 2636
rect 1063 2616 1067 2636
rect 1085 2596 1089 2636
rect 1131 2616 1135 2636
rect 1191 2596 1195 2636
rect 1211 2596 1215 2636
rect 1231 2596 1235 2636
rect 1291 2616 1295 2636
rect 1353 2596 1357 2636
rect 1363 2596 1367 2636
rect 1431 2596 1435 2636
rect 1453 2616 1457 2636
rect 1463 2616 1467 2636
rect 1483 2616 1487 2636
rect 1491 2616 1495 2636
rect 1537 2616 1541 2636
rect 1559 2616 1563 2636
rect 1569 2616 1573 2636
rect 1591 2616 1595 2636
rect 1601 2616 1605 2636
rect 1621 2596 1625 2636
rect 1671 2596 1675 2636
rect 1691 2596 1695 2636
rect 1711 2596 1715 2636
rect 1771 2596 1775 2636
rect 1793 2616 1797 2636
rect 1803 2616 1807 2636
rect 1823 2616 1827 2636
rect 1831 2616 1835 2636
rect 1877 2616 1881 2636
rect 1899 2616 1903 2636
rect 1909 2616 1913 2636
rect 1931 2616 1935 2636
rect 1941 2616 1945 2636
rect 1961 2596 1965 2636
rect 2011 2596 2015 2636
rect 2031 2596 2035 2636
rect 2051 2596 2055 2636
rect 2071 2596 2075 2636
rect 2091 2596 2095 2636
rect 2111 2596 2115 2636
rect 2131 2596 2135 2636
rect 2151 2596 2155 2636
rect 2215 2596 2219 2636
rect 2235 2616 2239 2636
rect 2245 2616 2249 2636
rect 2267 2616 2271 2636
rect 2277 2616 2281 2636
rect 2299 2616 2303 2636
rect 2345 2616 2349 2636
rect 2353 2616 2357 2636
rect 2373 2616 2377 2636
rect 2383 2616 2387 2636
rect 2405 2596 2409 2636
rect 2473 2596 2477 2636
rect 2483 2596 2487 2636
rect 2531 2616 2535 2636
rect 2605 2596 2609 2636
rect 2625 2596 2629 2636
rect 2645 2596 2649 2636
rect 2691 2616 2695 2636
rect 2773 2596 2777 2636
rect 2783 2596 2787 2636
rect 2845 2596 2849 2636
rect 2865 2596 2869 2636
rect 2885 2596 2889 2636
rect 2931 2596 2935 2636
rect 2941 2596 2945 2636
rect 2961 2596 2965 2636
rect 3031 2596 3035 2636
rect 3051 2596 3055 2636
rect 3071 2596 3075 2636
rect 3153 2596 3157 2636
rect 3163 2596 3167 2636
rect 3211 2596 3215 2636
rect 3221 2596 3225 2636
rect 3241 2596 3245 2636
rect 3348 2576 3352 2636
rect 3356 2576 3360 2636
rect 3364 2576 3368 2636
rect 3411 2616 3415 2636
rect 3473 2596 3477 2636
rect 3483 2596 3487 2636
rect 3551 2596 3555 2636
rect 3561 2596 3565 2636
rect 3581 2596 3585 2636
rect 3651 2616 3655 2636
rect 3673 2596 3677 2636
rect 3731 2616 3735 2636
rect 3815 2596 3819 2636
rect 3835 2596 3839 2636
rect 3845 2596 3849 2636
rect 3926 2596 3930 2636
rect 3934 2596 3938 2636
rect 3954 2596 3958 2636
rect 3962 2596 3966 2636
rect 4033 2596 4037 2636
rect 4043 2596 4047 2636
rect 4113 2596 4117 2636
rect 4123 2596 4127 2636
rect 4171 2596 4175 2636
rect 4191 2596 4195 2636
rect 4211 2596 4215 2636
rect 4273 2596 4277 2636
rect 4283 2596 4287 2636
rect 4388 2576 4392 2636
rect 4396 2576 4400 2636
rect 4404 2576 4408 2636
rect 4488 2576 4492 2636
rect 4496 2576 4500 2636
rect 4504 2576 4508 2636
rect 4554 2596 4558 2636
rect 4562 2596 4566 2636
rect 4584 2616 4588 2636
rect 4688 2576 4692 2636
rect 4696 2576 4700 2636
rect 4704 2576 4708 2636
rect 35 2184 39 2224
rect 55 2184 59 2204
rect 65 2184 69 2204
rect 87 2184 91 2204
rect 97 2184 101 2204
rect 119 2184 123 2204
rect 165 2184 169 2204
rect 173 2184 177 2204
rect 193 2184 197 2204
rect 203 2184 207 2204
rect 225 2184 229 2224
rect 271 2184 275 2224
rect 291 2184 295 2224
rect 311 2184 315 2224
rect 374 2184 378 2224
rect 382 2184 386 2224
rect 402 2184 406 2224
rect 410 2184 414 2224
rect 491 2184 495 2204
rect 513 2184 517 2224
rect 573 2184 577 2224
rect 583 2184 587 2224
rect 665 2184 669 2204
rect 711 2184 715 2204
rect 731 2184 735 2204
rect 812 2184 816 2204
rect 834 2184 838 2224
rect 842 2184 846 2224
rect 891 2184 895 2204
rect 911 2184 915 2204
rect 971 2184 975 2204
rect 991 2184 995 2204
rect 1051 2184 1055 2204
rect 1111 2184 1115 2224
rect 1133 2184 1137 2204
rect 1143 2184 1147 2204
rect 1163 2184 1167 2204
rect 1171 2184 1175 2204
rect 1217 2184 1221 2204
rect 1239 2184 1243 2204
rect 1249 2184 1253 2204
rect 1271 2184 1275 2204
rect 1281 2184 1285 2204
rect 1301 2184 1305 2224
rect 1351 2184 1355 2224
rect 1371 2184 1375 2224
rect 1391 2184 1395 2224
rect 1451 2184 1455 2224
rect 1473 2184 1477 2204
rect 1483 2184 1487 2204
rect 1503 2184 1507 2204
rect 1511 2184 1515 2204
rect 1557 2184 1561 2204
rect 1579 2184 1583 2204
rect 1589 2184 1593 2204
rect 1611 2184 1615 2204
rect 1621 2184 1625 2204
rect 1641 2184 1645 2224
rect 1705 2184 1709 2204
rect 1725 2184 1729 2204
rect 1792 2184 1796 2204
rect 1814 2184 1818 2224
rect 1822 2184 1826 2224
rect 1871 2184 1875 2224
rect 1945 2184 1949 2204
rect 1965 2184 1969 2204
rect 2011 2184 2015 2224
rect 2031 2184 2035 2224
rect 2051 2184 2055 2224
rect 2071 2184 2075 2224
rect 2091 2184 2095 2224
rect 2111 2184 2115 2224
rect 2131 2184 2135 2224
rect 2151 2184 2155 2224
rect 2211 2184 2215 2224
rect 2231 2184 2235 2224
rect 2251 2184 2255 2224
rect 2315 2184 2319 2224
rect 2335 2184 2339 2204
rect 2345 2184 2349 2204
rect 2367 2184 2371 2204
rect 2377 2184 2381 2204
rect 2399 2184 2403 2204
rect 2445 2184 2449 2204
rect 2453 2184 2457 2204
rect 2473 2184 2477 2204
rect 2483 2184 2487 2204
rect 2505 2184 2509 2224
rect 2573 2184 2577 2224
rect 2583 2184 2587 2224
rect 2633 2184 2637 2224
rect 2643 2184 2647 2224
rect 2713 2184 2717 2224
rect 2723 2184 2727 2224
rect 2805 2184 2809 2224
rect 2825 2184 2829 2224
rect 2845 2184 2849 2224
rect 2905 2184 2909 2224
rect 2925 2184 2929 2224
rect 2945 2184 2949 2224
rect 2995 2184 2999 2224
rect 3015 2184 3019 2204
rect 3025 2184 3029 2204
rect 3047 2184 3051 2204
rect 3057 2184 3061 2204
rect 3079 2184 3083 2204
rect 3125 2184 3129 2204
rect 3133 2184 3137 2204
rect 3153 2184 3157 2204
rect 3163 2184 3167 2204
rect 3185 2184 3189 2224
rect 3231 2184 3235 2224
rect 3251 2184 3255 2224
rect 3271 2184 3275 2224
rect 3333 2184 3337 2224
rect 3343 2184 3347 2224
rect 3413 2184 3417 2224
rect 3423 2184 3427 2224
rect 3513 2184 3517 2224
rect 3523 2184 3527 2224
rect 3585 2184 3589 2224
rect 3645 2184 3649 2224
rect 3705 2184 3709 2204
rect 3751 2184 3755 2224
rect 3771 2184 3775 2224
rect 3791 2184 3795 2224
rect 3863 2184 3867 2224
rect 3885 2184 3889 2204
rect 3931 2184 3935 2224
rect 3991 2184 3995 2224
rect 4001 2184 4005 2224
rect 4021 2184 4025 2224
rect 4105 2184 4109 2224
rect 4125 2184 4129 2224
rect 4145 2184 4149 2224
rect 4228 2184 4232 2244
rect 4236 2184 4240 2244
rect 4244 2184 4248 2244
rect 4294 2184 4298 2224
rect 4302 2184 4306 2224
rect 4324 2184 4328 2204
rect 4405 2184 4409 2224
rect 4425 2184 4429 2224
rect 4445 2184 4449 2224
rect 4491 2184 4495 2224
rect 4511 2184 4515 2224
rect 4531 2184 4535 2224
rect 4605 2184 4609 2224
rect 4625 2184 4629 2224
rect 4645 2184 4649 2224
rect 4694 2184 4698 2224
rect 4702 2184 4706 2224
rect 4724 2184 4728 2204
rect 31 2116 35 2156
rect 51 2116 55 2156
rect 71 2116 75 2156
rect 91 2116 95 2156
rect 111 2116 115 2156
rect 131 2116 135 2156
rect 151 2116 155 2156
rect 171 2116 175 2156
rect 253 2116 257 2156
rect 263 2116 267 2156
rect 325 2116 329 2156
rect 345 2116 349 2156
rect 365 2116 369 2156
rect 414 2116 418 2156
rect 422 2116 426 2156
rect 442 2116 446 2156
rect 450 2116 454 2156
rect 535 2116 539 2156
rect 555 2136 559 2156
rect 565 2136 569 2156
rect 587 2136 591 2156
rect 597 2136 601 2156
rect 619 2136 623 2156
rect 665 2136 669 2156
rect 673 2136 677 2156
rect 693 2136 697 2156
rect 703 2136 707 2156
rect 725 2116 729 2156
rect 793 2116 797 2156
rect 803 2116 807 2156
rect 865 2116 869 2156
rect 885 2136 889 2156
rect 905 2136 909 2156
rect 953 2116 957 2156
rect 963 2116 967 2156
rect 1031 2136 1035 2156
rect 1051 2136 1055 2156
rect 1111 2116 1115 2156
rect 1131 2116 1135 2156
rect 1151 2116 1155 2156
rect 1213 2116 1217 2156
rect 1223 2116 1227 2156
rect 1291 2136 1295 2156
rect 1311 2136 1315 2156
rect 1371 2116 1375 2156
rect 1393 2136 1397 2156
rect 1403 2136 1407 2156
rect 1423 2136 1427 2156
rect 1431 2136 1435 2156
rect 1477 2136 1481 2156
rect 1499 2136 1503 2156
rect 1509 2136 1513 2156
rect 1531 2136 1535 2156
rect 1541 2136 1545 2156
rect 1561 2116 1565 2156
rect 1632 2136 1636 2156
rect 1654 2116 1658 2156
rect 1662 2116 1666 2156
rect 1723 2116 1727 2156
rect 1745 2136 1749 2156
rect 1791 2116 1795 2156
rect 1813 2136 1817 2156
rect 1823 2136 1827 2156
rect 1843 2136 1847 2156
rect 1851 2136 1855 2156
rect 1897 2136 1901 2156
rect 1919 2136 1923 2156
rect 1929 2136 1933 2156
rect 1951 2136 1955 2156
rect 1961 2136 1965 2156
rect 1981 2116 1985 2156
rect 2045 2136 2049 2156
rect 2113 2116 2117 2156
rect 2123 2116 2127 2156
rect 2171 2136 2175 2156
rect 2193 2116 2197 2156
rect 2253 2116 2257 2156
rect 2263 2116 2267 2156
rect 2345 2116 2349 2156
rect 2365 2116 2369 2156
rect 2385 2116 2389 2156
rect 2453 2116 2457 2156
rect 2463 2116 2467 2156
rect 2533 2116 2537 2156
rect 2543 2116 2547 2156
rect 2605 2116 2609 2156
rect 2625 2116 2629 2156
rect 2645 2116 2649 2156
rect 2705 2116 2709 2156
rect 2725 2116 2729 2156
rect 2745 2116 2749 2156
rect 2795 2116 2799 2156
rect 2815 2136 2819 2156
rect 2825 2136 2829 2156
rect 2847 2136 2851 2156
rect 2857 2136 2861 2156
rect 2879 2136 2883 2156
rect 2925 2136 2929 2156
rect 2933 2136 2937 2156
rect 2953 2136 2957 2156
rect 2963 2136 2967 2156
rect 2985 2116 2989 2156
rect 3031 2116 3035 2156
rect 3041 2116 3045 2156
rect 3061 2116 3065 2156
rect 3145 2116 3149 2156
rect 3165 2116 3169 2156
rect 3185 2116 3189 2156
rect 3245 2116 3249 2156
rect 3265 2116 3269 2156
rect 3285 2116 3289 2156
rect 3333 2116 3337 2156
rect 3343 2116 3347 2156
rect 3425 2116 3429 2156
rect 3445 2116 3449 2156
rect 3465 2116 3469 2156
rect 3512 2096 3516 2156
rect 3520 2096 3524 2156
rect 3528 2096 3532 2156
rect 3611 2136 3615 2156
rect 3672 2096 3676 2156
rect 3680 2096 3684 2156
rect 3688 2096 3692 2156
rect 3773 2116 3777 2156
rect 3783 2116 3787 2156
rect 3851 2136 3855 2156
rect 3873 2116 3877 2156
rect 3931 2116 3935 2156
rect 3951 2116 3955 2156
rect 3971 2116 3975 2156
rect 4053 2116 4057 2156
rect 4063 2116 4067 2156
rect 4133 2116 4137 2156
rect 4143 2116 4147 2156
rect 4213 2116 4217 2156
rect 4223 2116 4227 2156
rect 4271 2116 4275 2156
rect 4281 2116 4285 2156
rect 4301 2116 4305 2156
rect 4374 2116 4378 2156
rect 4382 2116 4386 2156
rect 4404 2136 4408 2156
rect 4492 2136 4496 2156
rect 4514 2116 4518 2156
rect 4522 2116 4526 2156
rect 4572 2096 4576 2156
rect 4580 2096 4584 2156
rect 4588 2096 4592 2156
rect 4672 2096 4676 2156
rect 4680 2096 4684 2156
rect 4688 2096 4692 2156
rect 35 1704 39 1744
rect 55 1704 59 1724
rect 65 1704 69 1724
rect 87 1704 91 1724
rect 97 1704 101 1724
rect 119 1704 123 1724
rect 165 1704 169 1724
rect 173 1704 177 1724
rect 193 1704 197 1724
rect 203 1704 207 1724
rect 225 1704 229 1744
rect 271 1704 275 1744
rect 291 1704 295 1744
rect 311 1704 315 1744
rect 385 1704 389 1744
rect 405 1704 409 1744
rect 425 1704 429 1744
rect 485 1704 489 1744
rect 505 1704 509 1744
rect 525 1704 529 1744
rect 585 1704 589 1744
rect 605 1704 609 1744
rect 625 1704 629 1744
rect 671 1704 675 1724
rect 731 1704 735 1724
rect 805 1704 809 1724
rect 825 1704 829 1724
rect 872 1704 876 1764
rect 880 1704 884 1764
rect 888 1704 892 1764
rect 975 1704 979 1744
rect 995 1704 999 1724
rect 1005 1704 1009 1724
rect 1027 1704 1031 1724
rect 1037 1704 1041 1724
rect 1059 1704 1063 1724
rect 1105 1704 1109 1724
rect 1113 1704 1117 1724
rect 1133 1704 1137 1724
rect 1143 1704 1147 1724
rect 1165 1704 1169 1744
rect 1213 1704 1217 1744
rect 1223 1704 1227 1744
rect 1305 1704 1309 1744
rect 1325 1704 1329 1744
rect 1345 1704 1349 1744
rect 1405 1704 1409 1744
rect 1425 1704 1429 1744
rect 1445 1704 1449 1744
rect 1465 1704 1469 1744
rect 1485 1704 1489 1744
rect 1505 1704 1509 1744
rect 1525 1704 1529 1744
rect 1545 1704 1549 1744
rect 1595 1704 1599 1744
rect 1615 1704 1619 1724
rect 1625 1704 1629 1724
rect 1647 1704 1651 1724
rect 1657 1704 1661 1724
rect 1679 1704 1683 1724
rect 1725 1704 1729 1724
rect 1733 1704 1737 1724
rect 1753 1704 1757 1724
rect 1763 1704 1767 1724
rect 1785 1704 1789 1744
rect 1852 1704 1856 1724
rect 1874 1704 1878 1744
rect 1882 1704 1886 1744
rect 1931 1704 1935 1724
rect 1951 1704 1955 1724
rect 2032 1704 2036 1724
rect 2054 1704 2058 1744
rect 2062 1704 2066 1744
rect 2125 1704 2129 1724
rect 2145 1704 2149 1724
rect 2194 1704 2198 1744
rect 2202 1704 2206 1744
rect 2224 1704 2228 1724
rect 2291 1704 2295 1744
rect 2313 1704 2317 1724
rect 2323 1704 2327 1724
rect 2343 1704 2347 1724
rect 2351 1704 2355 1724
rect 2397 1704 2401 1724
rect 2419 1704 2423 1724
rect 2429 1704 2433 1724
rect 2451 1704 2455 1724
rect 2461 1704 2465 1724
rect 2481 1704 2485 1744
rect 2535 1704 2539 1744
rect 2555 1704 2559 1724
rect 2565 1704 2569 1724
rect 2587 1704 2591 1724
rect 2597 1704 2601 1724
rect 2619 1704 2623 1724
rect 2665 1704 2669 1724
rect 2673 1704 2677 1724
rect 2693 1704 2697 1724
rect 2703 1704 2707 1724
rect 2725 1704 2729 1744
rect 2775 1704 2779 1744
rect 2795 1704 2799 1724
rect 2805 1704 2809 1724
rect 2827 1704 2831 1724
rect 2837 1704 2841 1724
rect 2859 1704 2863 1724
rect 2905 1704 2909 1724
rect 2913 1704 2917 1724
rect 2933 1704 2937 1724
rect 2943 1704 2947 1724
rect 2965 1704 2969 1744
rect 3025 1704 3029 1744
rect 3093 1704 3097 1744
rect 3103 1704 3107 1744
rect 3165 1704 3169 1744
rect 3214 1704 3218 1744
rect 3222 1704 3226 1744
rect 3244 1704 3248 1724
rect 3311 1704 3315 1724
rect 3331 1704 3335 1724
rect 3415 1704 3419 1744
rect 3435 1704 3439 1744
rect 3445 1704 3449 1744
rect 3491 1704 3495 1744
rect 3586 1704 3590 1744
rect 3594 1704 3598 1744
rect 3614 1704 3618 1744
rect 3622 1704 3626 1744
rect 3685 1704 3689 1744
rect 3745 1704 3749 1724
rect 3765 1704 3769 1724
rect 3811 1704 3815 1724
rect 3833 1704 3837 1744
rect 3891 1704 3895 1744
rect 3901 1704 3905 1744
rect 3921 1704 3925 1744
rect 4026 1704 4030 1744
rect 4034 1704 4038 1744
rect 4054 1704 4058 1744
rect 4062 1704 4066 1744
rect 4114 1704 4118 1744
rect 4122 1704 4126 1744
rect 4142 1704 4146 1744
rect 4150 1704 4154 1744
rect 4233 1704 4237 1744
rect 4243 1704 4247 1744
rect 4311 1704 4315 1744
rect 4321 1704 4325 1744
rect 4341 1704 4345 1744
rect 4414 1704 4418 1744
rect 4422 1704 4426 1744
rect 4442 1704 4446 1744
rect 4450 1704 4454 1744
rect 4545 1704 4549 1724
rect 4591 1704 4595 1744
rect 4611 1704 4615 1744
rect 4631 1704 4635 1744
rect 4691 1704 4695 1724
rect 31 1636 35 1676
rect 51 1636 55 1676
rect 71 1636 75 1676
rect 91 1636 95 1676
rect 111 1636 115 1676
rect 131 1636 135 1676
rect 151 1636 155 1676
rect 171 1636 175 1676
rect 245 1656 249 1676
rect 265 1656 269 1676
rect 323 1636 327 1676
rect 345 1656 349 1676
rect 395 1636 399 1676
rect 415 1656 419 1676
rect 425 1656 429 1676
rect 447 1656 451 1676
rect 457 1656 461 1676
rect 479 1656 483 1676
rect 525 1656 529 1676
rect 533 1656 537 1676
rect 553 1656 557 1676
rect 563 1656 567 1676
rect 585 1636 589 1676
rect 635 1636 639 1676
rect 655 1656 659 1676
rect 665 1656 669 1676
rect 687 1656 691 1676
rect 697 1656 701 1676
rect 719 1656 723 1676
rect 765 1656 769 1676
rect 773 1656 777 1676
rect 793 1656 797 1676
rect 803 1656 807 1676
rect 825 1636 829 1676
rect 871 1636 875 1676
rect 893 1656 897 1676
rect 903 1656 907 1676
rect 923 1656 927 1676
rect 931 1656 935 1676
rect 977 1656 981 1676
rect 999 1656 1003 1676
rect 1009 1656 1013 1676
rect 1031 1656 1035 1676
rect 1041 1656 1045 1676
rect 1061 1636 1065 1676
rect 1133 1636 1137 1676
rect 1143 1636 1147 1676
rect 1205 1636 1209 1676
rect 1225 1636 1229 1676
rect 1245 1636 1249 1676
rect 1291 1636 1295 1676
rect 1313 1656 1317 1676
rect 1323 1656 1327 1676
rect 1343 1656 1347 1676
rect 1351 1656 1355 1676
rect 1397 1656 1401 1676
rect 1419 1656 1423 1676
rect 1429 1656 1433 1676
rect 1451 1656 1455 1676
rect 1461 1656 1465 1676
rect 1481 1636 1485 1676
rect 1535 1636 1539 1676
rect 1555 1656 1559 1676
rect 1565 1656 1569 1676
rect 1587 1656 1591 1676
rect 1597 1656 1601 1676
rect 1619 1656 1623 1676
rect 1665 1656 1669 1676
rect 1673 1656 1677 1676
rect 1693 1656 1697 1676
rect 1703 1656 1707 1676
rect 1725 1636 1729 1676
rect 1792 1656 1796 1676
rect 1814 1636 1818 1676
rect 1822 1636 1826 1676
rect 1871 1656 1875 1676
rect 1891 1656 1895 1676
rect 1955 1636 1959 1676
rect 1975 1656 1979 1676
rect 1985 1656 1989 1676
rect 2007 1656 2011 1676
rect 2017 1656 2021 1676
rect 2039 1656 2043 1676
rect 2085 1656 2089 1676
rect 2093 1656 2097 1676
rect 2113 1656 2117 1676
rect 2123 1656 2127 1676
rect 2145 1636 2149 1676
rect 2205 1656 2209 1676
rect 2225 1656 2229 1676
rect 2293 1636 2297 1676
rect 2303 1636 2307 1676
rect 2351 1636 2355 1676
rect 2371 1636 2375 1676
rect 2391 1636 2395 1676
rect 2451 1636 2455 1676
rect 2473 1656 2477 1676
rect 2483 1656 2487 1676
rect 2503 1656 2507 1676
rect 2511 1656 2515 1676
rect 2557 1656 2561 1676
rect 2579 1656 2583 1676
rect 2589 1656 2593 1676
rect 2611 1656 2615 1676
rect 2621 1656 2625 1676
rect 2641 1636 2645 1676
rect 2695 1636 2699 1676
rect 2715 1656 2719 1676
rect 2725 1656 2729 1676
rect 2747 1656 2751 1676
rect 2757 1656 2761 1676
rect 2779 1656 2783 1676
rect 2825 1656 2829 1676
rect 2833 1656 2837 1676
rect 2853 1656 2857 1676
rect 2863 1656 2867 1676
rect 2885 1636 2889 1676
rect 2931 1636 2935 1676
rect 2993 1636 2997 1676
rect 3003 1636 3007 1676
rect 3093 1636 3097 1676
rect 3103 1636 3107 1676
rect 3151 1636 3155 1676
rect 3171 1636 3175 1676
rect 3191 1636 3195 1676
rect 3253 1636 3257 1676
rect 3263 1636 3267 1676
rect 3353 1636 3357 1676
rect 3363 1636 3367 1676
rect 3425 1636 3429 1676
rect 3445 1636 3449 1676
rect 3465 1636 3469 1676
rect 3512 1616 3516 1676
rect 3520 1616 3524 1676
rect 3528 1616 3532 1676
rect 3625 1636 3629 1676
rect 3645 1636 3649 1676
rect 3665 1636 3669 1676
rect 3685 1636 3689 1676
rect 3731 1656 3735 1676
rect 3792 1616 3796 1676
rect 3800 1616 3804 1676
rect 3808 1616 3812 1676
rect 3894 1636 3898 1676
rect 3902 1636 3906 1676
rect 3924 1656 3928 1676
rect 3991 1636 3995 1676
rect 4011 1636 4015 1676
rect 4031 1636 4035 1676
rect 4113 1636 4117 1676
rect 4123 1636 4127 1676
rect 4174 1636 4178 1676
rect 4182 1636 4186 1676
rect 4204 1656 4208 1676
rect 4271 1636 4275 1676
rect 4291 1636 4295 1676
rect 4311 1636 4315 1676
rect 4371 1656 4375 1676
rect 4431 1656 4435 1676
rect 4451 1656 4455 1676
rect 4513 1636 4517 1676
rect 4523 1636 4527 1676
rect 4593 1636 4597 1676
rect 4603 1636 4607 1676
rect 4673 1636 4677 1676
rect 4683 1636 4687 1676
rect 31 1224 35 1264
rect 53 1224 57 1244
rect 63 1224 67 1244
rect 83 1224 87 1244
rect 91 1224 95 1244
rect 137 1224 141 1244
rect 159 1224 163 1244
rect 169 1224 173 1244
rect 191 1224 195 1244
rect 201 1224 205 1244
rect 221 1224 225 1264
rect 275 1224 279 1264
rect 295 1224 299 1244
rect 305 1224 309 1244
rect 327 1224 331 1244
rect 337 1224 341 1244
rect 359 1224 363 1244
rect 405 1224 409 1244
rect 413 1224 417 1244
rect 433 1224 437 1244
rect 443 1224 447 1244
rect 465 1224 469 1264
rect 513 1224 517 1264
rect 523 1224 527 1264
rect 605 1224 609 1264
rect 625 1224 629 1264
rect 645 1224 649 1264
rect 705 1224 709 1264
rect 725 1224 729 1264
rect 745 1224 749 1264
rect 803 1224 807 1264
rect 825 1224 829 1244
rect 873 1224 877 1264
rect 883 1224 887 1264
rect 965 1224 969 1264
rect 985 1224 989 1264
rect 1005 1224 1009 1264
rect 1065 1224 1069 1244
rect 1111 1224 1115 1264
rect 1131 1224 1135 1264
rect 1151 1224 1155 1264
rect 1171 1224 1175 1264
rect 1253 1224 1257 1264
rect 1263 1224 1267 1264
rect 1325 1224 1329 1264
rect 1345 1224 1349 1264
rect 1365 1224 1369 1264
rect 1433 1224 1437 1264
rect 1443 1224 1447 1264
rect 1505 1224 1509 1264
rect 1525 1224 1529 1264
rect 1545 1224 1549 1264
rect 1591 1224 1595 1244
rect 1613 1224 1617 1264
rect 1673 1224 1677 1264
rect 1683 1224 1687 1264
rect 1765 1224 1769 1264
rect 1785 1224 1789 1264
rect 1805 1224 1809 1264
rect 1851 1224 1855 1264
rect 1873 1224 1877 1244
rect 1883 1224 1887 1244
rect 1903 1224 1907 1244
rect 1911 1224 1915 1244
rect 1957 1224 1961 1244
rect 1979 1224 1983 1244
rect 1989 1224 1993 1244
rect 2011 1224 2015 1244
rect 2021 1224 2025 1244
rect 2041 1224 2045 1264
rect 2091 1224 2095 1244
rect 2151 1224 2155 1264
rect 2171 1224 2175 1264
rect 2191 1224 2195 1264
rect 2273 1224 2277 1264
rect 2283 1224 2287 1264
rect 2345 1224 2349 1244
rect 2365 1224 2369 1244
rect 2425 1224 2429 1244
rect 2471 1224 2475 1244
rect 2491 1224 2495 1244
rect 2551 1224 2555 1264
rect 2573 1224 2577 1244
rect 2583 1224 2587 1244
rect 2603 1224 2607 1244
rect 2611 1224 2615 1244
rect 2657 1224 2661 1244
rect 2679 1224 2683 1244
rect 2689 1224 2693 1244
rect 2711 1224 2715 1244
rect 2721 1224 2725 1244
rect 2741 1224 2745 1264
rect 2791 1224 2795 1244
rect 2811 1224 2815 1244
rect 2885 1224 2889 1264
rect 2931 1224 2935 1264
rect 2951 1224 2955 1264
rect 2971 1224 2975 1264
rect 3031 1224 3035 1264
rect 3051 1224 3055 1264
rect 3071 1224 3075 1264
rect 3131 1224 3135 1264
rect 3151 1224 3155 1264
rect 3171 1224 3175 1264
rect 3231 1224 3235 1264
rect 3241 1224 3245 1264
rect 3261 1224 3265 1264
rect 3345 1224 3349 1244
rect 3365 1224 3369 1244
rect 3412 1224 3416 1284
rect 3420 1224 3424 1284
rect 3428 1224 3432 1284
rect 3525 1224 3529 1264
rect 3545 1224 3549 1264
rect 3565 1224 3569 1264
rect 3611 1224 3615 1264
rect 3631 1224 3635 1264
rect 3651 1224 3655 1264
rect 3733 1224 3737 1264
rect 3743 1224 3747 1264
rect 3813 1224 3817 1264
rect 3823 1224 3827 1264
rect 3871 1224 3875 1264
rect 3881 1224 3885 1264
rect 3901 1224 3905 1264
rect 3985 1224 3989 1264
rect 4005 1224 4009 1264
rect 4025 1224 4029 1264
rect 4071 1224 4075 1244
rect 4153 1224 4157 1264
rect 4163 1224 4167 1264
rect 4233 1224 4237 1264
rect 4243 1224 4247 1264
rect 4305 1224 4309 1244
rect 4325 1224 4329 1244
rect 4385 1224 4389 1264
rect 4405 1224 4409 1264
rect 4425 1224 4429 1264
rect 4471 1224 4475 1264
rect 4491 1224 4495 1264
rect 4511 1224 4515 1264
rect 4592 1224 4596 1244
rect 4614 1224 4618 1264
rect 4622 1224 4626 1264
rect 4673 1224 4677 1264
rect 4683 1224 4687 1264
rect 31 1176 35 1196
rect 113 1156 117 1196
rect 123 1156 127 1196
rect 185 1156 189 1196
rect 205 1156 209 1196
rect 225 1156 229 1196
rect 274 1156 278 1196
rect 282 1156 286 1196
rect 302 1156 306 1196
rect 310 1156 314 1196
rect 412 1176 416 1196
rect 434 1156 438 1196
rect 442 1156 446 1196
rect 505 1156 509 1196
rect 525 1176 529 1196
rect 545 1176 549 1196
rect 591 1176 595 1196
rect 611 1176 615 1196
rect 695 1156 699 1196
rect 715 1156 719 1196
rect 725 1156 729 1196
rect 783 1156 787 1196
rect 805 1176 809 1196
rect 865 1176 869 1196
rect 885 1176 889 1196
rect 945 1176 949 1196
rect 1005 1176 1009 1196
rect 1051 1176 1055 1196
rect 1071 1176 1075 1196
rect 1131 1176 1135 1196
rect 1205 1176 1209 1196
rect 1225 1176 1229 1196
rect 1274 1156 1278 1196
rect 1282 1156 1286 1196
rect 1304 1176 1308 1196
rect 1375 1156 1379 1196
rect 1395 1176 1399 1196
rect 1405 1176 1409 1196
rect 1427 1176 1431 1196
rect 1437 1176 1441 1196
rect 1459 1176 1463 1196
rect 1505 1176 1509 1196
rect 1513 1176 1517 1196
rect 1533 1176 1537 1196
rect 1543 1176 1547 1196
rect 1565 1156 1569 1196
rect 1625 1176 1629 1196
rect 1673 1156 1677 1196
rect 1683 1156 1687 1196
rect 1751 1176 1755 1196
rect 1771 1176 1775 1196
rect 1835 1156 1839 1196
rect 1855 1176 1859 1196
rect 1865 1176 1869 1196
rect 1887 1176 1891 1196
rect 1897 1176 1901 1196
rect 1919 1176 1923 1196
rect 1965 1176 1969 1196
rect 1973 1176 1977 1196
rect 1993 1176 1997 1196
rect 2003 1176 2007 1196
rect 2025 1156 2029 1196
rect 2085 1176 2089 1196
rect 2131 1176 2135 1196
rect 2151 1176 2155 1196
rect 2211 1176 2215 1196
rect 2231 1176 2235 1196
rect 2305 1176 2309 1196
rect 2351 1156 2355 1196
rect 2373 1176 2377 1196
rect 2383 1176 2387 1196
rect 2403 1176 2407 1196
rect 2411 1176 2415 1196
rect 2457 1176 2461 1196
rect 2479 1176 2483 1196
rect 2489 1176 2493 1196
rect 2511 1176 2515 1196
rect 2521 1176 2525 1196
rect 2541 1156 2545 1196
rect 2591 1176 2595 1196
rect 2651 1156 2655 1196
rect 2671 1156 2675 1196
rect 2691 1156 2695 1196
rect 2751 1156 2755 1196
rect 2771 1156 2775 1196
rect 2791 1156 2795 1196
rect 2811 1156 2815 1196
rect 2871 1176 2875 1196
rect 2891 1176 2895 1196
rect 2973 1156 2977 1196
rect 2983 1156 2987 1196
rect 3031 1156 3035 1196
rect 3041 1156 3045 1196
rect 3061 1156 3065 1196
rect 3131 1156 3135 1196
rect 3151 1156 3155 1196
rect 3171 1156 3175 1196
rect 3231 1176 3235 1196
rect 3251 1176 3255 1196
rect 3271 1156 3275 1196
rect 3353 1156 3357 1196
rect 3363 1156 3367 1196
rect 3433 1156 3437 1196
rect 3443 1156 3447 1196
rect 3493 1156 3497 1196
rect 3503 1156 3507 1196
rect 3573 1156 3577 1196
rect 3583 1156 3587 1196
rect 3651 1156 3655 1196
rect 3671 1156 3675 1196
rect 3691 1156 3695 1196
rect 3788 1136 3792 1196
rect 3796 1136 3800 1196
rect 3804 1136 3808 1196
rect 3854 1156 3858 1196
rect 3862 1156 3866 1196
rect 3884 1176 3888 1196
rect 3965 1176 3969 1196
rect 4048 1136 4052 1196
rect 4056 1136 4060 1196
rect 4064 1136 4068 1196
rect 4114 1156 4118 1196
rect 4122 1156 4126 1196
rect 4144 1176 4148 1196
rect 4211 1176 4215 1196
rect 4292 1176 4296 1196
rect 4314 1156 4318 1196
rect 4322 1156 4326 1196
rect 4385 1156 4389 1196
rect 4405 1156 4409 1196
rect 4425 1156 4429 1196
rect 4471 1156 4475 1196
rect 4491 1156 4495 1196
rect 4511 1156 4515 1196
rect 4571 1176 4575 1196
rect 4591 1176 4595 1196
rect 4673 1156 4677 1196
rect 4683 1156 4687 1196
rect 4745 1176 4749 1196
rect 35 744 39 784
rect 55 744 59 764
rect 65 744 69 764
rect 87 744 91 764
rect 97 744 101 764
rect 119 744 123 764
rect 165 744 169 764
rect 173 744 177 764
rect 193 744 197 764
rect 203 744 207 764
rect 225 744 229 784
rect 273 744 277 784
rect 283 744 287 784
rect 365 744 369 784
rect 385 744 389 784
rect 405 744 409 784
rect 455 744 459 784
rect 475 744 479 764
rect 485 744 489 764
rect 507 744 511 764
rect 517 744 521 764
rect 539 744 543 764
rect 585 744 589 764
rect 593 744 597 764
rect 613 744 617 764
rect 623 744 627 764
rect 645 744 649 784
rect 693 744 697 784
rect 703 744 707 784
rect 785 744 789 784
rect 805 744 809 784
rect 825 744 829 784
rect 885 744 889 784
rect 905 744 909 784
rect 925 744 929 784
rect 985 744 989 764
rect 1045 744 1049 764
rect 1065 744 1069 764
rect 1111 744 1115 764
rect 1131 744 1135 764
rect 1213 744 1217 784
rect 1223 744 1227 784
rect 1293 744 1297 784
rect 1303 744 1307 784
rect 1373 744 1377 784
rect 1383 744 1387 784
rect 1452 744 1456 764
rect 1474 744 1478 784
rect 1482 744 1486 784
rect 1555 744 1559 784
rect 1575 744 1579 784
rect 1585 744 1589 784
rect 1634 744 1638 784
rect 1642 744 1646 784
rect 1664 744 1668 764
rect 1731 744 1735 784
rect 1751 744 1755 784
rect 1771 744 1775 784
rect 1791 744 1795 784
rect 1811 744 1815 784
rect 1831 744 1835 784
rect 1851 744 1855 784
rect 1871 744 1875 784
rect 1953 744 1957 784
rect 1963 744 1967 784
rect 2025 744 2029 764
rect 2045 744 2049 764
rect 2091 744 2095 784
rect 2111 744 2115 784
rect 2131 744 2135 784
rect 2191 744 2195 784
rect 2211 744 2215 784
rect 2231 744 2235 784
rect 2291 744 2295 784
rect 2311 744 2315 784
rect 2331 744 2335 784
rect 2393 744 2397 784
rect 2403 744 2407 784
rect 2485 744 2489 764
rect 2531 744 2535 784
rect 2553 744 2557 764
rect 2563 744 2567 764
rect 2583 744 2587 764
rect 2591 744 2595 764
rect 2637 744 2641 764
rect 2659 744 2663 764
rect 2669 744 2673 764
rect 2691 744 2695 764
rect 2701 744 2705 764
rect 2721 744 2725 784
rect 2785 744 2789 784
rect 2805 744 2809 784
rect 2825 744 2829 784
rect 2885 744 2889 764
rect 2931 744 2935 764
rect 2992 744 2996 804
rect 3000 744 3004 804
rect 3008 744 3012 804
rect 3091 744 3095 764
rect 3173 744 3177 784
rect 3183 744 3187 784
rect 3231 744 3235 764
rect 3251 744 3255 764
rect 3271 744 3275 784
rect 3333 744 3337 784
rect 3343 744 3347 784
rect 3413 744 3417 784
rect 3423 744 3427 784
rect 3505 744 3509 764
rect 3525 744 3529 764
rect 3573 744 3577 784
rect 3583 744 3587 784
rect 3688 744 3692 804
rect 3696 744 3700 804
rect 3704 744 3708 804
rect 3788 744 3792 804
rect 3796 744 3800 804
rect 3804 744 3808 804
rect 3853 744 3857 784
rect 3863 744 3867 784
rect 3968 744 3972 804
rect 3976 744 3980 804
rect 3984 744 3988 804
rect 4045 744 4049 764
rect 4105 744 4109 784
rect 4125 744 4129 784
rect 4145 744 4149 784
rect 4205 744 4209 784
rect 4225 744 4229 784
rect 4245 744 4249 784
rect 4312 744 4316 764
rect 4334 744 4338 784
rect 4342 744 4346 784
rect 4392 744 4396 804
rect 4400 744 4404 804
rect 4408 744 4412 804
rect 4528 744 4532 804
rect 4536 744 4540 804
rect 4544 744 4548 804
rect 4612 744 4616 764
rect 4634 744 4638 784
rect 4642 744 4646 784
rect 4692 744 4696 804
rect 4700 744 4704 804
rect 4708 744 4712 804
rect 35 676 39 716
rect 55 696 59 716
rect 65 696 69 716
rect 87 696 91 716
rect 97 696 101 716
rect 119 696 123 716
rect 165 696 169 716
rect 173 696 177 716
rect 193 696 197 716
rect 203 696 207 716
rect 225 676 229 716
rect 271 696 275 716
rect 331 676 335 716
rect 351 676 355 716
rect 371 676 375 716
rect 433 676 437 716
rect 443 676 447 716
rect 511 696 515 716
rect 533 676 537 716
rect 605 696 609 716
rect 651 676 655 716
rect 673 696 677 716
rect 683 696 687 716
rect 703 696 707 716
rect 711 696 715 716
rect 757 696 761 716
rect 779 696 783 716
rect 789 696 793 716
rect 811 696 815 716
rect 821 696 825 716
rect 841 676 845 716
rect 891 676 895 716
rect 911 676 915 716
rect 931 676 935 716
rect 1005 696 1009 716
rect 1025 696 1029 716
rect 1071 696 1075 716
rect 1091 696 1095 716
rect 1111 676 1115 716
rect 1185 676 1189 716
rect 1205 676 1209 716
rect 1225 676 1229 716
rect 1295 676 1299 716
rect 1315 676 1319 716
rect 1325 676 1329 716
rect 1371 696 1375 716
rect 1391 696 1395 716
rect 1451 696 1455 716
rect 1473 676 1477 716
rect 1535 676 1539 716
rect 1555 696 1559 716
rect 1565 696 1569 716
rect 1587 696 1591 716
rect 1597 696 1601 716
rect 1619 696 1623 716
rect 1665 696 1669 716
rect 1673 696 1677 716
rect 1693 696 1697 716
rect 1703 696 1707 716
rect 1725 676 1729 716
rect 1771 696 1775 716
rect 1793 676 1797 716
rect 1865 696 1869 716
rect 1885 696 1889 716
rect 1945 696 1949 716
rect 1965 696 1969 716
rect 2025 696 2029 716
rect 2071 696 2075 716
rect 2091 696 2095 716
rect 2151 676 2155 716
rect 2173 696 2177 716
rect 2183 696 2187 716
rect 2203 696 2207 716
rect 2211 696 2215 716
rect 2257 696 2261 716
rect 2279 696 2283 716
rect 2289 696 2293 716
rect 2311 696 2315 716
rect 2321 696 2325 716
rect 2341 676 2345 716
rect 2394 676 2398 716
rect 2402 676 2406 716
rect 2422 676 2426 716
rect 2430 676 2434 716
rect 2525 676 2529 716
rect 2545 696 2549 716
rect 2565 696 2569 716
rect 2632 696 2636 716
rect 2654 676 2658 716
rect 2662 676 2666 716
rect 2732 696 2736 716
rect 2754 676 2758 716
rect 2762 676 2766 716
rect 2811 696 2815 716
rect 2885 676 2889 716
rect 2905 676 2909 716
rect 2925 676 2929 716
rect 2971 676 2975 716
rect 2991 676 2995 716
rect 3011 676 3015 716
rect 3073 676 3077 716
rect 3083 676 3087 716
rect 3165 696 3169 716
rect 3211 696 3215 716
rect 3308 656 3312 716
rect 3316 656 3320 716
rect 3324 656 3328 716
rect 3385 696 3389 716
rect 3405 696 3409 716
rect 3451 676 3455 716
rect 3471 676 3475 716
rect 3491 676 3495 716
rect 3554 676 3558 716
rect 3562 676 3566 716
rect 3584 696 3588 716
rect 3672 696 3676 716
rect 3694 676 3698 716
rect 3702 676 3706 716
rect 3786 676 3790 716
rect 3794 676 3798 716
rect 3814 676 3818 716
rect 3822 676 3826 716
rect 3908 656 3912 716
rect 3916 656 3920 716
rect 3924 656 3928 716
rect 4008 656 4012 716
rect 4016 656 4020 716
rect 4024 656 4028 716
rect 4071 696 4075 716
rect 4132 656 4136 716
rect 4140 656 4144 716
rect 4148 656 4152 716
rect 4232 656 4236 716
rect 4240 656 4244 716
rect 4248 656 4252 716
rect 4368 656 4372 716
rect 4376 656 4380 716
rect 4384 656 4388 716
rect 4468 656 4472 716
rect 4476 656 4480 716
rect 4484 656 4488 716
rect 4531 696 4535 716
rect 4605 676 4609 716
rect 4625 676 4629 716
rect 4645 676 4649 716
rect 4691 676 4695 716
rect 4711 676 4715 716
rect 4731 676 4735 716
rect 35 264 39 304
rect 55 264 59 284
rect 65 264 69 284
rect 87 264 91 284
rect 97 264 101 284
rect 119 264 123 284
rect 165 264 169 284
rect 173 264 177 284
rect 193 264 197 284
rect 203 264 207 284
rect 225 264 229 304
rect 273 264 277 304
rect 283 264 287 304
rect 365 264 369 304
rect 385 264 389 304
rect 405 264 409 304
rect 451 264 455 284
rect 513 264 517 304
rect 523 264 527 304
rect 605 264 609 304
rect 625 264 629 304
rect 645 264 649 304
rect 691 264 695 304
rect 711 264 715 304
rect 731 264 735 304
rect 791 264 795 304
rect 811 264 815 304
rect 831 264 835 304
rect 905 264 909 304
rect 925 264 929 304
rect 945 264 949 304
rect 991 264 995 284
rect 1053 264 1057 304
rect 1063 264 1067 304
rect 1152 264 1156 284
rect 1174 264 1178 304
rect 1182 264 1186 304
rect 1245 264 1249 284
rect 1305 264 1309 304
rect 1325 264 1329 304
rect 1345 264 1349 304
rect 1405 264 1409 284
rect 1425 264 1429 284
rect 1471 264 1475 304
rect 1491 264 1495 304
rect 1511 264 1515 304
rect 1573 264 1577 304
rect 1583 264 1587 304
rect 1651 264 1655 304
rect 1673 264 1677 284
rect 1683 264 1687 284
rect 1703 264 1707 284
rect 1711 264 1715 284
rect 1757 264 1761 284
rect 1779 264 1783 284
rect 1789 264 1793 284
rect 1811 264 1815 284
rect 1821 264 1825 284
rect 1841 264 1845 304
rect 1913 264 1917 304
rect 1923 264 1927 304
rect 1985 264 1989 304
rect 2005 264 2009 304
rect 2025 264 2029 304
rect 2075 264 2079 304
rect 2095 264 2099 284
rect 2105 264 2109 284
rect 2127 264 2131 284
rect 2137 264 2141 284
rect 2159 264 2163 284
rect 2205 264 2209 284
rect 2213 264 2217 284
rect 2233 264 2237 284
rect 2243 264 2247 284
rect 2265 264 2269 304
rect 2325 264 2329 284
rect 2371 264 2375 284
rect 2391 264 2395 284
rect 2451 264 2455 284
rect 2533 264 2537 304
rect 2543 264 2547 304
rect 2591 264 2595 304
rect 2613 264 2617 284
rect 2623 264 2627 284
rect 2643 264 2647 284
rect 2651 264 2655 284
rect 2697 264 2701 284
rect 2719 264 2723 284
rect 2729 264 2733 284
rect 2751 264 2755 284
rect 2761 264 2765 284
rect 2781 264 2785 304
rect 2833 264 2837 304
rect 2843 264 2847 304
rect 2914 264 2918 304
rect 2922 264 2926 304
rect 2942 264 2946 304
rect 2950 264 2954 304
rect 3031 264 3035 284
rect 3051 264 3055 284
rect 3111 264 3115 284
rect 3208 264 3212 324
rect 3216 264 3220 324
rect 3224 264 3228 324
rect 3308 264 3312 324
rect 3316 264 3320 324
rect 3324 264 3328 324
rect 3371 264 3375 304
rect 3391 264 3395 304
rect 3411 264 3415 304
rect 3485 264 3489 284
rect 3533 264 3537 304
rect 3543 264 3547 304
rect 3613 264 3617 304
rect 3623 264 3627 304
rect 3691 264 3695 304
rect 3711 264 3715 304
rect 3731 264 3735 304
rect 3805 264 3809 284
rect 3825 264 3829 284
rect 3885 264 3889 284
rect 3905 264 3909 284
rect 3951 264 3955 304
rect 3961 264 3965 304
rect 3981 264 3985 304
rect 4051 264 4055 284
rect 4071 264 4075 284
rect 4152 264 4156 284
rect 4174 264 4178 304
rect 4182 264 4186 304
rect 4268 264 4272 324
rect 4276 264 4280 324
rect 4284 264 4288 324
rect 4334 264 4338 304
rect 4342 264 4346 304
rect 4364 264 4368 284
rect 4431 264 4435 284
rect 4505 264 4509 304
rect 4525 264 4529 304
rect 4545 264 4549 304
rect 4591 264 4595 284
rect 4651 264 4655 284
rect 4711 264 4715 284
rect 35 196 39 236
rect 55 216 59 236
rect 65 216 69 236
rect 87 216 91 236
rect 97 216 101 236
rect 119 216 123 236
rect 165 216 169 236
rect 173 216 177 236
rect 193 216 197 236
rect 203 216 207 236
rect 225 196 229 236
rect 274 196 278 236
rect 282 196 286 236
rect 302 196 306 236
rect 310 196 314 236
rect 391 216 395 236
rect 411 216 415 236
rect 472 176 476 236
rect 480 176 484 236
rect 488 176 492 236
rect 585 196 589 236
rect 605 216 609 236
rect 625 216 629 236
rect 692 216 696 236
rect 714 196 718 236
rect 722 196 726 236
rect 771 196 775 236
rect 793 216 797 236
rect 803 216 807 236
rect 823 216 827 236
rect 831 216 835 236
rect 877 216 881 236
rect 899 216 903 236
rect 909 216 913 236
rect 931 216 935 236
rect 941 216 945 236
rect 961 196 965 236
rect 1025 196 1029 236
rect 1045 196 1049 236
rect 1065 196 1069 236
rect 1125 216 1129 236
rect 1185 216 1189 236
rect 1205 216 1209 236
rect 1265 216 1269 236
rect 1325 196 1329 236
rect 1345 196 1349 236
rect 1365 196 1369 236
rect 1425 216 1429 236
rect 1485 216 1489 236
rect 1531 216 1535 236
rect 1551 216 1555 236
rect 1632 216 1636 236
rect 1654 196 1658 236
rect 1662 196 1666 236
rect 1715 196 1719 236
rect 1735 216 1739 236
rect 1745 216 1749 236
rect 1767 216 1771 236
rect 1777 216 1781 236
rect 1799 216 1803 236
rect 1845 216 1849 236
rect 1853 216 1857 236
rect 1873 216 1877 236
rect 1883 216 1887 236
rect 1905 196 1909 236
rect 1965 196 1969 236
rect 1985 196 1989 236
rect 2005 196 2009 236
rect 2051 216 2055 236
rect 2111 216 2115 236
rect 2131 216 2135 236
rect 2191 216 2195 236
rect 2211 216 2215 236
rect 2285 216 2289 236
rect 2305 216 2309 236
rect 2351 216 2355 236
rect 2371 216 2375 236
rect 2445 216 2449 236
rect 2491 196 2495 236
rect 2513 216 2517 236
rect 2523 216 2527 236
rect 2543 216 2547 236
rect 2551 216 2555 236
rect 2597 216 2601 236
rect 2619 216 2623 236
rect 2629 216 2633 236
rect 2651 216 2655 236
rect 2661 216 2665 236
rect 2681 196 2685 236
rect 2731 196 2735 236
rect 2753 216 2757 236
rect 2763 216 2767 236
rect 2783 216 2787 236
rect 2791 216 2795 236
rect 2837 216 2841 236
rect 2859 216 2863 236
rect 2869 216 2873 236
rect 2891 216 2895 236
rect 2901 216 2905 236
rect 2921 196 2925 236
rect 2971 196 2975 236
rect 2991 196 2995 236
rect 3011 196 3015 236
rect 3031 196 3035 236
rect 3105 196 3109 236
rect 3125 216 3129 236
rect 3145 216 3149 236
rect 3191 196 3195 236
rect 3211 196 3215 236
rect 3231 196 3235 236
rect 3305 216 3309 236
rect 3353 196 3357 236
rect 3363 196 3367 236
rect 3468 176 3472 236
rect 3476 176 3480 236
rect 3484 176 3488 236
rect 3545 216 3549 236
rect 3612 216 3616 236
rect 3634 196 3638 236
rect 3642 196 3646 236
rect 3705 216 3709 236
rect 3725 216 3729 236
rect 3771 216 3775 236
rect 3831 196 3835 236
rect 3851 196 3855 236
rect 3871 196 3875 236
rect 3931 216 3935 236
rect 3951 216 3955 236
rect 4048 176 4052 236
rect 4056 176 4060 236
rect 4064 176 4068 236
rect 4113 196 4117 236
rect 4123 196 4127 236
rect 4228 176 4232 236
rect 4236 176 4240 236
rect 4244 176 4248 236
rect 4313 196 4317 236
rect 4323 196 4327 236
rect 4408 176 4412 236
rect 4416 176 4420 236
rect 4424 176 4428 236
rect 4473 196 4477 236
rect 4483 196 4487 236
rect 4552 176 4556 236
rect 4560 176 4564 236
rect 4568 176 4572 236
rect 4672 216 4676 236
rect 4694 196 4698 236
rect 4702 196 4706 236
<< ptransistor >>
rect 43 4344 47 4424
rect 65 4344 69 4384
rect 125 4344 129 4384
rect 145 4344 149 4384
rect 210 4344 214 4384
rect 232 4344 236 4424
rect 240 4344 244 4424
rect 291 4344 295 4384
rect 313 4344 317 4424
rect 397 4344 401 4424
rect 405 4344 409 4424
rect 477 4344 481 4424
rect 485 4344 489 4424
rect 531 4344 535 4384
rect 553 4344 557 4424
rect 625 4344 629 4384
rect 671 4344 675 4424
rect 679 4344 683 4424
rect 751 4344 755 4384
rect 811 4344 815 4424
rect 833 4344 837 4364
rect 841 4344 845 4364
rect 861 4344 865 4384
rect 869 4344 873 4384
rect 915 4344 919 4384
rect 935 4344 939 4384
rect 947 4344 951 4384
rect 967 4344 971 4384
rect 981 4344 985 4384
rect 1001 4344 1005 4424
rect 1056 4344 1060 4424
rect 1064 4344 1068 4424
rect 1086 4344 1090 4384
rect 1151 4344 1155 4424
rect 1173 4344 1177 4364
rect 1181 4344 1185 4364
rect 1201 4344 1205 4384
rect 1209 4344 1213 4384
rect 1255 4344 1259 4384
rect 1275 4344 1279 4384
rect 1287 4344 1291 4384
rect 1307 4344 1311 4384
rect 1321 4344 1325 4384
rect 1341 4344 1345 4424
rect 1396 4344 1400 4424
rect 1404 4344 1408 4424
rect 1426 4344 1430 4384
rect 1495 4344 1499 4424
rect 1515 4344 1519 4384
rect 1529 4344 1533 4384
rect 1549 4344 1553 4384
rect 1561 4344 1565 4384
rect 1581 4344 1585 4384
rect 1627 4344 1631 4384
rect 1635 4344 1639 4384
rect 1655 4344 1659 4364
rect 1663 4344 1667 4364
rect 1685 4344 1689 4424
rect 1731 4344 1735 4384
rect 1751 4344 1755 4384
rect 1811 4344 1815 4424
rect 1833 4344 1837 4364
rect 1841 4344 1845 4364
rect 1861 4344 1865 4384
rect 1869 4344 1873 4384
rect 1915 4344 1919 4384
rect 1935 4344 1939 4384
rect 1947 4344 1951 4384
rect 1967 4344 1971 4384
rect 1981 4344 1985 4384
rect 2001 4344 2005 4424
rect 2051 4344 2055 4424
rect 2061 4344 2065 4424
rect 2091 4344 2095 4424
rect 2101 4344 2105 4424
rect 2185 4344 2189 4384
rect 2205 4344 2209 4384
rect 2225 4344 2229 4384
rect 2290 4344 2294 4384
rect 2312 4344 2316 4424
rect 2320 4344 2324 4424
rect 2385 4344 2389 4384
rect 2431 4344 2435 4424
rect 2439 4344 2443 4424
rect 2525 4344 2529 4384
rect 2576 4344 2580 4424
rect 2584 4344 2588 4424
rect 2606 4344 2610 4384
rect 2671 4344 2675 4384
rect 2693 4344 2697 4424
rect 2751 4344 2755 4384
rect 2773 4344 2777 4424
rect 2843 4344 2847 4424
rect 2865 4344 2869 4384
rect 2925 4344 2929 4384
rect 2945 4344 2949 4384
rect 2965 4344 2969 4384
rect 3021 4344 3025 4424
rect 3043 4344 3047 4384
rect 3065 4344 3069 4384
rect 3123 4344 3127 4424
rect 3145 4344 3149 4384
rect 3205 4344 3209 4384
rect 3225 4344 3229 4384
rect 3245 4344 3249 4384
rect 3291 4344 3295 4384
rect 3311 4344 3315 4384
rect 3371 4344 3375 4424
rect 3391 4344 3395 4424
rect 3411 4344 3415 4424
rect 3471 4344 3475 4384
rect 3531 4344 3535 4384
rect 3551 4344 3555 4384
rect 3611 4344 3615 4384
rect 3631 4344 3635 4384
rect 3651 4344 3655 4384
rect 3711 4344 3715 4424
rect 3731 4344 3735 4424
rect 3751 4344 3755 4424
rect 3816 4344 3820 4424
rect 3824 4344 3828 4424
rect 3846 4344 3850 4384
rect 3930 4344 3934 4384
rect 3952 4344 3956 4424
rect 3960 4344 3964 4424
rect 4025 4344 4029 4384
rect 4045 4344 4049 4384
rect 4065 4344 4069 4384
rect 4125 4344 4129 4384
rect 4145 4344 4149 4384
rect 4165 4344 4169 4384
rect 4211 4344 4215 4424
rect 4231 4344 4235 4424
rect 4251 4344 4255 4424
rect 4311 4344 4315 4384
rect 4331 4344 4335 4384
rect 4405 4344 4409 4424
rect 4425 4344 4429 4424
rect 4445 4344 4449 4424
rect 4505 4344 4509 4384
rect 4551 4344 4555 4384
rect 4571 4344 4575 4384
rect 4591 4344 4595 4384
rect 4651 4344 4655 4384
rect 4671 4344 4675 4384
rect 4691 4344 4695 4384
rect 50 4276 54 4316
rect 72 4236 76 4316
rect 80 4236 84 4316
rect 141 4236 145 4316
rect 163 4276 167 4316
rect 185 4276 189 4316
rect 231 4236 235 4316
rect 239 4236 243 4316
rect 325 4236 329 4316
rect 345 4236 349 4316
rect 365 4236 369 4316
rect 411 4276 415 4316
rect 433 4276 437 4316
rect 455 4236 459 4316
rect 525 4236 529 4316
rect 545 4236 549 4316
rect 565 4236 569 4316
rect 611 4276 615 4316
rect 631 4276 635 4316
rect 651 4276 655 4316
rect 711 4236 715 4316
rect 731 4236 735 4316
rect 751 4236 755 4316
rect 811 4276 815 4316
rect 833 4276 837 4316
rect 855 4236 859 4316
rect 930 4276 934 4316
rect 952 4236 956 4316
rect 960 4236 964 4316
rect 1025 4276 1029 4316
rect 1071 4236 1075 4316
rect 1079 4236 1083 4316
rect 1151 4236 1155 4316
rect 1159 4236 1163 4316
rect 1231 4236 1235 4316
rect 1239 4236 1243 4316
rect 1311 4276 1315 4316
rect 1371 4236 1375 4316
rect 1393 4296 1397 4316
rect 1401 4296 1405 4316
rect 1421 4276 1425 4316
rect 1429 4276 1433 4316
rect 1475 4276 1479 4316
rect 1495 4276 1499 4316
rect 1507 4276 1511 4316
rect 1527 4276 1531 4316
rect 1541 4276 1545 4316
rect 1561 4236 1565 4316
rect 1616 4236 1620 4316
rect 1624 4236 1628 4316
rect 1646 4276 1650 4316
rect 1711 4236 1715 4316
rect 1719 4236 1723 4316
rect 1805 4276 1809 4316
rect 1851 4236 1855 4316
rect 1873 4296 1877 4316
rect 1881 4296 1885 4316
rect 1901 4276 1905 4316
rect 1909 4276 1913 4316
rect 1955 4276 1959 4316
rect 1975 4276 1979 4316
rect 1987 4276 1991 4316
rect 2007 4276 2011 4316
rect 2021 4276 2025 4316
rect 2041 4236 2045 4316
rect 2105 4276 2109 4316
rect 2125 4276 2129 4316
rect 2171 4236 2175 4316
rect 2181 4236 2185 4316
rect 2201 4236 2205 4316
rect 2285 4236 2289 4316
rect 2305 4236 2309 4316
rect 2325 4236 2329 4316
rect 2345 4236 2349 4316
rect 2391 4276 2395 4316
rect 2411 4276 2415 4316
rect 2490 4276 2494 4316
rect 2512 4236 2516 4316
rect 2520 4236 2524 4316
rect 2597 4236 2601 4316
rect 2605 4236 2609 4316
rect 2651 4236 2655 4316
rect 2671 4236 2675 4316
rect 2691 4236 2695 4316
rect 2765 4236 2769 4316
rect 2785 4236 2789 4316
rect 2805 4236 2809 4316
rect 2851 4276 2855 4316
rect 2873 4236 2877 4316
rect 2945 4276 2949 4316
rect 2965 4276 2969 4316
rect 2985 4276 2989 4316
rect 3045 4276 3049 4316
rect 3065 4276 3069 4316
rect 3085 4276 3089 4316
rect 3131 4276 3135 4316
rect 3151 4276 3155 4316
rect 3225 4276 3229 4316
rect 3285 4276 3289 4316
rect 3305 4276 3309 4316
rect 3325 4276 3329 4316
rect 3385 4276 3389 4316
rect 3405 4276 3409 4316
rect 3425 4276 3429 4316
rect 3485 4276 3489 4316
rect 3505 4276 3509 4316
rect 3525 4276 3529 4316
rect 3585 4276 3589 4316
rect 3605 4276 3609 4316
rect 3625 4276 3629 4316
rect 3671 4276 3675 4316
rect 3691 4276 3695 4316
rect 3711 4276 3715 4316
rect 3771 4236 3775 4316
rect 3791 4236 3795 4316
rect 3811 4236 3815 4316
rect 3876 4236 3880 4316
rect 3884 4236 3888 4316
rect 3906 4276 3910 4316
rect 3971 4276 3975 4316
rect 4031 4236 4035 4316
rect 4051 4236 4055 4316
rect 4071 4236 4075 4316
rect 4145 4276 4149 4316
rect 4165 4276 4169 4316
rect 4185 4276 4189 4316
rect 4231 4276 4235 4316
rect 4251 4276 4255 4316
rect 4271 4276 4275 4316
rect 4331 4236 4335 4316
rect 4351 4236 4355 4316
rect 4371 4236 4375 4316
rect 4436 4236 4440 4316
rect 4444 4236 4448 4316
rect 4466 4276 4470 4316
rect 4531 4236 4535 4316
rect 4551 4236 4555 4316
rect 4571 4236 4575 4316
rect 4591 4236 4595 4316
rect 4677 4236 4681 4316
rect 4685 4236 4689 4316
rect 45 3864 49 3904
rect 65 3864 69 3904
rect 125 3864 129 3904
rect 145 3864 149 3904
rect 217 3864 221 3944
rect 225 3864 229 3944
rect 276 3864 280 3944
rect 284 3864 288 3944
rect 306 3864 310 3904
rect 385 3864 389 3904
rect 445 3864 449 3904
rect 517 3864 521 3944
rect 525 3864 529 3944
rect 571 3864 575 3904
rect 593 3864 597 3904
rect 615 3864 619 3944
rect 676 3864 680 3944
rect 684 3864 688 3944
rect 706 3864 710 3904
rect 771 3864 775 3904
rect 836 3864 840 3944
rect 844 3864 848 3944
rect 866 3864 870 3904
rect 931 3864 935 3904
rect 951 3864 955 3904
rect 1025 3864 1029 3904
rect 1097 3864 1101 3944
rect 1105 3864 1109 3944
rect 1151 3864 1155 3904
rect 1211 3864 1215 3944
rect 1219 3864 1223 3944
rect 1291 3864 1295 3904
rect 1377 3864 1381 3944
rect 1385 3864 1389 3944
rect 1445 3864 1449 3904
rect 1496 3864 1500 3944
rect 1504 3864 1508 3944
rect 1526 3864 1530 3904
rect 1591 3864 1595 3944
rect 1601 3864 1605 3944
rect 1631 3864 1635 3944
rect 1641 3864 1645 3944
rect 1711 3864 1715 3904
rect 1731 3864 1735 3904
rect 1805 3864 1809 3944
rect 1825 3864 1829 3944
rect 1845 3864 1849 3944
rect 1891 3864 1895 3904
rect 1911 3864 1915 3904
rect 1931 3864 1935 3904
rect 2010 3864 2014 3904
rect 2032 3864 2036 3944
rect 2040 3864 2044 3944
rect 2105 3864 2109 3904
rect 2165 3864 2169 3904
rect 2185 3864 2189 3904
rect 2205 3864 2209 3904
rect 2265 3864 2269 3904
rect 2285 3864 2289 3904
rect 2305 3864 2309 3904
rect 2365 3864 2369 3944
rect 2385 3864 2389 3944
rect 2405 3864 2409 3944
rect 2465 3864 2469 3904
rect 2530 3864 2534 3904
rect 2552 3864 2556 3944
rect 2560 3864 2564 3944
rect 2625 3864 2629 3904
rect 2645 3864 2649 3904
rect 2665 3864 2669 3904
rect 2725 3864 2729 3944
rect 2745 3864 2749 3944
rect 2765 3864 2769 3944
rect 2830 3864 2834 3904
rect 2852 3864 2856 3944
rect 2860 3864 2864 3944
rect 2916 3864 2920 3944
rect 2924 3864 2928 3944
rect 2946 3864 2950 3904
rect 3025 3864 3029 3904
rect 3045 3864 3049 3904
rect 3065 3864 3069 3904
rect 3125 3864 3129 3904
rect 3176 3864 3180 3944
rect 3184 3864 3188 3944
rect 3206 3864 3210 3904
rect 3271 3864 3275 3944
rect 3291 3864 3295 3944
rect 3311 3864 3315 3944
rect 3376 3864 3380 3944
rect 3384 3864 3388 3944
rect 3406 3864 3410 3904
rect 3490 3864 3494 3904
rect 3512 3864 3516 3944
rect 3520 3864 3524 3944
rect 3590 3864 3594 3904
rect 3612 3864 3616 3944
rect 3620 3864 3624 3944
rect 3685 3864 3689 3944
rect 3705 3864 3709 3944
rect 3725 3864 3729 3944
rect 3785 3864 3789 3904
rect 3805 3864 3809 3904
rect 3825 3864 3829 3904
rect 3885 3864 3889 3904
rect 3905 3864 3909 3904
rect 3965 3864 3969 3904
rect 3985 3864 3989 3904
rect 4031 3864 4035 3904
rect 4051 3864 4055 3904
rect 4125 3864 4129 3904
rect 4145 3864 4149 3904
rect 4165 3864 4169 3904
rect 4230 3864 4234 3904
rect 4252 3864 4256 3944
rect 4260 3864 4264 3944
rect 4316 3864 4320 3944
rect 4324 3864 4328 3944
rect 4346 3864 4350 3904
rect 4425 3864 4429 3904
rect 4485 3864 4489 3904
rect 4505 3864 4509 3904
rect 4525 3864 4529 3904
rect 4585 3864 4589 3904
rect 4605 3864 4609 3904
rect 4625 3864 4629 3904
rect 4671 3864 4675 3944
rect 4691 3864 4695 3944
rect 4711 3864 4715 3944
rect 50 3796 54 3836
rect 72 3756 76 3836
rect 80 3756 84 3836
rect 145 3796 149 3836
rect 191 3756 195 3836
rect 213 3816 217 3836
rect 221 3816 225 3836
rect 241 3796 245 3836
rect 249 3796 253 3836
rect 295 3796 299 3836
rect 315 3796 319 3836
rect 327 3796 331 3836
rect 347 3796 351 3836
rect 361 3796 365 3836
rect 381 3756 385 3836
rect 450 3796 454 3836
rect 472 3756 476 3836
rect 480 3756 484 3836
rect 531 3796 535 3836
rect 553 3796 557 3836
rect 575 3756 579 3836
rect 655 3756 659 3836
rect 675 3756 679 3836
rect 685 3756 689 3836
rect 745 3796 749 3836
rect 765 3796 769 3836
rect 815 3756 819 3836
rect 835 3796 839 3836
rect 849 3796 853 3836
rect 869 3796 873 3836
rect 881 3796 885 3836
rect 901 3796 905 3836
rect 947 3796 951 3836
rect 955 3796 959 3836
rect 975 3816 979 3836
rect 983 3816 987 3836
rect 1005 3756 1009 3836
rect 1063 3756 1067 3836
rect 1085 3796 1089 3836
rect 1131 3756 1135 3836
rect 1153 3816 1157 3836
rect 1161 3816 1165 3836
rect 1181 3796 1185 3836
rect 1189 3796 1193 3836
rect 1235 3796 1239 3836
rect 1255 3796 1259 3836
rect 1267 3796 1271 3836
rect 1287 3796 1291 3836
rect 1301 3796 1305 3836
rect 1321 3756 1325 3836
rect 1376 3756 1380 3836
rect 1384 3756 1388 3836
rect 1406 3796 1410 3836
rect 1471 3796 1475 3836
rect 1491 3796 1495 3836
rect 1551 3796 1555 3836
rect 1571 3796 1575 3836
rect 1631 3796 1635 3836
rect 1653 3756 1657 3836
rect 1711 3756 1715 3836
rect 1733 3816 1737 3836
rect 1741 3816 1745 3836
rect 1761 3796 1765 3836
rect 1769 3796 1773 3836
rect 1815 3796 1819 3836
rect 1835 3796 1839 3836
rect 1847 3796 1851 3836
rect 1867 3796 1871 3836
rect 1881 3796 1885 3836
rect 1901 3756 1905 3836
rect 1965 3796 1969 3836
rect 2025 3756 2029 3836
rect 2045 3756 2049 3836
rect 2065 3756 2069 3836
rect 2125 3796 2129 3836
rect 2171 3796 2175 3836
rect 2191 3796 2195 3836
rect 2211 3796 2215 3836
rect 2290 3796 2294 3836
rect 2312 3756 2316 3836
rect 2320 3756 2324 3836
rect 2385 3796 2389 3836
rect 2405 3796 2409 3836
rect 2425 3796 2429 3836
rect 2485 3756 2489 3836
rect 2505 3756 2509 3836
rect 2525 3756 2529 3836
rect 2585 3796 2589 3836
rect 2605 3796 2609 3836
rect 2625 3796 2629 3836
rect 2671 3756 2675 3836
rect 2691 3756 2695 3836
rect 2711 3756 2715 3836
rect 2785 3756 2789 3836
rect 2805 3756 2809 3836
rect 2825 3756 2829 3836
rect 2885 3796 2889 3836
rect 2945 3796 2949 3836
rect 3005 3796 3009 3836
rect 3025 3796 3029 3836
rect 3045 3796 3049 3836
rect 3105 3756 3109 3836
rect 3125 3756 3129 3836
rect 3145 3756 3149 3836
rect 3205 3796 3209 3836
rect 3225 3796 3229 3836
rect 3245 3796 3249 3836
rect 3305 3796 3309 3836
rect 3370 3796 3374 3836
rect 3392 3756 3396 3836
rect 3400 3756 3404 3836
rect 3465 3796 3469 3836
rect 3485 3796 3489 3836
rect 3531 3796 3535 3836
rect 3553 3796 3557 3836
rect 3575 3756 3579 3836
rect 3645 3756 3649 3836
rect 3665 3756 3669 3836
rect 3685 3756 3689 3836
rect 3745 3796 3749 3836
rect 3765 3796 3769 3836
rect 3785 3796 3789 3836
rect 3845 3796 3849 3836
rect 3891 3756 3895 3836
rect 3911 3756 3915 3836
rect 3931 3756 3935 3836
rect 4010 3796 4014 3836
rect 4032 3756 4036 3836
rect 4040 3756 4044 3836
rect 4096 3756 4100 3836
rect 4104 3756 4108 3836
rect 4126 3796 4130 3836
rect 4191 3756 4195 3836
rect 4211 3756 4215 3836
rect 4231 3756 4235 3836
rect 4305 3756 4309 3836
rect 4325 3756 4329 3836
rect 4345 3756 4349 3836
rect 4391 3796 4395 3836
rect 4411 3796 4415 3836
rect 4431 3796 4435 3836
rect 4505 3796 4509 3836
rect 4565 3796 4569 3836
rect 4585 3796 4589 3836
rect 4605 3796 4609 3836
rect 4651 3796 4655 3836
rect 4671 3796 4675 3836
rect 4691 3796 4695 3836
rect 35 3384 39 3464
rect 55 3384 59 3424
rect 69 3384 73 3424
rect 89 3384 93 3424
rect 101 3384 105 3424
rect 121 3384 125 3424
rect 167 3384 171 3424
rect 175 3384 179 3424
rect 195 3384 199 3404
rect 203 3384 207 3404
rect 225 3384 229 3464
rect 285 3384 289 3424
rect 305 3384 309 3424
rect 370 3384 374 3424
rect 392 3384 396 3464
rect 400 3384 404 3464
rect 465 3384 469 3424
rect 485 3384 489 3424
rect 545 3384 549 3424
rect 565 3384 569 3424
rect 585 3384 589 3424
rect 645 3384 649 3424
rect 710 3384 714 3424
rect 732 3384 736 3464
rect 740 3384 744 3464
rect 810 3384 814 3424
rect 832 3384 836 3464
rect 840 3384 844 3464
rect 891 3384 895 3424
rect 977 3384 981 3464
rect 985 3384 989 3464
rect 1031 3384 1035 3464
rect 1053 3384 1057 3404
rect 1061 3384 1065 3404
rect 1081 3384 1085 3424
rect 1089 3384 1093 3424
rect 1135 3384 1139 3424
rect 1155 3384 1159 3424
rect 1167 3384 1171 3424
rect 1187 3384 1191 3424
rect 1201 3384 1205 3424
rect 1221 3384 1225 3464
rect 1271 3384 1275 3424
rect 1331 3384 1335 3464
rect 1339 3384 1343 3464
rect 1416 3384 1420 3464
rect 1424 3384 1428 3464
rect 1446 3384 1450 3424
rect 1511 3384 1515 3424
rect 1531 3384 1535 3424
rect 1603 3384 1607 3464
rect 1625 3384 1629 3424
rect 1685 3384 1689 3424
rect 1731 3384 1735 3464
rect 1753 3384 1757 3404
rect 1761 3384 1765 3404
rect 1781 3384 1785 3424
rect 1789 3384 1793 3424
rect 1835 3384 1839 3424
rect 1855 3384 1859 3424
rect 1867 3384 1871 3424
rect 1887 3384 1891 3424
rect 1901 3384 1905 3424
rect 1921 3384 1925 3464
rect 1971 3384 1975 3464
rect 1981 3384 1985 3464
rect 2011 3384 2015 3464
rect 2021 3384 2025 3464
rect 2091 3384 2095 3424
rect 2111 3384 2115 3424
rect 2185 3384 2189 3464
rect 2205 3384 2209 3464
rect 2225 3384 2229 3464
rect 2285 3384 2289 3424
rect 2305 3384 2309 3424
rect 2325 3384 2329 3424
rect 2385 3384 2389 3424
rect 2445 3384 2449 3424
rect 2465 3384 2469 3424
rect 2485 3384 2489 3424
rect 2545 3384 2549 3424
rect 2565 3384 2569 3424
rect 2585 3384 2589 3424
rect 2650 3384 2654 3424
rect 2672 3384 2676 3464
rect 2680 3384 2684 3464
rect 2736 3384 2740 3464
rect 2744 3384 2748 3464
rect 2766 3384 2770 3424
rect 2831 3384 2835 3424
rect 2851 3384 2855 3424
rect 2916 3384 2920 3464
rect 2924 3384 2928 3464
rect 2946 3384 2950 3424
rect 3011 3384 3015 3464
rect 3019 3384 3023 3464
rect 3110 3384 3114 3424
rect 3132 3384 3136 3464
rect 3140 3384 3144 3464
rect 3191 3384 3195 3464
rect 3211 3384 3215 3464
rect 3231 3384 3235 3464
rect 3251 3384 3255 3464
rect 3311 3384 3315 3424
rect 3331 3384 3335 3424
rect 3391 3384 3395 3424
rect 3411 3384 3415 3424
rect 3471 3384 3475 3424
rect 3491 3384 3495 3424
rect 3551 3384 3555 3464
rect 3559 3384 3563 3464
rect 3631 3384 3635 3424
rect 3651 3384 3655 3424
rect 3711 3384 3715 3424
rect 3731 3384 3735 3424
rect 3805 3384 3809 3424
rect 3825 3384 3829 3424
rect 3897 3384 3901 3464
rect 3905 3384 3909 3464
rect 3951 3384 3955 3424
rect 3971 3384 3975 3424
rect 4031 3384 4035 3424
rect 4051 3384 4055 3424
rect 4116 3384 4120 3464
rect 4124 3384 4128 3464
rect 4146 3384 4150 3424
rect 4225 3384 4229 3424
rect 4245 3384 4249 3424
rect 4265 3384 4269 3424
rect 4311 3384 4315 3424
rect 4331 3384 4335 3424
rect 4351 3384 4355 3424
rect 4411 3384 4415 3464
rect 4431 3384 4435 3464
rect 4451 3384 4455 3464
rect 4511 3384 4515 3424
rect 4585 3384 4589 3424
rect 4605 3384 4609 3424
rect 4625 3384 4629 3424
rect 4671 3384 4675 3424
rect 4691 3384 4695 3424
rect 4711 3384 4715 3424
rect 35 3276 39 3356
rect 55 3316 59 3356
rect 69 3316 73 3356
rect 89 3316 93 3356
rect 101 3316 105 3356
rect 121 3316 125 3356
rect 167 3316 171 3356
rect 175 3316 179 3356
rect 195 3336 199 3356
rect 203 3336 207 3356
rect 225 3276 229 3356
rect 285 3276 289 3356
rect 305 3276 309 3356
rect 325 3276 329 3356
rect 345 3276 349 3356
rect 391 3316 395 3356
rect 411 3316 415 3356
rect 476 3276 480 3356
rect 484 3276 488 3356
rect 506 3316 510 3356
rect 576 3276 580 3356
rect 584 3276 588 3356
rect 606 3316 610 3356
rect 685 3316 689 3356
rect 705 3316 709 3356
rect 751 3316 755 3356
rect 825 3276 829 3356
rect 845 3276 849 3356
rect 865 3276 869 3356
rect 885 3276 889 3356
rect 905 3276 909 3356
rect 925 3276 929 3356
rect 945 3276 949 3356
rect 965 3276 969 3356
rect 1011 3276 1015 3356
rect 1031 3276 1035 3356
rect 1051 3276 1055 3356
rect 1071 3276 1075 3356
rect 1091 3276 1095 3356
rect 1111 3276 1115 3356
rect 1131 3276 1135 3356
rect 1151 3276 1155 3356
rect 1225 3316 1229 3356
rect 1271 3276 1275 3356
rect 1293 3336 1297 3356
rect 1301 3336 1305 3356
rect 1321 3316 1325 3356
rect 1329 3316 1333 3356
rect 1375 3316 1379 3356
rect 1395 3316 1399 3356
rect 1407 3316 1411 3356
rect 1427 3316 1431 3356
rect 1441 3316 1445 3356
rect 1461 3276 1465 3356
rect 1516 3276 1520 3356
rect 1524 3276 1528 3356
rect 1546 3316 1550 3356
rect 1630 3316 1634 3356
rect 1652 3276 1656 3356
rect 1660 3276 1664 3356
rect 1730 3316 1734 3356
rect 1752 3276 1756 3356
rect 1760 3276 1764 3356
rect 1825 3316 1829 3356
rect 1890 3316 1894 3356
rect 1912 3276 1916 3356
rect 1920 3276 1924 3356
rect 1990 3316 1994 3356
rect 2012 3276 2016 3356
rect 2020 3276 2024 3356
rect 2071 3276 2075 3356
rect 2093 3336 2097 3356
rect 2101 3336 2105 3356
rect 2121 3316 2125 3356
rect 2129 3316 2133 3356
rect 2175 3316 2179 3356
rect 2195 3316 2199 3356
rect 2207 3316 2211 3356
rect 2227 3316 2231 3356
rect 2241 3316 2245 3356
rect 2261 3276 2265 3356
rect 2325 3316 2329 3356
rect 2385 3316 2389 3356
rect 2445 3316 2449 3356
rect 2465 3316 2469 3356
rect 2485 3316 2489 3356
rect 2531 3276 2535 3356
rect 2551 3276 2555 3356
rect 2571 3276 2575 3356
rect 2645 3316 2649 3356
rect 2710 3316 2714 3356
rect 2732 3276 2736 3356
rect 2740 3276 2744 3356
rect 2791 3276 2795 3356
rect 2799 3276 2803 3356
rect 2876 3276 2880 3356
rect 2884 3276 2888 3356
rect 2906 3316 2910 3356
rect 2971 3316 2975 3356
rect 2991 3316 2995 3356
rect 3051 3316 3055 3356
rect 3071 3316 3075 3356
rect 3145 3276 3149 3356
rect 3165 3276 3169 3356
rect 3185 3276 3189 3356
rect 3245 3316 3249 3356
rect 3265 3316 3269 3356
rect 3285 3316 3289 3356
rect 3350 3316 3354 3356
rect 3372 3276 3376 3356
rect 3380 3276 3384 3356
rect 3441 3276 3445 3356
rect 3463 3316 3467 3356
rect 3485 3316 3489 3356
rect 3531 3316 3535 3356
rect 3551 3316 3555 3356
rect 3621 3276 3625 3356
rect 3643 3316 3647 3356
rect 3665 3316 3669 3356
rect 3725 3276 3729 3356
rect 3745 3276 3749 3356
rect 3765 3276 3769 3356
rect 3785 3276 3789 3356
rect 3845 3316 3849 3356
rect 3865 3316 3869 3356
rect 3916 3276 3920 3356
rect 3924 3276 3928 3356
rect 3946 3316 3950 3356
rect 4011 3316 4015 3356
rect 4031 3316 4035 3356
rect 4101 3276 4105 3356
rect 4123 3316 4127 3356
rect 4145 3316 4149 3356
rect 4191 3316 4195 3356
rect 4211 3316 4215 3356
rect 4271 3316 4275 3356
rect 4293 3316 4297 3356
rect 4315 3276 4319 3356
rect 4371 3276 4375 3356
rect 4391 3276 4395 3356
rect 4411 3276 4415 3356
rect 4476 3276 4480 3356
rect 4484 3276 4488 3356
rect 4506 3316 4510 3356
rect 4576 3276 4580 3356
rect 4584 3276 4588 3356
rect 4606 3316 4610 3356
rect 4685 3316 4689 3356
rect 4705 3316 4709 3356
rect 4725 3316 4729 3356
rect 35 2904 39 2984
rect 55 2904 59 2944
rect 69 2904 73 2944
rect 89 2904 93 2944
rect 101 2904 105 2944
rect 121 2904 125 2944
rect 167 2904 171 2944
rect 175 2904 179 2944
rect 195 2904 199 2924
rect 203 2904 207 2924
rect 225 2904 229 2984
rect 290 2904 294 2944
rect 312 2904 316 2984
rect 320 2904 324 2984
rect 385 2904 389 2944
rect 405 2904 409 2944
rect 451 2904 455 2984
rect 473 2904 477 2924
rect 481 2904 485 2924
rect 501 2904 505 2944
rect 509 2904 513 2944
rect 555 2904 559 2944
rect 575 2904 579 2944
rect 587 2904 591 2944
rect 607 2904 611 2944
rect 621 2904 625 2944
rect 641 2904 645 2984
rect 695 2904 699 2984
rect 715 2904 719 2944
rect 729 2904 733 2944
rect 749 2904 753 2944
rect 761 2904 765 2944
rect 781 2904 785 2944
rect 827 2904 831 2944
rect 835 2904 839 2944
rect 855 2904 859 2924
rect 863 2904 867 2924
rect 885 2904 889 2984
rect 931 2904 935 2944
rect 1017 2904 1021 2984
rect 1025 2904 1029 2984
rect 1085 2904 1089 2944
rect 1105 2904 1109 2944
rect 1156 2904 1160 2984
rect 1164 2904 1168 2984
rect 1186 2904 1190 2944
rect 1251 2904 1255 2984
rect 1271 2904 1275 2984
rect 1291 2904 1295 2984
rect 1355 2904 1359 2984
rect 1375 2904 1379 2944
rect 1389 2904 1393 2944
rect 1409 2904 1413 2944
rect 1421 2904 1425 2944
rect 1441 2904 1445 2944
rect 1487 2904 1491 2944
rect 1495 2904 1499 2944
rect 1515 2904 1519 2924
rect 1523 2904 1527 2924
rect 1545 2904 1549 2984
rect 1617 2904 1621 2984
rect 1625 2904 1629 2984
rect 1685 2904 1689 2944
rect 1705 2904 1709 2944
rect 1756 2904 1760 2984
rect 1764 2904 1768 2984
rect 1786 2904 1790 2944
rect 1870 2904 1874 2944
rect 1892 2904 1896 2984
rect 1900 2904 1904 2984
rect 1951 2904 1955 2984
rect 1973 2904 1977 2924
rect 1981 2904 1985 2924
rect 2001 2904 2005 2944
rect 2009 2904 2013 2944
rect 2055 2904 2059 2944
rect 2075 2904 2079 2944
rect 2087 2904 2091 2944
rect 2107 2904 2111 2944
rect 2121 2904 2125 2944
rect 2141 2904 2145 2984
rect 2217 2904 2221 2984
rect 2225 2904 2229 2984
rect 2285 2904 2289 2944
rect 2345 2904 2349 2944
rect 2365 2904 2369 2944
rect 2385 2904 2389 2944
rect 2445 2904 2449 2984
rect 2465 2904 2469 2984
rect 2485 2904 2489 2984
rect 2545 2904 2549 2944
rect 2565 2904 2569 2944
rect 2585 2904 2589 2944
rect 2650 2904 2654 2944
rect 2672 2904 2676 2984
rect 2680 2904 2684 2984
rect 2757 2904 2761 2984
rect 2765 2904 2769 2984
rect 2811 2904 2815 2944
rect 2831 2904 2835 2944
rect 2891 2904 2895 2944
rect 2911 2904 2915 2944
rect 2971 2904 2975 2984
rect 2991 2904 2995 2984
rect 3011 2904 3015 2984
rect 3031 2904 3035 2984
rect 3091 2904 3095 2944
rect 3111 2904 3115 2944
rect 3176 2904 3180 2984
rect 3184 2904 3188 2984
rect 3206 2904 3210 2944
rect 3271 2904 3275 2984
rect 3331 2904 3335 2944
rect 3353 2904 3357 2944
rect 3375 2904 3379 2984
rect 3443 2904 3447 2984
rect 3465 2904 3469 2944
rect 3523 2904 3527 2984
rect 3545 2904 3549 2944
rect 3591 2904 3595 2944
rect 3611 2904 3615 2944
rect 3676 2904 3680 2984
rect 3684 2904 3688 2984
rect 3706 2904 3710 2944
rect 3783 2904 3787 2984
rect 3805 2904 3809 2944
rect 3856 2904 3860 2984
rect 3864 2904 3868 2984
rect 3886 2904 3890 2944
rect 3951 2904 3955 2944
rect 3971 2904 3975 2944
rect 3991 2904 3995 2944
rect 4051 2904 4055 2944
rect 4073 2904 4077 2984
rect 4145 2904 4149 2984
rect 4165 2904 4169 2984
rect 4185 2904 4189 2984
rect 4231 2904 4235 2944
rect 4251 2904 4255 2944
rect 4271 2904 4275 2944
rect 4345 2904 4349 2984
rect 4365 2904 4369 2984
rect 4385 2904 4389 2984
rect 4445 2904 4449 2944
rect 4465 2904 4469 2944
rect 4485 2904 4489 2944
rect 4545 2904 4549 2944
rect 4610 2904 4614 2944
rect 4632 2904 4636 2984
rect 4640 2904 4644 2984
rect 4696 2904 4700 2984
rect 4704 2904 4708 2984
rect 4726 2904 4730 2944
rect 35 2796 39 2876
rect 55 2836 59 2876
rect 69 2836 73 2876
rect 89 2836 93 2876
rect 101 2836 105 2876
rect 121 2836 125 2876
rect 167 2836 171 2876
rect 175 2836 179 2876
rect 195 2856 199 2876
rect 203 2856 207 2876
rect 225 2796 229 2876
rect 285 2796 289 2876
rect 305 2796 309 2876
rect 325 2796 329 2876
rect 345 2796 349 2876
rect 391 2836 395 2876
rect 411 2836 415 2876
rect 490 2836 494 2876
rect 512 2796 516 2876
rect 520 2796 524 2876
rect 583 2796 587 2876
rect 605 2836 609 2876
rect 651 2836 655 2876
rect 671 2836 675 2876
rect 750 2836 754 2876
rect 772 2796 776 2876
rect 780 2796 784 2876
rect 857 2796 861 2876
rect 865 2796 869 2876
rect 925 2836 929 2876
rect 945 2836 949 2876
rect 991 2836 995 2876
rect 1065 2836 1069 2876
rect 1085 2836 1089 2876
rect 1131 2796 1135 2876
rect 1139 2796 1143 2876
rect 1223 2796 1227 2876
rect 1245 2836 1249 2876
rect 1295 2796 1299 2876
rect 1315 2836 1319 2876
rect 1329 2836 1333 2876
rect 1349 2836 1353 2876
rect 1361 2836 1365 2876
rect 1381 2836 1385 2876
rect 1427 2836 1431 2876
rect 1435 2836 1439 2876
rect 1455 2856 1459 2876
rect 1463 2856 1467 2876
rect 1485 2796 1489 2876
rect 1531 2836 1535 2876
rect 1551 2836 1555 2876
rect 1630 2836 1634 2876
rect 1652 2796 1656 2876
rect 1660 2796 1664 2876
rect 1730 2836 1734 2876
rect 1752 2796 1756 2876
rect 1760 2796 1764 2876
rect 1837 2796 1841 2876
rect 1845 2796 1849 2876
rect 1905 2796 1909 2876
rect 1925 2796 1929 2876
rect 1945 2796 1949 2876
rect 2003 2796 2007 2876
rect 2025 2836 2029 2876
rect 2085 2836 2089 2876
rect 2105 2836 2109 2876
rect 2125 2836 2129 2876
rect 2171 2836 2175 2876
rect 2193 2796 2197 2876
rect 2255 2796 2259 2876
rect 2275 2836 2279 2876
rect 2289 2836 2293 2876
rect 2309 2836 2313 2876
rect 2321 2836 2325 2876
rect 2341 2836 2345 2876
rect 2387 2836 2391 2876
rect 2395 2836 2399 2876
rect 2415 2856 2419 2876
rect 2423 2856 2427 2876
rect 2445 2796 2449 2876
rect 2510 2836 2514 2876
rect 2532 2796 2536 2876
rect 2540 2796 2544 2876
rect 2610 2836 2614 2876
rect 2632 2796 2636 2876
rect 2640 2796 2644 2876
rect 2696 2796 2700 2876
rect 2704 2796 2708 2876
rect 2726 2836 2730 2876
rect 2791 2836 2795 2876
rect 2811 2836 2815 2876
rect 2871 2836 2875 2876
rect 2891 2836 2895 2876
rect 2956 2796 2960 2876
rect 2964 2796 2968 2876
rect 2986 2836 2990 2876
rect 3056 2796 3060 2876
rect 3064 2796 3068 2876
rect 3086 2836 3090 2876
rect 3151 2836 3155 2876
rect 3171 2836 3175 2876
rect 3250 2836 3254 2876
rect 3272 2796 3276 2876
rect 3280 2796 3284 2876
rect 3345 2836 3349 2876
rect 3365 2836 3369 2876
rect 3411 2836 3415 2876
rect 3431 2836 3435 2876
rect 3451 2836 3455 2876
rect 3530 2836 3534 2876
rect 3552 2796 3556 2876
rect 3560 2796 3564 2876
rect 3616 2796 3620 2876
rect 3624 2796 3628 2876
rect 3646 2836 3650 2876
rect 3725 2836 3729 2876
rect 3745 2836 3749 2876
rect 3810 2836 3814 2876
rect 3832 2796 3836 2876
rect 3840 2796 3844 2876
rect 3891 2836 3895 2876
rect 3911 2836 3915 2876
rect 3931 2836 3935 2876
rect 3991 2836 3995 2876
rect 4065 2796 4069 2876
rect 4085 2796 4089 2876
rect 4105 2796 4109 2876
rect 4125 2796 4129 2876
rect 4171 2836 4175 2876
rect 4191 2836 4195 2876
rect 4211 2836 4215 2876
rect 4276 2796 4280 2876
rect 4284 2796 4288 2876
rect 4306 2836 4310 2876
rect 4371 2836 4375 2876
rect 4393 2836 4397 2876
rect 4415 2796 4419 2876
rect 4471 2796 4475 2876
rect 4491 2796 4495 2876
rect 4511 2796 4515 2876
rect 4531 2796 4535 2876
rect 4591 2836 4595 2876
rect 4651 2796 4655 2876
rect 4671 2796 4675 2876
rect 4691 2796 4695 2876
rect 35 2424 39 2504
rect 55 2424 59 2464
rect 69 2424 73 2464
rect 89 2424 93 2464
rect 101 2424 105 2464
rect 121 2424 125 2464
rect 167 2424 171 2464
rect 175 2424 179 2464
rect 195 2424 199 2444
rect 203 2424 207 2444
rect 225 2424 229 2504
rect 290 2424 294 2464
rect 312 2424 316 2504
rect 320 2424 324 2504
rect 371 2424 375 2464
rect 393 2424 397 2504
rect 451 2424 455 2464
rect 471 2424 475 2464
rect 550 2424 554 2464
rect 572 2424 576 2504
rect 580 2424 584 2504
rect 631 2424 635 2464
rect 653 2424 657 2504
rect 730 2424 734 2464
rect 752 2424 756 2504
rect 760 2424 764 2504
rect 811 2424 815 2504
rect 819 2424 823 2504
rect 895 2424 899 2504
rect 915 2424 919 2464
rect 929 2424 933 2464
rect 949 2424 953 2464
rect 961 2424 965 2464
rect 981 2424 985 2464
rect 1027 2424 1031 2464
rect 1035 2424 1039 2464
rect 1055 2424 1059 2444
rect 1063 2424 1067 2444
rect 1085 2424 1089 2504
rect 1131 2424 1135 2464
rect 1196 2424 1200 2504
rect 1204 2424 1208 2504
rect 1226 2424 1230 2464
rect 1291 2424 1295 2464
rect 1351 2424 1355 2464
rect 1371 2424 1375 2464
rect 1431 2424 1435 2504
rect 1453 2424 1457 2444
rect 1461 2424 1465 2444
rect 1481 2424 1485 2464
rect 1489 2424 1493 2464
rect 1535 2424 1539 2464
rect 1555 2424 1559 2464
rect 1567 2424 1571 2464
rect 1587 2424 1591 2464
rect 1601 2424 1605 2464
rect 1621 2424 1625 2504
rect 1676 2424 1680 2504
rect 1684 2424 1688 2504
rect 1706 2424 1710 2464
rect 1771 2424 1775 2504
rect 1793 2424 1797 2444
rect 1801 2424 1805 2444
rect 1821 2424 1825 2464
rect 1829 2424 1833 2464
rect 1875 2424 1879 2464
rect 1895 2424 1899 2464
rect 1907 2424 1911 2464
rect 1927 2424 1931 2464
rect 1941 2424 1945 2464
rect 1961 2424 1965 2504
rect 2011 2424 2015 2504
rect 2031 2424 2035 2504
rect 2051 2424 2055 2504
rect 2071 2424 2075 2504
rect 2091 2424 2095 2504
rect 2111 2424 2115 2504
rect 2131 2424 2135 2504
rect 2151 2424 2155 2504
rect 2215 2424 2219 2504
rect 2235 2424 2239 2464
rect 2249 2424 2253 2464
rect 2269 2424 2273 2464
rect 2281 2424 2285 2464
rect 2301 2424 2305 2464
rect 2347 2424 2351 2464
rect 2355 2424 2359 2464
rect 2375 2424 2379 2444
rect 2383 2424 2387 2444
rect 2405 2424 2409 2504
rect 2465 2424 2469 2464
rect 2485 2424 2489 2464
rect 2531 2424 2535 2464
rect 2610 2424 2614 2464
rect 2632 2424 2636 2504
rect 2640 2424 2644 2504
rect 2691 2424 2695 2464
rect 2765 2424 2769 2464
rect 2785 2424 2789 2464
rect 2850 2424 2854 2464
rect 2872 2424 2876 2504
rect 2880 2424 2884 2504
rect 2931 2424 2935 2464
rect 2953 2424 2957 2464
rect 2975 2424 2979 2504
rect 3036 2424 3040 2504
rect 3044 2424 3048 2504
rect 3066 2424 3070 2464
rect 3145 2424 3149 2464
rect 3165 2424 3169 2464
rect 3211 2424 3215 2464
rect 3233 2424 3237 2464
rect 3255 2424 3259 2504
rect 3325 2424 3329 2464
rect 3345 2424 3349 2464
rect 3365 2424 3369 2464
rect 3411 2424 3415 2464
rect 3471 2424 3475 2464
rect 3491 2424 3495 2464
rect 3551 2424 3555 2464
rect 3573 2424 3577 2464
rect 3595 2424 3599 2504
rect 3651 2424 3655 2464
rect 3673 2424 3677 2504
rect 3731 2424 3735 2464
rect 3801 2424 3805 2504
rect 3823 2424 3827 2464
rect 3845 2424 3849 2464
rect 3905 2424 3909 2504
rect 3925 2424 3929 2504
rect 3945 2424 3949 2504
rect 3965 2424 3969 2504
rect 4025 2424 4029 2464
rect 4045 2424 4049 2464
rect 4105 2424 4109 2464
rect 4125 2424 4129 2464
rect 4176 2424 4180 2504
rect 4184 2424 4188 2504
rect 4206 2424 4210 2464
rect 4271 2424 4275 2464
rect 4291 2424 4295 2464
rect 4365 2424 4369 2464
rect 4385 2424 4389 2464
rect 4405 2424 4409 2464
rect 4465 2424 4469 2464
rect 4485 2424 4489 2464
rect 4505 2424 4509 2464
rect 4551 2424 4555 2504
rect 4571 2424 4575 2504
rect 4591 2424 4595 2504
rect 4665 2424 4669 2464
rect 4685 2424 4689 2464
rect 4705 2424 4709 2464
rect 35 2316 39 2396
rect 55 2356 59 2396
rect 69 2356 73 2396
rect 89 2356 93 2396
rect 101 2356 105 2396
rect 121 2356 125 2396
rect 167 2356 171 2396
rect 175 2356 179 2396
rect 195 2376 199 2396
rect 203 2376 207 2396
rect 225 2316 229 2396
rect 276 2316 280 2396
rect 284 2316 288 2396
rect 306 2356 310 2396
rect 371 2316 375 2396
rect 391 2316 395 2396
rect 411 2316 415 2396
rect 431 2316 435 2396
rect 491 2356 495 2396
rect 513 2316 517 2396
rect 571 2356 575 2396
rect 591 2356 595 2396
rect 665 2356 669 2396
rect 711 2316 715 2396
rect 719 2316 723 2396
rect 805 2316 809 2396
rect 825 2316 829 2396
rect 845 2316 849 2396
rect 891 2316 895 2396
rect 899 2316 903 2396
rect 971 2316 975 2396
rect 979 2316 983 2396
rect 1051 2356 1055 2396
rect 1111 2316 1115 2396
rect 1133 2376 1137 2396
rect 1141 2376 1145 2396
rect 1161 2356 1165 2396
rect 1169 2356 1173 2396
rect 1215 2356 1219 2396
rect 1235 2356 1239 2396
rect 1247 2356 1251 2396
rect 1267 2356 1271 2396
rect 1281 2356 1285 2396
rect 1301 2316 1305 2396
rect 1356 2316 1360 2396
rect 1364 2316 1368 2396
rect 1386 2356 1390 2396
rect 1451 2316 1455 2396
rect 1473 2376 1477 2396
rect 1481 2376 1485 2396
rect 1501 2356 1505 2396
rect 1509 2356 1513 2396
rect 1555 2356 1559 2396
rect 1575 2356 1579 2396
rect 1587 2356 1591 2396
rect 1607 2356 1611 2396
rect 1621 2356 1625 2396
rect 1641 2316 1645 2396
rect 1717 2316 1721 2396
rect 1725 2316 1729 2396
rect 1785 2316 1789 2396
rect 1805 2316 1809 2396
rect 1825 2316 1829 2396
rect 1871 2316 1875 2396
rect 1957 2316 1961 2396
rect 1965 2316 1969 2396
rect 2011 2316 2015 2396
rect 2031 2316 2035 2396
rect 2051 2316 2055 2396
rect 2071 2316 2075 2396
rect 2091 2316 2095 2396
rect 2111 2316 2115 2396
rect 2131 2316 2135 2396
rect 2151 2316 2155 2396
rect 2216 2316 2220 2396
rect 2224 2316 2228 2396
rect 2246 2356 2250 2396
rect 2315 2316 2319 2396
rect 2335 2356 2339 2396
rect 2349 2356 2353 2396
rect 2369 2356 2373 2396
rect 2381 2356 2385 2396
rect 2401 2356 2405 2396
rect 2447 2356 2451 2396
rect 2455 2356 2459 2396
rect 2475 2376 2479 2396
rect 2483 2376 2487 2396
rect 2505 2316 2509 2396
rect 2565 2356 2569 2396
rect 2585 2356 2589 2396
rect 2631 2356 2635 2396
rect 2651 2356 2655 2396
rect 2711 2356 2715 2396
rect 2731 2356 2735 2396
rect 2810 2356 2814 2396
rect 2832 2316 2836 2396
rect 2840 2316 2844 2396
rect 2910 2356 2914 2396
rect 2932 2316 2936 2396
rect 2940 2316 2944 2396
rect 2995 2316 2999 2396
rect 3015 2356 3019 2396
rect 3029 2356 3033 2396
rect 3049 2356 3053 2396
rect 3061 2356 3065 2396
rect 3081 2356 3085 2396
rect 3127 2356 3131 2396
rect 3135 2356 3139 2396
rect 3155 2376 3159 2396
rect 3163 2376 3167 2396
rect 3185 2316 3189 2396
rect 3236 2316 3240 2396
rect 3244 2316 3248 2396
rect 3266 2356 3270 2396
rect 3331 2356 3335 2396
rect 3351 2356 3355 2396
rect 3411 2356 3415 2396
rect 3431 2356 3435 2396
rect 3505 2356 3509 2396
rect 3525 2356 3529 2396
rect 3585 2316 3589 2396
rect 3645 2316 3649 2396
rect 3705 2356 3709 2396
rect 3756 2316 3760 2396
rect 3764 2316 3768 2396
rect 3786 2356 3790 2396
rect 3863 2316 3867 2396
rect 3885 2356 3889 2396
rect 3931 2316 3935 2396
rect 3991 2356 3995 2396
rect 4013 2356 4017 2396
rect 4035 2316 4039 2396
rect 4110 2356 4114 2396
rect 4132 2316 4136 2396
rect 4140 2316 4144 2396
rect 4205 2356 4209 2396
rect 4225 2356 4229 2396
rect 4245 2356 4249 2396
rect 4291 2316 4295 2396
rect 4311 2316 4315 2396
rect 4331 2316 4335 2396
rect 4410 2356 4414 2396
rect 4432 2316 4436 2396
rect 4440 2316 4444 2396
rect 4496 2316 4500 2396
rect 4504 2316 4508 2396
rect 4526 2356 4530 2396
rect 4610 2356 4614 2396
rect 4632 2316 4636 2396
rect 4640 2316 4644 2396
rect 4691 2316 4695 2396
rect 4711 2316 4715 2396
rect 4731 2316 4735 2396
rect 31 1944 35 2024
rect 51 1944 55 2024
rect 71 1944 75 2024
rect 91 1944 95 2024
rect 111 1944 115 2024
rect 131 1944 135 2024
rect 151 1944 155 2024
rect 171 1944 175 2024
rect 245 1944 249 1984
rect 265 1944 269 1984
rect 330 1944 334 1984
rect 352 1944 356 2024
rect 360 1944 364 2024
rect 411 1944 415 2024
rect 431 1944 435 2024
rect 451 1944 455 2024
rect 471 1944 475 2024
rect 535 1944 539 2024
rect 555 1944 559 1984
rect 569 1944 573 1984
rect 589 1944 593 1984
rect 601 1944 605 1984
rect 621 1944 625 1984
rect 667 1944 671 1984
rect 675 1944 679 1984
rect 695 1944 699 1964
rect 703 1944 707 1964
rect 725 1944 729 2024
rect 785 1944 789 1984
rect 805 1944 809 1984
rect 875 1944 879 2024
rect 895 1944 899 2024
rect 905 1944 909 2024
rect 951 1944 955 1984
rect 971 1944 975 1984
rect 1031 1944 1035 2024
rect 1039 1944 1043 2024
rect 1116 1944 1120 2024
rect 1124 1944 1128 2024
rect 1146 1944 1150 1984
rect 1211 1944 1215 1984
rect 1231 1944 1235 1984
rect 1291 1944 1295 2024
rect 1299 1944 1303 2024
rect 1371 1944 1375 2024
rect 1393 1944 1397 1964
rect 1401 1944 1405 1964
rect 1421 1944 1425 1984
rect 1429 1944 1433 1984
rect 1475 1944 1479 1984
rect 1495 1944 1499 1984
rect 1507 1944 1511 1984
rect 1527 1944 1531 1984
rect 1541 1944 1545 1984
rect 1561 1944 1565 2024
rect 1625 1944 1629 2024
rect 1645 1944 1649 2024
rect 1665 1944 1669 2024
rect 1723 1944 1727 2024
rect 1745 1944 1749 1984
rect 1791 1944 1795 2024
rect 1813 1944 1817 1964
rect 1821 1944 1825 1964
rect 1841 1944 1845 1984
rect 1849 1944 1853 1984
rect 1895 1944 1899 1984
rect 1915 1944 1919 1984
rect 1927 1944 1931 1984
rect 1947 1944 1951 1984
rect 1961 1944 1965 1984
rect 1981 1944 1985 2024
rect 2045 1944 2049 1984
rect 2105 1944 2109 1984
rect 2125 1944 2129 1984
rect 2171 1944 2175 1984
rect 2193 1944 2197 2024
rect 2251 1944 2255 1984
rect 2271 1944 2275 1984
rect 2350 1944 2354 1984
rect 2372 1944 2376 2024
rect 2380 1944 2384 2024
rect 2445 1944 2449 1984
rect 2465 1944 2469 1984
rect 2525 1944 2529 1984
rect 2545 1944 2549 1984
rect 2610 1944 2614 1984
rect 2632 1944 2636 2024
rect 2640 1944 2644 2024
rect 2710 1944 2714 1984
rect 2732 1944 2736 2024
rect 2740 1944 2744 2024
rect 2795 1944 2799 2024
rect 2815 1944 2819 1984
rect 2829 1944 2833 1984
rect 2849 1944 2853 1984
rect 2861 1944 2865 1984
rect 2881 1944 2885 1984
rect 2927 1944 2931 1984
rect 2935 1944 2939 1984
rect 2955 1944 2959 1964
rect 2963 1944 2967 1964
rect 2985 1944 2989 2024
rect 3031 1944 3035 1984
rect 3053 1944 3057 1984
rect 3075 1944 3079 2024
rect 3150 1944 3154 1984
rect 3172 1944 3176 2024
rect 3180 1944 3184 2024
rect 3250 1944 3254 1984
rect 3272 1944 3276 2024
rect 3280 1944 3284 2024
rect 3331 1944 3335 1984
rect 3351 1944 3355 1984
rect 3430 1944 3434 1984
rect 3452 1944 3456 2024
rect 3460 1944 3464 2024
rect 3511 1944 3515 1984
rect 3531 1944 3535 1984
rect 3551 1944 3555 1984
rect 3611 1944 3615 1984
rect 3671 1944 3675 1984
rect 3691 1944 3695 1984
rect 3711 1944 3715 1984
rect 3771 1944 3775 1984
rect 3791 1944 3795 1984
rect 3851 1944 3855 1984
rect 3873 1944 3877 2024
rect 3936 1944 3940 2024
rect 3944 1944 3948 2024
rect 3966 1944 3970 1984
rect 4045 1944 4049 1984
rect 4065 1944 4069 1984
rect 4125 1944 4129 1984
rect 4145 1944 4149 1984
rect 4205 1944 4209 1984
rect 4225 1944 4229 1984
rect 4271 1944 4275 1984
rect 4293 1944 4297 1984
rect 4315 1944 4319 2024
rect 4371 1944 4375 2024
rect 4391 1944 4395 2024
rect 4411 1944 4415 2024
rect 4485 1944 4489 2024
rect 4505 1944 4509 2024
rect 4525 1944 4529 2024
rect 4571 1944 4575 1984
rect 4591 1944 4595 1984
rect 4611 1944 4615 1984
rect 4671 1944 4675 1984
rect 4691 1944 4695 1984
rect 4711 1944 4715 1984
rect 35 1836 39 1916
rect 55 1876 59 1916
rect 69 1876 73 1916
rect 89 1876 93 1916
rect 101 1876 105 1916
rect 121 1876 125 1916
rect 167 1876 171 1916
rect 175 1876 179 1916
rect 195 1896 199 1916
rect 203 1896 207 1916
rect 225 1836 229 1916
rect 276 1836 280 1916
rect 284 1836 288 1916
rect 306 1876 310 1916
rect 390 1876 394 1916
rect 412 1836 416 1916
rect 420 1836 424 1916
rect 490 1876 494 1916
rect 512 1836 516 1916
rect 520 1836 524 1916
rect 590 1876 594 1916
rect 612 1836 616 1916
rect 620 1836 624 1916
rect 671 1876 675 1916
rect 731 1876 735 1916
rect 817 1836 821 1916
rect 825 1836 829 1916
rect 871 1876 875 1916
rect 891 1876 895 1916
rect 911 1876 915 1916
rect 975 1836 979 1916
rect 995 1876 999 1916
rect 1009 1876 1013 1916
rect 1029 1876 1033 1916
rect 1041 1876 1045 1916
rect 1061 1876 1065 1916
rect 1107 1876 1111 1916
rect 1115 1876 1119 1916
rect 1135 1896 1139 1916
rect 1143 1896 1147 1916
rect 1165 1836 1169 1916
rect 1211 1876 1215 1916
rect 1231 1876 1235 1916
rect 1310 1876 1314 1916
rect 1332 1836 1336 1916
rect 1340 1836 1344 1916
rect 1405 1836 1409 1916
rect 1425 1836 1429 1916
rect 1445 1836 1449 1916
rect 1465 1836 1469 1916
rect 1485 1836 1489 1916
rect 1505 1836 1509 1916
rect 1525 1836 1529 1916
rect 1545 1836 1549 1916
rect 1595 1836 1599 1916
rect 1615 1876 1619 1916
rect 1629 1876 1633 1916
rect 1649 1876 1653 1916
rect 1661 1876 1665 1916
rect 1681 1876 1685 1916
rect 1727 1876 1731 1916
rect 1735 1876 1739 1916
rect 1755 1896 1759 1916
rect 1763 1896 1767 1916
rect 1785 1836 1789 1916
rect 1845 1836 1849 1916
rect 1865 1836 1869 1916
rect 1885 1836 1889 1916
rect 1931 1836 1935 1916
rect 1939 1836 1943 1916
rect 2025 1836 2029 1916
rect 2045 1836 2049 1916
rect 2065 1836 2069 1916
rect 2137 1836 2141 1916
rect 2145 1836 2149 1916
rect 2191 1836 2195 1916
rect 2211 1836 2215 1916
rect 2231 1836 2235 1916
rect 2291 1836 2295 1916
rect 2313 1896 2317 1916
rect 2321 1896 2325 1916
rect 2341 1876 2345 1916
rect 2349 1876 2353 1916
rect 2395 1876 2399 1916
rect 2415 1876 2419 1916
rect 2427 1876 2431 1916
rect 2447 1876 2451 1916
rect 2461 1876 2465 1916
rect 2481 1836 2485 1916
rect 2535 1836 2539 1916
rect 2555 1876 2559 1916
rect 2569 1876 2573 1916
rect 2589 1876 2593 1916
rect 2601 1876 2605 1916
rect 2621 1876 2625 1916
rect 2667 1876 2671 1916
rect 2675 1876 2679 1916
rect 2695 1896 2699 1916
rect 2703 1896 2707 1916
rect 2725 1836 2729 1916
rect 2775 1836 2779 1916
rect 2795 1876 2799 1916
rect 2809 1876 2813 1916
rect 2829 1876 2833 1916
rect 2841 1876 2845 1916
rect 2861 1876 2865 1916
rect 2907 1876 2911 1916
rect 2915 1876 2919 1916
rect 2935 1896 2939 1916
rect 2943 1896 2947 1916
rect 2965 1836 2969 1916
rect 3025 1836 3029 1916
rect 3085 1876 3089 1916
rect 3105 1876 3109 1916
rect 3165 1836 3169 1916
rect 3211 1836 3215 1916
rect 3231 1836 3235 1916
rect 3251 1836 3255 1916
rect 3311 1836 3315 1916
rect 3319 1836 3323 1916
rect 3401 1836 3405 1916
rect 3423 1876 3427 1916
rect 3445 1876 3449 1916
rect 3491 1836 3495 1916
rect 3565 1836 3569 1916
rect 3585 1836 3589 1916
rect 3605 1836 3609 1916
rect 3625 1836 3629 1916
rect 3685 1836 3689 1916
rect 3757 1836 3761 1916
rect 3765 1836 3769 1916
rect 3811 1876 3815 1916
rect 3833 1836 3837 1916
rect 3891 1876 3895 1916
rect 3913 1876 3917 1916
rect 3935 1836 3939 1916
rect 4005 1836 4009 1916
rect 4025 1836 4029 1916
rect 4045 1836 4049 1916
rect 4065 1836 4069 1916
rect 4111 1836 4115 1916
rect 4131 1836 4135 1916
rect 4151 1836 4155 1916
rect 4171 1836 4175 1916
rect 4231 1876 4235 1916
rect 4251 1876 4255 1916
rect 4311 1876 4315 1916
rect 4333 1876 4337 1916
rect 4355 1836 4359 1916
rect 4411 1836 4415 1916
rect 4431 1836 4435 1916
rect 4451 1836 4455 1916
rect 4471 1836 4475 1916
rect 4545 1876 4549 1916
rect 4596 1836 4600 1916
rect 4604 1836 4608 1916
rect 4626 1876 4630 1916
rect 4691 1876 4695 1916
rect 31 1464 35 1544
rect 51 1464 55 1544
rect 71 1464 75 1544
rect 91 1464 95 1544
rect 111 1464 115 1544
rect 131 1464 135 1544
rect 151 1464 155 1544
rect 171 1464 175 1544
rect 257 1464 261 1544
rect 265 1464 269 1544
rect 323 1464 327 1544
rect 345 1464 349 1504
rect 395 1464 399 1544
rect 415 1464 419 1504
rect 429 1464 433 1504
rect 449 1464 453 1504
rect 461 1464 465 1504
rect 481 1464 485 1504
rect 527 1464 531 1504
rect 535 1464 539 1504
rect 555 1464 559 1484
rect 563 1464 567 1484
rect 585 1464 589 1544
rect 635 1464 639 1544
rect 655 1464 659 1504
rect 669 1464 673 1504
rect 689 1464 693 1504
rect 701 1464 705 1504
rect 721 1464 725 1504
rect 767 1464 771 1504
rect 775 1464 779 1504
rect 795 1464 799 1484
rect 803 1464 807 1484
rect 825 1464 829 1544
rect 871 1464 875 1544
rect 893 1464 897 1484
rect 901 1464 905 1484
rect 921 1464 925 1504
rect 929 1464 933 1504
rect 975 1464 979 1504
rect 995 1464 999 1504
rect 1007 1464 1011 1504
rect 1027 1464 1031 1504
rect 1041 1464 1045 1504
rect 1061 1464 1065 1544
rect 1125 1464 1129 1504
rect 1145 1464 1149 1504
rect 1210 1464 1214 1504
rect 1232 1464 1236 1544
rect 1240 1464 1244 1544
rect 1291 1464 1295 1544
rect 1313 1464 1317 1484
rect 1321 1464 1325 1484
rect 1341 1464 1345 1504
rect 1349 1464 1353 1504
rect 1395 1464 1399 1504
rect 1415 1464 1419 1504
rect 1427 1464 1431 1504
rect 1447 1464 1451 1504
rect 1461 1464 1465 1504
rect 1481 1464 1485 1544
rect 1535 1464 1539 1544
rect 1555 1464 1559 1504
rect 1569 1464 1573 1504
rect 1589 1464 1593 1504
rect 1601 1464 1605 1504
rect 1621 1464 1625 1504
rect 1667 1464 1671 1504
rect 1675 1464 1679 1504
rect 1695 1464 1699 1484
rect 1703 1464 1707 1484
rect 1725 1464 1729 1544
rect 1785 1464 1789 1544
rect 1805 1464 1809 1544
rect 1825 1464 1829 1544
rect 1871 1464 1875 1544
rect 1879 1464 1883 1544
rect 1955 1464 1959 1544
rect 1975 1464 1979 1504
rect 1989 1464 1993 1504
rect 2009 1464 2013 1504
rect 2021 1464 2025 1504
rect 2041 1464 2045 1504
rect 2087 1464 2091 1504
rect 2095 1464 2099 1504
rect 2115 1464 2119 1484
rect 2123 1464 2127 1484
rect 2145 1464 2149 1544
rect 2217 1464 2221 1544
rect 2225 1464 2229 1544
rect 2285 1464 2289 1504
rect 2305 1464 2309 1504
rect 2356 1464 2360 1544
rect 2364 1464 2368 1544
rect 2386 1464 2390 1504
rect 2451 1464 2455 1544
rect 2473 1464 2477 1484
rect 2481 1464 2485 1484
rect 2501 1464 2505 1504
rect 2509 1464 2513 1504
rect 2555 1464 2559 1504
rect 2575 1464 2579 1504
rect 2587 1464 2591 1504
rect 2607 1464 2611 1504
rect 2621 1464 2625 1504
rect 2641 1464 2645 1544
rect 2695 1464 2699 1544
rect 2715 1464 2719 1504
rect 2729 1464 2733 1504
rect 2749 1464 2753 1504
rect 2761 1464 2765 1504
rect 2781 1464 2785 1504
rect 2827 1464 2831 1504
rect 2835 1464 2839 1504
rect 2855 1464 2859 1484
rect 2863 1464 2867 1484
rect 2885 1464 2889 1544
rect 2931 1464 2935 1544
rect 2991 1464 2995 1504
rect 3011 1464 3015 1504
rect 3085 1464 3089 1504
rect 3105 1464 3109 1504
rect 3156 1464 3160 1544
rect 3164 1464 3168 1544
rect 3186 1464 3190 1504
rect 3251 1464 3255 1504
rect 3271 1464 3275 1504
rect 3345 1464 3349 1504
rect 3365 1464 3369 1504
rect 3430 1464 3434 1504
rect 3452 1464 3456 1544
rect 3460 1464 3464 1544
rect 3511 1464 3515 1504
rect 3531 1464 3535 1504
rect 3551 1464 3555 1504
rect 3635 1464 3639 1544
rect 3645 1464 3649 1544
rect 3675 1464 3679 1544
rect 3685 1464 3689 1544
rect 3731 1464 3735 1504
rect 3791 1464 3795 1504
rect 3811 1464 3815 1504
rect 3831 1464 3835 1504
rect 3891 1464 3895 1544
rect 3911 1464 3915 1544
rect 3931 1464 3935 1544
rect 3996 1464 4000 1544
rect 4004 1464 4008 1544
rect 4026 1464 4030 1504
rect 4105 1464 4109 1504
rect 4125 1464 4129 1504
rect 4171 1464 4175 1544
rect 4191 1464 4195 1544
rect 4211 1464 4215 1544
rect 4276 1464 4280 1544
rect 4284 1464 4288 1544
rect 4306 1464 4310 1504
rect 4371 1464 4375 1504
rect 4431 1464 4435 1544
rect 4439 1464 4443 1544
rect 4511 1464 4515 1504
rect 4531 1464 4535 1504
rect 4591 1464 4595 1504
rect 4611 1464 4615 1504
rect 4671 1464 4675 1504
rect 4691 1464 4695 1504
rect 31 1356 35 1436
rect 53 1416 57 1436
rect 61 1416 65 1436
rect 81 1396 85 1436
rect 89 1396 93 1436
rect 135 1396 139 1436
rect 155 1396 159 1436
rect 167 1396 171 1436
rect 187 1396 191 1436
rect 201 1396 205 1436
rect 221 1356 225 1436
rect 275 1356 279 1436
rect 295 1396 299 1436
rect 309 1396 313 1436
rect 329 1396 333 1436
rect 341 1396 345 1436
rect 361 1396 365 1436
rect 407 1396 411 1436
rect 415 1396 419 1436
rect 435 1416 439 1436
rect 443 1416 447 1436
rect 465 1356 469 1436
rect 511 1396 515 1436
rect 531 1396 535 1436
rect 610 1396 614 1436
rect 632 1356 636 1436
rect 640 1356 644 1436
rect 710 1396 714 1436
rect 732 1356 736 1436
rect 740 1356 744 1436
rect 803 1356 807 1436
rect 825 1396 829 1436
rect 871 1396 875 1436
rect 891 1396 895 1436
rect 970 1396 974 1436
rect 992 1356 996 1436
rect 1000 1356 1004 1436
rect 1065 1396 1069 1436
rect 1111 1356 1115 1436
rect 1131 1356 1135 1436
rect 1151 1356 1155 1436
rect 1171 1356 1175 1436
rect 1245 1396 1249 1436
rect 1265 1396 1269 1436
rect 1330 1396 1334 1436
rect 1352 1356 1356 1436
rect 1360 1356 1364 1436
rect 1425 1396 1429 1436
rect 1445 1396 1449 1436
rect 1510 1396 1514 1436
rect 1532 1356 1536 1436
rect 1540 1356 1544 1436
rect 1591 1396 1595 1436
rect 1613 1356 1617 1436
rect 1671 1396 1675 1436
rect 1691 1396 1695 1436
rect 1770 1396 1774 1436
rect 1792 1356 1796 1436
rect 1800 1356 1804 1436
rect 1851 1356 1855 1436
rect 1873 1416 1877 1436
rect 1881 1416 1885 1436
rect 1901 1396 1905 1436
rect 1909 1396 1913 1436
rect 1955 1396 1959 1436
rect 1975 1396 1979 1436
rect 1987 1396 1991 1436
rect 2007 1396 2011 1436
rect 2021 1396 2025 1436
rect 2041 1356 2045 1436
rect 2091 1396 2095 1436
rect 2156 1356 2160 1436
rect 2164 1356 2168 1436
rect 2186 1396 2190 1436
rect 2265 1396 2269 1436
rect 2285 1396 2289 1436
rect 2357 1356 2361 1436
rect 2365 1356 2369 1436
rect 2425 1396 2429 1436
rect 2471 1356 2475 1436
rect 2479 1356 2483 1436
rect 2551 1356 2555 1436
rect 2573 1416 2577 1436
rect 2581 1416 2585 1436
rect 2601 1396 2605 1436
rect 2609 1396 2613 1436
rect 2655 1396 2659 1436
rect 2675 1396 2679 1436
rect 2687 1396 2691 1436
rect 2707 1396 2711 1436
rect 2721 1396 2725 1436
rect 2741 1356 2745 1436
rect 2791 1356 2795 1436
rect 2799 1356 2803 1436
rect 2885 1356 2889 1436
rect 2936 1356 2940 1436
rect 2944 1356 2948 1436
rect 2966 1396 2970 1436
rect 3036 1356 3040 1436
rect 3044 1356 3048 1436
rect 3066 1396 3070 1436
rect 3136 1356 3140 1436
rect 3144 1356 3148 1436
rect 3166 1396 3170 1436
rect 3231 1396 3235 1436
rect 3253 1396 3257 1436
rect 3275 1356 3279 1436
rect 3357 1356 3361 1436
rect 3365 1356 3369 1436
rect 3411 1396 3415 1436
rect 3431 1396 3435 1436
rect 3451 1396 3455 1436
rect 3530 1396 3534 1436
rect 3552 1356 3556 1436
rect 3560 1356 3564 1436
rect 3616 1356 3620 1436
rect 3624 1356 3628 1436
rect 3646 1396 3650 1436
rect 3725 1396 3729 1436
rect 3745 1396 3749 1436
rect 3805 1396 3809 1436
rect 3825 1396 3829 1436
rect 3871 1396 3875 1436
rect 3893 1396 3897 1436
rect 3915 1356 3919 1436
rect 3990 1396 3994 1436
rect 4012 1356 4016 1436
rect 4020 1356 4024 1436
rect 4071 1396 4075 1436
rect 4145 1396 4149 1436
rect 4165 1396 4169 1436
rect 4225 1396 4229 1436
rect 4245 1396 4249 1436
rect 4317 1356 4321 1436
rect 4325 1356 4329 1436
rect 4390 1396 4394 1436
rect 4412 1356 4416 1436
rect 4420 1356 4424 1436
rect 4476 1356 4480 1436
rect 4484 1356 4488 1436
rect 4506 1396 4510 1436
rect 4585 1356 4589 1436
rect 4605 1356 4609 1436
rect 4625 1356 4629 1436
rect 4671 1396 4675 1436
rect 4691 1396 4695 1436
rect 31 984 35 1024
rect 105 984 109 1024
rect 125 984 129 1024
rect 190 984 194 1024
rect 212 984 216 1064
rect 220 984 224 1064
rect 271 984 275 1064
rect 291 984 295 1064
rect 311 984 315 1064
rect 331 984 335 1064
rect 405 984 409 1064
rect 425 984 429 1064
rect 445 984 449 1064
rect 515 984 519 1064
rect 535 984 539 1064
rect 545 984 549 1064
rect 591 984 595 1064
rect 599 984 603 1064
rect 681 984 685 1064
rect 703 984 707 1024
rect 725 984 729 1024
rect 783 984 787 1064
rect 805 984 809 1024
rect 877 984 881 1064
rect 885 984 889 1064
rect 945 984 949 1024
rect 1005 984 1009 1024
rect 1051 984 1055 1064
rect 1059 984 1063 1064
rect 1131 984 1135 1024
rect 1217 984 1221 1064
rect 1225 984 1229 1064
rect 1271 984 1275 1064
rect 1291 984 1295 1064
rect 1311 984 1315 1064
rect 1375 984 1379 1064
rect 1395 984 1399 1024
rect 1409 984 1413 1024
rect 1429 984 1433 1024
rect 1441 984 1445 1024
rect 1461 984 1465 1024
rect 1507 984 1511 1024
rect 1515 984 1519 1024
rect 1535 984 1539 1004
rect 1543 984 1547 1004
rect 1565 984 1569 1064
rect 1625 984 1629 1024
rect 1671 984 1675 1024
rect 1691 984 1695 1024
rect 1751 984 1755 1064
rect 1759 984 1763 1064
rect 1835 984 1839 1064
rect 1855 984 1859 1024
rect 1869 984 1873 1024
rect 1889 984 1893 1024
rect 1901 984 1905 1024
rect 1921 984 1925 1024
rect 1967 984 1971 1024
rect 1975 984 1979 1024
rect 1995 984 1999 1004
rect 2003 984 2007 1004
rect 2025 984 2029 1064
rect 2085 984 2089 1024
rect 2131 984 2135 1064
rect 2139 984 2143 1064
rect 2211 984 2215 1064
rect 2219 984 2223 1064
rect 2305 984 2309 1024
rect 2351 984 2355 1064
rect 2373 984 2377 1004
rect 2381 984 2385 1004
rect 2401 984 2405 1024
rect 2409 984 2413 1024
rect 2455 984 2459 1024
rect 2475 984 2479 1024
rect 2487 984 2491 1024
rect 2507 984 2511 1024
rect 2521 984 2525 1024
rect 2541 984 2545 1064
rect 2591 984 2595 1024
rect 2656 984 2660 1064
rect 2664 984 2668 1064
rect 2686 984 2690 1024
rect 2751 984 2755 1064
rect 2761 984 2765 1064
rect 2791 984 2795 1064
rect 2801 984 2805 1064
rect 2871 984 2875 1064
rect 2879 984 2883 1064
rect 2965 984 2969 1024
rect 2985 984 2989 1024
rect 3031 984 3035 1024
rect 3053 984 3057 1024
rect 3075 984 3079 1064
rect 3136 984 3140 1064
rect 3144 984 3148 1064
rect 3166 984 3170 1024
rect 3231 984 3235 1064
rect 3241 984 3245 1064
rect 3261 984 3265 1064
rect 3345 984 3349 1024
rect 3365 984 3369 1024
rect 3425 984 3429 1024
rect 3445 984 3449 1024
rect 3491 984 3495 1024
rect 3511 984 3515 1024
rect 3571 984 3575 1024
rect 3591 984 3595 1024
rect 3656 984 3660 1064
rect 3664 984 3668 1064
rect 3686 984 3690 1024
rect 3765 984 3769 1024
rect 3785 984 3789 1024
rect 3805 984 3809 1024
rect 3851 984 3855 1064
rect 3871 984 3875 1064
rect 3891 984 3895 1064
rect 3965 984 3969 1024
rect 4025 984 4029 1024
rect 4045 984 4049 1024
rect 4065 984 4069 1024
rect 4111 984 4115 1064
rect 4131 984 4135 1064
rect 4151 984 4155 1064
rect 4211 984 4215 1024
rect 4285 984 4289 1064
rect 4305 984 4309 1064
rect 4325 984 4329 1064
rect 4390 984 4394 1024
rect 4412 984 4416 1064
rect 4420 984 4424 1064
rect 4476 984 4480 1064
rect 4484 984 4488 1064
rect 4506 984 4510 1024
rect 4571 984 4575 1064
rect 4579 984 4583 1064
rect 4665 984 4669 1024
rect 4685 984 4689 1024
rect 4745 984 4749 1024
rect 35 876 39 956
rect 55 916 59 956
rect 69 916 73 956
rect 89 916 93 956
rect 101 916 105 956
rect 121 916 125 956
rect 167 916 171 956
rect 175 916 179 956
rect 195 936 199 956
rect 203 936 207 956
rect 225 876 229 956
rect 271 916 275 956
rect 291 916 295 956
rect 370 916 374 956
rect 392 876 396 956
rect 400 876 404 956
rect 455 876 459 956
rect 475 916 479 956
rect 489 916 493 956
rect 509 916 513 956
rect 521 916 525 956
rect 541 916 545 956
rect 587 916 591 956
rect 595 916 599 956
rect 615 936 619 956
rect 623 936 627 956
rect 645 876 649 956
rect 691 916 695 956
rect 711 916 715 956
rect 790 916 794 956
rect 812 876 816 956
rect 820 876 824 956
rect 890 916 894 956
rect 912 876 916 956
rect 920 876 924 956
rect 985 916 989 956
rect 1057 876 1061 956
rect 1065 876 1069 956
rect 1111 876 1115 956
rect 1119 876 1123 956
rect 1205 916 1209 956
rect 1225 916 1229 956
rect 1285 916 1289 956
rect 1305 916 1309 956
rect 1365 916 1369 956
rect 1385 916 1389 956
rect 1445 876 1449 956
rect 1465 876 1469 956
rect 1485 876 1489 956
rect 1541 876 1545 956
rect 1563 916 1567 956
rect 1585 916 1589 956
rect 1631 876 1635 956
rect 1651 876 1655 956
rect 1671 876 1675 956
rect 1731 876 1735 956
rect 1751 876 1755 956
rect 1771 876 1775 956
rect 1791 876 1795 956
rect 1811 876 1815 956
rect 1831 876 1835 956
rect 1851 876 1855 956
rect 1871 876 1875 956
rect 1945 916 1949 956
rect 1965 916 1969 956
rect 2037 876 2041 956
rect 2045 876 2049 956
rect 2096 876 2100 956
rect 2104 876 2108 956
rect 2126 916 2130 956
rect 2196 876 2200 956
rect 2204 876 2208 956
rect 2226 916 2230 956
rect 2296 876 2300 956
rect 2304 876 2308 956
rect 2326 916 2330 956
rect 2391 916 2395 956
rect 2411 916 2415 956
rect 2485 916 2489 956
rect 2531 876 2535 956
rect 2553 936 2557 956
rect 2561 936 2565 956
rect 2581 916 2585 956
rect 2589 916 2593 956
rect 2635 916 2639 956
rect 2655 916 2659 956
rect 2667 916 2671 956
rect 2687 916 2691 956
rect 2701 916 2705 956
rect 2721 876 2725 956
rect 2790 916 2794 956
rect 2812 876 2816 956
rect 2820 876 2824 956
rect 2885 916 2889 956
rect 2931 916 2935 956
rect 2991 916 2995 956
rect 3011 916 3015 956
rect 3031 916 3035 956
rect 3091 916 3095 956
rect 3165 916 3169 956
rect 3185 916 3189 956
rect 3231 876 3235 956
rect 3241 876 3245 956
rect 3261 876 3265 956
rect 3331 916 3335 956
rect 3351 916 3355 956
rect 3411 916 3415 956
rect 3431 916 3435 956
rect 3517 876 3521 956
rect 3525 876 3529 956
rect 3571 916 3575 956
rect 3591 916 3595 956
rect 3665 916 3669 956
rect 3685 916 3689 956
rect 3705 916 3709 956
rect 3765 916 3769 956
rect 3785 916 3789 956
rect 3805 916 3809 956
rect 3851 916 3855 956
rect 3871 916 3875 956
rect 3945 916 3949 956
rect 3965 916 3969 956
rect 3985 916 3989 956
rect 4045 916 4049 956
rect 4110 916 4114 956
rect 4132 876 4136 956
rect 4140 876 4144 956
rect 4210 916 4214 956
rect 4232 876 4236 956
rect 4240 876 4244 956
rect 4305 876 4309 956
rect 4325 876 4329 956
rect 4345 876 4349 956
rect 4391 916 4395 956
rect 4411 916 4415 956
rect 4431 916 4435 956
rect 4505 916 4509 956
rect 4525 916 4529 956
rect 4545 916 4549 956
rect 4605 876 4609 956
rect 4625 876 4629 956
rect 4645 876 4649 956
rect 4691 916 4695 956
rect 4711 916 4715 956
rect 4731 916 4735 956
rect 35 504 39 584
rect 55 504 59 544
rect 69 504 73 544
rect 89 504 93 544
rect 101 504 105 544
rect 121 504 125 544
rect 167 504 171 544
rect 175 504 179 544
rect 195 504 199 524
rect 203 504 207 524
rect 225 504 229 584
rect 271 504 275 544
rect 336 504 340 584
rect 344 504 348 584
rect 366 504 370 544
rect 431 504 435 544
rect 451 504 455 544
rect 511 504 515 544
rect 533 504 537 584
rect 605 504 609 544
rect 651 504 655 584
rect 673 504 677 524
rect 681 504 685 524
rect 701 504 705 544
rect 709 504 713 544
rect 755 504 759 544
rect 775 504 779 544
rect 787 504 791 544
rect 807 504 811 544
rect 821 504 825 544
rect 841 504 845 584
rect 896 504 900 584
rect 904 504 908 584
rect 926 504 930 544
rect 1017 504 1021 584
rect 1025 504 1029 584
rect 1071 504 1075 584
rect 1081 504 1085 584
rect 1101 504 1105 584
rect 1190 504 1194 544
rect 1212 504 1216 584
rect 1220 504 1224 584
rect 1281 504 1285 584
rect 1303 504 1307 544
rect 1325 504 1329 544
rect 1371 504 1375 584
rect 1379 504 1383 584
rect 1451 504 1455 544
rect 1473 504 1477 584
rect 1535 504 1539 584
rect 1555 504 1559 544
rect 1569 504 1573 544
rect 1589 504 1593 544
rect 1601 504 1605 544
rect 1621 504 1625 544
rect 1667 504 1671 544
rect 1675 504 1679 544
rect 1695 504 1699 524
rect 1703 504 1707 524
rect 1725 504 1729 584
rect 1771 504 1775 544
rect 1793 504 1797 584
rect 1877 504 1881 584
rect 1885 504 1889 584
rect 1957 504 1961 584
rect 1965 504 1969 584
rect 2025 504 2029 544
rect 2071 504 2075 584
rect 2079 504 2083 584
rect 2151 504 2155 584
rect 2173 504 2177 524
rect 2181 504 2185 524
rect 2201 504 2205 544
rect 2209 504 2213 544
rect 2255 504 2259 544
rect 2275 504 2279 544
rect 2287 504 2291 544
rect 2307 504 2311 544
rect 2321 504 2325 544
rect 2341 504 2345 584
rect 2391 504 2395 584
rect 2411 504 2415 584
rect 2431 504 2435 584
rect 2451 504 2455 584
rect 2535 504 2539 584
rect 2555 504 2559 584
rect 2565 504 2569 584
rect 2625 504 2629 584
rect 2645 504 2649 584
rect 2665 504 2669 584
rect 2725 504 2729 584
rect 2745 504 2749 584
rect 2765 504 2769 584
rect 2811 504 2815 544
rect 2890 504 2894 544
rect 2912 504 2916 584
rect 2920 504 2924 584
rect 2976 504 2980 584
rect 2984 504 2988 584
rect 3006 504 3010 544
rect 3071 504 3075 544
rect 3091 504 3095 544
rect 3165 504 3169 544
rect 3211 504 3215 544
rect 3285 504 3289 544
rect 3305 504 3309 544
rect 3325 504 3329 544
rect 3397 504 3401 584
rect 3405 504 3409 584
rect 3456 504 3460 584
rect 3464 504 3468 584
rect 3486 504 3490 544
rect 3551 504 3555 584
rect 3571 504 3575 584
rect 3591 504 3595 584
rect 3665 504 3669 584
rect 3685 504 3689 584
rect 3705 504 3709 584
rect 3765 504 3769 584
rect 3785 504 3789 584
rect 3805 504 3809 584
rect 3825 504 3829 584
rect 3885 504 3889 544
rect 3905 504 3909 544
rect 3925 504 3929 544
rect 3985 504 3989 544
rect 4005 504 4009 544
rect 4025 504 4029 544
rect 4071 504 4075 544
rect 4131 504 4135 544
rect 4151 504 4155 544
rect 4171 504 4175 544
rect 4231 504 4235 544
rect 4251 504 4255 544
rect 4271 504 4275 544
rect 4345 504 4349 544
rect 4365 504 4369 544
rect 4385 504 4389 544
rect 4445 504 4449 544
rect 4465 504 4469 544
rect 4485 504 4489 544
rect 4531 504 4535 544
rect 4610 504 4614 544
rect 4632 504 4636 584
rect 4640 504 4644 584
rect 4696 504 4700 584
rect 4704 504 4708 584
rect 4726 504 4730 544
rect 35 396 39 476
rect 55 436 59 476
rect 69 436 73 476
rect 89 436 93 476
rect 101 436 105 476
rect 121 436 125 476
rect 167 436 171 476
rect 175 436 179 476
rect 195 456 199 476
rect 203 456 207 476
rect 225 396 229 476
rect 271 436 275 476
rect 291 436 295 476
rect 370 436 374 476
rect 392 396 396 476
rect 400 396 404 476
rect 451 436 455 476
rect 511 436 515 476
rect 531 436 535 476
rect 610 436 614 476
rect 632 396 636 476
rect 640 396 644 476
rect 696 396 700 476
rect 704 396 708 476
rect 726 436 730 476
rect 796 396 800 476
rect 804 396 808 476
rect 826 436 830 476
rect 910 436 914 476
rect 932 396 936 476
rect 940 396 944 476
rect 991 436 995 476
rect 1051 436 1055 476
rect 1071 436 1075 476
rect 1145 396 1149 476
rect 1165 396 1169 476
rect 1185 396 1189 476
rect 1245 436 1249 476
rect 1310 436 1314 476
rect 1332 396 1336 476
rect 1340 396 1344 476
rect 1417 396 1421 476
rect 1425 396 1429 476
rect 1476 396 1480 476
rect 1484 396 1488 476
rect 1506 436 1510 476
rect 1571 436 1575 476
rect 1591 436 1595 476
rect 1651 396 1655 476
rect 1673 456 1677 476
rect 1681 456 1685 476
rect 1701 436 1705 476
rect 1709 436 1713 476
rect 1755 436 1759 476
rect 1775 436 1779 476
rect 1787 436 1791 476
rect 1807 436 1811 476
rect 1821 436 1825 476
rect 1841 396 1845 476
rect 1905 436 1909 476
rect 1925 436 1929 476
rect 1990 436 1994 476
rect 2012 396 2016 476
rect 2020 396 2024 476
rect 2075 396 2079 476
rect 2095 436 2099 476
rect 2109 436 2113 476
rect 2129 436 2133 476
rect 2141 436 2145 476
rect 2161 436 2165 476
rect 2207 436 2211 476
rect 2215 436 2219 476
rect 2235 456 2239 476
rect 2243 456 2247 476
rect 2265 396 2269 476
rect 2325 436 2329 476
rect 2371 396 2375 476
rect 2379 396 2383 476
rect 2451 436 2455 476
rect 2525 436 2529 476
rect 2545 436 2549 476
rect 2591 396 2595 476
rect 2613 456 2617 476
rect 2621 456 2625 476
rect 2641 436 2645 476
rect 2649 436 2653 476
rect 2695 436 2699 476
rect 2715 436 2719 476
rect 2727 436 2731 476
rect 2747 436 2751 476
rect 2761 436 2765 476
rect 2781 396 2785 476
rect 2831 436 2835 476
rect 2851 436 2855 476
rect 2911 396 2915 476
rect 2931 396 2935 476
rect 2951 396 2955 476
rect 2971 396 2975 476
rect 3031 396 3035 476
rect 3039 396 3043 476
rect 3111 436 3115 476
rect 3185 436 3189 476
rect 3205 436 3209 476
rect 3225 436 3229 476
rect 3285 436 3289 476
rect 3305 436 3309 476
rect 3325 436 3329 476
rect 3376 396 3380 476
rect 3384 396 3388 476
rect 3406 436 3410 476
rect 3485 436 3489 476
rect 3531 436 3535 476
rect 3551 436 3555 476
rect 3611 436 3615 476
rect 3631 436 3635 476
rect 3696 396 3700 476
rect 3704 396 3708 476
rect 3726 436 3730 476
rect 3817 396 3821 476
rect 3825 396 3829 476
rect 3897 396 3901 476
rect 3905 396 3909 476
rect 3951 436 3955 476
rect 3973 436 3977 476
rect 3995 396 3999 476
rect 4051 396 4055 476
rect 4059 396 4063 476
rect 4145 396 4149 476
rect 4165 396 4169 476
rect 4185 396 4189 476
rect 4245 436 4249 476
rect 4265 436 4269 476
rect 4285 436 4289 476
rect 4331 396 4335 476
rect 4351 396 4355 476
rect 4371 396 4375 476
rect 4431 436 4435 476
rect 4510 436 4514 476
rect 4532 396 4536 476
rect 4540 396 4544 476
rect 4591 436 4595 476
rect 4651 436 4655 476
rect 4711 436 4715 476
rect 35 24 39 104
rect 55 24 59 64
rect 69 24 73 64
rect 89 24 93 64
rect 101 24 105 64
rect 121 24 125 64
rect 167 24 171 64
rect 175 24 179 64
rect 195 24 199 44
rect 203 24 207 44
rect 225 24 229 104
rect 271 24 275 104
rect 291 24 295 104
rect 311 24 315 104
rect 331 24 335 104
rect 391 24 395 104
rect 399 24 403 104
rect 471 24 475 64
rect 491 24 495 64
rect 511 24 515 64
rect 595 24 599 104
rect 615 24 619 104
rect 625 24 629 104
rect 685 24 689 104
rect 705 24 709 104
rect 725 24 729 104
rect 771 24 775 104
rect 793 24 797 44
rect 801 24 805 44
rect 821 24 825 64
rect 829 24 833 64
rect 875 24 879 64
rect 895 24 899 64
rect 907 24 911 64
rect 927 24 931 64
rect 941 24 945 64
rect 961 24 965 104
rect 1030 24 1034 64
rect 1052 24 1056 104
rect 1060 24 1064 104
rect 1125 24 1129 64
rect 1197 24 1201 104
rect 1205 24 1209 104
rect 1265 24 1269 64
rect 1330 24 1334 64
rect 1352 24 1356 104
rect 1360 24 1364 104
rect 1425 24 1429 64
rect 1485 24 1489 64
rect 1531 24 1535 104
rect 1539 24 1543 104
rect 1625 24 1629 104
rect 1645 24 1649 104
rect 1665 24 1669 104
rect 1715 24 1719 104
rect 1735 24 1739 64
rect 1749 24 1753 64
rect 1769 24 1773 64
rect 1781 24 1785 64
rect 1801 24 1805 64
rect 1847 24 1851 64
rect 1855 24 1859 64
rect 1875 24 1879 44
rect 1883 24 1887 44
rect 1905 24 1909 104
rect 1970 24 1974 64
rect 1992 24 1996 104
rect 2000 24 2004 104
rect 2051 24 2055 64
rect 2111 24 2115 104
rect 2119 24 2123 104
rect 2191 24 2195 104
rect 2199 24 2203 104
rect 2297 24 2301 104
rect 2305 24 2309 104
rect 2351 24 2355 104
rect 2359 24 2363 104
rect 2445 24 2449 64
rect 2491 24 2495 104
rect 2513 24 2517 44
rect 2521 24 2525 44
rect 2541 24 2545 64
rect 2549 24 2553 64
rect 2595 24 2599 64
rect 2615 24 2619 64
rect 2627 24 2631 64
rect 2647 24 2651 64
rect 2661 24 2665 64
rect 2681 24 2685 104
rect 2731 24 2735 104
rect 2753 24 2757 44
rect 2761 24 2765 44
rect 2781 24 2785 64
rect 2789 24 2793 64
rect 2835 24 2839 64
rect 2855 24 2859 64
rect 2867 24 2871 64
rect 2887 24 2891 64
rect 2901 24 2905 64
rect 2921 24 2925 104
rect 2971 24 2975 104
rect 2981 24 2985 104
rect 3011 24 3015 104
rect 3021 24 3025 104
rect 3115 24 3119 104
rect 3135 24 3139 104
rect 3145 24 3149 104
rect 3196 24 3200 104
rect 3204 24 3208 104
rect 3226 24 3230 64
rect 3305 24 3309 64
rect 3351 24 3355 64
rect 3371 24 3375 64
rect 3445 24 3449 64
rect 3465 24 3469 64
rect 3485 24 3489 64
rect 3545 24 3549 64
rect 3605 24 3609 104
rect 3625 24 3629 104
rect 3645 24 3649 104
rect 3717 24 3721 104
rect 3725 24 3729 104
rect 3771 24 3775 64
rect 3836 24 3840 104
rect 3844 24 3848 104
rect 3866 24 3870 64
rect 3931 24 3935 104
rect 3939 24 3943 104
rect 4025 24 4029 64
rect 4045 24 4049 64
rect 4065 24 4069 64
rect 4111 24 4115 64
rect 4131 24 4135 64
rect 4205 24 4209 64
rect 4225 24 4229 64
rect 4245 24 4249 64
rect 4305 24 4309 64
rect 4325 24 4329 64
rect 4385 24 4389 64
rect 4405 24 4409 64
rect 4425 24 4429 64
rect 4471 24 4475 64
rect 4491 24 4495 64
rect 4551 24 4555 64
rect 4571 24 4575 64
rect 4591 24 4595 64
rect 4665 24 4669 104
rect 4685 24 4689 104
rect 4705 24 4709 104
<< ndiffusion >>
rect 41 4516 43 4556
rect 47 4516 49 4556
rect 61 4536 65 4556
rect 69 4536 71 4556
rect 131 4516 133 4556
rect 137 4516 143 4556
rect 147 4516 149 4556
rect 203 4516 205 4556
rect 209 4516 211 4556
rect 223 4516 225 4556
rect 229 4528 231 4556
rect 243 4528 245 4556
rect 229 4516 245 4528
rect 249 4516 251 4556
rect 289 4536 291 4556
rect 295 4536 299 4556
rect 311 4516 313 4556
rect 317 4516 319 4556
rect 383 4536 385 4556
rect 389 4536 391 4556
rect 403 4536 405 4556
rect 409 4536 411 4556
rect 463 4536 465 4556
rect 469 4536 471 4556
rect 483 4536 485 4556
rect 489 4536 491 4556
rect 529 4536 531 4556
rect 535 4536 539 4556
rect 551 4516 553 4556
rect 557 4516 559 4556
rect 623 4536 625 4556
rect 629 4536 631 4556
rect 669 4536 671 4556
rect 675 4536 677 4556
rect 689 4536 691 4556
rect 695 4536 697 4556
rect 749 4536 751 4556
rect 755 4536 757 4556
rect 809 4516 811 4556
rect 815 4536 819 4556
rect 831 4536 833 4556
rect 837 4536 843 4556
rect 847 4536 849 4556
rect 861 4536 863 4556
rect 867 4536 871 4556
rect 875 4536 877 4556
rect 915 4536 917 4556
rect 921 4536 925 4556
rect 937 4536 939 4556
rect 943 4536 949 4556
rect 953 4536 955 4556
rect 967 4536 971 4556
rect 975 4536 981 4556
rect 985 4536 987 4556
rect 999 4536 1001 4556
rect 815 4516 828 4536
rect 991 4516 1001 4536
rect 1005 4516 1007 4556
rect 1049 4516 1051 4556
rect 1055 4528 1057 4556
rect 1069 4528 1071 4556
rect 1055 4516 1071 4528
rect 1075 4516 1077 4556
rect 1089 4516 1091 4556
rect 1095 4516 1097 4556
rect 1149 4516 1151 4556
rect 1155 4536 1159 4556
rect 1171 4536 1173 4556
rect 1177 4536 1183 4556
rect 1187 4536 1189 4556
rect 1201 4536 1203 4556
rect 1207 4536 1211 4556
rect 1215 4536 1217 4556
rect 1255 4536 1257 4556
rect 1261 4536 1265 4556
rect 1277 4536 1279 4556
rect 1283 4536 1289 4556
rect 1293 4536 1295 4556
rect 1307 4536 1311 4556
rect 1315 4536 1321 4556
rect 1325 4536 1327 4556
rect 1339 4536 1341 4556
rect 1155 4516 1168 4536
rect 1331 4516 1341 4536
rect 1345 4516 1347 4556
rect 1389 4516 1391 4556
rect 1395 4528 1397 4556
rect 1409 4528 1411 4556
rect 1395 4516 1411 4528
rect 1415 4516 1417 4556
rect 1429 4516 1431 4556
rect 1435 4516 1437 4556
rect 1493 4516 1495 4556
rect 1499 4536 1501 4556
rect 1513 4536 1515 4556
rect 1519 4536 1525 4556
rect 1529 4536 1533 4556
rect 1545 4536 1547 4556
rect 1551 4536 1557 4556
rect 1561 4536 1563 4556
rect 1575 4536 1579 4556
rect 1583 4536 1585 4556
rect 1623 4536 1625 4556
rect 1629 4536 1633 4556
rect 1637 4536 1639 4556
rect 1651 4536 1653 4556
rect 1657 4536 1663 4556
rect 1667 4536 1669 4556
rect 1681 4536 1685 4556
rect 1499 4516 1509 4536
rect 1672 4516 1685 4536
rect 1689 4516 1691 4556
rect 1731 4516 1733 4556
rect 1737 4516 1743 4556
rect 1747 4516 1749 4556
rect 1809 4516 1811 4556
rect 1815 4536 1819 4556
rect 1831 4536 1833 4556
rect 1837 4536 1843 4556
rect 1847 4536 1849 4556
rect 1861 4536 1863 4556
rect 1867 4536 1871 4556
rect 1875 4536 1877 4556
rect 1915 4536 1917 4556
rect 1921 4536 1925 4556
rect 1937 4536 1939 4556
rect 1943 4536 1949 4556
rect 1953 4536 1955 4556
rect 1967 4536 1971 4556
rect 1975 4536 1981 4556
rect 1985 4536 1987 4556
rect 1999 4536 2001 4556
rect 1815 4516 1828 4536
rect 1991 4516 2001 4536
rect 2005 4516 2007 4556
rect 2049 4516 2051 4556
rect 2055 4526 2057 4556
rect 2069 4526 2071 4556
rect 2055 4516 2071 4526
rect 2075 4516 2077 4556
rect 2089 4516 2091 4556
rect 2095 4544 2111 4556
rect 2095 4516 2097 4544
rect 2109 4516 2111 4544
rect 2115 4516 2117 4556
rect 2206 4498 2208 4556
rect 2194 4496 2208 4498
rect 2212 4496 2216 4556
rect 2220 4496 2224 4556
rect 2228 4496 2230 4556
rect 2283 4516 2285 4556
rect 2289 4516 2291 4556
rect 2303 4516 2305 4556
rect 2309 4528 2311 4556
rect 2323 4528 2325 4556
rect 2309 4516 2325 4528
rect 2329 4516 2331 4556
rect 2383 4536 2385 4556
rect 2389 4536 2391 4556
rect 2429 4536 2431 4556
rect 2435 4536 2437 4556
rect 2449 4536 2451 4556
rect 2455 4536 2457 4556
rect 2523 4536 2525 4556
rect 2529 4536 2531 4556
rect 2569 4516 2571 4556
rect 2575 4528 2577 4556
rect 2589 4528 2591 4556
rect 2575 4516 2591 4528
rect 2595 4516 2597 4556
rect 2609 4516 2611 4556
rect 2615 4516 2617 4556
rect 2669 4536 2671 4556
rect 2675 4536 2679 4556
rect 2691 4516 2693 4556
rect 2697 4516 2699 4556
rect 2749 4536 2751 4556
rect 2755 4536 2759 4556
rect 2771 4516 2773 4556
rect 2777 4516 2779 4556
rect 2841 4516 2843 4556
rect 2847 4516 2849 4556
rect 2861 4536 2865 4556
rect 2869 4536 2871 4556
rect 2946 4498 2948 4556
rect 2934 4496 2948 4498
rect 2952 4496 2956 4556
rect 2960 4496 2964 4556
rect 2968 4496 2970 4556
rect 3033 4516 3035 4556
rect 3039 4516 3041 4556
rect 3053 4516 3055 4556
rect 3059 4516 3065 4556
rect 3069 4516 3071 4556
rect 3121 4516 3123 4556
rect 3127 4516 3129 4556
rect 3141 4536 3145 4556
rect 3149 4536 3151 4556
rect 3226 4498 3228 4556
rect 3214 4496 3228 4498
rect 3232 4496 3236 4556
rect 3240 4496 3244 4556
rect 3248 4496 3250 4556
rect 3291 4516 3293 4556
rect 3297 4516 3303 4556
rect 3307 4516 3309 4556
rect 3372 4516 3374 4556
rect 3378 4516 3382 4556
rect 3386 4516 3388 4556
rect 3400 4536 3404 4556
rect 3408 4536 3410 4556
rect 3469 4536 3471 4556
rect 3475 4536 3477 4556
rect 3531 4516 3533 4556
rect 3537 4516 3543 4556
rect 3547 4516 3549 4556
rect 3610 4496 3612 4556
rect 3616 4496 3620 4556
rect 3624 4496 3628 4556
rect 3632 4498 3634 4556
rect 3712 4516 3714 4556
rect 3718 4516 3722 4556
rect 3726 4516 3728 4556
rect 3740 4536 3744 4556
rect 3748 4536 3750 4556
rect 3632 4496 3646 4498
rect 3809 4516 3811 4556
rect 3815 4528 3817 4556
rect 3829 4528 3831 4556
rect 3815 4516 3831 4528
rect 3835 4516 3837 4556
rect 3849 4516 3851 4556
rect 3855 4516 3857 4556
rect 3923 4516 3925 4556
rect 3929 4516 3931 4556
rect 3943 4516 3945 4556
rect 3949 4528 3951 4556
rect 3963 4528 3965 4556
rect 3949 4516 3965 4528
rect 3969 4516 3971 4556
rect 4046 4498 4048 4556
rect 4034 4496 4048 4498
rect 4052 4496 4056 4556
rect 4060 4496 4064 4556
rect 4068 4496 4070 4556
rect 4146 4498 4148 4556
rect 4134 4496 4148 4498
rect 4152 4496 4156 4556
rect 4160 4496 4164 4556
rect 4168 4496 4170 4556
rect 4212 4516 4214 4556
rect 4218 4516 4222 4556
rect 4226 4516 4228 4556
rect 4240 4536 4244 4556
rect 4248 4536 4250 4556
rect 4311 4516 4313 4556
rect 4317 4516 4323 4556
rect 4327 4516 4329 4556
rect 4410 4536 4412 4556
rect 4416 4536 4420 4556
rect 4432 4516 4434 4556
rect 4438 4516 4442 4556
rect 4446 4516 4448 4556
rect 4503 4536 4505 4556
rect 4509 4536 4511 4556
rect 4550 4496 4552 4556
rect 4556 4496 4560 4556
rect 4564 4496 4568 4556
rect 4572 4498 4574 4556
rect 4572 4496 4586 4498
rect 4650 4496 4652 4556
rect 4656 4496 4660 4556
rect 4664 4496 4668 4556
rect 4672 4498 4674 4556
rect 4672 4496 4686 4498
rect 43 4104 45 4144
rect 49 4104 51 4144
rect 63 4104 65 4144
rect 69 4132 85 4144
rect 69 4104 71 4132
rect 83 4104 85 4132
rect 89 4104 91 4144
rect 153 4104 155 4144
rect 159 4104 161 4144
rect 173 4104 175 4144
rect 179 4104 185 4144
rect 189 4104 191 4144
rect 229 4104 231 4124
rect 235 4104 237 4124
rect 249 4104 251 4124
rect 255 4104 257 4124
rect 330 4104 332 4124
rect 336 4104 340 4124
rect 352 4104 354 4144
rect 358 4104 362 4144
rect 366 4104 368 4144
rect 409 4104 411 4144
rect 415 4104 421 4144
rect 425 4104 427 4144
rect 439 4104 441 4144
rect 445 4104 447 4144
rect 530 4104 532 4124
rect 536 4104 540 4124
rect 552 4104 554 4144
rect 558 4104 562 4144
rect 566 4104 568 4144
rect 610 4104 612 4164
rect 616 4104 620 4164
rect 624 4104 628 4164
rect 632 4162 646 4164
rect 632 4104 634 4162
rect 712 4104 714 4144
rect 718 4104 722 4144
rect 726 4104 728 4144
rect 740 4104 744 4124
rect 748 4104 750 4124
rect 809 4104 811 4144
rect 815 4104 821 4144
rect 825 4104 827 4144
rect 839 4104 841 4144
rect 845 4104 847 4144
rect 923 4104 925 4144
rect 929 4104 931 4144
rect 943 4104 945 4144
rect 949 4132 965 4144
rect 949 4104 951 4132
rect 963 4104 965 4132
rect 969 4104 971 4144
rect 1023 4104 1025 4124
rect 1029 4104 1031 4124
rect 1069 4104 1071 4124
rect 1075 4104 1077 4124
rect 1089 4104 1091 4124
rect 1095 4104 1097 4124
rect 1149 4104 1151 4124
rect 1155 4104 1157 4124
rect 1169 4104 1171 4124
rect 1175 4104 1177 4124
rect 1229 4104 1231 4124
rect 1235 4104 1237 4124
rect 1249 4104 1251 4124
rect 1255 4104 1257 4124
rect 1309 4104 1311 4124
rect 1315 4104 1317 4124
rect 1369 4104 1371 4144
rect 1375 4124 1388 4144
rect 1551 4124 1561 4144
rect 1375 4104 1379 4124
rect 1391 4104 1393 4124
rect 1397 4104 1403 4124
rect 1407 4104 1409 4124
rect 1421 4104 1423 4124
rect 1427 4104 1431 4124
rect 1435 4104 1437 4124
rect 1475 4104 1477 4124
rect 1481 4104 1485 4124
rect 1497 4104 1499 4124
rect 1503 4104 1509 4124
rect 1513 4104 1515 4124
rect 1527 4104 1531 4124
rect 1535 4104 1541 4124
rect 1545 4104 1547 4124
rect 1559 4104 1561 4124
rect 1565 4104 1567 4144
rect 1609 4104 1611 4144
rect 1615 4132 1631 4144
rect 1615 4104 1617 4132
rect 1629 4104 1631 4132
rect 1635 4104 1637 4144
rect 1649 4104 1651 4144
rect 1655 4104 1657 4144
rect 1709 4104 1711 4124
rect 1715 4104 1717 4124
rect 1729 4104 1731 4124
rect 1735 4104 1737 4124
rect 1803 4104 1805 4124
rect 1809 4104 1811 4124
rect 1849 4104 1851 4144
rect 1855 4124 1868 4144
rect 2031 4124 2041 4144
rect 1855 4104 1859 4124
rect 1871 4104 1873 4124
rect 1877 4104 1883 4124
rect 1887 4104 1889 4124
rect 1901 4104 1903 4124
rect 1907 4104 1911 4124
rect 1915 4104 1917 4124
rect 1955 4104 1957 4124
rect 1961 4104 1965 4124
rect 1977 4104 1979 4124
rect 1983 4104 1989 4124
rect 1993 4104 1995 4124
rect 2007 4104 2011 4124
rect 2015 4104 2021 4124
rect 2025 4104 2027 4124
rect 2039 4104 2041 4124
rect 2045 4104 2047 4144
rect 2111 4104 2113 4144
rect 2117 4104 2123 4144
rect 2127 4104 2129 4144
rect 2199 4124 2211 4144
rect 2169 4104 2171 4124
rect 2175 4104 2177 4124
rect 2189 4104 2191 4124
rect 2195 4104 2197 4124
rect 2209 4104 2211 4124
rect 2215 4104 2217 4144
rect 2304 4104 2306 4144
rect 2310 4104 2314 4144
rect 2318 4104 2320 4144
rect 2332 4104 2334 4144
rect 2338 4104 2342 4144
rect 2346 4104 2348 4144
rect 2391 4104 2393 4144
rect 2397 4104 2403 4144
rect 2407 4104 2409 4144
rect 2483 4104 2485 4144
rect 2489 4104 2491 4144
rect 2503 4104 2505 4144
rect 2509 4132 2525 4144
rect 2509 4104 2511 4132
rect 2523 4104 2525 4132
rect 2529 4104 2531 4144
rect 2583 4104 2585 4124
rect 2589 4104 2591 4124
rect 2603 4104 2605 4124
rect 2609 4104 2611 4124
rect 2652 4104 2654 4144
rect 2658 4104 2662 4144
rect 2666 4104 2668 4144
rect 2680 4104 2684 4124
rect 2688 4104 2690 4124
rect 2770 4104 2772 4124
rect 2776 4104 2780 4124
rect 2792 4104 2794 4144
rect 2798 4104 2802 4144
rect 2806 4104 2808 4144
rect 2954 4162 2968 4164
rect 2849 4104 2851 4124
rect 2855 4104 2859 4124
rect 2871 4104 2873 4144
rect 2877 4104 2879 4144
rect 2966 4104 2968 4162
rect 2972 4104 2976 4164
rect 2980 4104 2984 4164
rect 2988 4104 2990 4164
rect 3054 4162 3068 4164
rect 3066 4104 3068 4162
rect 3072 4104 3076 4164
rect 3080 4104 3084 4164
rect 3088 4104 3090 4164
rect 3131 4104 3133 4144
rect 3137 4104 3143 4144
rect 3147 4104 3149 4144
rect 3294 4162 3308 4164
rect 3223 4104 3225 4124
rect 3229 4104 3231 4124
rect 3306 4104 3308 4162
rect 3312 4104 3316 4164
rect 3320 4104 3324 4164
rect 3328 4104 3330 4164
rect 3394 4162 3408 4164
rect 3406 4104 3408 4162
rect 3412 4104 3416 4164
rect 3420 4104 3424 4164
rect 3428 4104 3430 4164
rect 3494 4162 3508 4164
rect 3506 4104 3508 4162
rect 3512 4104 3516 4164
rect 3520 4104 3524 4164
rect 3528 4104 3530 4164
rect 3594 4162 3608 4164
rect 3606 4104 3608 4162
rect 3612 4104 3616 4164
rect 3620 4104 3624 4164
rect 3628 4104 3630 4164
rect 3670 4104 3672 4164
rect 3676 4104 3680 4164
rect 3684 4104 3688 4164
rect 3692 4162 3706 4164
rect 3692 4104 3694 4162
rect 3772 4104 3774 4144
rect 3778 4104 3782 4144
rect 3786 4104 3788 4144
rect 3800 4104 3804 4124
rect 3808 4104 3810 4124
rect 3869 4104 3871 4144
rect 3875 4132 3891 4144
rect 3875 4104 3877 4132
rect 3889 4104 3891 4132
rect 3895 4104 3897 4144
rect 3909 4104 3911 4144
rect 3915 4104 3917 4144
rect 3969 4104 3971 4124
rect 3975 4104 3977 4124
rect 4032 4104 4034 4144
rect 4038 4104 4042 4144
rect 4046 4104 4048 4144
rect 4154 4162 4168 4164
rect 4060 4104 4064 4124
rect 4068 4104 4070 4124
rect 4166 4104 4168 4162
rect 4172 4104 4176 4164
rect 4180 4104 4184 4164
rect 4188 4104 4190 4164
rect 4230 4104 4232 4164
rect 4236 4104 4240 4164
rect 4244 4104 4248 4164
rect 4252 4162 4266 4164
rect 4252 4104 4254 4162
rect 4332 4104 4334 4144
rect 4338 4104 4342 4144
rect 4346 4104 4348 4144
rect 4360 4104 4364 4124
rect 4368 4104 4370 4124
rect 4429 4104 4431 4144
rect 4435 4132 4451 4144
rect 4435 4104 4437 4132
rect 4449 4104 4451 4132
rect 4455 4104 4457 4144
rect 4469 4104 4471 4144
rect 4475 4104 4477 4144
rect 4532 4104 4534 4144
rect 4538 4104 4542 4144
rect 4546 4104 4548 4144
rect 4560 4104 4562 4144
rect 4566 4104 4570 4144
rect 4574 4104 4576 4144
rect 4663 4104 4665 4124
rect 4669 4104 4671 4124
rect 4683 4104 4685 4124
rect 4689 4104 4691 4124
rect 51 4036 53 4076
rect 57 4036 63 4076
rect 67 4036 69 4076
rect 131 4036 133 4076
rect 137 4036 143 4076
rect 147 4036 149 4076
rect 203 4056 205 4076
rect 209 4056 211 4076
rect 223 4056 225 4076
rect 229 4056 231 4076
rect 269 4036 271 4076
rect 275 4048 277 4076
rect 289 4048 291 4076
rect 275 4036 291 4048
rect 295 4036 297 4076
rect 309 4036 311 4076
rect 315 4036 317 4076
rect 383 4056 385 4076
rect 389 4056 391 4076
rect 443 4056 445 4076
rect 449 4056 451 4076
rect 503 4056 505 4076
rect 509 4056 511 4076
rect 523 4056 525 4076
rect 529 4056 531 4076
rect 569 4036 571 4076
rect 575 4036 581 4076
rect 585 4036 587 4076
rect 599 4036 601 4076
rect 605 4036 607 4076
rect 669 4036 671 4076
rect 675 4048 677 4076
rect 689 4048 691 4076
rect 675 4036 691 4048
rect 695 4036 697 4076
rect 709 4036 711 4076
rect 715 4036 717 4076
rect 769 4056 771 4076
rect 775 4056 777 4076
rect 829 4036 831 4076
rect 835 4048 837 4076
rect 849 4048 851 4076
rect 835 4036 851 4048
rect 855 4036 857 4076
rect 869 4036 871 4076
rect 875 4036 877 4076
rect 931 4036 933 4076
rect 937 4036 943 4076
rect 947 4036 949 4076
rect 1023 4056 1025 4076
rect 1029 4056 1031 4076
rect 1083 4056 1085 4076
rect 1089 4056 1091 4076
rect 1103 4056 1105 4076
rect 1109 4056 1111 4076
rect 1149 4056 1151 4076
rect 1155 4056 1157 4076
rect 1209 4056 1211 4076
rect 1215 4056 1217 4076
rect 1229 4056 1231 4076
rect 1235 4056 1237 4076
rect 1289 4056 1291 4076
rect 1295 4056 1297 4076
rect 1363 4056 1365 4076
rect 1369 4056 1371 4076
rect 1383 4056 1385 4076
rect 1389 4056 1391 4076
rect 1443 4056 1445 4076
rect 1449 4056 1451 4076
rect 1489 4036 1491 4076
rect 1495 4048 1497 4076
rect 1509 4048 1511 4076
rect 1495 4036 1511 4048
rect 1515 4036 1517 4076
rect 1529 4036 1531 4076
rect 1535 4036 1537 4076
rect 1589 4036 1591 4076
rect 1595 4046 1597 4076
rect 1609 4046 1611 4076
rect 1595 4036 1611 4046
rect 1615 4036 1617 4076
rect 1629 4036 1631 4076
rect 1635 4064 1651 4076
rect 1635 4036 1637 4064
rect 1649 4036 1651 4064
rect 1655 4036 1657 4076
rect 1711 4036 1713 4076
rect 1717 4036 1723 4076
rect 1727 4036 1729 4076
rect 1810 4056 1812 4076
rect 1816 4056 1820 4076
rect 1832 4036 1834 4076
rect 1838 4036 1842 4076
rect 1846 4036 1848 4076
rect 1890 4016 1892 4076
rect 1896 4016 1900 4076
rect 1904 4016 1908 4076
rect 1912 4018 1914 4076
rect 2003 4036 2005 4076
rect 2009 4036 2011 4076
rect 2023 4036 2025 4076
rect 2029 4048 2031 4076
rect 2043 4048 2045 4076
rect 2029 4036 2045 4048
rect 2049 4036 2051 4076
rect 2103 4056 2105 4076
rect 2109 4056 2111 4076
rect 1912 4016 1926 4018
rect 2186 4018 2188 4076
rect 2174 4016 2188 4018
rect 2192 4016 2196 4076
rect 2200 4016 2204 4076
rect 2208 4016 2210 4076
rect 2286 4018 2288 4076
rect 2274 4016 2288 4018
rect 2292 4016 2296 4076
rect 2300 4016 2304 4076
rect 2308 4016 2310 4076
rect 2370 4056 2372 4076
rect 2376 4056 2380 4076
rect 2392 4036 2394 4076
rect 2398 4036 2402 4076
rect 2406 4036 2408 4076
rect 2463 4056 2465 4076
rect 2469 4056 2471 4076
rect 2523 4036 2525 4076
rect 2529 4036 2531 4076
rect 2543 4036 2545 4076
rect 2549 4048 2551 4076
rect 2563 4048 2565 4076
rect 2549 4036 2565 4048
rect 2569 4036 2571 4076
rect 2646 4018 2648 4076
rect 2634 4016 2648 4018
rect 2652 4016 2656 4076
rect 2660 4016 2664 4076
rect 2668 4016 2670 4076
rect 2730 4056 2732 4076
rect 2736 4056 2740 4076
rect 2752 4036 2754 4076
rect 2758 4036 2762 4076
rect 2766 4036 2768 4076
rect 2823 4036 2825 4076
rect 2829 4036 2831 4076
rect 2843 4036 2845 4076
rect 2849 4048 2851 4076
rect 2863 4048 2865 4076
rect 2849 4036 2865 4048
rect 2869 4036 2871 4076
rect 2909 4036 2911 4076
rect 2915 4048 2917 4076
rect 2929 4048 2931 4076
rect 2915 4036 2931 4048
rect 2935 4036 2937 4076
rect 2949 4036 2951 4076
rect 2955 4036 2957 4076
rect 3046 4018 3048 4076
rect 3034 4016 3048 4018
rect 3052 4016 3056 4076
rect 3060 4016 3064 4076
rect 3068 4016 3070 4076
rect 3123 4056 3125 4076
rect 3129 4056 3131 4076
rect 3169 4036 3171 4076
rect 3175 4048 3177 4076
rect 3189 4048 3191 4076
rect 3175 4036 3191 4048
rect 3195 4036 3197 4076
rect 3209 4036 3211 4076
rect 3215 4036 3217 4076
rect 3272 4036 3274 4076
rect 3278 4036 3282 4076
rect 3286 4036 3288 4076
rect 3300 4056 3304 4076
rect 3308 4056 3310 4076
rect 3369 4036 3371 4076
rect 3375 4048 3377 4076
rect 3389 4048 3391 4076
rect 3375 4036 3391 4048
rect 3395 4036 3397 4076
rect 3409 4036 3411 4076
rect 3415 4036 3417 4076
rect 3483 4036 3485 4076
rect 3489 4036 3491 4076
rect 3503 4036 3505 4076
rect 3509 4048 3511 4076
rect 3523 4048 3525 4076
rect 3509 4036 3525 4048
rect 3529 4036 3531 4076
rect 3583 4036 3585 4076
rect 3589 4036 3591 4076
rect 3603 4036 3605 4076
rect 3609 4048 3611 4076
rect 3623 4048 3625 4076
rect 3609 4036 3625 4048
rect 3629 4036 3631 4076
rect 3690 4056 3692 4076
rect 3696 4056 3700 4076
rect 3712 4036 3714 4076
rect 3718 4036 3722 4076
rect 3726 4036 3728 4076
rect 3806 4018 3808 4076
rect 3794 4016 3808 4018
rect 3812 4016 3816 4076
rect 3820 4016 3824 4076
rect 3828 4016 3830 4076
rect 3891 4036 3893 4076
rect 3897 4036 3903 4076
rect 3907 4036 3909 4076
rect 3971 4036 3973 4076
rect 3977 4036 3983 4076
rect 3987 4036 3989 4076
rect 4031 4036 4033 4076
rect 4037 4036 4043 4076
rect 4047 4036 4049 4076
rect 4146 4018 4148 4076
rect 4134 4016 4148 4018
rect 4152 4016 4156 4076
rect 4160 4016 4164 4076
rect 4168 4016 4170 4076
rect 4223 4036 4225 4076
rect 4229 4036 4231 4076
rect 4243 4036 4245 4076
rect 4249 4048 4251 4076
rect 4263 4048 4265 4076
rect 4249 4036 4265 4048
rect 4269 4036 4271 4076
rect 4309 4036 4311 4076
rect 4315 4048 4317 4076
rect 4329 4048 4331 4076
rect 4315 4036 4331 4048
rect 4335 4036 4337 4076
rect 4349 4036 4351 4076
rect 4355 4036 4357 4076
rect 4423 4056 4425 4076
rect 4429 4056 4431 4076
rect 4506 4018 4508 4076
rect 4494 4016 4508 4018
rect 4512 4016 4516 4076
rect 4520 4016 4524 4076
rect 4528 4016 4530 4076
rect 4606 4018 4608 4076
rect 4594 4016 4608 4018
rect 4612 4016 4616 4076
rect 4620 4016 4624 4076
rect 4628 4016 4630 4076
rect 4672 4036 4674 4076
rect 4678 4036 4682 4076
rect 4686 4036 4688 4076
rect 4700 4056 4704 4076
rect 4708 4056 4710 4076
rect 43 3624 45 3664
rect 49 3624 51 3664
rect 63 3624 65 3664
rect 69 3652 85 3664
rect 69 3624 71 3652
rect 83 3624 85 3652
rect 89 3624 91 3664
rect 143 3624 145 3644
rect 149 3624 151 3644
rect 189 3624 191 3664
rect 195 3644 208 3664
rect 371 3644 381 3664
rect 195 3624 199 3644
rect 211 3624 213 3644
rect 217 3624 223 3644
rect 227 3624 229 3644
rect 241 3624 243 3644
rect 247 3624 251 3644
rect 255 3624 257 3644
rect 295 3624 297 3644
rect 301 3624 305 3644
rect 317 3624 319 3644
rect 323 3624 329 3644
rect 333 3624 335 3644
rect 347 3624 351 3644
rect 355 3624 361 3644
rect 365 3624 367 3644
rect 379 3624 381 3644
rect 385 3624 387 3664
rect 443 3624 445 3664
rect 449 3624 451 3664
rect 463 3624 465 3664
rect 469 3652 485 3664
rect 469 3624 471 3652
rect 483 3624 485 3652
rect 489 3624 491 3664
rect 529 3624 531 3664
rect 535 3624 541 3664
rect 545 3624 547 3664
rect 559 3624 561 3664
rect 565 3624 567 3664
rect 643 3624 645 3664
rect 649 3644 661 3664
rect 649 3624 651 3644
rect 663 3624 665 3644
rect 669 3624 671 3644
rect 683 3624 685 3644
rect 689 3624 691 3644
rect 751 3624 753 3664
rect 757 3624 763 3664
rect 767 3624 769 3664
rect 813 3624 815 3664
rect 819 3644 829 3664
rect 992 3644 1005 3664
rect 819 3624 821 3644
rect 833 3624 835 3644
rect 839 3624 845 3644
rect 849 3624 853 3644
rect 865 3624 867 3644
rect 871 3624 877 3644
rect 881 3624 883 3644
rect 895 3624 899 3644
rect 903 3624 905 3644
rect 943 3624 945 3644
rect 949 3624 953 3644
rect 957 3624 959 3644
rect 971 3624 973 3644
rect 977 3624 983 3644
rect 987 3624 989 3644
rect 1001 3624 1005 3644
rect 1009 3624 1011 3664
rect 1061 3624 1063 3664
rect 1067 3624 1069 3664
rect 1081 3624 1085 3644
rect 1089 3624 1091 3644
rect 1129 3624 1131 3664
rect 1135 3644 1148 3664
rect 1311 3644 1321 3664
rect 1135 3624 1139 3644
rect 1151 3624 1153 3644
rect 1157 3624 1163 3644
rect 1167 3624 1169 3644
rect 1181 3624 1183 3644
rect 1187 3624 1191 3644
rect 1195 3624 1197 3644
rect 1235 3624 1237 3644
rect 1241 3624 1245 3644
rect 1257 3624 1259 3644
rect 1263 3624 1269 3644
rect 1273 3624 1275 3644
rect 1287 3624 1291 3644
rect 1295 3624 1301 3644
rect 1305 3624 1307 3644
rect 1319 3624 1321 3644
rect 1325 3624 1327 3664
rect 1369 3624 1371 3664
rect 1375 3652 1391 3664
rect 1375 3624 1377 3652
rect 1389 3624 1391 3652
rect 1395 3624 1397 3664
rect 1409 3624 1411 3664
rect 1415 3624 1417 3664
rect 1471 3624 1473 3664
rect 1477 3624 1483 3664
rect 1487 3624 1489 3664
rect 1551 3624 1553 3664
rect 1557 3624 1563 3664
rect 1567 3624 1569 3664
rect 1629 3624 1631 3644
rect 1635 3624 1639 3644
rect 1651 3624 1653 3664
rect 1657 3624 1659 3664
rect 1709 3624 1711 3664
rect 1715 3644 1728 3664
rect 1891 3644 1901 3664
rect 1715 3624 1719 3644
rect 1731 3624 1733 3644
rect 1737 3624 1743 3644
rect 1747 3624 1749 3644
rect 1761 3624 1763 3644
rect 1767 3624 1771 3644
rect 1775 3624 1777 3644
rect 1815 3624 1817 3644
rect 1821 3624 1825 3644
rect 1837 3624 1839 3644
rect 1843 3624 1849 3644
rect 1853 3624 1855 3644
rect 1867 3624 1871 3644
rect 1875 3624 1881 3644
rect 1885 3624 1887 3644
rect 1899 3624 1901 3644
rect 1905 3624 1907 3664
rect 1963 3624 1965 3644
rect 1969 3624 1971 3644
rect 2030 3624 2032 3644
rect 2036 3624 2040 3644
rect 2052 3624 2054 3664
rect 2058 3624 2062 3664
rect 2066 3624 2068 3664
rect 2123 3624 2125 3644
rect 2129 3624 2131 3644
rect 2170 3624 2172 3684
rect 2176 3624 2180 3684
rect 2184 3624 2188 3684
rect 2192 3682 2206 3684
rect 2192 3624 2194 3682
rect 2394 3682 2408 3684
rect 2283 3624 2285 3664
rect 2289 3624 2291 3664
rect 2303 3624 2305 3664
rect 2309 3652 2325 3664
rect 2309 3624 2311 3652
rect 2323 3624 2325 3652
rect 2329 3624 2331 3664
rect 2406 3624 2408 3682
rect 2412 3624 2416 3684
rect 2420 3624 2424 3684
rect 2428 3624 2430 3684
rect 2594 3682 2608 3684
rect 2490 3624 2492 3644
rect 2496 3624 2500 3644
rect 2512 3624 2514 3664
rect 2518 3624 2522 3664
rect 2526 3624 2528 3664
rect 2606 3624 2608 3682
rect 2612 3624 2616 3684
rect 2620 3624 2624 3684
rect 2628 3624 2630 3684
rect 2672 3624 2674 3664
rect 2678 3624 2682 3664
rect 2686 3624 2688 3664
rect 2700 3624 2704 3644
rect 2708 3624 2710 3644
rect 2790 3624 2792 3644
rect 2796 3624 2800 3644
rect 2812 3624 2814 3664
rect 2818 3624 2822 3664
rect 2826 3624 2828 3664
rect 3014 3682 3028 3684
rect 2883 3624 2885 3644
rect 2889 3624 2891 3644
rect 2943 3624 2945 3644
rect 2949 3624 2951 3644
rect 3026 3624 3028 3682
rect 3032 3624 3036 3684
rect 3040 3624 3044 3684
rect 3048 3624 3050 3684
rect 3214 3682 3228 3684
rect 3110 3624 3112 3644
rect 3116 3624 3120 3644
rect 3132 3624 3134 3664
rect 3138 3624 3142 3664
rect 3146 3624 3148 3664
rect 3226 3624 3228 3682
rect 3232 3624 3236 3684
rect 3240 3624 3244 3684
rect 3248 3624 3250 3684
rect 3303 3624 3305 3644
rect 3309 3624 3311 3644
rect 3363 3624 3365 3664
rect 3369 3624 3371 3664
rect 3383 3624 3385 3664
rect 3389 3652 3405 3664
rect 3389 3624 3391 3652
rect 3403 3624 3405 3652
rect 3409 3624 3411 3664
rect 3471 3624 3473 3664
rect 3477 3624 3483 3664
rect 3487 3624 3489 3664
rect 3529 3624 3531 3664
rect 3535 3624 3541 3664
rect 3545 3624 3547 3664
rect 3559 3624 3561 3664
rect 3565 3624 3567 3664
rect 3754 3682 3768 3684
rect 3650 3624 3652 3644
rect 3656 3624 3660 3644
rect 3672 3624 3674 3664
rect 3678 3624 3682 3664
rect 3686 3624 3688 3664
rect 3766 3624 3768 3682
rect 3772 3624 3776 3684
rect 3780 3624 3784 3684
rect 3788 3624 3790 3684
rect 3843 3624 3845 3644
rect 3849 3624 3851 3644
rect 3892 3624 3894 3664
rect 3898 3624 3902 3664
rect 3906 3624 3908 3664
rect 3920 3624 3924 3644
rect 3928 3624 3930 3644
rect 4003 3624 4005 3664
rect 4009 3624 4011 3664
rect 4023 3624 4025 3664
rect 4029 3652 4045 3664
rect 4029 3624 4031 3652
rect 4043 3624 4045 3652
rect 4049 3624 4051 3664
rect 4089 3624 4091 3664
rect 4095 3652 4111 3664
rect 4095 3624 4097 3652
rect 4109 3624 4111 3652
rect 4115 3624 4117 3664
rect 4129 3624 4131 3664
rect 4135 3624 4137 3664
rect 4192 3624 4194 3664
rect 4198 3624 4202 3664
rect 4206 3624 4208 3664
rect 4220 3624 4224 3644
rect 4228 3624 4230 3644
rect 4310 3624 4312 3644
rect 4316 3624 4320 3644
rect 4332 3624 4334 3664
rect 4338 3624 4342 3664
rect 4346 3624 4348 3664
rect 4390 3624 4392 3684
rect 4396 3624 4400 3684
rect 4404 3624 4408 3684
rect 4412 3682 4426 3684
rect 4412 3624 4414 3682
rect 4574 3682 4588 3684
rect 4503 3624 4505 3644
rect 4509 3624 4511 3644
rect 4586 3624 4588 3682
rect 4592 3624 4596 3684
rect 4600 3624 4604 3684
rect 4608 3624 4610 3684
rect 4650 3624 4652 3684
rect 4656 3624 4660 3684
rect 4664 3624 4668 3684
rect 4672 3682 4686 3684
rect 4672 3624 4674 3682
rect 33 3556 35 3596
rect 39 3576 41 3596
rect 53 3576 55 3596
rect 59 3576 65 3596
rect 69 3576 73 3596
rect 85 3576 87 3596
rect 91 3576 97 3596
rect 101 3576 103 3596
rect 115 3576 119 3596
rect 123 3576 125 3596
rect 163 3576 165 3596
rect 169 3576 173 3596
rect 177 3576 179 3596
rect 191 3576 193 3596
rect 197 3576 203 3596
rect 207 3576 209 3596
rect 221 3576 225 3596
rect 39 3556 49 3576
rect 212 3556 225 3576
rect 229 3556 231 3596
rect 291 3556 293 3596
rect 297 3556 303 3596
rect 307 3556 309 3596
rect 363 3556 365 3596
rect 369 3556 371 3596
rect 383 3556 385 3596
rect 389 3568 391 3596
rect 403 3568 405 3596
rect 389 3556 405 3568
rect 409 3556 411 3596
rect 471 3556 473 3596
rect 477 3556 483 3596
rect 487 3556 489 3596
rect 566 3538 568 3596
rect 554 3536 568 3538
rect 572 3536 576 3596
rect 580 3536 584 3596
rect 588 3536 590 3596
rect 643 3576 645 3596
rect 649 3576 651 3596
rect 703 3556 705 3596
rect 709 3556 711 3596
rect 723 3556 725 3596
rect 729 3568 731 3596
rect 743 3568 745 3596
rect 729 3556 745 3568
rect 749 3556 751 3596
rect 803 3556 805 3596
rect 809 3556 811 3596
rect 823 3556 825 3596
rect 829 3568 831 3596
rect 843 3568 845 3596
rect 829 3556 845 3568
rect 849 3556 851 3596
rect 889 3576 891 3596
rect 895 3576 897 3596
rect 963 3576 965 3596
rect 969 3576 971 3596
rect 983 3576 985 3596
rect 989 3576 991 3596
rect 1029 3556 1031 3596
rect 1035 3576 1039 3596
rect 1051 3576 1053 3596
rect 1057 3576 1063 3596
rect 1067 3576 1069 3596
rect 1081 3576 1083 3596
rect 1087 3576 1091 3596
rect 1095 3576 1097 3596
rect 1135 3576 1137 3596
rect 1141 3576 1145 3596
rect 1157 3576 1159 3596
rect 1163 3576 1169 3596
rect 1173 3576 1175 3596
rect 1187 3576 1191 3596
rect 1195 3576 1201 3596
rect 1205 3576 1207 3596
rect 1219 3576 1221 3596
rect 1035 3556 1048 3576
rect 1211 3556 1221 3576
rect 1225 3556 1227 3596
rect 1269 3576 1271 3596
rect 1275 3576 1277 3596
rect 1329 3576 1331 3596
rect 1335 3576 1337 3596
rect 1349 3576 1351 3596
rect 1355 3576 1357 3596
rect 1409 3556 1411 3596
rect 1415 3568 1417 3596
rect 1429 3568 1431 3596
rect 1415 3556 1431 3568
rect 1435 3556 1437 3596
rect 1449 3556 1451 3596
rect 1455 3556 1457 3596
rect 1511 3556 1513 3596
rect 1517 3556 1523 3596
rect 1527 3556 1529 3596
rect 1601 3556 1603 3596
rect 1607 3556 1609 3596
rect 1621 3576 1625 3596
rect 1629 3576 1631 3596
rect 1683 3576 1685 3596
rect 1689 3576 1691 3596
rect 1729 3556 1731 3596
rect 1735 3576 1739 3596
rect 1751 3576 1753 3596
rect 1757 3576 1763 3596
rect 1767 3576 1769 3596
rect 1781 3576 1783 3596
rect 1787 3576 1791 3596
rect 1795 3576 1797 3596
rect 1835 3576 1837 3596
rect 1841 3576 1845 3596
rect 1857 3576 1859 3596
rect 1863 3576 1869 3596
rect 1873 3576 1875 3596
rect 1887 3576 1891 3596
rect 1895 3576 1901 3596
rect 1905 3576 1907 3596
rect 1919 3576 1921 3596
rect 1735 3556 1748 3576
rect 1911 3556 1921 3576
rect 1925 3556 1927 3596
rect 1969 3556 1971 3596
rect 1975 3566 1977 3596
rect 1989 3566 1991 3596
rect 1975 3556 1991 3566
rect 1995 3556 1997 3596
rect 2009 3556 2011 3596
rect 2015 3584 2031 3596
rect 2015 3556 2017 3584
rect 2029 3556 2031 3584
rect 2035 3556 2037 3596
rect 2091 3556 2093 3596
rect 2097 3556 2103 3596
rect 2107 3556 2109 3596
rect 2190 3576 2192 3596
rect 2196 3576 2200 3596
rect 2212 3556 2214 3596
rect 2218 3556 2222 3596
rect 2226 3556 2228 3596
rect 2306 3538 2308 3596
rect 2294 3536 2308 3538
rect 2312 3536 2316 3596
rect 2320 3536 2324 3596
rect 2328 3536 2330 3596
rect 2383 3576 2385 3596
rect 2389 3576 2391 3596
rect 2466 3538 2468 3596
rect 2454 3536 2468 3538
rect 2472 3536 2476 3596
rect 2480 3536 2484 3596
rect 2488 3536 2490 3596
rect 2566 3538 2568 3596
rect 2554 3536 2568 3538
rect 2572 3536 2576 3596
rect 2580 3536 2584 3596
rect 2588 3536 2590 3596
rect 2643 3556 2645 3596
rect 2649 3556 2651 3596
rect 2663 3556 2665 3596
rect 2669 3568 2671 3596
rect 2683 3568 2685 3596
rect 2669 3556 2685 3568
rect 2689 3556 2691 3596
rect 2729 3556 2731 3596
rect 2735 3568 2737 3596
rect 2749 3568 2751 3596
rect 2735 3556 2751 3568
rect 2755 3556 2757 3596
rect 2769 3556 2771 3596
rect 2775 3556 2777 3596
rect 2831 3556 2833 3596
rect 2837 3556 2843 3596
rect 2847 3556 2849 3596
rect 2909 3556 2911 3596
rect 2915 3568 2917 3596
rect 2929 3568 2931 3596
rect 2915 3556 2931 3568
rect 2935 3556 2937 3596
rect 2949 3556 2951 3596
rect 2955 3556 2957 3596
rect 3009 3576 3011 3596
rect 3015 3576 3017 3596
rect 3029 3576 3031 3596
rect 3035 3576 3037 3596
rect 3103 3556 3105 3596
rect 3109 3556 3111 3596
rect 3123 3556 3125 3596
rect 3129 3568 3131 3596
rect 3143 3568 3145 3596
rect 3129 3556 3145 3568
rect 3149 3556 3151 3596
rect 3192 3556 3194 3596
rect 3198 3556 3202 3596
rect 3206 3556 3208 3596
rect 3220 3556 3222 3596
rect 3226 3556 3230 3596
rect 3234 3556 3236 3596
rect 3311 3556 3313 3596
rect 3317 3556 3323 3596
rect 3327 3556 3329 3596
rect 3391 3556 3393 3596
rect 3397 3556 3403 3596
rect 3407 3556 3409 3596
rect 3471 3556 3473 3596
rect 3477 3556 3483 3596
rect 3487 3556 3489 3596
rect 3549 3576 3551 3596
rect 3555 3576 3557 3596
rect 3569 3576 3571 3596
rect 3575 3576 3577 3596
rect 3631 3556 3633 3596
rect 3637 3556 3643 3596
rect 3647 3556 3649 3596
rect 3711 3556 3713 3596
rect 3717 3556 3723 3596
rect 3727 3556 3729 3596
rect 3811 3556 3813 3596
rect 3817 3556 3823 3596
rect 3827 3556 3829 3596
rect 3883 3576 3885 3596
rect 3889 3576 3891 3596
rect 3903 3576 3905 3596
rect 3909 3576 3911 3596
rect 3951 3556 3953 3596
rect 3957 3556 3963 3596
rect 3967 3556 3969 3596
rect 4031 3556 4033 3596
rect 4037 3556 4043 3596
rect 4047 3556 4049 3596
rect 4109 3556 4111 3596
rect 4115 3568 4117 3596
rect 4129 3568 4131 3596
rect 4115 3556 4131 3568
rect 4135 3556 4137 3596
rect 4149 3556 4151 3596
rect 4155 3556 4157 3596
rect 4246 3538 4248 3596
rect 4234 3536 4248 3538
rect 4252 3536 4256 3596
rect 4260 3536 4264 3596
rect 4268 3536 4270 3596
rect 4310 3536 4312 3596
rect 4316 3536 4320 3596
rect 4324 3536 4328 3596
rect 4332 3538 4334 3596
rect 4412 3556 4414 3596
rect 4418 3556 4422 3596
rect 4426 3556 4428 3596
rect 4440 3576 4444 3596
rect 4448 3576 4450 3596
rect 4509 3576 4511 3596
rect 4515 3576 4517 3596
rect 4332 3536 4346 3538
rect 4606 3538 4608 3596
rect 4594 3536 4608 3538
rect 4612 3536 4616 3596
rect 4620 3536 4624 3596
rect 4628 3536 4630 3596
rect 4670 3536 4672 3596
rect 4676 3536 4680 3596
rect 4684 3536 4688 3596
rect 4692 3538 4694 3596
rect 4692 3536 4706 3538
rect 33 3144 35 3184
rect 39 3164 49 3184
rect 212 3164 225 3184
rect 39 3144 41 3164
rect 53 3144 55 3164
rect 59 3144 65 3164
rect 69 3144 73 3164
rect 85 3144 87 3164
rect 91 3144 97 3164
rect 101 3144 103 3164
rect 115 3144 119 3164
rect 123 3144 125 3164
rect 163 3144 165 3164
rect 169 3144 173 3164
rect 177 3144 179 3164
rect 191 3144 193 3164
rect 197 3144 203 3164
rect 207 3144 209 3164
rect 221 3144 225 3164
rect 229 3144 231 3184
rect 304 3144 306 3184
rect 310 3144 314 3184
rect 318 3144 320 3184
rect 332 3144 334 3184
rect 338 3144 342 3184
rect 346 3144 348 3184
rect 391 3144 393 3184
rect 397 3144 403 3184
rect 407 3144 409 3184
rect 469 3144 471 3184
rect 475 3172 491 3184
rect 475 3144 477 3172
rect 489 3144 491 3172
rect 495 3144 497 3184
rect 509 3144 511 3184
rect 515 3144 517 3184
rect 569 3144 571 3184
rect 575 3172 591 3184
rect 575 3144 577 3172
rect 589 3144 591 3172
rect 595 3144 597 3184
rect 609 3144 611 3184
rect 615 3144 617 3184
rect 691 3144 693 3184
rect 697 3144 703 3184
rect 707 3144 709 3184
rect 749 3144 751 3164
rect 755 3144 757 3164
rect 823 3144 825 3184
rect 829 3144 831 3184
rect 843 3144 845 3184
rect 849 3144 851 3184
rect 863 3144 865 3184
rect 869 3144 871 3184
rect 883 3144 885 3184
rect 889 3144 891 3184
rect 903 3144 905 3184
rect 909 3144 911 3184
rect 923 3144 925 3184
rect 929 3144 931 3184
rect 943 3144 945 3184
rect 949 3144 951 3184
rect 963 3144 965 3184
rect 969 3144 971 3184
rect 1009 3144 1011 3184
rect 1015 3144 1017 3184
rect 1029 3144 1031 3184
rect 1035 3144 1037 3184
rect 1049 3144 1051 3184
rect 1055 3144 1057 3184
rect 1069 3144 1071 3184
rect 1075 3144 1077 3184
rect 1089 3144 1091 3184
rect 1095 3144 1097 3184
rect 1109 3144 1111 3184
rect 1115 3144 1117 3184
rect 1129 3144 1131 3184
rect 1135 3144 1137 3184
rect 1149 3144 1151 3184
rect 1155 3144 1157 3184
rect 1223 3144 1225 3164
rect 1229 3144 1231 3164
rect 1269 3144 1271 3184
rect 1275 3164 1288 3184
rect 1451 3164 1461 3184
rect 1275 3144 1279 3164
rect 1291 3144 1293 3164
rect 1297 3144 1303 3164
rect 1307 3144 1309 3164
rect 1321 3144 1323 3164
rect 1327 3144 1331 3164
rect 1335 3144 1337 3164
rect 1375 3144 1377 3164
rect 1381 3144 1385 3164
rect 1397 3144 1399 3164
rect 1403 3144 1409 3164
rect 1413 3144 1415 3164
rect 1427 3144 1431 3164
rect 1435 3144 1441 3164
rect 1445 3144 1447 3164
rect 1459 3144 1461 3164
rect 1465 3144 1467 3184
rect 1509 3144 1511 3184
rect 1515 3172 1531 3184
rect 1515 3144 1517 3172
rect 1529 3144 1531 3172
rect 1535 3144 1537 3184
rect 1549 3144 1551 3184
rect 1555 3144 1557 3184
rect 1623 3144 1625 3184
rect 1629 3144 1631 3184
rect 1643 3144 1645 3184
rect 1649 3172 1665 3184
rect 1649 3144 1651 3172
rect 1663 3144 1665 3172
rect 1669 3144 1671 3184
rect 1723 3144 1725 3184
rect 1729 3144 1731 3184
rect 1743 3144 1745 3184
rect 1749 3172 1765 3184
rect 1749 3144 1751 3172
rect 1763 3144 1765 3172
rect 1769 3144 1771 3184
rect 1823 3144 1825 3164
rect 1829 3144 1831 3164
rect 1883 3144 1885 3184
rect 1889 3144 1891 3184
rect 1903 3144 1905 3184
rect 1909 3172 1925 3184
rect 1909 3144 1911 3172
rect 1923 3144 1925 3172
rect 1929 3144 1931 3184
rect 1983 3144 1985 3184
rect 1989 3144 1991 3184
rect 2003 3144 2005 3184
rect 2009 3172 2025 3184
rect 2009 3144 2011 3172
rect 2023 3144 2025 3172
rect 2029 3144 2031 3184
rect 2069 3144 2071 3184
rect 2075 3164 2088 3184
rect 2251 3164 2261 3184
rect 2075 3144 2079 3164
rect 2091 3144 2093 3164
rect 2097 3144 2103 3164
rect 2107 3144 2109 3164
rect 2121 3144 2123 3164
rect 2127 3144 2131 3164
rect 2135 3144 2137 3164
rect 2175 3144 2177 3164
rect 2181 3144 2185 3164
rect 2197 3144 2199 3164
rect 2203 3144 2209 3164
rect 2213 3144 2215 3164
rect 2227 3144 2231 3164
rect 2235 3144 2241 3164
rect 2245 3144 2247 3164
rect 2259 3144 2261 3164
rect 2265 3144 2267 3184
rect 2454 3202 2468 3204
rect 2323 3144 2325 3164
rect 2329 3144 2331 3164
rect 2383 3144 2385 3164
rect 2389 3144 2391 3164
rect 2466 3144 2468 3202
rect 2472 3144 2476 3204
rect 2480 3144 2484 3204
rect 2488 3144 2490 3204
rect 2532 3144 2534 3184
rect 2538 3144 2542 3184
rect 2546 3144 2548 3184
rect 2560 3144 2564 3164
rect 2568 3144 2570 3164
rect 2643 3144 2645 3164
rect 2649 3144 2651 3164
rect 2703 3144 2705 3184
rect 2709 3144 2711 3184
rect 2723 3144 2725 3184
rect 2729 3172 2745 3184
rect 2729 3144 2731 3172
rect 2743 3144 2745 3172
rect 2749 3144 2751 3184
rect 2789 3144 2791 3164
rect 2795 3144 2797 3164
rect 2809 3144 2811 3164
rect 2815 3144 2817 3164
rect 2869 3144 2871 3184
rect 2875 3172 2891 3184
rect 2875 3144 2877 3172
rect 2889 3144 2891 3172
rect 2895 3144 2897 3184
rect 2909 3144 2911 3184
rect 2915 3144 2917 3184
rect 2971 3144 2973 3184
rect 2977 3144 2983 3184
rect 2987 3144 2989 3184
rect 3051 3144 3053 3184
rect 3057 3144 3063 3184
rect 3067 3144 3069 3184
rect 3254 3202 3268 3204
rect 3150 3144 3152 3164
rect 3156 3144 3160 3164
rect 3172 3144 3174 3184
rect 3178 3144 3182 3184
rect 3186 3144 3188 3184
rect 3266 3144 3268 3202
rect 3272 3144 3276 3204
rect 3280 3144 3284 3204
rect 3288 3144 3290 3204
rect 3343 3144 3345 3184
rect 3349 3144 3351 3184
rect 3363 3144 3365 3184
rect 3369 3172 3385 3184
rect 3369 3144 3371 3172
rect 3383 3144 3385 3172
rect 3389 3144 3391 3184
rect 3453 3144 3455 3184
rect 3459 3144 3461 3184
rect 3473 3144 3475 3184
rect 3479 3144 3485 3184
rect 3489 3144 3491 3184
rect 3531 3144 3533 3184
rect 3537 3144 3543 3184
rect 3547 3144 3549 3184
rect 3633 3144 3635 3184
rect 3639 3144 3641 3184
rect 3653 3144 3655 3184
rect 3659 3144 3665 3184
rect 3669 3144 3671 3184
rect 3744 3144 3746 3184
rect 3750 3144 3754 3184
rect 3758 3144 3760 3184
rect 3772 3144 3774 3184
rect 3778 3144 3782 3184
rect 3786 3144 3788 3184
rect 3851 3144 3853 3184
rect 3857 3144 3863 3184
rect 3867 3144 3869 3184
rect 3909 3144 3911 3184
rect 3915 3172 3931 3184
rect 3915 3144 3917 3172
rect 3929 3144 3931 3172
rect 3935 3144 3937 3184
rect 3949 3144 3951 3184
rect 3955 3144 3957 3184
rect 4011 3144 4013 3184
rect 4017 3144 4023 3184
rect 4027 3144 4029 3184
rect 4113 3144 4115 3184
rect 4119 3144 4121 3184
rect 4133 3144 4135 3184
rect 4139 3144 4145 3184
rect 4149 3144 4151 3184
rect 4191 3144 4193 3184
rect 4197 3144 4203 3184
rect 4207 3144 4209 3184
rect 4269 3144 4271 3184
rect 4275 3144 4281 3184
rect 4285 3144 4287 3184
rect 4299 3144 4301 3184
rect 4305 3144 4307 3184
rect 4372 3144 4374 3184
rect 4378 3144 4382 3184
rect 4386 3144 4388 3184
rect 4694 3202 4708 3204
rect 4400 3144 4404 3164
rect 4408 3144 4410 3164
rect 4469 3144 4471 3184
rect 4475 3172 4491 3184
rect 4475 3144 4477 3172
rect 4489 3144 4491 3172
rect 4495 3144 4497 3184
rect 4509 3144 4511 3184
rect 4515 3144 4517 3184
rect 4569 3144 4571 3184
rect 4575 3172 4591 3184
rect 4575 3144 4577 3172
rect 4589 3144 4591 3172
rect 4595 3144 4597 3184
rect 4609 3144 4611 3184
rect 4615 3144 4617 3184
rect 4706 3144 4708 3202
rect 4712 3144 4716 3204
rect 4720 3144 4724 3204
rect 4728 3144 4730 3204
rect 33 3076 35 3116
rect 39 3096 41 3116
rect 53 3096 55 3116
rect 59 3096 65 3116
rect 69 3096 73 3116
rect 85 3096 87 3116
rect 91 3096 97 3116
rect 101 3096 103 3116
rect 115 3096 119 3116
rect 123 3096 125 3116
rect 163 3096 165 3116
rect 169 3096 173 3116
rect 177 3096 179 3116
rect 191 3096 193 3116
rect 197 3096 203 3116
rect 207 3096 209 3116
rect 221 3096 225 3116
rect 39 3076 49 3096
rect 212 3076 225 3096
rect 229 3076 231 3116
rect 283 3076 285 3116
rect 289 3076 291 3116
rect 303 3076 305 3116
rect 309 3088 311 3116
rect 323 3088 325 3116
rect 309 3076 325 3088
rect 329 3076 331 3116
rect 391 3076 393 3116
rect 397 3076 403 3116
rect 407 3076 409 3116
rect 449 3076 451 3116
rect 455 3096 459 3116
rect 471 3096 473 3116
rect 477 3096 483 3116
rect 487 3096 489 3116
rect 501 3096 503 3116
rect 507 3096 511 3116
rect 515 3096 517 3116
rect 555 3096 557 3116
rect 561 3096 565 3116
rect 577 3096 579 3116
rect 583 3096 589 3116
rect 593 3096 595 3116
rect 607 3096 611 3116
rect 615 3096 621 3116
rect 625 3096 627 3116
rect 639 3096 641 3116
rect 455 3076 468 3096
rect 631 3076 641 3096
rect 645 3076 647 3116
rect 693 3076 695 3116
rect 699 3096 701 3116
rect 713 3096 715 3116
rect 719 3096 725 3116
rect 729 3096 733 3116
rect 745 3096 747 3116
rect 751 3096 757 3116
rect 761 3096 763 3116
rect 775 3096 779 3116
rect 783 3096 785 3116
rect 823 3096 825 3116
rect 829 3096 833 3116
rect 837 3096 839 3116
rect 851 3096 853 3116
rect 857 3096 863 3116
rect 867 3096 869 3116
rect 881 3096 885 3116
rect 699 3076 709 3096
rect 872 3076 885 3096
rect 889 3076 891 3116
rect 929 3096 931 3116
rect 935 3096 937 3116
rect 1003 3096 1005 3116
rect 1009 3096 1011 3116
rect 1023 3096 1025 3116
rect 1029 3096 1031 3116
rect 1091 3076 1093 3116
rect 1097 3076 1103 3116
rect 1107 3076 1109 3116
rect 1149 3076 1151 3116
rect 1155 3088 1157 3116
rect 1169 3088 1171 3116
rect 1155 3076 1171 3088
rect 1175 3076 1177 3116
rect 1189 3076 1191 3116
rect 1195 3076 1197 3116
rect 1252 3076 1254 3116
rect 1258 3076 1262 3116
rect 1266 3076 1268 3116
rect 1280 3096 1284 3116
rect 1288 3096 1290 3116
rect 1353 3076 1355 3116
rect 1359 3096 1361 3116
rect 1373 3096 1375 3116
rect 1379 3096 1385 3116
rect 1389 3096 1393 3116
rect 1405 3096 1407 3116
rect 1411 3096 1417 3116
rect 1421 3096 1423 3116
rect 1435 3096 1439 3116
rect 1443 3096 1445 3116
rect 1483 3096 1485 3116
rect 1489 3096 1493 3116
rect 1497 3096 1499 3116
rect 1511 3096 1513 3116
rect 1517 3096 1523 3116
rect 1527 3096 1529 3116
rect 1541 3096 1545 3116
rect 1359 3076 1369 3096
rect 1532 3076 1545 3096
rect 1549 3076 1551 3116
rect 1603 3096 1605 3116
rect 1609 3096 1611 3116
rect 1623 3096 1625 3116
rect 1629 3096 1631 3116
rect 1691 3076 1693 3116
rect 1697 3076 1703 3116
rect 1707 3076 1709 3116
rect 1749 3076 1751 3116
rect 1755 3088 1757 3116
rect 1769 3088 1771 3116
rect 1755 3076 1771 3088
rect 1775 3076 1777 3116
rect 1789 3076 1791 3116
rect 1795 3076 1797 3116
rect 1863 3076 1865 3116
rect 1869 3076 1871 3116
rect 1883 3076 1885 3116
rect 1889 3088 1891 3116
rect 1903 3088 1905 3116
rect 1889 3076 1905 3088
rect 1909 3076 1911 3116
rect 1949 3076 1951 3116
rect 1955 3096 1959 3116
rect 1971 3096 1973 3116
rect 1977 3096 1983 3116
rect 1987 3096 1989 3116
rect 2001 3096 2003 3116
rect 2007 3096 2011 3116
rect 2015 3096 2017 3116
rect 2055 3096 2057 3116
rect 2061 3096 2065 3116
rect 2077 3096 2079 3116
rect 2083 3096 2089 3116
rect 2093 3096 2095 3116
rect 2107 3096 2111 3116
rect 2115 3096 2121 3116
rect 2125 3096 2127 3116
rect 2139 3096 2141 3116
rect 1955 3076 1968 3096
rect 2131 3076 2141 3096
rect 2145 3076 2147 3116
rect 2203 3096 2205 3116
rect 2209 3096 2211 3116
rect 2223 3096 2225 3116
rect 2229 3096 2231 3116
rect 2283 3096 2285 3116
rect 2289 3096 2291 3116
rect 2366 3058 2368 3116
rect 2354 3056 2368 3058
rect 2372 3056 2376 3116
rect 2380 3056 2384 3116
rect 2388 3056 2390 3116
rect 2450 3096 2452 3116
rect 2456 3096 2460 3116
rect 2472 3076 2474 3116
rect 2478 3076 2482 3116
rect 2486 3076 2488 3116
rect 2566 3058 2568 3116
rect 2554 3056 2568 3058
rect 2572 3056 2576 3116
rect 2580 3056 2584 3116
rect 2588 3056 2590 3116
rect 2643 3076 2645 3116
rect 2649 3076 2651 3116
rect 2663 3076 2665 3116
rect 2669 3088 2671 3116
rect 2683 3088 2685 3116
rect 2669 3076 2685 3088
rect 2689 3076 2691 3116
rect 2743 3096 2745 3116
rect 2749 3096 2751 3116
rect 2763 3096 2765 3116
rect 2769 3096 2771 3116
rect 2811 3076 2813 3116
rect 2817 3076 2823 3116
rect 2827 3076 2829 3116
rect 2891 3076 2893 3116
rect 2897 3076 2903 3116
rect 2907 3076 2909 3116
rect 2972 3076 2974 3116
rect 2978 3076 2982 3116
rect 2986 3076 2988 3116
rect 3000 3076 3002 3116
rect 3006 3076 3010 3116
rect 3014 3076 3016 3116
rect 3091 3076 3093 3116
rect 3097 3076 3103 3116
rect 3107 3076 3109 3116
rect 3169 3076 3171 3116
rect 3175 3088 3177 3116
rect 3189 3088 3191 3116
rect 3175 3076 3191 3088
rect 3195 3076 3197 3116
rect 3209 3076 3211 3116
rect 3215 3076 3217 3116
rect 3269 3076 3271 3116
rect 3275 3076 3277 3116
rect 3329 3076 3331 3116
rect 3335 3076 3341 3116
rect 3345 3076 3347 3116
rect 3359 3076 3361 3116
rect 3365 3076 3367 3116
rect 3441 3076 3443 3116
rect 3447 3076 3449 3116
rect 3461 3096 3465 3116
rect 3469 3096 3471 3116
rect 3521 3076 3523 3116
rect 3527 3076 3529 3116
rect 3541 3096 3545 3116
rect 3549 3096 3551 3116
rect 3591 3076 3593 3116
rect 3597 3076 3603 3116
rect 3607 3076 3609 3116
rect 3669 3076 3671 3116
rect 3675 3088 3677 3116
rect 3689 3088 3691 3116
rect 3675 3076 3691 3088
rect 3695 3076 3697 3116
rect 3709 3076 3711 3116
rect 3715 3076 3717 3116
rect 3781 3076 3783 3116
rect 3787 3076 3789 3116
rect 3801 3096 3805 3116
rect 3809 3096 3811 3116
rect 3849 3076 3851 3116
rect 3855 3088 3857 3116
rect 3869 3088 3871 3116
rect 3855 3076 3871 3088
rect 3875 3076 3877 3116
rect 3889 3076 3891 3116
rect 3895 3076 3897 3116
rect 3950 3056 3952 3116
rect 3956 3056 3960 3116
rect 3964 3056 3968 3116
rect 3972 3058 3974 3116
rect 4049 3096 4051 3116
rect 4055 3096 4059 3116
rect 3972 3056 3986 3058
rect 4071 3076 4073 3116
rect 4077 3076 4079 3116
rect 4150 3096 4152 3116
rect 4156 3096 4160 3116
rect 4172 3076 4174 3116
rect 4178 3076 4182 3116
rect 4186 3076 4188 3116
rect 4230 3056 4232 3116
rect 4236 3056 4240 3116
rect 4244 3056 4248 3116
rect 4252 3058 4254 3116
rect 4350 3096 4352 3116
rect 4356 3096 4360 3116
rect 4252 3056 4266 3058
rect 4372 3076 4374 3116
rect 4378 3076 4382 3116
rect 4386 3076 4388 3116
rect 4466 3058 4468 3116
rect 4454 3056 4468 3058
rect 4472 3056 4476 3116
rect 4480 3056 4484 3116
rect 4488 3056 4490 3116
rect 4543 3096 4545 3116
rect 4549 3096 4551 3116
rect 4603 3076 4605 3116
rect 4609 3076 4611 3116
rect 4623 3076 4625 3116
rect 4629 3088 4631 3116
rect 4643 3088 4645 3116
rect 4629 3076 4645 3088
rect 4649 3076 4651 3116
rect 4689 3076 4691 3116
rect 4695 3088 4697 3116
rect 4709 3088 4711 3116
rect 4695 3076 4711 3088
rect 4715 3076 4717 3116
rect 4729 3076 4731 3116
rect 4735 3076 4737 3116
rect 33 2664 35 2704
rect 39 2684 49 2704
rect 212 2684 225 2704
rect 39 2664 41 2684
rect 53 2664 55 2684
rect 59 2664 65 2684
rect 69 2664 73 2684
rect 85 2664 87 2684
rect 91 2664 97 2684
rect 101 2664 103 2684
rect 115 2664 119 2684
rect 123 2664 125 2684
rect 163 2664 165 2684
rect 169 2664 173 2684
rect 177 2664 179 2684
rect 191 2664 193 2684
rect 197 2664 203 2684
rect 207 2664 209 2684
rect 221 2664 225 2684
rect 229 2664 231 2704
rect 304 2664 306 2704
rect 310 2664 314 2704
rect 318 2664 320 2704
rect 332 2664 334 2704
rect 338 2664 342 2704
rect 346 2664 348 2704
rect 391 2664 393 2704
rect 397 2664 403 2704
rect 407 2664 409 2704
rect 483 2664 485 2704
rect 489 2664 491 2704
rect 503 2664 505 2704
rect 509 2692 525 2704
rect 509 2664 511 2692
rect 523 2664 525 2692
rect 529 2664 531 2704
rect 581 2664 583 2704
rect 587 2664 589 2704
rect 601 2664 605 2684
rect 609 2664 611 2684
rect 651 2664 653 2704
rect 657 2664 663 2704
rect 667 2664 669 2704
rect 743 2664 745 2704
rect 749 2664 751 2704
rect 763 2664 765 2704
rect 769 2692 785 2704
rect 769 2664 771 2692
rect 783 2664 785 2692
rect 789 2664 791 2704
rect 843 2664 845 2684
rect 849 2664 851 2684
rect 863 2664 865 2684
rect 869 2664 871 2684
rect 931 2664 933 2704
rect 937 2664 943 2704
rect 947 2664 949 2704
rect 989 2664 991 2684
rect 995 2664 997 2684
rect 1071 2664 1073 2704
rect 1077 2664 1083 2704
rect 1087 2664 1089 2704
rect 1129 2664 1131 2684
rect 1135 2664 1137 2684
rect 1149 2664 1151 2684
rect 1155 2664 1157 2684
rect 1221 2664 1223 2704
rect 1227 2664 1229 2704
rect 1241 2664 1245 2684
rect 1249 2664 1251 2684
rect 1293 2664 1295 2704
rect 1299 2684 1309 2704
rect 1472 2684 1485 2704
rect 1299 2664 1301 2684
rect 1313 2664 1315 2684
rect 1319 2664 1325 2684
rect 1329 2664 1333 2684
rect 1345 2664 1347 2684
rect 1351 2664 1357 2684
rect 1361 2664 1363 2684
rect 1375 2664 1379 2684
rect 1383 2664 1385 2684
rect 1423 2664 1425 2684
rect 1429 2664 1433 2684
rect 1437 2664 1439 2684
rect 1451 2664 1453 2684
rect 1457 2664 1463 2684
rect 1467 2664 1469 2684
rect 1481 2664 1485 2684
rect 1489 2664 1491 2704
rect 1531 2664 1533 2704
rect 1537 2664 1543 2704
rect 1547 2664 1549 2704
rect 1623 2664 1625 2704
rect 1629 2664 1631 2704
rect 1643 2664 1645 2704
rect 1649 2692 1665 2704
rect 1649 2664 1651 2692
rect 1663 2664 1665 2692
rect 1669 2664 1671 2704
rect 1723 2664 1725 2704
rect 1729 2664 1731 2704
rect 1743 2664 1745 2704
rect 1749 2692 1765 2704
rect 1749 2664 1751 2692
rect 1763 2664 1765 2692
rect 1769 2664 1771 2704
rect 1823 2664 1825 2684
rect 1829 2664 1831 2684
rect 1843 2664 1845 2684
rect 1849 2664 1851 2684
rect 1910 2664 1912 2684
rect 1916 2664 1920 2684
rect 1932 2664 1934 2704
rect 1938 2664 1942 2704
rect 1946 2664 1948 2704
rect 2001 2664 2003 2704
rect 2007 2664 2009 2704
rect 2094 2722 2108 2724
rect 2021 2664 2025 2684
rect 2029 2664 2031 2684
rect 2106 2664 2108 2722
rect 2112 2664 2116 2724
rect 2120 2664 2124 2724
rect 2128 2664 2130 2724
rect 2169 2664 2171 2684
rect 2175 2664 2179 2684
rect 2191 2664 2193 2704
rect 2197 2664 2199 2704
rect 2253 2664 2255 2704
rect 2259 2684 2269 2704
rect 2432 2684 2445 2704
rect 2259 2664 2261 2684
rect 2273 2664 2275 2684
rect 2279 2664 2285 2684
rect 2289 2664 2293 2684
rect 2305 2664 2307 2684
rect 2311 2664 2317 2684
rect 2321 2664 2323 2684
rect 2335 2664 2339 2684
rect 2343 2664 2345 2684
rect 2383 2664 2385 2684
rect 2389 2664 2393 2684
rect 2397 2664 2399 2684
rect 2411 2664 2413 2684
rect 2417 2664 2423 2684
rect 2427 2664 2429 2684
rect 2441 2664 2445 2684
rect 2449 2664 2451 2704
rect 2503 2664 2505 2704
rect 2509 2664 2511 2704
rect 2523 2664 2525 2704
rect 2529 2692 2545 2704
rect 2529 2664 2531 2692
rect 2543 2664 2545 2692
rect 2549 2664 2551 2704
rect 2603 2664 2605 2704
rect 2609 2664 2611 2704
rect 2623 2664 2625 2704
rect 2629 2692 2645 2704
rect 2629 2664 2631 2692
rect 2643 2664 2645 2692
rect 2649 2664 2651 2704
rect 2689 2664 2691 2704
rect 2695 2692 2711 2704
rect 2695 2664 2697 2692
rect 2709 2664 2711 2692
rect 2715 2664 2717 2704
rect 2729 2664 2731 2704
rect 2735 2664 2737 2704
rect 2791 2664 2793 2704
rect 2797 2664 2803 2704
rect 2807 2664 2809 2704
rect 2871 2664 2873 2704
rect 2877 2664 2883 2704
rect 2887 2664 2889 2704
rect 2949 2664 2951 2704
rect 2955 2692 2971 2704
rect 2955 2664 2957 2692
rect 2969 2664 2971 2692
rect 2975 2664 2977 2704
rect 2989 2664 2991 2704
rect 2995 2664 2997 2704
rect 3049 2664 3051 2704
rect 3055 2692 3071 2704
rect 3055 2664 3057 2692
rect 3069 2664 3071 2692
rect 3075 2664 3077 2704
rect 3089 2664 3091 2704
rect 3095 2664 3097 2704
rect 3151 2664 3153 2704
rect 3157 2664 3163 2704
rect 3167 2664 3169 2704
rect 3243 2664 3245 2704
rect 3249 2664 3251 2704
rect 3263 2664 3265 2704
rect 3269 2692 3285 2704
rect 3269 2664 3271 2692
rect 3283 2664 3285 2692
rect 3289 2664 3291 2704
rect 3351 2664 3353 2704
rect 3357 2664 3363 2704
rect 3367 2664 3369 2704
rect 3410 2664 3412 2724
rect 3416 2664 3420 2724
rect 3424 2664 3428 2724
rect 3432 2722 3446 2724
rect 3432 2664 3434 2722
rect 3523 2664 3525 2704
rect 3529 2664 3531 2704
rect 3543 2664 3545 2704
rect 3549 2692 3565 2704
rect 3549 2664 3551 2692
rect 3563 2664 3565 2692
rect 3569 2664 3571 2704
rect 3609 2664 3611 2704
rect 3615 2692 3631 2704
rect 3615 2664 3617 2692
rect 3629 2664 3631 2692
rect 3635 2664 3637 2704
rect 3649 2664 3651 2704
rect 3655 2664 3657 2704
rect 3731 2664 3733 2704
rect 3737 2664 3743 2704
rect 3747 2664 3749 2704
rect 3803 2664 3805 2704
rect 3809 2664 3811 2704
rect 3823 2664 3825 2704
rect 3829 2692 3845 2704
rect 3829 2664 3831 2692
rect 3843 2664 3845 2692
rect 3849 2664 3851 2704
rect 3890 2664 3892 2724
rect 3896 2664 3900 2724
rect 3904 2664 3908 2724
rect 3912 2722 3926 2724
rect 3912 2664 3914 2722
rect 3989 2664 3991 2684
rect 3995 2664 3997 2684
rect 4084 2664 4086 2704
rect 4090 2664 4094 2704
rect 4098 2664 4100 2704
rect 4112 2664 4114 2704
rect 4118 2664 4122 2704
rect 4126 2664 4128 2704
rect 4170 2664 4172 2724
rect 4176 2664 4180 2724
rect 4184 2664 4188 2724
rect 4192 2722 4206 2724
rect 4192 2664 4194 2722
rect 4269 2664 4271 2704
rect 4275 2692 4291 2704
rect 4275 2664 4277 2692
rect 4289 2664 4291 2692
rect 4295 2664 4297 2704
rect 4309 2664 4311 2704
rect 4315 2664 4317 2704
rect 4369 2664 4371 2704
rect 4375 2664 4381 2704
rect 4385 2664 4387 2704
rect 4399 2664 4401 2704
rect 4405 2664 4407 2704
rect 4472 2664 4474 2704
rect 4478 2664 4482 2704
rect 4486 2664 4488 2704
rect 4500 2664 4502 2704
rect 4506 2664 4510 2704
rect 4514 2664 4516 2704
rect 4589 2664 4591 2684
rect 4595 2664 4597 2684
rect 4652 2664 4654 2704
rect 4658 2664 4662 2704
rect 4666 2664 4668 2704
rect 4680 2664 4684 2684
rect 4688 2664 4690 2684
rect 33 2596 35 2636
rect 39 2616 41 2636
rect 53 2616 55 2636
rect 59 2616 65 2636
rect 69 2616 73 2636
rect 85 2616 87 2636
rect 91 2616 97 2636
rect 101 2616 103 2636
rect 115 2616 119 2636
rect 123 2616 125 2636
rect 163 2616 165 2636
rect 169 2616 173 2636
rect 177 2616 179 2636
rect 191 2616 193 2636
rect 197 2616 203 2636
rect 207 2616 209 2636
rect 221 2616 225 2636
rect 39 2596 49 2616
rect 212 2596 225 2616
rect 229 2596 231 2636
rect 283 2596 285 2636
rect 289 2596 291 2636
rect 303 2596 305 2636
rect 309 2608 311 2636
rect 323 2608 325 2636
rect 309 2596 325 2608
rect 329 2596 331 2636
rect 369 2616 371 2636
rect 375 2616 379 2636
rect 391 2596 393 2636
rect 397 2596 399 2636
rect 451 2596 453 2636
rect 457 2596 463 2636
rect 467 2596 469 2636
rect 543 2596 545 2636
rect 549 2596 551 2636
rect 563 2596 565 2636
rect 569 2608 571 2636
rect 583 2608 585 2636
rect 569 2596 585 2608
rect 589 2596 591 2636
rect 629 2616 631 2636
rect 635 2616 639 2636
rect 651 2596 653 2636
rect 657 2596 659 2636
rect 723 2596 725 2636
rect 729 2596 731 2636
rect 743 2596 745 2636
rect 749 2608 751 2636
rect 763 2608 765 2636
rect 749 2596 765 2608
rect 769 2596 771 2636
rect 809 2616 811 2636
rect 815 2616 817 2636
rect 829 2616 831 2636
rect 835 2616 837 2636
rect 893 2596 895 2636
rect 899 2616 901 2636
rect 913 2616 915 2636
rect 919 2616 925 2636
rect 929 2616 933 2636
rect 945 2616 947 2636
rect 951 2616 957 2636
rect 961 2616 963 2636
rect 975 2616 979 2636
rect 983 2616 985 2636
rect 1023 2616 1025 2636
rect 1029 2616 1033 2636
rect 1037 2616 1039 2636
rect 1051 2616 1053 2636
rect 1057 2616 1063 2636
rect 1067 2616 1069 2636
rect 1081 2616 1085 2636
rect 899 2596 909 2616
rect 1072 2596 1085 2616
rect 1089 2596 1091 2636
rect 1129 2616 1131 2636
rect 1135 2616 1137 2636
rect 1189 2596 1191 2636
rect 1195 2608 1197 2636
rect 1209 2608 1211 2636
rect 1195 2596 1211 2608
rect 1215 2596 1217 2636
rect 1229 2596 1231 2636
rect 1235 2596 1237 2636
rect 1289 2616 1291 2636
rect 1295 2616 1297 2636
rect 1351 2596 1353 2636
rect 1357 2596 1363 2636
rect 1367 2596 1369 2636
rect 1429 2596 1431 2636
rect 1435 2616 1439 2636
rect 1451 2616 1453 2636
rect 1457 2616 1463 2636
rect 1467 2616 1469 2636
rect 1481 2616 1483 2636
rect 1487 2616 1491 2636
rect 1495 2616 1497 2636
rect 1535 2616 1537 2636
rect 1541 2616 1545 2636
rect 1557 2616 1559 2636
rect 1563 2616 1569 2636
rect 1573 2616 1575 2636
rect 1587 2616 1591 2636
rect 1595 2616 1601 2636
rect 1605 2616 1607 2636
rect 1619 2616 1621 2636
rect 1435 2596 1448 2616
rect 1611 2596 1621 2616
rect 1625 2596 1627 2636
rect 1669 2596 1671 2636
rect 1675 2608 1677 2636
rect 1689 2608 1691 2636
rect 1675 2596 1691 2608
rect 1695 2596 1697 2636
rect 1709 2596 1711 2636
rect 1715 2596 1717 2636
rect 1769 2596 1771 2636
rect 1775 2616 1779 2636
rect 1791 2616 1793 2636
rect 1797 2616 1803 2636
rect 1807 2616 1809 2636
rect 1821 2616 1823 2636
rect 1827 2616 1831 2636
rect 1835 2616 1837 2636
rect 1875 2616 1877 2636
rect 1881 2616 1885 2636
rect 1897 2616 1899 2636
rect 1903 2616 1909 2636
rect 1913 2616 1915 2636
rect 1927 2616 1931 2636
rect 1935 2616 1941 2636
rect 1945 2616 1947 2636
rect 1959 2616 1961 2636
rect 1775 2596 1788 2616
rect 1951 2596 1961 2616
rect 1965 2596 1967 2636
rect 2009 2596 2011 2636
rect 2015 2596 2017 2636
rect 2029 2596 2031 2636
rect 2035 2596 2037 2636
rect 2049 2596 2051 2636
rect 2055 2596 2057 2636
rect 2069 2596 2071 2636
rect 2075 2596 2077 2636
rect 2089 2596 2091 2636
rect 2095 2596 2097 2636
rect 2109 2596 2111 2636
rect 2115 2596 2117 2636
rect 2129 2596 2131 2636
rect 2135 2596 2137 2636
rect 2149 2596 2151 2636
rect 2155 2596 2157 2636
rect 2213 2596 2215 2636
rect 2219 2616 2221 2636
rect 2233 2616 2235 2636
rect 2239 2616 2245 2636
rect 2249 2616 2253 2636
rect 2265 2616 2267 2636
rect 2271 2616 2277 2636
rect 2281 2616 2283 2636
rect 2295 2616 2299 2636
rect 2303 2616 2305 2636
rect 2343 2616 2345 2636
rect 2349 2616 2353 2636
rect 2357 2616 2359 2636
rect 2371 2616 2373 2636
rect 2377 2616 2383 2636
rect 2387 2616 2389 2636
rect 2401 2616 2405 2636
rect 2219 2596 2229 2616
rect 2392 2596 2405 2616
rect 2409 2596 2411 2636
rect 2471 2596 2473 2636
rect 2477 2596 2483 2636
rect 2487 2596 2489 2636
rect 2529 2616 2531 2636
rect 2535 2616 2537 2636
rect 2603 2596 2605 2636
rect 2609 2596 2611 2636
rect 2623 2596 2625 2636
rect 2629 2608 2631 2636
rect 2643 2608 2645 2636
rect 2629 2596 2645 2608
rect 2649 2596 2651 2636
rect 2689 2616 2691 2636
rect 2695 2616 2697 2636
rect 2771 2596 2773 2636
rect 2777 2596 2783 2636
rect 2787 2596 2789 2636
rect 2843 2596 2845 2636
rect 2849 2596 2851 2636
rect 2863 2596 2865 2636
rect 2869 2608 2871 2636
rect 2883 2608 2885 2636
rect 2869 2596 2885 2608
rect 2889 2596 2891 2636
rect 2929 2596 2931 2636
rect 2935 2596 2941 2636
rect 2945 2596 2947 2636
rect 2959 2596 2961 2636
rect 2965 2596 2967 2636
rect 3029 2596 3031 2636
rect 3035 2608 3037 2636
rect 3049 2608 3051 2636
rect 3035 2596 3051 2608
rect 3055 2596 3057 2636
rect 3069 2596 3071 2636
rect 3075 2596 3077 2636
rect 3151 2596 3153 2636
rect 3157 2596 3163 2636
rect 3167 2596 3169 2636
rect 3209 2596 3211 2636
rect 3215 2596 3221 2636
rect 3225 2596 3227 2636
rect 3239 2596 3241 2636
rect 3245 2596 3247 2636
rect 3346 2578 3348 2636
rect 3334 2576 3348 2578
rect 3352 2576 3356 2636
rect 3360 2576 3364 2636
rect 3368 2576 3370 2636
rect 3409 2616 3411 2636
rect 3415 2616 3417 2636
rect 3471 2596 3473 2636
rect 3477 2596 3483 2636
rect 3487 2596 3489 2636
rect 3549 2596 3551 2636
rect 3555 2596 3561 2636
rect 3565 2596 3567 2636
rect 3579 2596 3581 2636
rect 3585 2596 3587 2636
rect 3649 2616 3651 2636
rect 3655 2616 3659 2636
rect 3671 2596 3673 2636
rect 3677 2596 3679 2636
rect 3729 2616 3731 2636
rect 3735 2616 3737 2636
rect 3813 2596 3815 2636
rect 3819 2596 3821 2636
rect 3833 2596 3835 2636
rect 3839 2596 3845 2636
rect 3849 2596 3851 2636
rect 3924 2596 3926 2636
rect 3930 2596 3934 2636
rect 3938 2596 3940 2636
rect 3952 2596 3954 2636
rect 3958 2596 3962 2636
rect 3966 2596 3968 2636
rect 4031 2596 4033 2636
rect 4037 2596 4043 2636
rect 4047 2596 4049 2636
rect 4111 2596 4113 2636
rect 4117 2596 4123 2636
rect 4127 2596 4129 2636
rect 4169 2596 4171 2636
rect 4175 2608 4177 2636
rect 4189 2608 4191 2636
rect 4175 2596 4191 2608
rect 4195 2596 4197 2636
rect 4209 2596 4211 2636
rect 4215 2596 4217 2636
rect 4271 2596 4273 2636
rect 4277 2596 4283 2636
rect 4287 2596 4289 2636
rect 4386 2578 4388 2636
rect 4374 2576 4388 2578
rect 4392 2576 4396 2636
rect 4400 2576 4404 2636
rect 4408 2576 4410 2636
rect 4486 2578 4488 2636
rect 4474 2576 4488 2578
rect 4492 2576 4496 2636
rect 4500 2576 4504 2636
rect 4508 2576 4510 2636
rect 4552 2596 4554 2636
rect 4558 2596 4562 2636
rect 4566 2596 4568 2636
rect 4580 2616 4584 2636
rect 4588 2616 4590 2636
rect 4686 2578 4688 2636
rect 4674 2576 4688 2578
rect 4692 2576 4696 2636
rect 4700 2576 4704 2636
rect 4708 2576 4710 2636
rect 33 2184 35 2224
rect 39 2204 49 2224
rect 212 2204 225 2224
rect 39 2184 41 2204
rect 53 2184 55 2204
rect 59 2184 65 2204
rect 69 2184 73 2204
rect 85 2184 87 2204
rect 91 2184 97 2204
rect 101 2184 103 2204
rect 115 2184 119 2204
rect 123 2184 125 2204
rect 163 2184 165 2204
rect 169 2184 173 2204
rect 177 2184 179 2204
rect 191 2184 193 2204
rect 197 2184 203 2204
rect 207 2184 209 2204
rect 221 2184 225 2204
rect 229 2184 231 2224
rect 269 2184 271 2224
rect 275 2212 291 2224
rect 275 2184 277 2212
rect 289 2184 291 2212
rect 295 2184 297 2224
rect 309 2184 311 2224
rect 315 2184 317 2224
rect 372 2184 374 2224
rect 378 2184 382 2224
rect 386 2184 388 2224
rect 400 2184 402 2224
rect 406 2184 410 2224
rect 414 2184 416 2224
rect 489 2184 491 2204
rect 495 2184 499 2204
rect 511 2184 513 2224
rect 517 2184 519 2224
rect 571 2184 573 2224
rect 577 2184 583 2224
rect 587 2184 589 2224
rect 663 2184 665 2204
rect 669 2184 671 2204
rect 709 2184 711 2204
rect 715 2184 717 2204
rect 729 2184 731 2204
rect 735 2184 737 2204
rect 810 2184 812 2204
rect 816 2184 820 2204
rect 832 2184 834 2224
rect 838 2184 842 2224
rect 846 2184 848 2224
rect 889 2184 891 2204
rect 895 2184 897 2204
rect 909 2184 911 2204
rect 915 2184 917 2204
rect 969 2184 971 2204
rect 975 2184 977 2204
rect 989 2184 991 2204
rect 995 2184 997 2204
rect 1049 2184 1051 2204
rect 1055 2184 1057 2204
rect 1109 2184 1111 2224
rect 1115 2204 1128 2224
rect 1291 2204 1301 2224
rect 1115 2184 1119 2204
rect 1131 2184 1133 2204
rect 1137 2184 1143 2204
rect 1147 2184 1149 2204
rect 1161 2184 1163 2204
rect 1167 2184 1171 2204
rect 1175 2184 1177 2204
rect 1215 2184 1217 2204
rect 1221 2184 1225 2204
rect 1237 2184 1239 2204
rect 1243 2184 1249 2204
rect 1253 2184 1255 2204
rect 1267 2184 1271 2204
rect 1275 2184 1281 2204
rect 1285 2184 1287 2204
rect 1299 2184 1301 2204
rect 1305 2184 1307 2224
rect 1349 2184 1351 2224
rect 1355 2212 1371 2224
rect 1355 2184 1357 2212
rect 1369 2184 1371 2212
rect 1375 2184 1377 2224
rect 1389 2184 1391 2224
rect 1395 2184 1397 2224
rect 1449 2184 1451 2224
rect 1455 2204 1468 2224
rect 1631 2204 1641 2224
rect 1455 2184 1459 2204
rect 1471 2184 1473 2204
rect 1477 2184 1483 2204
rect 1487 2184 1489 2204
rect 1501 2184 1503 2204
rect 1507 2184 1511 2204
rect 1515 2184 1517 2204
rect 1555 2184 1557 2204
rect 1561 2184 1565 2204
rect 1577 2184 1579 2204
rect 1583 2184 1589 2204
rect 1593 2184 1595 2204
rect 1607 2184 1611 2204
rect 1615 2184 1621 2204
rect 1625 2184 1627 2204
rect 1639 2184 1641 2204
rect 1645 2184 1647 2224
rect 1703 2184 1705 2204
rect 1709 2184 1711 2204
rect 1723 2184 1725 2204
rect 1729 2184 1731 2204
rect 1790 2184 1792 2204
rect 1796 2184 1800 2204
rect 1812 2184 1814 2224
rect 1818 2184 1822 2224
rect 1826 2184 1828 2224
rect 1869 2184 1871 2224
rect 1875 2184 1877 2224
rect 1943 2184 1945 2204
rect 1949 2184 1951 2204
rect 1963 2184 1965 2204
rect 1969 2184 1971 2204
rect 2009 2184 2011 2224
rect 2015 2184 2017 2224
rect 2029 2184 2031 2224
rect 2035 2184 2037 2224
rect 2049 2184 2051 2224
rect 2055 2184 2057 2224
rect 2069 2184 2071 2224
rect 2075 2184 2077 2224
rect 2089 2184 2091 2224
rect 2095 2184 2097 2224
rect 2109 2184 2111 2224
rect 2115 2184 2117 2224
rect 2129 2184 2131 2224
rect 2135 2184 2137 2224
rect 2149 2184 2151 2224
rect 2155 2184 2157 2224
rect 2209 2184 2211 2224
rect 2215 2212 2231 2224
rect 2215 2184 2217 2212
rect 2229 2184 2231 2212
rect 2235 2184 2237 2224
rect 2249 2184 2251 2224
rect 2255 2184 2257 2224
rect 2313 2184 2315 2224
rect 2319 2204 2329 2224
rect 2492 2204 2505 2224
rect 2319 2184 2321 2204
rect 2333 2184 2335 2204
rect 2339 2184 2345 2204
rect 2349 2184 2353 2204
rect 2365 2184 2367 2204
rect 2371 2184 2377 2204
rect 2381 2184 2383 2204
rect 2395 2184 2399 2204
rect 2403 2184 2405 2204
rect 2443 2184 2445 2204
rect 2449 2184 2453 2204
rect 2457 2184 2459 2204
rect 2471 2184 2473 2204
rect 2477 2184 2483 2204
rect 2487 2184 2489 2204
rect 2501 2184 2505 2204
rect 2509 2184 2511 2224
rect 2571 2184 2573 2224
rect 2577 2184 2583 2224
rect 2587 2184 2589 2224
rect 2631 2184 2633 2224
rect 2637 2184 2643 2224
rect 2647 2184 2649 2224
rect 2711 2184 2713 2224
rect 2717 2184 2723 2224
rect 2727 2184 2729 2224
rect 2803 2184 2805 2224
rect 2809 2184 2811 2224
rect 2823 2184 2825 2224
rect 2829 2212 2845 2224
rect 2829 2184 2831 2212
rect 2843 2184 2845 2212
rect 2849 2184 2851 2224
rect 2903 2184 2905 2224
rect 2909 2184 2911 2224
rect 2923 2184 2925 2224
rect 2929 2212 2945 2224
rect 2929 2184 2931 2212
rect 2943 2184 2945 2212
rect 2949 2184 2951 2224
rect 2993 2184 2995 2224
rect 2999 2204 3009 2224
rect 3172 2204 3185 2224
rect 2999 2184 3001 2204
rect 3013 2184 3015 2204
rect 3019 2184 3025 2204
rect 3029 2184 3033 2204
rect 3045 2184 3047 2204
rect 3051 2184 3057 2204
rect 3061 2184 3063 2204
rect 3075 2184 3079 2204
rect 3083 2184 3085 2204
rect 3123 2184 3125 2204
rect 3129 2184 3133 2204
rect 3137 2184 3139 2204
rect 3151 2184 3153 2204
rect 3157 2184 3163 2204
rect 3167 2184 3169 2204
rect 3181 2184 3185 2204
rect 3189 2184 3191 2224
rect 3229 2184 3231 2224
rect 3235 2212 3251 2224
rect 3235 2184 3237 2212
rect 3249 2184 3251 2212
rect 3255 2184 3257 2224
rect 3269 2184 3271 2224
rect 3275 2184 3277 2224
rect 3331 2184 3333 2224
rect 3337 2184 3343 2224
rect 3347 2184 3349 2224
rect 3411 2184 3413 2224
rect 3417 2184 3423 2224
rect 3427 2184 3429 2224
rect 3511 2184 3513 2224
rect 3517 2184 3523 2224
rect 3527 2184 3529 2224
rect 3583 2184 3585 2224
rect 3589 2184 3591 2224
rect 3643 2184 3645 2224
rect 3649 2184 3651 2224
rect 3703 2184 3705 2204
rect 3709 2184 3711 2204
rect 3749 2184 3751 2224
rect 3755 2212 3771 2224
rect 3755 2184 3757 2212
rect 3769 2184 3771 2212
rect 3775 2184 3777 2224
rect 3789 2184 3791 2224
rect 3795 2184 3797 2224
rect 3861 2184 3863 2224
rect 3867 2184 3869 2224
rect 4214 2242 4228 2244
rect 3881 2184 3885 2204
rect 3889 2184 3891 2204
rect 3929 2184 3931 2224
rect 3935 2184 3937 2224
rect 3989 2184 3991 2224
rect 3995 2184 4001 2224
rect 4005 2184 4007 2224
rect 4019 2184 4021 2224
rect 4025 2184 4027 2224
rect 4103 2184 4105 2224
rect 4109 2184 4111 2224
rect 4123 2184 4125 2224
rect 4129 2212 4145 2224
rect 4129 2184 4131 2212
rect 4143 2184 4145 2212
rect 4149 2184 4151 2224
rect 4226 2184 4228 2242
rect 4232 2184 4236 2244
rect 4240 2184 4244 2244
rect 4248 2184 4250 2244
rect 4292 2184 4294 2224
rect 4298 2184 4302 2224
rect 4306 2184 4308 2224
rect 4320 2184 4324 2204
rect 4328 2184 4330 2204
rect 4403 2184 4405 2224
rect 4409 2184 4411 2224
rect 4423 2184 4425 2224
rect 4429 2212 4445 2224
rect 4429 2184 4431 2212
rect 4443 2184 4445 2212
rect 4449 2184 4451 2224
rect 4489 2184 4491 2224
rect 4495 2212 4511 2224
rect 4495 2184 4497 2212
rect 4509 2184 4511 2212
rect 4515 2184 4517 2224
rect 4529 2184 4531 2224
rect 4535 2184 4537 2224
rect 4603 2184 4605 2224
rect 4609 2184 4611 2224
rect 4623 2184 4625 2224
rect 4629 2212 4645 2224
rect 4629 2184 4631 2212
rect 4643 2184 4645 2212
rect 4649 2184 4651 2224
rect 4692 2184 4694 2224
rect 4698 2184 4702 2224
rect 4706 2184 4708 2224
rect 4720 2184 4724 2204
rect 4728 2184 4730 2204
rect 29 2116 31 2156
rect 35 2116 37 2156
rect 49 2116 51 2156
rect 55 2116 57 2156
rect 69 2116 71 2156
rect 75 2116 77 2156
rect 89 2116 91 2156
rect 95 2116 97 2156
rect 109 2116 111 2156
rect 115 2116 117 2156
rect 129 2116 131 2156
rect 135 2116 137 2156
rect 149 2116 151 2156
rect 155 2116 157 2156
rect 169 2116 171 2156
rect 175 2116 177 2156
rect 251 2116 253 2156
rect 257 2116 263 2156
rect 267 2116 269 2156
rect 323 2116 325 2156
rect 329 2116 331 2156
rect 343 2116 345 2156
rect 349 2128 351 2156
rect 363 2128 365 2156
rect 349 2116 365 2128
rect 369 2116 371 2156
rect 412 2116 414 2156
rect 418 2116 422 2156
rect 426 2116 428 2156
rect 440 2116 442 2156
rect 446 2116 450 2156
rect 454 2116 456 2156
rect 533 2116 535 2156
rect 539 2136 541 2156
rect 553 2136 555 2156
rect 559 2136 565 2156
rect 569 2136 573 2156
rect 585 2136 587 2156
rect 591 2136 597 2156
rect 601 2136 603 2156
rect 615 2136 619 2156
rect 623 2136 625 2156
rect 663 2136 665 2156
rect 669 2136 673 2156
rect 677 2136 679 2156
rect 691 2136 693 2156
rect 697 2136 703 2156
rect 707 2136 709 2156
rect 721 2136 725 2156
rect 539 2116 549 2136
rect 712 2116 725 2136
rect 729 2116 731 2156
rect 791 2116 793 2156
rect 797 2116 803 2156
rect 807 2116 809 2156
rect 863 2116 865 2156
rect 869 2136 871 2156
rect 883 2136 885 2156
rect 889 2136 891 2156
rect 903 2136 905 2156
rect 909 2136 911 2156
rect 869 2116 881 2136
rect 951 2116 953 2156
rect 957 2116 963 2156
rect 967 2116 969 2156
rect 1029 2136 1031 2156
rect 1035 2136 1037 2156
rect 1049 2136 1051 2156
rect 1055 2136 1057 2156
rect 1109 2116 1111 2156
rect 1115 2128 1117 2156
rect 1129 2128 1131 2156
rect 1115 2116 1131 2128
rect 1135 2116 1137 2156
rect 1149 2116 1151 2156
rect 1155 2116 1157 2156
rect 1211 2116 1213 2156
rect 1217 2116 1223 2156
rect 1227 2116 1229 2156
rect 1289 2136 1291 2156
rect 1295 2136 1297 2156
rect 1309 2136 1311 2156
rect 1315 2136 1317 2156
rect 1369 2116 1371 2156
rect 1375 2136 1379 2156
rect 1391 2136 1393 2156
rect 1397 2136 1403 2156
rect 1407 2136 1409 2156
rect 1421 2136 1423 2156
rect 1427 2136 1431 2156
rect 1435 2136 1437 2156
rect 1475 2136 1477 2156
rect 1481 2136 1485 2156
rect 1497 2136 1499 2156
rect 1503 2136 1509 2156
rect 1513 2136 1515 2156
rect 1527 2136 1531 2156
rect 1535 2136 1541 2156
rect 1545 2136 1547 2156
rect 1559 2136 1561 2156
rect 1375 2116 1388 2136
rect 1551 2116 1561 2136
rect 1565 2116 1567 2156
rect 1630 2136 1632 2156
rect 1636 2136 1640 2156
rect 1652 2116 1654 2156
rect 1658 2116 1662 2156
rect 1666 2116 1668 2156
rect 1721 2116 1723 2156
rect 1727 2116 1729 2156
rect 1741 2136 1745 2156
rect 1749 2136 1751 2156
rect 1789 2116 1791 2156
rect 1795 2136 1799 2156
rect 1811 2136 1813 2156
rect 1817 2136 1823 2156
rect 1827 2136 1829 2156
rect 1841 2136 1843 2156
rect 1847 2136 1851 2156
rect 1855 2136 1857 2156
rect 1895 2136 1897 2156
rect 1901 2136 1905 2156
rect 1917 2136 1919 2156
rect 1923 2136 1929 2156
rect 1933 2136 1935 2156
rect 1947 2136 1951 2156
rect 1955 2136 1961 2156
rect 1965 2136 1967 2156
rect 1979 2136 1981 2156
rect 1795 2116 1808 2136
rect 1971 2116 1981 2136
rect 1985 2116 1987 2156
rect 2043 2136 2045 2156
rect 2049 2136 2051 2156
rect 2111 2116 2113 2156
rect 2117 2116 2123 2156
rect 2127 2116 2129 2156
rect 2169 2136 2171 2156
rect 2175 2136 2179 2156
rect 2191 2116 2193 2156
rect 2197 2116 2199 2156
rect 2251 2116 2253 2156
rect 2257 2116 2263 2156
rect 2267 2116 2269 2156
rect 2343 2116 2345 2156
rect 2349 2116 2351 2156
rect 2363 2116 2365 2156
rect 2369 2128 2371 2156
rect 2383 2128 2385 2156
rect 2369 2116 2385 2128
rect 2389 2116 2391 2156
rect 2451 2116 2453 2156
rect 2457 2116 2463 2156
rect 2467 2116 2469 2156
rect 2531 2116 2533 2156
rect 2537 2116 2543 2156
rect 2547 2116 2549 2156
rect 2603 2116 2605 2156
rect 2609 2116 2611 2156
rect 2623 2116 2625 2156
rect 2629 2128 2631 2156
rect 2643 2128 2645 2156
rect 2629 2116 2645 2128
rect 2649 2116 2651 2156
rect 2703 2116 2705 2156
rect 2709 2116 2711 2156
rect 2723 2116 2725 2156
rect 2729 2128 2731 2156
rect 2743 2128 2745 2156
rect 2729 2116 2745 2128
rect 2749 2116 2751 2156
rect 2793 2116 2795 2156
rect 2799 2136 2801 2156
rect 2813 2136 2815 2156
rect 2819 2136 2825 2156
rect 2829 2136 2833 2156
rect 2845 2136 2847 2156
rect 2851 2136 2857 2156
rect 2861 2136 2863 2156
rect 2875 2136 2879 2156
rect 2883 2136 2885 2156
rect 2923 2136 2925 2156
rect 2929 2136 2933 2156
rect 2937 2136 2939 2156
rect 2951 2136 2953 2156
rect 2957 2136 2963 2156
rect 2967 2136 2969 2156
rect 2981 2136 2985 2156
rect 2799 2116 2809 2136
rect 2972 2116 2985 2136
rect 2989 2116 2991 2156
rect 3029 2116 3031 2156
rect 3035 2116 3041 2156
rect 3045 2116 3047 2156
rect 3059 2116 3061 2156
rect 3065 2116 3067 2156
rect 3143 2116 3145 2156
rect 3149 2116 3151 2156
rect 3163 2116 3165 2156
rect 3169 2128 3171 2156
rect 3183 2128 3185 2156
rect 3169 2116 3185 2128
rect 3189 2116 3191 2156
rect 3243 2116 3245 2156
rect 3249 2116 3251 2156
rect 3263 2116 3265 2156
rect 3269 2128 3271 2156
rect 3283 2128 3285 2156
rect 3269 2116 3285 2128
rect 3289 2116 3291 2156
rect 3331 2116 3333 2156
rect 3337 2116 3343 2156
rect 3347 2116 3349 2156
rect 3423 2116 3425 2156
rect 3429 2116 3431 2156
rect 3443 2116 3445 2156
rect 3449 2128 3451 2156
rect 3463 2128 3465 2156
rect 3449 2116 3465 2128
rect 3469 2116 3471 2156
rect 3510 2096 3512 2156
rect 3516 2096 3520 2156
rect 3524 2096 3528 2156
rect 3532 2098 3534 2156
rect 3609 2136 3611 2156
rect 3615 2136 3617 2156
rect 3532 2096 3546 2098
rect 3670 2096 3672 2156
rect 3676 2096 3680 2156
rect 3684 2096 3688 2156
rect 3692 2098 3694 2156
rect 3771 2116 3773 2156
rect 3777 2116 3783 2156
rect 3787 2116 3789 2156
rect 3849 2136 3851 2156
rect 3855 2136 3859 2156
rect 3692 2096 3706 2098
rect 3871 2116 3873 2156
rect 3877 2116 3879 2156
rect 3929 2116 3931 2156
rect 3935 2128 3937 2156
rect 3949 2128 3951 2156
rect 3935 2116 3951 2128
rect 3955 2116 3957 2156
rect 3969 2116 3971 2156
rect 3975 2116 3977 2156
rect 4051 2116 4053 2156
rect 4057 2116 4063 2156
rect 4067 2116 4069 2156
rect 4131 2116 4133 2156
rect 4137 2116 4143 2156
rect 4147 2116 4149 2156
rect 4211 2116 4213 2156
rect 4217 2116 4223 2156
rect 4227 2116 4229 2156
rect 4269 2116 4271 2156
rect 4275 2116 4281 2156
rect 4285 2116 4287 2156
rect 4299 2116 4301 2156
rect 4305 2116 4307 2156
rect 4372 2116 4374 2156
rect 4378 2116 4382 2156
rect 4386 2116 4388 2156
rect 4400 2136 4404 2156
rect 4408 2136 4410 2156
rect 4490 2136 4492 2156
rect 4496 2136 4500 2156
rect 4512 2116 4514 2156
rect 4518 2116 4522 2156
rect 4526 2116 4528 2156
rect 4570 2096 4572 2156
rect 4576 2096 4580 2156
rect 4584 2096 4588 2156
rect 4592 2098 4594 2156
rect 4592 2096 4606 2098
rect 4670 2096 4672 2156
rect 4676 2096 4680 2156
rect 4684 2096 4688 2156
rect 4692 2098 4694 2156
rect 4692 2096 4706 2098
rect 33 1704 35 1744
rect 39 1724 49 1744
rect 212 1724 225 1744
rect 39 1704 41 1724
rect 53 1704 55 1724
rect 59 1704 65 1724
rect 69 1704 73 1724
rect 85 1704 87 1724
rect 91 1704 97 1724
rect 101 1704 103 1724
rect 115 1704 119 1724
rect 123 1704 125 1724
rect 163 1704 165 1724
rect 169 1704 173 1724
rect 177 1704 179 1724
rect 191 1704 193 1724
rect 197 1704 203 1724
rect 207 1704 209 1724
rect 221 1704 225 1724
rect 229 1704 231 1744
rect 269 1704 271 1744
rect 275 1732 291 1744
rect 275 1704 277 1732
rect 289 1704 291 1732
rect 295 1704 297 1744
rect 309 1704 311 1744
rect 315 1704 317 1744
rect 383 1704 385 1744
rect 389 1704 391 1744
rect 403 1704 405 1744
rect 409 1732 425 1744
rect 409 1704 411 1732
rect 423 1704 425 1732
rect 429 1704 431 1744
rect 483 1704 485 1744
rect 489 1704 491 1744
rect 503 1704 505 1744
rect 509 1732 525 1744
rect 509 1704 511 1732
rect 523 1704 525 1732
rect 529 1704 531 1744
rect 583 1704 585 1744
rect 589 1704 591 1744
rect 603 1704 605 1744
rect 609 1732 625 1744
rect 609 1704 611 1732
rect 623 1704 625 1732
rect 629 1704 631 1744
rect 669 1704 671 1724
rect 675 1704 677 1724
rect 729 1704 731 1724
rect 735 1704 737 1724
rect 803 1704 805 1724
rect 809 1704 811 1724
rect 823 1704 825 1724
rect 829 1704 831 1724
rect 870 1704 872 1764
rect 876 1704 880 1764
rect 884 1704 888 1764
rect 892 1762 906 1764
rect 892 1704 894 1762
rect 973 1704 975 1744
rect 979 1724 989 1744
rect 1152 1724 1165 1744
rect 979 1704 981 1724
rect 993 1704 995 1724
rect 999 1704 1005 1724
rect 1009 1704 1013 1724
rect 1025 1704 1027 1724
rect 1031 1704 1037 1724
rect 1041 1704 1043 1724
rect 1055 1704 1059 1724
rect 1063 1704 1065 1724
rect 1103 1704 1105 1724
rect 1109 1704 1113 1724
rect 1117 1704 1119 1724
rect 1131 1704 1133 1724
rect 1137 1704 1143 1724
rect 1147 1704 1149 1724
rect 1161 1704 1165 1724
rect 1169 1704 1171 1744
rect 1211 1704 1213 1744
rect 1217 1704 1223 1744
rect 1227 1704 1229 1744
rect 1303 1704 1305 1744
rect 1309 1704 1311 1744
rect 1323 1704 1325 1744
rect 1329 1732 1345 1744
rect 1329 1704 1331 1732
rect 1343 1704 1345 1732
rect 1349 1704 1351 1744
rect 1403 1704 1405 1744
rect 1409 1704 1411 1744
rect 1423 1704 1425 1744
rect 1429 1704 1431 1744
rect 1443 1704 1445 1744
rect 1449 1704 1451 1744
rect 1463 1704 1465 1744
rect 1469 1704 1471 1744
rect 1483 1704 1485 1744
rect 1489 1704 1491 1744
rect 1503 1704 1505 1744
rect 1509 1704 1511 1744
rect 1523 1704 1525 1744
rect 1529 1704 1531 1744
rect 1543 1704 1545 1744
rect 1549 1704 1551 1744
rect 1593 1704 1595 1744
rect 1599 1724 1609 1744
rect 1772 1724 1785 1744
rect 1599 1704 1601 1724
rect 1613 1704 1615 1724
rect 1619 1704 1625 1724
rect 1629 1704 1633 1724
rect 1645 1704 1647 1724
rect 1651 1704 1657 1724
rect 1661 1704 1663 1724
rect 1675 1704 1679 1724
rect 1683 1704 1685 1724
rect 1723 1704 1725 1724
rect 1729 1704 1733 1724
rect 1737 1704 1739 1724
rect 1751 1704 1753 1724
rect 1757 1704 1763 1724
rect 1767 1704 1769 1724
rect 1781 1704 1785 1724
rect 1789 1704 1791 1744
rect 1850 1704 1852 1724
rect 1856 1704 1860 1724
rect 1872 1704 1874 1744
rect 1878 1704 1882 1744
rect 1886 1704 1888 1744
rect 1929 1704 1931 1724
rect 1935 1704 1937 1724
rect 1949 1704 1951 1724
rect 1955 1704 1957 1724
rect 2030 1704 2032 1724
rect 2036 1704 2040 1724
rect 2052 1704 2054 1744
rect 2058 1704 2062 1744
rect 2066 1704 2068 1744
rect 2123 1704 2125 1724
rect 2129 1704 2131 1724
rect 2143 1704 2145 1724
rect 2149 1704 2151 1724
rect 2192 1704 2194 1744
rect 2198 1704 2202 1744
rect 2206 1704 2208 1744
rect 2220 1704 2224 1724
rect 2228 1704 2230 1724
rect 2289 1704 2291 1744
rect 2295 1724 2308 1744
rect 2471 1724 2481 1744
rect 2295 1704 2299 1724
rect 2311 1704 2313 1724
rect 2317 1704 2323 1724
rect 2327 1704 2329 1724
rect 2341 1704 2343 1724
rect 2347 1704 2351 1724
rect 2355 1704 2357 1724
rect 2395 1704 2397 1724
rect 2401 1704 2405 1724
rect 2417 1704 2419 1724
rect 2423 1704 2429 1724
rect 2433 1704 2435 1724
rect 2447 1704 2451 1724
rect 2455 1704 2461 1724
rect 2465 1704 2467 1724
rect 2479 1704 2481 1724
rect 2485 1704 2487 1744
rect 2533 1704 2535 1744
rect 2539 1724 2549 1744
rect 2712 1724 2725 1744
rect 2539 1704 2541 1724
rect 2553 1704 2555 1724
rect 2559 1704 2565 1724
rect 2569 1704 2573 1724
rect 2585 1704 2587 1724
rect 2591 1704 2597 1724
rect 2601 1704 2603 1724
rect 2615 1704 2619 1724
rect 2623 1704 2625 1724
rect 2663 1704 2665 1724
rect 2669 1704 2673 1724
rect 2677 1704 2679 1724
rect 2691 1704 2693 1724
rect 2697 1704 2703 1724
rect 2707 1704 2709 1724
rect 2721 1704 2725 1724
rect 2729 1704 2731 1744
rect 2773 1704 2775 1744
rect 2779 1724 2789 1744
rect 2952 1724 2965 1744
rect 2779 1704 2781 1724
rect 2793 1704 2795 1724
rect 2799 1704 2805 1724
rect 2809 1704 2813 1724
rect 2825 1704 2827 1724
rect 2831 1704 2837 1724
rect 2841 1704 2843 1724
rect 2855 1704 2859 1724
rect 2863 1704 2865 1724
rect 2903 1704 2905 1724
rect 2909 1704 2913 1724
rect 2917 1704 2919 1724
rect 2931 1704 2933 1724
rect 2937 1704 2943 1724
rect 2947 1704 2949 1724
rect 2961 1704 2965 1724
rect 2969 1704 2971 1744
rect 3023 1704 3025 1744
rect 3029 1704 3031 1744
rect 3091 1704 3093 1744
rect 3097 1704 3103 1744
rect 3107 1704 3109 1744
rect 3163 1704 3165 1744
rect 3169 1704 3171 1744
rect 3212 1704 3214 1744
rect 3218 1704 3222 1744
rect 3226 1704 3228 1744
rect 3240 1704 3244 1724
rect 3248 1704 3250 1724
rect 3309 1704 3311 1724
rect 3315 1704 3317 1724
rect 3329 1704 3331 1724
rect 3335 1704 3337 1724
rect 3413 1704 3415 1744
rect 3419 1704 3421 1744
rect 3433 1704 3435 1744
rect 3439 1704 3445 1744
rect 3449 1704 3451 1744
rect 3489 1704 3491 1744
rect 3495 1704 3497 1744
rect 3584 1704 3586 1744
rect 3590 1704 3594 1744
rect 3598 1704 3600 1744
rect 3612 1704 3614 1744
rect 3618 1704 3622 1744
rect 3626 1704 3628 1744
rect 3683 1704 3685 1744
rect 3689 1704 3691 1744
rect 3743 1704 3745 1724
rect 3749 1704 3751 1724
rect 3763 1704 3765 1724
rect 3769 1704 3771 1724
rect 3809 1704 3811 1724
rect 3815 1704 3819 1724
rect 3831 1704 3833 1744
rect 3837 1704 3839 1744
rect 3889 1704 3891 1744
rect 3895 1704 3901 1744
rect 3905 1704 3907 1744
rect 3919 1704 3921 1744
rect 3925 1704 3927 1744
rect 4024 1704 4026 1744
rect 4030 1704 4034 1744
rect 4038 1704 4040 1744
rect 4052 1704 4054 1744
rect 4058 1704 4062 1744
rect 4066 1704 4068 1744
rect 4112 1704 4114 1744
rect 4118 1704 4122 1744
rect 4126 1704 4128 1744
rect 4140 1704 4142 1744
rect 4146 1704 4150 1744
rect 4154 1704 4156 1744
rect 4231 1704 4233 1744
rect 4237 1704 4243 1744
rect 4247 1704 4249 1744
rect 4309 1704 4311 1744
rect 4315 1704 4321 1744
rect 4325 1704 4327 1744
rect 4339 1704 4341 1744
rect 4345 1704 4347 1744
rect 4412 1704 4414 1744
rect 4418 1704 4422 1744
rect 4426 1704 4428 1744
rect 4440 1704 4442 1744
rect 4446 1704 4450 1744
rect 4454 1704 4456 1744
rect 4543 1704 4545 1724
rect 4549 1704 4551 1724
rect 4589 1704 4591 1744
rect 4595 1732 4611 1744
rect 4595 1704 4597 1732
rect 4609 1704 4611 1732
rect 4615 1704 4617 1744
rect 4629 1704 4631 1744
rect 4635 1704 4637 1744
rect 4689 1704 4691 1724
rect 4695 1704 4697 1724
rect 29 1636 31 1676
rect 35 1636 37 1676
rect 49 1636 51 1676
rect 55 1636 57 1676
rect 69 1636 71 1676
rect 75 1636 77 1676
rect 89 1636 91 1676
rect 95 1636 97 1676
rect 109 1636 111 1676
rect 115 1636 117 1676
rect 129 1636 131 1676
rect 135 1636 137 1676
rect 149 1636 151 1676
rect 155 1636 157 1676
rect 169 1636 171 1676
rect 175 1636 177 1676
rect 243 1656 245 1676
rect 249 1656 251 1676
rect 263 1656 265 1676
rect 269 1656 271 1676
rect 321 1636 323 1676
rect 327 1636 329 1676
rect 341 1656 345 1676
rect 349 1656 351 1676
rect 393 1636 395 1676
rect 399 1656 401 1676
rect 413 1656 415 1676
rect 419 1656 425 1676
rect 429 1656 433 1676
rect 445 1656 447 1676
rect 451 1656 457 1676
rect 461 1656 463 1676
rect 475 1656 479 1676
rect 483 1656 485 1676
rect 523 1656 525 1676
rect 529 1656 533 1676
rect 537 1656 539 1676
rect 551 1656 553 1676
rect 557 1656 563 1676
rect 567 1656 569 1676
rect 581 1656 585 1676
rect 399 1636 409 1656
rect 572 1636 585 1656
rect 589 1636 591 1676
rect 633 1636 635 1676
rect 639 1656 641 1676
rect 653 1656 655 1676
rect 659 1656 665 1676
rect 669 1656 673 1676
rect 685 1656 687 1676
rect 691 1656 697 1676
rect 701 1656 703 1676
rect 715 1656 719 1676
rect 723 1656 725 1676
rect 763 1656 765 1676
rect 769 1656 773 1676
rect 777 1656 779 1676
rect 791 1656 793 1676
rect 797 1656 803 1676
rect 807 1656 809 1676
rect 821 1656 825 1676
rect 639 1636 649 1656
rect 812 1636 825 1656
rect 829 1636 831 1676
rect 869 1636 871 1676
rect 875 1656 879 1676
rect 891 1656 893 1676
rect 897 1656 903 1676
rect 907 1656 909 1676
rect 921 1656 923 1676
rect 927 1656 931 1676
rect 935 1656 937 1676
rect 975 1656 977 1676
rect 981 1656 985 1676
rect 997 1656 999 1676
rect 1003 1656 1009 1676
rect 1013 1656 1015 1676
rect 1027 1656 1031 1676
rect 1035 1656 1041 1676
rect 1045 1656 1047 1676
rect 1059 1656 1061 1676
rect 875 1636 888 1656
rect 1051 1636 1061 1656
rect 1065 1636 1067 1676
rect 1131 1636 1133 1676
rect 1137 1636 1143 1676
rect 1147 1636 1149 1676
rect 1203 1636 1205 1676
rect 1209 1636 1211 1676
rect 1223 1636 1225 1676
rect 1229 1648 1231 1676
rect 1243 1648 1245 1676
rect 1229 1636 1245 1648
rect 1249 1636 1251 1676
rect 1289 1636 1291 1676
rect 1295 1656 1299 1676
rect 1311 1656 1313 1676
rect 1317 1656 1323 1676
rect 1327 1656 1329 1676
rect 1341 1656 1343 1676
rect 1347 1656 1351 1676
rect 1355 1656 1357 1676
rect 1395 1656 1397 1676
rect 1401 1656 1405 1676
rect 1417 1656 1419 1676
rect 1423 1656 1429 1676
rect 1433 1656 1435 1676
rect 1447 1656 1451 1676
rect 1455 1656 1461 1676
rect 1465 1656 1467 1676
rect 1479 1656 1481 1676
rect 1295 1636 1308 1656
rect 1471 1636 1481 1656
rect 1485 1636 1487 1676
rect 1533 1636 1535 1676
rect 1539 1656 1541 1676
rect 1553 1656 1555 1676
rect 1559 1656 1565 1676
rect 1569 1656 1573 1676
rect 1585 1656 1587 1676
rect 1591 1656 1597 1676
rect 1601 1656 1603 1676
rect 1615 1656 1619 1676
rect 1623 1656 1625 1676
rect 1663 1656 1665 1676
rect 1669 1656 1673 1676
rect 1677 1656 1679 1676
rect 1691 1656 1693 1676
rect 1697 1656 1703 1676
rect 1707 1656 1709 1676
rect 1721 1656 1725 1676
rect 1539 1636 1549 1656
rect 1712 1636 1725 1656
rect 1729 1636 1731 1676
rect 1790 1656 1792 1676
rect 1796 1656 1800 1676
rect 1812 1636 1814 1676
rect 1818 1636 1822 1676
rect 1826 1636 1828 1676
rect 1869 1656 1871 1676
rect 1875 1656 1877 1676
rect 1889 1656 1891 1676
rect 1895 1656 1897 1676
rect 1953 1636 1955 1676
rect 1959 1656 1961 1676
rect 1973 1656 1975 1676
rect 1979 1656 1985 1676
rect 1989 1656 1993 1676
rect 2005 1656 2007 1676
rect 2011 1656 2017 1676
rect 2021 1656 2023 1676
rect 2035 1656 2039 1676
rect 2043 1656 2045 1676
rect 2083 1656 2085 1676
rect 2089 1656 2093 1676
rect 2097 1656 2099 1676
rect 2111 1656 2113 1676
rect 2117 1656 2123 1676
rect 2127 1656 2129 1676
rect 2141 1656 2145 1676
rect 1959 1636 1969 1656
rect 2132 1636 2145 1656
rect 2149 1636 2151 1676
rect 2203 1656 2205 1676
rect 2209 1656 2211 1676
rect 2223 1656 2225 1676
rect 2229 1656 2231 1676
rect 2291 1636 2293 1676
rect 2297 1636 2303 1676
rect 2307 1636 2309 1676
rect 2349 1636 2351 1676
rect 2355 1648 2357 1676
rect 2369 1648 2371 1676
rect 2355 1636 2371 1648
rect 2375 1636 2377 1676
rect 2389 1636 2391 1676
rect 2395 1636 2397 1676
rect 2449 1636 2451 1676
rect 2455 1656 2459 1676
rect 2471 1656 2473 1676
rect 2477 1656 2483 1676
rect 2487 1656 2489 1676
rect 2501 1656 2503 1676
rect 2507 1656 2511 1676
rect 2515 1656 2517 1676
rect 2555 1656 2557 1676
rect 2561 1656 2565 1676
rect 2577 1656 2579 1676
rect 2583 1656 2589 1676
rect 2593 1656 2595 1676
rect 2607 1656 2611 1676
rect 2615 1656 2621 1676
rect 2625 1656 2627 1676
rect 2639 1656 2641 1676
rect 2455 1636 2468 1656
rect 2631 1636 2641 1656
rect 2645 1636 2647 1676
rect 2693 1636 2695 1676
rect 2699 1656 2701 1676
rect 2713 1656 2715 1676
rect 2719 1656 2725 1676
rect 2729 1656 2733 1676
rect 2745 1656 2747 1676
rect 2751 1656 2757 1676
rect 2761 1656 2763 1676
rect 2775 1656 2779 1676
rect 2783 1656 2785 1676
rect 2823 1656 2825 1676
rect 2829 1656 2833 1676
rect 2837 1656 2839 1676
rect 2851 1656 2853 1676
rect 2857 1656 2863 1676
rect 2867 1656 2869 1676
rect 2881 1656 2885 1676
rect 2699 1636 2709 1656
rect 2872 1636 2885 1656
rect 2889 1636 2891 1676
rect 2929 1636 2931 1676
rect 2935 1636 2937 1676
rect 2991 1636 2993 1676
rect 2997 1636 3003 1676
rect 3007 1636 3009 1676
rect 3091 1636 3093 1676
rect 3097 1636 3103 1676
rect 3107 1636 3109 1676
rect 3149 1636 3151 1676
rect 3155 1648 3157 1676
rect 3169 1648 3171 1676
rect 3155 1636 3171 1648
rect 3175 1636 3177 1676
rect 3189 1636 3191 1676
rect 3195 1636 3197 1676
rect 3251 1636 3253 1676
rect 3257 1636 3263 1676
rect 3267 1636 3269 1676
rect 3351 1636 3353 1676
rect 3357 1636 3363 1676
rect 3367 1636 3369 1676
rect 3423 1636 3425 1676
rect 3429 1636 3431 1676
rect 3443 1636 3445 1676
rect 3449 1648 3451 1676
rect 3463 1648 3465 1676
rect 3449 1636 3465 1648
rect 3469 1636 3471 1676
rect 3510 1616 3512 1676
rect 3516 1616 3520 1676
rect 3524 1616 3528 1676
rect 3532 1618 3534 1676
rect 3623 1636 3625 1676
rect 3629 1664 3645 1676
rect 3629 1636 3631 1664
rect 3643 1636 3645 1664
rect 3649 1636 3651 1676
rect 3663 1636 3665 1676
rect 3669 1646 3671 1676
rect 3683 1646 3685 1676
rect 3669 1636 3685 1646
rect 3689 1636 3691 1676
rect 3729 1656 3731 1676
rect 3735 1656 3737 1676
rect 3532 1616 3546 1618
rect 3790 1616 3792 1676
rect 3796 1616 3800 1676
rect 3804 1616 3808 1676
rect 3812 1618 3814 1676
rect 3892 1636 3894 1676
rect 3898 1636 3902 1676
rect 3906 1636 3908 1676
rect 3920 1656 3924 1676
rect 3928 1656 3930 1676
rect 3812 1616 3826 1618
rect 3989 1636 3991 1676
rect 3995 1648 3997 1676
rect 4009 1648 4011 1676
rect 3995 1636 4011 1648
rect 4015 1636 4017 1676
rect 4029 1636 4031 1676
rect 4035 1636 4037 1676
rect 4111 1636 4113 1676
rect 4117 1636 4123 1676
rect 4127 1636 4129 1676
rect 4172 1636 4174 1676
rect 4178 1636 4182 1676
rect 4186 1636 4188 1676
rect 4200 1656 4204 1676
rect 4208 1656 4210 1676
rect 4269 1636 4271 1676
rect 4275 1648 4277 1676
rect 4289 1648 4291 1676
rect 4275 1636 4291 1648
rect 4295 1636 4297 1676
rect 4309 1636 4311 1676
rect 4315 1636 4317 1676
rect 4369 1656 4371 1676
rect 4375 1656 4377 1676
rect 4429 1656 4431 1676
rect 4435 1656 4437 1676
rect 4449 1656 4451 1676
rect 4455 1656 4457 1676
rect 4511 1636 4513 1676
rect 4517 1636 4523 1676
rect 4527 1636 4529 1676
rect 4591 1636 4593 1676
rect 4597 1636 4603 1676
rect 4607 1636 4609 1676
rect 4671 1636 4673 1676
rect 4677 1636 4683 1676
rect 4687 1636 4689 1676
rect 29 1224 31 1264
rect 35 1244 48 1264
rect 211 1244 221 1264
rect 35 1224 39 1244
rect 51 1224 53 1244
rect 57 1224 63 1244
rect 67 1224 69 1244
rect 81 1224 83 1244
rect 87 1224 91 1244
rect 95 1224 97 1244
rect 135 1224 137 1244
rect 141 1224 145 1244
rect 157 1224 159 1244
rect 163 1224 169 1244
rect 173 1224 175 1244
rect 187 1224 191 1244
rect 195 1224 201 1244
rect 205 1224 207 1244
rect 219 1224 221 1244
rect 225 1224 227 1264
rect 273 1224 275 1264
rect 279 1244 289 1264
rect 452 1244 465 1264
rect 279 1224 281 1244
rect 293 1224 295 1244
rect 299 1224 305 1244
rect 309 1224 313 1244
rect 325 1224 327 1244
rect 331 1224 337 1244
rect 341 1224 343 1244
rect 355 1224 359 1244
rect 363 1224 365 1244
rect 403 1224 405 1244
rect 409 1224 413 1244
rect 417 1224 419 1244
rect 431 1224 433 1244
rect 437 1224 443 1244
rect 447 1224 449 1244
rect 461 1224 465 1244
rect 469 1224 471 1264
rect 511 1224 513 1264
rect 517 1224 523 1264
rect 527 1224 529 1264
rect 603 1224 605 1264
rect 609 1224 611 1264
rect 623 1224 625 1264
rect 629 1252 645 1264
rect 629 1224 631 1252
rect 643 1224 645 1252
rect 649 1224 651 1264
rect 703 1224 705 1264
rect 709 1224 711 1264
rect 723 1224 725 1264
rect 729 1252 745 1264
rect 729 1224 731 1252
rect 743 1224 745 1252
rect 749 1224 751 1264
rect 801 1224 803 1264
rect 807 1224 809 1264
rect 821 1224 825 1244
rect 829 1224 831 1244
rect 871 1224 873 1264
rect 877 1224 883 1264
rect 887 1224 889 1264
rect 963 1224 965 1264
rect 969 1224 971 1264
rect 983 1224 985 1264
rect 989 1252 1005 1264
rect 989 1224 991 1252
rect 1003 1224 1005 1252
rect 1009 1224 1011 1264
rect 1063 1224 1065 1244
rect 1069 1224 1071 1244
rect 1109 1224 1111 1264
rect 1115 1224 1117 1264
rect 1129 1224 1131 1264
rect 1135 1224 1137 1264
rect 1149 1224 1151 1264
rect 1155 1224 1157 1264
rect 1169 1224 1171 1264
rect 1175 1224 1177 1264
rect 1251 1224 1253 1264
rect 1257 1224 1263 1264
rect 1267 1224 1269 1264
rect 1323 1224 1325 1264
rect 1329 1224 1331 1264
rect 1343 1224 1345 1264
rect 1349 1252 1365 1264
rect 1349 1224 1351 1252
rect 1363 1224 1365 1252
rect 1369 1224 1371 1264
rect 1431 1224 1433 1264
rect 1437 1224 1443 1264
rect 1447 1224 1449 1264
rect 1503 1224 1505 1264
rect 1509 1224 1511 1264
rect 1523 1224 1525 1264
rect 1529 1252 1545 1264
rect 1529 1224 1531 1252
rect 1543 1224 1545 1252
rect 1549 1224 1551 1264
rect 1589 1224 1591 1244
rect 1595 1224 1599 1244
rect 1611 1224 1613 1264
rect 1617 1224 1619 1264
rect 1671 1224 1673 1264
rect 1677 1224 1683 1264
rect 1687 1224 1689 1264
rect 1763 1224 1765 1264
rect 1769 1224 1771 1264
rect 1783 1224 1785 1264
rect 1789 1252 1805 1264
rect 1789 1224 1791 1252
rect 1803 1224 1805 1252
rect 1809 1224 1811 1264
rect 1849 1224 1851 1264
rect 1855 1244 1868 1264
rect 2031 1244 2041 1264
rect 1855 1224 1859 1244
rect 1871 1224 1873 1244
rect 1877 1224 1883 1244
rect 1887 1224 1889 1244
rect 1901 1224 1903 1244
rect 1907 1224 1911 1244
rect 1915 1224 1917 1244
rect 1955 1224 1957 1244
rect 1961 1224 1965 1244
rect 1977 1224 1979 1244
rect 1983 1224 1989 1244
rect 1993 1224 1995 1244
rect 2007 1224 2011 1244
rect 2015 1224 2021 1244
rect 2025 1224 2027 1244
rect 2039 1224 2041 1244
rect 2045 1224 2047 1264
rect 2089 1224 2091 1244
rect 2095 1224 2097 1244
rect 2149 1224 2151 1264
rect 2155 1252 2171 1264
rect 2155 1224 2157 1252
rect 2169 1224 2171 1252
rect 2175 1224 2177 1264
rect 2189 1224 2191 1264
rect 2195 1224 2197 1264
rect 2271 1224 2273 1264
rect 2277 1224 2283 1264
rect 2287 1224 2289 1264
rect 2343 1224 2345 1244
rect 2349 1224 2351 1244
rect 2363 1224 2365 1244
rect 2369 1224 2371 1244
rect 2423 1224 2425 1244
rect 2429 1224 2431 1244
rect 2469 1224 2471 1244
rect 2475 1224 2477 1244
rect 2489 1224 2491 1244
rect 2495 1224 2497 1244
rect 2549 1224 2551 1264
rect 2555 1244 2568 1264
rect 2731 1244 2741 1264
rect 2555 1224 2559 1244
rect 2571 1224 2573 1244
rect 2577 1224 2583 1244
rect 2587 1224 2589 1244
rect 2601 1224 2603 1244
rect 2607 1224 2611 1244
rect 2615 1224 2617 1244
rect 2655 1224 2657 1244
rect 2661 1224 2665 1244
rect 2677 1224 2679 1244
rect 2683 1224 2689 1244
rect 2693 1224 2695 1244
rect 2707 1224 2711 1244
rect 2715 1224 2721 1244
rect 2725 1224 2727 1244
rect 2739 1224 2741 1244
rect 2745 1224 2747 1264
rect 2789 1224 2791 1244
rect 2795 1224 2797 1244
rect 2809 1224 2811 1244
rect 2815 1224 2817 1244
rect 2883 1224 2885 1264
rect 2889 1224 2891 1264
rect 2929 1224 2931 1264
rect 2935 1252 2951 1264
rect 2935 1224 2937 1252
rect 2949 1224 2951 1252
rect 2955 1224 2957 1264
rect 2969 1224 2971 1264
rect 2975 1224 2977 1264
rect 3029 1224 3031 1264
rect 3035 1252 3051 1264
rect 3035 1224 3037 1252
rect 3049 1224 3051 1252
rect 3055 1224 3057 1264
rect 3069 1224 3071 1264
rect 3075 1224 3077 1264
rect 3129 1224 3131 1264
rect 3135 1252 3151 1264
rect 3135 1224 3137 1252
rect 3149 1224 3151 1252
rect 3155 1224 3157 1264
rect 3169 1224 3171 1264
rect 3175 1224 3177 1264
rect 3229 1224 3231 1264
rect 3235 1224 3241 1264
rect 3245 1224 3247 1264
rect 3259 1224 3261 1264
rect 3265 1224 3267 1264
rect 3343 1224 3345 1244
rect 3349 1224 3351 1244
rect 3363 1224 3365 1244
rect 3369 1224 3371 1244
rect 3410 1224 3412 1284
rect 3416 1224 3420 1284
rect 3424 1224 3428 1284
rect 3432 1282 3446 1284
rect 3432 1224 3434 1282
rect 3523 1224 3525 1264
rect 3529 1224 3531 1264
rect 3543 1224 3545 1264
rect 3549 1252 3565 1264
rect 3549 1224 3551 1252
rect 3563 1224 3565 1252
rect 3569 1224 3571 1264
rect 3609 1224 3611 1264
rect 3615 1252 3631 1264
rect 3615 1224 3617 1252
rect 3629 1224 3631 1252
rect 3635 1224 3637 1264
rect 3649 1224 3651 1264
rect 3655 1224 3657 1264
rect 3731 1224 3733 1264
rect 3737 1224 3743 1264
rect 3747 1224 3749 1264
rect 3811 1224 3813 1264
rect 3817 1224 3823 1264
rect 3827 1224 3829 1264
rect 3869 1224 3871 1264
rect 3875 1224 3881 1264
rect 3885 1224 3887 1264
rect 3899 1224 3901 1264
rect 3905 1224 3907 1264
rect 3983 1224 3985 1264
rect 3989 1224 3991 1264
rect 4003 1224 4005 1264
rect 4009 1252 4025 1264
rect 4009 1224 4011 1252
rect 4023 1224 4025 1252
rect 4029 1224 4031 1264
rect 4069 1224 4071 1244
rect 4075 1224 4077 1244
rect 4151 1224 4153 1264
rect 4157 1224 4163 1264
rect 4167 1224 4169 1264
rect 4231 1224 4233 1264
rect 4237 1224 4243 1264
rect 4247 1224 4249 1264
rect 4303 1224 4305 1244
rect 4309 1224 4311 1244
rect 4323 1224 4325 1244
rect 4329 1224 4331 1244
rect 4383 1224 4385 1264
rect 4389 1224 4391 1264
rect 4403 1224 4405 1264
rect 4409 1252 4425 1264
rect 4409 1224 4411 1252
rect 4423 1224 4425 1252
rect 4429 1224 4431 1264
rect 4469 1224 4471 1264
rect 4475 1252 4491 1264
rect 4475 1224 4477 1252
rect 4489 1224 4491 1252
rect 4495 1224 4497 1264
rect 4509 1224 4511 1264
rect 4515 1224 4517 1264
rect 4590 1224 4592 1244
rect 4596 1224 4600 1244
rect 4612 1224 4614 1264
rect 4618 1224 4622 1264
rect 4626 1224 4628 1264
rect 4671 1224 4673 1264
rect 4677 1224 4683 1264
rect 4687 1224 4689 1264
rect 29 1176 31 1196
rect 35 1176 37 1196
rect 111 1156 113 1196
rect 117 1156 123 1196
rect 127 1156 129 1196
rect 183 1156 185 1196
rect 189 1156 191 1196
rect 203 1156 205 1196
rect 209 1168 211 1196
rect 223 1168 225 1196
rect 209 1156 225 1168
rect 229 1156 231 1196
rect 272 1156 274 1196
rect 278 1156 282 1196
rect 286 1156 288 1196
rect 300 1156 302 1196
rect 306 1156 310 1196
rect 314 1156 316 1196
rect 410 1176 412 1196
rect 416 1176 420 1196
rect 432 1156 434 1196
rect 438 1156 442 1196
rect 446 1156 448 1196
rect 503 1156 505 1196
rect 509 1176 511 1196
rect 523 1176 525 1196
rect 529 1176 531 1196
rect 543 1176 545 1196
rect 549 1176 551 1196
rect 589 1176 591 1196
rect 595 1176 597 1196
rect 609 1176 611 1196
rect 615 1176 617 1196
rect 509 1156 521 1176
rect 693 1156 695 1196
rect 699 1156 701 1196
rect 713 1156 715 1196
rect 719 1156 725 1196
rect 729 1156 731 1196
rect 781 1156 783 1196
rect 787 1156 789 1196
rect 801 1176 805 1196
rect 809 1176 811 1196
rect 863 1176 865 1196
rect 869 1176 871 1196
rect 883 1176 885 1196
rect 889 1176 891 1196
rect 943 1176 945 1196
rect 949 1176 951 1196
rect 1003 1176 1005 1196
rect 1009 1176 1011 1196
rect 1049 1176 1051 1196
rect 1055 1176 1057 1196
rect 1069 1176 1071 1196
rect 1075 1176 1077 1196
rect 1129 1176 1131 1196
rect 1135 1176 1137 1196
rect 1203 1176 1205 1196
rect 1209 1176 1211 1196
rect 1223 1176 1225 1196
rect 1229 1176 1231 1196
rect 1272 1156 1274 1196
rect 1278 1156 1282 1196
rect 1286 1156 1288 1196
rect 1300 1176 1304 1196
rect 1308 1176 1310 1196
rect 1373 1156 1375 1196
rect 1379 1176 1381 1196
rect 1393 1176 1395 1196
rect 1399 1176 1405 1196
rect 1409 1176 1413 1196
rect 1425 1176 1427 1196
rect 1431 1176 1437 1196
rect 1441 1176 1443 1196
rect 1455 1176 1459 1196
rect 1463 1176 1465 1196
rect 1503 1176 1505 1196
rect 1509 1176 1513 1196
rect 1517 1176 1519 1196
rect 1531 1176 1533 1196
rect 1537 1176 1543 1196
rect 1547 1176 1549 1196
rect 1561 1176 1565 1196
rect 1379 1156 1389 1176
rect 1552 1156 1565 1176
rect 1569 1156 1571 1196
rect 1623 1176 1625 1196
rect 1629 1176 1631 1196
rect 1671 1156 1673 1196
rect 1677 1156 1683 1196
rect 1687 1156 1689 1196
rect 1749 1176 1751 1196
rect 1755 1176 1757 1196
rect 1769 1176 1771 1196
rect 1775 1176 1777 1196
rect 1833 1156 1835 1196
rect 1839 1176 1841 1196
rect 1853 1176 1855 1196
rect 1859 1176 1865 1196
rect 1869 1176 1873 1196
rect 1885 1176 1887 1196
rect 1891 1176 1897 1196
rect 1901 1176 1903 1196
rect 1915 1176 1919 1196
rect 1923 1176 1925 1196
rect 1963 1176 1965 1196
rect 1969 1176 1973 1196
rect 1977 1176 1979 1196
rect 1991 1176 1993 1196
rect 1997 1176 2003 1196
rect 2007 1176 2009 1196
rect 2021 1176 2025 1196
rect 1839 1156 1849 1176
rect 2012 1156 2025 1176
rect 2029 1156 2031 1196
rect 2083 1176 2085 1196
rect 2089 1176 2091 1196
rect 2129 1176 2131 1196
rect 2135 1176 2137 1196
rect 2149 1176 2151 1196
rect 2155 1176 2157 1196
rect 2209 1176 2211 1196
rect 2215 1176 2217 1196
rect 2229 1176 2231 1196
rect 2235 1176 2237 1196
rect 2303 1176 2305 1196
rect 2309 1176 2311 1196
rect 2349 1156 2351 1196
rect 2355 1176 2359 1196
rect 2371 1176 2373 1196
rect 2377 1176 2383 1196
rect 2387 1176 2389 1196
rect 2401 1176 2403 1196
rect 2407 1176 2411 1196
rect 2415 1176 2417 1196
rect 2455 1176 2457 1196
rect 2461 1176 2465 1196
rect 2477 1176 2479 1196
rect 2483 1176 2489 1196
rect 2493 1176 2495 1196
rect 2507 1176 2511 1196
rect 2515 1176 2521 1196
rect 2525 1176 2527 1196
rect 2539 1176 2541 1196
rect 2355 1156 2368 1176
rect 2531 1156 2541 1176
rect 2545 1156 2547 1196
rect 2589 1176 2591 1196
rect 2595 1176 2597 1196
rect 2649 1156 2651 1196
rect 2655 1168 2657 1196
rect 2669 1168 2671 1196
rect 2655 1156 2671 1168
rect 2675 1156 2677 1196
rect 2689 1156 2691 1196
rect 2695 1156 2697 1196
rect 2749 1156 2751 1196
rect 2755 1166 2757 1196
rect 2769 1166 2771 1196
rect 2755 1156 2771 1166
rect 2775 1156 2777 1196
rect 2789 1156 2791 1196
rect 2795 1184 2811 1196
rect 2795 1156 2797 1184
rect 2809 1156 2811 1184
rect 2815 1156 2817 1196
rect 2869 1176 2871 1196
rect 2875 1176 2877 1196
rect 2889 1176 2891 1196
rect 2895 1176 2897 1196
rect 2971 1156 2973 1196
rect 2977 1156 2983 1196
rect 2987 1156 2989 1196
rect 3029 1156 3031 1196
rect 3035 1156 3041 1196
rect 3045 1156 3047 1196
rect 3059 1156 3061 1196
rect 3065 1156 3067 1196
rect 3129 1156 3131 1196
rect 3135 1168 3137 1196
rect 3149 1168 3151 1196
rect 3135 1156 3151 1168
rect 3155 1156 3157 1196
rect 3169 1156 3171 1196
rect 3175 1156 3177 1196
rect 3229 1176 3231 1196
rect 3235 1176 3237 1196
rect 3249 1176 3251 1196
rect 3255 1176 3257 1196
rect 3269 1176 3271 1196
rect 3259 1156 3271 1176
rect 3275 1156 3277 1196
rect 3351 1156 3353 1196
rect 3357 1156 3363 1196
rect 3367 1156 3369 1196
rect 3431 1156 3433 1196
rect 3437 1156 3443 1196
rect 3447 1156 3449 1196
rect 3491 1156 3493 1196
rect 3497 1156 3503 1196
rect 3507 1156 3509 1196
rect 3571 1156 3573 1196
rect 3577 1156 3583 1196
rect 3587 1156 3589 1196
rect 3649 1156 3651 1196
rect 3655 1168 3657 1196
rect 3669 1168 3671 1196
rect 3655 1156 3671 1168
rect 3675 1156 3677 1196
rect 3689 1156 3691 1196
rect 3695 1156 3697 1196
rect 3786 1138 3788 1196
rect 3774 1136 3788 1138
rect 3792 1136 3796 1196
rect 3800 1136 3804 1196
rect 3808 1136 3810 1196
rect 3852 1156 3854 1196
rect 3858 1156 3862 1196
rect 3866 1156 3868 1196
rect 3880 1176 3884 1196
rect 3888 1176 3890 1196
rect 3963 1176 3965 1196
rect 3969 1176 3971 1196
rect 4046 1138 4048 1196
rect 4034 1136 4048 1138
rect 4052 1136 4056 1196
rect 4060 1136 4064 1196
rect 4068 1136 4070 1196
rect 4112 1156 4114 1196
rect 4118 1156 4122 1196
rect 4126 1156 4128 1196
rect 4140 1176 4144 1196
rect 4148 1176 4150 1196
rect 4209 1176 4211 1196
rect 4215 1176 4217 1196
rect 4290 1176 4292 1196
rect 4296 1176 4300 1196
rect 4312 1156 4314 1196
rect 4318 1156 4322 1196
rect 4326 1156 4328 1196
rect 4383 1156 4385 1196
rect 4389 1156 4391 1196
rect 4403 1156 4405 1196
rect 4409 1168 4411 1196
rect 4423 1168 4425 1196
rect 4409 1156 4425 1168
rect 4429 1156 4431 1196
rect 4469 1156 4471 1196
rect 4475 1168 4477 1196
rect 4489 1168 4491 1196
rect 4475 1156 4491 1168
rect 4495 1156 4497 1196
rect 4509 1156 4511 1196
rect 4515 1156 4517 1196
rect 4569 1176 4571 1196
rect 4575 1176 4577 1196
rect 4589 1176 4591 1196
rect 4595 1176 4597 1196
rect 4671 1156 4673 1196
rect 4677 1156 4683 1196
rect 4687 1156 4689 1196
rect 4743 1176 4745 1196
rect 4749 1176 4751 1196
rect 33 744 35 784
rect 39 764 49 784
rect 212 764 225 784
rect 39 744 41 764
rect 53 744 55 764
rect 59 744 65 764
rect 69 744 73 764
rect 85 744 87 764
rect 91 744 97 764
rect 101 744 103 764
rect 115 744 119 764
rect 123 744 125 764
rect 163 744 165 764
rect 169 744 173 764
rect 177 744 179 764
rect 191 744 193 764
rect 197 744 203 764
rect 207 744 209 764
rect 221 744 225 764
rect 229 744 231 784
rect 271 744 273 784
rect 277 744 283 784
rect 287 744 289 784
rect 363 744 365 784
rect 369 744 371 784
rect 383 744 385 784
rect 389 772 405 784
rect 389 744 391 772
rect 403 744 405 772
rect 409 744 411 784
rect 453 744 455 784
rect 459 764 469 784
rect 632 764 645 784
rect 459 744 461 764
rect 473 744 475 764
rect 479 744 485 764
rect 489 744 493 764
rect 505 744 507 764
rect 511 744 517 764
rect 521 744 523 764
rect 535 744 539 764
rect 543 744 545 764
rect 583 744 585 764
rect 589 744 593 764
rect 597 744 599 764
rect 611 744 613 764
rect 617 744 623 764
rect 627 744 629 764
rect 641 744 645 764
rect 649 744 651 784
rect 691 744 693 784
rect 697 744 703 784
rect 707 744 709 784
rect 783 744 785 784
rect 789 744 791 784
rect 803 744 805 784
rect 809 772 825 784
rect 809 744 811 772
rect 823 744 825 772
rect 829 744 831 784
rect 883 744 885 784
rect 889 744 891 784
rect 903 744 905 784
rect 909 772 925 784
rect 909 744 911 772
rect 923 744 925 772
rect 929 744 931 784
rect 983 744 985 764
rect 989 744 991 764
rect 1043 744 1045 764
rect 1049 744 1051 764
rect 1063 744 1065 764
rect 1069 744 1071 764
rect 1109 744 1111 764
rect 1115 744 1117 764
rect 1129 744 1131 764
rect 1135 744 1137 764
rect 1211 744 1213 784
rect 1217 744 1223 784
rect 1227 744 1229 784
rect 1291 744 1293 784
rect 1297 744 1303 784
rect 1307 744 1309 784
rect 1371 744 1373 784
rect 1377 744 1383 784
rect 1387 744 1389 784
rect 1450 744 1452 764
rect 1456 744 1460 764
rect 1472 744 1474 784
rect 1478 744 1482 784
rect 1486 744 1488 784
rect 1553 744 1555 784
rect 1559 744 1561 784
rect 1573 744 1575 784
rect 1579 744 1585 784
rect 1589 744 1591 784
rect 1632 744 1634 784
rect 1638 744 1642 784
rect 1646 744 1648 784
rect 1660 744 1664 764
rect 1668 744 1670 764
rect 1729 744 1731 784
rect 1735 744 1737 784
rect 1749 744 1751 784
rect 1755 744 1757 784
rect 1769 744 1771 784
rect 1775 744 1777 784
rect 1789 744 1791 784
rect 1795 744 1797 784
rect 1809 744 1811 784
rect 1815 744 1817 784
rect 1829 744 1831 784
rect 1835 744 1837 784
rect 1849 744 1851 784
rect 1855 744 1857 784
rect 1869 744 1871 784
rect 1875 744 1877 784
rect 1951 744 1953 784
rect 1957 744 1963 784
rect 1967 744 1969 784
rect 2023 744 2025 764
rect 2029 744 2031 764
rect 2043 744 2045 764
rect 2049 744 2051 764
rect 2089 744 2091 784
rect 2095 772 2111 784
rect 2095 744 2097 772
rect 2109 744 2111 772
rect 2115 744 2117 784
rect 2129 744 2131 784
rect 2135 744 2137 784
rect 2189 744 2191 784
rect 2195 772 2211 784
rect 2195 744 2197 772
rect 2209 744 2211 772
rect 2215 744 2217 784
rect 2229 744 2231 784
rect 2235 744 2237 784
rect 2289 744 2291 784
rect 2295 772 2311 784
rect 2295 744 2297 772
rect 2309 744 2311 772
rect 2315 744 2317 784
rect 2329 744 2331 784
rect 2335 744 2337 784
rect 2391 744 2393 784
rect 2397 744 2403 784
rect 2407 744 2409 784
rect 2483 744 2485 764
rect 2489 744 2491 764
rect 2529 744 2531 784
rect 2535 764 2548 784
rect 2711 764 2721 784
rect 2535 744 2539 764
rect 2551 744 2553 764
rect 2557 744 2563 764
rect 2567 744 2569 764
rect 2581 744 2583 764
rect 2587 744 2591 764
rect 2595 744 2597 764
rect 2635 744 2637 764
rect 2641 744 2645 764
rect 2657 744 2659 764
rect 2663 744 2669 764
rect 2673 744 2675 764
rect 2687 744 2691 764
rect 2695 744 2701 764
rect 2705 744 2707 764
rect 2719 744 2721 764
rect 2725 744 2727 784
rect 2783 744 2785 784
rect 2789 744 2791 784
rect 2803 744 2805 784
rect 2809 772 2825 784
rect 2809 744 2811 772
rect 2823 744 2825 772
rect 2829 744 2831 784
rect 2883 744 2885 764
rect 2889 744 2891 764
rect 2929 744 2931 764
rect 2935 744 2937 764
rect 2990 744 2992 804
rect 2996 744 3000 804
rect 3004 744 3008 804
rect 3012 802 3026 804
rect 3012 744 3014 802
rect 3089 744 3091 764
rect 3095 744 3097 764
rect 3171 744 3173 784
rect 3177 744 3183 784
rect 3187 744 3189 784
rect 3259 764 3271 784
rect 3229 744 3231 764
rect 3235 744 3237 764
rect 3249 744 3251 764
rect 3255 744 3257 764
rect 3269 744 3271 764
rect 3275 744 3277 784
rect 3331 744 3333 784
rect 3337 744 3343 784
rect 3347 744 3349 784
rect 3411 744 3413 784
rect 3417 744 3423 784
rect 3427 744 3429 784
rect 3674 802 3688 804
rect 3503 744 3505 764
rect 3509 744 3511 764
rect 3523 744 3525 764
rect 3529 744 3531 764
rect 3571 744 3573 784
rect 3577 744 3583 784
rect 3587 744 3589 784
rect 3686 744 3688 802
rect 3692 744 3696 804
rect 3700 744 3704 804
rect 3708 744 3710 804
rect 3774 802 3788 804
rect 3786 744 3788 802
rect 3792 744 3796 804
rect 3800 744 3804 804
rect 3808 744 3810 804
rect 3954 802 3968 804
rect 3851 744 3853 784
rect 3857 744 3863 784
rect 3867 744 3869 784
rect 3966 744 3968 802
rect 3972 744 3976 804
rect 3980 744 3984 804
rect 3988 744 3990 804
rect 4043 744 4045 764
rect 4049 744 4051 764
rect 4103 744 4105 784
rect 4109 744 4111 784
rect 4123 744 4125 784
rect 4129 772 4145 784
rect 4129 744 4131 772
rect 4143 744 4145 772
rect 4149 744 4151 784
rect 4203 744 4205 784
rect 4209 744 4211 784
rect 4223 744 4225 784
rect 4229 772 4245 784
rect 4229 744 4231 772
rect 4243 744 4245 772
rect 4249 744 4251 784
rect 4310 744 4312 764
rect 4316 744 4320 764
rect 4332 744 4334 784
rect 4338 744 4342 784
rect 4346 744 4348 784
rect 4390 744 4392 804
rect 4396 744 4400 804
rect 4404 744 4408 804
rect 4412 802 4426 804
rect 4412 744 4414 802
rect 4514 802 4528 804
rect 4526 744 4528 802
rect 4532 744 4536 804
rect 4540 744 4544 804
rect 4548 744 4550 804
rect 4610 744 4612 764
rect 4616 744 4620 764
rect 4632 744 4634 784
rect 4638 744 4642 784
rect 4646 744 4648 784
rect 4690 744 4692 804
rect 4696 744 4700 804
rect 4704 744 4708 804
rect 4712 802 4726 804
rect 4712 744 4714 802
rect 33 676 35 716
rect 39 696 41 716
rect 53 696 55 716
rect 59 696 65 716
rect 69 696 73 716
rect 85 696 87 716
rect 91 696 97 716
rect 101 696 103 716
rect 115 696 119 716
rect 123 696 125 716
rect 163 696 165 716
rect 169 696 173 716
rect 177 696 179 716
rect 191 696 193 716
rect 197 696 203 716
rect 207 696 209 716
rect 221 696 225 716
rect 39 676 49 696
rect 212 676 225 696
rect 229 676 231 716
rect 269 696 271 716
rect 275 696 277 716
rect 329 676 331 716
rect 335 688 337 716
rect 349 688 351 716
rect 335 676 351 688
rect 355 676 357 716
rect 369 676 371 716
rect 375 676 377 716
rect 431 676 433 716
rect 437 676 443 716
rect 447 676 449 716
rect 509 696 511 716
rect 515 696 519 716
rect 531 676 533 716
rect 537 676 539 716
rect 603 696 605 716
rect 609 696 611 716
rect 649 676 651 716
rect 655 696 659 716
rect 671 696 673 716
rect 677 696 683 716
rect 687 696 689 716
rect 701 696 703 716
rect 707 696 711 716
rect 715 696 717 716
rect 755 696 757 716
rect 761 696 765 716
rect 777 696 779 716
rect 783 696 789 716
rect 793 696 795 716
rect 807 696 811 716
rect 815 696 821 716
rect 825 696 827 716
rect 839 696 841 716
rect 655 676 668 696
rect 831 676 841 696
rect 845 676 847 716
rect 889 676 891 716
rect 895 688 897 716
rect 909 688 911 716
rect 895 676 911 688
rect 915 676 917 716
rect 929 676 931 716
rect 935 676 937 716
rect 1003 696 1005 716
rect 1009 696 1011 716
rect 1023 696 1025 716
rect 1029 696 1031 716
rect 1069 696 1071 716
rect 1075 696 1077 716
rect 1089 696 1091 716
rect 1095 696 1097 716
rect 1109 696 1111 716
rect 1099 676 1111 696
rect 1115 676 1117 716
rect 1183 676 1185 716
rect 1189 676 1191 716
rect 1203 676 1205 716
rect 1209 688 1211 716
rect 1223 688 1225 716
rect 1209 676 1225 688
rect 1229 676 1231 716
rect 1293 676 1295 716
rect 1299 676 1301 716
rect 1313 676 1315 716
rect 1319 676 1325 716
rect 1329 676 1331 716
rect 1369 696 1371 716
rect 1375 696 1377 716
rect 1389 696 1391 716
rect 1395 696 1397 716
rect 1449 696 1451 716
rect 1455 696 1459 716
rect 1471 676 1473 716
rect 1477 676 1479 716
rect 1533 676 1535 716
rect 1539 696 1541 716
rect 1553 696 1555 716
rect 1559 696 1565 716
rect 1569 696 1573 716
rect 1585 696 1587 716
rect 1591 696 1597 716
rect 1601 696 1603 716
rect 1615 696 1619 716
rect 1623 696 1625 716
rect 1663 696 1665 716
rect 1669 696 1673 716
rect 1677 696 1679 716
rect 1691 696 1693 716
rect 1697 696 1703 716
rect 1707 696 1709 716
rect 1721 696 1725 716
rect 1539 676 1549 696
rect 1712 676 1725 696
rect 1729 676 1731 716
rect 1769 696 1771 716
rect 1775 696 1779 716
rect 1791 676 1793 716
rect 1797 676 1799 716
rect 1863 696 1865 716
rect 1869 696 1871 716
rect 1883 696 1885 716
rect 1889 696 1891 716
rect 1943 696 1945 716
rect 1949 696 1951 716
rect 1963 696 1965 716
rect 1969 696 1971 716
rect 2023 696 2025 716
rect 2029 696 2031 716
rect 2069 696 2071 716
rect 2075 696 2077 716
rect 2089 696 2091 716
rect 2095 696 2097 716
rect 2149 676 2151 716
rect 2155 696 2159 716
rect 2171 696 2173 716
rect 2177 696 2183 716
rect 2187 696 2189 716
rect 2201 696 2203 716
rect 2207 696 2211 716
rect 2215 696 2217 716
rect 2255 696 2257 716
rect 2261 696 2265 716
rect 2277 696 2279 716
rect 2283 696 2289 716
rect 2293 696 2295 716
rect 2307 696 2311 716
rect 2315 696 2321 716
rect 2325 696 2327 716
rect 2339 696 2341 716
rect 2155 676 2168 696
rect 2331 676 2341 696
rect 2345 676 2347 716
rect 2392 676 2394 716
rect 2398 676 2402 716
rect 2406 676 2408 716
rect 2420 676 2422 716
rect 2426 676 2430 716
rect 2434 676 2436 716
rect 2523 676 2525 716
rect 2529 696 2531 716
rect 2543 696 2545 716
rect 2549 696 2551 716
rect 2563 696 2565 716
rect 2569 696 2571 716
rect 2630 696 2632 716
rect 2636 696 2640 716
rect 2529 676 2541 696
rect 2652 676 2654 716
rect 2658 676 2662 716
rect 2666 676 2668 716
rect 2730 696 2732 716
rect 2736 696 2740 716
rect 2752 676 2754 716
rect 2758 676 2762 716
rect 2766 676 2768 716
rect 2809 696 2811 716
rect 2815 696 2817 716
rect 2883 676 2885 716
rect 2889 676 2891 716
rect 2903 676 2905 716
rect 2909 688 2911 716
rect 2923 688 2925 716
rect 2909 676 2925 688
rect 2929 676 2931 716
rect 2969 676 2971 716
rect 2975 688 2977 716
rect 2989 688 2991 716
rect 2975 676 2991 688
rect 2995 676 2997 716
rect 3009 676 3011 716
rect 3015 676 3017 716
rect 3071 676 3073 716
rect 3077 676 3083 716
rect 3087 676 3089 716
rect 3163 696 3165 716
rect 3169 696 3171 716
rect 3209 696 3211 716
rect 3215 696 3217 716
rect 3306 658 3308 716
rect 3294 656 3308 658
rect 3312 656 3316 716
rect 3320 656 3324 716
rect 3328 656 3330 716
rect 3383 696 3385 716
rect 3389 696 3391 716
rect 3403 696 3405 716
rect 3409 696 3411 716
rect 3449 676 3451 716
rect 3455 688 3457 716
rect 3469 688 3471 716
rect 3455 676 3471 688
rect 3475 676 3477 716
rect 3489 676 3491 716
rect 3495 676 3497 716
rect 3552 676 3554 716
rect 3558 676 3562 716
rect 3566 676 3568 716
rect 3580 696 3584 716
rect 3588 696 3590 716
rect 3670 696 3672 716
rect 3676 696 3680 716
rect 3692 676 3694 716
rect 3698 676 3702 716
rect 3706 676 3708 716
rect 3784 676 3786 716
rect 3790 676 3794 716
rect 3798 676 3800 716
rect 3812 676 3814 716
rect 3818 676 3822 716
rect 3826 676 3828 716
rect 3906 658 3908 716
rect 3894 656 3908 658
rect 3912 656 3916 716
rect 3920 656 3924 716
rect 3928 656 3930 716
rect 4006 658 4008 716
rect 3994 656 4008 658
rect 4012 656 4016 716
rect 4020 656 4024 716
rect 4028 656 4030 716
rect 4069 696 4071 716
rect 4075 696 4077 716
rect 4130 656 4132 716
rect 4136 656 4140 716
rect 4144 656 4148 716
rect 4152 658 4154 716
rect 4152 656 4166 658
rect 4230 656 4232 716
rect 4236 656 4240 716
rect 4244 656 4248 716
rect 4252 658 4254 716
rect 4252 656 4266 658
rect 4366 658 4368 716
rect 4354 656 4368 658
rect 4372 656 4376 716
rect 4380 656 4384 716
rect 4388 656 4390 716
rect 4466 658 4468 716
rect 4454 656 4468 658
rect 4472 656 4476 716
rect 4480 656 4484 716
rect 4488 656 4490 716
rect 4529 696 4531 716
rect 4535 696 4537 716
rect 4603 676 4605 716
rect 4609 676 4611 716
rect 4623 676 4625 716
rect 4629 688 4631 716
rect 4643 688 4645 716
rect 4629 676 4645 688
rect 4649 676 4651 716
rect 4689 676 4691 716
rect 4695 688 4697 716
rect 4709 688 4711 716
rect 4695 676 4711 688
rect 4715 676 4717 716
rect 4729 676 4731 716
rect 4735 676 4737 716
rect 33 264 35 304
rect 39 284 49 304
rect 212 284 225 304
rect 39 264 41 284
rect 53 264 55 284
rect 59 264 65 284
rect 69 264 73 284
rect 85 264 87 284
rect 91 264 97 284
rect 101 264 103 284
rect 115 264 119 284
rect 123 264 125 284
rect 163 264 165 284
rect 169 264 173 284
rect 177 264 179 284
rect 191 264 193 284
rect 197 264 203 284
rect 207 264 209 284
rect 221 264 225 284
rect 229 264 231 304
rect 271 264 273 304
rect 277 264 283 304
rect 287 264 289 304
rect 363 264 365 304
rect 369 264 371 304
rect 383 264 385 304
rect 389 292 405 304
rect 389 264 391 292
rect 403 264 405 292
rect 409 264 411 304
rect 449 264 451 284
rect 455 264 457 284
rect 511 264 513 304
rect 517 264 523 304
rect 527 264 529 304
rect 603 264 605 304
rect 609 264 611 304
rect 623 264 625 304
rect 629 292 645 304
rect 629 264 631 292
rect 643 264 645 292
rect 649 264 651 304
rect 689 264 691 304
rect 695 292 711 304
rect 695 264 697 292
rect 709 264 711 292
rect 715 264 717 304
rect 729 264 731 304
rect 735 264 737 304
rect 789 264 791 304
rect 795 292 811 304
rect 795 264 797 292
rect 809 264 811 292
rect 815 264 817 304
rect 829 264 831 304
rect 835 264 837 304
rect 903 264 905 304
rect 909 264 911 304
rect 923 264 925 304
rect 929 292 945 304
rect 929 264 931 292
rect 943 264 945 292
rect 949 264 951 304
rect 989 264 991 284
rect 995 264 997 284
rect 1051 264 1053 304
rect 1057 264 1063 304
rect 1067 264 1069 304
rect 1150 264 1152 284
rect 1156 264 1160 284
rect 1172 264 1174 304
rect 1178 264 1182 304
rect 1186 264 1188 304
rect 1243 264 1245 284
rect 1249 264 1251 284
rect 1303 264 1305 304
rect 1309 264 1311 304
rect 1323 264 1325 304
rect 1329 292 1345 304
rect 1329 264 1331 292
rect 1343 264 1345 292
rect 1349 264 1351 304
rect 1403 264 1405 284
rect 1409 264 1411 284
rect 1423 264 1425 284
rect 1429 264 1431 284
rect 1469 264 1471 304
rect 1475 292 1491 304
rect 1475 264 1477 292
rect 1489 264 1491 292
rect 1495 264 1497 304
rect 1509 264 1511 304
rect 1515 264 1517 304
rect 1571 264 1573 304
rect 1577 264 1583 304
rect 1587 264 1589 304
rect 1649 264 1651 304
rect 1655 284 1668 304
rect 1831 284 1841 304
rect 1655 264 1659 284
rect 1671 264 1673 284
rect 1677 264 1683 284
rect 1687 264 1689 284
rect 1701 264 1703 284
rect 1707 264 1711 284
rect 1715 264 1717 284
rect 1755 264 1757 284
rect 1761 264 1765 284
rect 1777 264 1779 284
rect 1783 264 1789 284
rect 1793 264 1795 284
rect 1807 264 1811 284
rect 1815 264 1821 284
rect 1825 264 1827 284
rect 1839 264 1841 284
rect 1845 264 1847 304
rect 1911 264 1913 304
rect 1917 264 1923 304
rect 1927 264 1929 304
rect 1983 264 1985 304
rect 1989 264 1991 304
rect 2003 264 2005 304
rect 2009 292 2025 304
rect 2009 264 2011 292
rect 2023 264 2025 292
rect 2029 264 2031 304
rect 2073 264 2075 304
rect 2079 284 2089 304
rect 2252 284 2265 304
rect 2079 264 2081 284
rect 2093 264 2095 284
rect 2099 264 2105 284
rect 2109 264 2113 284
rect 2125 264 2127 284
rect 2131 264 2137 284
rect 2141 264 2143 284
rect 2155 264 2159 284
rect 2163 264 2165 284
rect 2203 264 2205 284
rect 2209 264 2213 284
rect 2217 264 2219 284
rect 2231 264 2233 284
rect 2237 264 2243 284
rect 2247 264 2249 284
rect 2261 264 2265 284
rect 2269 264 2271 304
rect 2323 264 2325 284
rect 2329 264 2331 284
rect 2369 264 2371 284
rect 2375 264 2377 284
rect 2389 264 2391 284
rect 2395 264 2397 284
rect 2449 264 2451 284
rect 2455 264 2457 284
rect 2531 264 2533 304
rect 2537 264 2543 304
rect 2547 264 2549 304
rect 2589 264 2591 304
rect 2595 284 2608 304
rect 2771 284 2781 304
rect 2595 264 2599 284
rect 2611 264 2613 284
rect 2617 264 2623 284
rect 2627 264 2629 284
rect 2641 264 2643 284
rect 2647 264 2651 284
rect 2655 264 2657 284
rect 2695 264 2697 284
rect 2701 264 2705 284
rect 2717 264 2719 284
rect 2723 264 2729 284
rect 2733 264 2735 284
rect 2747 264 2751 284
rect 2755 264 2761 284
rect 2765 264 2767 284
rect 2779 264 2781 284
rect 2785 264 2787 304
rect 2831 264 2833 304
rect 2837 264 2843 304
rect 2847 264 2849 304
rect 2912 264 2914 304
rect 2918 264 2922 304
rect 2926 264 2928 304
rect 2940 264 2942 304
rect 2946 264 2950 304
rect 2954 264 2956 304
rect 3194 322 3208 324
rect 3029 264 3031 284
rect 3035 264 3037 284
rect 3049 264 3051 284
rect 3055 264 3057 284
rect 3109 264 3111 284
rect 3115 264 3117 284
rect 3206 264 3208 322
rect 3212 264 3216 324
rect 3220 264 3224 324
rect 3228 264 3230 324
rect 3294 322 3308 324
rect 3306 264 3308 322
rect 3312 264 3316 324
rect 3320 264 3324 324
rect 3328 264 3330 324
rect 3369 264 3371 304
rect 3375 292 3391 304
rect 3375 264 3377 292
rect 3389 264 3391 292
rect 3395 264 3397 304
rect 3409 264 3411 304
rect 3415 264 3417 304
rect 3483 264 3485 284
rect 3489 264 3491 284
rect 3531 264 3533 304
rect 3537 264 3543 304
rect 3547 264 3549 304
rect 3611 264 3613 304
rect 3617 264 3623 304
rect 3627 264 3629 304
rect 3689 264 3691 304
rect 3695 292 3711 304
rect 3695 264 3697 292
rect 3709 264 3711 292
rect 3715 264 3717 304
rect 3729 264 3731 304
rect 3735 264 3737 304
rect 3803 264 3805 284
rect 3809 264 3811 284
rect 3823 264 3825 284
rect 3829 264 3831 284
rect 3883 264 3885 284
rect 3889 264 3891 284
rect 3903 264 3905 284
rect 3909 264 3911 284
rect 3949 264 3951 304
rect 3955 264 3961 304
rect 3965 264 3967 304
rect 3979 264 3981 304
rect 3985 264 3987 304
rect 4254 322 4268 324
rect 4049 264 4051 284
rect 4055 264 4057 284
rect 4069 264 4071 284
rect 4075 264 4077 284
rect 4150 264 4152 284
rect 4156 264 4160 284
rect 4172 264 4174 304
rect 4178 264 4182 304
rect 4186 264 4188 304
rect 4266 264 4268 322
rect 4272 264 4276 324
rect 4280 264 4284 324
rect 4288 264 4290 324
rect 4332 264 4334 304
rect 4338 264 4342 304
rect 4346 264 4348 304
rect 4360 264 4364 284
rect 4368 264 4370 284
rect 4429 264 4431 284
rect 4435 264 4437 284
rect 4503 264 4505 304
rect 4509 264 4511 304
rect 4523 264 4525 304
rect 4529 292 4545 304
rect 4529 264 4531 292
rect 4543 264 4545 292
rect 4549 264 4551 304
rect 4589 264 4591 284
rect 4595 264 4597 284
rect 4649 264 4651 284
rect 4655 264 4657 284
rect 4709 264 4711 284
rect 4715 264 4717 284
rect 33 196 35 236
rect 39 216 41 236
rect 53 216 55 236
rect 59 216 65 236
rect 69 216 73 236
rect 85 216 87 236
rect 91 216 97 236
rect 101 216 103 236
rect 115 216 119 236
rect 123 216 125 236
rect 163 216 165 236
rect 169 216 173 236
rect 177 216 179 236
rect 191 216 193 236
rect 197 216 203 236
rect 207 216 209 236
rect 221 216 225 236
rect 39 196 49 216
rect 212 196 225 216
rect 229 196 231 236
rect 272 196 274 236
rect 278 196 282 236
rect 286 196 288 236
rect 300 196 302 236
rect 306 196 310 236
rect 314 196 316 236
rect 389 216 391 236
rect 395 216 397 236
rect 409 216 411 236
rect 415 216 417 236
rect 470 176 472 236
rect 476 176 480 236
rect 484 176 488 236
rect 492 178 494 236
rect 583 196 585 236
rect 589 216 591 236
rect 603 216 605 236
rect 609 216 611 236
rect 623 216 625 236
rect 629 216 631 236
rect 690 216 692 236
rect 696 216 700 236
rect 589 196 601 216
rect 492 176 506 178
rect 712 196 714 236
rect 718 196 722 236
rect 726 196 728 236
rect 769 196 771 236
rect 775 216 779 236
rect 791 216 793 236
rect 797 216 803 236
rect 807 216 809 236
rect 821 216 823 236
rect 827 216 831 236
rect 835 216 837 236
rect 875 216 877 236
rect 881 216 885 236
rect 897 216 899 236
rect 903 216 909 236
rect 913 216 915 236
rect 927 216 931 236
rect 935 216 941 236
rect 945 216 947 236
rect 959 216 961 236
rect 775 196 788 216
rect 951 196 961 216
rect 965 196 967 236
rect 1023 196 1025 236
rect 1029 196 1031 236
rect 1043 196 1045 236
rect 1049 208 1051 236
rect 1063 208 1065 236
rect 1049 196 1065 208
rect 1069 196 1071 236
rect 1123 216 1125 236
rect 1129 216 1131 236
rect 1183 216 1185 236
rect 1189 216 1191 236
rect 1203 216 1205 236
rect 1209 216 1211 236
rect 1263 216 1265 236
rect 1269 216 1271 236
rect 1323 196 1325 236
rect 1329 196 1331 236
rect 1343 196 1345 236
rect 1349 208 1351 236
rect 1363 208 1365 236
rect 1349 196 1365 208
rect 1369 196 1371 236
rect 1423 216 1425 236
rect 1429 216 1431 236
rect 1483 216 1485 236
rect 1489 216 1491 236
rect 1529 216 1531 236
rect 1535 216 1537 236
rect 1549 216 1551 236
rect 1555 216 1557 236
rect 1630 216 1632 236
rect 1636 216 1640 236
rect 1652 196 1654 236
rect 1658 196 1662 236
rect 1666 196 1668 236
rect 1713 196 1715 236
rect 1719 216 1721 236
rect 1733 216 1735 236
rect 1739 216 1745 236
rect 1749 216 1753 236
rect 1765 216 1767 236
rect 1771 216 1777 236
rect 1781 216 1783 236
rect 1795 216 1799 236
rect 1803 216 1805 236
rect 1843 216 1845 236
rect 1849 216 1853 236
rect 1857 216 1859 236
rect 1871 216 1873 236
rect 1877 216 1883 236
rect 1887 216 1889 236
rect 1901 216 1905 236
rect 1719 196 1729 216
rect 1892 196 1905 216
rect 1909 196 1911 236
rect 1963 196 1965 236
rect 1969 196 1971 236
rect 1983 196 1985 236
rect 1989 208 1991 236
rect 2003 208 2005 236
rect 1989 196 2005 208
rect 2009 196 2011 236
rect 2049 216 2051 236
rect 2055 216 2057 236
rect 2109 216 2111 236
rect 2115 216 2117 236
rect 2129 216 2131 236
rect 2135 216 2137 236
rect 2189 216 2191 236
rect 2195 216 2197 236
rect 2209 216 2211 236
rect 2215 216 2217 236
rect 2283 216 2285 236
rect 2289 216 2291 236
rect 2303 216 2305 236
rect 2309 216 2311 236
rect 2349 216 2351 236
rect 2355 216 2357 236
rect 2369 216 2371 236
rect 2375 216 2377 236
rect 2443 216 2445 236
rect 2449 216 2451 236
rect 2489 196 2491 236
rect 2495 216 2499 236
rect 2511 216 2513 236
rect 2517 216 2523 236
rect 2527 216 2529 236
rect 2541 216 2543 236
rect 2547 216 2551 236
rect 2555 216 2557 236
rect 2595 216 2597 236
rect 2601 216 2605 236
rect 2617 216 2619 236
rect 2623 216 2629 236
rect 2633 216 2635 236
rect 2647 216 2651 236
rect 2655 216 2661 236
rect 2665 216 2667 236
rect 2679 216 2681 236
rect 2495 196 2508 216
rect 2671 196 2681 216
rect 2685 196 2687 236
rect 2729 196 2731 236
rect 2735 216 2739 236
rect 2751 216 2753 236
rect 2757 216 2763 236
rect 2767 216 2769 236
rect 2781 216 2783 236
rect 2787 216 2791 236
rect 2795 216 2797 236
rect 2835 216 2837 236
rect 2841 216 2845 236
rect 2857 216 2859 236
rect 2863 216 2869 236
rect 2873 216 2875 236
rect 2887 216 2891 236
rect 2895 216 2901 236
rect 2905 216 2907 236
rect 2919 216 2921 236
rect 2735 196 2748 216
rect 2911 196 2921 216
rect 2925 196 2927 236
rect 2969 196 2971 236
rect 2975 206 2977 236
rect 2989 206 2991 236
rect 2975 196 2991 206
rect 2995 196 2997 236
rect 3009 196 3011 236
rect 3015 224 3031 236
rect 3015 196 3017 224
rect 3029 196 3031 224
rect 3035 196 3037 236
rect 3103 196 3105 236
rect 3109 216 3111 236
rect 3123 216 3125 236
rect 3129 216 3131 236
rect 3143 216 3145 236
rect 3149 216 3151 236
rect 3109 196 3121 216
rect 3189 196 3191 236
rect 3195 208 3197 236
rect 3209 208 3211 236
rect 3195 196 3211 208
rect 3215 196 3217 236
rect 3229 196 3231 236
rect 3235 196 3237 236
rect 3303 216 3305 236
rect 3309 216 3311 236
rect 3351 196 3353 236
rect 3357 196 3363 236
rect 3367 196 3369 236
rect 3466 178 3468 236
rect 3454 176 3468 178
rect 3472 176 3476 236
rect 3480 176 3484 236
rect 3488 176 3490 236
rect 3543 216 3545 236
rect 3549 216 3551 236
rect 3610 216 3612 236
rect 3616 216 3620 236
rect 3632 196 3634 236
rect 3638 196 3642 236
rect 3646 196 3648 236
rect 3703 216 3705 236
rect 3709 216 3711 236
rect 3723 216 3725 236
rect 3729 216 3731 236
rect 3769 216 3771 236
rect 3775 216 3777 236
rect 3829 196 3831 236
rect 3835 208 3837 236
rect 3849 208 3851 236
rect 3835 196 3851 208
rect 3855 196 3857 236
rect 3869 196 3871 236
rect 3875 196 3877 236
rect 3929 216 3931 236
rect 3935 216 3937 236
rect 3949 216 3951 236
rect 3955 216 3957 236
rect 4046 178 4048 236
rect 4034 176 4048 178
rect 4052 176 4056 236
rect 4060 176 4064 236
rect 4068 176 4070 236
rect 4111 196 4113 236
rect 4117 196 4123 236
rect 4127 196 4129 236
rect 4226 178 4228 236
rect 4214 176 4228 178
rect 4232 176 4236 236
rect 4240 176 4244 236
rect 4248 176 4250 236
rect 4311 196 4313 236
rect 4317 196 4323 236
rect 4327 196 4329 236
rect 4406 178 4408 236
rect 4394 176 4408 178
rect 4412 176 4416 236
rect 4420 176 4424 236
rect 4428 176 4430 236
rect 4471 196 4473 236
rect 4477 196 4483 236
rect 4487 196 4489 236
rect 4550 176 4552 236
rect 4556 176 4560 236
rect 4564 176 4568 236
rect 4572 178 4574 236
rect 4670 216 4672 236
rect 4676 216 4680 236
rect 4572 176 4586 178
rect 4692 196 4694 236
rect 4698 196 4702 236
rect 4706 196 4708 236
<< pdiffusion >>
rect 41 4344 43 4424
rect 47 4344 49 4424
rect 61 4344 65 4384
rect 69 4344 71 4384
rect 123 4344 125 4384
rect 129 4344 131 4384
rect 143 4344 145 4384
rect 149 4344 151 4384
rect 208 4344 210 4384
rect 214 4344 218 4384
rect 230 4344 232 4424
rect 236 4344 240 4424
rect 244 4344 246 4424
rect 289 4344 291 4384
rect 295 4344 299 4384
rect 311 4344 313 4424
rect 317 4344 319 4424
rect 395 4344 397 4424
rect 401 4344 405 4424
rect 409 4344 411 4424
rect 475 4344 477 4424
rect 481 4344 485 4424
rect 489 4344 491 4424
rect 529 4344 531 4384
rect 535 4344 539 4384
rect 551 4344 553 4424
rect 557 4344 559 4424
rect 623 4344 625 4384
rect 629 4344 631 4384
rect 669 4344 671 4424
rect 675 4344 679 4424
rect 683 4344 685 4424
rect 749 4344 751 4384
rect 755 4344 757 4384
rect 809 4344 811 4424
rect 815 4364 824 4424
rect 992 4384 1001 4424
rect 850 4364 861 4384
rect 815 4344 817 4364
rect 829 4344 833 4364
rect 837 4344 841 4364
rect 845 4344 847 4364
rect 859 4344 861 4364
rect 865 4344 869 4384
rect 873 4344 875 4384
rect 913 4344 915 4384
rect 919 4344 921 4384
rect 933 4344 935 4384
rect 939 4344 947 4384
rect 951 4344 953 4384
rect 965 4344 967 4384
rect 971 4344 981 4384
rect 985 4344 987 4384
rect 999 4344 1001 4384
rect 1005 4344 1007 4424
rect 1054 4344 1056 4424
rect 1060 4344 1064 4424
rect 1068 4344 1070 4424
rect 1082 4344 1086 4384
rect 1090 4344 1092 4384
rect 1149 4344 1151 4424
rect 1155 4364 1164 4424
rect 1332 4384 1341 4424
rect 1190 4364 1201 4384
rect 1155 4344 1157 4364
rect 1169 4344 1173 4364
rect 1177 4344 1181 4364
rect 1185 4344 1187 4364
rect 1199 4344 1201 4364
rect 1205 4344 1209 4384
rect 1213 4344 1215 4384
rect 1253 4344 1255 4384
rect 1259 4344 1261 4384
rect 1273 4344 1275 4384
rect 1279 4344 1287 4384
rect 1291 4344 1293 4384
rect 1305 4344 1307 4384
rect 1311 4344 1321 4384
rect 1325 4344 1327 4384
rect 1339 4344 1341 4384
rect 1345 4344 1347 4424
rect 1394 4344 1396 4424
rect 1400 4344 1404 4424
rect 1408 4344 1410 4424
rect 1422 4344 1426 4384
rect 1430 4344 1432 4384
rect 1493 4344 1495 4424
rect 1499 4384 1508 4424
rect 1499 4344 1501 4384
rect 1513 4344 1515 4384
rect 1519 4344 1529 4384
rect 1533 4344 1535 4384
rect 1547 4344 1549 4384
rect 1553 4344 1561 4384
rect 1565 4344 1567 4384
rect 1579 4344 1581 4384
rect 1585 4344 1587 4384
rect 1625 4344 1627 4384
rect 1631 4344 1635 4384
rect 1639 4364 1650 4384
rect 1676 4364 1685 4424
rect 1639 4344 1641 4364
rect 1653 4344 1655 4364
rect 1659 4344 1663 4364
rect 1667 4344 1671 4364
rect 1683 4344 1685 4364
rect 1689 4344 1691 4424
rect 1729 4344 1731 4384
rect 1735 4344 1737 4384
rect 1749 4344 1751 4384
rect 1755 4344 1757 4384
rect 1809 4344 1811 4424
rect 1815 4364 1824 4424
rect 1992 4384 2001 4424
rect 1850 4364 1861 4384
rect 1815 4344 1817 4364
rect 1829 4344 1833 4364
rect 1837 4344 1841 4364
rect 1845 4344 1847 4364
rect 1859 4344 1861 4364
rect 1865 4344 1869 4384
rect 1873 4344 1875 4384
rect 1913 4344 1915 4384
rect 1919 4344 1921 4384
rect 1933 4344 1935 4384
rect 1939 4344 1947 4384
rect 1951 4344 1953 4384
rect 1965 4344 1967 4384
rect 1971 4344 1981 4384
rect 1985 4344 1987 4384
rect 1999 4344 2001 4384
rect 2005 4344 2007 4424
rect 2049 4344 2051 4424
rect 2055 4344 2061 4424
rect 2065 4344 2067 4424
rect 2089 4344 2091 4424
rect 2095 4344 2101 4424
rect 2105 4344 2107 4424
rect 2183 4344 2185 4384
rect 2189 4380 2205 4384
rect 2189 4344 2191 4380
rect 2203 4344 2205 4380
rect 2209 4344 2211 4384
rect 2223 4344 2225 4384
rect 2229 4344 2231 4384
rect 2288 4344 2290 4384
rect 2294 4344 2298 4384
rect 2310 4344 2312 4424
rect 2316 4344 2320 4424
rect 2324 4344 2326 4424
rect 2383 4344 2385 4384
rect 2389 4344 2391 4384
rect 2429 4344 2431 4424
rect 2435 4344 2439 4424
rect 2443 4344 2445 4424
rect 2523 4344 2525 4384
rect 2529 4344 2531 4384
rect 2574 4344 2576 4424
rect 2580 4344 2584 4424
rect 2588 4344 2590 4424
rect 2602 4344 2606 4384
rect 2610 4344 2612 4384
rect 2669 4344 2671 4384
rect 2675 4344 2679 4384
rect 2691 4344 2693 4424
rect 2697 4344 2699 4424
rect 2749 4344 2751 4384
rect 2755 4344 2759 4384
rect 2771 4344 2773 4424
rect 2777 4344 2779 4424
rect 2841 4344 2843 4424
rect 2847 4344 2849 4424
rect 2861 4344 2865 4384
rect 2869 4344 2871 4384
rect 2923 4344 2925 4384
rect 2929 4380 2945 4384
rect 2929 4344 2931 4380
rect 2943 4344 2945 4380
rect 2949 4344 2951 4384
rect 2963 4344 2965 4384
rect 2969 4344 2971 4384
rect 3019 4344 3021 4424
rect 3025 4344 3027 4424
rect 3039 4344 3043 4384
rect 3047 4344 3051 4384
rect 3063 4344 3065 4384
rect 3069 4344 3071 4384
rect 3121 4344 3123 4424
rect 3127 4344 3129 4424
rect 3357 4416 3371 4424
rect 3141 4344 3145 4384
rect 3149 4344 3151 4384
rect 3203 4344 3205 4384
rect 3209 4380 3225 4384
rect 3209 4344 3211 4380
rect 3223 4344 3225 4380
rect 3229 4344 3231 4384
rect 3243 4344 3245 4384
rect 3249 4344 3251 4384
rect 3289 4344 3291 4384
rect 3295 4344 3297 4384
rect 3309 4344 3311 4384
rect 3315 4344 3317 4384
rect 3369 4344 3371 4416
rect 3375 4412 3391 4424
rect 3375 4344 3377 4412
rect 3389 4344 3391 4412
rect 3395 4344 3397 4424
rect 3409 4344 3411 4424
rect 3415 4344 3417 4424
rect 3697 4416 3711 4424
rect 3469 4344 3471 4384
rect 3475 4344 3477 4384
rect 3529 4344 3531 4384
rect 3535 4344 3537 4384
rect 3549 4344 3551 4384
rect 3555 4344 3557 4384
rect 3609 4344 3611 4384
rect 3615 4344 3617 4384
rect 3629 4344 3631 4384
rect 3635 4380 3651 4384
rect 3635 4344 3637 4380
rect 3649 4344 3651 4380
rect 3655 4344 3657 4384
rect 3709 4344 3711 4416
rect 3715 4412 3731 4424
rect 3715 4344 3717 4412
rect 3729 4344 3731 4412
rect 3735 4344 3737 4424
rect 3749 4344 3751 4424
rect 3755 4344 3757 4424
rect 3814 4344 3816 4424
rect 3820 4344 3824 4424
rect 3828 4344 3830 4424
rect 3842 4344 3846 4384
rect 3850 4344 3852 4384
rect 3928 4344 3930 4384
rect 3934 4344 3938 4384
rect 3950 4344 3952 4424
rect 3956 4344 3960 4424
rect 3964 4344 3966 4424
rect 4197 4416 4211 4424
rect 4023 4344 4025 4384
rect 4029 4380 4045 4384
rect 4029 4344 4031 4380
rect 4043 4344 4045 4380
rect 4049 4344 4051 4384
rect 4063 4344 4065 4384
rect 4069 4344 4071 4384
rect 4123 4344 4125 4384
rect 4129 4380 4145 4384
rect 4129 4344 4131 4380
rect 4143 4344 4145 4380
rect 4149 4344 4151 4384
rect 4163 4344 4165 4384
rect 4169 4344 4171 4384
rect 4209 4344 4211 4416
rect 4215 4412 4231 4424
rect 4215 4344 4217 4412
rect 4229 4344 4231 4412
rect 4235 4344 4237 4424
rect 4249 4344 4251 4424
rect 4255 4344 4257 4424
rect 4309 4344 4311 4384
rect 4315 4344 4317 4384
rect 4329 4344 4331 4384
rect 4335 4344 4337 4384
rect 4403 4344 4405 4424
rect 4409 4344 4411 4424
rect 4423 4344 4425 4424
rect 4429 4412 4445 4424
rect 4429 4344 4431 4412
rect 4443 4344 4445 4412
rect 4449 4416 4463 4424
rect 4449 4344 4451 4416
rect 4503 4344 4505 4384
rect 4509 4344 4511 4384
rect 4549 4344 4551 4384
rect 4555 4344 4557 4384
rect 4569 4344 4571 4384
rect 4575 4380 4591 4384
rect 4575 4344 4577 4380
rect 4589 4344 4591 4380
rect 4595 4344 4597 4384
rect 4649 4344 4651 4384
rect 4655 4344 4657 4384
rect 4669 4344 4671 4384
rect 4675 4380 4691 4384
rect 4675 4344 4677 4380
rect 4689 4344 4691 4380
rect 4695 4344 4697 4384
rect 48 4276 50 4316
rect 54 4276 58 4316
rect 70 4236 72 4316
rect 76 4236 80 4316
rect 84 4236 86 4316
rect 139 4236 141 4316
rect 145 4236 147 4316
rect 159 4276 163 4316
rect 167 4276 171 4316
rect 183 4276 185 4316
rect 189 4276 191 4316
rect 229 4236 231 4316
rect 235 4236 239 4316
rect 243 4236 245 4316
rect 323 4236 325 4316
rect 329 4236 331 4316
rect 343 4236 345 4316
rect 349 4248 351 4316
rect 363 4248 365 4316
rect 349 4236 365 4248
rect 369 4244 371 4316
rect 409 4276 411 4316
rect 415 4276 417 4316
rect 429 4276 433 4316
rect 437 4276 441 4316
rect 369 4236 383 4244
rect 453 4236 455 4316
rect 459 4236 461 4316
rect 523 4236 525 4316
rect 529 4236 531 4316
rect 543 4236 545 4316
rect 549 4248 551 4316
rect 563 4248 565 4316
rect 549 4236 565 4248
rect 569 4244 571 4316
rect 609 4276 611 4316
rect 615 4276 617 4316
rect 629 4276 631 4316
rect 635 4280 637 4316
rect 649 4280 651 4316
rect 635 4276 651 4280
rect 655 4276 657 4316
rect 569 4236 583 4244
rect 709 4244 711 4316
rect 697 4236 711 4244
rect 715 4248 717 4316
rect 729 4248 731 4316
rect 715 4236 731 4248
rect 735 4236 737 4316
rect 749 4236 751 4316
rect 755 4236 757 4316
rect 809 4276 811 4316
rect 815 4276 817 4316
rect 829 4276 833 4316
rect 837 4276 841 4316
rect 853 4236 855 4316
rect 859 4236 861 4316
rect 928 4276 930 4316
rect 934 4276 938 4316
rect 950 4236 952 4316
rect 956 4236 960 4316
rect 964 4236 966 4316
rect 1023 4276 1025 4316
rect 1029 4276 1031 4316
rect 1069 4236 1071 4316
rect 1075 4236 1079 4316
rect 1083 4236 1085 4316
rect 1149 4236 1151 4316
rect 1155 4236 1159 4316
rect 1163 4236 1165 4316
rect 1229 4236 1231 4316
rect 1235 4236 1239 4316
rect 1243 4236 1245 4316
rect 1309 4276 1311 4316
rect 1315 4276 1317 4316
rect 1369 4236 1371 4316
rect 1375 4296 1377 4316
rect 1389 4296 1393 4316
rect 1397 4296 1401 4316
rect 1405 4296 1407 4316
rect 1419 4296 1421 4316
rect 1375 4236 1384 4296
rect 1410 4276 1421 4296
rect 1425 4276 1429 4316
rect 1433 4276 1435 4316
rect 1473 4276 1475 4316
rect 1479 4276 1481 4316
rect 1493 4276 1495 4316
rect 1499 4276 1507 4316
rect 1511 4276 1513 4316
rect 1525 4276 1527 4316
rect 1531 4276 1541 4316
rect 1545 4276 1547 4316
rect 1559 4276 1561 4316
rect 1552 4236 1561 4276
rect 1565 4236 1567 4316
rect 1614 4236 1616 4316
rect 1620 4236 1624 4316
rect 1628 4236 1630 4316
rect 1642 4276 1646 4316
rect 1650 4276 1652 4316
rect 1709 4236 1711 4316
rect 1715 4236 1719 4316
rect 1723 4236 1725 4316
rect 1803 4276 1805 4316
rect 1809 4276 1811 4316
rect 1849 4236 1851 4316
rect 1855 4296 1857 4316
rect 1869 4296 1873 4316
rect 1877 4296 1881 4316
rect 1885 4296 1887 4316
rect 1899 4296 1901 4316
rect 1855 4236 1864 4296
rect 1890 4276 1901 4296
rect 1905 4276 1909 4316
rect 1913 4276 1915 4316
rect 1953 4276 1955 4316
rect 1959 4276 1961 4316
rect 1973 4276 1975 4316
rect 1979 4276 1987 4316
rect 1991 4276 1993 4316
rect 2005 4276 2007 4316
rect 2011 4276 2021 4316
rect 2025 4276 2027 4316
rect 2039 4276 2041 4316
rect 2032 4236 2041 4276
rect 2045 4236 2047 4316
rect 2103 4276 2105 4316
rect 2109 4276 2111 4316
rect 2123 4276 2125 4316
rect 2129 4276 2131 4316
rect 2169 4236 2171 4316
rect 2175 4236 2181 4316
rect 2185 4237 2187 4316
rect 2199 4237 2201 4316
rect 2185 4236 2201 4237
rect 2205 4237 2207 4316
rect 2205 4236 2219 4237
rect 2283 4236 2285 4316
rect 2289 4304 2305 4316
rect 2289 4236 2291 4304
rect 2303 4236 2305 4304
rect 2309 4238 2311 4316
rect 2323 4238 2325 4316
rect 2309 4236 2325 4238
rect 2329 4250 2331 4316
rect 2343 4250 2345 4316
rect 2329 4236 2345 4250
rect 2349 4238 2351 4316
rect 2389 4276 2391 4316
rect 2395 4276 2397 4316
rect 2409 4276 2411 4316
rect 2415 4276 2417 4316
rect 2488 4276 2490 4316
rect 2494 4276 2498 4316
rect 2349 4236 2363 4238
rect 2510 4236 2512 4316
rect 2516 4236 2520 4316
rect 2524 4236 2526 4316
rect 2595 4236 2597 4316
rect 2601 4236 2605 4316
rect 2609 4236 2611 4316
rect 2649 4244 2651 4316
rect 2637 4236 2651 4244
rect 2655 4248 2657 4316
rect 2669 4248 2671 4316
rect 2655 4236 2671 4248
rect 2675 4236 2677 4316
rect 2689 4236 2691 4316
rect 2695 4236 2697 4316
rect 2763 4236 2765 4316
rect 2769 4236 2771 4316
rect 2783 4236 2785 4316
rect 2789 4248 2791 4316
rect 2803 4248 2805 4316
rect 2789 4236 2805 4248
rect 2809 4244 2811 4316
rect 2849 4276 2851 4316
rect 2855 4276 2859 4316
rect 2809 4236 2823 4244
rect 2871 4236 2873 4316
rect 2877 4236 2879 4316
rect 2943 4276 2945 4316
rect 2949 4280 2951 4316
rect 2963 4280 2965 4316
rect 2949 4276 2965 4280
rect 2969 4276 2971 4316
rect 2983 4276 2985 4316
rect 2989 4276 2991 4316
rect 3043 4276 3045 4316
rect 3049 4280 3051 4316
rect 3063 4280 3065 4316
rect 3049 4276 3065 4280
rect 3069 4276 3071 4316
rect 3083 4276 3085 4316
rect 3089 4276 3091 4316
rect 3129 4276 3131 4316
rect 3135 4276 3137 4316
rect 3149 4276 3151 4316
rect 3155 4276 3157 4316
rect 3223 4276 3225 4316
rect 3229 4276 3231 4316
rect 3283 4276 3285 4316
rect 3289 4280 3291 4316
rect 3303 4280 3305 4316
rect 3289 4276 3305 4280
rect 3309 4276 3311 4316
rect 3323 4276 3325 4316
rect 3329 4276 3331 4316
rect 3383 4276 3385 4316
rect 3389 4280 3391 4316
rect 3403 4280 3405 4316
rect 3389 4276 3405 4280
rect 3409 4276 3411 4316
rect 3423 4276 3425 4316
rect 3429 4276 3431 4316
rect 3483 4276 3485 4316
rect 3489 4280 3491 4316
rect 3503 4280 3505 4316
rect 3489 4276 3505 4280
rect 3509 4276 3511 4316
rect 3523 4276 3525 4316
rect 3529 4276 3531 4316
rect 3583 4276 3585 4316
rect 3589 4280 3591 4316
rect 3603 4280 3605 4316
rect 3589 4276 3605 4280
rect 3609 4276 3611 4316
rect 3623 4276 3625 4316
rect 3629 4276 3631 4316
rect 3669 4276 3671 4316
rect 3675 4276 3677 4316
rect 3689 4276 3691 4316
rect 3695 4280 3697 4316
rect 3709 4280 3711 4316
rect 3695 4276 3711 4280
rect 3715 4276 3717 4316
rect 3769 4244 3771 4316
rect 3757 4236 3771 4244
rect 3775 4248 3777 4316
rect 3789 4248 3791 4316
rect 3775 4236 3791 4248
rect 3795 4236 3797 4316
rect 3809 4236 3811 4316
rect 3815 4236 3817 4316
rect 3874 4236 3876 4316
rect 3880 4236 3884 4316
rect 3888 4236 3890 4316
rect 3902 4276 3906 4316
rect 3910 4276 3912 4316
rect 3969 4276 3971 4316
rect 3975 4276 3977 4316
rect 4029 4244 4031 4316
rect 4017 4236 4031 4244
rect 4035 4248 4037 4316
rect 4049 4248 4051 4316
rect 4035 4236 4051 4248
rect 4055 4236 4057 4316
rect 4069 4236 4071 4316
rect 4075 4236 4077 4316
rect 4143 4276 4145 4316
rect 4149 4280 4151 4316
rect 4163 4280 4165 4316
rect 4149 4276 4165 4280
rect 4169 4276 4171 4316
rect 4183 4276 4185 4316
rect 4189 4276 4191 4316
rect 4229 4276 4231 4316
rect 4235 4276 4237 4316
rect 4249 4276 4251 4316
rect 4255 4280 4257 4316
rect 4269 4280 4271 4316
rect 4255 4276 4271 4280
rect 4275 4276 4277 4316
rect 4329 4244 4331 4316
rect 4317 4236 4331 4244
rect 4335 4248 4337 4316
rect 4349 4248 4351 4316
rect 4335 4236 4351 4248
rect 4355 4236 4357 4316
rect 4369 4236 4371 4316
rect 4375 4236 4377 4316
rect 4434 4236 4436 4316
rect 4440 4236 4444 4316
rect 4448 4236 4450 4316
rect 4462 4276 4466 4316
rect 4470 4276 4472 4316
rect 4529 4238 4531 4316
rect 4517 4236 4531 4238
rect 4535 4250 4537 4316
rect 4549 4250 4551 4316
rect 4535 4236 4551 4250
rect 4555 4238 4557 4316
rect 4569 4238 4571 4316
rect 4555 4236 4571 4238
rect 4575 4304 4591 4316
rect 4575 4236 4577 4304
rect 4589 4236 4591 4304
rect 4595 4236 4597 4316
rect 4675 4236 4677 4316
rect 4681 4236 4685 4316
rect 4689 4236 4691 4316
rect 43 3864 45 3904
rect 49 3864 51 3904
rect 63 3864 65 3904
rect 69 3864 71 3904
rect 123 3864 125 3904
rect 129 3864 131 3904
rect 143 3864 145 3904
rect 149 3864 151 3904
rect 215 3864 217 3944
rect 221 3864 225 3944
rect 229 3864 231 3944
rect 274 3864 276 3944
rect 280 3864 284 3944
rect 288 3864 290 3944
rect 302 3864 306 3904
rect 310 3864 312 3904
rect 383 3864 385 3904
rect 389 3864 391 3904
rect 443 3864 445 3904
rect 449 3864 451 3904
rect 515 3864 517 3944
rect 521 3864 525 3944
rect 529 3864 531 3944
rect 569 3864 571 3904
rect 575 3864 577 3904
rect 589 3864 593 3904
rect 597 3864 601 3904
rect 613 3864 615 3944
rect 619 3864 621 3944
rect 674 3864 676 3944
rect 680 3864 684 3944
rect 688 3864 690 3944
rect 702 3864 706 3904
rect 710 3864 712 3904
rect 769 3864 771 3904
rect 775 3864 777 3904
rect 834 3864 836 3944
rect 840 3864 844 3944
rect 848 3864 850 3944
rect 862 3864 866 3904
rect 870 3864 872 3904
rect 929 3864 931 3904
rect 935 3864 937 3904
rect 949 3864 951 3904
rect 955 3864 957 3904
rect 1023 3864 1025 3904
rect 1029 3864 1031 3904
rect 1095 3864 1097 3944
rect 1101 3864 1105 3944
rect 1109 3864 1111 3944
rect 1149 3864 1151 3904
rect 1155 3864 1157 3904
rect 1209 3864 1211 3944
rect 1215 3864 1219 3944
rect 1223 3864 1225 3944
rect 1289 3864 1291 3904
rect 1295 3864 1297 3904
rect 1375 3864 1377 3944
rect 1381 3864 1385 3944
rect 1389 3864 1391 3944
rect 1443 3864 1445 3904
rect 1449 3864 1451 3904
rect 1494 3864 1496 3944
rect 1500 3864 1504 3944
rect 1508 3864 1510 3944
rect 1522 3864 1526 3904
rect 1530 3864 1532 3904
rect 1589 3864 1591 3944
rect 1595 3864 1601 3944
rect 1605 3864 1607 3944
rect 1629 3864 1631 3944
rect 1635 3864 1641 3944
rect 1645 3864 1647 3944
rect 1709 3864 1711 3904
rect 1715 3864 1717 3904
rect 1729 3864 1731 3904
rect 1735 3864 1737 3904
rect 1803 3864 1805 3944
rect 1809 3864 1811 3944
rect 1823 3864 1825 3944
rect 1829 3932 1845 3944
rect 1829 3864 1831 3932
rect 1843 3864 1845 3932
rect 1849 3936 1863 3944
rect 1849 3864 1851 3936
rect 1889 3864 1891 3904
rect 1895 3864 1897 3904
rect 1909 3864 1911 3904
rect 1915 3900 1931 3904
rect 1915 3864 1917 3900
rect 1929 3864 1931 3900
rect 1935 3864 1937 3904
rect 2008 3864 2010 3904
rect 2014 3864 2018 3904
rect 2030 3864 2032 3944
rect 2036 3864 2040 3944
rect 2044 3864 2046 3944
rect 2103 3864 2105 3904
rect 2109 3864 2111 3904
rect 2163 3864 2165 3904
rect 2169 3900 2185 3904
rect 2169 3864 2171 3900
rect 2183 3864 2185 3900
rect 2189 3864 2191 3904
rect 2203 3864 2205 3904
rect 2209 3864 2211 3904
rect 2263 3864 2265 3904
rect 2269 3900 2285 3904
rect 2269 3864 2271 3900
rect 2283 3864 2285 3900
rect 2289 3864 2291 3904
rect 2303 3864 2305 3904
rect 2309 3864 2311 3904
rect 2363 3864 2365 3944
rect 2369 3864 2371 3944
rect 2383 3864 2385 3944
rect 2389 3932 2405 3944
rect 2389 3864 2391 3932
rect 2403 3864 2405 3932
rect 2409 3936 2423 3944
rect 2409 3864 2411 3936
rect 2463 3864 2465 3904
rect 2469 3864 2471 3904
rect 2528 3864 2530 3904
rect 2534 3864 2538 3904
rect 2550 3864 2552 3944
rect 2556 3864 2560 3944
rect 2564 3864 2566 3944
rect 2623 3864 2625 3904
rect 2629 3900 2645 3904
rect 2629 3864 2631 3900
rect 2643 3864 2645 3900
rect 2649 3864 2651 3904
rect 2663 3864 2665 3904
rect 2669 3864 2671 3904
rect 2723 3864 2725 3944
rect 2729 3864 2731 3944
rect 2743 3864 2745 3944
rect 2749 3932 2765 3944
rect 2749 3864 2751 3932
rect 2763 3864 2765 3932
rect 2769 3936 2783 3944
rect 2769 3864 2771 3936
rect 2828 3864 2830 3904
rect 2834 3864 2838 3904
rect 2850 3864 2852 3944
rect 2856 3864 2860 3944
rect 2864 3864 2866 3944
rect 2914 3864 2916 3944
rect 2920 3864 2924 3944
rect 2928 3864 2930 3944
rect 2942 3864 2946 3904
rect 2950 3864 2952 3904
rect 3023 3864 3025 3904
rect 3029 3900 3045 3904
rect 3029 3864 3031 3900
rect 3043 3864 3045 3900
rect 3049 3864 3051 3904
rect 3063 3864 3065 3904
rect 3069 3864 3071 3904
rect 3123 3864 3125 3904
rect 3129 3864 3131 3904
rect 3174 3864 3176 3944
rect 3180 3864 3184 3944
rect 3188 3864 3190 3944
rect 3257 3936 3271 3944
rect 3202 3864 3206 3904
rect 3210 3864 3212 3904
rect 3269 3864 3271 3936
rect 3275 3932 3291 3944
rect 3275 3864 3277 3932
rect 3289 3864 3291 3932
rect 3295 3864 3297 3944
rect 3309 3864 3311 3944
rect 3315 3864 3317 3944
rect 3374 3864 3376 3944
rect 3380 3864 3384 3944
rect 3388 3864 3390 3944
rect 3402 3864 3406 3904
rect 3410 3864 3412 3904
rect 3488 3864 3490 3904
rect 3494 3864 3498 3904
rect 3510 3864 3512 3944
rect 3516 3864 3520 3944
rect 3524 3864 3526 3944
rect 3588 3864 3590 3904
rect 3594 3864 3598 3904
rect 3610 3864 3612 3944
rect 3616 3864 3620 3944
rect 3624 3864 3626 3944
rect 3683 3864 3685 3944
rect 3689 3864 3691 3944
rect 3703 3864 3705 3944
rect 3709 3932 3725 3944
rect 3709 3864 3711 3932
rect 3723 3864 3725 3932
rect 3729 3936 3743 3944
rect 3729 3864 3731 3936
rect 3783 3864 3785 3904
rect 3789 3900 3805 3904
rect 3789 3864 3791 3900
rect 3803 3864 3805 3900
rect 3809 3864 3811 3904
rect 3823 3864 3825 3904
rect 3829 3864 3831 3904
rect 3883 3864 3885 3904
rect 3889 3864 3891 3904
rect 3903 3864 3905 3904
rect 3909 3864 3911 3904
rect 3963 3864 3965 3904
rect 3969 3864 3971 3904
rect 3983 3864 3985 3904
rect 3989 3864 3991 3904
rect 4029 3864 4031 3904
rect 4035 3864 4037 3904
rect 4049 3864 4051 3904
rect 4055 3864 4057 3904
rect 4123 3864 4125 3904
rect 4129 3900 4145 3904
rect 4129 3864 4131 3900
rect 4143 3864 4145 3900
rect 4149 3864 4151 3904
rect 4163 3864 4165 3904
rect 4169 3864 4171 3904
rect 4228 3864 4230 3904
rect 4234 3864 4238 3904
rect 4250 3864 4252 3944
rect 4256 3864 4260 3944
rect 4264 3864 4266 3944
rect 4314 3864 4316 3944
rect 4320 3864 4324 3944
rect 4328 3864 4330 3944
rect 4657 3936 4671 3944
rect 4342 3864 4346 3904
rect 4350 3864 4352 3904
rect 4423 3864 4425 3904
rect 4429 3864 4431 3904
rect 4483 3864 4485 3904
rect 4489 3900 4505 3904
rect 4489 3864 4491 3900
rect 4503 3864 4505 3900
rect 4509 3864 4511 3904
rect 4523 3864 4525 3904
rect 4529 3864 4531 3904
rect 4583 3864 4585 3904
rect 4589 3900 4605 3904
rect 4589 3864 4591 3900
rect 4603 3864 4605 3900
rect 4609 3864 4611 3904
rect 4623 3864 4625 3904
rect 4629 3864 4631 3904
rect 4669 3864 4671 3936
rect 4675 3932 4691 3944
rect 4675 3864 4677 3932
rect 4689 3864 4691 3932
rect 4695 3864 4697 3944
rect 4709 3864 4711 3944
rect 4715 3864 4717 3944
rect 48 3796 50 3836
rect 54 3796 58 3836
rect 70 3756 72 3836
rect 76 3756 80 3836
rect 84 3756 86 3836
rect 143 3796 145 3836
rect 149 3796 151 3836
rect 189 3756 191 3836
rect 195 3816 197 3836
rect 209 3816 213 3836
rect 217 3816 221 3836
rect 225 3816 227 3836
rect 239 3816 241 3836
rect 195 3756 204 3816
rect 230 3796 241 3816
rect 245 3796 249 3836
rect 253 3796 255 3836
rect 293 3796 295 3836
rect 299 3796 301 3836
rect 313 3796 315 3836
rect 319 3796 327 3836
rect 331 3796 333 3836
rect 345 3796 347 3836
rect 351 3796 361 3836
rect 365 3796 367 3836
rect 379 3796 381 3836
rect 372 3756 381 3796
rect 385 3756 387 3836
rect 448 3796 450 3836
rect 454 3796 458 3836
rect 470 3756 472 3836
rect 476 3756 480 3836
rect 484 3756 486 3836
rect 529 3796 531 3836
rect 535 3796 537 3836
rect 549 3796 553 3836
rect 557 3796 561 3836
rect 573 3756 575 3836
rect 579 3756 581 3836
rect 653 3757 655 3836
rect 641 3756 655 3757
rect 659 3757 661 3836
rect 673 3757 675 3836
rect 659 3756 675 3757
rect 679 3756 685 3836
rect 689 3756 691 3836
rect 743 3796 745 3836
rect 749 3796 751 3836
rect 763 3796 765 3836
rect 769 3796 771 3836
rect 813 3756 815 3836
rect 819 3796 821 3836
rect 833 3796 835 3836
rect 839 3796 849 3836
rect 853 3796 855 3836
rect 867 3796 869 3836
rect 873 3796 881 3836
rect 885 3796 887 3836
rect 899 3796 901 3836
rect 905 3796 907 3836
rect 945 3796 947 3836
rect 951 3796 955 3836
rect 959 3816 961 3836
rect 973 3816 975 3836
rect 979 3816 983 3836
rect 987 3816 991 3836
rect 1003 3816 1005 3836
rect 959 3796 970 3816
rect 819 3756 828 3796
rect 996 3756 1005 3816
rect 1009 3756 1011 3836
rect 1061 3756 1063 3836
rect 1067 3756 1069 3836
rect 1081 3796 1085 3836
rect 1089 3796 1091 3836
rect 1129 3756 1131 3836
rect 1135 3816 1137 3836
rect 1149 3816 1153 3836
rect 1157 3816 1161 3836
rect 1165 3816 1167 3836
rect 1179 3816 1181 3836
rect 1135 3756 1144 3816
rect 1170 3796 1181 3816
rect 1185 3796 1189 3836
rect 1193 3796 1195 3836
rect 1233 3796 1235 3836
rect 1239 3796 1241 3836
rect 1253 3796 1255 3836
rect 1259 3796 1267 3836
rect 1271 3796 1273 3836
rect 1285 3796 1287 3836
rect 1291 3796 1301 3836
rect 1305 3796 1307 3836
rect 1319 3796 1321 3836
rect 1312 3756 1321 3796
rect 1325 3756 1327 3836
rect 1374 3756 1376 3836
rect 1380 3756 1384 3836
rect 1388 3756 1390 3836
rect 1402 3796 1406 3836
rect 1410 3796 1412 3836
rect 1469 3796 1471 3836
rect 1475 3796 1477 3836
rect 1489 3796 1491 3836
rect 1495 3796 1497 3836
rect 1549 3796 1551 3836
rect 1555 3796 1557 3836
rect 1569 3796 1571 3836
rect 1575 3796 1577 3836
rect 1629 3796 1631 3836
rect 1635 3796 1639 3836
rect 1651 3756 1653 3836
rect 1657 3756 1659 3836
rect 1709 3756 1711 3836
rect 1715 3816 1717 3836
rect 1729 3816 1733 3836
rect 1737 3816 1741 3836
rect 1745 3816 1747 3836
rect 1759 3816 1761 3836
rect 1715 3756 1724 3816
rect 1750 3796 1761 3816
rect 1765 3796 1769 3836
rect 1773 3796 1775 3836
rect 1813 3796 1815 3836
rect 1819 3796 1821 3836
rect 1833 3796 1835 3836
rect 1839 3796 1847 3836
rect 1851 3796 1853 3836
rect 1865 3796 1867 3836
rect 1871 3796 1881 3836
rect 1885 3796 1887 3836
rect 1899 3796 1901 3836
rect 1892 3756 1901 3796
rect 1905 3756 1907 3836
rect 1963 3796 1965 3836
rect 1969 3796 1971 3836
rect 2023 3756 2025 3836
rect 2029 3756 2031 3836
rect 2043 3756 2045 3836
rect 2049 3768 2051 3836
rect 2063 3768 2065 3836
rect 2049 3756 2065 3768
rect 2069 3764 2071 3836
rect 2123 3796 2125 3836
rect 2129 3796 2131 3836
rect 2169 3796 2171 3836
rect 2175 3796 2177 3836
rect 2189 3796 2191 3836
rect 2195 3800 2197 3836
rect 2209 3800 2211 3836
rect 2195 3796 2211 3800
rect 2215 3796 2217 3836
rect 2288 3796 2290 3836
rect 2294 3796 2298 3836
rect 2069 3756 2083 3764
rect 2310 3756 2312 3836
rect 2316 3756 2320 3836
rect 2324 3756 2326 3836
rect 2383 3796 2385 3836
rect 2389 3800 2391 3836
rect 2403 3800 2405 3836
rect 2389 3796 2405 3800
rect 2409 3796 2411 3836
rect 2423 3796 2425 3836
rect 2429 3796 2431 3836
rect 2483 3756 2485 3836
rect 2489 3756 2491 3836
rect 2503 3756 2505 3836
rect 2509 3768 2511 3836
rect 2523 3768 2525 3836
rect 2509 3756 2525 3768
rect 2529 3764 2531 3836
rect 2583 3796 2585 3836
rect 2589 3800 2591 3836
rect 2603 3800 2605 3836
rect 2589 3796 2605 3800
rect 2609 3796 2611 3836
rect 2623 3796 2625 3836
rect 2629 3796 2631 3836
rect 2529 3756 2543 3764
rect 2669 3764 2671 3836
rect 2657 3756 2671 3764
rect 2675 3768 2677 3836
rect 2689 3768 2691 3836
rect 2675 3756 2691 3768
rect 2695 3756 2697 3836
rect 2709 3756 2711 3836
rect 2715 3756 2717 3836
rect 2783 3756 2785 3836
rect 2789 3756 2791 3836
rect 2803 3756 2805 3836
rect 2809 3768 2811 3836
rect 2823 3768 2825 3836
rect 2809 3756 2825 3768
rect 2829 3764 2831 3836
rect 2883 3796 2885 3836
rect 2889 3796 2891 3836
rect 2943 3796 2945 3836
rect 2949 3796 2951 3836
rect 3003 3796 3005 3836
rect 3009 3800 3011 3836
rect 3023 3800 3025 3836
rect 3009 3796 3025 3800
rect 3029 3796 3031 3836
rect 3043 3796 3045 3836
rect 3049 3796 3051 3836
rect 2829 3756 2843 3764
rect 3103 3756 3105 3836
rect 3109 3756 3111 3836
rect 3123 3756 3125 3836
rect 3129 3768 3131 3836
rect 3143 3768 3145 3836
rect 3129 3756 3145 3768
rect 3149 3764 3151 3836
rect 3203 3796 3205 3836
rect 3209 3800 3211 3836
rect 3223 3800 3225 3836
rect 3209 3796 3225 3800
rect 3229 3796 3231 3836
rect 3243 3796 3245 3836
rect 3249 3796 3251 3836
rect 3303 3796 3305 3836
rect 3309 3796 3311 3836
rect 3368 3796 3370 3836
rect 3374 3796 3378 3836
rect 3149 3756 3163 3764
rect 3390 3756 3392 3836
rect 3396 3756 3400 3836
rect 3404 3756 3406 3836
rect 3463 3796 3465 3836
rect 3469 3796 3471 3836
rect 3483 3796 3485 3836
rect 3489 3796 3491 3836
rect 3529 3796 3531 3836
rect 3535 3796 3537 3836
rect 3549 3796 3553 3836
rect 3557 3796 3561 3836
rect 3573 3756 3575 3836
rect 3579 3756 3581 3836
rect 3643 3756 3645 3836
rect 3649 3756 3651 3836
rect 3663 3756 3665 3836
rect 3669 3768 3671 3836
rect 3683 3768 3685 3836
rect 3669 3756 3685 3768
rect 3689 3764 3691 3836
rect 3743 3796 3745 3836
rect 3749 3800 3751 3836
rect 3763 3800 3765 3836
rect 3749 3796 3765 3800
rect 3769 3796 3771 3836
rect 3783 3796 3785 3836
rect 3789 3796 3791 3836
rect 3843 3796 3845 3836
rect 3849 3796 3851 3836
rect 3689 3756 3703 3764
rect 3889 3764 3891 3836
rect 3877 3756 3891 3764
rect 3895 3768 3897 3836
rect 3909 3768 3911 3836
rect 3895 3756 3911 3768
rect 3915 3756 3917 3836
rect 3929 3756 3931 3836
rect 3935 3756 3937 3836
rect 4008 3796 4010 3836
rect 4014 3796 4018 3836
rect 4030 3756 4032 3836
rect 4036 3756 4040 3836
rect 4044 3756 4046 3836
rect 4094 3756 4096 3836
rect 4100 3756 4104 3836
rect 4108 3756 4110 3836
rect 4122 3796 4126 3836
rect 4130 3796 4132 3836
rect 4189 3764 4191 3836
rect 4177 3756 4191 3764
rect 4195 3768 4197 3836
rect 4209 3768 4211 3836
rect 4195 3756 4211 3768
rect 4215 3756 4217 3836
rect 4229 3756 4231 3836
rect 4235 3756 4237 3836
rect 4303 3756 4305 3836
rect 4309 3756 4311 3836
rect 4323 3756 4325 3836
rect 4329 3768 4331 3836
rect 4343 3768 4345 3836
rect 4329 3756 4345 3768
rect 4349 3764 4351 3836
rect 4389 3796 4391 3836
rect 4395 3796 4397 3836
rect 4409 3796 4411 3836
rect 4415 3800 4417 3836
rect 4429 3800 4431 3836
rect 4415 3796 4431 3800
rect 4435 3796 4437 3836
rect 4503 3796 4505 3836
rect 4509 3796 4511 3836
rect 4563 3796 4565 3836
rect 4569 3800 4571 3836
rect 4583 3800 4585 3836
rect 4569 3796 4585 3800
rect 4589 3796 4591 3836
rect 4603 3796 4605 3836
rect 4609 3796 4611 3836
rect 4649 3796 4651 3836
rect 4655 3796 4657 3836
rect 4669 3796 4671 3836
rect 4675 3800 4677 3836
rect 4689 3800 4691 3836
rect 4675 3796 4691 3800
rect 4695 3796 4697 3836
rect 4349 3756 4363 3764
rect 33 3384 35 3464
rect 39 3424 48 3464
rect 39 3384 41 3424
rect 53 3384 55 3424
rect 59 3384 69 3424
rect 73 3384 75 3424
rect 87 3384 89 3424
rect 93 3384 101 3424
rect 105 3384 107 3424
rect 119 3384 121 3424
rect 125 3384 127 3424
rect 165 3384 167 3424
rect 171 3384 175 3424
rect 179 3404 190 3424
rect 216 3404 225 3464
rect 179 3384 181 3404
rect 193 3384 195 3404
rect 199 3384 203 3404
rect 207 3384 211 3404
rect 223 3384 225 3404
rect 229 3384 231 3464
rect 283 3384 285 3424
rect 289 3384 291 3424
rect 303 3384 305 3424
rect 309 3384 311 3424
rect 368 3384 370 3424
rect 374 3384 378 3424
rect 390 3384 392 3464
rect 396 3384 400 3464
rect 404 3384 406 3464
rect 463 3384 465 3424
rect 469 3384 471 3424
rect 483 3384 485 3424
rect 489 3384 491 3424
rect 543 3384 545 3424
rect 549 3420 565 3424
rect 549 3384 551 3420
rect 563 3384 565 3420
rect 569 3384 571 3424
rect 583 3384 585 3424
rect 589 3384 591 3424
rect 643 3384 645 3424
rect 649 3384 651 3424
rect 708 3384 710 3424
rect 714 3384 718 3424
rect 730 3384 732 3464
rect 736 3384 740 3464
rect 744 3384 746 3464
rect 808 3384 810 3424
rect 814 3384 818 3424
rect 830 3384 832 3464
rect 836 3384 840 3464
rect 844 3384 846 3464
rect 889 3384 891 3424
rect 895 3384 897 3424
rect 975 3384 977 3464
rect 981 3384 985 3464
rect 989 3384 991 3464
rect 1029 3384 1031 3464
rect 1035 3404 1044 3464
rect 1212 3424 1221 3464
rect 1070 3404 1081 3424
rect 1035 3384 1037 3404
rect 1049 3384 1053 3404
rect 1057 3384 1061 3404
rect 1065 3384 1067 3404
rect 1079 3384 1081 3404
rect 1085 3384 1089 3424
rect 1093 3384 1095 3424
rect 1133 3384 1135 3424
rect 1139 3384 1141 3424
rect 1153 3384 1155 3424
rect 1159 3384 1167 3424
rect 1171 3384 1173 3424
rect 1185 3384 1187 3424
rect 1191 3384 1201 3424
rect 1205 3384 1207 3424
rect 1219 3384 1221 3424
rect 1225 3384 1227 3464
rect 1269 3384 1271 3424
rect 1275 3384 1277 3424
rect 1329 3384 1331 3464
rect 1335 3384 1339 3464
rect 1343 3384 1345 3464
rect 1414 3384 1416 3464
rect 1420 3384 1424 3464
rect 1428 3384 1430 3464
rect 1442 3384 1446 3424
rect 1450 3384 1452 3424
rect 1509 3384 1511 3424
rect 1515 3384 1517 3424
rect 1529 3384 1531 3424
rect 1535 3384 1537 3424
rect 1601 3384 1603 3464
rect 1607 3384 1609 3464
rect 1621 3384 1625 3424
rect 1629 3384 1631 3424
rect 1683 3384 1685 3424
rect 1689 3384 1691 3424
rect 1729 3384 1731 3464
rect 1735 3404 1744 3464
rect 1912 3424 1921 3464
rect 1770 3404 1781 3424
rect 1735 3384 1737 3404
rect 1749 3384 1753 3404
rect 1757 3384 1761 3404
rect 1765 3384 1767 3404
rect 1779 3384 1781 3404
rect 1785 3384 1789 3424
rect 1793 3384 1795 3424
rect 1833 3384 1835 3424
rect 1839 3384 1841 3424
rect 1853 3384 1855 3424
rect 1859 3384 1867 3424
rect 1871 3384 1873 3424
rect 1885 3384 1887 3424
rect 1891 3384 1901 3424
rect 1905 3384 1907 3424
rect 1919 3384 1921 3424
rect 1925 3384 1927 3464
rect 1969 3384 1971 3464
rect 1975 3384 1981 3464
rect 1985 3384 1987 3464
rect 2009 3384 2011 3464
rect 2015 3384 2021 3464
rect 2025 3384 2027 3464
rect 2089 3384 2091 3424
rect 2095 3384 2097 3424
rect 2109 3384 2111 3424
rect 2115 3384 2117 3424
rect 2183 3384 2185 3464
rect 2189 3384 2191 3464
rect 2203 3384 2205 3464
rect 2209 3452 2225 3464
rect 2209 3384 2211 3452
rect 2223 3384 2225 3452
rect 2229 3456 2243 3464
rect 2229 3384 2231 3456
rect 2283 3384 2285 3424
rect 2289 3420 2305 3424
rect 2289 3384 2291 3420
rect 2303 3384 2305 3420
rect 2309 3384 2311 3424
rect 2323 3384 2325 3424
rect 2329 3384 2331 3424
rect 2383 3384 2385 3424
rect 2389 3384 2391 3424
rect 2443 3384 2445 3424
rect 2449 3420 2465 3424
rect 2449 3384 2451 3420
rect 2463 3384 2465 3420
rect 2469 3384 2471 3424
rect 2483 3384 2485 3424
rect 2489 3384 2491 3424
rect 2543 3384 2545 3424
rect 2549 3420 2565 3424
rect 2549 3384 2551 3420
rect 2563 3384 2565 3420
rect 2569 3384 2571 3424
rect 2583 3384 2585 3424
rect 2589 3384 2591 3424
rect 2648 3384 2650 3424
rect 2654 3384 2658 3424
rect 2670 3384 2672 3464
rect 2676 3384 2680 3464
rect 2684 3384 2686 3464
rect 2734 3384 2736 3464
rect 2740 3384 2744 3464
rect 2748 3384 2750 3464
rect 2762 3384 2766 3424
rect 2770 3384 2772 3424
rect 2829 3384 2831 3424
rect 2835 3384 2837 3424
rect 2849 3384 2851 3424
rect 2855 3384 2857 3424
rect 2914 3384 2916 3464
rect 2920 3384 2924 3464
rect 2928 3384 2930 3464
rect 2942 3384 2946 3424
rect 2950 3384 2952 3424
rect 3009 3384 3011 3464
rect 3015 3384 3019 3464
rect 3023 3384 3025 3464
rect 3108 3384 3110 3424
rect 3114 3384 3118 3424
rect 3130 3384 3132 3464
rect 3136 3384 3140 3464
rect 3144 3384 3146 3464
rect 3177 3462 3191 3464
rect 3189 3384 3191 3462
rect 3195 3450 3211 3464
rect 3195 3384 3197 3450
rect 3209 3384 3211 3450
rect 3215 3462 3231 3464
rect 3215 3384 3217 3462
rect 3229 3384 3231 3462
rect 3235 3396 3237 3464
rect 3249 3396 3251 3464
rect 3235 3384 3251 3396
rect 3255 3384 3257 3464
rect 3309 3384 3311 3424
rect 3315 3384 3317 3424
rect 3329 3384 3331 3424
rect 3335 3384 3337 3424
rect 3389 3384 3391 3424
rect 3395 3384 3397 3424
rect 3409 3384 3411 3424
rect 3415 3384 3417 3424
rect 3469 3384 3471 3424
rect 3475 3384 3477 3424
rect 3489 3384 3491 3424
rect 3495 3384 3497 3424
rect 3549 3384 3551 3464
rect 3555 3384 3559 3464
rect 3563 3384 3565 3464
rect 3629 3384 3631 3424
rect 3635 3384 3637 3424
rect 3649 3384 3651 3424
rect 3655 3384 3657 3424
rect 3709 3384 3711 3424
rect 3715 3384 3717 3424
rect 3729 3384 3731 3424
rect 3735 3384 3737 3424
rect 3803 3384 3805 3424
rect 3809 3384 3811 3424
rect 3823 3384 3825 3424
rect 3829 3384 3831 3424
rect 3895 3384 3897 3464
rect 3901 3384 3905 3464
rect 3909 3384 3911 3464
rect 3949 3384 3951 3424
rect 3955 3384 3957 3424
rect 3969 3384 3971 3424
rect 3975 3384 3977 3424
rect 4029 3384 4031 3424
rect 4035 3384 4037 3424
rect 4049 3384 4051 3424
rect 4055 3384 4057 3424
rect 4114 3384 4116 3464
rect 4120 3384 4124 3464
rect 4128 3384 4130 3464
rect 4397 3456 4411 3464
rect 4142 3384 4146 3424
rect 4150 3384 4152 3424
rect 4223 3384 4225 3424
rect 4229 3420 4245 3424
rect 4229 3384 4231 3420
rect 4243 3384 4245 3420
rect 4249 3384 4251 3424
rect 4263 3384 4265 3424
rect 4269 3384 4271 3424
rect 4309 3384 4311 3424
rect 4315 3384 4317 3424
rect 4329 3384 4331 3424
rect 4335 3420 4351 3424
rect 4335 3384 4337 3420
rect 4349 3384 4351 3420
rect 4355 3384 4357 3424
rect 4409 3384 4411 3456
rect 4415 3452 4431 3464
rect 4415 3384 4417 3452
rect 4429 3384 4431 3452
rect 4435 3384 4437 3464
rect 4449 3384 4451 3464
rect 4455 3384 4457 3464
rect 4509 3384 4511 3424
rect 4515 3384 4517 3424
rect 4583 3384 4585 3424
rect 4589 3420 4605 3424
rect 4589 3384 4591 3420
rect 4603 3384 4605 3420
rect 4609 3384 4611 3424
rect 4623 3384 4625 3424
rect 4629 3384 4631 3424
rect 4669 3384 4671 3424
rect 4675 3384 4677 3424
rect 4689 3384 4691 3424
rect 4695 3420 4711 3424
rect 4695 3384 4697 3420
rect 4709 3384 4711 3420
rect 4715 3384 4717 3424
rect 33 3276 35 3356
rect 39 3316 41 3356
rect 53 3316 55 3356
rect 59 3316 69 3356
rect 73 3316 75 3356
rect 87 3316 89 3356
rect 93 3316 101 3356
rect 105 3316 107 3356
rect 119 3316 121 3356
rect 125 3316 127 3356
rect 165 3316 167 3356
rect 171 3316 175 3356
rect 179 3336 181 3356
rect 193 3336 195 3356
rect 199 3336 203 3356
rect 207 3336 211 3356
rect 223 3336 225 3356
rect 179 3316 190 3336
rect 39 3276 48 3316
rect 216 3276 225 3336
rect 229 3276 231 3356
rect 283 3276 285 3356
rect 289 3344 305 3356
rect 289 3276 291 3344
rect 303 3276 305 3344
rect 309 3278 311 3356
rect 323 3278 325 3356
rect 309 3276 325 3278
rect 329 3290 331 3356
rect 343 3290 345 3356
rect 329 3276 345 3290
rect 349 3278 351 3356
rect 389 3316 391 3356
rect 395 3316 397 3356
rect 409 3316 411 3356
rect 415 3316 417 3356
rect 349 3276 363 3278
rect 474 3276 476 3356
rect 480 3276 484 3356
rect 488 3276 490 3356
rect 502 3316 506 3356
rect 510 3316 512 3356
rect 574 3276 576 3356
rect 580 3276 584 3356
rect 588 3276 590 3356
rect 602 3316 606 3356
rect 610 3316 612 3356
rect 683 3316 685 3356
rect 689 3316 691 3356
rect 703 3316 705 3356
rect 709 3316 711 3356
rect 749 3316 751 3356
rect 755 3316 757 3356
rect 823 3276 825 3356
rect 829 3276 831 3356
rect 843 3276 845 3356
rect 849 3276 851 3356
rect 863 3276 865 3356
rect 869 3276 871 3356
rect 883 3276 885 3356
rect 889 3276 891 3356
rect 903 3276 905 3356
rect 909 3276 911 3356
rect 923 3276 925 3356
rect 929 3276 931 3356
rect 943 3276 945 3356
rect 949 3276 951 3356
rect 963 3276 965 3356
rect 969 3276 971 3356
rect 1009 3276 1011 3356
rect 1015 3276 1017 3356
rect 1029 3276 1031 3356
rect 1035 3276 1037 3356
rect 1049 3276 1051 3356
rect 1055 3276 1057 3356
rect 1069 3276 1071 3356
rect 1075 3276 1077 3356
rect 1089 3276 1091 3356
rect 1095 3276 1097 3356
rect 1109 3276 1111 3356
rect 1115 3276 1117 3356
rect 1129 3276 1131 3356
rect 1135 3276 1137 3356
rect 1149 3276 1151 3356
rect 1155 3276 1157 3356
rect 1223 3316 1225 3356
rect 1229 3316 1231 3356
rect 1269 3276 1271 3356
rect 1275 3336 1277 3356
rect 1289 3336 1293 3356
rect 1297 3336 1301 3356
rect 1305 3336 1307 3356
rect 1319 3336 1321 3356
rect 1275 3276 1284 3336
rect 1310 3316 1321 3336
rect 1325 3316 1329 3356
rect 1333 3316 1335 3356
rect 1373 3316 1375 3356
rect 1379 3316 1381 3356
rect 1393 3316 1395 3356
rect 1399 3316 1407 3356
rect 1411 3316 1413 3356
rect 1425 3316 1427 3356
rect 1431 3316 1441 3356
rect 1445 3316 1447 3356
rect 1459 3316 1461 3356
rect 1452 3276 1461 3316
rect 1465 3276 1467 3356
rect 1514 3276 1516 3356
rect 1520 3276 1524 3356
rect 1528 3276 1530 3356
rect 1542 3316 1546 3356
rect 1550 3316 1552 3356
rect 1628 3316 1630 3356
rect 1634 3316 1638 3356
rect 1650 3276 1652 3356
rect 1656 3276 1660 3356
rect 1664 3276 1666 3356
rect 1728 3316 1730 3356
rect 1734 3316 1738 3356
rect 1750 3276 1752 3356
rect 1756 3276 1760 3356
rect 1764 3276 1766 3356
rect 1823 3316 1825 3356
rect 1829 3316 1831 3356
rect 1888 3316 1890 3356
rect 1894 3316 1898 3356
rect 1910 3276 1912 3356
rect 1916 3276 1920 3356
rect 1924 3276 1926 3356
rect 1988 3316 1990 3356
rect 1994 3316 1998 3356
rect 2010 3276 2012 3356
rect 2016 3276 2020 3356
rect 2024 3276 2026 3356
rect 2069 3276 2071 3356
rect 2075 3336 2077 3356
rect 2089 3336 2093 3356
rect 2097 3336 2101 3356
rect 2105 3336 2107 3356
rect 2119 3336 2121 3356
rect 2075 3276 2084 3336
rect 2110 3316 2121 3336
rect 2125 3316 2129 3356
rect 2133 3316 2135 3356
rect 2173 3316 2175 3356
rect 2179 3316 2181 3356
rect 2193 3316 2195 3356
rect 2199 3316 2207 3356
rect 2211 3316 2213 3356
rect 2225 3316 2227 3356
rect 2231 3316 2241 3356
rect 2245 3316 2247 3356
rect 2259 3316 2261 3356
rect 2252 3276 2261 3316
rect 2265 3276 2267 3356
rect 2323 3316 2325 3356
rect 2329 3316 2331 3356
rect 2383 3316 2385 3356
rect 2389 3316 2391 3356
rect 2443 3316 2445 3356
rect 2449 3320 2451 3356
rect 2463 3320 2465 3356
rect 2449 3316 2465 3320
rect 2469 3316 2471 3356
rect 2483 3316 2485 3356
rect 2489 3316 2491 3356
rect 2529 3284 2531 3356
rect 2517 3276 2531 3284
rect 2535 3288 2537 3356
rect 2549 3288 2551 3356
rect 2535 3276 2551 3288
rect 2555 3276 2557 3356
rect 2569 3276 2571 3356
rect 2575 3276 2577 3356
rect 2643 3316 2645 3356
rect 2649 3316 2651 3356
rect 2708 3316 2710 3356
rect 2714 3316 2718 3356
rect 2730 3276 2732 3356
rect 2736 3276 2740 3356
rect 2744 3276 2746 3356
rect 2789 3276 2791 3356
rect 2795 3276 2799 3356
rect 2803 3276 2805 3356
rect 2874 3276 2876 3356
rect 2880 3276 2884 3356
rect 2888 3276 2890 3356
rect 2902 3316 2906 3356
rect 2910 3316 2912 3356
rect 2969 3316 2971 3356
rect 2975 3316 2977 3356
rect 2989 3316 2991 3356
rect 2995 3316 2997 3356
rect 3049 3316 3051 3356
rect 3055 3316 3057 3356
rect 3069 3316 3071 3356
rect 3075 3316 3077 3356
rect 3143 3276 3145 3356
rect 3149 3276 3151 3356
rect 3163 3276 3165 3356
rect 3169 3288 3171 3356
rect 3183 3288 3185 3356
rect 3169 3276 3185 3288
rect 3189 3284 3191 3356
rect 3243 3316 3245 3356
rect 3249 3320 3251 3356
rect 3263 3320 3265 3356
rect 3249 3316 3265 3320
rect 3269 3316 3271 3356
rect 3283 3316 3285 3356
rect 3289 3316 3291 3356
rect 3348 3316 3350 3356
rect 3354 3316 3358 3356
rect 3189 3276 3203 3284
rect 3370 3276 3372 3356
rect 3376 3276 3380 3356
rect 3384 3276 3386 3356
rect 3439 3276 3441 3356
rect 3445 3276 3447 3356
rect 3459 3316 3463 3356
rect 3467 3316 3471 3356
rect 3483 3316 3485 3356
rect 3489 3316 3491 3356
rect 3529 3316 3531 3356
rect 3535 3316 3537 3356
rect 3549 3316 3551 3356
rect 3555 3316 3557 3356
rect 3619 3276 3621 3356
rect 3625 3276 3627 3356
rect 3639 3316 3643 3356
rect 3647 3316 3651 3356
rect 3663 3316 3665 3356
rect 3669 3316 3671 3356
rect 3723 3276 3725 3356
rect 3729 3344 3745 3356
rect 3729 3276 3731 3344
rect 3743 3276 3745 3344
rect 3749 3278 3751 3356
rect 3763 3278 3765 3356
rect 3749 3276 3765 3278
rect 3769 3290 3771 3356
rect 3783 3290 3785 3356
rect 3769 3276 3785 3290
rect 3789 3278 3791 3356
rect 3843 3316 3845 3356
rect 3849 3316 3851 3356
rect 3863 3316 3865 3356
rect 3869 3316 3871 3356
rect 3789 3276 3803 3278
rect 3914 3276 3916 3356
rect 3920 3276 3924 3356
rect 3928 3276 3930 3356
rect 3942 3316 3946 3356
rect 3950 3316 3952 3356
rect 4009 3316 4011 3356
rect 4015 3316 4017 3356
rect 4029 3316 4031 3356
rect 4035 3316 4037 3356
rect 4099 3276 4101 3356
rect 4105 3276 4107 3356
rect 4119 3316 4123 3356
rect 4127 3316 4131 3356
rect 4143 3316 4145 3356
rect 4149 3316 4151 3356
rect 4189 3316 4191 3356
rect 4195 3316 4197 3356
rect 4209 3316 4211 3356
rect 4215 3316 4217 3356
rect 4269 3316 4271 3356
rect 4275 3316 4277 3356
rect 4289 3316 4293 3356
rect 4297 3316 4301 3356
rect 4313 3276 4315 3356
rect 4319 3276 4321 3356
rect 4369 3284 4371 3356
rect 4357 3276 4371 3284
rect 4375 3288 4377 3356
rect 4389 3288 4391 3356
rect 4375 3276 4391 3288
rect 4395 3276 4397 3356
rect 4409 3276 4411 3356
rect 4415 3276 4417 3356
rect 4474 3276 4476 3356
rect 4480 3276 4484 3356
rect 4488 3276 4490 3356
rect 4502 3316 4506 3356
rect 4510 3316 4512 3356
rect 4574 3276 4576 3356
rect 4580 3276 4584 3356
rect 4588 3276 4590 3356
rect 4602 3316 4606 3356
rect 4610 3316 4612 3356
rect 4683 3316 4685 3356
rect 4689 3320 4691 3356
rect 4703 3320 4705 3356
rect 4689 3316 4705 3320
rect 4709 3316 4711 3356
rect 4723 3316 4725 3356
rect 4729 3316 4731 3356
rect 33 2904 35 2984
rect 39 2944 48 2984
rect 39 2904 41 2944
rect 53 2904 55 2944
rect 59 2904 69 2944
rect 73 2904 75 2944
rect 87 2904 89 2944
rect 93 2904 101 2944
rect 105 2904 107 2944
rect 119 2904 121 2944
rect 125 2904 127 2944
rect 165 2904 167 2944
rect 171 2904 175 2944
rect 179 2924 190 2944
rect 216 2924 225 2984
rect 179 2904 181 2924
rect 193 2904 195 2924
rect 199 2904 203 2924
rect 207 2904 211 2924
rect 223 2904 225 2924
rect 229 2904 231 2984
rect 288 2904 290 2944
rect 294 2904 298 2944
rect 310 2904 312 2984
rect 316 2904 320 2984
rect 324 2904 326 2984
rect 383 2904 385 2944
rect 389 2904 391 2944
rect 403 2904 405 2944
rect 409 2904 411 2944
rect 449 2904 451 2984
rect 455 2924 464 2984
rect 632 2944 641 2984
rect 490 2924 501 2944
rect 455 2904 457 2924
rect 469 2904 473 2924
rect 477 2904 481 2924
rect 485 2904 487 2924
rect 499 2904 501 2924
rect 505 2904 509 2944
rect 513 2904 515 2944
rect 553 2904 555 2944
rect 559 2904 561 2944
rect 573 2904 575 2944
rect 579 2904 587 2944
rect 591 2904 593 2944
rect 605 2904 607 2944
rect 611 2904 621 2944
rect 625 2904 627 2944
rect 639 2904 641 2944
rect 645 2904 647 2984
rect 693 2904 695 2984
rect 699 2944 708 2984
rect 699 2904 701 2944
rect 713 2904 715 2944
rect 719 2904 729 2944
rect 733 2904 735 2944
rect 747 2904 749 2944
rect 753 2904 761 2944
rect 765 2904 767 2944
rect 779 2904 781 2944
rect 785 2904 787 2944
rect 825 2904 827 2944
rect 831 2904 835 2944
rect 839 2924 850 2944
rect 876 2924 885 2984
rect 839 2904 841 2924
rect 853 2904 855 2924
rect 859 2904 863 2924
rect 867 2904 871 2924
rect 883 2904 885 2924
rect 889 2904 891 2984
rect 929 2904 931 2944
rect 935 2904 937 2944
rect 1015 2904 1017 2984
rect 1021 2904 1025 2984
rect 1029 2904 1031 2984
rect 1083 2904 1085 2944
rect 1089 2904 1091 2944
rect 1103 2904 1105 2944
rect 1109 2904 1111 2944
rect 1154 2904 1156 2984
rect 1160 2904 1164 2984
rect 1168 2904 1170 2984
rect 1237 2976 1251 2984
rect 1182 2904 1186 2944
rect 1190 2904 1192 2944
rect 1249 2904 1251 2976
rect 1255 2972 1271 2984
rect 1255 2904 1257 2972
rect 1269 2904 1271 2972
rect 1275 2904 1277 2984
rect 1289 2904 1291 2984
rect 1295 2904 1297 2984
rect 1353 2904 1355 2984
rect 1359 2944 1368 2984
rect 1359 2904 1361 2944
rect 1373 2904 1375 2944
rect 1379 2904 1389 2944
rect 1393 2904 1395 2944
rect 1407 2904 1409 2944
rect 1413 2904 1421 2944
rect 1425 2904 1427 2944
rect 1439 2904 1441 2944
rect 1445 2904 1447 2944
rect 1485 2904 1487 2944
rect 1491 2904 1495 2944
rect 1499 2924 1510 2944
rect 1536 2924 1545 2984
rect 1499 2904 1501 2924
rect 1513 2904 1515 2924
rect 1519 2904 1523 2924
rect 1527 2904 1531 2924
rect 1543 2904 1545 2924
rect 1549 2904 1551 2984
rect 1615 2904 1617 2984
rect 1621 2904 1625 2984
rect 1629 2904 1631 2984
rect 1683 2904 1685 2944
rect 1689 2904 1691 2944
rect 1703 2904 1705 2944
rect 1709 2904 1711 2944
rect 1754 2904 1756 2984
rect 1760 2904 1764 2984
rect 1768 2904 1770 2984
rect 1782 2904 1786 2944
rect 1790 2904 1792 2944
rect 1868 2904 1870 2944
rect 1874 2904 1878 2944
rect 1890 2904 1892 2984
rect 1896 2904 1900 2984
rect 1904 2904 1906 2984
rect 1949 2904 1951 2984
rect 1955 2924 1964 2984
rect 2132 2944 2141 2984
rect 1990 2924 2001 2944
rect 1955 2904 1957 2924
rect 1969 2904 1973 2924
rect 1977 2904 1981 2924
rect 1985 2904 1987 2924
rect 1999 2904 2001 2924
rect 2005 2904 2009 2944
rect 2013 2904 2015 2944
rect 2053 2904 2055 2944
rect 2059 2904 2061 2944
rect 2073 2904 2075 2944
rect 2079 2904 2087 2944
rect 2091 2904 2093 2944
rect 2105 2904 2107 2944
rect 2111 2904 2121 2944
rect 2125 2904 2127 2944
rect 2139 2904 2141 2944
rect 2145 2904 2147 2984
rect 2215 2904 2217 2984
rect 2221 2904 2225 2984
rect 2229 2904 2231 2984
rect 2283 2904 2285 2944
rect 2289 2904 2291 2944
rect 2343 2904 2345 2944
rect 2349 2940 2365 2944
rect 2349 2904 2351 2940
rect 2363 2904 2365 2940
rect 2369 2904 2371 2944
rect 2383 2904 2385 2944
rect 2389 2904 2391 2944
rect 2443 2904 2445 2984
rect 2449 2904 2451 2984
rect 2463 2904 2465 2984
rect 2469 2972 2485 2984
rect 2469 2904 2471 2972
rect 2483 2904 2485 2972
rect 2489 2976 2503 2984
rect 2489 2904 2491 2976
rect 2543 2904 2545 2944
rect 2549 2940 2565 2944
rect 2549 2904 2551 2940
rect 2563 2904 2565 2940
rect 2569 2904 2571 2944
rect 2583 2904 2585 2944
rect 2589 2904 2591 2944
rect 2648 2904 2650 2944
rect 2654 2904 2658 2944
rect 2670 2904 2672 2984
rect 2676 2904 2680 2984
rect 2684 2904 2686 2984
rect 2755 2904 2757 2984
rect 2761 2904 2765 2984
rect 2769 2904 2771 2984
rect 2957 2982 2971 2984
rect 2809 2904 2811 2944
rect 2815 2904 2817 2944
rect 2829 2904 2831 2944
rect 2835 2904 2837 2944
rect 2889 2904 2891 2944
rect 2895 2904 2897 2944
rect 2909 2904 2911 2944
rect 2915 2904 2917 2944
rect 2969 2904 2971 2982
rect 2975 2970 2991 2984
rect 2975 2904 2977 2970
rect 2989 2904 2991 2970
rect 2995 2982 3011 2984
rect 2995 2904 2997 2982
rect 3009 2904 3011 2982
rect 3015 2916 3017 2984
rect 3029 2916 3031 2984
rect 3015 2904 3031 2916
rect 3035 2904 3037 2984
rect 3089 2904 3091 2944
rect 3095 2904 3097 2944
rect 3109 2904 3111 2944
rect 3115 2904 3117 2944
rect 3174 2904 3176 2984
rect 3180 2904 3184 2984
rect 3188 2904 3190 2984
rect 3202 2904 3206 2944
rect 3210 2904 3212 2944
rect 3269 2904 3271 2984
rect 3275 2904 3277 2984
rect 3329 2904 3331 2944
rect 3335 2904 3337 2944
rect 3349 2904 3353 2944
rect 3357 2904 3361 2944
rect 3373 2904 3375 2984
rect 3379 2904 3381 2984
rect 3441 2904 3443 2984
rect 3447 2904 3449 2984
rect 3461 2904 3465 2944
rect 3469 2904 3471 2944
rect 3521 2904 3523 2984
rect 3527 2904 3529 2984
rect 3541 2904 3545 2944
rect 3549 2904 3551 2944
rect 3589 2904 3591 2944
rect 3595 2904 3597 2944
rect 3609 2904 3611 2944
rect 3615 2904 3617 2944
rect 3674 2904 3676 2984
rect 3680 2904 3684 2984
rect 3688 2904 3690 2984
rect 3702 2904 3706 2944
rect 3710 2904 3712 2944
rect 3781 2904 3783 2984
rect 3787 2904 3789 2984
rect 3801 2904 3805 2944
rect 3809 2904 3811 2944
rect 3854 2904 3856 2984
rect 3860 2904 3864 2984
rect 3868 2904 3870 2984
rect 3882 2904 3886 2944
rect 3890 2904 3892 2944
rect 3949 2904 3951 2944
rect 3955 2904 3957 2944
rect 3969 2904 3971 2944
rect 3975 2940 3991 2944
rect 3975 2904 3977 2940
rect 3989 2904 3991 2940
rect 3995 2904 3997 2944
rect 4049 2904 4051 2944
rect 4055 2904 4059 2944
rect 4071 2904 4073 2984
rect 4077 2904 4079 2984
rect 4143 2904 4145 2984
rect 4149 2904 4151 2984
rect 4163 2904 4165 2984
rect 4169 2972 4185 2984
rect 4169 2904 4171 2972
rect 4183 2904 4185 2972
rect 4189 2976 4203 2984
rect 4189 2904 4191 2976
rect 4229 2904 4231 2944
rect 4235 2904 4237 2944
rect 4249 2904 4251 2944
rect 4255 2940 4271 2944
rect 4255 2904 4257 2940
rect 4269 2904 4271 2940
rect 4275 2904 4277 2944
rect 4343 2904 4345 2984
rect 4349 2904 4351 2984
rect 4363 2904 4365 2984
rect 4369 2972 4385 2984
rect 4369 2904 4371 2972
rect 4383 2904 4385 2972
rect 4389 2976 4403 2984
rect 4389 2904 4391 2976
rect 4443 2904 4445 2944
rect 4449 2940 4465 2944
rect 4449 2904 4451 2940
rect 4463 2904 4465 2940
rect 4469 2904 4471 2944
rect 4483 2904 4485 2944
rect 4489 2904 4491 2944
rect 4543 2904 4545 2944
rect 4549 2904 4551 2944
rect 4608 2904 4610 2944
rect 4614 2904 4618 2944
rect 4630 2904 4632 2984
rect 4636 2904 4640 2984
rect 4644 2904 4646 2984
rect 4694 2904 4696 2984
rect 4700 2904 4704 2984
rect 4708 2904 4710 2984
rect 4722 2904 4726 2944
rect 4730 2904 4732 2944
rect 33 2796 35 2876
rect 39 2836 41 2876
rect 53 2836 55 2876
rect 59 2836 69 2876
rect 73 2836 75 2876
rect 87 2836 89 2876
rect 93 2836 101 2876
rect 105 2836 107 2876
rect 119 2836 121 2876
rect 125 2836 127 2876
rect 165 2836 167 2876
rect 171 2836 175 2876
rect 179 2856 181 2876
rect 193 2856 195 2876
rect 199 2856 203 2876
rect 207 2856 211 2876
rect 223 2856 225 2876
rect 179 2836 190 2856
rect 39 2796 48 2836
rect 216 2796 225 2856
rect 229 2796 231 2876
rect 283 2796 285 2876
rect 289 2864 305 2876
rect 289 2796 291 2864
rect 303 2796 305 2864
rect 309 2798 311 2876
rect 323 2798 325 2876
rect 309 2796 325 2798
rect 329 2810 331 2876
rect 343 2810 345 2876
rect 329 2796 345 2810
rect 349 2798 351 2876
rect 389 2836 391 2876
rect 395 2836 397 2876
rect 409 2836 411 2876
rect 415 2836 417 2876
rect 488 2836 490 2876
rect 494 2836 498 2876
rect 349 2796 363 2798
rect 510 2796 512 2876
rect 516 2796 520 2876
rect 524 2796 526 2876
rect 581 2796 583 2876
rect 587 2796 589 2876
rect 601 2836 605 2876
rect 609 2836 611 2876
rect 649 2836 651 2876
rect 655 2836 657 2876
rect 669 2836 671 2876
rect 675 2836 677 2876
rect 748 2836 750 2876
rect 754 2836 758 2876
rect 770 2796 772 2876
rect 776 2796 780 2876
rect 784 2796 786 2876
rect 855 2796 857 2876
rect 861 2796 865 2876
rect 869 2796 871 2876
rect 923 2836 925 2876
rect 929 2836 931 2876
rect 943 2836 945 2876
rect 949 2836 951 2876
rect 989 2836 991 2876
rect 995 2836 997 2876
rect 1063 2836 1065 2876
rect 1069 2836 1071 2876
rect 1083 2836 1085 2876
rect 1089 2836 1091 2876
rect 1129 2796 1131 2876
rect 1135 2796 1139 2876
rect 1143 2796 1145 2876
rect 1221 2796 1223 2876
rect 1227 2796 1229 2876
rect 1241 2836 1245 2876
rect 1249 2836 1251 2876
rect 1293 2796 1295 2876
rect 1299 2836 1301 2876
rect 1313 2836 1315 2876
rect 1319 2836 1329 2876
rect 1333 2836 1335 2876
rect 1347 2836 1349 2876
rect 1353 2836 1361 2876
rect 1365 2836 1367 2876
rect 1379 2836 1381 2876
rect 1385 2836 1387 2876
rect 1425 2836 1427 2876
rect 1431 2836 1435 2876
rect 1439 2856 1441 2876
rect 1453 2856 1455 2876
rect 1459 2856 1463 2876
rect 1467 2856 1471 2876
rect 1483 2856 1485 2876
rect 1439 2836 1450 2856
rect 1299 2796 1308 2836
rect 1476 2796 1485 2856
rect 1489 2796 1491 2876
rect 1529 2836 1531 2876
rect 1535 2836 1537 2876
rect 1549 2836 1551 2876
rect 1555 2836 1557 2876
rect 1628 2836 1630 2876
rect 1634 2836 1638 2876
rect 1650 2796 1652 2876
rect 1656 2796 1660 2876
rect 1664 2796 1666 2876
rect 1728 2836 1730 2876
rect 1734 2836 1738 2876
rect 1750 2796 1752 2876
rect 1756 2796 1760 2876
rect 1764 2796 1766 2876
rect 1835 2796 1837 2876
rect 1841 2796 1845 2876
rect 1849 2796 1851 2876
rect 1903 2796 1905 2876
rect 1909 2796 1911 2876
rect 1923 2796 1925 2876
rect 1929 2808 1931 2876
rect 1943 2808 1945 2876
rect 1929 2796 1945 2808
rect 1949 2804 1951 2876
rect 1949 2796 1963 2804
rect 2001 2796 2003 2876
rect 2007 2796 2009 2876
rect 2021 2836 2025 2876
rect 2029 2836 2031 2876
rect 2083 2836 2085 2876
rect 2089 2840 2091 2876
rect 2103 2840 2105 2876
rect 2089 2836 2105 2840
rect 2109 2836 2111 2876
rect 2123 2836 2125 2876
rect 2129 2836 2131 2876
rect 2169 2836 2171 2876
rect 2175 2836 2179 2876
rect 2191 2796 2193 2876
rect 2197 2796 2199 2876
rect 2253 2796 2255 2876
rect 2259 2836 2261 2876
rect 2273 2836 2275 2876
rect 2279 2836 2289 2876
rect 2293 2836 2295 2876
rect 2307 2836 2309 2876
rect 2313 2836 2321 2876
rect 2325 2836 2327 2876
rect 2339 2836 2341 2876
rect 2345 2836 2347 2876
rect 2385 2836 2387 2876
rect 2391 2836 2395 2876
rect 2399 2856 2401 2876
rect 2413 2856 2415 2876
rect 2419 2856 2423 2876
rect 2427 2856 2431 2876
rect 2443 2856 2445 2876
rect 2399 2836 2410 2856
rect 2259 2796 2268 2836
rect 2436 2796 2445 2856
rect 2449 2796 2451 2876
rect 2508 2836 2510 2876
rect 2514 2836 2518 2876
rect 2530 2796 2532 2876
rect 2536 2796 2540 2876
rect 2544 2796 2546 2876
rect 2608 2836 2610 2876
rect 2614 2836 2618 2876
rect 2630 2796 2632 2876
rect 2636 2796 2640 2876
rect 2644 2796 2646 2876
rect 2694 2796 2696 2876
rect 2700 2796 2704 2876
rect 2708 2796 2710 2876
rect 2722 2836 2726 2876
rect 2730 2836 2732 2876
rect 2789 2836 2791 2876
rect 2795 2836 2797 2876
rect 2809 2836 2811 2876
rect 2815 2836 2817 2876
rect 2869 2836 2871 2876
rect 2875 2836 2877 2876
rect 2889 2836 2891 2876
rect 2895 2836 2897 2876
rect 2954 2796 2956 2876
rect 2960 2796 2964 2876
rect 2968 2796 2970 2876
rect 2982 2836 2986 2876
rect 2990 2836 2992 2876
rect 3054 2796 3056 2876
rect 3060 2796 3064 2876
rect 3068 2796 3070 2876
rect 3082 2836 3086 2876
rect 3090 2836 3092 2876
rect 3149 2836 3151 2876
rect 3155 2836 3157 2876
rect 3169 2836 3171 2876
rect 3175 2836 3177 2876
rect 3248 2836 3250 2876
rect 3254 2836 3258 2876
rect 3270 2796 3272 2876
rect 3276 2796 3280 2876
rect 3284 2796 3286 2876
rect 3343 2836 3345 2876
rect 3349 2836 3351 2876
rect 3363 2836 3365 2876
rect 3369 2836 3371 2876
rect 3409 2836 3411 2876
rect 3415 2836 3417 2876
rect 3429 2836 3431 2876
rect 3435 2840 3437 2876
rect 3449 2840 3451 2876
rect 3435 2836 3451 2840
rect 3455 2836 3457 2876
rect 3528 2836 3530 2876
rect 3534 2836 3538 2876
rect 3550 2796 3552 2876
rect 3556 2796 3560 2876
rect 3564 2796 3566 2876
rect 3614 2796 3616 2876
rect 3620 2796 3624 2876
rect 3628 2796 3630 2876
rect 3642 2836 3646 2876
rect 3650 2836 3652 2876
rect 3723 2836 3725 2876
rect 3729 2836 3731 2876
rect 3743 2836 3745 2876
rect 3749 2836 3751 2876
rect 3808 2836 3810 2876
rect 3814 2836 3818 2876
rect 3830 2796 3832 2876
rect 3836 2796 3840 2876
rect 3844 2796 3846 2876
rect 3889 2836 3891 2876
rect 3895 2836 3897 2876
rect 3909 2836 3911 2876
rect 3915 2840 3917 2876
rect 3929 2840 3931 2876
rect 3915 2836 3931 2840
rect 3935 2836 3937 2876
rect 3989 2836 3991 2876
rect 3995 2836 3997 2876
rect 4063 2796 4065 2876
rect 4069 2864 4085 2876
rect 4069 2796 4071 2864
rect 4083 2796 4085 2864
rect 4089 2798 4091 2876
rect 4103 2798 4105 2876
rect 4089 2796 4105 2798
rect 4109 2810 4111 2876
rect 4123 2810 4125 2876
rect 4109 2796 4125 2810
rect 4129 2798 4131 2876
rect 4169 2836 4171 2876
rect 4175 2836 4177 2876
rect 4189 2836 4191 2876
rect 4195 2840 4197 2876
rect 4209 2840 4211 2876
rect 4195 2836 4211 2840
rect 4215 2836 4217 2876
rect 4129 2796 4143 2798
rect 4274 2796 4276 2876
rect 4280 2796 4284 2876
rect 4288 2796 4290 2876
rect 4302 2836 4306 2876
rect 4310 2836 4312 2876
rect 4369 2836 4371 2876
rect 4375 2836 4377 2876
rect 4389 2836 4393 2876
rect 4397 2836 4401 2876
rect 4413 2796 4415 2876
rect 4419 2796 4421 2876
rect 4469 2798 4471 2876
rect 4457 2796 4471 2798
rect 4475 2810 4477 2876
rect 4489 2810 4491 2876
rect 4475 2796 4491 2810
rect 4495 2798 4497 2876
rect 4509 2798 4511 2876
rect 4495 2796 4511 2798
rect 4515 2864 4531 2876
rect 4515 2796 4517 2864
rect 4529 2796 4531 2864
rect 4535 2796 4537 2876
rect 4589 2836 4591 2876
rect 4595 2836 4597 2876
rect 4649 2804 4651 2876
rect 4637 2796 4651 2804
rect 4655 2808 4657 2876
rect 4669 2808 4671 2876
rect 4655 2796 4671 2808
rect 4675 2796 4677 2876
rect 4689 2796 4691 2876
rect 4695 2796 4697 2876
rect 33 2424 35 2504
rect 39 2464 48 2504
rect 39 2424 41 2464
rect 53 2424 55 2464
rect 59 2424 69 2464
rect 73 2424 75 2464
rect 87 2424 89 2464
rect 93 2424 101 2464
rect 105 2424 107 2464
rect 119 2424 121 2464
rect 125 2424 127 2464
rect 165 2424 167 2464
rect 171 2424 175 2464
rect 179 2444 190 2464
rect 216 2444 225 2504
rect 179 2424 181 2444
rect 193 2424 195 2444
rect 199 2424 203 2444
rect 207 2424 211 2444
rect 223 2424 225 2444
rect 229 2424 231 2504
rect 288 2424 290 2464
rect 294 2424 298 2464
rect 310 2424 312 2504
rect 316 2424 320 2504
rect 324 2424 326 2504
rect 369 2424 371 2464
rect 375 2424 379 2464
rect 391 2424 393 2504
rect 397 2424 399 2504
rect 449 2424 451 2464
rect 455 2424 457 2464
rect 469 2424 471 2464
rect 475 2424 477 2464
rect 548 2424 550 2464
rect 554 2424 558 2464
rect 570 2424 572 2504
rect 576 2424 580 2504
rect 584 2424 586 2504
rect 629 2424 631 2464
rect 635 2424 639 2464
rect 651 2424 653 2504
rect 657 2424 659 2504
rect 728 2424 730 2464
rect 734 2424 738 2464
rect 750 2424 752 2504
rect 756 2424 760 2504
rect 764 2424 766 2504
rect 809 2424 811 2504
rect 815 2424 819 2504
rect 823 2424 825 2504
rect 893 2424 895 2504
rect 899 2464 908 2504
rect 899 2424 901 2464
rect 913 2424 915 2464
rect 919 2424 929 2464
rect 933 2424 935 2464
rect 947 2424 949 2464
rect 953 2424 961 2464
rect 965 2424 967 2464
rect 979 2424 981 2464
rect 985 2424 987 2464
rect 1025 2424 1027 2464
rect 1031 2424 1035 2464
rect 1039 2444 1050 2464
rect 1076 2444 1085 2504
rect 1039 2424 1041 2444
rect 1053 2424 1055 2444
rect 1059 2424 1063 2444
rect 1067 2424 1071 2444
rect 1083 2424 1085 2444
rect 1089 2424 1091 2504
rect 1129 2424 1131 2464
rect 1135 2424 1137 2464
rect 1194 2424 1196 2504
rect 1200 2424 1204 2504
rect 1208 2424 1210 2504
rect 1222 2424 1226 2464
rect 1230 2424 1232 2464
rect 1289 2424 1291 2464
rect 1295 2424 1297 2464
rect 1349 2424 1351 2464
rect 1355 2424 1357 2464
rect 1369 2424 1371 2464
rect 1375 2424 1377 2464
rect 1429 2424 1431 2504
rect 1435 2444 1444 2504
rect 1612 2464 1621 2504
rect 1470 2444 1481 2464
rect 1435 2424 1437 2444
rect 1449 2424 1453 2444
rect 1457 2424 1461 2444
rect 1465 2424 1467 2444
rect 1479 2424 1481 2444
rect 1485 2424 1489 2464
rect 1493 2424 1495 2464
rect 1533 2424 1535 2464
rect 1539 2424 1541 2464
rect 1553 2424 1555 2464
rect 1559 2424 1567 2464
rect 1571 2424 1573 2464
rect 1585 2424 1587 2464
rect 1591 2424 1601 2464
rect 1605 2424 1607 2464
rect 1619 2424 1621 2464
rect 1625 2424 1627 2504
rect 1674 2424 1676 2504
rect 1680 2424 1684 2504
rect 1688 2424 1690 2504
rect 1702 2424 1706 2464
rect 1710 2424 1712 2464
rect 1769 2424 1771 2504
rect 1775 2444 1784 2504
rect 1952 2464 1961 2504
rect 1810 2444 1821 2464
rect 1775 2424 1777 2444
rect 1789 2424 1793 2444
rect 1797 2424 1801 2444
rect 1805 2424 1807 2444
rect 1819 2424 1821 2444
rect 1825 2424 1829 2464
rect 1833 2424 1835 2464
rect 1873 2424 1875 2464
rect 1879 2424 1881 2464
rect 1893 2424 1895 2464
rect 1899 2424 1907 2464
rect 1911 2424 1913 2464
rect 1925 2424 1927 2464
rect 1931 2424 1941 2464
rect 1945 2424 1947 2464
rect 1959 2424 1961 2464
rect 1965 2424 1967 2504
rect 2009 2424 2011 2504
rect 2015 2424 2017 2504
rect 2029 2424 2031 2504
rect 2035 2424 2037 2504
rect 2049 2424 2051 2504
rect 2055 2424 2057 2504
rect 2069 2424 2071 2504
rect 2075 2424 2077 2504
rect 2089 2424 2091 2504
rect 2095 2424 2097 2504
rect 2109 2424 2111 2504
rect 2115 2424 2117 2504
rect 2129 2424 2131 2504
rect 2135 2424 2137 2504
rect 2149 2424 2151 2504
rect 2155 2424 2157 2504
rect 2213 2424 2215 2504
rect 2219 2464 2228 2504
rect 2219 2424 2221 2464
rect 2233 2424 2235 2464
rect 2239 2424 2249 2464
rect 2253 2424 2255 2464
rect 2267 2424 2269 2464
rect 2273 2424 2281 2464
rect 2285 2424 2287 2464
rect 2299 2424 2301 2464
rect 2305 2424 2307 2464
rect 2345 2424 2347 2464
rect 2351 2424 2355 2464
rect 2359 2444 2370 2464
rect 2396 2444 2405 2504
rect 2359 2424 2361 2444
rect 2373 2424 2375 2444
rect 2379 2424 2383 2444
rect 2387 2424 2391 2444
rect 2403 2424 2405 2444
rect 2409 2424 2411 2504
rect 2463 2424 2465 2464
rect 2469 2424 2471 2464
rect 2483 2424 2485 2464
rect 2489 2424 2491 2464
rect 2529 2424 2531 2464
rect 2535 2424 2537 2464
rect 2608 2424 2610 2464
rect 2614 2424 2618 2464
rect 2630 2424 2632 2504
rect 2636 2424 2640 2504
rect 2644 2424 2646 2504
rect 2689 2424 2691 2464
rect 2695 2424 2697 2464
rect 2763 2424 2765 2464
rect 2769 2424 2771 2464
rect 2783 2424 2785 2464
rect 2789 2424 2791 2464
rect 2848 2424 2850 2464
rect 2854 2424 2858 2464
rect 2870 2424 2872 2504
rect 2876 2424 2880 2504
rect 2884 2424 2886 2504
rect 2929 2424 2931 2464
rect 2935 2424 2937 2464
rect 2949 2424 2953 2464
rect 2957 2424 2961 2464
rect 2973 2424 2975 2504
rect 2979 2424 2981 2504
rect 3034 2424 3036 2504
rect 3040 2424 3044 2504
rect 3048 2424 3050 2504
rect 3062 2424 3066 2464
rect 3070 2424 3072 2464
rect 3143 2424 3145 2464
rect 3149 2424 3151 2464
rect 3163 2424 3165 2464
rect 3169 2424 3171 2464
rect 3209 2424 3211 2464
rect 3215 2424 3217 2464
rect 3229 2424 3233 2464
rect 3237 2424 3241 2464
rect 3253 2424 3255 2504
rect 3259 2424 3261 2504
rect 3323 2424 3325 2464
rect 3329 2460 3345 2464
rect 3329 2424 3331 2460
rect 3343 2424 3345 2460
rect 3349 2424 3351 2464
rect 3363 2424 3365 2464
rect 3369 2424 3371 2464
rect 3409 2424 3411 2464
rect 3415 2424 3417 2464
rect 3469 2424 3471 2464
rect 3475 2424 3477 2464
rect 3489 2424 3491 2464
rect 3495 2424 3497 2464
rect 3549 2424 3551 2464
rect 3555 2424 3557 2464
rect 3569 2424 3573 2464
rect 3577 2424 3581 2464
rect 3593 2424 3595 2504
rect 3599 2424 3601 2504
rect 3649 2424 3651 2464
rect 3655 2424 3659 2464
rect 3671 2424 3673 2504
rect 3677 2424 3679 2504
rect 3729 2424 3731 2464
rect 3735 2424 3737 2464
rect 3799 2424 3801 2504
rect 3805 2424 3807 2504
rect 3819 2424 3823 2464
rect 3827 2424 3831 2464
rect 3843 2424 3845 2464
rect 3849 2424 3851 2464
rect 3903 2424 3905 2504
rect 3909 2436 3911 2504
rect 3923 2436 3925 2504
rect 3909 2424 3925 2436
rect 3929 2502 3945 2504
rect 3929 2424 3931 2502
rect 3943 2424 3945 2502
rect 3949 2490 3965 2504
rect 3949 2424 3951 2490
rect 3963 2424 3965 2490
rect 3969 2502 3983 2504
rect 3969 2424 3971 2502
rect 4023 2424 4025 2464
rect 4029 2424 4031 2464
rect 4043 2424 4045 2464
rect 4049 2424 4051 2464
rect 4103 2424 4105 2464
rect 4109 2424 4111 2464
rect 4123 2424 4125 2464
rect 4129 2424 4131 2464
rect 4174 2424 4176 2504
rect 4180 2424 4184 2504
rect 4188 2424 4190 2504
rect 4537 2496 4551 2504
rect 4202 2424 4206 2464
rect 4210 2424 4212 2464
rect 4269 2424 4271 2464
rect 4275 2424 4277 2464
rect 4289 2424 4291 2464
rect 4295 2424 4297 2464
rect 4363 2424 4365 2464
rect 4369 2460 4385 2464
rect 4369 2424 4371 2460
rect 4383 2424 4385 2460
rect 4389 2424 4391 2464
rect 4403 2424 4405 2464
rect 4409 2424 4411 2464
rect 4463 2424 4465 2464
rect 4469 2460 4485 2464
rect 4469 2424 4471 2460
rect 4483 2424 4485 2460
rect 4489 2424 4491 2464
rect 4503 2424 4505 2464
rect 4509 2424 4511 2464
rect 4549 2424 4551 2496
rect 4555 2492 4571 2504
rect 4555 2424 4557 2492
rect 4569 2424 4571 2492
rect 4575 2424 4577 2504
rect 4589 2424 4591 2504
rect 4595 2424 4597 2504
rect 4663 2424 4665 2464
rect 4669 2460 4685 2464
rect 4669 2424 4671 2460
rect 4683 2424 4685 2460
rect 4689 2424 4691 2464
rect 4703 2424 4705 2464
rect 4709 2424 4711 2464
rect 33 2316 35 2396
rect 39 2356 41 2396
rect 53 2356 55 2396
rect 59 2356 69 2396
rect 73 2356 75 2396
rect 87 2356 89 2396
rect 93 2356 101 2396
rect 105 2356 107 2396
rect 119 2356 121 2396
rect 125 2356 127 2396
rect 165 2356 167 2396
rect 171 2356 175 2396
rect 179 2376 181 2396
rect 193 2376 195 2396
rect 199 2376 203 2396
rect 207 2376 211 2396
rect 223 2376 225 2396
rect 179 2356 190 2376
rect 39 2316 48 2356
rect 216 2316 225 2376
rect 229 2316 231 2396
rect 274 2316 276 2396
rect 280 2316 284 2396
rect 288 2316 290 2396
rect 302 2356 306 2396
rect 310 2356 312 2396
rect 369 2318 371 2396
rect 357 2316 371 2318
rect 375 2330 377 2396
rect 389 2330 391 2396
rect 375 2316 391 2330
rect 395 2318 397 2396
rect 409 2318 411 2396
rect 395 2316 411 2318
rect 415 2384 431 2396
rect 415 2316 417 2384
rect 429 2316 431 2384
rect 435 2316 437 2396
rect 489 2356 491 2396
rect 495 2356 499 2396
rect 511 2316 513 2396
rect 517 2316 519 2396
rect 569 2356 571 2396
rect 575 2356 577 2396
rect 589 2356 591 2396
rect 595 2356 597 2396
rect 663 2356 665 2396
rect 669 2356 671 2396
rect 709 2316 711 2396
rect 715 2316 719 2396
rect 723 2316 725 2396
rect 803 2316 805 2396
rect 809 2316 811 2396
rect 823 2316 825 2396
rect 829 2328 831 2396
rect 843 2328 845 2396
rect 829 2316 845 2328
rect 849 2324 851 2396
rect 849 2316 863 2324
rect 889 2316 891 2396
rect 895 2316 899 2396
rect 903 2316 905 2396
rect 969 2316 971 2396
rect 975 2316 979 2396
rect 983 2316 985 2396
rect 1049 2356 1051 2396
rect 1055 2356 1057 2396
rect 1109 2316 1111 2396
rect 1115 2376 1117 2396
rect 1129 2376 1133 2396
rect 1137 2376 1141 2396
rect 1145 2376 1147 2396
rect 1159 2376 1161 2396
rect 1115 2316 1124 2376
rect 1150 2356 1161 2376
rect 1165 2356 1169 2396
rect 1173 2356 1175 2396
rect 1213 2356 1215 2396
rect 1219 2356 1221 2396
rect 1233 2356 1235 2396
rect 1239 2356 1247 2396
rect 1251 2356 1253 2396
rect 1265 2356 1267 2396
rect 1271 2356 1281 2396
rect 1285 2356 1287 2396
rect 1299 2356 1301 2396
rect 1292 2316 1301 2356
rect 1305 2316 1307 2396
rect 1354 2316 1356 2396
rect 1360 2316 1364 2396
rect 1368 2316 1370 2396
rect 1382 2356 1386 2396
rect 1390 2356 1392 2396
rect 1449 2316 1451 2396
rect 1455 2376 1457 2396
rect 1469 2376 1473 2396
rect 1477 2376 1481 2396
rect 1485 2376 1487 2396
rect 1499 2376 1501 2396
rect 1455 2316 1464 2376
rect 1490 2356 1501 2376
rect 1505 2356 1509 2396
rect 1513 2356 1515 2396
rect 1553 2356 1555 2396
rect 1559 2356 1561 2396
rect 1573 2356 1575 2396
rect 1579 2356 1587 2396
rect 1591 2356 1593 2396
rect 1605 2356 1607 2396
rect 1611 2356 1621 2396
rect 1625 2356 1627 2396
rect 1639 2356 1641 2396
rect 1632 2316 1641 2356
rect 1645 2316 1647 2396
rect 1715 2316 1717 2396
rect 1721 2316 1725 2396
rect 1729 2316 1731 2396
rect 1783 2316 1785 2396
rect 1789 2316 1791 2396
rect 1803 2316 1805 2396
rect 1809 2328 1811 2396
rect 1823 2328 1825 2396
rect 1809 2316 1825 2328
rect 1829 2324 1831 2396
rect 1829 2316 1843 2324
rect 1869 2316 1871 2396
rect 1875 2316 1877 2396
rect 1955 2316 1957 2396
rect 1961 2316 1965 2396
rect 1969 2316 1971 2396
rect 2009 2316 2011 2396
rect 2015 2316 2017 2396
rect 2029 2316 2031 2396
rect 2035 2316 2037 2396
rect 2049 2316 2051 2396
rect 2055 2316 2057 2396
rect 2069 2316 2071 2396
rect 2075 2316 2077 2396
rect 2089 2316 2091 2396
rect 2095 2316 2097 2396
rect 2109 2316 2111 2396
rect 2115 2316 2117 2396
rect 2129 2316 2131 2396
rect 2135 2316 2137 2396
rect 2149 2316 2151 2396
rect 2155 2316 2157 2396
rect 2214 2316 2216 2396
rect 2220 2316 2224 2396
rect 2228 2316 2230 2396
rect 2242 2356 2246 2396
rect 2250 2356 2252 2396
rect 2313 2316 2315 2396
rect 2319 2356 2321 2396
rect 2333 2356 2335 2396
rect 2339 2356 2349 2396
rect 2353 2356 2355 2396
rect 2367 2356 2369 2396
rect 2373 2356 2381 2396
rect 2385 2356 2387 2396
rect 2399 2356 2401 2396
rect 2405 2356 2407 2396
rect 2445 2356 2447 2396
rect 2451 2356 2455 2396
rect 2459 2376 2461 2396
rect 2473 2376 2475 2396
rect 2479 2376 2483 2396
rect 2487 2376 2491 2396
rect 2503 2376 2505 2396
rect 2459 2356 2470 2376
rect 2319 2316 2328 2356
rect 2496 2316 2505 2376
rect 2509 2316 2511 2396
rect 2563 2356 2565 2396
rect 2569 2356 2571 2396
rect 2583 2356 2585 2396
rect 2589 2356 2591 2396
rect 2629 2356 2631 2396
rect 2635 2356 2637 2396
rect 2649 2356 2651 2396
rect 2655 2356 2657 2396
rect 2709 2356 2711 2396
rect 2715 2356 2717 2396
rect 2729 2356 2731 2396
rect 2735 2356 2737 2396
rect 2808 2356 2810 2396
rect 2814 2356 2818 2396
rect 2830 2316 2832 2396
rect 2836 2316 2840 2396
rect 2844 2316 2846 2396
rect 2908 2356 2910 2396
rect 2914 2356 2918 2396
rect 2930 2316 2932 2396
rect 2936 2316 2940 2396
rect 2944 2316 2946 2396
rect 2993 2316 2995 2396
rect 2999 2356 3001 2396
rect 3013 2356 3015 2396
rect 3019 2356 3029 2396
rect 3033 2356 3035 2396
rect 3047 2356 3049 2396
rect 3053 2356 3061 2396
rect 3065 2356 3067 2396
rect 3079 2356 3081 2396
rect 3085 2356 3087 2396
rect 3125 2356 3127 2396
rect 3131 2356 3135 2396
rect 3139 2376 3141 2396
rect 3153 2376 3155 2396
rect 3159 2376 3163 2396
rect 3167 2376 3171 2396
rect 3183 2376 3185 2396
rect 3139 2356 3150 2376
rect 2999 2316 3008 2356
rect 3176 2316 3185 2376
rect 3189 2316 3191 2396
rect 3234 2316 3236 2396
rect 3240 2316 3244 2396
rect 3248 2316 3250 2396
rect 3262 2356 3266 2396
rect 3270 2356 3272 2396
rect 3329 2356 3331 2396
rect 3335 2356 3337 2396
rect 3349 2356 3351 2396
rect 3355 2356 3357 2396
rect 3409 2356 3411 2396
rect 3415 2356 3417 2396
rect 3429 2356 3431 2396
rect 3435 2356 3437 2396
rect 3503 2356 3505 2396
rect 3509 2356 3511 2396
rect 3523 2356 3525 2396
rect 3529 2356 3531 2396
rect 3583 2316 3585 2396
rect 3589 2316 3591 2396
rect 3643 2316 3645 2396
rect 3649 2316 3651 2396
rect 3703 2356 3705 2396
rect 3709 2356 3711 2396
rect 3754 2316 3756 2396
rect 3760 2316 3764 2396
rect 3768 2316 3770 2396
rect 3782 2356 3786 2396
rect 3790 2356 3792 2396
rect 3861 2316 3863 2396
rect 3867 2316 3869 2396
rect 3881 2356 3885 2396
rect 3889 2356 3891 2396
rect 3929 2316 3931 2396
rect 3935 2316 3937 2396
rect 3989 2356 3991 2396
rect 3995 2356 3997 2396
rect 4009 2356 4013 2396
rect 4017 2356 4021 2396
rect 4033 2316 4035 2396
rect 4039 2316 4041 2396
rect 4108 2356 4110 2396
rect 4114 2356 4118 2396
rect 4130 2316 4132 2396
rect 4136 2316 4140 2396
rect 4144 2316 4146 2396
rect 4203 2356 4205 2396
rect 4209 2360 4211 2396
rect 4223 2360 4225 2396
rect 4209 2356 4225 2360
rect 4229 2356 4231 2396
rect 4243 2356 4245 2396
rect 4249 2356 4251 2396
rect 4289 2324 4291 2396
rect 4277 2316 4291 2324
rect 4295 2328 4297 2396
rect 4309 2328 4311 2396
rect 4295 2316 4311 2328
rect 4315 2316 4317 2396
rect 4329 2316 4331 2396
rect 4335 2316 4337 2396
rect 4408 2356 4410 2396
rect 4414 2356 4418 2396
rect 4430 2316 4432 2396
rect 4436 2316 4440 2396
rect 4444 2316 4446 2396
rect 4494 2316 4496 2396
rect 4500 2316 4504 2396
rect 4508 2316 4510 2396
rect 4522 2356 4526 2396
rect 4530 2356 4532 2396
rect 4608 2356 4610 2396
rect 4614 2356 4618 2396
rect 4630 2316 4632 2396
rect 4636 2316 4640 2396
rect 4644 2316 4646 2396
rect 4689 2324 4691 2396
rect 4677 2316 4691 2324
rect 4695 2328 4697 2396
rect 4709 2328 4711 2396
rect 4695 2316 4711 2328
rect 4715 2316 4717 2396
rect 4729 2316 4731 2396
rect 4735 2316 4737 2396
rect 29 1944 31 2024
rect 35 1944 37 2024
rect 49 1944 51 2024
rect 55 1944 57 2024
rect 69 1944 71 2024
rect 75 1944 77 2024
rect 89 1944 91 2024
rect 95 1944 97 2024
rect 109 1944 111 2024
rect 115 1944 117 2024
rect 129 1944 131 2024
rect 135 1944 137 2024
rect 149 1944 151 2024
rect 155 1944 157 2024
rect 169 1944 171 2024
rect 175 1944 177 2024
rect 243 1944 245 1984
rect 249 1944 251 1984
rect 263 1944 265 1984
rect 269 1944 271 1984
rect 328 1944 330 1984
rect 334 1944 338 1984
rect 350 1944 352 2024
rect 356 1944 360 2024
rect 364 1944 366 2024
rect 397 2022 411 2024
rect 409 1944 411 2022
rect 415 2010 431 2024
rect 415 1944 417 2010
rect 429 1944 431 2010
rect 435 2022 451 2024
rect 435 1944 437 2022
rect 449 1944 451 2022
rect 455 1956 457 2024
rect 469 1956 471 2024
rect 455 1944 471 1956
rect 475 1944 477 2024
rect 533 1944 535 2024
rect 539 1984 548 2024
rect 539 1944 541 1984
rect 553 1944 555 1984
rect 559 1944 569 1984
rect 573 1944 575 1984
rect 587 1944 589 1984
rect 593 1944 601 1984
rect 605 1944 607 1984
rect 619 1944 621 1984
rect 625 1944 627 1984
rect 665 1944 667 1984
rect 671 1944 675 1984
rect 679 1964 690 1984
rect 716 1964 725 2024
rect 679 1944 681 1964
rect 693 1944 695 1964
rect 699 1944 703 1964
rect 707 1944 711 1964
rect 723 1944 725 1964
rect 729 1944 731 2024
rect 861 2023 875 2024
rect 783 1944 785 1984
rect 789 1944 791 1984
rect 803 1944 805 1984
rect 809 1944 811 1984
rect 873 1944 875 2023
rect 879 2023 895 2024
rect 879 1944 881 2023
rect 893 1944 895 2023
rect 899 1944 905 2024
rect 909 1944 911 2024
rect 949 1944 951 1984
rect 955 1944 957 1984
rect 969 1944 971 1984
rect 975 1944 977 1984
rect 1029 1944 1031 2024
rect 1035 1944 1039 2024
rect 1043 1944 1045 2024
rect 1114 1944 1116 2024
rect 1120 1944 1124 2024
rect 1128 1944 1130 2024
rect 1142 1944 1146 1984
rect 1150 1944 1152 1984
rect 1209 1944 1211 1984
rect 1215 1944 1217 1984
rect 1229 1944 1231 1984
rect 1235 1944 1237 1984
rect 1289 1944 1291 2024
rect 1295 1944 1299 2024
rect 1303 1944 1305 2024
rect 1369 1944 1371 2024
rect 1375 1964 1384 2024
rect 1552 1984 1561 2024
rect 1410 1964 1421 1984
rect 1375 1944 1377 1964
rect 1389 1944 1393 1964
rect 1397 1944 1401 1964
rect 1405 1944 1407 1964
rect 1419 1944 1421 1964
rect 1425 1944 1429 1984
rect 1433 1944 1435 1984
rect 1473 1944 1475 1984
rect 1479 1944 1481 1984
rect 1493 1944 1495 1984
rect 1499 1944 1507 1984
rect 1511 1944 1513 1984
rect 1525 1944 1527 1984
rect 1531 1944 1541 1984
rect 1545 1944 1547 1984
rect 1559 1944 1561 1984
rect 1565 1944 1567 2024
rect 1623 1944 1625 2024
rect 1629 1944 1631 2024
rect 1643 1944 1645 2024
rect 1649 2012 1665 2024
rect 1649 1944 1651 2012
rect 1663 1944 1665 2012
rect 1669 2016 1683 2024
rect 1669 1944 1671 2016
rect 1721 1944 1723 2024
rect 1727 1944 1729 2024
rect 1741 1944 1745 1984
rect 1749 1944 1751 1984
rect 1789 1944 1791 2024
rect 1795 1964 1804 2024
rect 1972 1984 1981 2024
rect 1830 1964 1841 1984
rect 1795 1944 1797 1964
rect 1809 1944 1813 1964
rect 1817 1944 1821 1964
rect 1825 1944 1827 1964
rect 1839 1944 1841 1964
rect 1845 1944 1849 1984
rect 1853 1944 1855 1984
rect 1893 1944 1895 1984
rect 1899 1944 1901 1984
rect 1913 1944 1915 1984
rect 1919 1944 1927 1984
rect 1931 1944 1933 1984
rect 1945 1944 1947 1984
rect 1951 1944 1961 1984
rect 1965 1944 1967 1984
rect 1979 1944 1981 1984
rect 1985 1944 1987 2024
rect 2043 1944 2045 1984
rect 2049 1944 2051 1984
rect 2103 1944 2105 1984
rect 2109 1944 2111 1984
rect 2123 1944 2125 1984
rect 2129 1944 2131 1984
rect 2169 1944 2171 1984
rect 2175 1944 2179 1984
rect 2191 1944 2193 2024
rect 2197 1944 2199 2024
rect 2249 1944 2251 1984
rect 2255 1944 2257 1984
rect 2269 1944 2271 1984
rect 2275 1944 2277 1984
rect 2348 1944 2350 1984
rect 2354 1944 2358 1984
rect 2370 1944 2372 2024
rect 2376 1944 2380 2024
rect 2384 1944 2386 2024
rect 2443 1944 2445 1984
rect 2449 1944 2451 1984
rect 2463 1944 2465 1984
rect 2469 1944 2471 1984
rect 2523 1944 2525 1984
rect 2529 1944 2531 1984
rect 2543 1944 2545 1984
rect 2549 1944 2551 1984
rect 2608 1944 2610 1984
rect 2614 1944 2618 1984
rect 2630 1944 2632 2024
rect 2636 1944 2640 2024
rect 2644 1944 2646 2024
rect 2708 1944 2710 1984
rect 2714 1944 2718 1984
rect 2730 1944 2732 2024
rect 2736 1944 2740 2024
rect 2744 1944 2746 2024
rect 2793 1944 2795 2024
rect 2799 1984 2808 2024
rect 2799 1944 2801 1984
rect 2813 1944 2815 1984
rect 2819 1944 2829 1984
rect 2833 1944 2835 1984
rect 2847 1944 2849 1984
rect 2853 1944 2861 1984
rect 2865 1944 2867 1984
rect 2879 1944 2881 1984
rect 2885 1944 2887 1984
rect 2925 1944 2927 1984
rect 2931 1944 2935 1984
rect 2939 1964 2950 1984
rect 2976 1964 2985 2024
rect 2939 1944 2941 1964
rect 2953 1944 2955 1964
rect 2959 1944 2963 1964
rect 2967 1944 2971 1964
rect 2983 1944 2985 1964
rect 2989 1944 2991 2024
rect 3029 1944 3031 1984
rect 3035 1944 3037 1984
rect 3049 1944 3053 1984
rect 3057 1944 3061 1984
rect 3073 1944 3075 2024
rect 3079 1944 3081 2024
rect 3148 1944 3150 1984
rect 3154 1944 3158 1984
rect 3170 1944 3172 2024
rect 3176 1944 3180 2024
rect 3184 1944 3186 2024
rect 3248 1944 3250 1984
rect 3254 1944 3258 1984
rect 3270 1944 3272 2024
rect 3276 1944 3280 2024
rect 3284 1944 3286 2024
rect 3329 1944 3331 1984
rect 3335 1944 3337 1984
rect 3349 1944 3351 1984
rect 3355 1944 3357 1984
rect 3428 1944 3430 1984
rect 3434 1944 3438 1984
rect 3450 1944 3452 2024
rect 3456 1944 3460 2024
rect 3464 1944 3466 2024
rect 3509 1944 3511 1984
rect 3515 1944 3517 1984
rect 3529 1944 3531 1984
rect 3535 1980 3551 1984
rect 3535 1944 3537 1980
rect 3549 1944 3551 1980
rect 3555 1944 3557 1984
rect 3609 1944 3611 1984
rect 3615 1944 3617 1984
rect 3669 1944 3671 1984
rect 3675 1944 3677 1984
rect 3689 1944 3691 1984
rect 3695 1980 3711 1984
rect 3695 1944 3697 1980
rect 3709 1944 3711 1980
rect 3715 1944 3717 1984
rect 3769 1944 3771 1984
rect 3775 1944 3777 1984
rect 3789 1944 3791 1984
rect 3795 1944 3797 1984
rect 3849 1944 3851 1984
rect 3855 1944 3859 1984
rect 3871 1944 3873 2024
rect 3877 1944 3879 2024
rect 3934 1944 3936 2024
rect 3940 1944 3944 2024
rect 3948 1944 3950 2024
rect 3962 1944 3966 1984
rect 3970 1944 3972 1984
rect 4043 1944 4045 1984
rect 4049 1944 4051 1984
rect 4063 1944 4065 1984
rect 4069 1944 4071 1984
rect 4123 1944 4125 1984
rect 4129 1944 4131 1984
rect 4143 1944 4145 1984
rect 4149 1944 4151 1984
rect 4203 1944 4205 1984
rect 4209 1944 4211 1984
rect 4223 1944 4225 1984
rect 4229 1944 4231 1984
rect 4269 1944 4271 1984
rect 4275 1944 4277 1984
rect 4289 1944 4293 1984
rect 4297 1944 4301 1984
rect 4313 1944 4315 2024
rect 4319 1944 4321 2024
rect 4357 2016 4371 2024
rect 4369 1944 4371 2016
rect 4375 2012 4391 2024
rect 4375 1944 4377 2012
rect 4389 1944 4391 2012
rect 4395 1944 4397 2024
rect 4409 1944 4411 2024
rect 4415 1944 4417 2024
rect 4483 1944 4485 2024
rect 4489 1944 4491 2024
rect 4503 1944 4505 2024
rect 4509 2012 4525 2024
rect 4509 1944 4511 2012
rect 4523 1944 4525 2012
rect 4529 2016 4543 2024
rect 4529 1944 4531 2016
rect 4569 1944 4571 1984
rect 4575 1944 4577 1984
rect 4589 1944 4591 1984
rect 4595 1980 4611 1984
rect 4595 1944 4597 1980
rect 4609 1944 4611 1980
rect 4615 1944 4617 1984
rect 4669 1944 4671 1984
rect 4675 1944 4677 1984
rect 4689 1944 4691 1984
rect 4695 1980 4711 1984
rect 4695 1944 4697 1980
rect 4709 1944 4711 1980
rect 4715 1944 4717 1984
rect 33 1836 35 1916
rect 39 1876 41 1916
rect 53 1876 55 1916
rect 59 1876 69 1916
rect 73 1876 75 1916
rect 87 1876 89 1916
rect 93 1876 101 1916
rect 105 1876 107 1916
rect 119 1876 121 1916
rect 125 1876 127 1916
rect 165 1876 167 1916
rect 171 1876 175 1916
rect 179 1896 181 1916
rect 193 1896 195 1916
rect 199 1896 203 1916
rect 207 1896 211 1916
rect 223 1896 225 1916
rect 179 1876 190 1896
rect 39 1836 48 1876
rect 216 1836 225 1896
rect 229 1836 231 1916
rect 274 1836 276 1916
rect 280 1836 284 1916
rect 288 1836 290 1916
rect 302 1876 306 1916
rect 310 1876 312 1916
rect 388 1876 390 1916
rect 394 1876 398 1916
rect 410 1836 412 1916
rect 416 1836 420 1916
rect 424 1836 426 1916
rect 488 1876 490 1916
rect 494 1876 498 1916
rect 510 1836 512 1916
rect 516 1836 520 1916
rect 524 1836 526 1916
rect 588 1876 590 1916
rect 594 1876 598 1916
rect 610 1836 612 1916
rect 616 1836 620 1916
rect 624 1836 626 1916
rect 669 1876 671 1916
rect 675 1876 677 1916
rect 729 1876 731 1916
rect 735 1876 737 1916
rect 815 1836 817 1916
rect 821 1836 825 1916
rect 829 1836 831 1916
rect 869 1876 871 1916
rect 875 1876 877 1916
rect 889 1876 891 1916
rect 895 1880 897 1916
rect 909 1880 911 1916
rect 895 1876 911 1880
rect 915 1876 917 1916
rect 973 1836 975 1916
rect 979 1876 981 1916
rect 993 1876 995 1916
rect 999 1876 1009 1916
rect 1013 1876 1015 1916
rect 1027 1876 1029 1916
rect 1033 1876 1041 1916
rect 1045 1876 1047 1916
rect 1059 1876 1061 1916
rect 1065 1876 1067 1916
rect 1105 1876 1107 1916
rect 1111 1876 1115 1916
rect 1119 1896 1121 1916
rect 1133 1896 1135 1916
rect 1139 1896 1143 1916
rect 1147 1896 1151 1916
rect 1163 1896 1165 1916
rect 1119 1876 1130 1896
rect 979 1836 988 1876
rect 1156 1836 1165 1896
rect 1169 1836 1171 1916
rect 1209 1876 1211 1916
rect 1215 1876 1217 1916
rect 1229 1876 1231 1916
rect 1235 1876 1237 1916
rect 1308 1876 1310 1916
rect 1314 1876 1318 1916
rect 1330 1836 1332 1916
rect 1336 1836 1340 1916
rect 1344 1836 1346 1916
rect 1403 1836 1405 1916
rect 1409 1836 1411 1916
rect 1423 1836 1425 1916
rect 1429 1836 1431 1916
rect 1443 1836 1445 1916
rect 1449 1836 1451 1916
rect 1463 1836 1465 1916
rect 1469 1836 1471 1916
rect 1483 1836 1485 1916
rect 1489 1836 1491 1916
rect 1503 1836 1505 1916
rect 1509 1836 1511 1916
rect 1523 1836 1525 1916
rect 1529 1836 1531 1916
rect 1543 1836 1545 1916
rect 1549 1836 1551 1916
rect 1593 1836 1595 1916
rect 1599 1876 1601 1916
rect 1613 1876 1615 1916
rect 1619 1876 1629 1916
rect 1633 1876 1635 1916
rect 1647 1876 1649 1916
rect 1653 1876 1661 1916
rect 1665 1876 1667 1916
rect 1679 1876 1681 1916
rect 1685 1876 1687 1916
rect 1725 1876 1727 1916
rect 1731 1876 1735 1916
rect 1739 1896 1741 1916
rect 1753 1896 1755 1916
rect 1759 1896 1763 1916
rect 1767 1896 1771 1916
rect 1783 1896 1785 1916
rect 1739 1876 1750 1896
rect 1599 1836 1608 1876
rect 1776 1836 1785 1896
rect 1789 1836 1791 1916
rect 1843 1836 1845 1916
rect 1849 1836 1851 1916
rect 1863 1836 1865 1916
rect 1869 1848 1871 1916
rect 1883 1848 1885 1916
rect 1869 1836 1885 1848
rect 1889 1844 1891 1916
rect 1889 1836 1903 1844
rect 1929 1836 1931 1916
rect 1935 1836 1939 1916
rect 1943 1836 1945 1916
rect 2023 1836 2025 1916
rect 2029 1836 2031 1916
rect 2043 1836 2045 1916
rect 2049 1848 2051 1916
rect 2063 1848 2065 1916
rect 2049 1836 2065 1848
rect 2069 1844 2071 1916
rect 2069 1836 2083 1844
rect 2135 1836 2137 1916
rect 2141 1836 2145 1916
rect 2149 1836 2151 1916
rect 2189 1844 2191 1916
rect 2177 1836 2191 1844
rect 2195 1848 2197 1916
rect 2209 1848 2211 1916
rect 2195 1836 2211 1848
rect 2215 1836 2217 1916
rect 2229 1836 2231 1916
rect 2235 1836 2237 1916
rect 2289 1836 2291 1916
rect 2295 1896 2297 1916
rect 2309 1896 2313 1916
rect 2317 1896 2321 1916
rect 2325 1896 2327 1916
rect 2339 1896 2341 1916
rect 2295 1836 2304 1896
rect 2330 1876 2341 1896
rect 2345 1876 2349 1916
rect 2353 1876 2355 1916
rect 2393 1876 2395 1916
rect 2399 1876 2401 1916
rect 2413 1876 2415 1916
rect 2419 1876 2427 1916
rect 2431 1876 2433 1916
rect 2445 1876 2447 1916
rect 2451 1876 2461 1916
rect 2465 1876 2467 1916
rect 2479 1876 2481 1916
rect 2472 1836 2481 1876
rect 2485 1836 2487 1916
rect 2533 1836 2535 1916
rect 2539 1876 2541 1916
rect 2553 1876 2555 1916
rect 2559 1876 2569 1916
rect 2573 1876 2575 1916
rect 2587 1876 2589 1916
rect 2593 1876 2601 1916
rect 2605 1876 2607 1916
rect 2619 1876 2621 1916
rect 2625 1876 2627 1916
rect 2665 1876 2667 1916
rect 2671 1876 2675 1916
rect 2679 1896 2681 1916
rect 2693 1896 2695 1916
rect 2699 1896 2703 1916
rect 2707 1896 2711 1916
rect 2723 1896 2725 1916
rect 2679 1876 2690 1896
rect 2539 1836 2548 1876
rect 2716 1836 2725 1896
rect 2729 1836 2731 1916
rect 2773 1836 2775 1916
rect 2779 1876 2781 1916
rect 2793 1876 2795 1916
rect 2799 1876 2809 1916
rect 2813 1876 2815 1916
rect 2827 1876 2829 1916
rect 2833 1876 2841 1916
rect 2845 1876 2847 1916
rect 2859 1876 2861 1916
rect 2865 1876 2867 1916
rect 2905 1876 2907 1916
rect 2911 1876 2915 1916
rect 2919 1896 2921 1916
rect 2933 1896 2935 1916
rect 2939 1896 2943 1916
rect 2947 1896 2951 1916
rect 2963 1896 2965 1916
rect 2919 1876 2930 1896
rect 2779 1836 2788 1876
rect 2956 1836 2965 1896
rect 2969 1836 2971 1916
rect 3023 1836 3025 1916
rect 3029 1836 3031 1916
rect 3083 1876 3085 1916
rect 3089 1876 3091 1916
rect 3103 1876 3105 1916
rect 3109 1876 3111 1916
rect 3163 1836 3165 1916
rect 3169 1836 3171 1916
rect 3209 1844 3211 1916
rect 3197 1836 3211 1844
rect 3215 1848 3217 1916
rect 3229 1848 3231 1916
rect 3215 1836 3231 1848
rect 3235 1836 3237 1916
rect 3249 1836 3251 1916
rect 3255 1836 3257 1916
rect 3309 1836 3311 1916
rect 3315 1836 3319 1916
rect 3323 1836 3325 1916
rect 3399 1836 3401 1916
rect 3405 1836 3407 1916
rect 3419 1876 3423 1916
rect 3427 1876 3431 1916
rect 3443 1876 3445 1916
rect 3449 1876 3451 1916
rect 3489 1836 3491 1916
rect 3495 1836 3497 1916
rect 3563 1836 3565 1916
rect 3569 1904 3585 1916
rect 3569 1836 3571 1904
rect 3583 1836 3585 1904
rect 3589 1838 3591 1916
rect 3603 1838 3605 1916
rect 3589 1836 3605 1838
rect 3609 1850 3611 1916
rect 3623 1850 3625 1916
rect 3609 1836 3625 1850
rect 3629 1838 3631 1916
rect 3629 1836 3643 1838
rect 3683 1836 3685 1916
rect 3689 1836 3691 1916
rect 3755 1836 3757 1916
rect 3761 1836 3765 1916
rect 3769 1836 3771 1916
rect 3809 1876 3811 1916
rect 3815 1876 3819 1916
rect 3831 1836 3833 1916
rect 3837 1836 3839 1916
rect 3889 1876 3891 1916
rect 3895 1876 3897 1916
rect 3909 1876 3913 1916
rect 3917 1876 3921 1916
rect 3933 1836 3935 1916
rect 3939 1836 3941 1916
rect 4003 1836 4005 1916
rect 4009 1904 4025 1916
rect 4009 1836 4011 1904
rect 4023 1836 4025 1904
rect 4029 1838 4031 1916
rect 4043 1838 4045 1916
rect 4029 1836 4045 1838
rect 4049 1850 4051 1916
rect 4063 1850 4065 1916
rect 4049 1836 4065 1850
rect 4069 1838 4071 1916
rect 4069 1836 4083 1838
rect 4109 1838 4111 1916
rect 4097 1836 4111 1838
rect 4115 1850 4117 1916
rect 4129 1850 4131 1916
rect 4115 1836 4131 1850
rect 4135 1838 4137 1916
rect 4149 1838 4151 1916
rect 4135 1836 4151 1838
rect 4155 1904 4171 1916
rect 4155 1836 4157 1904
rect 4169 1836 4171 1904
rect 4175 1836 4177 1916
rect 4229 1876 4231 1916
rect 4235 1876 4237 1916
rect 4249 1876 4251 1916
rect 4255 1876 4257 1916
rect 4309 1876 4311 1916
rect 4315 1876 4317 1916
rect 4329 1876 4333 1916
rect 4337 1876 4341 1916
rect 4353 1836 4355 1916
rect 4359 1836 4361 1916
rect 4409 1838 4411 1916
rect 4397 1836 4411 1838
rect 4415 1850 4417 1916
rect 4429 1850 4431 1916
rect 4415 1836 4431 1850
rect 4435 1838 4437 1916
rect 4449 1838 4451 1916
rect 4435 1836 4451 1838
rect 4455 1904 4471 1916
rect 4455 1836 4457 1904
rect 4469 1836 4471 1904
rect 4475 1836 4477 1916
rect 4543 1876 4545 1916
rect 4549 1876 4551 1916
rect 4594 1836 4596 1916
rect 4600 1836 4604 1916
rect 4608 1836 4610 1916
rect 4622 1876 4626 1916
rect 4630 1876 4632 1916
rect 4689 1876 4691 1916
rect 4695 1876 4697 1916
rect 29 1464 31 1544
rect 35 1464 37 1544
rect 49 1464 51 1544
rect 55 1464 57 1544
rect 69 1464 71 1544
rect 75 1464 77 1544
rect 89 1464 91 1544
rect 95 1464 97 1544
rect 109 1464 111 1544
rect 115 1464 117 1544
rect 129 1464 131 1544
rect 135 1464 137 1544
rect 149 1464 151 1544
rect 155 1464 157 1544
rect 169 1464 171 1544
rect 175 1464 177 1544
rect 255 1464 257 1544
rect 261 1464 265 1544
rect 269 1464 271 1544
rect 321 1464 323 1544
rect 327 1464 329 1544
rect 341 1464 345 1504
rect 349 1464 351 1504
rect 393 1464 395 1544
rect 399 1504 408 1544
rect 399 1464 401 1504
rect 413 1464 415 1504
rect 419 1464 429 1504
rect 433 1464 435 1504
rect 447 1464 449 1504
rect 453 1464 461 1504
rect 465 1464 467 1504
rect 479 1464 481 1504
rect 485 1464 487 1504
rect 525 1464 527 1504
rect 531 1464 535 1504
rect 539 1484 550 1504
rect 576 1484 585 1544
rect 539 1464 541 1484
rect 553 1464 555 1484
rect 559 1464 563 1484
rect 567 1464 571 1484
rect 583 1464 585 1484
rect 589 1464 591 1544
rect 633 1464 635 1544
rect 639 1504 648 1544
rect 639 1464 641 1504
rect 653 1464 655 1504
rect 659 1464 669 1504
rect 673 1464 675 1504
rect 687 1464 689 1504
rect 693 1464 701 1504
rect 705 1464 707 1504
rect 719 1464 721 1504
rect 725 1464 727 1504
rect 765 1464 767 1504
rect 771 1464 775 1504
rect 779 1484 790 1504
rect 816 1484 825 1544
rect 779 1464 781 1484
rect 793 1464 795 1484
rect 799 1464 803 1484
rect 807 1464 811 1484
rect 823 1464 825 1484
rect 829 1464 831 1544
rect 869 1464 871 1544
rect 875 1484 884 1544
rect 1052 1504 1061 1544
rect 910 1484 921 1504
rect 875 1464 877 1484
rect 889 1464 893 1484
rect 897 1464 901 1484
rect 905 1464 907 1484
rect 919 1464 921 1484
rect 925 1464 929 1504
rect 933 1464 935 1504
rect 973 1464 975 1504
rect 979 1464 981 1504
rect 993 1464 995 1504
rect 999 1464 1007 1504
rect 1011 1464 1013 1504
rect 1025 1464 1027 1504
rect 1031 1464 1041 1504
rect 1045 1464 1047 1504
rect 1059 1464 1061 1504
rect 1065 1464 1067 1544
rect 1123 1464 1125 1504
rect 1129 1464 1131 1504
rect 1143 1464 1145 1504
rect 1149 1464 1151 1504
rect 1208 1464 1210 1504
rect 1214 1464 1218 1504
rect 1230 1464 1232 1544
rect 1236 1464 1240 1544
rect 1244 1464 1246 1544
rect 1289 1464 1291 1544
rect 1295 1484 1304 1544
rect 1472 1504 1481 1544
rect 1330 1484 1341 1504
rect 1295 1464 1297 1484
rect 1309 1464 1313 1484
rect 1317 1464 1321 1484
rect 1325 1464 1327 1484
rect 1339 1464 1341 1484
rect 1345 1464 1349 1504
rect 1353 1464 1355 1504
rect 1393 1464 1395 1504
rect 1399 1464 1401 1504
rect 1413 1464 1415 1504
rect 1419 1464 1427 1504
rect 1431 1464 1433 1504
rect 1445 1464 1447 1504
rect 1451 1464 1461 1504
rect 1465 1464 1467 1504
rect 1479 1464 1481 1504
rect 1485 1464 1487 1544
rect 1533 1464 1535 1544
rect 1539 1504 1548 1544
rect 1539 1464 1541 1504
rect 1553 1464 1555 1504
rect 1559 1464 1569 1504
rect 1573 1464 1575 1504
rect 1587 1464 1589 1504
rect 1593 1464 1601 1504
rect 1605 1464 1607 1504
rect 1619 1464 1621 1504
rect 1625 1464 1627 1504
rect 1665 1464 1667 1504
rect 1671 1464 1675 1504
rect 1679 1484 1690 1504
rect 1716 1484 1725 1544
rect 1679 1464 1681 1484
rect 1693 1464 1695 1484
rect 1699 1464 1703 1484
rect 1707 1464 1711 1484
rect 1723 1464 1725 1484
rect 1729 1464 1731 1544
rect 1783 1464 1785 1544
rect 1789 1464 1791 1544
rect 1803 1464 1805 1544
rect 1809 1532 1825 1544
rect 1809 1464 1811 1532
rect 1823 1464 1825 1532
rect 1829 1536 1843 1544
rect 1829 1464 1831 1536
rect 1869 1464 1871 1544
rect 1875 1464 1879 1544
rect 1883 1464 1885 1544
rect 1953 1464 1955 1544
rect 1959 1504 1968 1544
rect 1959 1464 1961 1504
rect 1973 1464 1975 1504
rect 1979 1464 1989 1504
rect 1993 1464 1995 1504
rect 2007 1464 2009 1504
rect 2013 1464 2021 1504
rect 2025 1464 2027 1504
rect 2039 1464 2041 1504
rect 2045 1464 2047 1504
rect 2085 1464 2087 1504
rect 2091 1464 2095 1504
rect 2099 1484 2110 1504
rect 2136 1484 2145 1544
rect 2099 1464 2101 1484
rect 2113 1464 2115 1484
rect 2119 1464 2123 1484
rect 2127 1464 2131 1484
rect 2143 1464 2145 1484
rect 2149 1464 2151 1544
rect 2215 1464 2217 1544
rect 2221 1464 2225 1544
rect 2229 1464 2231 1544
rect 2283 1464 2285 1504
rect 2289 1464 2291 1504
rect 2303 1464 2305 1504
rect 2309 1464 2311 1504
rect 2354 1464 2356 1544
rect 2360 1464 2364 1544
rect 2368 1464 2370 1544
rect 2382 1464 2386 1504
rect 2390 1464 2392 1504
rect 2449 1464 2451 1544
rect 2455 1484 2464 1544
rect 2632 1504 2641 1544
rect 2490 1484 2501 1504
rect 2455 1464 2457 1484
rect 2469 1464 2473 1484
rect 2477 1464 2481 1484
rect 2485 1464 2487 1484
rect 2499 1464 2501 1484
rect 2505 1464 2509 1504
rect 2513 1464 2515 1504
rect 2553 1464 2555 1504
rect 2559 1464 2561 1504
rect 2573 1464 2575 1504
rect 2579 1464 2587 1504
rect 2591 1464 2593 1504
rect 2605 1464 2607 1504
rect 2611 1464 2621 1504
rect 2625 1464 2627 1504
rect 2639 1464 2641 1504
rect 2645 1464 2647 1544
rect 2693 1464 2695 1544
rect 2699 1504 2708 1544
rect 2699 1464 2701 1504
rect 2713 1464 2715 1504
rect 2719 1464 2729 1504
rect 2733 1464 2735 1504
rect 2747 1464 2749 1504
rect 2753 1464 2761 1504
rect 2765 1464 2767 1504
rect 2779 1464 2781 1504
rect 2785 1464 2787 1504
rect 2825 1464 2827 1504
rect 2831 1464 2835 1504
rect 2839 1484 2850 1504
rect 2876 1484 2885 1544
rect 2839 1464 2841 1484
rect 2853 1464 2855 1484
rect 2859 1464 2863 1484
rect 2867 1464 2871 1484
rect 2883 1464 2885 1484
rect 2889 1464 2891 1544
rect 2929 1464 2931 1544
rect 2935 1464 2937 1544
rect 2989 1464 2991 1504
rect 2995 1464 2997 1504
rect 3009 1464 3011 1504
rect 3015 1464 3017 1504
rect 3083 1464 3085 1504
rect 3089 1464 3091 1504
rect 3103 1464 3105 1504
rect 3109 1464 3111 1504
rect 3154 1464 3156 1544
rect 3160 1464 3164 1544
rect 3168 1464 3170 1544
rect 3182 1464 3186 1504
rect 3190 1464 3192 1504
rect 3249 1464 3251 1504
rect 3255 1464 3257 1504
rect 3269 1464 3271 1504
rect 3275 1464 3277 1504
rect 3343 1464 3345 1504
rect 3349 1464 3351 1504
rect 3363 1464 3365 1504
rect 3369 1464 3371 1504
rect 3428 1464 3430 1504
rect 3434 1464 3438 1504
rect 3450 1464 3452 1544
rect 3456 1464 3460 1544
rect 3464 1464 3466 1544
rect 3509 1464 3511 1504
rect 3515 1464 3517 1504
rect 3529 1464 3531 1504
rect 3535 1500 3551 1504
rect 3535 1464 3537 1500
rect 3549 1464 3551 1500
rect 3555 1464 3557 1504
rect 3633 1464 3635 1544
rect 3639 1464 3645 1544
rect 3649 1464 3651 1544
rect 3673 1464 3675 1544
rect 3679 1464 3685 1544
rect 3689 1464 3691 1544
rect 3877 1536 3891 1544
rect 3729 1464 3731 1504
rect 3735 1464 3737 1504
rect 3789 1464 3791 1504
rect 3795 1464 3797 1504
rect 3809 1464 3811 1504
rect 3815 1500 3831 1504
rect 3815 1464 3817 1500
rect 3829 1464 3831 1500
rect 3835 1464 3837 1504
rect 3889 1464 3891 1536
rect 3895 1532 3911 1544
rect 3895 1464 3897 1532
rect 3909 1464 3911 1532
rect 3915 1464 3917 1544
rect 3929 1464 3931 1544
rect 3935 1464 3937 1544
rect 3994 1464 3996 1544
rect 4000 1464 4004 1544
rect 4008 1464 4010 1544
rect 4157 1536 4171 1544
rect 4022 1464 4026 1504
rect 4030 1464 4032 1504
rect 4103 1464 4105 1504
rect 4109 1464 4111 1504
rect 4123 1464 4125 1504
rect 4129 1464 4131 1504
rect 4169 1464 4171 1536
rect 4175 1532 4191 1544
rect 4175 1464 4177 1532
rect 4189 1464 4191 1532
rect 4195 1464 4197 1544
rect 4209 1464 4211 1544
rect 4215 1464 4217 1544
rect 4274 1464 4276 1544
rect 4280 1464 4284 1544
rect 4288 1464 4290 1544
rect 4302 1464 4306 1504
rect 4310 1464 4312 1504
rect 4369 1464 4371 1504
rect 4375 1464 4377 1504
rect 4429 1464 4431 1544
rect 4435 1464 4439 1544
rect 4443 1464 4445 1544
rect 4509 1464 4511 1504
rect 4515 1464 4517 1504
rect 4529 1464 4531 1504
rect 4535 1464 4537 1504
rect 4589 1464 4591 1504
rect 4595 1464 4597 1504
rect 4609 1464 4611 1504
rect 4615 1464 4617 1504
rect 4669 1464 4671 1504
rect 4675 1464 4677 1504
rect 4689 1464 4691 1504
rect 4695 1464 4697 1504
rect 29 1356 31 1436
rect 35 1416 37 1436
rect 49 1416 53 1436
rect 57 1416 61 1436
rect 65 1416 67 1436
rect 79 1416 81 1436
rect 35 1356 44 1416
rect 70 1396 81 1416
rect 85 1396 89 1436
rect 93 1396 95 1436
rect 133 1396 135 1436
rect 139 1396 141 1436
rect 153 1396 155 1436
rect 159 1396 167 1436
rect 171 1396 173 1436
rect 185 1396 187 1436
rect 191 1396 201 1436
rect 205 1396 207 1436
rect 219 1396 221 1436
rect 212 1356 221 1396
rect 225 1356 227 1436
rect 273 1356 275 1436
rect 279 1396 281 1436
rect 293 1396 295 1436
rect 299 1396 309 1436
rect 313 1396 315 1436
rect 327 1396 329 1436
rect 333 1396 341 1436
rect 345 1396 347 1436
rect 359 1396 361 1436
rect 365 1396 367 1436
rect 405 1396 407 1436
rect 411 1396 415 1436
rect 419 1416 421 1436
rect 433 1416 435 1436
rect 439 1416 443 1436
rect 447 1416 451 1436
rect 463 1416 465 1436
rect 419 1396 430 1416
rect 279 1356 288 1396
rect 456 1356 465 1416
rect 469 1356 471 1436
rect 509 1396 511 1436
rect 515 1396 517 1436
rect 529 1396 531 1436
rect 535 1396 537 1436
rect 608 1396 610 1436
rect 614 1396 618 1436
rect 630 1356 632 1436
rect 636 1356 640 1436
rect 644 1356 646 1436
rect 708 1396 710 1436
rect 714 1396 718 1436
rect 730 1356 732 1436
rect 736 1356 740 1436
rect 744 1356 746 1436
rect 801 1356 803 1436
rect 807 1356 809 1436
rect 821 1396 825 1436
rect 829 1396 831 1436
rect 869 1396 871 1436
rect 875 1396 877 1436
rect 889 1396 891 1436
rect 895 1396 897 1436
rect 968 1396 970 1436
rect 974 1396 978 1436
rect 990 1356 992 1436
rect 996 1356 1000 1436
rect 1004 1356 1006 1436
rect 1063 1396 1065 1436
rect 1069 1396 1071 1436
rect 1109 1356 1111 1436
rect 1115 1356 1117 1436
rect 1129 1356 1131 1436
rect 1135 1356 1137 1436
rect 1149 1356 1151 1436
rect 1155 1356 1157 1436
rect 1169 1356 1171 1436
rect 1175 1356 1177 1436
rect 1243 1396 1245 1436
rect 1249 1396 1251 1436
rect 1263 1396 1265 1436
rect 1269 1396 1271 1436
rect 1328 1396 1330 1436
rect 1334 1396 1338 1436
rect 1350 1356 1352 1436
rect 1356 1356 1360 1436
rect 1364 1356 1366 1436
rect 1423 1396 1425 1436
rect 1429 1396 1431 1436
rect 1443 1396 1445 1436
rect 1449 1396 1451 1436
rect 1508 1396 1510 1436
rect 1514 1396 1518 1436
rect 1530 1356 1532 1436
rect 1536 1356 1540 1436
rect 1544 1356 1546 1436
rect 1589 1396 1591 1436
rect 1595 1396 1599 1436
rect 1611 1356 1613 1436
rect 1617 1356 1619 1436
rect 1669 1396 1671 1436
rect 1675 1396 1677 1436
rect 1689 1396 1691 1436
rect 1695 1396 1697 1436
rect 1768 1396 1770 1436
rect 1774 1396 1778 1436
rect 1790 1356 1792 1436
rect 1796 1356 1800 1436
rect 1804 1356 1806 1436
rect 1849 1356 1851 1436
rect 1855 1416 1857 1436
rect 1869 1416 1873 1436
rect 1877 1416 1881 1436
rect 1885 1416 1887 1436
rect 1899 1416 1901 1436
rect 1855 1356 1864 1416
rect 1890 1396 1901 1416
rect 1905 1396 1909 1436
rect 1913 1396 1915 1436
rect 1953 1396 1955 1436
rect 1959 1396 1961 1436
rect 1973 1396 1975 1436
rect 1979 1396 1987 1436
rect 1991 1396 1993 1436
rect 2005 1396 2007 1436
rect 2011 1396 2021 1436
rect 2025 1396 2027 1436
rect 2039 1396 2041 1436
rect 2032 1356 2041 1396
rect 2045 1356 2047 1436
rect 2089 1396 2091 1436
rect 2095 1396 2097 1436
rect 2154 1356 2156 1436
rect 2160 1356 2164 1436
rect 2168 1356 2170 1436
rect 2182 1396 2186 1436
rect 2190 1396 2192 1436
rect 2263 1396 2265 1436
rect 2269 1396 2271 1436
rect 2283 1396 2285 1436
rect 2289 1396 2291 1436
rect 2355 1356 2357 1436
rect 2361 1356 2365 1436
rect 2369 1356 2371 1436
rect 2423 1396 2425 1436
rect 2429 1396 2431 1436
rect 2469 1356 2471 1436
rect 2475 1356 2479 1436
rect 2483 1356 2485 1436
rect 2549 1356 2551 1436
rect 2555 1416 2557 1436
rect 2569 1416 2573 1436
rect 2577 1416 2581 1436
rect 2585 1416 2587 1436
rect 2599 1416 2601 1436
rect 2555 1356 2564 1416
rect 2590 1396 2601 1416
rect 2605 1396 2609 1436
rect 2613 1396 2615 1436
rect 2653 1396 2655 1436
rect 2659 1396 2661 1436
rect 2673 1396 2675 1436
rect 2679 1396 2687 1436
rect 2691 1396 2693 1436
rect 2705 1396 2707 1436
rect 2711 1396 2721 1436
rect 2725 1396 2727 1436
rect 2739 1396 2741 1436
rect 2732 1356 2741 1396
rect 2745 1356 2747 1436
rect 2789 1356 2791 1436
rect 2795 1356 2799 1436
rect 2803 1356 2805 1436
rect 2883 1356 2885 1436
rect 2889 1356 2891 1436
rect 2934 1356 2936 1436
rect 2940 1356 2944 1436
rect 2948 1356 2950 1436
rect 2962 1396 2966 1436
rect 2970 1396 2972 1436
rect 3034 1356 3036 1436
rect 3040 1356 3044 1436
rect 3048 1356 3050 1436
rect 3062 1396 3066 1436
rect 3070 1396 3072 1436
rect 3134 1356 3136 1436
rect 3140 1356 3144 1436
rect 3148 1356 3150 1436
rect 3162 1396 3166 1436
rect 3170 1396 3172 1436
rect 3229 1396 3231 1436
rect 3235 1396 3237 1436
rect 3249 1396 3253 1436
rect 3257 1396 3261 1436
rect 3273 1356 3275 1436
rect 3279 1356 3281 1436
rect 3355 1356 3357 1436
rect 3361 1356 3365 1436
rect 3369 1356 3371 1436
rect 3409 1396 3411 1436
rect 3415 1396 3417 1436
rect 3429 1396 3431 1436
rect 3435 1400 3437 1436
rect 3449 1400 3451 1436
rect 3435 1396 3451 1400
rect 3455 1396 3457 1436
rect 3528 1396 3530 1436
rect 3534 1396 3538 1436
rect 3550 1356 3552 1436
rect 3556 1356 3560 1436
rect 3564 1356 3566 1436
rect 3614 1356 3616 1436
rect 3620 1356 3624 1436
rect 3628 1356 3630 1436
rect 3642 1396 3646 1436
rect 3650 1396 3652 1436
rect 3723 1396 3725 1436
rect 3729 1396 3731 1436
rect 3743 1396 3745 1436
rect 3749 1396 3751 1436
rect 3803 1396 3805 1436
rect 3809 1396 3811 1436
rect 3823 1396 3825 1436
rect 3829 1396 3831 1436
rect 3869 1396 3871 1436
rect 3875 1396 3877 1436
rect 3889 1396 3893 1436
rect 3897 1396 3901 1436
rect 3913 1356 3915 1436
rect 3919 1356 3921 1436
rect 3988 1396 3990 1436
rect 3994 1396 3998 1436
rect 4010 1356 4012 1436
rect 4016 1356 4020 1436
rect 4024 1356 4026 1436
rect 4069 1396 4071 1436
rect 4075 1396 4077 1436
rect 4143 1396 4145 1436
rect 4149 1396 4151 1436
rect 4163 1396 4165 1436
rect 4169 1396 4171 1436
rect 4223 1396 4225 1436
rect 4229 1396 4231 1436
rect 4243 1396 4245 1436
rect 4249 1396 4251 1436
rect 4315 1356 4317 1436
rect 4321 1356 4325 1436
rect 4329 1356 4331 1436
rect 4388 1396 4390 1436
rect 4394 1396 4398 1436
rect 4410 1356 4412 1436
rect 4416 1356 4420 1436
rect 4424 1356 4426 1436
rect 4474 1356 4476 1436
rect 4480 1356 4484 1436
rect 4488 1356 4490 1436
rect 4502 1396 4506 1436
rect 4510 1396 4512 1436
rect 4583 1356 4585 1436
rect 4589 1356 4591 1436
rect 4603 1356 4605 1436
rect 4609 1368 4611 1436
rect 4623 1368 4625 1436
rect 4609 1356 4625 1368
rect 4629 1364 4631 1436
rect 4669 1396 4671 1436
rect 4675 1396 4677 1436
rect 4689 1396 4691 1436
rect 4695 1396 4697 1436
rect 4629 1356 4643 1364
rect 29 984 31 1024
rect 35 984 37 1024
rect 103 984 105 1024
rect 109 984 111 1024
rect 123 984 125 1024
rect 129 984 131 1024
rect 188 984 190 1024
rect 194 984 198 1024
rect 210 984 212 1064
rect 216 984 220 1064
rect 224 984 226 1064
rect 257 1062 271 1064
rect 269 984 271 1062
rect 275 1050 291 1064
rect 275 984 277 1050
rect 289 984 291 1050
rect 295 1062 311 1064
rect 295 984 297 1062
rect 309 984 311 1062
rect 315 996 317 1064
rect 329 996 331 1064
rect 315 984 331 996
rect 335 984 337 1064
rect 403 984 405 1064
rect 409 984 411 1064
rect 423 984 425 1064
rect 429 1052 445 1064
rect 429 984 431 1052
rect 443 984 445 1052
rect 449 1056 463 1064
rect 449 984 451 1056
rect 501 1063 515 1064
rect 513 984 515 1063
rect 519 1063 535 1064
rect 519 984 521 1063
rect 533 984 535 1063
rect 539 984 545 1064
rect 549 984 551 1064
rect 589 984 591 1064
rect 595 984 599 1064
rect 603 984 605 1064
rect 679 984 681 1064
rect 685 984 687 1064
rect 699 984 703 1024
rect 707 984 711 1024
rect 723 984 725 1024
rect 729 984 731 1024
rect 781 984 783 1064
rect 787 984 789 1064
rect 801 984 805 1024
rect 809 984 811 1024
rect 875 984 877 1064
rect 881 984 885 1064
rect 889 984 891 1064
rect 943 984 945 1024
rect 949 984 951 1024
rect 1003 984 1005 1024
rect 1009 984 1011 1024
rect 1049 984 1051 1064
rect 1055 984 1059 1064
rect 1063 984 1065 1064
rect 1129 984 1131 1024
rect 1135 984 1137 1024
rect 1215 984 1217 1064
rect 1221 984 1225 1064
rect 1229 984 1231 1064
rect 1257 1056 1271 1064
rect 1269 984 1271 1056
rect 1275 1052 1291 1064
rect 1275 984 1277 1052
rect 1289 984 1291 1052
rect 1295 984 1297 1064
rect 1309 984 1311 1064
rect 1315 984 1317 1064
rect 1373 984 1375 1064
rect 1379 1024 1388 1064
rect 1379 984 1381 1024
rect 1393 984 1395 1024
rect 1399 984 1409 1024
rect 1413 984 1415 1024
rect 1427 984 1429 1024
rect 1433 984 1441 1024
rect 1445 984 1447 1024
rect 1459 984 1461 1024
rect 1465 984 1467 1024
rect 1505 984 1507 1024
rect 1511 984 1515 1024
rect 1519 1004 1530 1024
rect 1556 1004 1565 1064
rect 1519 984 1521 1004
rect 1533 984 1535 1004
rect 1539 984 1543 1004
rect 1547 984 1551 1004
rect 1563 984 1565 1004
rect 1569 984 1571 1064
rect 1623 984 1625 1024
rect 1629 984 1631 1024
rect 1669 984 1671 1024
rect 1675 984 1677 1024
rect 1689 984 1691 1024
rect 1695 984 1697 1024
rect 1749 984 1751 1064
rect 1755 984 1759 1064
rect 1763 984 1765 1064
rect 1833 984 1835 1064
rect 1839 1024 1848 1064
rect 1839 984 1841 1024
rect 1853 984 1855 1024
rect 1859 984 1869 1024
rect 1873 984 1875 1024
rect 1887 984 1889 1024
rect 1893 984 1901 1024
rect 1905 984 1907 1024
rect 1919 984 1921 1024
rect 1925 984 1927 1024
rect 1965 984 1967 1024
rect 1971 984 1975 1024
rect 1979 1004 1990 1024
rect 2016 1004 2025 1064
rect 1979 984 1981 1004
rect 1993 984 1995 1004
rect 1999 984 2003 1004
rect 2007 984 2011 1004
rect 2023 984 2025 1004
rect 2029 984 2031 1064
rect 2083 984 2085 1024
rect 2089 984 2091 1024
rect 2129 984 2131 1064
rect 2135 984 2139 1064
rect 2143 984 2145 1064
rect 2209 984 2211 1064
rect 2215 984 2219 1064
rect 2223 984 2225 1064
rect 2303 984 2305 1024
rect 2309 984 2311 1024
rect 2349 984 2351 1064
rect 2355 1004 2364 1064
rect 2532 1024 2541 1064
rect 2390 1004 2401 1024
rect 2355 984 2357 1004
rect 2369 984 2373 1004
rect 2377 984 2381 1004
rect 2385 984 2387 1004
rect 2399 984 2401 1004
rect 2405 984 2409 1024
rect 2413 984 2415 1024
rect 2453 984 2455 1024
rect 2459 984 2461 1024
rect 2473 984 2475 1024
rect 2479 984 2487 1024
rect 2491 984 2493 1024
rect 2505 984 2507 1024
rect 2511 984 2521 1024
rect 2525 984 2527 1024
rect 2539 984 2541 1024
rect 2545 984 2547 1064
rect 2589 984 2591 1024
rect 2595 984 2597 1024
rect 2654 984 2656 1064
rect 2660 984 2664 1064
rect 2668 984 2670 1064
rect 2682 984 2686 1024
rect 2690 984 2692 1024
rect 2749 984 2751 1064
rect 2755 984 2761 1064
rect 2765 984 2767 1064
rect 2789 984 2791 1064
rect 2795 984 2801 1064
rect 2805 984 2807 1064
rect 2869 984 2871 1064
rect 2875 984 2879 1064
rect 2883 984 2885 1064
rect 2963 984 2965 1024
rect 2969 984 2971 1024
rect 2983 984 2985 1024
rect 2989 984 2991 1024
rect 3029 984 3031 1024
rect 3035 984 3037 1024
rect 3049 984 3053 1024
rect 3057 984 3061 1024
rect 3073 984 3075 1064
rect 3079 984 3081 1064
rect 3134 984 3136 1064
rect 3140 984 3144 1064
rect 3148 984 3150 1064
rect 3162 984 3166 1024
rect 3170 984 3172 1024
rect 3229 984 3231 1064
rect 3235 984 3241 1064
rect 3245 1063 3261 1064
rect 3245 984 3247 1063
rect 3259 984 3261 1063
rect 3265 1063 3279 1064
rect 3265 984 3267 1063
rect 3343 984 3345 1024
rect 3349 984 3351 1024
rect 3363 984 3365 1024
rect 3369 984 3371 1024
rect 3423 984 3425 1024
rect 3429 984 3431 1024
rect 3443 984 3445 1024
rect 3449 984 3451 1024
rect 3489 984 3491 1024
rect 3495 984 3497 1024
rect 3509 984 3511 1024
rect 3515 984 3517 1024
rect 3569 984 3571 1024
rect 3575 984 3577 1024
rect 3589 984 3591 1024
rect 3595 984 3597 1024
rect 3654 984 3656 1064
rect 3660 984 3664 1064
rect 3668 984 3670 1064
rect 3837 1056 3851 1064
rect 3682 984 3686 1024
rect 3690 984 3692 1024
rect 3763 984 3765 1024
rect 3769 1020 3785 1024
rect 3769 984 3771 1020
rect 3783 984 3785 1020
rect 3789 984 3791 1024
rect 3803 984 3805 1024
rect 3809 984 3811 1024
rect 3849 984 3851 1056
rect 3855 1052 3871 1064
rect 3855 984 3857 1052
rect 3869 984 3871 1052
rect 3875 984 3877 1064
rect 3889 984 3891 1064
rect 3895 984 3897 1064
rect 4097 1056 4111 1064
rect 3963 984 3965 1024
rect 3969 984 3971 1024
rect 4023 984 4025 1024
rect 4029 1020 4045 1024
rect 4029 984 4031 1020
rect 4043 984 4045 1020
rect 4049 984 4051 1024
rect 4063 984 4065 1024
rect 4069 984 4071 1024
rect 4109 984 4111 1056
rect 4115 1052 4131 1064
rect 4115 984 4117 1052
rect 4129 984 4131 1052
rect 4135 984 4137 1064
rect 4149 984 4151 1064
rect 4155 984 4157 1064
rect 4209 984 4211 1024
rect 4215 984 4217 1024
rect 4283 984 4285 1064
rect 4289 984 4291 1064
rect 4303 984 4305 1064
rect 4309 1052 4325 1064
rect 4309 984 4311 1052
rect 4323 984 4325 1052
rect 4329 1056 4343 1064
rect 4329 984 4331 1056
rect 4388 984 4390 1024
rect 4394 984 4398 1024
rect 4410 984 4412 1064
rect 4416 984 4420 1064
rect 4424 984 4426 1064
rect 4474 984 4476 1064
rect 4480 984 4484 1064
rect 4488 984 4490 1064
rect 4502 984 4506 1024
rect 4510 984 4512 1024
rect 4569 984 4571 1064
rect 4575 984 4579 1064
rect 4583 984 4585 1064
rect 4663 984 4665 1024
rect 4669 984 4671 1024
rect 4683 984 4685 1024
rect 4689 984 4691 1024
rect 4743 984 4745 1024
rect 4749 984 4751 1024
rect 33 876 35 956
rect 39 916 41 956
rect 53 916 55 956
rect 59 916 69 956
rect 73 916 75 956
rect 87 916 89 956
rect 93 916 101 956
rect 105 916 107 956
rect 119 916 121 956
rect 125 916 127 956
rect 165 916 167 956
rect 171 916 175 956
rect 179 936 181 956
rect 193 936 195 956
rect 199 936 203 956
rect 207 936 211 956
rect 223 936 225 956
rect 179 916 190 936
rect 39 876 48 916
rect 216 876 225 936
rect 229 876 231 956
rect 269 916 271 956
rect 275 916 277 956
rect 289 916 291 956
rect 295 916 297 956
rect 368 916 370 956
rect 374 916 378 956
rect 390 876 392 956
rect 396 876 400 956
rect 404 876 406 956
rect 453 876 455 956
rect 459 916 461 956
rect 473 916 475 956
rect 479 916 489 956
rect 493 916 495 956
rect 507 916 509 956
rect 513 916 521 956
rect 525 916 527 956
rect 539 916 541 956
rect 545 916 547 956
rect 585 916 587 956
rect 591 916 595 956
rect 599 936 601 956
rect 613 936 615 956
rect 619 936 623 956
rect 627 936 631 956
rect 643 936 645 956
rect 599 916 610 936
rect 459 876 468 916
rect 636 876 645 936
rect 649 876 651 956
rect 689 916 691 956
rect 695 916 697 956
rect 709 916 711 956
rect 715 916 717 956
rect 788 916 790 956
rect 794 916 798 956
rect 810 876 812 956
rect 816 876 820 956
rect 824 876 826 956
rect 888 916 890 956
rect 894 916 898 956
rect 910 876 912 956
rect 916 876 920 956
rect 924 876 926 956
rect 983 916 985 956
rect 989 916 991 956
rect 1055 876 1057 956
rect 1061 876 1065 956
rect 1069 876 1071 956
rect 1109 876 1111 956
rect 1115 876 1119 956
rect 1123 876 1125 956
rect 1203 916 1205 956
rect 1209 916 1211 956
rect 1223 916 1225 956
rect 1229 916 1231 956
rect 1283 916 1285 956
rect 1289 916 1291 956
rect 1303 916 1305 956
rect 1309 916 1311 956
rect 1363 916 1365 956
rect 1369 916 1371 956
rect 1383 916 1385 956
rect 1389 916 1391 956
rect 1443 876 1445 956
rect 1449 876 1451 956
rect 1463 876 1465 956
rect 1469 888 1471 956
rect 1483 888 1485 956
rect 1469 876 1485 888
rect 1489 884 1491 956
rect 1489 876 1503 884
rect 1539 876 1541 956
rect 1545 876 1547 956
rect 1559 916 1563 956
rect 1567 916 1571 956
rect 1583 916 1585 956
rect 1589 916 1591 956
rect 1629 884 1631 956
rect 1617 876 1631 884
rect 1635 888 1637 956
rect 1649 888 1651 956
rect 1635 876 1651 888
rect 1655 876 1657 956
rect 1669 876 1671 956
rect 1675 876 1677 956
rect 1729 876 1731 956
rect 1735 876 1737 956
rect 1749 876 1751 956
rect 1755 876 1757 956
rect 1769 876 1771 956
rect 1775 876 1777 956
rect 1789 876 1791 956
rect 1795 876 1797 956
rect 1809 876 1811 956
rect 1815 876 1817 956
rect 1829 876 1831 956
rect 1835 876 1837 956
rect 1849 876 1851 956
rect 1855 876 1857 956
rect 1869 876 1871 956
rect 1875 876 1877 956
rect 1943 916 1945 956
rect 1949 916 1951 956
rect 1963 916 1965 956
rect 1969 916 1971 956
rect 2035 876 2037 956
rect 2041 876 2045 956
rect 2049 876 2051 956
rect 2094 876 2096 956
rect 2100 876 2104 956
rect 2108 876 2110 956
rect 2122 916 2126 956
rect 2130 916 2132 956
rect 2194 876 2196 956
rect 2200 876 2204 956
rect 2208 876 2210 956
rect 2222 916 2226 956
rect 2230 916 2232 956
rect 2294 876 2296 956
rect 2300 876 2304 956
rect 2308 876 2310 956
rect 2322 916 2326 956
rect 2330 916 2332 956
rect 2389 916 2391 956
rect 2395 916 2397 956
rect 2409 916 2411 956
rect 2415 916 2417 956
rect 2483 916 2485 956
rect 2489 916 2491 956
rect 2529 876 2531 956
rect 2535 936 2537 956
rect 2549 936 2553 956
rect 2557 936 2561 956
rect 2565 936 2567 956
rect 2579 936 2581 956
rect 2535 876 2544 936
rect 2570 916 2581 936
rect 2585 916 2589 956
rect 2593 916 2595 956
rect 2633 916 2635 956
rect 2639 916 2641 956
rect 2653 916 2655 956
rect 2659 916 2667 956
rect 2671 916 2673 956
rect 2685 916 2687 956
rect 2691 916 2701 956
rect 2705 916 2707 956
rect 2719 916 2721 956
rect 2712 876 2721 916
rect 2725 876 2727 956
rect 2788 916 2790 956
rect 2794 916 2798 956
rect 2810 876 2812 956
rect 2816 876 2820 956
rect 2824 876 2826 956
rect 2883 916 2885 956
rect 2889 916 2891 956
rect 2929 916 2931 956
rect 2935 916 2937 956
rect 2989 916 2991 956
rect 2995 916 2997 956
rect 3009 916 3011 956
rect 3015 920 3017 956
rect 3029 920 3031 956
rect 3015 916 3031 920
rect 3035 916 3037 956
rect 3089 916 3091 956
rect 3095 916 3097 956
rect 3163 916 3165 956
rect 3169 916 3171 956
rect 3183 916 3185 956
rect 3189 916 3191 956
rect 3229 876 3231 956
rect 3235 876 3241 956
rect 3245 877 3247 956
rect 3259 877 3261 956
rect 3245 876 3261 877
rect 3265 877 3267 956
rect 3329 916 3331 956
rect 3335 916 3337 956
rect 3349 916 3351 956
rect 3355 916 3357 956
rect 3409 916 3411 956
rect 3415 916 3417 956
rect 3429 916 3431 956
rect 3435 916 3437 956
rect 3265 876 3279 877
rect 3515 876 3517 956
rect 3521 876 3525 956
rect 3529 876 3531 956
rect 3569 916 3571 956
rect 3575 916 3577 956
rect 3589 916 3591 956
rect 3595 916 3597 956
rect 3663 916 3665 956
rect 3669 920 3671 956
rect 3683 920 3685 956
rect 3669 916 3685 920
rect 3689 916 3691 956
rect 3703 916 3705 956
rect 3709 916 3711 956
rect 3763 916 3765 956
rect 3769 920 3771 956
rect 3783 920 3785 956
rect 3769 916 3785 920
rect 3789 916 3791 956
rect 3803 916 3805 956
rect 3809 916 3811 956
rect 3849 916 3851 956
rect 3855 916 3857 956
rect 3869 916 3871 956
rect 3875 916 3877 956
rect 3943 916 3945 956
rect 3949 920 3951 956
rect 3963 920 3965 956
rect 3949 916 3965 920
rect 3969 916 3971 956
rect 3983 916 3985 956
rect 3989 916 3991 956
rect 4043 916 4045 956
rect 4049 916 4051 956
rect 4108 916 4110 956
rect 4114 916 4118 956
rect 4130 876 4132 956
rect 4136 876 4140 956
rect 4144 876 4146 956
rect 4208 916 4210 956
rect 4214 916 4218 956
rect 4230 876 4232 956
rect 4236 876 4240 956
rect 4244 876 4246 956
rect 4303 876 4305 956
rect 4309 876 4311 956
rect 4323 876 4325 956
rect 4329 888 4331 956
rect 4343 888 4345 956
rect 4329 876 4345 888
rect 4349 884 4351 956
rect 4389 916 4391 956
rect 4395 916 4397 956
rect 4409 916 4411 956
rect 4415 920 4417 956
rect 4429 920 4431 956
rect 4415 916 4431 920
rect 4435 916 4437 956
rect 4503 916 4505 956
rect 4509 920 4511 956
rect 4523 920 4525 956
rect 4509 916 4525 920
rect 4529 916 4531 956
rect 4543 916 4545 956
rect 4549 916 4551 956
rect 4349 876 4363 884
rect 4603 876 4605 956
rect 4609 876 4611 956
rect 4623 876 4625 956
rect 4629 888 4631 956
rect 4643 888 4645 956
rect 4629 876 4645 888
rect 4649 884 4651 956
rect 4689 916 4691 956
rect 4695 916 4697 956
rect 4709 916 4711 956
rect 4715 920 4717 956
rect 4729 920 4731 956
rect 4715 916 4731 920
rect 4735 916 4737 956
rect 4649 876 4663 884
rect 33 504 35 584
rect 39 544 48 584
rect 39 504 41 544
rect 53 504 55 544
rect 59 504 69 544
rect 73 504 75 544
rect 87 504 89 544
rect 93 504 101 544
rect 105 504 107 544
rect 119 504 121 544
rect 125 504 127 544
rect 165 504 167 544
rect 171 504 175 544
rect 179 524 190 544
rect 216 524 225 584
rect 179 504 181 524
rect 193 504 195 524
rect 199 504 203 524
rect 207 504 211 524
rect 223 504 225 524
rect 229 504 231 584
rect 269 504 271 544
rect 275 504 277 544
rect 334 504 336 584
rect 340 504 344 584
rect 348 504 350 584
rect 362 504 366 544
rect 370 504 372 544
rect 429 504 431 544
rect 435 504 437 544
rect 449 504 451 544
rect 455 504 457 544
rect 509 504 511 544
rect 515 504 519 544
rect 531 504 533 584
rect 537 504 539 584
rect 603 504 605 544
rect 609 504 611 544
rect 649 504 651 584
rect 655 524 664 584
rect 832 544 841 584
rect 690 524 701 544
rect 655 504 657 524
rect 669 504 673 524
rect 677 504 681 524
rect 685 504 687 524
rect 699 504 701 524
rect 705 504 709 544
rect 713 504 715 544
rect 753 504 755 544
rect 759 504 761 544
rect 773 504 775 544
rect 779 504 787 544
rect 791 504 793 544
rect 805 504 807 544
rect 811 504 821 544
rect 825 504 827 544
rect 839 504 841 544
rect 845 504 847 584
rect 894 504 896 584
rect 900 504 904 584
rect 908 504 910 584
rect 922 504 926 544
rect 930 504 932 544
rect 1015 504 1017 584
rect 1021 504 1025 584
rect 1029 504 1031 584
rect 1069 504 1071 584
rect 1075 504 1081 584
rect 1085 583 1101 584
rect 1085 504 1087 583
rect 1099 504 1101 583
rect 1105 583 1119 584
rect 1105 504 1107 583
rect 1188 504 1190 544
rect 1194 504 1198 544
rect 1210 504 1212 584
rect 1216 504 1220 584
rect 1224 504 1226 584
rect 1279 504 1281 584
rect 1285 504 1287 584
rect 1299 504 1303 544
rect 1307 504 1311 544
rect 1323 504 1325 544
rect 1329 504 1331 544
rect 1369 504 1371 584
rect 1375 504 1379 584
rect 1383 504 1385 584
rect 1449 504 1451 544
rect 1455 504 1459 544
rect 1471 504 1473 584
rect 1477 504 1479 584
rect 1533 504 1535 584
rect 1539 544 1548 584
rect 1539 504 1541 544
rect 1553 504 1555 544
rect 1559 504 1569 544
rect 1573 504 1575 544
rect 1587 504 1589 544
rect 1593 504 1601 544
rect 1605 504 1607 544
rect 1619 504 1621 544
rect 1625 504 1627 544
rect 1665 504 1667 544
rect 1671 504 1675 544
rect 1679 524 1690 544
rect 1716 524 1725 584
rect 1679 504 1681 524
rect 1693 504 1695 524
rect 1699 504 1703 524
rect 1707 504 1711 524
rect 1723 504 1725 524
rect 1729 504 1731 584
rect 1769 504 1771 544
rect 1775 504 1779 544
rect 1791 504 1793 584
rect 1797 504 1799 584
rect 1875 504 1877 584
rect 1881 504 1885 584
rect 1889 504 1891 584
rect 1955 504 1957 584
rect 1961 504 1965 584
rect 1969 504 1971 584
rect 2023 504 2025 544
rect 2029 504 2031 544
rect 2069 504 2071 584
rect 2075 504 2079 584
rect 2083 504 2085 584
rect 2149 504 2151 584
rect 2155 524 2164 584
rect 2332 544 2341 584
rect 2190 524 2201 544
rect 2155 504 2157 524
rect 2169 504 2173 524
rect 2177 504 2181 524
rect 2185 504 2187 524
rect 2199 504 2201 524
rect 2205 504 2209 544
rect 2213 504 2215 544
rect 2253 504 2255 544
rect 2259 504 2261 544
rect 2273 504 2275 544
rect 2279 504 2287 544
rect 2291 504 2293 544
rect 2305 504 2307 544
rect 2311 504 2321 544
rect 2325 504 2327 544
rect 2339 504 2341 544
rect 2345 504 2347 584
rect 2377 582 2391 584
rect 2389 504 2391 582
rect 2395 570 2411 584
rect 2395 504 2397 570
rect 2409 504 2411 570
rect 2415 582 2431 584
rect 2415 504 2417 582
rect 2429 504 2431 582
rect 2435 516 2437 584
rect 2449 516 2451 584
rect 2435 504 2451 516
rect 2455 504 2457 584
rect 2521 583 2535 584
rect 2533 504 2535 583
rect 2539 583 2555 584
rect 2539 504 2541 583
rect 2553 504 2555 583
rect 2559 504 2565 584
rect 2569 504 2571 584
rect 2623 504 2625 584
rect 2629 504 2631 584
rect 2643 504 2645 584
rect 2649 572 2665 584
rect 2649 504 2651 572
rect 2663 504 2665 572
rect 2669 576 2683 584
rect 2669 504 2671 576
rect 2723 504 2725 584
rect 2729 504 2731 584
rect 2743 504 2745 584
rect 2749 572 2765 584
rect 2749 504 2751 572
rect 2763 504 2765 572
rect 2769 576 2783 584
rect 2769 504 2771 576
rect 2809 504 2811 544
rect 2815 504 2817 544
rect 2888 504 2890 544
rect 2894 504 2898 544
rect 2910 504 2912 584
rect 2916 504 2920 584
rect 2924 504 2926 584
rect 2974 504 2976 584
rect 2980 504 2984 584
rect 2988 504 2990 584
rect 3002 504 3006 544
rect 3010 504 3012 544
rect 3069 504 3071 544
rect 3075 504 3077 544
rect 3089 504 3091 544
rect 3095 504 3097 544
rect 3163 504 3165 544
rect 3169 504 3171 544
rect 3209 504 3211 544
rect 3215 504 3217 544
rect 3283 504 3285 544
rect 3289 540 3305 544
rect 3289 504 3291 540
rect 3303 504 3305 540
rect 3309 504 3311 544
rect 3323 504 3325 544
rect 3329 504 3331 544
rect 3395 504 3397 584
rect 3401 504 3405 584
rect 3409 504 3411 584
rect 3454 504 3456 584
rect 3460 504 3464 584
rect 3468 504 3470 584
rect 3537 576 3551 584
rect 3482 504 3486 544
rect 3490 504 3492 544
rect 3549 504 3551 576
rect 3555 572 3571 584
rect 3555 504 3557 572
rect 3569 504 3571 572
rect 3575 504 3577 584
rect 3589 504 3591 584
rect 3595 504 3597 584
rect 3663 504 3665 584
rect 3669 504 3671 584
rect 3683 504 3685 584
rect 3689 572 3705 584
rect 3689 504 3691 572
rect 3703 504 3705 572
rect 3709 576 3723 584
rect 3709 504 3711 576
rect 3763 504 3765 584
rect 3769 516 3771 584
rect 3783 516 3785 584
rect 3769 504 3785 516
rect 3789 582 3805 584
rect 3789 504 3791 582
rect 3803 504 3805 582
rect 3809 570 3825 584
rect 3809 504 3811 570
rect 3823 504 3825 570
rect 3829 582 3843 584
rect 3829 504 3831 582
rect 3883 504 3885 544
rect 3889 540 3905 544
rect 3889 504 3891 540
rect 3903 504 3905 540
rect 3909 504 3911 544
rect 3923 504 3925 544
rect 3929 504 3931 544
rect 3983 504 3985 544
rect 3989 540 4005 544
rect 3989 504 3991 540
rect 4003 504 4005 540
rect 4009 504 4011 544
rect 4023 504 4025 544
rect 4029 504 4031 544
rect 4069 504 4071 544
rect 4075 504 4077 544
rect 4129 504 4131 544
rect 4135 504 4137 544
rect 4149 504 4151 544
rect 4155 540 4171 544
rect 4155 504 4157 540
rect 4169 504 4171 540
rect 4175 504 4177 544
rect 4229 504 4231 544
rect 4235 504 4237 544
rect 4249 504 4251 544
rect 4255 540 4271 544
rect 4255 504 4257 540
rect 4269 504 4271 540
rect 4275 504 4277 544
rect 4343 504 4345 544
rect 4349 540 4365 544
rect 4349 504 4351 540
rect 4363 504 4365 540
rect 4369 504 4371 544
rect 4383 504 4385 544
rect 4389 504 4391 544
rect 4443 504 4445 544
rect 4449 540 4465 544
rect 4449 504 4451 540
rect 4463 504 4465 540
rect 4469 504 4471 544
rect 4483 504 4485 544
rect 4489 504 4491 544
rect 4529 504 4531 544
rect 4535 504 4537 544
rect 4608 504 4610 544
rect 4614 504 4618 544
rect 4630 504 4632 584
rect 4636 504 4640 584
rect 4644 504 4646 584
rect 4694 504 4696 584
rect 4700 504 4704 584
rect 4708 504 4710 584
rect 4722 504 4726 544
rect 4730 504 4732 544
rect 33 396 35 476
rect 39 436 41 476
rect 53 436 55 476
rect 59 436 69 476
rect 73 436 75 476
rect 87 436 89 476
rect 93 436 101 476
rect 105 436 107 476
rect 119 436 121 476
rect 125 436 127 476
rect 165 436 167 476
rect 171 436 175 476
rect 179 456 181 476
rect 193 456 195 476
rect 199 456 203 476
rect 207 456 211 476
rect 223 456 225 476
rect 179 436 190 456
rect 39 396 48 436
rect 216 396 225 456
rect 229 396 231 476
rect 269 436 271 476
rect 275 436 277 476
rect 289 436 291 476
rect 295 436 297 476
rect 368 436 370 476
rect 374 436 378 476
rect 390 396 392 476
rect 396 396 400 476
rect 404 396 406 476
rect 449 436 451 476
rect 455 436 457 476
rect 509 436 511 476
rect 515 436 517 476
rect 529 436 531 476
rect 535 436 537 476
rect 608 436 610 476
rect 614 436 618 476
rect 630 396 632 476
rect 636 396 640 476
rect 644 396 646 476
rect 694 396 696 476
rect 700 396 704 476
rect 708 396 710 476
rect 722 436 726 476
rect 730 436 732 476
rect 794 396 796 476
rect 800 396 804 476
rect 808 396 810 476
rect 822 436 826 476
rect 830 436 832 476
rect 908 436 910 476
rect 914 436 918 476
rect 930 396 932 476
rect 936 396 940 476
rect 944 396 946 476
rect 989 436 991 476
rect 995 436 997 476
rect 1049 436 1051 476
rect 1055 436 1057 476
rect 1069 436 1071 476
rect 1075 436 1077 476
rect 1143 396 1145 476
rect 1149 396 1151 476
rect 1163 396 1165 476
rect 1169 408 1171 476
rect 1183 408 1185 476
rect 1169 396 1185 408
rect 1189 404 1191 476
rect 1243 436 1245 476
rect 1249 436 1251 476
rect 1308 436 1310 476
rect 1314 436 1318 476
rect 1189 396 1203 404
rect 1330 396 1332 476
rect 1336 396 1340 476
rect 1344 396 1346 476
rect 1415 396 1417 476
rect 1421 396 1425 476
rect 1429 396 1431 476
rect 1474 396 1476 476
rect 1480 396 1484 476
rect 1488 396 1490 476
rect 1502 436 1506 476
rect 1510 436 1512 476
rect 1569 436 1571 476
rect 1575 436 1577 476
rect 1589 436 1591 476
rect 1595 436 1597 476
rect 1649 396 1651 476
rect 1655 456 1657 476
rect 1669 456 1673 476
rect 1677 456 1681 476
rect 1685 456 1687 476
rect 1699 456 1701 476
rect 1655 396 1664 456
rect 1690 436 1701 456
rect 1705 436 1709 476
rect 1713 436 1715 476
rect 1753 436 1755 476
rect 1759 436 1761 476
rect 1773 436 1775 476
rect 1779 436 1787 476
rect 1791 436 1793 476
rect 1805 436 1807 476
rect 1811 436 1821 476
rect 1825 436 1827 476
rect 1839 436 1841 476
rect 1832 396 1841 436
rect 1845 396 1847 476
rect 1903 436 1905 476
rect 1909 436 1911 476
rect 1923 436 1925 476
rect 1929 436 1931 476
rect 1988 436 1990 476
rect 1994 436 1998 476
rect 2010 396 2012 476
rect 2016 396 2020 476
rect 2024 396 2026 476
rect 2073 396 2075 476
rect 2079 436 2081 476
rect 2093 436 2095 476
rect 2099 436 2109 476
rect 2113 436 2115 476
rect 2127 436 2129 476
rect 2133 436 2141 476
rect 2145 436 2147 476
rect 2159 436 2161 476
rect 2165 436 2167 476
rect 2205 436 2207 476
rect 2211 436 2215 476
rect 2219 456 2221 476
rect 2233 456 2235 476
rect 2239 456 2243 476
rect 2247 456 2251 476
rect 2263 456 2265 476
rect 2219 436 2230 456
rect 2079 396 2088 436
rect 2256 396 2265 456
rect 2269 396 2271 476
rect 2323 436 2325 476
rect 2329 436 2331 476
rect 2369 396 2371 476
rect 2375 396 2379 476
rect 2383 396 2385 476
rect 2449 436 2451 476
rect 2455 436 2457 476
rect 2523 436 2525 476
rect 2529 436 2531 476
rect 2543 436 2545 476
rect 2549 436 2551 476
rect 2589 396 2591 476
rect 2595 456 2597 476
rect 2609 456 2613 476
rect 2617 456 2621 476
rect 2625 456 2627 476
rect 2639 456 2641 476
rect 2595 396 2604 456
rect 2630 436 2641 456
rect 2645 436 2649 476
rect 2653 436 2655 476
rect 2693 436 2695 476
rect 2699 436 2701 476
rect 2713 436 2715 476
rect 2719 436 2727 476
rect 2731 436 2733 476
rect 2745 436 2747 476
rect 2751 436 2761 476
rect 2765 436 2767 476
rect 2779 436 2781 476
rect 2772 396 2781 436
rect 2785 396 2787 476
rect 2829 436 2831 476
rect 2835 436 2837 476
rect 2849 436 2851 476
rect 2855 436 2857 476
rect 2909 398 2911 476
rect 2897 396 2911 398
rect 2915 410 2917 476
rect 2929 410 2931 476
rect 2915 396 2931 410
rect 2935 398 2937 476
rect 2949 398 2951 476
rect 2935 396 2951 398
rect 2955 464 2971 476
rect 2955 396 2957 464
rect 2969 396 2971 464
rect 2975 396 2977 476
rect 3029 396 3031 476
rect 3035 396 3039 476
rect 3043 396 3045 476
rect 3109 436 3111 476
rect 3115 436 3117 476
rect 3183 436 3185 476
rect 3189 440 3191 476
rect 3203 440 3205 476
rect 3189 436 3205 440
rect 3209 436 3211 476
rect 3223 436 3225 476
rect 3229 436 3231 476
rect 3283 436 3285 476
rect 3289 440 3291 476
rect 3303 440 3305 476
rect 3289 436 3305 440
rect 3309 436 3311 476
rect 3323 436 3325 476
rect 3329 436 3331 476
rect 3374 396 3376 476
rect 3380 396 3384 476
rect 3388 396 3390 476
rect 3402 436 3406 476
rect 3410 436 3412 476
rect 3483 436 3485 476
rect 3489 436 3491 476
rect 3529 436 3531 476
rect 3535 436 3537 476
rect 3549 436 3551 476
rect 3555 436 3557 476
rect 3609 436 3611 476
rect 3615 436 3617 476
rect 3629 436 3631 476
rect 3635 436 3637 476
rect 3694 396 3696 476
rect 3700 396 3704 476
rect 3708 396 3710 476
rect 3722 436 3726 476
rect 3730 436 3732 476
rect 3815 396 3817 476
rect 3821 396 3825 476
rect 3829 396 3831 476
rect 3895 396 3897 476
rect 3901 396 3905 476
rect 3909 396 3911 476
rect 3949 436 3951 476
rect 3955 436 3957 476
rect 3969 436 3973 476
rect 3977 436 3981 476
rect 3993 396 3995 476
rect 3999 396 4001 476
rect 4049 396 4051 476
rect 4055 396 4059 476
rect 4063 396 4065 476
rect 4143 396 4145 476
rect 4149 396 4151 476
rect 4163 396 4165 476
rect 4169 408 4171 476
rect 4183 408 4185 476
rect 4169 396 4185 408
rect 4189 404 4191 476
rect 4243 436 4245 476
rect 4249 440 4251 476
rect 4263 440 4265 476
rect 4249 436 4265 440
rect 4269 436 4271 476
rect 4283 436 4285 476
rect 4289 436 4291 476
rect 4189 396 4203 404
rect 4329 404 4331 476
rect 4317 396 4331 404
rect 4335 408 4337 476
rect 4349 408 4351 476
rect 4335 396 4351 408
rect 4355 396 4357 476
rect 4369 396 4371 476
rect 4375 396 4377 476
rect 4429 436 4431 476
rect 4435 436 4437 476
rect 4508 436 4510 476
rect 4514 436 4518 476
rect 4530 396 4532 476
rect 4536 396 4540 476
rect 4544 396 4546 476
rect 4589 436 4591 476
rect 4595 436 4597 476
rect 4649 436 4651 476
rect 4655 436 4657 476
rect 4709 436 4711 476
rect 4715 436 4717 476
rect 33 24 35 104
rect 39 64 48 104
rect 39 24 41 64
rect 53 24 55 64
rect 59 24 69 64
rect 73 24 75 64
rect 87 24 89 64
rect 93 24 101 64
rect 105 24 107 64
rect 119 24 121 64
rect 125 24 127 64
rect 165 24 167 64
rect 171 24 175 64
rect 179 44 190 64
rect 216 44 225 104
rect 179 24 181 44
rect 193 24 195 44
rect 199 24 203 44
rect 207 24 211 44
rect 223 24 225 44
rect 229 24 231 104
rect 257 102 271 104
rect 269 24 271 102
rect 275 90 291 104
rect 275 24 277 90
rect 289 24 291 90
rect 295 102 311 104
rect 295 24 297 102
rect 309 24 311 102
rect 315 36 317 104
rect 329 36 331 104
rect 315 24 331 36
rect 335 24 337 104
rect 389 24 391 104
rect 395 24 399 104
rect 403 24 405 104
rect 581 103 595 104
rect 469 24 471 64
rect 475 24 477 64
rect 489 24 491 64
rect 495 60 511 64
rect 495 24 497 60
rect 509 24 511 60
rect 515 24 517 64
rect 593 24 595 103
rect 599 103 615 104
rect 599 24 601 103
rect 613 24 615 103
rect 619 24 625 104
rect 629 24 631 104
rect 683 24 685 104
rect 689 24 691 104
rect 703 24 705 104
rect 709 92 725 104
rect 709 24 711 92
rect 723 24 725 92
rect 729 96 743 104
rect 729 24 731 96
rect 769 24 771 104
rect 775 44 784 104
rect 952 64 961 104
rect 810 44 821 64
rect 775 24 777 44
rect 789 24 793 44
rect 797 24 801 44
rect 805 24 807 44
rect 819 24 821 44
rect 825 24 829 64
rect 833 24 835 64
rect 873 24 875 64
rect 879 24 881 64
rect 893 24 895 64
rect 899 24 907 64
rect 911 24 913 64
rect 925 24 927 64
rect 931 24 941 64
rect 945 24 947 64
rect 959 24 961 64
rect 965 24 967 104
rect 1028 24 1030 64
rect 1034 24 1038 64
rect 1050 24 1052 104
rect 1056 24 1060 104
rect 1064 24 1066 104
rect 1123 24 1125 64
rect 1129 24 1131 64
rect 1195 24 1197 104
rect 1201 24 1205 104
rect 1209 24 1211 104
rect 1263 24 1265 64
rect 1269 24 1271 64
rect 1328 24 1330 64
rect 1334 24 1338 64
rect 1350 24 1352 104
rect 1356 24 1360 104
rect 1364 24 1366 104
rect 1423 24 1425 64
rect 1429 24 1431 64
rect 1483 24 1485 64
rect 1489 24 1491 64
rect 1529 24 1531 104
rect 1535 24 1539 104
rect 1543 24 1545 104
rect 1623 24 1625 104
rect 1629 24 1631 104
rect 1643 24 1645 104
rect 1649 92 1665 104
rect 1649 24 1651 92
rect 1663 24 1665 92
rect 1669 96 1683 104
rect 1669 24 1671 96
rect 1713 24 1715 104
rect 1719 64 1728 104
rect 1719 24 1721 64
rect 1733 24 1735 64
rect 1739 24 1749 64
rect 1753 24 1755 64
rect 1767 24 1769 64
rect 1773 24 1781 64
rect 1785 24 1787 64
rect 1799 24 1801 64
rect 1805 24 1807 64
rect 1845 24 1847 64
rect 1851 24 1855 64
rect 1859 44 1870 64
rect 1896 44 1905 104
rect 1859 24 1861 44
rect 1873 24 1875 44
rect 1879 24 1883 44
rect 1887 24 1891 44
rect 1903 24 1905 44
rect 1909 24 1911 104
rect 1968 24 1970 64
rect 1974 24 1978 64
rect 1990 24 1992 104
rect 1996 24 2000 104
rect 2004 24 2006 104
rect 2049 24 2051 64
rect 2055 24 2057 64
rect 2109 24 2111 104
rect 2115 24 2119 104
rect 2123 24 2125 104
rect 2189 24 2191 104
rect 2195 24 2199 104
rect 2203 24 2205 104
rect 2295 24 2297 104
rect 2301 24 2305 104
rect 2309 24 2311 104
rect 2349 24 2351 104
rect 2355 24 2359 104
rect 2363 24 2365 104
rect 2443 24 2445 64
rect 2449 24 2451 64
rect 2489 24 2491 104
rect 2495 44 2504 104
rect 2672 64 2681 104
rect 2530 44 2541 64
rect 2495 24 2497 44
rect 2509 24 2513 44
rect 2517 24 2521 44
rect 2525 24 2527 44
rect 2539 24 2541 44
rect 2545 24 2549 64
rect 2553 24 2555 64
rect 2593 24 2595 64
rect 2599 24 2601 64
rect 2613 24 2615 64
rect 2619 24 2627 64
rect 2631 24 2633 64
rect 2645 24 2647 64
rect 2651 24 2661 64
rect 2665 24 2667 64
rect 2679 24 2681 64
rect 2685 24 2687 104
rect 2729 24 2731 104
rect 2735 44 2744 104
rect 2912 64 2921 104
rect 2770 44 2781 64
rect 2735 24 2737 44
rect 2749 24 2753 44
rect 2757 24 2761 44
rect 2765 24 2767 44
rect 2779 24 2781 44
rect 2785 24 2789 64
rect 2793 24 2795 64
rect 2833 24 2835 64
rect 2839 24 2841 64
rect 2853 24 2855 64
rect 2859 24 2867 64
rect 2871 24 2873 64
rect 2885 24 2887 64
rect 2891 24 2901 64
rect 2905 24 2907 64
rect 2919 24 2921 64
rect 2925 24 2927 104
rect 2969 24 2971 104
rect 2975 24 2981 104
rect 2985 24 2987 104
rect 3009 24 3011 104
rect 3015 24 3021 104
rect 3025 24 3027 104
rect 3101 103 3115 104
rect 3113 24 3115 103
rect 3119 103 3135 104
rect 3119 24 3121 103
rect 3133 24 3135 103
rect 3139 24 3145 104
rect 3149 24 3151 104
rect 3194 24 3196 104
rect 3200 24 3204 104
rect 3208 24 3210 104
rect 3222 24 3226 64
rect 3230 24 3232 64
rect 3303 24 3305 64
rect 3309 24 3311 64
rect 3349 24 3351 64
rect 3355 24 3357 64
rect 3369 24 3371 64
rect 3375 24 3377 64
rect 3443 24 3445 64
rect 3449 60 3465 64
rect 3449 24 3451 60
rect 3463 24 3465 60
rect 3469 24 3471 64
rect 3483 24 3485 64
rect 3489 24 3491 64
rect 3543 24 3545 64
rect 3549 24 3551 64
rect 3603 24 3605 104
rect 3609 24 3611 104
rect 3623 24 3625 104
rect 3629 92 3645 104
rect 3629 24 3631 92
rect 3643 24 3645 92
rect 3649 96 3663 104
rect 3649 24 3651 96
rect 3715 24 3717 104
rect 3721 24 3725 104
rect 3729 24 3731 104
rect 3769 24 3771 64
rect 3775 24 3777 64
rect 3834 24 3836 104
rect 3840 24 3844 104
rect 3848 24 3850 104
rect 3862 24 3866 64
rect 3870 24 3872 64
rect 3929 24 3931 104
rect 3935 24 3939 104
rect 3943 24 3945 104
rect 4023 24 4025 64
rect 4029 60 4045 64
rect 4029 24 4031 60
rect 4043 24 4045 60
rect 4049 24 4051 64
rect 4063 24 4065 64
rect 4069 24 4071 64
rect 4109 24 4111 64
rect 4115 24 4117 64
rect 4129 24 4131 64
rect 4135 24 4137 64
rect 4203 24 4205 64
rect 4209 60 4225 64
rect 4209 24 4211 60
rect 4223 24 4225 60
rect 4229 24 4231 64
rect 4243 24 4245 64
rect 4249 24 4251 64
rect 4303 24 4305 64
rect 4309 24 4311 64
rect 4323 24 4325 64
rect 4329 24 4331 64
rect 4383 24 4385 64
rect 4389 60 4405 64
rect 4389 24 4391 60
rect 4403 24 4405 60
rect 4409 24 4411 64
rect 4423 24 4425 64
rect 4429 24 4431 64
rect 4469 24 4471 64
rect 4475 24 4477 64
rect 4489 24 4491 64
rect 4495 24 4497 64
rect 4549 24 4551 64
rect 4555 24 4557 64
rect 4569 24 4571 64
rect 4575 60 4591 64
rect 4575 24 4577 60
rect 4589 24 4591 60
rect 4595 24 4597 64
rect 4663 24 4665 104
rect 4669 24 4671 104
rect 4683 24 4685 104
rect 4689 92 4705 104
rect 4689 24 4691 92
rect 4703 24 4705 92
rect 4709 96 4723 104
rect 4709 24 4711 96
<< ndcontact >>
rect 29 4516 41 4556
rect 49 4516 61 4556
rect 71 4536 83 4556
rect 119 4516 131 4556
rect 149 4516 161 4556
rect 191 4516 203 4556
rect 211 4516 223 4556
rect 231 4528 243 4556
rect 251 4516 263 4556
rect 277 4536 289 4556
rect 299 4516 311 4556
rect 319 4516 331 4556
rect 371 4536 383 4556
rect 391 4536 403 4556
rect 411 4536 423 4556
rect 451 4536 463 4556
rect 471 4536 483 4556
rect 491 4536 503 4556
rect 517 4536 529 4556
rect 539 4516 551 4556
rect 559 4516 571 4556
rect 611 4536 623 4556
rect 631 4536 643 4556
rect 657 4536 669 4556
rect 677 4536 689 4556
rect 697 4536 709 4556
rect 737 4536 749 4556
rect 757 4536 769 4556
rect 797 4516 809 4556
rect 819 4536 831 4556
rect 849 4536 861 4556
rect 877 4536 889 4556
rect 903 4536 915 4556
rect 925 4536 937 4556
rect 955 4536 967 4556
rect 987 4536 999 4556
rect 1007 4516 1019 4556
rect 1037 4516 1049 4556
rect 1057 4528 1069 4556
rect 1077 4516 1089 4556
rect 1097 4516 1109 4556
rect 1137 4516 1149 4556
rect 1159 4536 1171 4556
rect 1189 4536 1201 4556
rect 1217 4536 1229 4556
rect 1243 4536 1255 4556
rect 1265 4536 1277 4556
rect 1295 4536 1307 4556
rect 1327 4536 1339 4556
rect 1347 4516 1359 4556
rect 1377 4516 1389 4556
rect 1397 4528 1409 4556
rect 1417 4516 1429 4556
rect 1437 4516 1449 4556
rect 1481 4516 1493 4556
rect 1501 4536 1513 4556
rect 1533 4536 1545 4556
rect 1563 4536 1575 4556
rect 1585 4536 1597 4556
rect 1611 4536 1623 4556
rect 1639 4536 1651 4556
rect 1669 4536 1681 4556
rect 1691 4516 1703 4556
rect 1719 4516 1731 4556
rect 1749 4516 1761 4556
rect 1797 4516 1809 4556
rect 1819 4536 1831 4556
rect 1849 4536 1861 4556
rect 1877 4536 1889 4556
rect 1903 4536 1915 4556
rect 1925 4536 1937 4556
rect 1955 4536 1967 4556
rect 1987 4536 1999 4556
rect 2007 4516 2019 4556
rect 2037 4516 2049 4556
rect 2057 4526 2069 4556
rect 2077 4516 2089 4556
rect 2097 4516 2109 4544
rect 2117 4516 2129 4556
rect 2194 4498 2206 4556
rect 2230 4496 2242 4556
rect 2271 4516 2283 4556
rect 2291 4516 2303 4556
rect 2311 4528 2323 4556
rect 2331 4516 2343 4556
rect 2371 4536 2383 4556
rect 2391 4536 2403 4556
rect 2417 4536 2429 4556
rect 2437 4536 2449 4556
rect 2457 4536 2469 4556
rect 2511 4536 2523 4556
rect 2531 4536 2543 4556
rect 2557 4516 2569 4556
rect 2577 4528 2589 4556
rect 2597 4516 2609 4556
rect 2617 4516 2629 4556
rect 2657 4536 2669 4556
rect 2679 4516 2691 4556
rect 2699 4516 2711 4556
rect 2737 4536 2749 4556
rect 2759 4516 2771 4556
rect 2779 4516 2791 4556
rect 2829 4516 2841 4556
rect 2849 4516 2861 4556
rect 2871 4536 2883 4556
rect 2934 4498 2946 4556
rect 2970 4496 2982 4556
rect 3021 4516 3033 4556
rect 3041 4516 3053 4556
rect 3071 4516 3083 4556
rect 3109 4516 3121 4556
rect 3129 4516 3141 4556
rect 3151 4536 3163 4556
rect 3214 4498 3226 4556
rect 3250 4496 3262 4556
rect 3279 4516 3291 4556
rect 3309 4516 3321 4556
rect 3360 4516 3372 4556
rect 3388 4516 3400 4556
rect 3410 4536 3422 4556
rect 3457 4536 3469 4556
rect 3477 4536 3489 4556
rect 3519 4516 3531 4556
rect 3549 4516 3561 4556
rect 3598 4496 3610 4556
rect 3634 4498 3646 4556
rect 3700 4516 3712 4556
rect 3728 4516 3740 4556
rect 3750 4536 3762 4556
rect 3797 4516 3809 4556
rect 3817 4528 3829 4556
rect 3837 4516 3849 4556
rect 3857 4516 3869 4556
rect 3911 4516 3923 4556
rect 3931 4516 3943 4556
rect 3951 4528 3963 4556
rect 3971 4516 3983 4556
rect 4034 4498 4046 4556
rect 4070 4496 4082 4556
rect 4134 4498 4146 4556
rect 4170 4496 4182 4556
rect 4200 4516 4212 4556
rect 4228 4516 4240 4556
rect 4250 4536 4262 4556
rect 4299 4516 4311 4556
rect 4329 4516 4341 4556
rect 4398 4536 4410 4556
rect 4420 4516 4432 4556
rect 4448 4516 4460 4556
rect 4491 4536 4503 4556
rect 4511 4536 4523 4556
rect 4538 4496 4550 4556
rect 4574 4498 4586 4556
rect 4638 4496 4650 4556
rect 4674 4498 4686 4556
rect 31 4104 43 4144
rect 51 4104 63 4144
rect 71 4104 83 4132
rect 91 4104 103 4144
rect 141 4104 153 4144
rect 161 4104 173 4144
rect 191 4104 203 4144
rect 217 4104 229 4124
rect 237 4104 249 4124
rect 257 4104 269 4124
rect 318 4104 330 4124
rect 340 4104 352 4144
rect 368 4104 380 4144
rect 397 4104 409 4144
rect 427 4104 439 4144
rect 447 4104 459 4144
rect 518 4104 530 4124
rect 540 4104 552 4144
rect 568 4104 580 4144
rect 598 4104 610 4164
rect 634 4104 646 4162
rect 700 4104 712 4144
rect 728 4104 740 4144
rect 750 4104 762 4124
rect 797 4104 809 4144
rect 827 4104 839 4144
rect 847 4104 859 4144
rect 911 4104 923 4144
rect 931 4104 943 4144
rect 951 4104 963 4132
rect 971 4104 983 4144
rect 1011 4104 1023 4124
rect 1031 4104 1043 4124
rect 1057 4104 1069 4124
rect 1077 4104 1089 4124
rect 1097 4104 1109 4124
rect 1137 4104 1149 4124
rect 1157 4104 1169 4124
rect 1177 4104 1189 4124
rect 1217 4104 1229 4124
rect 1237 4104 1249 4124
rect 1257 4104 1269 4124
rect 1297 4104 1309 4124
rect 1317 4104 1329 4124
rect 1357 4104 1369 4144
rect 1379 4104 1391 4124
rect 1409 4104 1421 4124
rect 1437 4104 1449 4124
rect 1463 4104 1475 4124
rect 1485 4104 1497 4124
rect 1515 4104 1527 4124
rect 1547 4104 1559 4124
rect 1567 4104 1579 4144
rect 1597 4104 1609 4144
rect 1617 4104 1629 4132
rect 1637 4104 1649 4144
rect 1657 4104 1669 4144
rect 1697 4104 1709 4124
rect 1717 4104 1729 4124
rect 1737 4104 1749 4124
rect 1791 4104 1803 4124
rect 1811 4104 1823 4124
rect 1837 4104 1849 4144
rect 1859 4104 1871 4124
rect 1889 4104 1901 4124
rect 1917 4104 1929 4124
rect 1943 4104 1955 4124
rect 1965 4104 1977 4124
rect 1995 4104 2007 4124
rect 2027 4104 2039 4124
rect 2047 4104 2059 4144
rect 2099 4104 2111 4144
rect 2129 4104 2141 4144
rect 2157 4104 2169 4124
rect 2177 4104 2189 4124
rect 2197 4104 2209 4124
rect 2217 4104 2229 4144
rect 2292 4104 2304 4144
rect 2320 4104 2332 4144
rect 2348 4104 2360 4144
rect 2379 4104 2391 4144
rect 2409 4104 2421 4144
rect 2471 4104 2483 4144
rect 2491 4104 2503 4144
rect 2511 4104 2523 4132
rect 2531 4104 2543 4144
rect 2571 4104 2583 4124
rect 2591 4104 2603 4124
rect 2611 4104 2623 4124
rect 2640 4104 2652 4144
rect 2668 4104 2680 4144
rect 2690 4104 2702 4124
rect 2758 4104 2770 4124
rect 2780 4104 2792 4144
rect 2808 4104 2820 4144
rect 2837 4104 2849 4124
rect 2859 4104 2871 4144
rect 2879 4104 2891 4144
rect 2954 4104 2966 4162
rect 2990 4104 3002 4164
rect 3054 4104 3066 4162
rect 3090 4104 3102 4164
rect 3119 4104 3131 4144
rect 3149 4104 3161 4144
rect 3211 4104 3223 4124
rect 3231 4104 3243 4124
rect 3294 4104 3306 4162
rect 3330 4104 3342 4164
rect 3394 4104 3406 4162
rect 3430 4104 3442 4164
rect 3494 4104 3506 4162
rect 3530 4104 3542 4164
rect 3594 4104 3606 4162
rect 3630 4104 3642 4164
rect 3658 4104 3670 4164
rect 3694 4104 3706 4162
rect 3760 4104 3772 4144
rect 3788 4104 3800 4144
rect 3810 4104 3822 4124
rect 3857 4104 3869 4144
rect 3877 4104 3889 4132
rect 3897 4104 3909 4144
rect 3917 4104 3929 4144
rect 3957 4104 3969 4124
rect 3977 4104 3989 4124
rect 4020 4104 4032 4144
rect 4048 4104 4060 4144
rect 4070 4104 4082 4124
rect 4154 4104 4166 4162
rect 4190 4104 4202 4164
rect 4218 4104 4230 4164
rect 4254 4104 4266 4162
rect 4320 4104 4332 4144
rect 4348 4104 4360 4144
rect 4370 4104 4382 4124
rect 4417 4104 4429 4144
rect 4437 4104 4449 4132
rect 4457 4104 4469 4144
rect 4477 4104 4489 4144
rect 4520 4104 4532 4144
rect 4548 4104 4560 4144
rect 4576 4104 4588 4144
rect 4651 4104 4663 4124
rect 4671 4104 4683 4124
rect 4691 4104 4703 4124
rect 39 4036 51 4076
rect 69 4036 81 4076
rect 119 4036 131 4076
rect 149 4036 161 4076
rect 191 4056 203 4076
rect 211 4056 223 4076
rect 231 4056 243 4076
rect 257 4036 269 4076
rect 277 4048 289 4076
rect 297 4036 309 4076
rect 317 4036 329 4076
rect 371 4056 383 4076
rect 391 4056 403 4076
rect 431 4056 443 4076
rect 451 4056 463 4076
rect 491 4056 503 4076
rect 511 4056 523 4076
rect 531 4056 543 4076
rect 557 4036 569 4076
rect 587 4036 599 4076
rect 607 4036 619 4076
rect 657 4036 669 4076
rect 677 4048 689 4076
rect 697 4036 709 4076
rect 717 4036 729 4076
rect 757 4056 769 4076
rect 777 4056 789 4076
rect 817 4036 829 4076
rect 837 4048 849 4076
rect 857 4036 869 4076
rect 877 4036 889 4076
rect 919 4036 931 4076
rect 949 4036 961 4076
rect 1011 4056 1023 4076
rect 1031 4056 1043 4076
rect 1071 4056 1083 4076
rect 1091 4056 1103 4076
rect 1111 4056 1123 4076
rect 1137 4056 1149 4076
rect 1157 4056 1169 4076
rect 1197 4056 1209 4076
rect 1217 4056 1229 4076
rect 1237 4056 1249 4076
rect 1277 4056 1289 4076
rect 1297 4056 1309 4076
rect 1351 4056 1363 4076
rect 1371 4056 1383 4076
rect 1391 4056 1403 4076
rect 1431 4056 1443 4076
rect 1451 4056 1463 4076
rect 1477 4036 1489 4076
rect 1497 4048 1509 4076
rect 1517 4036 1529 4076
rect 1537 4036 1549 4076
rect 1577 4036 1589 4076
rect 1597 4046 1609 4076
rect 1617 4036 1629 4076
rect 1637 4036 1649 4064
rect 1657 4036 1669 4076
rect 1699 4036 1711 4076
rect 1729 4036 1741 4076
rect 1798 4056 1810 4076
rect 1820 4036 1832 4076
rect 1848 4036 1860 4076
rect 1878 4016 1890 4076
rect 1914 4018 1926 4076
rect 1991 4036 2003 4076
rect 2011 4036 2023 4076
rect 2031 4048 2043 4076
rect 2051 4036 2063 4076
rect 2091 4056 2103 4076
rect 2111 4056 2123 4076
rect 2174 4018 2186 4076
rect 2210 4016 2222 4076
rect 2274 4018 2286 4076
rect 2310 4016 2322 4076
rect 2358 4056 2370 4076
rect 2380 4036 2392 4076
rect 2408 4036 2420 4076
rect 2451 4056 2463 4076
rect 2471 4056 2483 4076
rect 2511 4036 2523 4076
rect 2531 4036 2543 4076
rect 2551 4048 2563 4076
rect 2571 4036 2583 4076
rect 2634 4018 2646 4076
rect 2670 4016 2682 4076
rect 2718 4056 2730 4076
rect 2740 4036 2752 4076
rect 2768 4036 2780 4076
rect 2811 4036 2823 4076
rect 2831 4036 2843 4076
rect 2851 4048 2863 4076
rect 2871 4036 2883 4076
rect 2897 4036 2909 4076
rect 2917 4048 2929 4076
rect 2937 4036 2949 4076
rect 2957 4036 2969 4076
rect 3034 4018 3046 4076
rect 3070 4016 3082 4076
rect 3111 4056 3123 4076
rect 3131 4056 3143 4076
rect 3157 4036 3169 4076
rect 3177 4048 3189 4076
rect 3197 4036 3209 4076
rect 3217 4036 3229 4076
rect 3260 4036 3272 4076
rect 3288 4036 3300 4076
rect 3310 4056 3322 4076
rect 3357 4036 3369 4076
rect 3377 4048 3389 4076
rect 3397 4036 3409 4076
rect 3417 4036 3429 4076
rect 3471 4036 3483 4076
rect 3491 4036 3503 4076
rect 3511 4048 3523 4076
rect 3531 4036 3543 4076
rect 3571 4036 3583 4076
rect 3591 4036 3603 4076
rect 3611 4048 3623 4076
rect 3631 4036 3643 4076
rect 3678 4056 3690 4076
rect 3700 4036 3712 4076
rect 3728 4036 3740 4076
rect 3794 4018 3806 4076
rect 3830 4016 3842 4076
rect 3879 4036 3891 4076
rect 3909 4036 3921 4076
rect 3959 4036 3971 4076
rect 3989 4036 4001 4076
rect 4019 4036 4031 4076
rect 4049 4036 4061 4076
rect 4134 4018 4146 4076
rect 4170 4016 4182 4076
rect 4211 4036 4223 4076
rect 4231 4036 4243 4076
rect 4251 4048 4263 4076
rect 4271 4036 4283 4076
rect 4297 4036 4309 4076
rect 4317 4048 4329 4076
rect 4337 4036 4349 4076
rect 4357 4036 4369 4076
rect 4411 4056 4423 4076
rect 4431 4056 4443 4076
rect 4494 4018 4506 4076
rect 4530 4016 4542 4076
rect 4594 4018 4606 4076
rect 4630 4016 4642 4076
rect 4660 4036 4672 4076
rect 4688 4036 4700 4076
rect 4710 4056 4722 4076
rect 31 3624 43 3664
rect 51 3624 63 3664
rect 71 3624 83 3652
rect 91 3624 103 3664
rect 131 3624 143 3644
rect 151 3624 163 3644
rect 177 3624 189 3664
rect 199 3624 211 3644
rect 229 3624 241 3644
rect 257 3624 269 3644
rect 283 3624 295 3644
rect 305 3624 317 3644
rect 335 3624 347 3644
rect 367 3624 379 3644
rect 387 3624 399 3664
rect 431 3624 443 3664
rect 451 3624 463 3664
rect 471 3624 483 3652
rect 491 3624 503 3664
rect 517 3624 529 3664
rect 547 3624 559 3664
rect 567 3624 579 3664
rect 631 3624 643 3664
rect 651 3624 663 3644
rect 671 3624 683 3644
rect 691 3624 703 3644
rect 739 3624 751 3664
rect 769 3624 781 3664
rect 801 3624 813 3664
rect 821 3624 833 3644
rect 853 3624 865 3644
rect 883 3624 895 3644
rect 905 3624 917 3644
rect 931 3624 943 3644
rect 959 3624 971 3644
rect 989 3624 1001 3644
rect 1011 3624 1023 3664
rect 1049 3624 1061 3664
rect 1069 3624 1081 3664
rect 1091 3624 1103 3644
rect 1117 3624 1129 3664
rect 1139 3624 1151 3644
rect 1169 3624 1181 3644
rect 1197 3624 1209 3644
rect 1223 3624 1235 3644
rect 1245 3624 1257 3644
rect 1275 3624 1287 3644
rect 1307 3624 1319 3644
rect 1327 3624 1339 3664
rect 1357 3624 1369 3664
rect 1377 3624 1389 3652
rect 1397 3624 1409 3664
rect 1417 3624 1429 3664
rect 1459 3624 1471 3664
rect 1489 3624 1501 3664
rect 1539 3624 1551 3664
rect 1569 3624 1581 3664
rect 1617 3624 1629 3644
rect 1639 3624 1651 3664
rect 1659 3624 1671 3664
rect 1697 3624 1709 3664
rect 1719 3624 1731 3644
rect 1749 3624 1761 3644
rect 1777 3624 1789 3644
rect 1803 3624 1815 3644
rect 1825 3624 1837 3644
rect 1855 3624 1867 3644
rect 1887 3624 1899 3644
rect 1907 3624 1919 3664
rect 1951 3624 1963 3644
rect 1971 3624 1983 3644
rect 2018 3624 2030 3644
rect 2040 3624 2052 3664
rect 2068 3624 2080 3664
rect 2111 3624 2123 3644
rect 2131 3624 2143 3644
rect 2158 3624 2170 3684
rect 2194 3624 2206 3682
rect 2271 3624 2283 3664
rect 2291 3624 2303 3664
rect 2311 3624 2323 3652
rect 2331 3624 2343 3664
rect 2394 3624 2406 3682
rect 2430 3624 2442 3684
rect 2478 3624 2490 3644
rect 2500 3624 2512 3664
rect 2528 3624 2540 3664
rect 2594 3624 2606 3682
rect 2630 3624 2642 3684
rect 2660 3624 2672 3664
rect 2688 3624 2700 3664
rect 2710 3624 2722 3644
rect 2778 3624 2790 3644
rect 2800 3624 2812 3664
rect 2828 3624 2840 3664
rect 2871 3624 2883 3644
rect 2891 3624 2903 3644
rect 2931 3624 2943 3644
rect 2951 3624 2963 3644
rect 3014 3624 3026 3682
rect 3050 3624 3062 3684
rect 3098 3624 3110 3644
rect 3120 3624 3132 3664
rect 3148 3624 3160 3664
rect 3214 3624 3226 3682
rect 3250 3624 3262 3684
rect 3291 3624 3303 3644
rect 3311 3624 3323 3644
rect 3351 3624 3363 3664
rect 3371 3624 3383 3664
rect 3391 3624 3403 3652
rect 3411 3624 3423 3664
rect 3459 3624 3471 3664
rect 3489 3624 3501 3664
rect 3517 3624 3529 3664
rect 3547 3624 3559 3664
rect 3567 3624 3579 3664
rect 3638 3624 3650 3644
rect 3660 3624 3672 3664
rect 3688 3624 3700 3664
rect 3754 3624 3766 3682
rect 3790 3624 3802 3684
rect 3831 3624 3843 3644
rect 3851 3624 3863 3644
rect 3880 3624 3892 3664
rect 3908 3624 3920 3664
rect 3930 3624 3942 3644
rect 3991 3624 4003 3664
rect 4011 3624 4023 3664
rect 4031 3624 4043 3652
rect 4051 3624 4063 3664
rect 4077 3624 4089 3664
rect 4097 3624 4109 3652
rect 4117 3624 4129 3664
rect 4137 3624 4149 3664
rect 4180 3624 4192 3664
rect 4208 3624 4220 3664
rect 4230 3624 4242 3644
rect 4298 3624 4310 3644
rect 4320 3624 4332 3664
rect 4348 3624 4360 3664
rect 4378 3624 4390 3684
rect 4414 3624 4426 3682
rect 4491 3624 4503 3644
rect 4511 3624 4523 3644
rect 4574 3624 4586 3682
rect 4610 3624 4622 3684
rect 4638 3624 4650 3684
rect 4674 3624 4686 3682
rect 21 3556 33 3596
rect 41 3576 53 3596
rect 73 3576 85 3596
rect 103 3576 115 3596
rect 125 3576 137 3596
rect 151 3576 163 3596
rect 179 3576 191 3596
rect 209 3576 221 3596
rect 231 3556 243 3596
rect 279 3556 291 3596
rect 309 3556 321 3596
rect 351 3556 363 3596
rect 371 3556 383 3596
rect 391 3568 403 3596
rect 411 3556 423 3596
rect 459 3556 471 3596
rect 489 3556 501 3596
rect 554 3538 566 3596
rect 590 3536 602 3596
rect 631 3576 643 3596
rect 651 3576 663 3596
rect 691 3556 703 3596
rect 711 3556 723 3596
rect 731 3568 743 3596
rect 751 3556 763 3596
rect 791 3556 803 3596
rect 811 3556 823 3596
rect 831 3568 843 3596
rect 851 3556 863 3596
rect 877 3576 889 3596
rect 897 3576 909 3596
rect 951 3576 963 3596
rect 971 3576 983 3596
rect 991 3576 1003 3596
rect 1017 3556 1029 3596
rect 1039 3576 1051 3596
rect 1069 3576 1081 3596
rect 1097 3576 1109 3596
rect 1123 3576 1135 3596
rect 1145 3576 1157 3596
rect 1175 3576 1187 3596
rect 1207 3576 1219 3596
rect 1227 3556 1239 3596
rect 1257 3576 1269 3596
rect 1277 3576 1289 3596
rect 1317 3576 1329 3596
rect 1337 3576 1349 3596
rect 1357 3576 1369 3596
rect 1397 3556 1409 3596
rect 1417 3568 1429 3596
rect 1437 3556 1449 3596
rect 1457 3556 1469 3596
rect 1499 3556 1511 3596
rect 1529 3556 1541 3596
rect 1589 3556 1601 3596
rect 1609 3556 1621 3596
rect 1631 3576 1643 3596
rect 1671 3576 1683 3596
rect 1691 3576 1703 3596
rect 1717 3556 1729 3596
rect 1739 3576 1751 3596
rect 1769 3576 1781 3596
rect 1797 3576 1809 3596
rect 1823 3576 1835 3596
rect 1845 3576 1857 3596
rect 1875 3576 1887 3596
rect 1907 3576 1919 3596
rect 1927 3556 1939 3596
rect 1957 3556 1969 3596
rect 1977 3566 1989 3596
rect 1997 3556 2009 3596
rect 2017 3556 2029 3584
rect 2037 3556 2049 3596
rect 2079 3556 2091 3596
rect 2109 3556 2121 3596
rect 2178 3576 2190 3596
rect 2200 3556 2212 3596
rect 2228 3556 2240 3596
rect 2294 3538 2306 3596
rect 2330 3536 2342 3596
rect 2371 3576 2383 3596
rect 2391 3576 2403 3596
rect 2454 3538 2466 3596
rect 2490 3536 2502 3596
rect 2554 3538 2566 3596
rect 2590 3536 2602 3596
rect 2631 3556 2643 3596
rect 2651 3556 2663 3596
rect 2671 3568 2683 3596
rect 2691 3556 2703 3596
rect 2717 3556 2729 3596
rect 2737 3568 2749 3596
rect 2757 3556 2769 3596
rect 2777 3556 2789 3596
rect 2819 3556 2831 3596
rect 2849 3556 2861 3596
rect 2897 3556 2909 3596
rect 2917 3568 2929 3596
rect 2937 3556 2949 3596
rect 2957 3556 2969 3596
rect 2997 3576 3009 3596
rect 3017 3576 3029 3596
rect 3037 3576 3049 3596
rect 3091 3556 3103 3596
rect 3111 3556 3123 3596
rect 3131 3568 3143 3596
rect 3151 3556 3163 3596
rect 3180 3556 3192 3596
rect 3208 3556 3220 3596
rect 3236 3556 3248 3596
rect 3299 3556 3311 3596
rect 3329 3556 3341 3596
rect 3379 3556 3391 3596
rect 3409 3556 3421 3596
rect 3459 3556 3471 3596
rect 3489 3556 3501 3596
rect 3537 3576 3549 3596
rect 3557 3576 3569 3596
rect 3577 3576 3589 3596
rect 3619 3556 3631 3596
rect 3649 3556 3661 3596
rect 3699 3556 3711 3596
rect 3729 3556 3741 3596
rect 3799 3556 3811 3596
rect 3829 3556 3841 3596
rect 3871 3576 3883 3596
rect 3891 3576 3903 3596
rect 3911 3576 3923 3596
rect 3939 3556 3951 3596
rect 3969 3556 3981 3596
rect 4019 3556 4031 3596
rect 4049 3556 4061 3596
rect 4097 3556 4109 3596
rect 4117 3568 4129 3596
rect 4137 3556 4149 3596
rect 4157 3556 4169 3596
rect 4234 3538 4246 3596
rect 4270 3536 4282 3596
rect 4298 3536 4310 3596
rect 4334 3538 4346 3596
rect 4400 3556 4412 3596
rect 4428 3556 4440 3596
rect 4450 3576 4462 3596
rect 4497 3576 4509 3596
rect 4517 3576 4529 3596
rect 4594 3538 4606 3596
rect 4630 3536 4642 3596
rect 4658 3536 4670 3596
rect 4694 3538 4706 3596
rect 21 3144 33 3184
rect 41 3144 53 3164
rect 73 3144 85 3164
rect 103 3144 115 3164
rect 125 3144 137 3164
rect 151 3144 163 3164
rect 179 3144 191 3164
rect 209 3144 221 3164
rect 231 3144 243 3184
rect 292 3144 304 3184
rect 320 3144 332 3184
rect 348 3144 360 3184
rect 379 3144 391 3184
rect 409 3144 421 3184
rect 457 3144 469 3184
rect 477 3144 489 3172
rect 497 3144 509 3184
rect 517 3144 529 3184
rect 557 3144 569 3184
rect 577 3144 589 3172
rect 597 3144 609 3184
rect 617 3144 629 3184
rect 679 3144 691 3184
rect 709 3144 721 3184
rect 737 3144 749 3164
rect 757 3144 769 3164
rect 811 3144 823 3184
rect 831 3144 843 3184
rect 851 3144 863 3184
rect 871 3144 883 3184
rect 891 3144 903 3184
rect 911 3144 923 3184
rect 931 3144 943 3184
rect 951 3144 963 3184
rect 971 3144 983 3184
rect 997 3144 1009 3184
rect 1017 3144 1029 3184
rect 1037 3144 1049 3184
rect 1057 3144 1069 3184
rect 1077 3144 1089 3184
rect 1097 3144 1109 3184
rect 1117 3144 1129 3184
rect 1137 3144 1149 3184
rect 1157 3144 1169 3184
rect 1211 3144 1223 3164
rect 1231 3144 1243 3164
rect 1257 3144 1269 3184
rect 1279 3144 1291 3164
rect 1309 3144 1321 3164
rect 1337 3144 1349 3164
rect 1363 3144 1375 3164
rect 1385 3144 1397 3164
rect 1415 3144 1427 3164
rect 1447 3144 1459 3164
rect 1467 3144 1479 3184
rect 1497 3144 1509 3184
rect 1517 3144 1529 3172
rect 1537 3144 1549 3184
rect 1557 3144 1569 3184
rect 1611 3144 1623 3184
rect 1631 3144 1643 3184
rect 1651 3144 1663 3172
rect 1671 3144 1683 3184
rect 1711 3144 1723 3184
rect 1731 3144 1743 3184
rect 1751 3144 1763 3172
rect 1771 3144 1783 3184
rect 1811 3144 1823 3164
rect 1831 3144 1843 3164
rect 1871 3144 1883 3184
rect 1891 3144 1903 3184
rect 1911 3144 1923 3172
rect 1931 3144 1943 3184
rect 1971 3144 1983 3184
rect 1991 3144 2003 3184
rect 2011 3144 2023 3172
rect 2031 3144 2043 3184
rect 2057 3144 2069 3184
rect 2079 3144 2091 3164
rect 2109 3144 2121 3164
rect 2137 3144 2149 3164
rect 2163 3144 2175 3164
rect 2185 3144 2197 3164
rect 2215 3144 2227 3164
rect 2247 3144 2259 3164
rect 2267 3144 2279 3184
rect 2311 3144 2323 3164
rect 2331 3144 2343 3164
rect 2371 3144 2383 3164
rect 2391 3144 2403 3164
rect 2454 3144 2466 3202
rect 2490 3144 2502 3204
rect 2520 3144 2532 3184
rect 2548 3144 2560 3184
rect 2570 3144 2582 3164
rect 2631 3144 2643 3164
rect 2651 3144 2663 3164
rect 2691 3144 2703 3184
rect 2711 3144 2723 3184
rect 2731 3144 2743 3172
rect 2751 3144 2763 3184
rect 2777 3144 2789 3164
rect 2797 3144 2809 3164
rect 2817 3144 2829 3164
rect 2857 3144 2869 3184
rect 2877 3144 2889 3172
rect 2897 3144 2909 3184
rect 2917 3144 2929 3184
rect 2959 3144 2971 3184
rect 2989 3144 3001 3184
rect 3039 3144 3051 3184
rect 3069 3144 3081 3184
rect 3138 3144 3150 3164
rect 3160 3144 3172 3184
rect 3188 3144 3200 3184
rect 3254 3144 3266 3202
rect 3290 3144 3302 3204
rect 3331 3144 3343 3184
rect 3351 3144 3363 3184
rect 3371 3144 3383 3172
rect 3391 3144 3403 3184
rect 3441 3144 3453 3184
rect 3461 3144 3473 3184
rect 3491 3144 3503 3184
rect 3519 3144 3531 3184
rect 3549 3144 3561 3184
rect 3621 3144 3633 3184
rect 3641 3144 3653 3184
rect 3671 3144 3683 3184
rect 3732 3144 3744 3184
rect 3760 3144 3772 3184
rect 3788 3144 3800 3184
rect 3839 3144 3851 3184
rect 3869 3144 3881 3184
rect 3897 3144 3909 3184
rect 3917 3144 3929 3172
rect 3937 3144 3949 3184
rect 3957 3144 3969 3184
rect 3999 3144 4011 3184
rect 4029 3144 4041 3184
rect 4101 3144 4113 3184
rect 4121 3144 4133 3184
rect 4151 3144 4163 3184
rect 4179 3144 4191 3184
rect 4209 3144 4221 3184
rect 4257 3144 4269 3184
rect 4287 3144 4299 3184
rect 4307 3144 4319 3184
rect 4360 3144 4372 3184
rect 4388 3144 4400 3184
rect 4410 3144 4422 3164
rect 4457 3144 4469 3184
rect 4477 3144 4489 3172
rect 4497 3144 4509 3184
rect 4517 3144 4529 3184
rect 4557 3144 4569 3184
rect 4577 3144 4589 3172
rect 4597 3144 4609 3184
rect 4617 3144 4629 3184
rect 4694 3144 4706 3202
rect 4730 3144 4742 3204
rect 21 3076 33 3116
rect 41 3096 53 3116
rect 73 3096 85 3116
rect 103 3096 115 3116
rect 125 3096 137 3116
rect 151 3096 163 3116
rect 179 3096 191 3116
rect 209 3096 221 3116
rect 231 3076 243 3116
rect 271 3076 283 3116
rect 291 3076 303 3116
rect 311 3088 323 3116
rect 331 3076 343 3116
rect 379 3076 391 3116
rect 409 3076 421 3116
rect 437 3076 449 3116
rect 459 3096 471 3116
rect 489 3096 501 3116
rect 517 3096 529 3116
rect 543 3096 555 3116
rect 565 3096 577 3116
rect 595 3096 607 3116
rect 627 3096 639 3116
rect 647 3076 659 3116
rect 681 3076 693 3116
rect 701 3096 713 3116
rect 733 3096 745 3116
rect 763 3096 775 3116
rect 785 3096 797 3116
rect 811 3096 823 3116
rect 839 3096 851 3116
rect 869 3096 881 3116
rect 891 3076 903 3116
rect 917 3096 929 3116
rect 937 3096 949 3116
rect 991 3096 1003 3116
rect 1011 3096 1023 3116
rect 1031 3096 1043 3116
rect 1079 3076 1091 3116
rect 1109 3076 1121 3116
rect 1137 3076 1149 3116
rect 1157 3088 1169 3116
rect 1177 3076 1189 3116
rect 1197 3076 1209 3116
rect 1240 3076 1252 3116
rect 1268 3076 1280 3116
rect 1290 3096 1302 3116
rect 1341 3076 1353 3116
rect 1361 3096 1373 3116
rect 1393 3096 1405 3116
rect 1423 3096 1435 3116
rect 1445 3096 1457 3116
rect 1471 3096 1483 3116
rect 1499 3096 1511 3116
rect 1529 3096 1541 3116
rect 1551 3076 1563 3116
rect 1591 3096 1603 3116
rect 1611 3096 1623 3116
rect 1631 3096 1643 3116
rect 1679 3076 1691 3116
rect 1709 3076 1721 3116
rect 1737 3076 1749 3116
rect 1757 3088 1769 3116
rect 1777 3076 1789 3116
rect 1797 3076 1809 3116
rect 1851 3076 1863 3116
rect 1871 3076 1883 3116
rect 1891 3088 1903 3116
rect 1911 3076 1923 3116
rect 1937 3076 1949 3116
rect 1959 3096 1971 3116
rect 1989 3096 2001 3116
rect 2017 3096 2029 3116
rect 2043 3096 2055 3116
rect 2065 3096 2077 3116
rect 2095 3096 2107 3116
rect 2127 3096 2139 3116
rect 2147 3076 2159 3116
rect 2191 3096 2203 3116
rect 2211 3096 2223 3116
rect 2231 3096 2243 3116
rect 2271 3096 2283 3116
rect 2291 3096 2303 3116
rect 2354 3058 2366 3116
rect 2390 3056 2402 3116
rect 2438 3096 2450 3116
rect 2460 3076 2472 3116
rect 2488 3076 2500 3116
rect 2554 3058 2566 3116
rect 2590 3056 2602 3116
rect 2631 3076 2643 3116
rect 2651 3076 2663 3116
rect 2671 3088 2683 3116
rect 2691 3076 2703 3116
rect 2731 3096 2743 3116
rect 2751 3096 2763 3116
rect 2771 3096 2783 3116
rect 2799 3076 2811 3116
rect 2829 3076 2841 3116
rect 2879 3076 2891 3116
rect 2909 3076 2921 3116
rect 2960 3076 2972 3116
rect 2988 3076 3000 3116
rect 3016 3076 3028 3116
rect 3079 3076 3091 3116
rect 3109 3076 3121 3116
rect 3157 3076 3169 3116
rect 3177 3088 3189 3116
rect 3197 3076 3209 3116
rect 3217 3076 3229 3116
rect 3257 3076 3269 3116
rect 3277 3076 3289 3116
rect 3317 3076 3329 3116
rect 3347 3076 3359 3116
rect 3367 3076 3379 3116
rect 3429 3076 3441 3116
rect 3449 3076 3461 3116
rect 3471 3096 3483 3116
rect 3509 3076 3521 3116
rect 3529 3076 3541 3116
rect 3551 3096 3563 3116
rect 3579 3076 3591 3116
rect 3609 3076 3621 3116
rect 3657 3076 3669 3116
rect 3677 3088 3689 3116
rect 3697 3076 3709 3116
rect 3717 3076 3729 3116
rect 3769 3076 3781 3116
rect 3789 3076 3801 3116
rect 3811 3096 3823 3116
rect 3837 3076 3849 3116
rect 3857 3088 3869 3116
rect 3877 3076 3889 3116
rect 3897 3076 3909 3116
rect 3938 3056 3950 3116
rect 3974 3058 3986 3116
rect 4037 3096 4049 3116
rect 4059 3076 4071 3116
rect 4079 3076 4091 3116
rect 4138 3096 4150 3116
rect 4160 3076 4172 3116
rect 4188 3076 4200 3116
rect 4218 3056 4230 3116
rect 4254 3058 4266 3116
rect 4338 3096 4350 3116
rect 4360 3076 4372 3116
rect 4388 3076 4400 3116
rect 4454 3058 4466 3116
rect 4490 3056 4502 3116
rect 4531 3096 4543 3116
rect 4551 3096 4563 3116
rect 4591 3076 4603 3116
rect 4611 3076 4623 3116
rect 4631 3088 4643 3116
rect 4651 3076 4663 3116
rect 4677 3076 4689 3116
rect 4697 3088 4709 3116
rect 4717 3076 4729 3116
rect 4737 3076 4749 3116
rect 21 2664 33 2704
rect 41 2664 53 2684
rect 73 2664 85 2684
rect 103 2664 115 2684
rect 125 2664 137 2684
rect 151 2664 163 2684
rect 179 2664 191 2684
rect 209 2664 221 2684
rect 231 2664 243 2704
rect 292 2664 304 2704
rect 320 2664 332 2704
rect 348 2664 360 2704
rect 379 2664 391 2704
rect 409 2664 421 2704
rect 471 2664 483 2704
rect 491 2664 503 2704
rect 511 2664 523 2692
rect 531 2664 543 2704
rect 569 2664 581 2704
rect 589 2664 601 2704
rect 611 2664 623 2684
rect 639 2664 651 2704
rect 669 2664 681 2704
rect 731 2664 743 2704
rect 751 2664 763 2704
rect 771 2664 783 2692
rect 791 2664 803 2704
rect 831 2664 843 2684
rect 851 2664 863 2684
rect 871 2664 883 2684
rect 919 2664 931 2704
rect 949 2664 961 2704
rect 977 2664 989 2684
rect 997 2664 1009 2684
rect 1059 2664 1071 2704
rect 1089 2664 1101 2704
rect 1117 2664 1129 2684
rect 1137 2664 1149 2684
rect 1157 2664 1169 2684
rect 1209 2664 1221 2704
rect 1229 2664 1241 2704
rect 1251 2664 1263 2684
rect 1281 2664 1293 2704
rect 1301 2664 1313 2684
rect 1333 2664 1345 2684
rect 1363 2664 1375 2684
rect 1385 2664 1397 2684
rect 1411 2664 1423 2684
rect 1439 2664 1451 2684
rect 1469 2664 1481 2684
rect 1491 2664 1503 2704
rect 1519 2664 1531 2704
rect 1549 2664 1561 2704
rect 1611 2664 1623 2704
rect 1631 2664 1643 2704
rect 1651 2664 1663 2692
rect 1671 2664 1683 2704
rect 1711 2664 1723 2704
rect 1731 2664 1743 2704
rect 1751 2664 1763 2692
rect 1771 2664 1783 2704
rect 1811 2664 1823 2684
rect 1831 2664 1843 2684
rect 1851 2664 1863 2684
rect 1898 2664 1910 2684
rect 1920 2664 1932 2704
rect 1948 2664 1960 2704
rect 1989 2664 2001 2704
rect 2009 2664 2021 2704
rect 2031 2664 2043 2684
rect 2094 2664 2106 2722
rect 2130 2664 2142 2724
rect 2157 2664 2169 2684
rect 2179 2664 2191 2704
rect 2199 2664 2211 2704
rect 2241 2664 2253 2704
rect 2261 2664 2273 2684
rect 2293 2664 2305 2684
rect 2323 2664 2335 2684
rect 2345 2664 2357 2684
rect 2371 2664 2383 2684
rect 2399 2664 2411 2684
rect 2429 2664 2441 2684
rect 2451 2664 2463 2704
rect 2491 2664 2503 2704
rect 2511 2664 2523 2704
rect 2531 2664 2543 2692
rect 2551 2664 2563 2704
rect 2591 2664 2603 2704
rect 2611 2664 2623 2704
rect 2631 2664 2643 2692
rect 2651 2664 2663 2704
rect 2677 2664 2689 2704
rect 2697 2664 2709 2692
rect 2717 2664 2729 2704
rect 2737 2664 2749 2704
rect 2779 2664 2791 2704
rect 2809 2664 2821 2704
rect 2859 2664 2871 2704
rect 2889 2664 2901 2704
rect 2937 2664 2949 2704
rect 2957 2664 2969 2692
rect 2977 2664 2989 2704
rect 2997 2664 3009 2704
rect 3037 2664 3049 2704
rect 3057 2664 3069 2692
rect 3077 2664 3089 2704
rect 3097 2664 3109 2704
rect 3139 2664 3151 2704
rect 3169 2664 3181 2704
rect 3231 2664 3243 2704
rect 3251 2664 3263 2704
rect 3271 2664 3283 2692
rect 3291 2664 3303 2704
rect 3339 2664 3351 2704
rect 3369 2664 3381 2704
rect 3398 2664 3410 2724
rect 3434 2664 3446 2722
rect 3511 2664 3523 2704
rect 3531 2664 3543 2704
rect 3551 2664 3563 2692
rect 3571 2664 3583 2704
rect 3597 2664 3609 2704
rect 3617 2664 3629 2692
rect 3637 2664 3649 2704
rect 3657 2664 3669 2704
rect 3719 2664 3731 2704
rect 3749 2664 3761 2704
rect 3791 2664 3803 2704
rect 3811 2664 3823 2704
rect 3831 2664 3843 2692
rect 3851 2664 3863 2704
rect 3878 2664 3890 2724
rect 3914 2664 3926 2722
rect 3977 2664 3989 2684
rect 3997 2664 4009 2684
rect 4072 2664 4084 2704
rect 4100 2664 4112 2704
rect 4128 2664 4140 2704
rect 4158 2664 4170 2724
rect 4194 2664 4206 2722
rect 4257 2664 4269 2704
rect 4277 2664 4289 2692
rect 4297 2664 4309 2704
rect 4317 2664 4329 2704
rect 4357 2664 4369 2704
rect 4387 2664 4399 2704
rect 4407 2664 4419 2704
rect 4460 2664 4472 2704
rect 4488 2664 4500 2704
rect 4516 2664 4528 2704
rect 4577 2664 4589 2684
rect 4597 2664 4609 2684
rect 4640 2664 4652 2704
rect 4668 2664 4680 2704
rect 4690 2664 4702 2684
rect 21 2596 33 2636
rect 41 2616 53 2636
rect 73 2616 85 2636
rect 103 2616 115 2636
rect 125 2616 137 2636
rect 151 2616 163 2636
rect 179 2616 191 2636
rect 209 2616 221 2636
rect 231 2596 243 2636
rect 271 2596 283 2636
rect 291 2596 303 2636
rect 311 2608 323 2636
rect 331 2596 343 2636
rect 357 2616 369 2636
rect 379 2596 391 2636
rect 399 2596 411 2636
rect 439 2596 451 2636
rect 469 2596 481 2636
rect 531 2596 543 2636
rect 551 2596 563 2636
rect 571 2608 583 2636
rect 591 2596 603 2636
rect 617 2616 629 2636
rect 639 2596 651 2636
rect 659 2596 671 2636
rect 711 2596 723 2636
rect 731 2596 743 2636
rect 751 2608 763 2636
rect 771 2596 783 2636
rect 797 2616 809 2636
rect 817 2616 829 2636
rect 837 2616 849 2636
rect 881 2596 893 2636
rect 901 2616 913 2636
rect 933 2616 945 2636
rect 963 2616 975 2636
rect 985 2616 997 2636
rect 1011 2616 1023 2636
rect 1039 2616 1051 2636
rect 1069 2616 1081 2636
rect 1091 2596 1103 2636
rect 1117 2616 1129 2636
rect 1137 2616 1149 2636
rect 1177 2596 1189 2636
rect 1197 2608 1209 2636
rect 1217 2596 1229 2636
rect 1237 2596 1249 2636
rect 1277 2616 1289 2636
rect 1297 2616 1309 2636
rect 1339 2596 1351 2636
rect 1369 2596 1381 2636
rect 1417 2596 1429 2636
rect 1439 2616 1451 2636
rect 1469 2616 1481 2636
rect 1497 2616 1509 2636
rect 1523 2616 1535 2636
rect 1545 2616 1557 2636
rect 1575 2616 1587 2636
rect 1607 2616 1619 2636
rect 1627 2596 1639 2636
rect 1657 2596 1669 2636
rect 1677 2608 1689 2636
rect 1697 2596 1709 2636
rect 1717 2596 1729 2636
rect 1757 2596 1769 2636
rect 1779 2616 1791 2636
rect 1809 2616 1821 2636
rect 1837 2616 1849 2636
rect 1863 2616 1875 2636
rect 1885 2616 1897 2636
rect 1915 2616 1927 2636
rect 1947 2616 1959 2636
rect 1967 2596 1979 2636
rect 1997 2596 2009 2636
rect 2017 2596 2029 2636
rect 2037 2596 2049 2636
rect 2057 2596 2069 2636
rect 2077 2596 2089 2636
rect 2097 2596 2109 2636
rect 2117 2596 2129 2636
rect 2137 2596 2149 2636
rect 2157 2596 2169 2636
rect 2201 2596 2213 2636
rect 2221 2616 2233 2636
rect 2253 2616 2265 2636
rect 2283 2616 2295 2636
rect 2305 2616 2317 2636
rect 2331 2616 2343 2636
rect 2359 2616 2371 2636
rect 2389 2616 2401 2636
rect 2411 2596 2423 2636
rect 2459 2596 2471 2636
rect 2489 2596 2501 2636
rect 2517 2616 2529 2636
rect 2537 2616 2549 2636
rect 2591 2596 2603 2636
rect 2611 2596 2623 2636
rect 2631 2608 2643 2636
rect 2651 2596 2663 2636
rect 2677 2616 2689 2636
rect 2697 2616 2709 2636
rect 2759 2596 2771 2636
rect 2789 2596 2801 2636
rect 2831 2596 2843 2636
rect 2851 2596 2863 2636
rect 2871 2608 2883 2636
rect 2891 2596 2903 2636
rect 2917 2596 2929 2636
rect 2947 2596 2959 2636
rect 2967 2596 2979 2636
rect 3017 2596 3029 2636
rect 3037 2608 3049 2636
rect 3057 2596 3069 2636
rect 3077 2596 3089 2636
rect 3139 2596 3151 2636
rect 3169 2596 3181 2636
rect 3197 2596 3209 2636
rect 3227 2596 3239 2636
rect 3247 2596 3259 2636
rect 3334 2578 3346 2636
rect 3370 2576 3382 2636
rect 3397 2616 3409 2636
rect 3417 2616 3429 2636
rect 3459 2596 3471 2636
rect 3489 2596 3501 2636
rect 3537 2596 3549 2636
rect 3567 2596 3579 2636
rect 3587 2596 3599 2636
rect 3637 2616 3649 2636
rect 3659 2596 3671 2636
rect 3679 2596 3691 2636
rect 3717 2616 3729 2636
rect 3737 2616 3749 2636
rect 3801 2596 3813 2636
rect 3821 2596 3833 2636
rect 3851 2596 3863 2636
rect 3912 2596 3924 2636
rect 3940 2596 3952 2636
rect 3968 2596 3980 2636
rect 4019 2596 4031 2636
rect 4049 2596 4061 2636
rect 4099 2596 4111 2636
rect 4129 2596 4141 2636
rect 4157 2596 4169 2636
rect 4177 2608 4189 2636
rect 4197 2596 4209 2636
rect 4217 2596 4229 2636
rect 4259 2596 4271 2636
rect 4289 2596 4301 2636
rect 4374 2578 4386 2636
rect 4410 2576 4422 2636
rect 4474 2578 4486 2636
rect 4510 2576 4522 2636
rect 4540 2596 4552 2636
rect 4568 2596 4580 2636
rect 4590 2616 4602 2636
rect 4674 2578 4686 2636
rect 4710 2576 4722 2636
rect 21 2184 33 2224
rect 41 2184 53 2204
rect 73 2184 85 2204
rect 103 2184 115 2204
rect 125 2184 137 2204
rect 151 2184 163 2204
rect 179 2184 191 2204
rect 209 2184 221 2204
rect 231 2184 243 2224
rect 257 2184 269 2224
rect 277 2184 289 2212
rect 297 2184 309 2224
rect 317 2184 329 2224
rect 360 2184 372 2224
rect 388 2184 400 2224
rect 416 2184 428 2224
rect 477 2184 489 2204
rect 499 2184 511 2224
rect 519 2184 531 2224
rect 559 2184 571 2224
rect 589 2184 601 2224
rect 651 2184 663 2204
rect 671 2184 683 2204
rect 697 2184 709 2204
rect 717 2184 729 2204
rect 737 2184 749 2204
rect 798 2184 810 2204
rect 820 2184 832 2224
rect 848 2184 860 2224
rect 877 2184 889 2204
rect 897 2184 909 2204
rect 917 2184 929 2204
rect 957 2184 969 2204
rect 977 2184 989 2204
rect 997 2184 1009 2204
rect 1037 2184 1049 2204
rect 1057 2184 1069 2204
rect 1097 2184 1109 2224
rect 1119 2184 1131 2204
rect 1149 2184 1161 2204
rect 1177 2184 1189 2204
rect 1203 2184 1215 2204
rect 1225 2184 1237 2204
rect 1255 2184 1267 2204
rect 1287 2184 1299 2204
rect 1307 2184 1319 2224
rect 1337 2184 1349 2224
rect 1357 2184 1369 2212
rect 1377 2184 1389 2224
rect 1397 2184 1409 2224
rect 1437 2184 1449 2224
rect 1459 2184 1471 2204
rect 1489 2184 1501 2204
rect 1517 2184 1529 2204
rect 1543 2184 1555 2204
rect 1565 2184 1577 2204
rect 1595 2184 1607 2204
rect 1627 2184 1639 2204
rect 1647 2184 1659 2224
rect 1691 2184 1703 2204
rect 1711 2184 1723 2204
rect 1731 2184 1743 2204
rect 1778 2184 1790 2204
rect 1800 2184 1812 2224
rect 1828 2184 1840 2224
rect 1857 2184 1869 2224
rect 1877 2184 1889 2224
rect 1931 2184 1943 2204
rect 1951 2184 1963 2204
rect 1971 2184 1983 2204
rect 1997 2184 2009 2224
rect 2017 2184 2029 2224
rect 2037 2184 2049 2224
rect 2057 2184 2069 2224
rect 2077 2184 2089 2224
rect 2097 2184 2109 2224
rect 2117 2184 2129 2224
rect 2137 2184 2149 2224
rect 2157 2184 2169 2224
rect 2197 2184 2209 2224
rect 2217 2184 2229 2212
rect 2237 2184 2249 2224
rect 2257 2184 2269 2224
rect 2301 2184 2313 2224
rect 2321 2184 2333 2204
rect 2353 2184 2365 2204
rect 2383 2184 2395 2204
rect 2405 2184 2417 2204
rect 2431 2184 2443 2204
rect 2459 2184 2471 2204
rect 2489 2184 2501 2204
rect 2511 2184 2523 2224
rect 2559 2184 2571 2224
rect 2589 2184 2601 2224
rect 2619 2184 2631 2224
rect 2649 2184 2661 2224
rect 2699 2184 2711 2224
rect 2729 2184 2741 2224
rect 2791 2184 2803 2224
rect 2811 2184 2823 2224
rect 2831 2184 2843 2212
rect 2851 2184 2863 2224
rect 2891 2184 2903 2224
rect 2911 2184 2923 2224
rect 2931 2184 2943 2212
rect 2951 2184 2963 2224
rect 2981 2184 2993 2224
rect 3001 2184 3013 2204
rect 3033 2184 3045 2204
rect 3063 2184 3075 2204
rect 3085 2184 3097 2204
rect 3111 2184 3123 2204
rect 3139 2184 3151 2204
rect 3169 2184 3181 2204
rect 3191 2184 3203 2224
rect 3217 2184 3229 2224
rect 3237 2184 3249 2212
rect 3257 2184 3269 2224
rect 3277 2184 3289 2224
rect 3319 2184 3331 2224
rect 3349 2184 3361 2224
rect 3399 2184 3411 2224
rect 3429 2184 3441 2224
rect 3499 2184 3511 2224
rect 3529 2184 3541 2224
rect 3571 2184 3583 2224
rect 3591 2184 3603 2224
rect 3631 2184 3643 2224
rect 3651 2184 3663 2224
rect 3691 2184 3703 2204
rect 3711 2184 3723 2204
rect 3737 2184 3749 2224
rect 3757 2184 3769 2212
rect 3777 2184 3789 2224
rect 3797 2184 3809 2224
rect 3849 2184 3861 2224
rect 3869 2184 3881 2224
rect 3891 2184 3903 2204
rect 3917 2184 3929 2224
rect 3937 2184 3949 2224
rect 3977 2184 3989 2224
rect 4007 2184 4019 2224
rect 4027 2184 4039 2224
rect 4091 2184 4103 2224
rect 4111 2184 4123 2224
rect 4131 2184 4143 2212
rect 4151 2184 4163 2224
rect 4214 2184 4226 2242
rect 4250 2184 4262 2244
rect 4280 2184 4292 2224
rect 4308 2184 4320 2224
rect 4330 2184 4342 2204
rect 4391 2184 4403 2224
rect 4411 2184 4423 2224
rect 4431 2184 4443 2212
rect 4451 2184 4463 2224
rect 4477 2184 4489 2224
rect 4497 2184 4509 2212
rect 4517 2184 4529 2224
rect 4537 2184 4549 2224
rect 4591 2184 4603 2224
rect 4611 2184 4623 2224
rect 4631 2184 4643 2212
rect 4651 2184 4663 2224
rect 4680 2184 4692 2224
rect 4708 2184 4720 2224
rect 4730 2184 4742 2204
rect 17 2116 29 2156
rect 37 2116 49 2156
rect 57 2116 69 2156
rect 77 2116 89 2156
rect 97 2116 109 2156
rect 117 2116 129 2156
rect 137 2116 149 2156
rect 157 2116 169 2156
rect 177 2116 189 2156
rect 239 2116 251 2156
rect 269 2116 281 2156
rect 311 2116 323 2156
rect 331 2116 343 2156
rect 351 2128 363 2156
rect 371 2116 383 2156
rect 400 2116 412 2156
rect 428 2116 440 2156
rect 456 2116 468 2156
rect 521 2116 533 2156
rect 541 2136 553 2156
rect 573 2136 585 2156
rect 603 2136 615 2156
rect 625 2136 637 2156
rect 651 2136 663 2156
rect 679 2136 691 2156
rect 709 2136 721 2156
rect 731 2116 743 2156
rect 779 2116 791 2156
rect 809 2116 821 2156
rect 851 2116 863 2156
rect 871 2136 883 2156
rect 891 2136 903 2156
rect 911 2136 923 2156
rect 939 2116 951 2156
rect 969 2116 981 2156
rect 1017 2136 1029 2156
rect 1037 2136 1049 2156
rect 1057 2136 1069 2156
rect 1097 2116 1109 2156
rect 1117 2128 1129 2156
rect 1137 2116 1149 2156
rect 1157 2116 1169 2156
rect 1199 2116 1211 2156
rect 1229 2116 1241 2156
rect 1277 2136 1289 2156
rect 1297 2136 1309 2156
rect 1317 2136 1329 2156
rect 1357 2116 1369 2156
rect 1379 2136 1391 2156
rect 1409 2136 1421 2156
rect 1437 2136 1449 2156
rect 1463 2136 1475 2156
rect 1485 2136 1497 2156
rect 1515 2136 1527 2156
rect 1547 2136 1559 2156
rect 1567 2116 1579 2156
rect 1618 2136 1630 2156
rect 1640 2116 1652 2156
rect 1668 2116 1680 2156
rect 1709 2116 1721 2156
rect 1729 2116 1741 2156
rect 1751 2136 1763 2156
rect 1777 2116 1789 2156
rect 1799 2136 1811 2156
rect 1829 2136 1841 2156
rect 1857 2136 1869 2156
rect 1883 2136 1895 2156
rect 1905 2136 1917 2156
rect 1935 2136 1947 2156
rect 1967 2136 1979 2156
rect 1987 2116 1999 2156
rect 2031 2136 2043 2156
rect 2051 2136 2063 2156
rect 2099 2116 2111 2156
rect 2129 2116 2141 2156
rect 2157 2136 2169 2156
rect 2179 2116 2191 2156
rect 2199 2116 2211 2156
rect 2239 2116 2251 2156
rect 2269 2116 2281 2156
rect 2331 2116 2343 2156
rect 2351 2116 2363 2156
rect 2371 2128 2383 2156
rect 2391 2116 2403 2156
rect 2439 2116 2451 2156
rect 2469 2116 2481 2156
rect 2519 2116 2531 2156
rect 2549 2116 2561 2156
rect 2591 2116 2603 2156
rect 2611 2116 2623 2156
rect 2631 2128 2643 2156
rect 2651 2116 2663 2156
rect 2691 2116 2703 2156
rect 2711 2116 2723 2156
rect 2731 2128 2743 2156
rect 2751 2116 2763 2156
rect 2781 2116 2793 2156
rect 2801 2136 2813 2156
rect 2833 2136 2845 2156
rect 2863 2136 2875 2156
rect 2885 2136 2897 2156
rect 2911 2136 2923 2156
rect 2939 2136 2951 2156
rect 2969 2136 2981 2156
rect 2991 2116 3003 2156
rect 3017 2116 3029 2156
rect 3047 2116 3059 2156
rect 3067 2116 3079 2156
rect 3131 2116 3143 2156
rect 3151 2116 3163 2156
rect 3171 2128 3183 2156
rect 3191 2116 3203 2156
rect 3231 2116 3243 2156
rect 3251 2116 3263 2156
rect 3271 2128 3283 2156
rect 3291 2116 3303 2156
rect 3319 2116 3331 2156
rect 3349 2116 3361 2156
rect 3411 2116 3423 2156
rect 3431 2116 3443 2156
rect 3451 2128 3463 2156
rect 3471 2116 3483 2156
rect 3498 2096 3510 2156
rect 3534 2098 3546 2156
rect 3597 2136 3609 2156
rect 3617 2136 3629 2156
rect 3658 2096 3670 2156
rect 3694 2098 3706 2156
rect 3759 2116 3771 2156
rect 3789 2116 3801 2156
rect 3837 2136 3849 2156
rect 3859 2116 3871 2156
rect 3879 2116 3891 2156
rect 3917 2116 3929 2156
rect 3937 2128 3949 2156
rect 3957 2116 3969 2156
rect 3977 2116 3989 2156
rect 4039 2116 4051 2156
rect 4069 2116 4081 2156
rect 4119 2116 4131 2156
rect 4149 2116 4161 2156
rect 4199 2116 4211 2156
rect 4229 2116 4241 2156
rect 4257 2116 4269 2156
rect 4287 2116 4299 2156
rect 4307 2116 4319 2156
rect 4360 2116 4372 2156
rect 4388 2116 4400 2156
rect 4410 2136 4422 2156
rect 4478 2136 4490 2156
rect 4500 2116 4512 2156
rect 4528 2116 4540 2156
rect 4558 2096 4570 2156
rect 4594 2098 4606 2156
rect 4658 2096 4670 2156
rect 4694 2098 4706 2156
rect 21 1704 33 1744
rect 41 1704 53 1724
rect 73 1704 85 1724
rect 103 1704 115 1724
rect 125 1704 137 1724
rect 151 1704 163 1724
rect 179 1704 191 1724
rect 209 1704 221 1724
rect 231 1704 243 1744
rect 257 1704 269 1744
rect 277 1704 289 1732
rect 297 1704 309 1744
rect 317 1704 329 1744
rect 371 1704 383 1744
rect 391 1704 403 1744
rect 411 1704 423 1732
rect 431 1704 443 1744
rect 471 1704 483 1744
rect 491 1704 503 1744
rect 511 1704 523 1732
rect 531 1704 543 1744
rect 571 1704 583 1744
rect 591 1704 603 1744
rect 611 1704 623 1732
rect 631 1704 643 1744
rect 657 1704 669 1724
rect 677 1704 689 1724
rect 717 1704 729 1724
rect 737 1704 749 1724
rect 791 1704 803 1724
rect 811 1704 823 1724
rect 831 1704 843 1724
rect 858 1704 870 1764
rect 894 1704 906 1762
rect 961 1704 973 1744
rect 981 1704 993 1724
rect 1013 1704 1025 1724
rect 1043 1704 1055 1724
rect 1065 1704 1077 1724
rect 1091 1704 1103 1724
rect 1119 1704 1131 1724
rect 1149 1704 1161 1724
rect 1171 1704 1183 1744
rect 1199 1704 1211 1744
rect 1229 1704 1241 1744
rect 1291 1704 1303 1744
rect 1311 1704 1323 1744
rect 1331 1704 1343 1732
rect 1351 1704 1363 1744
rect 1391 1704 1403 1744
rect 1411 1704 1423 1744
rect 1431 1704 1443 1744
rect 1451 1704 1463 1744
rect 1471 1704 1483 1744
rect 1491 1704 1503 1744
rect 1511 1704 1523 1744
rect 1531 1704 1543 1744
rect 1551 1704 1563 1744
rect 1581 1704 1593 1744
rect 1601 1704 1613 1724
rect 1633 1704 1645 1724
rect 1663 1704 1675 1724
rect 1685 1704 1697 1724
rect 1711 1704 1723 1724
rect 1739 1704 1751 1724
rect 1769 1704 1781 1724
rect 1791 1704 1803 1744
rect 1838 1704 1850 1724
rect 1860 1704 1872 1744
rect 1888 1704 1900 1744
rect 1917 1704 1929 1724
rect 1937 1704 1949 1724
rect 1957 1704 1969 1724
rect 2018 1704 2030 1724
rect 2040 1704 2052 1744
rect 2068 1704 2080 1744
rect 2111 1704 2123 1724
rect 2131 1704 2143 1724
rect 2151 1704 2163 1724
rect 2180 1704 2192 1744
rect 2208 1704 2220 1744
rect 2230 1704 2242 1724
rect 2277 1704 2289 1744
rect 2299 1704 2311 1724
rect 2329 1704 2341 1724
rect 2357 1704 2369 1724
rect 2383 1704 2395 1724
rect 2405 1704 2417 1724
rect 2435 1704 2447 1724
rect 2467 1704 2479 1724
rect 2487 1704 2499 1744
rect 2521 1704 2533 1744
rect 2541 1704 2553 1724
rect 2573 1704 2585 1724
rect 2603 1704 2615 1724
rect 2625 1704 2637 1724
rect 2651 1704 2663 1724
rect 2679 1704 2691 1724
rect 2709 1704 2721 1724
rect 2731 1704 2743 1744
rect 2761 1704 2773 1744
rect 2781 1704 2793 1724
rect 2813 1704 2825 1724
rect 2843 1704 2855 1724
rect 2865 1704 2877 1724
rect 2891 1704 2903 1724
rect 2919 1704 2931 1724
rect 2949 1704 2961 1724
rect 2971 1704 2983 1744
rect 3011 1704 3023 1744
rect 3031 1704 3043 1744
rect 3079 1704 3091 1744
rect 3109 1704 3121 1744
rect 3151 1704 3163 1744
rect 3171 1704 3183 1744
rect 3200 1704 3212 1744
rect 3228 1704 3240 1744
rect 3250 1704 3262 1724
rect 3297 1704 3309 1724
rect 3317 1704 3329 1724
rect 3337 1704 3349 1724
rect 3401 1704 3413 1744
rect 3421 1704 3433 1744
rect 3451 1704 3463 1744
rect 3477 1704 3489 1744
rect 3497 1704 3509 1744
rect 3572 1704 3584 1744
rect 3600 1704 3612 1744
rect 3628 1704 3640 1744
rect 3671 1704 3683 1744
rect 3691 1704 3703 1744
rect 3731 1704 3743 1724
rect 3751 1704 3763 1724
rect 3771 1704 3783 1724
rect 3797 1704 3809 1724
rect 3819 1704 3831 1744
rect 3839 1704 3851 1744
rect 3877 1704 3889 1744
rect 3907 1704 3919 1744
rect 3927 1704 3939 1744
rect 4012 1704 4024 1744
rect 4040 1704 4052 1744
rect 4068 1704 4080 1744
rect 4100 1704 4112 1744
rect 4128 1704 4140 1744
rect 4156 1704 4168 1744
rect 4219 1704 4231 1744
rect 4249 1704 4261 1744
rect 4297 1704 4309 1744
rect 4327 1704 4339 1744
rect 4347 1704 4359 1744
rect 4400 1704 4412 1744
rect 4428 1704 4440 1744
rect 4456 1704 4468 1744
rect 4531 1704 4543 1724
rect 4551 1704 4563 1724
rect 4577 1704 4589 1744
rect 4597 1704 4609 1732
rect 4617 1704 4629 1744
rect 4637 1704 4649 1744
rect 4677 1704 4689 1724
rect 4697 1704 4709 1724
rect 17 1636 29 1676
rect 37 1636 49 1676
rect 57 1636 69 1676
rect 77 1636 89 1676
rect 97 1636 109 1676
rect 117 1636 129 1676
rect 137 1636 149 1676
rect 157 1636 169 1676
rect 177 1636 189 1676
rect 231 1656 243 1676
rect 251 1656 263 1676
rect 271 1656 283 1676
rect 309 1636 321 1676
rect 329 1636 341 1676
rect 351 1656 363 1676
rect 381 1636 393 1676
rect 401 1656 413 1676
rect 433 1656 445 1676
rect 463 1656 475 1676
rect 485 1656 497 1676
rect 511 1656 523 1676
rect 539 1656 551 1676
rect 569 1656 581 1676
rect 591 1636 603 1676
rect 621 1636 633 1676
rect 641 1656 653 1676
rect 673 1656 685 1676
rect 703 1656 715 1676
rect 725 1656 737 1676
rect 751 1656 763 1676
rect 779 1656 791 1676
rect 809 1656 821 1676
rect 831 1636 843 1676
rect 857 1636 869 1676
rect 879 1656 891 1676
rect 909 1656 921 1676
rect 937 1656 949 1676
rect 963 1656 975 1676
rect 985 1656 997 1676
rect 1015 1656 1027 1676
rect 1047 1656 1059 1676
rect 1067 1636 1079 1676
rect 1119 1636 1131 1676
rect 1149 1636 1161 1676
rect 1191 1636 1203 1676
rect 1211 1636 1223 1676
rect 1231 1648 1243 1676
rect 1251 1636 1263 1676
rect 1277 1636 1289 1676
rect 1299 1656 1311 1676
rect 1329 1656 1341 1676
rect 1357 1656 1369 1676
rect 1383 1656 1395 1676
rect 1405 1656 1417 1676
rect 1435 1656 1447 1676
rect 1467 1656 1479 1676
rect 1487 1636 1499 1676
rect 1521 1636 1533 1676
rect 1541 1656 1553 1676
rect 1573 1656 1585 1676
rect 1603 1656 1615 1676
rect 1625 1656 1637 1676
rect 1651 1656 1663 1676
rect 1679 1656 1691 1676
rect 1709 1656 1721 1676
rect 1731 1636 1743 1676
rect 1778 1656 1790 1676
rect 1800 1636 1812 1676
rect 1828 1636 1840 1676
rect 1857 1656 1869 1676
rect 1877 1656 1889 1676
rect 1897 1656 1909 1676
rect 1941 1636 1953 1676
rect 1961 1656 1973 1676
rect 1993 1656 2005 1676
rect 2023 1656 2035 1676
rect 2045 1656 2057 1676
rect 2071 1656 2083 1676
rect 2099 1656 2111 1676
rect 2129 1656 2141 1676
rect 2151 1636 2163 1676
rect 2191 1656 2203 1676
rect 2211 1656 2223 1676
rect 2231 1656 2243 1676
rect 2279 1636 2291 1676
rect 2309 1636 2321 1676
rect 2337 1636 2349 1676
rect 2357 1648 2369 1676
rect 2377 1636 2389 1676
rect 2397 1636 2409 1676
rect 2437 1636 2449 1676
rect 2459 1656 2471 1676
rect 2489 1656 2501 1676
rect 2517 1656 2529 1676
rect 2543 1656 2555 1676
rect 2565 1656 2577 1676
rect 2595 1656 2607 1676
rect 2627 1656 2639 1676
rect 2647 1636 2659 1676
rect 2681 1636 2693 1676
rect 2701 1656 2713 1676
rect 2733 1656 2745 1676
rect 2763 1656 2775 1676
rect 2785 1656 2797 1676
rect 2811 1656 2823 1676
rect 2839 1656 2851 1676
rect 2869 1656 2881 1676
rect 2891 1636 2903 1676
rect 2917 1636 2929 1676
rect 2937 1636 2949 1676
rect 2979 1636 2991 1676
rect 3009 1636 3021 1676
rect 3079 1636 3091 1676
rect 3109 1636 3121 1676
rect 3137 1636 3149 1676
rect 3157 1648 3169 1676
rect 3177 1636 3189 1676
rect 3197 1636 3209 1676
rect 3239 1636 3251 1676
rect 3269 1636 3281 1676
rect 3339 1636 3351 1676
rect 3369 1636 3381 1676
rect 3411 1636 3423 1676
rect 3431 1636 3443 1676
rect 3451 1648 3463 1676
rect 3471 1636 3483 1676
rect 3498 1616 3510 1676
rect 3534 1618 3546 1676
rect 3611 1636 3623 1676
rect 3631 1636 3643 1664
rect 3651 1636 3663 1676
rect 3671 1646 3683 1676
rect 3691 1636 3703 1676
rect 3717 1656 3729 1676
rect 3737 1656 3749 1676
rect 3778 1616 3790 1676
rect 3814 1618 3826 1676
rect 3880 1636 3892 1676
rect 3908 1636 3920 1676
rect 3930 1656 3942 1676
rect 3977 1636 3989 1676
rect 3997 1648 4009 1676
rect 4017 1636 4029 1676
rect 4037 1636 4049 1676
rect 4099 1636 4111 1676
rect 4129 1636 4141 1676
rect 4160 1636 4172 1676
rect 4188 1636 4200 1676
rect 4210 1656 4222 1676
rect 4257 1636 4269 1676
rect 4277 1648 4289 1676
rect 4297 1636 4309 1676
rect 4317 1636 4329 1676
rect 4357 1656 4369 1676
rect 4377 1656 4389 1676
rect 4417 1656 4429 1676
rect 4437 1656 4449 1676
rect 4457 1656 4469 1676
rect 4499 1636 4511 1676
rect 4529 1636 4541 1676
rect 4579 1636 4591 1676
rect 4609 1636 4621 1676
rect 4659 1636 4671 1676
rect 4689 1636 4701 1676
rect 17 1224 29 1264
rect 39 1224 51 1244
rect 69 1224 81 1244
rect 97 1224 109 1244
rect 123 1224 135 1244
rect 145 1224 157 1244
rect 175 1224 187 1244
rect 207 1224 219 1244
rect 227 1224 239 1264
rect 261 1224 273 1264
rect 281 1224 293 1244
rect 313 1224 325 1244
rect 343 1224 355 1244
rect 365 1224 377 1244
rect 391 1224 403 1244
rect 419 1224 431 1244
rect 449 1224 461 1244
rect 471 1224 483 1264
rect 499 1224 511 1264
rect 529 1224 541 1264
rect 591 1224 603 1264
rect 611 1224 623 1264
rect 631 1224 643 1252
rect 651 1224 663 1264
rect 691 1224 703 1264
rect 711 1224 723 1264
rect 731 1224 743 1252
rect 751 1224 763 1264
rect 789 1224 801 1264
rect 809 1224 821 1264
rect 831 1224 843 1244
rect 859 1224 871 1264
rect 889 1224 901 1264
rect 951 1224 963 1264
rect 971 1224 983 1264
rect 991 1224 1003 1252
rect 1011 1224 1023 1264
rect 1051 1224 1063 1244
rect 1071 1224 1083 1244
rect 1097 1224 1109 1264
rect 1117 1224 1129 1264
rect 1137 1224 1149 1264
rect 1157 1224 1169 1264
rect 1177 1224 1189 1264
rect 1239 1224 1251 1264
rect 1269 1224 1281 1264
rect 1311 1224 1323 1264
rect 1331 1224 1343 1264
rect 1351 1224 1363 1252
rect 1371 1224 1383 1264
rect 1419 1224 1431 1264
rect 1449 1224 1461 1264
rect 1491 1224 1503 1264
rect 1511 1224 1523 1264
rect 1531 1224 1543 1252
rect 1551 1224 1563 1264
rect 1577 1224 1589 1244
rect 1599 1224 1611 1264
rect 1619 1224 1631 1264
rect 1659 1224 1671 1264
rect 1689 1224 1701 1264
rect 1751 1224 1763 1264
rect 1771 1224 1783 1264
rect 1791 1224 1803 1252
rect 1811 1224 1823 1264
rect 1837 1224 1849 1264
rect 1859 1224 1871 1244
rect 1889 1224 1901 1244
rect 1917 1224 1929 1244
rect 1943 1224 1955 1244
rect 1965 1224 1977 1244
rect 1995 1224 2007 1244
rect 2027 1224 2039 1244
rect 2047 1224 2059 1264
rect 2077 1224 2089 1244
rect 2097 1224 2109 1244
rect 2137 1224 2149 1264
rect 2157 1224 2169 1252
rect 2177 1224 2189 1264
rect 2197 1224 2209 1264
rect 2259 1224 2271 1264
rect 2289 1224 2301 1264
rect 2331 1224 2343 1244
rect 2351 1224 2363 1244
rect 2371 1224 2383 1244
rect 2411 1224 2423 1244
rect 2431 1224 2443 1244
rect 2457 1224 2469 1244
rect 2477 1224 2489 1244
rect 2497 1224 2509 1244
rect 2537 1224 2549 1264
rect 2559 1224 2571 1244
rect 2589 1224 2601 1244
rect 2617 1224 2629 1244
rect 2643 1224 2655 1244
rect 2665 1224 2677 1244
rect 2695 1224 2707 1244
rect 2727 1224 2739 1244
rect 2747 1224 2759 1264
rect 2777 1224 2789 1244
rect 2797 1224 2809 1244
rect 2817 1224 2829 1244
rect 2871 1224 2883 1264
rect 2891 1224 2903 1264
rect 2917 1224 2929 1264
rect 2937 1224 2949 1252
rect 2957 1224 2969 1264
rect 2977 1224 2989 1264
rect 3017 1224 3029 1264
rect 3037 1224 3049 1252
rect 3057 1224 3069 1264
rect 3077 1224 3089 1264
rect 3117 1224 3129 1264
rect 3137 1224 3149 1252
rect 3157 1224 3169 1264
rect 3177 1224 3189 1264
rect 3217 1224 3229 1264
rect 3247 1224 3259 1264
rect 3267 1224 3279 1264
rect 3331 1224 3343 1244
rect 3351 1224 3363 1244
rect 3371 1224 3383 1244
rect 3398 1224 3410 1284
rect 3434 1224 3446 1282
rect 3511 1224 3523 1264
rect 3531 1224 3543 1264
rect 3551 1224 3563 1252
rect 3571 1224 3583 1264
rect 3597 1224 3609 1264
rect 3617 1224 3629 1252
rect 3637 1224 3649 1264
rect 3657 1224 3669 1264
rect 3719 1224 3731 1264
rect 3749 1224 3761 1264
rect 3799 1224 3811 1264
rect 3829 1224 3841 1264
rect 3857 1224 3869 1264
rect 3887 1224 3899 1264
rect 3907 1224 3919 1264
rect 3971 1224 3983 1264
rect 3991 1224 4003 1264
rect 4011 1224 4023 1252
rect 4031 1224 4043 1264
rect 4057 1224 4069 1244
rect 4077 1224 4089 1244
rect 4139 1224 4151 1264
rect 4169 1224 4181 1264
rect 4219 1224 4231 1264
rect 4249 1224 4261 1264
rect 4291 1224 4303 1244
rect 4311 1224 4323 1244
rect 4331 1224 4343 1244
rect 4371 1224 4383 1264
rect 4391 1224 4403 1264
rect 4411 1224 4423 1252
rect 4431 1224 4443 1264
rect 4457 1224 4469 1264
rect 4477 1224 4489 1252
rect 4497 1224 4509 1264
rect 4517 1224 4529 1264
rect 4578 1224 4590 1244
rect 4600 1224 4612 1264
rect 4628 1224 4640 1264
rect 4659 1224 4671 1264
rect 4689 1224 4701 1264
rect 17 1176 29 1196
rect 37 1176 49 1196
rect 99 1156 111 1196
rect 129 1156 141 1196
rect 171 1156 183 1196
rect 191 1156 203 1196
rect 211 1168 223 1196
rect 231 1156 243 1196
rect 260 1156 272 1196
rect 288 1156 300 1196
rect 316 1156 328 1196
rect 398 1176 410 1196
rect 420 1156 432 1196
rect 448 1156 460 1196
rect 491 1156 503 1196
rect 511 1176 523 1196
rect 531 1176 543 1196
rect 551 1176 563 1196
rect 577 1176 589 1196
rect 597 1176 609 1196
rect 617 1176 629 1196
rect 681 1156 693 1196
rect 701 1156 713 1196
rect 731 1156 743 1196
rect 769 1156 781 1196
rect 789 1156 801 1196
rect 811 1176 823 1196
rect 851 1176 863 1196
rect 871 1176 883 1196
rect 891 1176 903 1196
rect 931 1176 943 1196
rect 951 1176 963 1196
rect 991 1176 1003 1196
rect 1011 1176 1023 1196
rect 1037 1176 1049 1196
rect 1057 1176 1069 1196
rect 1077 1176 1089 1196
rect 1117 1176 1129 1196
rect 1137 1176 1149 1196
rect 1191 1176 1203 1196
rect 1211 1176 1223 1196
rect 1231 1176 1243 1196
rect 1260 1156 1272 1196
rect 1288 1156 1300 1196
rect 1310 1176 1322 1196
rect 1361 1156 1373 1196
rect 1381 1176 1393 1196
rect 1413 1176 1425 1196
rect 1443 1176 1455 1196
rect 1465 1176 1477 1196
rect 1491 1176 1503 1196
rect 1519 1176 1531 1196
rect 1549 1176 1561 1196
rect 1571 1156 1583 1196
rect 1611 1176 1623 1196
rect 1631 1176 1643 1196
rect 1659 1156 1671 1196
rect 1689 1156 1701 1196
rect 1737 1176 1749 1196
rect 1757 1176 1769 1196
rect 1777 1176 1789 1196
rect 1821 1156 1833 1196
rect 1841 1176 1853 1196
rect 1873 1176 1885 1196
rect 1903 1176 1915 1196
rect 1925 1176 1937 1196
rect 1951 1176 1963 1196
rect 1979 1176 1991 1196
rect 2009 1176 2021 1196
rect 2031 1156 2043 1196
rect 2071 1176 2083 1196
rect 2091 1176 2103 1196
rect 2117 1176 2129 1196
rect 2137 1176 2149 1196
rect 2157 1176 2169 1196
rect 2197 1176 2209 1196
rect 2217 1176 2229 1196
rect 2237 1176 2249 1196
rect 2291 1176 2303 1196
rect 2311 1176 2323 1196
rect 2337 1156 2349 1196
rect 2359 1176 2371 1196
rect 2389 1176 2401 1196
rect 2417 1176 2429 1196
rect 2443 1176 2455 1196
rect 2465 1176 2477 1196
rect 2495 1176 2507 1196
rect 2527 1176 2539 1196
rect 2547 1156 2559 1196
rect 2577 1176 2589 1196
rect 2597 1176 2609 1196
rect 2637 1156 2649 1196
rect 2657 1168 2669 1196
rect 2677 1156 2689 1196
rect 2697 1156 2709 1196
rect 2737 1156 2749 1196
rect 2757 1166 2769 1196
rect 2777 1156 2789 1196
rect 2797 1156 2809 1184
rect 2817 1156 2829 1196
rect 2857 1176 2869 1196
rect 2877 1176 2889 1196
rect 2897 1176 2909 1196
rect 2959 1156 2971 1196
rect 2989 1156 3001 1196
rect 3017 1156 3029 1196
rect 3047 1156 3059 1196
rect 3067 1156 3079 1196
rect 3117 1156 3129 1196
rect 3137 1168 3149 1196
rect 3157 1156 3169 1196
rect 3177 1156 3189 1196
rect 3217 1176 3229 1196
rect 3237 1176 3249 1196
rect 3257 1176 3269 1196
rect 3277 1156 3289 1196
rect 3339 1156 3351 1196
rect 3369 1156 3381 1196
rect 3419 1156 3431 1196
rect 3449 1156 3461 1196
rect 3479 1156 3491 1196
rect 3509 1156 3521 1196
rect 3559 1156 3571 1196
rect 3589 1156 3601 1196
rect 3637 1156 3649 1196
rect 3657 1168 3669 1196
rect 3677 1156 3689 1196
rect 3697 1156 3709 1196
rect 3774 1138 3786 1196
rect 3810 1136 3822 1196
rect 3840 1156 3852 1196
rect 3868 1156 3880 1196
rect 3890 1176 3902 1196
rect 3951 1176 3963 1196
rect 3971 1176 3983 1196
rect 4034 1138 4046 1196
rect 4070 1136 4082 1196
rect 4100 1156 4112 1196
rect 4128 1156 4140 1196
rect 4150 1176 4162 1196
rect 4197 1176 4209 1196
rect 4217 1176 4229 1196
rect 4278 1176 4290 1196
rect 4300 1156 4312 1196
rect 4328 1156 4340 1196
rect 4371 1156 4383 1196
rect 4391 1156 4403 1196
rect 4411 1168 4423 1196
rect 4431 1156 4443 1196
rect 4457 1156 4469 1196
rect 4477 1168 4489 1196
rect 4497 1156 4509 1196
rect 4517 1156 4529 1196
rect 4557 1176 4569 1196
rect 4577 1176 4589 1196
rect 4597 1176 4609 1196
rect 4659 1156 4671 1196
rect 4689 1156 4701 1196
rect 4731 1176 4743 1196
rect 4751 1176 4763 1196
rect 21 744 33 784
rect 41 744 53 764
rect 73 744 85 764
rect 103 744 115 764
rect 125 744 137 764
rect 151 744 163 764
rect 179 744 191 764
rect 209 744 221 764
rect 231 744 243 784
rect 259 744 271 784
rect 289 744 301 784
rect 351 744 363 784
rect 371 744 383 784
rect 391 744 403 772
rect 411 744 423 784
rect 441 744 453 784
rect 461 744 473 764
rect 493 744 505 764
rect 523 744 535 764
rect 545 744 557 764
rect 571 744 583 764
rect 599 744 611 764
rect 629 744 641 764
rect 651 744 663 784
rect 679 744 691 784
rect 709 744 721 784
rect 771 744 783 784
rect 791 744 803 784
rect 811 744 823 772
rect 831 744 843 784
rect 871 744 883 784
rect 891 744 903 784
rect 911 744 923 772
rect 931 744 943 784
rect 971 744 983 764
rect 991 744 1003 764
rect 1031 744 1043 764
rect 1051 744 1063 764
rect 1071 744 1083 764
rect 1097 744 1109 764
rect 1117 744 1129 764
rect 1137 744 1149 764
rect 1199 744 1211 784
rect 1229 744 1241 784
rect 1279 744 1291 784
rect 1309 744 1321 784
rect 1359 744 1371 784
rect 1389 744 1401 784
rect 1438 744 1450 764
rect 1460 744 1472 784
rect 1488 744 1500 784
rect 1541 744 1553 784
rect 1561 744 1573 784
rect 1591 744 1603 784
rect 1620 744 1632 784
rect 1648 744 1660 784
rect 1670 744 1682 764
rect 1717 744 1729 784
rect 1737 744 1749 784
rect 1757 744 1769 784
rect 1777 744 1789 784
rect 1797 744 1809 784
rect 1817 744 1829 784
rect 1837 744 1849 784
rect 1857 744 1869 784
rect 1877 744 1889 784
rect 1939 744 1951 784
rect 1969 744 1981 784
rect 2011 744 2023 764
rect 2031 744 2043 764
rect 2051 744 2063 764
rect 2077 744 2089 784
rect 2097 744 2109 772
rect 2117 744 2129 784
rect 2137 744 2149 784
rect 2177 744 2189 784
rect 2197 744 2209 772
rect 2217 744 2229 784
rect 2237 744 2249 784
rect 2277 744 2289 784
rect 2297 744 2309 772
rect 2317 744 2329 784
rect 2337 744 2349 784
rect 2379 744 2391 784
rect 2409 744 2421 784
rect 2471 744 2483 764
rect 2491 744 2503 764
rect 2517 744 2529 784
rect 2539 744 2551 764
rect 2569 744 2581 764
rect 2597 744 2609 764
rect 2623 744 2635 764
rect 2645 744 2657 764
rect 2675 744 2687 764
rect 2707 744 2719 764
rect 2727 744 2739 784
rect 2771 744 2783 784
rect 2791 744 2803 784
rect 2811 744 2823 772
rect 2831 744 2843 784
rect 2871 744 2883 764
rect 2891 744 2903 764
rect 2917 744 2929 764
rect 2937 744 2949 764
rect 2978 744 2990 804
rect 3014 744 3026 802
rect 3077 744 3089 764
rect 3097 744 3109 764
rect 3159 744 3171 784
rect 3189 744 3201 784
rect 3217 744 3229 764
rect 3237 744 3249 764
rect 3257 744 3269 764
rect 3277 744 3289 784
rect 3319 744 3331 784
rect 3349 744 3361 784
rect 3399 744 3411 784
rect 3429 744 3441 784
rect 3491 744 3503 764
rect 3511 744 3523 764
rect 3531 744 3543 764
rect 3559 744 3571 784
rect 3589 744 3601 784
rect 3674 744 3686 802
rect 3710 744 3722 804
rect 3774 744 3786 802
rect 3810 744 3822 804
rect 3839 744 3851 784
rect 3869 744 3881 784
rect 3954 744 3966 802
rect 3990 744 4002 804
rect 4031 744 4043 764
rect 4051 744 4063 764
rect 4091 744 4103 784
rect 4111 744 4123 784
rect 4131 744 4143 772
rect 4151 744 4163 784
rect 4191 744 4203 784
rect 4211 744 4223 784
rect 4231 744 4243 772
rect 4251 744 4263 784
rect 4298 744 4310 764
rect 4320 744 4332 784
rect 4348 744 4360 784
rect 4378 744 4390 804
rect 4414 744 4426 802
rect 4514 744 4526 802
rect 4550 744 4562 804
rect 4598 744 4610 764
rect 4620 744 4632 784
rect 4648 744 4660 784
rect 4678 744 4690 804
rect 4714 744 4726 802
rect 21 676 33 716
rect 41 696 53 716
rect 73 696 85 716
rect 103 696 115 716
rect 125 696 137 716
rect 151 696 163 716
rect 179 696 191 716
rect 209 696 221 716
rect 231 676 243 716
rect 257 696 269 716
rect 277 696 289 716
rect 317 676 329 716
rect 337 688 349 716
rect 357 676 369 716
rect 377 676 389 716
rect 419 676 431 716
rect 449 676 461 716
rect 497 696 509 716
rect 519 676 531 716
rect 539 676 551 716
rect 591 696 603 716
rect 611 696 623 716
rect 637 676 649 716
rect 659 696 671 716
rect 689 696 701 716
rect 717 696 729 716
rect 743 696 755 716
rect 765 696 777 716
rect 795 696 807 716
rect 827 696 839 716
rect 847 676 859 716
rect 877 676 889 716
rect 897 688 909 716
rect 917 676 929 716
rect 937 676 949 716
rect 991 696 1003 716
rect 1011 696 1023 716
rect 1031 696 1043 716
rect 1057 696 1069 716
rect 1077 696 1089 716
rect 1097 696 1109 716
rect 1117 676 1129 716
rect 1171 676 1183 716
rect 1191 676 1203 716
rect 1211 688 1223 716
rect 1231 676 1243 716
rect 1281 676 1293 716
rect 1301 676 1313 716
rect 1331 676 1343 716
rect 1357 696 1369 716
rect 1377 696 1389 716
rect 1397 696 1409 716
rect 1437 696 1449 716
rect 1459 676 1471 716
rect 1479 676 1491 716
rect 1521 676 1533 716
rect 1541 696 1553 716
rect 1573 696 1585 716
rect 1603 696 1615 716
rect 1625 696 1637 716
rect 1651 696 1663 716
rect 1679 696 1691 716
rect 1709 696 1721 716
rect 1731 676 1743 716
rect 1757 696 1769 716
rect 1779 676 1791 716
rect 1799 676 1811 716
rect 1851 696 1863 716
rect 1871 696 1883 716
rect 1891 696 1903 716
rect 1931 696 1943 716
rect 1951 696 1963 716
rect 1971 696 1983 716
rect 2011 696 2023 716
rect 2031 696 2043 716
rect 2057 696 2069 716
rect 2077 696 2089 716
rect 2097 696 2109 716
rect 2137 676 2149 716
rect 2159 696 2171 716
rect 2189 696 2201 716
rect 2217 696 2229 716
rect 2243 696 2255 716
rect 2265 696 2277 716
rect 2295 696 2307 716
rect 2327 696 2339 716
rect 2347 676 2359 716
rect 2380 676 2392 716
rect 2408 676 2420 716
rect 2436 676 2448 716
rect 2511 676 2523 716
rect 2531 696 2543 716
rect 2551 696 2563 716
rect 2571 696 2583 716
rect 2618 696 2630 716
rect 2640 676 2652 716
rect 2668 676 2680 716
rect 2718 696 2730 716
rect 2740 676 2752 716
rect 2768 676 2780 716
rect 2797 696 2809 716
rect 2817 696 2829 716
rect 2871 676 2883 716
rect 2891 676 2903 716
rect 2911 688 2923 716
rect 2931 676 2943 716
rect 2957 676 2969 716
rect 2977 688 2989 716
rect 2997 676 3009 716
rect 3017 676 3029 716
rect 3059 676 3071 716
rect 3089 676 3101 716
rect 3151 696 3163 716
rect 3171 696 3183 716
rect 3197 696 3209 716
rect 3217 696 3229 716
rect 3294 658 3306 716
rect 3330 656 3342 716
rect 3371 696 3383 716
rect 3391 696 3403 716
rect 3411 696 3423 716
rect 3437 676 3449 716
rect 3457 688 3469 716
rect 3477 676 3489 716
rect 3497 676 3509 716
rect 3540 676 3552 716
rect 3568 676 3580 716
rect 3590 696 3602 716
rect 3658 696 3670 716
rect 3680 676 3692 716
rect 3708 676 3720 716
rect 3772 676 3784 716
rect 3800 676 3812 716
rect 3828 676 3840 716
rect 3894 658 3906 716
rect 3930 656 3942 716
rect 3994 658 4006 716
rect 4030 656 4042 716
rect 4057 696 4069 716
rect 4077 696 4089 716
rect 4118 656 4130 716
rect 4154 658 4166 716
rect 4218 656 4230 716
rect 4254 658 4266 716
rect 4354 658 4366 716
rect 4390 656 4402 716
rect 4454 658 4466 716
rect 4490 656 4502 716
rect 4517 696 4529 716
rect 4537 696 4549 716
rect 4591 676 4603 716
rect 4611 676 4623 716
rect 4631 688 4643 716
rect 4651 676 4663 716
rect 4677 676 4689 716
rect 4697 688 4709 716
rect 4717 676 4729 716
rect 4737 676 4749 716
rect 21 264 33 304
rect 41 264 53 284
rect 73 264 85 284
rect 103 264 115 284
rect 125 264 137 284
rect 151 264 163 284
rect 179 264 191 284
rect 209 264 221 284
rect 231 264 243 304
rect 259 264 271 304
rect 289 264 301 304
rect 351 264 363 304
rect 371 264 383 304
rect 391 264 403 292
rect 411 264 423 304
rect 437 264 449 284
rect 457 264 469 284
rect 499 264 511 304
rect 529 264 541 304
rect 591 264 603 304
rect 611 264 623 304
rect 631 264 643 292
rect 651 264 663 304
rect 677 264 689 304
rect 697 264 709 292
rect 717 264 729 304
rect 737 264 749 304
rect 777 264 789 304
rect 797 264 809 292
rect 817 264 829 304
rect 837 264 849 304
rect 891 264 903 304
rect 911 264 923 304
rect 931 264 943 292
rect 951 264 963 304
rect 977 264 989 284
rect 997 264 1009 284
rect 1039 264 1051 304
rect 1069 264 1081 304
rect 1138 264 1150 284
rect 1160 264 1172 304
rect 1188 264 1200 304
rect 1231 264 1243 284
rect 1251 264 1263 284
rect 1291 264 1303 304
rect 1311 264 1323 304
rect 1331 264 1343 292
rect 1351 264 1363 304
rect 1391 264 1403 284
rect 1411 264 1423 284
rect 1431 264 1443 284
rect 1457 264 1469 304
rect 1477 264 1489 292
rect 1497 264 1509 304
rect 1517 264 1529 304
rect 1559 264 1571 304
rect 1589 264 1601 304
rect 1637 264 1649 304
rect 1659 264 1671 284
rect 1689 264 1701 284
rect 1717 264 1729 284
rect 1743 264 1755 284
rect 1765 264 1777 284
rect 1795 264 1807 284
rect 1827 264 1839 284
rect 1847 264 1859 304
rect 1899 264 1911 304
rect 1929 264 1941 304
rect 1971 264 1983 304
rect 1991 264 2003 304
rect 2011 264 2023 292
rect 2031 264 2043 304
rect 2061 264 2073 304
rect 2081 264 2093 284
rect 2113 264 2125 284
rect 2143 264 2155 284
rect 2165 264 2177 284
rect 2191 264 2203 284
rect 2219 264 2231 284
rect 2249 264 2261 284
rect 2271 264 2283 304
rect 2311 264 2323 284
rect 2331 264 2343 284
rect 2357 264 2369 284
rect 2377 264 2389 284
rect 2397 264 2409 284
rect 2437 264 2449 284
rect 2457 264 2469 284
rect 2519 264 2531 304
rect 2549 264 2561 304
rect 2577 264 2589 304
rect 2599 264 2611 284
rect 2629 264 2641 284
rect 2657 264 2669 284
rect 2683 264 2695 284
rect 2705 264 2717 284
rect 2735 264 2747 284
rect 2767 264 2779 284
rect 2787 264 2799 304
rect 2819 264 2831 304
rect 2849 264 2861 304
rect 2900 264 2912 304
rect 2928 264 2940 304
rect 2956 264 2968 304
rect 3017 264 3029 284
rect 3037 264 3049 284
rect 3057 264 3069 284
rect 3097 264 3109 284
rect 3117 264 3129 284
rect 3194 264 3206 322
rect 3230 264 3242 324
rect 3294 264 3306 322
rect 3330 264 3342 324
rect 3357 264 3369 304
rect 3377 264 3389 292
rect 3397 264 3409 304
rect 3417 264 3429 304
rect 3471 264 3483 284
rect 3491 264 3503 284
rect 3519 264 3531 304
rect 3549 264 3561 304
rect 3599 264 3611 304
rect 3629 264 3641 304
rect 3677 264 3689 304
rect 3697 264 3709 292
rect 3717 264 3729 304
rect 3737 264 3749 304
rect 3791 264 3803 284
rect 3811 264 3823 284
rect 3831 264 3843 284
rect 3871 264 3883 284
rect 3891 264 3903 284
rect 3911 264 3923 284
rect 3937 264 3949 304
rect 3967 264 3979 304
rect 3987 264 3999 304
rect 4037 264 4049 284
rect 4057 264 4069 284
rect 4077 264 4089 284
rect 4138 264 4150 284
rect 4160 264 4172 304
rect 4188 264 4200 304
rect 4254 264 4266 322
rect 4290 264 4302 324
rect 4320 264 4332 304
rect 4348 264 4360 304
rect 4370 264 4382 284
rect 4417 264 4429 284
rect 4437 264 4449 284
rect 4491 264 4503 304
rect 4511 264 4523 304
rect 4531 264 4543 292
rect 4551 264 4563 304
rect 4577 264 4589 284
rect 4597 264 4609 284
rect 4637 264 4649 284
rect 4657 264 4669 284
rect 4697 264 4709 284
rect 4717 264 4729 284
rect 21 196 33 236
rect 41 216 53 236
rect 73 216 85 236
rect 103 216 115 236
rect 125 216 137 236
rect 151 216 163 236
rect 179 216 191 236
rect 209 216 221 236
rect 231 196 243 236
rect 260 196 272 236
rect 288 196 300 236
rect 316 196 328 236
rect 377 216 389 236
rect 397 216 409 236
rect 417 216 429 236
rect 458 176 470 236
rect 494 178 506 236
rect 571 196 583 236
rect 591 216 603 236
rect 611 216 623 236
rect 631 216 643 236
rect 678 216 690 236
rect 700 196 712 236
rect 728 196 740 236
rect 757 196 769 236
rect 779 216 791 236
rect 809 216 821 236
rect 837 216 849 236
rect 863 216 875 236
rect 885 216 897 236
rect 915 216 927 236
rect 947 216 959 236
rect 967 196 979 236
rect 1011 196 1023 236
rect 1031 196 1043 236
rect 1051 208 1063 236
rect 1071 196 1083 236
rect 1111 216 1123 236
rect 1131 216 1143 236
rect 1171 216 1183 236
rect 1191 216 1203 236
rect 1211 216 1223 236
rect 1251 216 1263 236
rect 1271 216 1283 236
rect 1311 196 1323 236
rect 1331 196 1343 236
rect 1351 208 1363 236
rect 1371 196 1383 236
rect 1411 216 1423 236
rect 1431 216 1443 236
rect 1471 216 1483 236
rect 1491 216 1503 236
rect 1517 216 1529 236
rect 1537 216 1549 236
rect 1557 216 1569 236
rect 1618 216 1630 236
rect 1640 196 1652 236
rect 1668 196 1680 236
rect 1701 196 1713 236
rect 1721 216 1733 236
rect 1753 216 1765 236
rect 1783 216 1795 236
rect 1805 216 1817 236
rect 1831 216 1843 236
rect 1859 216 1871 236
rect 1889 216 1901 236
rect 1911 196 1923 236
rect 1951 196 1963 236
rect 1971 196 1983 236
rect 1991 208 2003 236
rect 2011 196 2023 236
rect 2037 216 2049 236
rect 2057 216 2069 236
rect 2097 216 2109 236
rect 2117 216 2129 236
rect 2137 216 2149 236
rect 2177 216 2189 236
rect 2197 216 2209 236
rect 2217 216 2229 236
rect 2271 216 2283 236
rect 2291 216 2303 236
rect 2311 216 2323 236
rect 2337 216 2349 236
rect 2357 216 2369 236
rect 2377 216 2389 236
rect 2431 216 2443 236
rect 2451 216 2463 236
rect 2477 196 2489 236
rect 2499 216 2511 236
rect 2529 216 2541 236
rect 2557 216 2569 236
rect 2583 216 2595 236
rect 2605 216 2617 236
rect 2635 216 2647 236
rect 2667 216 2679 236
rect 2687 196 2699 236
rect 2717 196 2729 236
rect 2739 216 2751 236
rect 2769 216 2781 236
rect 2797 216 2809 236
rect 2823 216 2835 236
rect 2845 216 2857 236
rect 2875 216 2887 236
rect 2907 216 2919 236
rect 2927 196 2939 236
rect 2957 196 2969 236
rect 2977 206 2989 236
rect 2997 196 3009 236
rect 3017 196 3029 224
rect 3037 196 3049 236
rect 3091 196 3103 236
rect 3111 216 3123 236
rect 3131 216 3143 236
rect 3151 216 3163 236
rect 3177 196 3189 236
rect 3197 208 3209 236
rect 3217 196 3229 236
rect 3237 196 3249 236
rect 3291 216 3303 236
rect 3311 216 3323 236
rect 3339 196 3351 236
rect 3369 196 3381 236
rect 3454 178 3466 236
rect 3490 176 3502 236
rect 3531 216 3543 236
rect 3551 216 3563 236
rect 3598 216 3610 236
rect 3620 196 3632 236
rect 3648 196 3660 236
rect 3691 216 3703 236
rect 3711 216 3723 236
rect 3731 216 3743 236
rect 3757 216 3769 236
rect 3777 216 3789 236
rect 3817 196 3829 236
rect 3837 208 3849 236
rect 3857 196 3869 236
rect 3877 196 3889 236
rect 3917 216 3929 236
rect 3937 216 3949 236
rect 3957 216 3969 236
rect 4034 178 4046 236
rect 4070 176 4082 236
rect 4099 196 4111 236
rect 4129 196 4141 236
rect 4214 178 4226 236
rect 4250 176 4262 236
rect 4299 196 4311 236
rect 4329 196 4341 236
rect 4394 178 4406 236
rect 4430 176 4442 236
rect 4459 196 4471 236
rect 4489 196 4501 236
rect 4538 176 4550 236
rect 4574 178 4586 236
rect 4658 216 4670 236
rect 4680 196 4692 236
rect 4708 196 4720 236
<< pdcontact >>
rect 29 4344 41 4424
rect 49 4344 61 4424
rect 71 4344 83 4384
rect 111 4344 123 4384
rect 131 4344 143 4384
rect 151 4344 163 4384
rect 196 4344 208 4384
rect 218 4344 230 4424
rect 246 4344 258 4424
rect 277 4344 289 4384
rect 299 4344 311 4424
rect 319 4344 331 4424
rect 383 4344 395 4424
rect 411 4344 423 4424
rect 463 4344 475 4424
rect 491 4344 503 4424
rect 517 4344 529 4384
rect 539 4344 551 4424
rect 559 4344 571 4424
rect 611 4344 623 4384
rect 631 4344 643 4384
rect 657 4344 669 4424
rect 685 4344 697 4424
rect 737 4344 749 4384
rect 757 4344 769 4384
rect 797 4344 809 4424
rect 817 4344 829 4364
rect 847 4344 859 4364
rect 875 4344 887 4384
rect 901 4344 913 4384
rect 921 4344 933 4384
rect 953 4344 965 4384
rect 987 4344 999 4384
rect 1007 4344 1019 4424
rect 1042 4344 1054 4424
rect 1070 4344 1082 4424
rect 1092 4344 1104 4384
rect 1137 4344 1149 4424
rect 1157 4344 1169 4364
rect 1187 4344 1199 4364
rect 1215 4344 1227 4384
rect 1241 4344 1253 4384
rect 1261 4344 1273 4384
rect 1293 4344 1305 4384
rect 1327 4344 1339 4384
rect 1347 4344 1359 4424
rect 1382 4344 1394 4424
rect 1410 4344 1422 4424
rect 1432 4344 1444 4384
rect 1481 4344 1493 4424
rect 1501 4344 1513 4384
rect 1535 4344 1547 4384
rect 1567 4344 1579 4384
rect 1587 4344 1599 4384
rect 1613 4344 1625 4384
rect 1641 4344 1653 4364
rect 1671 4344 1683 4364
rect 1691 4344 1703 4424
rect 1717 4344 1729 4384
rect 1737 4344 1749 4384
rect 1757 4344 1769 4384
rect 1797 4344 1809 4424
rect 1817 4344 1829 4364
rect 1847 4344 1859 4364
rect 1875 4344 1887 4384
rect 1901 4344 1913 4384
rect 1921 4344 1933 4384
rect 1953 4344 1965 4384
rect 1987 4344 1999 4384
rect 2007 4344 2019 4424
rect 2037 4344 2049 4424
rect 2067 4344 2089 4424
rect 2107 4344 2119 4424
rect 2171 4344 2183 4384
rect 2191 4344 2203 4380
rect 2211 4344 2223 4384
rect 2231 4344 2243 4384
rect 2276 4344 2288 4384
rect 2298 4344 2310 4424
rect 2326 4344 2338 4424
rect 2371 4344 2383 4384
rect 2391 4344 2403 4384
rect 2417 4344 2429 4424
rect 2445 4344 2457 4424
rect 2511 4344 2523 4384
rect 2531 4344 2543 4384
rect 2562 4344 2574 4424
rect 2590 4344 2602 4424
rect 2612 4344 2624 4384
rect 2657 4344 2669 4384
rect 2679 4344 2691 4424
rect 2699 4344 2711 4424
rect 2737 4344 2749 4384
rect 2759 4344 2771 4424
rect 2779 4344 2791 4424
rect 2829 4344 2841 4424
rect 2849 4344 2861 4424
rect 2871 4344 2883 4384
rect 2911 4344 2923 4384
rect 2931 4344 2943 4380
rect 2951 4344 2963 4384
rect 2971 4344 2983 4384
rect 3007 4344 3019 4424
rect 3027 4344 3039 4424
rect 3051 4344 3063 4384
rect 3071 4344 3083 4384
rect 3109 4344 3121 4424
rect 3129 4344 3141 4424
rect 3151 4344 3163 4384
rect 3191 4344 3203 4384
rect 3211 4344 3223 4380
rect 3231 4344 3243 4384
rect 3251 4344 3263 4384
rect 3277 4344 3289 4384
rect 3297 4344 3309 4384
rect 3317 4344 3329 4384
rect 3357 4344 3369 4416
rect 3377 4344 3389 4412
rect 3397 4344 3409 4424
rect 3417 4344 3429 4424
rect 3457 4344 3469 4384
rect 3477 4344 3489 4384
rect 3517 4344 3529 4384
rect 3537 4344 3549 4384
rect 3557 4344 3569 4384
rect 3597 4344 3609 4384
rect 3617 4344 3629 4384
rect 3637 4344 3649 4380
rect 3657 4344 3669 4384
rect 3697 4344 3709 4416
rect 3717 4344 3729 4412
rect 3737 4344 3749 4424
rect 3757 4344 3769 4424
rect 3802 4344 3814 4424
rect 3830 4344 3842 4424
rect 3852 4344 3864 4384
rect 3916 4344 3928 4384
rect 3938 4344 3950 4424
rect 3966 4344 3978 4424
rect 4011 4344 4023 4384
rect 4031 4344 4043 4380
rect 4051 4344 4063 4384
rect 4071 4344 4083 4384
rect 4111 4344 4123 4384
rect 4131 4344 4143 4380
rect 4151 4344 4163 4384
rect 4171 4344 4183 4384
rect 4197 4344 4209 4416
rect 4217 4344 4229 4412
rect 4237 4344 4249 4424
rect 4257 4344 4269 4424
rect 4297 4344 4309 4384
rect 4317 4344 4329 4384
rect 4337 4344 4349 4384
rect 4391 4344 4403 4424
rect 4411 4344 4423 4424
rect 4431 4344 4443 4412
rect 4451 4344 4463 4416
rect 4491 4344 4503 4384
rect 4511 4344 4523 4384
rect 4537 4344 4549 4384
rect 4557 4344 4569 4384
rect 4577 4344 4589 4380
rect 4597 4344 4609 4384
rect 4637 4344 4649 4384
rect 4657 4344 4669 4384
rect 4677 4344 4689 4380
rect 4697 4344 4709 4384
rect 36 4276 48 4316
rect 58 4236 70 4316
rect 86 4236 98 4316
rect 127 4236 139 4316
rect 147 4236 159 4316
rect 171 4276 183 4316
rect 191 4276 203 4316
rect 217 4236 229 4316
rect 245 4236 257 4316
rect 311 4236 323 4316
rect 331 4236 343 4316
rect 351 4248 363 4316
rect 371 4244 383 4316
rect 397 4276 409 4316
rect 417 4276 429 4316
rect 441 4236 453 4316
rect 461 4236 473 4316
rect 511 4236 523 4316
rect 531 4236 543 4316
rect 551 4248 563 4316
rect 571 4244 583 4316
rect 597 4276 609 4316
rect 617 4276 629 4316
rect 637 4280 649 4316
rect 657 4276 669 4316
rect 697 4244 709 4316
rect 717 4248 729 4316
rect 737 4236 749 4316
rect 757 4236 769 4316
rect 797 4276 809 4316
rect 817 4276 829 4316
rect 841 4236 853 4316
rect 861 4236 873 4316
rect 916 4276 928 4316
rect 938 4236 950 4316
rect 966 4236 978 4316
rect 1011 4276 1023 4316
rect 1031 4276 1043 4316
rect 1057 4236 1069 4316
rect 1085 4236 1097 4316
rect 1137 4236 1149 4316
rect 1165 4236 1177 4316
rect 1217 4236 1229 4316
rect 1245 4236 1257 4316
rect 1297 4276 1309 4316
rect 1317 4276 1329 4316
rect 1357 4236 1369 4316
rect 1377 4296 1389 4316
rect 1407 4296 1419 4316
rect 1435 4276 1447 4316
rect 1461 4276 1473 4316
rect 1481 4276 1493 4316
rect 1513 4276 1525 4316
rect 1547 4276 1559 4316
rect 1567 4236 1579 4316
rect 1602 4236 1614 4316
rect 1630 4236 1642 4316
rect 1652 4276 1664 4316
rect 1697 4236 1709 4316
rect 1725 4236 1737 4316
rect 1791 4276 1803 4316
rect 1811 4276 1823 4316
rect 1837 4236 1849 4316
rect 1857 4296 1869 4316
rect 1887 4296 1899 4316
rect 1915 4276 1927 4316
rect 1941 4276 1953 4316
rect 1961 4276 1973 4316
rect 1993 4276 2005 4316
rect 2027 4276 2039 4316
rect 2047 4236 2059 4316
rect 2091 4276 2103 4316
rect 2111 4276 2123 4316
rect 2131 4276 2143 4316
rect 2157 4236 2169 4316
rect 2187 4237 2199 4316
rect 2207 4237 2219 4316
rect 2271 4236 2283 4316
rect 2291 4236 2303 4304
rect 2311 4238 2323 4316
rect 2331 4250 2343 4316
rect 2351 4238 2363 4316
rect 2377 4276 2389 4316
rect 2397 4276 2409 4316
rect 2417 4276 2429 4316
rect 2476 4276 2488 4316
rect 2498 4236 2510 4316
rect 2526 4236 2538 4316
rect 2583 4236 2595 4316
rect 2611 4236 2623 4316
rect 2637 4244 2649 4316
rect 2657 4248 2669 4316
rect 2677 4236 2689 4316
rect 2697 4236 2709 4316
rect 2751 4236 2763 4316
rect 2771 4236 2783 4316
rect 2791 4248 2803 4316
rect 2811 4244 2823 4316
rect 2837 4276 2849 4316
rect 2859 4236 2871 4316
rect 2879 4236 2891 4316
rect 2931 4276 2943 4316
rect 2951 4280 2963 4316
rect 2971 4276 2983 4316
rect 2991 4276 3003 4316
rect 3031 4276 3043 4316
rect 3051 4280 3063 4316
rect 3071 4276 3083 4316
rect 3091 4276 3103 4316
rect 3117 4276 3129 4316
rect 3137 4276 3149 4316
rect 3157 4276 3169 4316
rect 3211 4276 3223 4316
rect 3231 4276 3243 4316
rect 3271 4276 3283 4316
rect 3291 4280 3303 4316
rect 3311 4276 3323 4316
rect 3331 4276 3343 4316
rect 3371 4276 3383 4316
rect 3391 4280 3403 4316
rect 3411 4276 3423 4316
rect 3431 4276 3443 4316
rect 3471 4276 3483 4316
rect 3491 4280 3503 4316
rect 3511 4276 3523 4316
rect 3531 4276 3543 4316
rect 3571 4276 3583 4316
rect 3591 4280 3603 4316
rect 3611 4276 3623 4316
rect 3631 4276 3643 4316
rect 3657 4276 3669 4316
rect 3677 4276 3689 4316
rect 3697 4280 3709 4316
rect 3717 4276 3729 4316
rect 3757 4244 3769 4316
rect 3777 4248 3789 4316
rect 3797 4236 3809 4316
rect 3817 4236 3829 4316
rect 3862 4236 3874 4316
rect 3890 4236 3902 4316
rect 3912 4276 3924 4316
rect 3957 4276 3969 4316
rect 3977 4276 3989 4316
rect 4017 4244 4029 4316
rect 4037 4248 4049 4316
rect 4057 4236 4069 4316
rect 4077 4236 4089 4316
rect 4131 4276 4143 4316
rect 4151 4280 4163 4316
rect 4171 4276 4183 4316
rect 4191 4276 4203 4316
rect 4217 4276 4229 4316
rect 4237 4276 4249 4316
rect 4257 4280 4269 4316
rect 4277 4276 4289 4316
rect 4317 4244 4329 4316
rect 4337 4248 4349 4316
rect 4357 4236 4369 4316
rect 4377 4236 4389 4316
rect 4422 4236 4434 4316
rect 4450 4236 4462 4316
rect 4472 4276 4484 4316
rect 4517 4238 4529 4316
rect 4537 4250 4549 4316
rect 4557 4238 4569 4316
rect 4577 4236 4589 4304
rect 4597 4236 4609 4316
rect 4663 4236 4675 4316
rect 4691 4236 4703 4316
rect 31 3864 43 3904
rect 51 3864 63 3904
rect 71 3864 83 3904
rect 111 3864 123 3904
rect 131 3864 143 3904
rect 151 3864 163 3904
rect 203 3864 215 3944
rect 231 3864 243 3944
rect 262 3864 274 3944
rect 290 3864 302 3944
rect 312 3864 324 3904
rect 371 3864 383 3904
rect 391 3864 403 3904
rect 431 3864 443 3904
rect 451 3864 463 3904
rect 503 3864 515 3944
rect 531 3864 543 3944
rect 557 3864 569 3904
rect 577 3864 589 3904
rect 601 3864 613 3944
rect 621 3864 633 3944
rect 662 3864 674 3944
rect 690 3864 702 3944
rect 712 3864 724 3904
rect 757 3864 769 3904
rect 777 3864 789 3904
rect 822 3864 834 3944
rect 850 3864 862 3944
rect 872 3864 884 3904
rect 917 3864 929 3904
rect 937 3864 949 3904
rect 957 3864 969 3904
rect 1011 3864 1023 3904
rect 1031 3864 1043 3904
rect 1083 3864 1095 3944
rect 1111 3864 1123 3944
rect 1137 3864 1149 3904
rect 1157 3864 1169 3904
rect 1197 3864 1209 3944
rect 1225 3864 1237 3944
rect 1277 3864 1289 3904
rect 1297 3864 1309 3904
rect 1363 3864 1375 3944
rect 1391 3864 1403 3944
rect 1431 3864 1443 3904
rect 1451 3864 1463 3904
rect 1482 3864 1494 3944
rect 1510 3864 1522 3944
rect 1532 3864 1544 3904
rect 1577 3864 1589 3944
rect 1607 3864 1629 3944
rect 1647 3864 1659 3944
rect 1697 3864 1709 3904
rect 1717 3864 1729 3904
rect 1737 3864 1749 3904
rect 1791 3864 1803 3944
rect 1811 3864 1823 3944
rect 1831 3864 1843 3932
rect 1851 3864 1863 3936
rect 1877 3864 1889 3904
rect 1897 3864 1909 3904
rect 1917 3864 1929 3900
rect 1937 3864 1949 3904
rect 1996 3864 2008 3904
rect 2018 3864 2030 3944
rect 2046 3864 2058 3944
rect 2091 3864 2103 3904
rect 2111 3864 2123 3904
rect 2151 3864 2163 3904
rect 2171 3864 2183 3900
rect 2191 3864 2203 3904
rect 2211 3864 2223 3904
rect 2251 3864 2263 3904
rect 2271 3864 2283 3900
rect 2291 3864 2303 3904
rect 2311 3864 2323 3904
rect 2351 3864 2363 3944
rect 2371 3864 2383 3944
rect 2391 3864 2403 3932
rect 2411 3864 2423 3936
rect 2451 3864 2463 3904
rect 2471 3864 2483 3904
rect 2516 3864 2528 3904
rect 2538 3864 2550 3944
rect 2566 3864 2578 3944
rect 2611 3864 2623 3904
rect 2631 3864 2643 3900
rect 2651 3864 2663 3904
rect 2671 3864 2683 3904
rect 2711 3864 2723 3944
rect 2731 3864 2743 3944
rect 2751 3864 2763 3932
rect 2771 3864 2783 3936
rect 2816 3864 2828 3904
rect 2838 3864 2850 3944
rect 2866 3864 2878 3944
rect 2902 3864 2914 3944
rect 2930 3864 2942 3944
rect 2952 3864 2964 3904
rect 3011 3864 3023 3904
rect 3031 3864 3043 3900
rect 3051 3864 3063 3904
rect 3071 3864 3083 3904
rect 3111 3864 3123 3904
rect 3131 3864 3143 3904
rect 3162 3864 3174 3944
rect 3190 3864 3202 3944
rect 3212 3864 3224 3904
rect 3257 3864 3269 3936
rect 3277 3864 3289 3932
rect 3297 3864 3309 3944
rect 3317 3864 3329 3944
rect 3362 3864 3374 3944
rect 3390 3864 3402 3944
rect 3412 3864 3424 3904
rect 3476 3864 3488 3904
rect 3498 3864 3510 3944
rect 3526 3864 3538 3944
rect 3576 3864 3588 3904
rect 3598 3864 3610 3944
rect 3626 3864 3638 3944
rect 3671 3864 3683 3944
rect 3691 3864 3703 3944
rect 3711 3864 3723 3932
rect 3731 3864 3743 3936
rect 3771 3864 3783 3904
rect 3791 3864 3803 3900
rect 3811 3864 3823 3904
rect 3831 3864 3843 3904
rect 3871 3864 3883 3904
rect 3891 3864 3903 3904
rect 3911 3864 3923 3904
rect 3951 3864 3963 3904
rect 3971 3864 3983 3904
rect 3991 3864 4003 3904
rect 4017 3864 4029 3904
rect 4037 3864 4049 3904
rect 4057 3864 4069 3904
rect 4111 3864 4123 3904
rect 4131 3864 4143 3900
rect 4151 3864 4163 3904
rect 4171 3864 4183 3904
rect 4216 3864 4228 3904
rect 4238 3864 4250 3944
rect 4266 3864 4278 3944
rect 4302 3864 4314 3944
rect 4330 3864 4342 3944
rect 4352 3864 4364 3904
rect 4411 3864 4423 3904
rect 4431 3864 4443 3904
rect 4471 3864 4483 3904
rect 4491 3864 4503 3900
rect 4511 3864 4523 3904
rect 4531 3864 4543 3904
rect 4571 3864 4583 3904
rect 4591 3864 4603 3900
rect 4611 3864 4623 3904
rect 4631 3864 4643 3904
rect 4657 3864 4669 3936
rect 4677 3864 4689 3932
rect 4697 3864 4709 3944
rect 4717 3864 4729 3944
rect 36 3796 48 3836
rect 58 3756 70 3836
rect 86 3756 98 3836
rect 131 3796 143 3836
rect 151 3796 163 3836
rect 177 3756 189 3836
rect 197 3816 209 3836
rect 227 3816 239 3836
rect 255 3796 267 3836
rect 281 3796 293 3836
rect 301 3796 313 3836
rect 333 3796 345 3836
rect 367 3796 379 3836
rect 387 3756 399 3836
rect 436 3796 448 3836
rect 458 3756 470 3836
rect 486 3756 498 3836
rect 517 3796 529 3836
rect 537 3796 549 3836
rect 561 3756 573 3836
rect 581 3756 593 3836
rect 641 3757 653 3836
rect 661 3757 673 3836
rect 691 3756 703 3836
rect 731 3796 743 3836
rect 751 3796 763 3836
rect 771 3796 783 3836
rect 801 3756 813 3836
rect 821 3796 833 3836
rect 855 3796 867 3836
rect 887 3796 899 3836
rect 907 3796 919 3836
rect 933 3796 945 3836
rect 961 3816 973 3836
rect 991 3816 1003 3836
rect 1011 3756 1023 3836
rect 1049 3756 1061 3836
rect 1069 3756 1081 3836
rect 1091 3796 1103 3836
rect 1117 3756 1129 3836
rect 1137 3816 1149 3836
rect 1167 3816 1179 3836
rect 1195 3796 1207 3836
rect 1221 3796 1233 3836
rect 1241 3796 1253 3836
rect 1273 3796 1285 3836
rect 1307 3796 1319 3836
rect 1327 3756 1339 3836
rect 1362 3756 1374 3836
rect 1390 3756 1402 3836
rect 1412 3796 1424 3836
rect 1457 3796 1469 3836
rect 1477 3796 1489 3836
rect 1497 3796 1509 3836
rect 1537 3796 1549 3836
rect 1557 3796 1569 3836
rect 1577 3796 1589 3836
rect 1617 3796 1629 3836
rect 1639 3756 1651 3836
rect 1659 3756 1671 3836
rect 1697 3756 1709 3836
rect 1717 3816 1729 3836
rect 1747 3816 1759 3836
rect 1775 3796 1787 3836
rect 1801 3796 1813 3836
rect 1821 3796 1833 3836
rect 1853 3796 1865 3836
rect 1887 3796 1899 3836
rect 1907 3756 1919 3836
rect 1951 3796 1963 3836
rect 1971 3796 1983 3836
rect 2011 3756 2023 3836
rect 2031 3756 2043 3836
rect 2051 3768 2063 3836
rect 2071 3764 2083 3836
rect 2111 3796 2123 3836
rect 2131 3796 2143 3836
rect 2157 3796 2169 3836
rect 2177 3796 2189 3836
rect 2197 3800 2209 3836
rect 2217 3796 2229 3836
rect 2276 3796 2288 3836
rect 2298 3756 2310 3836
rect 2326 3756 2338 3836
rect 2371 3796 2383 3836
rect 2391 3800 2403 3836
rect 2411 3796 2423 3836
rect 2431 3796 2443 3836
rect 2471 3756 2483 3836
rect 2491 3756 2503 3836
rect 2511 3768 2523 3836
rect 2531 3764 2543 3836
rect 2571 3796 2583 3836
rect 2591 3800 2603 3836
rect 2611 3796 2623 3836
rect 2631 3796 2643 3836
rect 2657 3764 2669 3836
rect 2677 3768 2689 3836
rect 2697 3756 2709 3836
rect 2717 3756 2729 3836
rect 2771 3756 2783 3836
rect 2791 3756 2803 3836
rect 2811 3768 2823 3836
rect 2831 3764 2843 3836
rect 2871 3796 2883 3836
rect 2891 3796 2903 3836
rect 2931 3796 2943 3836
rect 2951 3796 2963 3836
rect 2991 3796 3003 3836
rect 3011 3800 3023 3836
rect 3031 3796 3043 3836
rect 3051 3796 3063 3836
rect 3091 3756 3103 3836
rect 3111 3756 3123 3836
rect 3131 3768 3143 3836
rect 3151 3764 3163 3836
rect 3191 3796 3203 3836
rect 3211 3800 3223 3836
rect 3231 3796 3243 3836
rect 3251 3796 3263 3836
rect 3291 3796 3303 3836
rect 3311 3796 3323 3836
rect 3356 3796 3368 3836
rect 3378 3756 3390 3836
rect 3406 3756 3418 3836
rect 3451 3796 3463 3836
rect 3471 3796 3483 3836
rect 3491 3796 3503 3836
rect 3517 3796 3529 3836
rect 3537 3796 3549 3836
rect 3561 3756 3573 3836
rect 3581 3756 3593 3836
rect 3631 3756 3643 3836
rect 3651 3756 3663 3836
rect 3671 3768 3683 3836
rect 3691 3764 3703 3836
rect 3731 3796 3743 3836
rect 3751 3800 3763 3836
rect 3771 3796 3783 3836
rect 3791 3796 3803 3836
rect 3831 3796 3843 3836
rect 3851 3796 3863 3836
rect 3877 3764 3889 3836
rect 3897 3768 3909 3836
rect 3917 3756 3929 3836
rect 3937 3756 3949 3836
rect 3996 3796 4008 3836
rect 4018 3756 4030 3836
rect 4046 3756 4058 3836
rect 4082 3756 4094 3836
rect 4110 3756 4122 3836
rect 4132 3796 4144 3836
rect 4177 3764 4189 3836
rect 4197 3768 4209 3836
rect 4217 3756 4229 3836
rect 4237 3756 4249 3836
rect 4291 3756 4303 3836
rect 4311 3756 4323 3836
rect 4331 3768 4343 3836
rect 4351 3764 4363 3836
rect 4377 3796 4389 3836
rect 4397 3796 4409 3836
rect 4417 3800 4429 3836
rect 4437 3796 4449 3836
rect 4491 3796 4503 3836
rect 4511 3796 4523 3836
rect 4551 3796 4563 3836
rect 4571 3800 4583 3836
rect 4591 3796 4603 3836
rect 4611 3796 4623 3836
rect 4637 3796 4649 3836
rect 4657 3796 4669 3836
rect 4677 3800 4689 3836
rect 4697 3796 4709 3836
rect 21 3384 33 3464
rect 41 3384 53 3424
rect 75 3384 87 3424
rect 107 3384 119 3424
rect 127 3384 139 3424
rect 153 3384 165 3424
rect 181 3384 193 3404
rect 211 3384 223 3404
rect 231 3384 243 3464
rect 271 3384 283 3424
rect 291 3384 303 3424
rect 311 3384 323 3424
rect 356 3384 368 3424
rect 378 3384 390 3464
rect 406 3384 418 3464
rect 451 3384 463 3424
rect 471 3384 483 3424
rect 491 3384 503 3424
rect 531 3384 543 3424
rect 551 3384 563 3420
rect 571 3384 583 3424
rect 591 3384 603 3424
rect 631 3384 643 3424
rect 651 3384 663 3424
rect 696 3384 708 3424
rect 718 3384 730 3464
rect 746 3384 758 3464
rect 796 3384 808 3424
rect 818 3384 830 3464
rect 846 3384 858 3464
rect 877 3384 889 3424
rect 897 3384 909 3424
rect 963 3384 975 3464
rect 991 3384 1003 3464
rect 1017 3384 1029 3464
rect 1037 3384 1049 3404
rect 1067 3384 1079 3404
rect 1095 3384 1107 3424
rect 1121 3384 1133 3424
rect 1141 3384 1153 3424
rect 1173 3384 1185 3424
rect 1207 3384 1219 3424
rect 1227 3384 1239 3464
rect 1257 3384 1269 3424
rect 1277 3384 1289 3424
rect 1317 3384 1329 3464
rect 1345 3384 1357 3464
rect 1402 3384 1414 3464
rect 1430 3384 1442 3464
rect 1452 3384 1464 3424
rect 1497 3384 1509 3424
rect 1517 3384 1529 3424
rect 1537 3384 1549 3424
rect 1589 3384 1601 3464
rect 1609 3384 1621 3464
rect 1631 3384 1643 3424
rect 1671 3384 1683 3424
rect 1691 3384 1703 3424
rect 1717 3384 1729 3464
rect 1737 3384 1749 3404
rect 1767 3384 1779 3404
rect 1795 3384 1807 3424
rect 1821 3384 1833 3424
rect 1841 3384 1853 3424
rect 1873 3384 1885 3424
rect 1907 3384 1919 3424
rect 1927 3384 1939 3464
rect 1957 3384 1969 3464
rect 1987 3384 2009 3464
rect 2027 3384 2039 3464
rect 2077 3384 2089 3424
rect 2097 3384 2109 3424
rect 2117 3384 2129 3424
rect 2171 3384 2183 3464
rect 2191 3384 2203 3464
rect 2211 3384 2223 3452
rect 2231 3384 2243 3456
rect 2271 3384 2283 3424
rect 2291 3384 2303 3420
rect 2311 3384 2323 3424
rect 2331 3384 2343 3424
rect 2371 3384 2383 3424
rect 2391 3384 2403 3424
rect 2431 3384 2443 3424
rect 2451 3384 2463 3420
rect 2471 3384 2483 3424
rect 2491 3384 2503 3424
rect 2531 3384 2543 3424
rect 2551 3384 2563 3420
rect 2571 3384 2583 3424
rect 2591 3384 2603 3424
rect 2636 3384 2648 3424
rect 2658 3384 2670 3464
rect 2686 3384 2698 3464
rect 2722 3384 2734 3464
rect 2750 3384 2762 3464
rect 2772 3384 2784 3424
rect 2817 3384 2829 3424
rect 2837 3384 2849 3424
rect 2857 3384 2869 3424
rect 2902 3384 2914 3464
rect 2930 3384 2942 3464
rect 2952 3384 2964 3424
rect 2997 3384 3009 3464
rect 3025 3384 3037 3464
rect 3096 3384 3108 3424
rect 3118 3384 3130 3464
rect 3146 3384 3158 3464
rect 3177 3384 3189 3462
rect 3197 3384 3209 3450
rect 3217 3384 3229 3462
rect 3237 3396 3249 3464
rect 3257 3384 3269 3464
rect 3297 3384 3309 3424
rect 3317 3384 3329 3424
rect 3337 3384 3349 3424
rect 3377 3384 3389 3424
rect 3397 3384 3409 3424
rect 3417 3384 3429 3424
rect 3457 3384 3469 3424
rect 3477 3384 3489 3424
rect 3497 3384 3509 3424
rect 3537 3384 3549 3464
rect 3565 3384 3577 3464
rect 3617 3384 3629 3424
rect 3637 3384 3649 3424
rect 3657 3384 3669 3424
rect 3697 3384 3709 3424
rect 3717 3384 3729 3424
rect 3737 3384 3749 3424
rect 3791 3384 3803 3424
rect 3811 3384 3823 3424
rect 3831 3384 3843 3424
rect 3883 3384 3895 3464
rect 3911 3384 3923 3464
rect 3937 3384 3949 3424
rect 3957 3384 3969 3424
rect 3977 3384 3989 3424
rect 4017 3384 4029 3424
rect 4037 3384 4049 3424
rect 4057 3384 4069 3424
rect 4102 3384 4114 3464
rect 4130 3384 4142 3464
rect 4152 3384 4164 3424
rect 4211 3384 4223 3424
rect 4231 3384 4243 3420
rect 4251 3384 4263 3424
rect 4271 3384 4283 3424
rect 4297 3384 4309 3424
rect 4317 3384 4329 3424
rect 4337 3384 4349 3420
rect 4357 3384 4369 3424
rect 4397 3384 4409 3456
rect 4417 3384 4429 3452
rect 4437 3384 4449 3464
rect 4457 3384 4469 3464
rect 4497 3384 4509 3424
rect 4517 3384 4529 3424
rect 4571 3384 4583 3424
rect 4591 3384 4603 3420
rect 4611 3384 4623 3424
rect 4631 3384 4643 3424
rect 4657 3384 4669 3424
rect 4677 3384 4689 3424
rect 4697 3384 4709 3420
rect 4717 3384 4729 3424
rect 21 3276 33 3356
rect 41 3316 53 3356
rect 75 3316 87 3356
rect 107 3316 119 3356
rect 127 3316 139 3356
rect 153 3316 165 3356
rect 181 3336 193 3356
rect 211 3336 223 3356
rect 231 3276 243 3356
rect 271 3276 283 3356
rect 291 3276 303 3344
rect 311 3278 323 3356
rect 331 3290 343 3356
rect 351 3278 363 3356
rect 377 3316 389 3356
rect 397 3316 409 3356
rect 417 3316 429 3356
rect 462 3276 474 3356
rect 490 3276 502 3356
rect 512 3316 524 3356
rect 562 3276 574 3356
rect 590 3276 602 3356
rect 612 3316 624 3356
rect 671 3316 683 3356
rect 691 3316 703 3356
rect 711 3316 723 3356
rect 737 3316 749 3356
rect 757 3316 769 3356
rect 811 3276 823 3356
rect 831 3276 843 3356
rect 851 3276 863 3356
rect 871 3276 883 3356
rect 891 3276 903 3356
rect 911 3276 923 3356
rect 931 3276 943 3356
rect 951 3276 963 3356
rect 971 3276 983 3356
rect 997 3276 1009 3356
rect 1017 3276 1029 3356
rect 1037 3276 1049 3356
rect 1057 3276 1069 3356
rect 1077 3276 1089 3356
rect 1097 3276 1109 3356
rect 1117 3276 1129 3356
rect 1137 3276 1149 3356
rect 1157 3276 1169 3356
rect 1211 3316 1223 3356
rect 1231 3316 1243 3356
rect 1257 3276 1269 3356
rect 1277 3336 1289 3356
rect 1307 3336 1319 3356
rect 1335 3316 1347 3356
rect 1361 3316 1373 3356
rect 1381 3316 1393 3356
rect 1413 3316 1425 3356
rect 1447 3316 1459 3356
rect 1467 3276 1479 3356
rect 1502 3276 1514 3356
rect 1530 3276 1542 3356
rect 1552 3316 1564 3356
rect 1616 3316 1628 3356
rect 1638 3276 1650 3356
rect 1666 3276 1678 3356
rect 1716 3316 1728 3356
rect 1738 3276 1750 3356
rect 1766 3276 1778 3356
rect 1811 3316 1823 3356
rect 1831 3316 1843 3356
rect 1876 3316 1888 3356
rect 1898 3276 1910 3356
rect 1926 3276 1938 3356
rect 1976 3316 1988 3356
rect 1998 3276 2010 3356
rect 2026 3276 2038 3356
rect 2057 3276 2069 3356
rect 2077 3336 2089 3356
rect 2107 3336 2119 3356
rect 2135 3316 2147 3356
rect 2161 3316 2173 3356
rect 2181 3316 2193 3356
rect 2213 3316 2225 3356
rect 2247 3316 2259 3356
rect 2267 3276 2279 3356
rect 2311 3316 2323 3356
rect 2331 3316 2343 3356
rect 2371 3316 2383 3356
rect 2391 3316 2403 3356
rect 2431 3316 2443 3356
rect 2451 3320 2463 3356
rect 2471 3316 2483 3356
rect 2491 3316 2503 3356
rect 2517 3284 2529 3356
rect 2537 3288 2549 3356
rect 2557 3276 2569 3356
rect 2577 3276 2589 3356
rect 2631 3316 2643 3356
rect 2651 3316 2663 3356
rect 2696 3316 2708 3356
rect 2718 3276 2730 3356
rect 2746 3276 2758 3356
rect 2777 3276 2789 3356
rect 2805 3276 2817 3356
rect 2862 3276 2874 3356
rect 2890 3276 2902 3356
rect 2912 3316 2924 3356
rect 2957 3316 2969 3356
rect 2977 3316 2989 3356
rect 2997 3316 3009 3356
rect 3037 3316 3049 3356
rect 3057 3316 3069 3356
rect 3077 3316 3089 3356
rect 3131 3276 3143 3356
rect 3151 3276 3163 3356
rect 3171 3288 3183 3356
rect 3191 3284 3203 3356
rect 3231 3316 3243 3356
rect 3251 3320 3263 3356
rect 3271 3316 3283 3356
rect 3291 3316 3303 3356
rect 3336 3316 3348 3356
rect 3358 3276 3370 3356
rect 3386 3276 3398 3356
rect 3427 3276 3439 3356
rect 3447 3276 3459 3356
rect 3471 3316 3483 3356
rect 3491 3316 3503 3356
rect 3517 3316 3529 3356
rect 3537 3316 3549 3356
rect 3557 3316 3569 3356
rect 3607 3276 3619 3356
rect 3627 3276 3639 3356
rect 3651 3316 3663 3356
rect 3671 3316 3683 3356
rect 3711 3276 3723 3356
rect 3731 3276 3743 3344
rect 3751 3278 3763 3356
rect 3771 3290 3783 3356
rect 3791 3278 3803 3356
rect 3831 3316 3843 3356
rect 3851 3316 3863 3356
rect 3871 3316 3883 3356
rect 3902 3276 3914 3356
rect 3930 3276 3942 3356
rect 3952 3316 3964 3356
rect 3997 3316 4009 3356
rect 4017 3316 4029 3356
rect 4037 3316 4049 3356
rect 4087 3276 4099 3356
rect 4107 3276 4119 3356
rect 4131 3316 4143 3356
rect 4151 3316 4163 3356
rect 4177 3316 4189 3356
rect 4197 3316 4209 3356
rect 4217 3316 4229 3356
rect 4257 3316 4269 3356
rect 4277 3316 4289 3356
rect 4301 3276 4313 3356
rect 4321 3276 4333 3356
rect 4357 3284 4369 3356
rect 4377 3288 4389 3356
rect 4397 3276 4409 3356
rect 4417 3276 4429 3356
rect 4462 3276 4474 3356
rect 4490 3276 4502 3356
rect 4512 3316 4524 3356
rect 4562 3276 4574 3356
rect 4590 3276 4602 3356
rect 4612 3316 4624 3356
rect 4671 3316 4683 3356
rect 4691 3320 4703 3356
rect 4711 3316 4723 3356
rect 4731 3316 4743 3356
rect 21 2904 33 2984
rect 41 2904 53 2944
rect 75 2904 87 2944
rect 107 2904 119 2944
rect 127 2904 139 2944
rect 153 2904 165 2944
rect 181 2904 193 2924
rect 211 2904 223 2924
rect 231 2904 243 2984
rect 276 2904 288 2944
rect 298 2904 310 2984
rect 326 2904 338 2984
rect 371 2904 383 2944
rect 391 2904 403 2944
rect 411 2904 423 2944
rect 437 2904 449 2984
rect 457 2904 469 2924
rect 487 2904 499 2924
rect 515 2904 527 2944
rect 541 2904 553 2944
rect 561 2904 573 2944
rect 593 2904 605 2944
rect 627 2904 639 2944
rect 647 2904 659 2984
rect 681 2904 693 2984
rect 701 2904 713 2944
rect 735 2904 747 2944
rect 767 2904 779 2944
rect 787 2904 799 2944
rect 813 2904 825 2944
rect 841 2904 853 2924
rect 871 2904 883 2924
rect 891 2904 903 2984
rect 917 2904 929 2944
rect 937 2904 949 2944
rect 1003 2904 1015 2984
rect 1031 2904 1043 2984
rect 1071 2904 1083 2944
rect 1091 2904 1103 2944
rect 1111 2904 1123 2944
rect 1142 2904 1154 2984
rect 1170 2904 1182 2984
rect 1192 2904 1204 2944
rect 1237 2904 1249 2976
rect 1257 2904 1269 2972
rect 1277 2904 1289 2984
rect 1297 2904 1309 2984
rect 1341 2904 1353 2984
rect 1361 2904 1373 2944
rect 1395 2904 1407 2944
rect 1427 2904 1439 2944
rect 1447 2904 1459 2944
rect 1473 2904 1485 2944
rect 1501 2904 1513 2924
rect 1531 2904 1543 2924
rect 1551 2904 1563 2984
rect 1603 2904 1615 2984
rect 1631 2904 1643 2984
rect 1671 2904 1683 2944
rect 1691 2904 1703 2944
rect 1711 2904 1723 2944
rect 1742 2904 1754 2984
rect 1770 2904 1782 2984
rect 1792 2904 1804 2944
rect 1856 2904 1868 2944
rect 1878 2904 1890 2984
rect 1906 2904 1918 2984
rect 1937 2904 1949 2984
rect 1957 2904 1969 2924
rect 1987 2904 1999 2924
rect 2015 2904 2027 2944
rect 2041 2904 2053 2944
rect 2061 2904 2073 2944
rect 2093 2904 2105 2944
rect 2127 2904 2139 2944
rect 2147 2904 2159 2984
rect 2203 2904 2215 2984
rect 2231 2904 2243 2984
rect 2271 2904 2283 2944
rect 2291 2904 2303 2944
rect 2331 2904 2343 2944
rect 2351 2904 2363 2940
rect 2371 2904 2383 2944
rect 2391 2904 2403 2944
rect 2431 2904 2443 2984
rect 2451 2904 2463 2984
rect 2471 2904 2483 2972
rect 2491 2904 2503 2976
rect 2531 2904 2543 2944
rect 2551 2904 2563 2940
rect 2571 2904 2583 2944
rect 2591 2904 2603 2944
rect 2636 2904 2648 2944
rect 2658 2904 2670 2984
rect 2686 2904 2698 2984
rect 2743 2904 2755 2984
rect 2771 2904 2783 2984
rect 2797 2904 2809 2944
rect 2817 2904 2829 2944
rect 2837 2904 2849 2944
rect 2877 2904 2889 2944
rect 2897 2904 2909 2944
rect 2917 2904 2929 2944
rect 2957 2904 2969 2982
rect 2977 2904 2989 2970
rect 2997 2904 3009 2982
rect 3017 2916 3029 2984
rect 3037 2904 3049 2984
rect 3077 2904 3089 2944
rect 3097 2904 3109 2944
rect 3117 2904 3129 2944
rect 3162 2904 3174 2984
rect 3190 2904 3202 2984
rect 3212 2904 3224 2944
rect 3257 2904 3269 2984
rect 3277 2904 3289 2984
rect 3317 2904 3329 2944
rect 3337 2904 3349 2944
rect 3361 2904 3373 2984
rect 3381 2904 3393 2984
rect 3429 2904 3441 2984
rect 3449 2904 3461 2984
rect 3471 2904 3483 2944
rect 3509 2904 3521 2984
rect 3529 2904 3541 2984
rect 3551 2904 3563 2944
rect 3577 2904 3589 2944
rect 3597 2904 3609 2944
rect 3617 2904 3629 2944
rect 3662 2904 3674 2984
rect 3690 2904 3702 2984
rect 3712 2904 3724 2944
rect 3769 2904 3781 2984
rect 3789 2904 3801 2984
rect 3811 2904 3823 2944
rect 3842 2904 3854 2984
rect 3870 2904 3882 2984
rect 3892 2904 3904 2944
rect 3937 2904 3949 2944
rect 3957 2904 3969 2944
rect 3977 2904 3989 2940
rect 3997 2904 4009 2944
rect 4037 2904 4049 2944
rect 4059 2904 4071 2984
rect 4079 2904 4091 2984
rect 4131 2904 4143 2984
rect 4151 2904 4163 2984
rect 4171 2904 4183 2972
rect 4191 2904 4203 2976
rect 4217 2904 4229 2944
rect 4237 2904 4249 2944
rect 4257 2904 4269 2940
rect 4277 2904 4289 2944
rect 4331 2904 4343 2984
rect 4351 2904 4363 2984
rect 4371 2904 4383 2972
rect 4391 2904 4403 2976
rect 4431 2904 4443 2944
rect 4451 2904 4463 2940
rect 4471 2904 4483 2944
rect 4491 2904 4503 2944
rect 4531 2904 4543 2944
rect 4551 2904 4563 2944
rect 4596 2904 4608 2944
rect 4618 2904 4630 2984
rect 4646 2904 4658 2984
rect 4682 2904 4694 2984
rect 4710 2904 4722 2984
rect 4732 2904 4744 2944
rect 21 2796 33 2876
rect 41 2836 53 2876
rect 75 2836 87 2876
rect 107 2836 119 2876
rect 127 2836 139 2876
rect 153 2836 165 2876
rect 181 2856 193 2876
rect 211 2856 223 2876
rect 231 2796 243 2876
rect 271 2796 283 2876
rect 291 2796 303 2864
rect 311 2798 323 2876
rect 331 2810 343 2876
rect 351 2798 363 2876
rect 377 2836 389 2876
rect 397 2836 409 2876
rect 417 2836 429 2876
rect 476 2836 488 2876
rect 498 2796 510 2876
rect 526 2796 538 2876
rect 569 2796 581 2876
rect 589 2796 601 2876
rect 611 2836 623 2876
rect 637 2836 649 2876
rect 657 2836 669 2876
rect 677 2836 689 2876
rect 736 2836 748 2876
rect 758 2796 770 2876
rect 786 2796 798 2876
rect 843 2796 855 2876
rect 871 2796 883 2876
rect 911 2836 923 2876
rect 931 2836 943 2876
rect 951 2836 963 2876
rect 977 2836 989 2876
rect 997 2836 1009 2876
rect 1051 2836 1063 2876
rect 1071 2836 1083 2876
rect 1091 2836 1103 2876
rect 1117 2796 1129 2876
rect 1145 2796 1157 2876
rect 1209 2796 1221 2876
rect 1229 2796 1241 2876
rect 1251 2836 1263 2876
rect 1281 2796 1293 2876
rect 1301 2836 1313 2876
rect 1335 2836 1347 2876
rect 1367 2836 1379 2876
rect 1387 2836 1399 2876
rect 1413 2836 1425 2876
rect 1441 2856 1453 2876
rect 1471 2856 1483 2876
rect 1491 2796 1503 2876
rect 1517 2836 1529 2876
rect 1537 2836 1549 2876
rect 1557 2836 1569 2876
rect 1616 2836 1628 2876
rect 1638 2796 1650 2876
rect 1666 2796 1678 2876
rect 1716 2836 1728 2876
rect 1738 2796 1750 2876
rect 1766 2796 1778 2876
rect 1823 2796 1835 2876
rect 1851 2796 1863 2876
rect 1891 2796 1903 2876
rect 1911 2796 1923 2876
rect 1931 2808 1943 2876
rect 1951 2804 1963 2876
rect 1989 2796 2001 2876
rect 2009 2796 2021 2876
rect 2031 2836 2043 2876
rect 2071 2836 2083 2876
rect 2091 2840 2103 2876
rect 2111 2836 2123 2876
rect 2131 2836 2143 2876
rect 2157 2836 2169 2876
rect 2179 2796 2191 2876
rect 2199 2796 2211 2876
rect 2241 2796 2253 2876
rect 2261 2836 2273 2876
rect 2295 2836 2307 2876
rect 2327 2836 2339 2876
rect 2347 2836 2359 2876
rect 2373 2836 2385 2876
rect 2401 2856 2413 2876
rect 2431 2856 2443 2876
rect 2451 2796 2463 2876
rect 2496 2836 2508 2876
rect 2518 2796 2530 2876
rect 2546 2796 2558 2876
rect 2596 2836 2608 2876
rect 2618 2796 2630 2876
rect 2646 2796 2658 2876
rect 2682 2796 2694 2876
rect 2710 2796 2722 2876
rect 2732 2836 2744 2876
rect 2777 2836 2789 2876
rect 2797 2836 2809 2876
rect 2817 2836 2829 2876
rect 2857 2836 2869 2876
rect 2877 2836 2889 2876
rect 2897 2836 2909 2876
rect 2942 2796 2954 2876
rect 2970 2796 2982 2876
rect 2992 2836 3004 2876
rect 3042 2796 3054 2876
rect 3070 2796 3082 2876
rect 3092 2836 3104 2876
rect 3137 2836 3149 2876
rect 3157 2836 3169 2876
rect 3177 2836 3189 2876
rect 3236 2836 3248 2876
rect 3258 2796 3270 2876
rect 3286 2796 3298 2876
rect 3331 2836 3343 2876
rect 3351 2836 3363 2876
rect 3371 2836 3383 2876
rect 3397 2836 3409 2876
rect 3417 2836 3429 2876
rect 3437 2840 3449 2876
rect 3457 2836 3469 2876
rect 3516 2836 3528 2876
rect 3538 2796 3550 2876
rect 3566 2796 3578 2876
rect 3602 2796 3614 2876
rect 3630 2796 3642 2876
rect 3652 2836 3664 2876
rect 3711 2836 3723 2876
rect 3731 2836 3743 2876
rect 3751 2836 3763 2876
rect 3796 2836 3808 2876
rect 3818 2796 3830 2876
rect 3846 2796 3858 2876
rect 3877 2836 3889 2876
rect 3897 2836 3909 2876
rect 3917 2840 3929 2876
rect 3937 2836 3949 2876
rect 3977 2836 3989 2876
rect 3997 2836 4009 2876
rect 4051 2796 4063 2876
rect 4071 2796 4083 2864
rect 4091 2798 4103 2876
rect 4111 2810 4123 2876
rect 4131 2798 4143 2876
rect 4157 2836 4169 2876
rect 4177 2836 4189 2876
rect 4197 2840 4209 2876
rect 4217 2836 4229 2876
rect 4262 2796 4274 2876
rect 4290 2796 4302 2876
rect 4312 2836 4324 2876
rect 4357 2836 4369 2876
rect 4377 2836 4389 2876
rect 4401 2796 4413 2876
rect 4421 2796 4433 2876
rect 4457 2798 4469 2876
rect 4477 2810 4489 2876
rect 4497 2798 4509 2876
rect 4517 2796 4529 2864
rect 4537 2796 4549 2876
rect 4577 2836 4589 2876
rect 4597 2836 4609 2876
rect 4637 2804 4649 2876
rect 4657 2808 4669 2876
rect 4677 2796 4689 2876
rect 4697 2796 4709 2876
rect 21 2424 33 2504
rect 41 2424 53 2464
rect 75 2424 87 2464
rect 107 2424 119 2464
rect 127 2424 139 2464
rect 153 2424 165 2464
rect 181 2424 193 2444
rect 211 2424 223 2444
rect 231 2424 243 2504
rect 276 2424 288 2464
rect 298 2424 310 2504
rect 326 2424 338 2504
rect 357 2424 369 2464
rect 379 2424 391 2504
rect 399 2424 411 2504
rect 437 2424 449 2464
rect 457 2424 469 2464
rect 477 2424 489 2464
rect 536 2424 548 2464
rect 558 2424 570 2504
rect 586 2424 598 2504
rect 617 2424 629 2464
rect 639 2424 651 2504
rect 659 2424 671 2504
rect 716 2424 728 2464
rect 738 2424 750 2504
rect 766 2424 778 2504
rect 797 2424 809 2504
rect 825 2424 837 2504
rect 881 2424 893 2504
rect 901 2424 913 2464
rect 935 2424 947 2464
rect 967 2424 979 2464
rect 987 2424 999 2464
rect 1013 2424 1025 2464
rect 1041 2424 1053 2444
rect 1071 2424 1083 2444
rect 1091 2424 1103 2504
rect 1117 2424 1129 2464
rect 1137 2424 1149 2464
rect 1182 2424 1194 2504
rect 1210 2424 1222 2504
rect 1232 2424 1244 2464
rect 1277 2424 1289 2464
rect 1297 2424 1309 2464
rect 1337 2424 1349 2464
rect 1357 2424 1369 2464
rect 1377 2424 1389 2464
rect 1417 2424 1429 2504
rect 1437 2424 1449 2444
rect 1467 2424 1479 2444
rect 1495 2424 1507 2464
rect 1521 2424 1533 2464
rect 1541 2424 1553 2464
rect 1573 2424 1585 2464
rect 1607 2424 1619 2464
rect 1627 2424 1639 2504
rect 1662 2424 1674 2504
rect 1690 2424 1702 2504
rect 1712 2424 1724 2464
rect 1757 2424 1769 2504
rect 1777 2424 1789 2444
rect 1807 2424 1819 2444
rect 1835 2424 1847 2464
rect 1861 2424 1873 2464
rect 1881 2424 1893 2464
rect 1913 2424 1925 2464
rect 1947 2424 1959 2464
rect 1967 2424 1979 2504
rect 1997 2424 2009 2504
rect 2017 2424 2029 2504
rect 2037 2424 2049 2504
rect 2057 2424 2069 2504
rect 2077 2424 2089 2504
rect 2097 2424 2109 2504
rect 2117 2424 2129 2504
rect 2137 2424 2149 2504
rect 2157 2424 2169 2504
rect 2201 2424 2213 2504
rect 2221 2424 2233 2464
rect 2255 2424 2267 2464
rect 2287 2424 2299 2464
rect 2307 2424 2319 2464
rect 2333 2424 2345 2464
rect 2361 2424 2373 2444
rect 2391 2424 2403 2444
rect 2411 2424 2423 2504
rect 2451 2424 2463 2464
rect 2471 2424 2483 2464
rect 2491 2424 2503 2464
rect 2517 2424 2529 2464
rect 2537 2424 2549 2464
rect 2596 2424 2608 2464
rect 2618 2424 2630 2504
rect 2646 2424 2658 2504
rect 2677 2424 2689 2464
rect 2697 2424 2709 2464
rect 2751 2424 2763 2464
rect 2771 2424 2783 2464
rect 2791 2424 2803 2464
rect 2836 2424 2848 2464
rect 2858 2424 2870 2504
rect 2886 2424 2898 2504
rect 2917 2424 2929 2464
rect 2937 2424 2949 2464
rect 2961 2424 2973 2504
rect 2981 2424 2993 2504
rect 3022 2424 3034 2504
rect 3050 2424 3062 2504
rect 3072 2424 3084 2464
rect 3131 2424 3143 2464
rect 3151 2424 3163 2464
rect 3171 2424 3183 2464
rect 3197 2424 3209 2464
rect 3217 2424 3229 2464
rect 3241 2424 3253 2504
rect 3261 2424 3273 2504
rect 3311 2424 3323 2464
rect 3331 2424 3343 2460
rect 3351 2424 3363 2464
rect 3371 2424 3383 2464
rect 3397 2424 3409 2464
rect 3417 2424 3429 2464
rect 3457 2424 3469 2464
rect 3477 2424 3489 2464
rect 3497 2424 3509 2464
rect 3537 2424 3549 2464
rect 3557 2424 3569 2464
rect 3581 2424 3593 2504
rect 3601 2424 3613 2504
rect 3637 2424 3649 2464
rect 3659 2424 3671 2504
rect 3679 2424 3691 2504
rect 3717 2424 3729 2464
rect 3737 2424 3749 2464
rect 3787 2424 3799 2504
rect 3807 2424 3819 2504
rect 3831 2424 3843 2464
rect 3851 2424 3863 2464
rect 3891 2424 3903 2504
rect 3911 2436 3923 2504
rect 3931 2424 3943 2502
rect 3951 2424 3963 2490
rect 3971 2424 3983 2502
rect 4011 2424 4023 2464
rect 4031 2424 4043 2464
rect 4051 2424 4063 2464
rect 4091 2424 4103 2464
rect 4111 2424 4123 2464
rect 4131 2424 4143 2464
rect 4162 2424 4174 2504
rect 4190 2424 4202 2504
rect 4212 2424 4224 2464
rect 4257 2424 4269 2464
rect 4277 2424 4289 2464
rect 4297 2424 4309 2464
rect 4351 2424 4363 2464
rect 4371 2424 4383 2460
rect 4391 2424 4403 2464
rect 4411 2424 4423 2464
rect 4451 2424 4463 2464
rect 4471 2424 4483 2460
rect 4491 2424 4503 2464
rect 4511 2424 4523 2464
rect 4537 2424 4549 2496
rect 4557 2424 4569 2492
rect 4577 2424 4589 2504
rect 4597 2424 4609 2504
rect 4651 2424 4663 2464
rect 4671 2424 4683 2460
rect 4691 2424 4703 2464
rect 4711 2424 4723 2464
rect 21 2316 33 2396
rect 41 2356 53 2396
rect 75 2356 87 2396
rect 107 2356 119 2396
rect 127 2356 139 2396
rect 153 2356 165 2396
rect 181 2376 193 2396
rect 211 2376 223 2396
rect 231 2316 243 2396
rect 262 2316 274 2396
rect 290 2316 302 2396
rect 312 2356 324 2396
rect 357 2318 369 2396
rect 377 2330 389 2396
rect 397 2318 409 2396
rect 417 2316 429 2384
rect 437 2316 449 2396
rect 477 2356 489 2396
rect 499 2316 511 2396
rect 519 2316 531 2396
rect 557 2356 569 2396
rect 577 2356 589 2396
rect 597 2356 609 2396
rect 651 2356 663 2396
rect 671 2356 683 2396
rect 697 2316 709 2396
rect 725 2316 737 2396
rect 791 2316 803 2396
rect 811 2316 823 2396
rect 831 2328 843 2396
rect 851 2324 863 2396
rect 877 2316 889 2396
rect 905 2316 917 2396
rect 957 2316 969 2396
rect 985 2316 997 2396
rect 1037 2356 1049 2396
rect 1057 2356 1069 2396
rect 1097 2316 1109 2396
rect 1117 2376 1129 2396
rect 1147 2376 1159 2396
rect 1175 2356 1187 2396
rect 1201 2356 1213 2396
rect 1221 2356 1233 2396
rect 1253 2356 1265 2396
rect 1287 2356 1299 2396
rect 1307 2316 1319 2396
rect 1342 2316 1354 2396
rect 1370 2316 1382 2396
rect 1392 2356 1404 2396
rect 1437 2316 1449 2396
rect 1457 2376 1469 2396
rect 1487 2376 1499 2396
rect 1515 2356 1527 2396
rect 1541 2356 1553 2396
rect 1561 2356 1573 2396
rect 1593 2356 1605 2396
rect 1627 2356 1639 2396
rect 1647 2316 1659 2396
rect 1703 2316 1715 2396
rect 1731 2316 1743 2396
rect 1771 2316 1783 2396
rect 1791 2316 1803 2396
rect 1811 2328 1823 2396
rect 1831 2324 1843 2396
rect 1857 2316 1869 2396
rect 1877 2316 1889 2396
rect 1943 2316 1955 2396
rect 1971 2316 1983 2396
rect 1997 2316 2009 2396
rect 2017 2316 2029 2396
rect 2037 2316 2049 2396
rect 2057 2316 2069 2396
rect 2077 2316 2089 2396
rect 2097 2316 2109 2396
rect 2117 2316 2129 2396
rect 2137 2316 2149 2396
rect 2157 2316 2169 2396
rect 2202 2316 2214 2396
rect 2230 2316 2242 2396
rect 2252 2356 2264 2396
rect 2301 2316 2313 2396
rect 2321 2356 2333 2396
rect 2355 2356 2367 2396
rect 2387 2356 2399 2396
rect 2407 2356 2419 2396
rect 2433 2356 2445 2396
rect 2461 2376 2473 2396
rect 2491 2376 2503 2396
rect 2511 2316 2523 2396
rect 2551 2356 2563 2396
rect 2571 2356 2583 2396
rect 2591 2356 2603 2396
rect 2617 2356 2629 2396
rect 2637 2356 2649 2396
rect 2657 2356 2669 2396
rect 2697 2356 2709 2396
rect 2717 2356 2729 2396
rect 2737 2356 2749 2396
rect 2796 2356 2808 2396
rect 2818 2316 2830 2396
rect 2846 2316 2858 2396
rect 2896 2356 2908 2396
rect 2918 2316 2930 2396
rect 2946 2316 2958 2396
rect 2981 2316 2993 2396
rect 3001 2356 3013 2396
rect 3035 2356 3047 2396
rect 3067 2356 3079 2396
rect 3087 2356 3099 2396
rect 3113 2356 3125 2396
rect 3141 2376 3153 2396
rect 3171 2376 3183 2396
rect 3191 2316 3203 2396
rect 3222 2316 3234 2396
rect 3250 2316 3262 2396
rect 3272 2356 3284 2396
rect 3317 2356 3329 2396
rect 3337 2356 3349 2396
rect 3357 2356 3369 2396
rect 3397 2356 3409 2396
rect 3417 2356 3429 2396
rect 3437 2356 3449 2396
rect 3491 2356 3503 2396
rect 3511 2356 3523 2396
rect 3531 2356 3543 2396
rect 3571 2316 3583 2396
rect 3591 2316 3603 2396
rect 3631 2316 3643 2396
rect 3651 2316 3663 2396
rect 3691 2356 3703 2396
rect 3711 2356 3723 2396
rect 3742 2316 3754 2396
rect 3770 2316 3782 2396
rect 3792 2356 3804 2396
rect 3849 2316 3861 2396
rect 3869 2316 3881 2396
rect 3891 2356 3903 2396
rect 3917 2316 3929 2396
rect 3937 2316 3949 2396
rect 3977 2356 3989 2396
rect 3997 2356 4009 2396
rect 4021 2316 4033 2396
rect 4041 2316 4053 2396
rect 4096 2356 4108 2396
rect 4118 2316 4130 2396
rect 4146 2316 4158 2396
rect 4191 2356 4203 2396
rect 4211 2360 4223 2396
rect 4231 2356 4243 2396
rect 4251 2356 4263 2396
rect 4277 2324 4289 2396
rect 4297 2328 4309 2396
rect 4317 2316 4329 2396
rect 4337 2316 4349 2396
rect 4396 2356 4408 2396
rect 4418 2316 4430 2396
rect 4446 2316 4458 2396
rect 4482 2316 4494 2396
rect 4510 2316 4522 2396
rect 4532 2356 4544 2396
rect 4596 2356 4608 2396
rect 4618 2316 4630 2396
rect 4646 2316 4658 2396
rect 4677 2324 4689 2396
rect 4697 2328 4709 2396
rect 4717 2316 4729 2396
rect 4737 2316 4749 2396
rect 17 1944 29 2024
rect 37 1944 49 2024
rect 57 1944 69 2024
rect 77 1944 89 2024
rect 97 1944 109 2024
rect 117 1944 129 2024
rect 137 1944 149 2024
rect 157 1944 169 2024
rect 177 1944 189 2024
rect 231 1944 243 1984
rect 251 1944 263 1984
rect 271 1944 283 1984
rect 316 1944 328 1984
rect 338 1944 350 2024
rect 366 1944 378 2024
rect 397 1944 409 2022
rect 417 1944 429 2010
rect 437 1944 449 2022
rect 457 1956 469 2024
rect 477 1944 489 2024
rect 521 1944 533 2024
rect 541 1944 553 1984
rect 575 1944 587 1984
rect 607 1944 619 1984
rect 627 1944 639 1984
rect 653 1944 665 1984
rect 681 1944 693 1964
rect 711 1944 723 1964
rect 731 1944 743 2024
rect 771 1944 783 1984
rect 791 1944 803 1984
rect 811 1944 823 1984
rect 861 1944 873 2023
rect 881 1944 893 2023
rect 911 1944 923 2024
rect 937 1944 949 1984
rect 957 1944 969 1984
rect 977 1944 989 1984
rect 1017 1944 1029 2024
rect 1045 1944 1057 2024
rect 1102 1944 1114 2024
rect 1130 1944 1142 2024
rect 1152 1944 1164 1984
rect 1197 1944 1209 1984
rect 1217 1944 1229 1984
rect 1237 1944 1249 1984
rect 1277 1944 1289 2024
rect 1305 1944 1317 2024
rect 1357 1944 1369 2024
rect 1377 1944 1389 1964
rect 1407 1944 1419 1964
rect 1435 1944 1447 1984
rect 1461 1944 1473 1984
rect 1481 1944 1493 1984
rect 1513 1944 1525 1984
rect 1547 1944 1559 1984
rect 1567 1944 1579 2024
rect 1611 1944 1623 2024
rect 1631 1944 1643 2024
rect 1651 1944 1663 2012
rect 1671 1944 1683 2016
rect 1709 1944 1721 2024
rect 1729 1944 1741 2024
rect 1751 1944 1763 1984
rect 1777 1944 1789 2024
rect 1797 1944 1809 1964
rect 1827 1944 1839 1964
rect 1855 1944 1867 1984
rect 1881 1944 1893 1984
rect 1901 1944 1913 1984
rect 1933 1944 1945 1984
rect 1967 1944 1979 1984
rect 1987 1944 1999 2024
rect 2031 1944 2043 1984
rect 2051 1944 2063 1984
rect 2091 1944 2103 1984
rect 2111 1944 2123 1984
rect 2131 1944 2143 1984
rect 2157 1944 2169 1984
rect 2179 1944 2191 2024
rect 2199 1944 2211 2024
rect 2237 1944 2249 1984
rect 2257 1944 2269 1984
rect 2277 1944 2289 1984
rect 2336 1944 2348 1984
rect 2358 1944 2370 2024
rect 2386 1944 2398 2024
rect 2431 1944 2443 1984
rect 2451 1944 2463 1984
rect 2471 1944 2483 1984
rect 2511 1944 2523 1984
rect 2531 1944 2543 1984
rect 2551 1944 2563 1984
rect 2596 1944 2608 1984
rect 2618 1944 2630 2024
rect 2646 1944 2658 2024
rect 2696 1944 2708 1984
rect 2718 1944 2730 2024
rect 2746 1944 2758 2024
rect 2781 1944 2793 2024
rect 2801 1944 2813 1984
rect 2835 1944 2847 1984
rect 2867 1944 2879 1984
rect 2887 1944 2899 1984
rect 2913 1944 2925 1984
rect 2941 1944 2953 1964
rect 2971 1944 2983 1964
rect 2991 1944 3003 2024
rect 3017 1944 3029 1984
rect 3037 1944 3049 1984
rect 3061 1944 3073 2024
rect 3081 1944 3093 2024
rect 3136 1944 3148 1984
rect 3158 1944 3170 2024
rect 3186 1944 3198 2024
rect 3236 1944 3248 1984
rect 3258 1944 3270 2024
rect 3286 1944 3298 2024
rect 3317 1944 3329 1984
rect 3337 1944 3349 1984
rect 3357 1944 3369 1984
rect 3416 1944 3428 1984
rect 3438 1944 3450 2024
rect 3466 1944 3478 2024
rect 3497 1944 3509 1984
rect 3517 1944 3529 1984
rect 3537 1944 3549 1980
rect 3557 1944 3569 1984
rect 3597 1944 3609 1984
rect 3617 1944 3629 1984
rect 3657 1944 3669 1984
rect 3677 1944 3689 1984
rect 3697 1944 3709 1980
rect 3717 1944 3729 1984
rect 3757 1944 3769 1984
rect 3777 1944 3789 1984
rect 3797 1944 3809 1984
rect 3837 1944 3849 1984
rect 3859 1944 3871 2024
rect 3879 1944 3891 2024
rect 3922 1944 3934 2024
rect 3950 1944 3962 2024
rect 3972 1944 3984 1984
rect 4031 1944 4043 1984
rect 4051 1944 4063 1984
rect 4071 1944 4083 1984
rect 4111 1944 4123 1984
rect 4131 1944 4143 1984
rect 4151 1944 4163 1984
rect 4191 1944 4203 1984
rect 4211 1944 4223 1984
rect 4231 1944 4243 1984
rect 4257 1944 4269 1984
rect 4277 1944 4289 1984
rect 4301 1944 4313 2024
rect 4321 1944 4333 2024
rect 4357 1944 4369 2016
rect 4377 1944 4389 2012
rect 4397 1944 4409 2024
rect 4417 1944 4429 2024
rect 4471 1944 4483 2024
rect 4491 1944 4503 2024
rect 4511 1944 4523 2012
rect 4531 1944 4543 2016
rect 4557 1944 4569 1984
rect 4577 1944 4589 1984
rect 4597 1944 4609 1980
rect 4617 1944 4629 1984
rect 4657 1944 4669 1984
rect 4677 1944 4689 1984
rect 4697 1944 4709 1980
rect 4717 1944 4729 1984
rect 21 1836 33 1916
rect 41 1876 53 1916
rect 75 1876 87 1916
rect 107 1876 119 1916
rect 127 1876 139 1916
rect 153 1876 165 1916
rect 181 1896 193 1916
rect 211 1896 223 1916
rect 231 1836 243 1916
rect 262 1836 274 1916
rect 290 1836 302 1916
rect 312 1876 324 1916
rect 376 1876 388 1916
rect 398 1836 410 1916
rect 426 1836 438 1916
rect 476 1876 488 1916
rect 498 1836 510 1916
rect 526 1836 538 1916
rect 576 1876 588 1916
rect 598 1836 610 1916
rect 626 1836 638 1916
rect 657 1876 669 1916
rect 677 1876 689 1916
rect 717 1876 729 1916
rect 737 1876 749 1916
rect 803 1836 815 1916
rect 831 1836 843 1916
rect 857 1876 869 1916
rect 877 1876 889 1916
rect 897 1880 909 1916
rect 917 1876 929 1916
rect 961 1836 973 1916
rect 981 1876 993 1916
rect 1015 1876 1027 1916
rect 1047 1876 1059 1916
rect 1067 1876 1079 1916
rect 1093 1876 1105 1916
rect 1121 1896 1133 1916
rect 1151 1896 1163 1916
rect 1171 1836 1183 1916
rect 1197 1876 1209 1916
rect 1217 1876 1229 1916
rect 1237 1876 1249 1916
rect 1296 1876 1308 1916
rect 1318 1836 1330 1916
rect 1346 1836 1358 1916
rect 1391 1836 1403 1916
rect 1411 1836 1423 1916
rect 1431 1836 1443 1916
rect 1451 1836 1463 1916
rect 1471 1836 1483 1916
rect 1491 1836 1503 1916
rect 1511 1836 1523 1916
rect 1531 1836 1543 1916
rect 1551 1836 1563 1916
rect 1581 1836 1593 1916
rect 1601 1876 1613 1916
rect 1635 1876 1647 1916
rect 1667 1876 1679 1916
rect 1687 1876 1699 1916
rect 1713 1876 1725 1916
rect 1741 1896 1753 1916
rect 1771 1896 1783 1916
rect 1791 1836 1803 1916
rect 1831 1836 1843 1916
rect 1851 1836 1863 1916
rect 1871 1848 1883 1916
rect 1891 1844 1903 1916
rect 1917 1836 1929 1916
rect 1945 1836 1957 1916
rect 2011 1836 2023 1916
rect 2031 1836 2043 1916
rect 2051 1848 2063 1916
rect 2071 1844 2083 1916
rect 2123 1836 2135 1916
rect 2151 1836 2163 1916
rect 2177 1844 2189 1916
rect 2197 1848 2209 1916
rect 2217 1836 2229 1916
rect 2237 1836 2249 1916
rect 2277 1836 2289 1916
rect 2297 1896 2309 1916
rect 2327 1896 2339 1916
rect 2355 1876 2367 1916
rect 2381 1876 2393 1916
rect 2401 1876 2413 1916
rect 2433 1876 2445 1916
rect 2467 1876 2479 1916
rect 2487 1836 2499 1916
rect 2521 1836 2533 1916
rect 2541 1876 2553 1916
rect 2575 1876 2587 1916
rect 2607 1876 2619 1916
rect 2627 1876 2639 1916
rect 2653 1876 2665 1916
rect 2681 1896 2693 1916
rect 2711 1896 2723 1916
rect 2731 1836 2743 1916
rect 2761 1836 2773 1916
rect 2781 1876 2793 1916
rect 2815 1876 2827 1916
rect 2847 1876 2859 1916
rect 2867 1876 2879 1916
rect 2893 1876 2905 1916
rect 2921 1896 2933 1916
rect 2951 1896 2963 1916
rect 2971 1836 2983 1916
rect 3011 1836 3023 1916
rect 3031 1836 3043 1916
rect 3071 1876 3083 1916
rect 3091 1876 3103 1916
rect 3111 1876 3123 1916
rect 3151 1836 3163 1916
rect 3171 1836 3183 1916
rect 3197 1844 3209 1916
rect 3217 1848 3229 1916
rect 3237 1836 3249 1916
rect 3257 1836 3269 1916
rect 3297 1836 3309 1916
rect 3325 1836 3337 1916
rect 3387 1836 3399 1916
rect 3407 1836 3419 1916
rect 3431 1876 3443 1916
rect 3451 1876 3463 1916
rect 3477 1836 3489 1916
rect 3497 1836 3509 1916
rect 3551 1836 3563 1916
rect 3571 1836 3583 1904
rect 3591 1838 3603 1916
rect 3611 1850 3623 1916
rect 3631 1838 3643 1916
rect 3671 1836 3683 1916
rect 3691 1836 3703 1916
rect 3743 1836 3755 1916
rect 3771 1836 3783 1916
rect 3797 1876 3809 1916
rect 3819 1836 3831 1916
rect 3839 1836 3851 1916
rect 3877 1876 3889 1916
rect 3897 1876 3909 1916
rect 3921 1836 3933 1916
rect 3941 1836 3953 1916
rect 3991 1836 4003 1916
rect 4011 1836 4023 1904
rect 4031 1838 4043 1916
rect 4051 1850 4063 1916
rect 4071 1838 4083 1916
rect 4097 1838 4109 1916
rect 4117 1850 4129 1916
rect 4137 1838 4149 1916
rect 4157 1836 4169 1904
rect 4177 1836 4189 1916
rect 4217 1876 4229 1916
rect 4237 1876 4249 1916
rect 4257 1876 4269 1916
rect 4297 1876 4309 1916
rect 4317 1876 4329 1916
rect 4341 1836 4353 1916
rect 4361 1836 4373 1916
rect 4397 1838 4409 1916
rect 4417 1850 4429 1916
rect 4437 1838 4449 1916
rect 4457 1836 4469 1904
rect 4477 1836 4489 1916
rect 4531 1876 4543 1916
rect 4551 1876 4563 1916
rect 4582 1836 4594 1916
rect 4610 1836 4622 1916
rect 4632 1876 4644 1916
rect 4677 1876 4689 1916
rect 4697 1876 4709 1916
rect 17 1464 29 1544
rect 37 1464 49 1544
rect 57 1464 69 1544
rect 77 1464 89 1544
rect 97 1464 109 1544
rect 117 1464 129 1544
rect 137 1464 149 1544
rect 157 1464 169 1544
rect 177 1464 189 1544
rect 243 1464 255 1544
rect 271 1464 283 1544
rect 309 1464 321 1544
rect 329 1464 341 1544
rect 351 1464 363 1504
rect 381 1464 393 1544
rect 401 1464 413 1504
rect 435 1464 447 1504
rect 467 1464 479 1504
rect 487 1464 499 1504
rect 513 1464 525 1504
rect 541 1464 553 1484
rect 571 1464 583 1484
rect 591 1464 603 1544
rect 621 1464 633 1544
rect 641 1464 653 1504
rect 675 1464 687 1504
rect 707 1464 719 1504
rect 727 1464 739 1504
rect 753 1464 765 1504
rect 781 1464 793 1484
rect 811 1464 823 1484
rect 831 1464 843 1544
rect 857 1464 869 1544
rect 877 1464 889 1484
rect 907 1464 919 1484
rect 935 1464 947 1504
rect 961 1464 973 1504
rect 981 1464 993 1504
rect 1013 1464 1025 1504
rect 1047 1464 1059 1504
rect 1067 1464 1079 1544
rect 1111 1464 1123 1504
rect 1131 1464 1143 1504
rect 1151 1464 1163 1504
rect 1196 1464 1208 1504
rect 1218 1464 1230 1544
rect 1246 1464 1258 1544
rect 1277 1464 1289 1544
rect 1297 1464 1309 1484
rect 1327 1464 1339 1484
rect 1355 1464 1367 1504
rect 1381 1464 1393 1504
rect 1401 1464 1413 1504
rect 1433 1464 1445 1504
rect 1467 1464 1479 1504
rect 1487 1464 1499 1544
rect 1521 1464 1533 1544
rect 1541 1464 1553 1504
rect 1575 1464 1587 1504
rect 1607 1464 1619 1504
rect 1627 1464 1639 1504
rect 1653 1464 1665 1504
rect 1681 1464 1693 1484
rect 1711 1464 1723 1484
rect 1731 1464 1743 1544
rect 1771 1464 1783 1544
rect 1791 1464 1803 1544
rect 1811 1464 1823 1532
rect 1831 1464 1843 1536
rect 1857 1464 1869 1544
rect 1885 1464 1897 1544
rect 1941 1464 1953 1544
rect 1961 1464 1973 1504
rect 1995 1464 2007 1504
rect 2027 1464 2039 1504
rect 2047 1464 2059 1504
rect 2073 1464 2085 1504
rect 2101 1464 2113 1484
rect 2131 1464 2143 1484
rect 2151 1464 2163 1544
rect 2203 1464 2215 1544
rect 2231 1464 2243 1544
rect 2271 1464 2283 1504
rect 2291 1464 2303 1504
rect 2311 1464 2323 1504
rect 2342 1464 2354 1544
rect 2370 1464 2382 1544
rect 2392 1464 2404 1504
rect 2437 1464 2449 1544
rect 2457 1464 2469 1484
rect 2487 1464 2499 1484
rect 2515 1464 2527 1504
rect 2541 1464 2553 1504
rect 2561 1464 2573 1504
rect 2593 1464 2605 1504
rect 2627 1464 2639 1504
rect 2647 1464 2659 1544
rect 2681 1464 2693 1544
rect 2701 1464 2713 1504
rect 2735 1464 2747 1504
rect 2767 1464 2779 1504
rect 2787 1464 2799 1504
rect 2813 1464 2825 1504
rect 2841 1464 2853 1484
rect 2871 1464 2883 1484
rect 2891 1464 2903 1544
rect 2917 1464 2929 1544
rect 2937 1464 2949 1544
rect 2977 1464 2989 1504
rect 2997 1464 3009 1504
rect 3017 1464 3029 1504
rect 3071 1464 3083 1504
rect 3091 1464 3103 1504
rect 3111 1464 3123 1504
rect 3142 1464 3154 1544
rect 3170 1464 3182 1544
rect 3192 1464 3204 1504
rect 3237 1464 3249 1504
rect 3257 1464 3269 1504
rect 3277 1464 3289 1504
rect 3331 1464 3343 1504
rect 3351 1464 3363 1504
rect 3371 1464 3383 1504
rect 3416 1464 3428 1504
rect 3438 1464 3450 1544
rect 3466 1464 3478 1544
rect 3497 1464 3509 1504
rect 3517 1464 3529 1504
rect 3537 1464 3549 1500
rect 3557 1464 3569 1504
rect 3621 1464 3633 1544
rect 3651 1464 3673 1544
rect 3691 1464 3703 1544
rect 3717 1464 3729 1504
rect 3737 1464 3749 1504
rect 3777 1464 3789 1504
rect 3797 1464 3809 1504
rect 3817 1464 3829 1500
rect 3837 1464 3849 1504
rect 3877 1464 3889 1536
rect 3897 1464 3909 1532
rect 3917 1464 3929 1544
rect 3937 1464 3949 1544
rect 3982 1464 3994 1544
rect 4010 1464 4022 1544
rect 4032 1464 4044 1504
rect 4091 1464 4103 1504
rect 4111 1464 4123 1504
rect 4131 1464 4143 1504
rect 4157 1464 4169 1536
rect 4177 1464 4189 1532
rect 4197 1464 4209 1544
rect 4217 1464 4229 1544
rect 4262 1464 4274 1544
rect 4290 1464 4302 1544
rect 4312 1464 4324 1504
rect 4357 1464 4369 1504
rect 4377 1464 4389 1504
rect 4417 1464 4429 1544
rect 4445 1464 4457 1544
rect 4497 1464 4509 1504
rect 4517 1464 4529 1504
rect 4537 1464 4549 1504
rect 4577 1464 4589 1504
rect 4597 1464 4609 1504
rect 4617 1464 4629 1504
rect 4657 1464 4669 1504
rect 4677 1464 4689 1504
rect 4697 1464 4709 1504
rect 17 1356 29 1436
rect 37 1416 49 1436
rect 67 1416 79 1436
rect 95 1396 107 1436
rect 121 1396 133 1436
rect 141 1396 153 1436
rect 173 1396 185 1436
rect 207 1396 219 1436
rect 227 1356 239 1436
rect 261 1356 273 1436
rect 281 1396 293 1436
rect 315 1396 327 1436
rect 347 1396 359 1436
rect 367 1396 379 1436
rect 393 1396 405 1436
rect 421 1416 433 1436
rect 451 1416 463 1436
rect 471 1356 483 1436
rect 497 1396 509 1436
rect 517 1396 529 1436
rect 537 1396 549 1436
rect 596 1396 608 1436
rect 618 1356 630 1436
rect 646 1356 658 1436
rect 696 1396 708 1436
rect 718 1356 730 1436
rect 746 1356 758 1436
rect 789 1356 801 1436
rect 809 1356 821 1436
rect 831 1396 843 1436
rect 857 1396 869 1436
rect 877 1396 889 1436
rect 897 1396 909 1436
rect 956 1396 968 1436
rect 978 1356 990 1436
rect 1006 1356 1018 1436
rect 1051 1396 1063 1436
rect 1071 1396 1083 1436
rect 1097 1356 1109 1436
rect 1117 1356 1129 1436
rect 1137 1356 1149 1436
rect 1157 1356 1169 1436
rect 1177 1356 1189 1436
rect 1231 1396 1243 1436
rect 1251 1396 1263 1436
rect 1271 1396 1283 1436
rect 1316 1396 1328 1436
rect 1338 1356 1350 1436
rect 1366 1356 1378 1436
rect 1411 1396 1423 1436
rect 1431 1396 1443 1436
rect 1451 1396 1463 1436
rect 1496 1396 1508 1436
rect 1518 1356 1530 1436
rect 1546 1356 1558 1436
rect 1577 1396 1589 1436
rect 1599 1356 1611 1436
rect 1619 1356 1631 1436
rect 1657 1396 1669 1436
rect 1677 1396 1689 1436
rect 1697 1396 1709 1436
rect 1756 1396 1768 1436
rect 1778 1356 1790 1436
rect 1806 1356 1818 1436
rect 1837 1356 1849 1436
rect 1857 1416 1869 1436
rect 1887 1416 1899 1436
rect 1915 1396 1927 1436
rect 1941 1396 1953 1436
rect 1961 1396 1973 1436
rect 1993 1396 2005 1436
rect 2027 1396 2039 1436
rect 2047 1356 2059 1436
rect 2077 1396 2089 1436
rect 2097 1396 2109 1436
rect 2142 1356 2154 1436
rect 2170 1356 2182 1436
rect 2192 1396 2204 1436
rect 2251 1396 2263 1436
rect 2271 1396 2283 1436
rect 2291 1396 2303 1436
rect 2343 1356 2355 1436
rect 2371 1356 2383 1436
rect 2411 1396 2423 1436
rect 2431 1396 2443 1436
rect 2457 1356 2469 1436
rect 2485 1356 2497 1436
rect 2537 1356 2549 1436
rect 2557 1416 2569 1436
rect 2587 1416 2599 1436
rect 2615 1396 2627 1436
rect 2641 1396 2653 1436
rect 2661 1396 2673 1436
rect 2693 1396 2705 1436
rect 2727 1396 2739 1436
rect 2747 1356 2759 1436
rect 2777 1356 2789 1436
rect 2805 1356 2817 1436
rect 2871 1356 2883 1436
rect 2891 1356 2903 1436
rect 2922 1356 2934 1436
rect 2950 1356 2962 1436
rect 2972 1396 2984 1436
rect 3022 1356 3034 1436
rect 3050 1356 3062 1436
rect 3072 1396 3084 1436
rect 3122 1356 3134 1436
rect 3150 1356 3162 1436
rect 3172 1396 3184 1436
rect 3217 1396 3229 1436
rect 3237 1396 3249 1436
rect 3261 1356 3273 1436
rect 3281 1356 3293 1436
rect 3343 1356 3355 1436
rect 3371 1356 3383 1436
rect 3397 1396 3409 1436
rect 3417 1396 3429 1436
rect 3437 1400 3449 1436
rect 3457 1396 3469 1436
rect 3516 1396 3528 1436
rect 3538 1356 3550 1436
rect 3566 1356 3578 1436
rect 3602 1356 3614 1436
rect 3630 1356 3642 1436
rect 3652 1396 3664 1436
rect 3711 1396 3723 1436
rect 3731 1396 3743 1436
rect 3751 1396 3763 1436
rect 3791 1396 3803 1436
rect 3811 1396 3823 1436
rect 3831 1396 3843 1436
rect 3857 1396 3869 1436
rect 3877 1396 3889 1436
rect 3901 1356 3913 1436
rect 3921 1356 3933 1436
rect 3976 1396 3988 1436
rect 3998 1356 4010 1436
rect 4026 1356 4038 1436
rect 4057 1396 4069 1436
rect 4077 1396 4089 1436
rect 4131 1396 4143 1436
rect 4151 1396 4163 1436
rect 4171 1396 4183 1436
rect 4211 1396 4223 1436
rect 4231 1396 4243 1436
rect 4251 1396 4263 1436
rect 4303 1356 4315 1436
rect 4331 1356 4343 1436
rect 4376 1396 4388 1436
rect 4398 1356 4410 1436
rect 4426 1356 4438 1436
rect 4462 1356 4474 1436
rect 4490 1356 4502 1436
rect 4512 1396 4524 1436
rect 4571 1356 4583 1436
rect 4591 1356 4603 1436
rect 4611 1368 4623 1436
rect 4631 1364 4643 1436
rect 4657 1396 4669 1436
rect 4677 1396 4689 1436
rect 4697 1396 4709 1436
rect 17 984 29 1024
rect 37 984 49 1024
rect 91 984 103 1024
rect 111 984 123 1024
rect 131 984 143 1024
rect 176 984 188 1024
rect 198 984 210 1064
rect 226 984 238 1064
rect 257 984 269 1062
rect 277 984 289 1050
rect 297 984 309 1062
rect 317 996 329 1064
rect 337 984 349 1064
rect 391 984 403 1064
rect 411 984 423 1064
rect 431 984 443 1052
rect 451 984 463 1056
rect 501 984 513 1063
rect 521 984 533 1063
rect 551 984 563 1064
rect 577 984 589 1064
rect 605 984 617 1064
rect 667 984 679 1064
rect 687 984 699 1064
rect 711 984 723 1024
rect 731 984 743 1024
rect 769 984 781 1064
rect 789 984 801 1064
rect 811 984 823 1024
rect 863 984 875 1064
rect 891 984 903 1064
rect 931 984 943 1024
rect 951 984 963 1024
rect 991 984 1003 1024
rect 1011 984 1023 1024
rect 1037 984 1049 1064
rect 1065 984 1077 1064
rect 1117 984 1129 1024
rect 1137 984 1149 1024
rect 1203 984 1215 1064
rect 1231 984 1243 1064
rect 1257 984 1269 1056
rect 1277 984 1289 1052
rect 1297 984 1309 1064
rect 1317 984 1329 1064
rect 1361 984 1373 1064
rect 1381 984 1393 1024
rect 1415 984 1427 1024
rect 1447 984 1459 1024
rect 1467 984 1479 1024
rect 1493 984 1505 1024
rect 1521 984 1533 1004
rect 1551 984 1563 1004
rect 1571 984 1583 1064
rect 1611 984 1623 1024
rect 1631 984 1643 1024
rect 1657 984 1669 1024
rect 1677 984 1689 1024
rect 1697 984 1709 1024
rect 1737 984 1749 1064
rect 1765 984 1777 1064
rect 1821 984 1833 1064
rect 1841 984 1853 1024
rect 1875 984 1887 1024
rect 1907 984 1919 1024
rect 1927 984 1939 1024
rect 1953 984 1965 1024
rect 1981 984 1993 1004
rect 2011 984 2023 1004
rect 2031 984 2043 1064
rect 2071 984 2083 1024
rect 2091 984 2103 1024
rect 2117 984 2129 1064
rect 2145 984 2157 1064
rect 2197 984 2209 1064
rect 2225 984 2237 1064
rect 2291 984 2303 1024
rect 2311 984 2323 1024
rect 2337 984 2349 1064
rect 2357 984 2369 1004
rect 2387 984 2399 1004
rect 2415 984 2427 1024
rect 2441 984 2453 1024
rect 2461 984 2473 1024
rect 2493 984 2505 1024
rect 2527 984 2539 1024
rect 2547 984 2559 1064
rect 2577 984 2589 1024
rect 2597 984 2609 1024
rect 2642 984 2654 1064
rect 2670 984 2682 1064
rect 2692 984 2704 1024
rect 2737 984 2749 1064
rect 2767 984 2789 1064
rect 2807 984 2819 1064
rect 2857 984 2869 1064
rect 2885 984 2897 1064
rect 2951 984 2963 1024
rect 2971 984 2983 1024
rect 2991 984 3003 1024
rect 3017 984 3029 1024
rect 3037 984 3049 1024
rect 3061 984 3073 1064
rect 3081 984 3093 1064
rect 3122 984 3134 1064
rect 3150 984 3162 1064
rect 3172 984 3184 1024
rect 3217 984 3229 1064
rect 3247 984 3259 1063
rect 3267 984 3279 1063
rect 3331 984 3343 1024
rect 3351 984 3363 1024
rect 3371 984 3383 1024
rect 3411 984 3423 1024
rect 3431 984 3443 1024
rect 3451 984 3463 1024
rect 3477 984 3489 1024
rect 3497 984 3509 1024
rect 3517 984 3529 1024
rect 3557 984 3569 1024
rect 3577 984 3589 1024
rect 3597 984 3609 1024
rect 3642 984 3654 1064
rect 3670 984 3682 1064
rect 3692 984 3704 1024
rect 3751 984 3763 1024
rect 3771 984 3783 1020
rect 3791 984 3803 1024
rect 3811 984 3823 1024
rect 3837 984 3849 1056
rect 3857 984 3869 1052
rect 3877 984 3889 1064
rect 3897 984 3909 1064
rect 3951 984 3963 1024
rect 3971 984 3983 1024
rect 4011 984 4023 1024
rect 4031 984 4043 1020
rect 4051 984 4063 1024
rect 4071 984 4083 1024
rect 4097 984 4109 1056
rect 4117 984 4129 1052
rect 4137 984 4149 1064
rect 4157 984 4169 1064
rect 4197 984 4209 1024
rect 4217 984 4229 1024
rect 4271 984 4283 1064
rect 4291 984 4303 1064
rect 4311 984 4323 1052
rect 4331 984 4343 1056
rect 4376 984 4388 1024
rect 4398 984 4410 1064
rect 4426 984 4438 1064
rect 4462 984 4474 1064
rect 4490 984 4502 1064
rect 4512 984 4524 1024
rect 4557 984 4569 1064
rect 4585 984 4597 1064
rect 4651 984 4663 1024
rect 4671 984 4683 1024
rect 4691 984 4703 1024
rect 4731 984 4743 1024
rect 4751 984 4763 1024
rect 21 876 33 956
rect 41 916 53 956
rect 75 916 87 956
rect 107 916 119 956
rect 127 916 139 956
rect 153 916 165 956
rect 181 936 193 956
rect 211 936 223 956
rect 231 876 243 956
rect 257 916 269 956
rect 277 916 289 956
rect 297 916 309 956
rect 356 916 368 956
rect 378 876 390 956
rect 406 876 418 956
rect 441 876 453 956
rect 461 916 473 956
rect 495 916 507 956
rect 527 916 539 956
rect 547 916 559 956
rect 573 916 585 956
rect 601 936 613 956
rect 631 936 643 956
rect 651 876 663 956
rect 677 916 689 956
rect 697 916 709 956
rect 717 916 729 956
rect 776 916 788 956
rect 798 876 810 956
rect 826 876 838 956
rect 876 916 888 956
rect 898 876 910 956
rect 926 876 938 956
rect 971 916 983 956
rect 991 916 1003 956
rect 1043 876 1055 956
rect 1071 876 1083 956
rect 1097 876 1109 956
rect 1125 876 1137 956
rect 1191 916 1203 956
rect 1211 916 1223 956
rect 1231 916 1243 956
rect 1271 916 1283 956
rect 1291 916 1303 956
rect 1311 916 1323 956
rect 1351 916 1363 956
rect 1371 916 1383 956
rect 1391 916 1403 956
rect 1431 876 1443 956
rect 1451 876 1463 956
rect 1471 888 1483 956
rect 1491 884 1503 956
rect 1527 876 1539 956
rect 1547 876 1559 956
rect 1571 916 1583 956
rect 1591 916 1603 956
rect 1617 884 1629 956
rect 1637 888 1649 956
rect 1657 876 1669 956
rect 1677 876 1689 956
rect 1717 876 1729 956
rect 1737 876 1749 956
rect 1757 876 1769 956
rect 1777 876 1789 956
rect 1797 876 1809 956
rect 1817 876 1829 956
rect 1837 876 1849 956
rect 1857 876 1869 956
rect 1877 876 1889 956
rect 1931 916 1943 956
rect 1951 916 1963 956
rect 1971 916 1983 956
rect 2023 876 2035 956
rect 2051 876 2063 956
rect 2082 876 2094 956
rect 2110 876 2122 956
rect 2132 916 2144 956
rect 2182 876 2194 956
rect 2210 876 2222 956
rect 2232 916 2244 956
rect 2282 876 2294 956
rect 2310 876 2322 956
rect 2332 916 2344 956
rect 2377 916 2389 956
rect 2397 916 2409 956
rect 2417 916 2429 956
rect 2471 916 2483 956
rect 2491 916 2503 956
rect 2517 876 2529 956
rect 2537 936 2549 956
rect 2567 936 2579 956
rect 2595 916 2607 956
rect 2621 916 2633 956
rect 2641 916 2653 956
rect 2673 916 2685 956
rect 2707 916 2719 956
rect 2727 876 2739 956
rect 2776 916 2788 956
rect 2798 876 2810 956
rect 2826 876 2838 956
rect 2871 916 2883 956
rect 2891 916 2903 956
rect 2917 916 2929 956
rect 2937 916 2949 956
rect 2977 916 2989 956
rect 2997 916 3009 956
rect 3017 920 3029 956
rect 3037 916 3049 956
rect 3077 916 3089 956
rect 3097 916 3109 956
rect 3151 916 3163 956
rect 3171 916 3183 956
rect 3191 916 3203 956
rect 3217 876 3229 956
rect 3247 877 3259 956
rect 3267 877 3279 956
rect 3317 916 3329 956
rect 3337 916 3349 956
rect 3357 916 3369 956
rect 3397 916 3409 956
rect 3417 916 3429 956
rect 3437 916 3449 956
rect 3503 876 3515 956
rect 3531 876 3543 956
rect 3557 916 3569 956
rect 3577 916 3589 956
rect 3597 916 3609 956
rect 3651 916 3663 956
rect 3671 920 3683 956
rect 3691 916 3703 956
rect 3711 916 3723 956
rect 3751 916 3763 956
rect 3771 920 3783 956
rect 3791 916 3803 956
rect 3811 916 3823 956
rect 3837 916 3849 956
rect 3857 916 3869 956
rect 3877 916 3889 956
rect 3931 916 3943 956
rect 3951 920 3963 956
rect 3971 916 3983 956
rect 3991 916 4003 956
rect 4031 916 4043 956
rect 4051 916 4063 956
rect 4096 916 4108 956
rect 4118 876 4130 956
rect 4146 876 4158 956
rect 4196 916 4208 956
rect 4218 876 4230 956
rect 4246 876 4258 956
rect 4291 876 4303 956
rect 4311 876 4323 956
rect 4331 888 4343 956
rect 4351 884 4363 956
rect 4377 916 4389 956
rect 4397 916 4409 956
rect 4417 920 4429 956
rect 4437 916 4449 956
rect 4491 916 4503 956
rect 4511 920 4523 956
rect 4531 916 4543 956
rect 4551 916 4563 956
rect 4591 876 4603 956
rect 4611 876 4623 956
rect 4631 888 4643 956
rect 4651 884 4663 956
rect 4677 916 4689 956
rect 4697 916 4709 956
rect 4717 920 4729 956
rect 4737 916 4749 956
rect 21 504 33 584
rect 41 504 53 544
rect 75 504 87 544
rect 107 504 119 544
rect 127 504 139 544
rect 153 504 165 544
rect 181 504 193 524
rect 211 504 223 524
rect 231 504 243 584
rect 257 504 269 544
rect 277 504 289 544
rect 322 504 334 584
rect 350 504 362 584
rect 372 504 384 544
rect 417 504 429 544
rect 437 504 449 544
rect 457 504 469 544
rect 497 504 509 544
rect 519 504 531 584
rect 539 504 551 584
rect 591 504 603 544
rect 611 504 623 544
rect 637 504 649 584
rect 657 504 669 524
rect 687 504 699 524
rect 715 504 727 544
rect 741 504 753 544
rect 761 504 773 544
rect 793 504 805 544
rect 827 504 839 544
rect 847 504 859 584
rect 882 504 894 584
rect 910 504 922 584
rect 932 504 944 544
rect 1003 504 1015 584
rect 1031 504 1043 584
rect 1057 504 1069 584
rect 1087 504 1099 583
rect 1107 504 1119 583
rect 1176 504 1188 544
rect 1198 504 1210 584
rect 1226 504 1238 584
rect 1267 504 1279 584
rect 1287 504 1299 584
rect 1311 504 1323 544
rect 1331 504 1343 544
rect 1357 504 1369 584
rect 1385 504 1397 584
rect 1437 504 1449 544
rect 1459 504 1471 584
rect 1479 504 1491 584
rect 1521 504 1533 584
rect 1541 504 1553 544
rect 1575 504 1587 544
rect 1607 504 1619 544
rect 1627 504 1639 544
rect 1653 504 1665 544
rect 1681 504 1693 524
rect 1711 504 1723 524
rect 1731 504 1743 584
rect 1757 504 1769 544
rect 1779 504 1791 584
rect 1799 504 1811 584
rect 1863 504 1875 584
rect 1891 504 1903 584
rect 1943 504 1955 584
rect 1971 504 1983 584
rect 2011 504 2023 544
rect 2031 504 2043 544
rect 2057 504 2069 584
rect 2085 504 2097 584
rect 2137 504 2149 584
rect 2157 504 2169 524
rect 2187 504 2199 524
rect 2215 504 2227 544
rect 2241 504 2253 544
rect 2261 504 2273 544
rect 2293 504 2305 544
rect 2327 504 2339 544
rect 2347 504 2359 584
rect 2377 504 2389 582
rect 2397 504 2409 570
rect 2417 504 2429 582
rect 2437 516 2449 584
rect 2457 504 2469 584
rect 2521 504 2533 583
rect 2541 504 2553 583
rect 2571 504 2583 584
rect 2611 504 2623 584
rect 2631 504 2643 584
rect 2651 504 2663 572
rect 2671 504 2683 576
rect 2711 504 2723 584
rect 2731 504 2743 584
rect 2751 504 2763 572
rect 2771 504 2783 576
rect 2797 504 2809 544
rect 2817 504 2829 544
rect 2876 504 2888 544
rect 2898 504 2910 584
rect 2926 504 2938 584
rect 2962 504 2974 584
rect 2990 504 3002 584
rect 3012 504 3024 544
rect 3057 504 3069 544
rect 3077 504 3089 544
rect 3097 504 3109 544
rect 3151 504 3163 544
rect 3171 504 3183 544
rect 3197 504 3209 544
rect 3217 504 3229 544
rect 3271 504 3283 544
rect 3291 504 3303 540
rect 3311 504 3323 544
rect 3331 504 3343 544
rect 3383 504 3395 584
rect 3411 504 3423 584
rect 3442 504 3454 584
rect 3470 504 3482 584
rect 3492 504 3504 544
rect 3537 504 3549 576
rect 3557 504 3569 572
rect 3577 504 3589 584
rect 3597 504 3609 584
rect 3651 504 3663 584
rect 3671 504 3683 584
rect 3691 504 3703 572
rect 3711 504 3723 576
rect 3751 504 3763 584
rect 3771 516 3783 584
rect 3791 504 3803 582
rect 3811 504 3823 570
rect 3831 504 3843 582
rect 3871 504 3883 544
rect 3891 504 3903 540
rect 3911 504 3923 544
rect 3931 504 3943 544
rect 3971 504 3983 544
rect 3991 504 4003 540
rect 4011 504 4023 544
rect 4031 504 4043 544
rect 4057 504 4069 544
rect 4077 504 4089 544
rect 4117 504 4129 544
rect 4137 504 4149 544
rect 4157 504 4169 540
rect 4177 504 4189 544
rect 4217 504 4229 544
rect 4237 504 4249 544
rect 4257 504 4269 540
rect 4277 504 4289 544
rect 4331 504 4343 544
rect 4351 504 4363 540
rect 4371 504 4383 544
rect 4391 504 4403 544
rect 4431 504 4443 544
rect 4451 504 4463 540
rect 4471 504 4483 544
rect 4491 504 4503 544
rect 4517 504 4529 544
rect 4537 504 4549 544
rect 4596 504 4608 544
rect 4618 504 4630 584
rect 4646 504 4658 584
rect 4682 504 4694 584
rect 4710 504 4722 584
rect 4732 504 4744 544
rect 21 396 33 476
rect 41 436 53 476
rect 75 436 87 476
rect 107 436 119 476
rect 127 436 139 476
rect 153 436 165 476
rect 181 456 193 476
rect 211 456 223 476
rect 231 396 243 476
rect 257 436 269 476
rect 277 436 289 476
rect 297 436 309 476
rect 356 436 368 476
rect 378 396 390 476
rect 406 396 418 476
rect 437 436 449 476
rect 457 436 469 476
rect 497 436 509 476
rect 517 436 529 476
rect 537 436 549 476
rect 596 436 608 476
rect 618 396 630 476
rect 646 396 658 476
rect 682 396 694 476
rect 710 396 722 476
rect 732 436 744 476
rect 782 396 794 476
rect 810 396 822 476
rect 832 436 844 476
rect 896 436 908 476
rect 918 396 930 476
rect 946 396 958 476
rect 977 436 989 476
rect 997 436 1009 476
rect 1037 436 1049 476
rect 1057 436 1069 476
rect 1077 436 1089 476
rect 1131 396 1143 476
rect 1151 396 1163 476
rect 1171 408 1183 476
rect 1191 404 1203 476
rect 1231 436 1243 476
rect 1251 436 1263 476
rect 1296 436 1308 476
rect 1318 396 1330 476
rect 1346 396 1358 476
rect 1403 396 1415 476
rect 1431 396 1443 476
rect 1462 396 1474 476
rect 1490 396 1502 476
rect 1512 436 1524 476
rect 1557 436 1569 476
rect 1577 436 1589 476
rect 1597 436 1609 476
rect 1637 396 1649 476
rect 1657 456 1669 476
rect 1687 456 1699 476
rect 1715 436 1727 476
rect 1741 436 1753 476
rect 1761 436 1773 476
rect 1793 436 1805 476
rect 1827 436 1839 476
rect 1847 396 1859 476
rect 1891 436 1903 476
rect 1911 436 1923 476
rect 1931 436 1943 476
rect 1976 436 1988 476
rect 1998 396 2010 476
rect 2026 396 2038 476
rect 2061 396 2073 476
rect 2081 436 2093 476
rect 2115 436 2127 476
rect 2147 436 2159 476
rect 2167 436 2179 476
rect 2193 436 2205 476
rect 2221 456 2233 476
rect 2251 456 2263 476
rect 2271 396 2283 476
rect 2311 436 2323 476
rect 2331 436 2343 476
rect 2357 396 2369 476
rect 2385 396 2397 476
rect 2437 436 2449 476
rect 2457 436 2469 476
rect 2511 436 2523 476
rect 2531 436 2543 476
rect 2551 436 2563 476
rect 2577 396 2589 476
rect 2597 456 2609 476
rect 2627 456 2639 476
rect 2655 436 2667 476
rect 2681 436 2693 476
rect 2701 436 2713 476
rect 2733 436 2745 476
rect 2767 436 2779 476
rect 2787 396 2799 476
rect 2817 436 2829 476
rect 2837 436 2849 476
rect 2857 436 2869 476
rect 2897 398 2909 476
rect 2917 410 2929 476
rect 2937 398 2949 476
rect 2957 396 2969 464
rect 2977 396 2989 476
rect 3017 396 3029 476
rect 3045 396 3057 476
rect 3097 436 3109 476
rect 3117 436 3129 476
rect 3171 436 3183 476
rect 3191 440 3203 476
rect 3211 436 3223 476
rect 3231 436 3243 476
rect 3271 436 3283 476
rect 3291 440 3303 476
rect 3311 436 3323 476
rect 3331 436 3343 476
rect 3362 396 3374 476
rect 3390 396 3402 476
rect 3412 436 3424 476
rect 3471 436 3483 476
rect 3491 436 3503 476
rect 3517 436 3529 476
rect 3537 436 3549 476
rect 3557 436 3569 476
rect 3597 436 3609 476
rect 3617 436 3629 476
rect 3637 436 3649 476
rect 3682 396 3694 476
rect 3710 396 3722 476
rect 3732 436 3744 476
rect 3803 396 3815 476
rect 3831 396 3843 476
rect 3883 396 3895 476
rect 3911 396 3923 476
rect 3937 436 3949 476
rect 3957 436 3969 476
rect 3981 396 3993 476
rect 4001 396 4013 476
rect 4037 396 4049 476
rect 4065 396 4077 476
rect 4131 396 4143 476
rect 4151 396 4163 476
rect 4171 408 4183 476
rect 4191 404 4203 476
rect 4231 436 4243 476
rect 4251 440 4263 476
rect 4271 436 4283 476
rect 4291 436 4303 476
rect 4317 404 4329 476
rect 4337 408 4349 476
rect 4357 396 4369 476
rect 4377 396 4389 476
rect 4417 436 4429 476
rect 4437 436 4449 476
rect 4496 436 4508 476
rect 4518 396 4530 476
rect 4546 396 4558 476
rect 4577 436 4589 476
rect 4597 436 4609 476
rect 4637 436 4649 476
rect 4657 436 4669 476
rect 4697 436 4709 476
rect 4717 436 4729 476
rect 21 24 33 104
rect 41 24 53 64
rect 75 24 87 64
rect 107 24 119 64
rect 127 24 139 64
rect 153 24 165 64
rect 181 24 193 44
rect 211 24 223 44
rect 231 24 243 104
rect 257 24 269 102
rect 277 24 289 90
rect 297 24 309 102
rect 317 36 329 104
rect 337 24 349 104
rect 377 24 389 104
rect 405 24 417 104
rect 457 24 469 64
rect 477 24 489 64
rect 497 24 509 60
rect 517 24 529 64
rect 581 24 593 103
rect 601 24 613 103
rect 631 24 643 104
rect 671 24 683 104
rect 691 24 703 104
rect 711 24 723 92
rect 731 24 743 96
rect 757 24 769 104
rect 777 24 789 44
rect 807 24 819 44
rect 835 24 847 64
rect 861 24 873 64
rect 881 24 893 64
rect 913 24 925 64
rect 947 24 959 64
rect 967 24 979 104
rect 1016 24 1028 64
rect 1038 24 1050 104
rect 1066 24 1078 104
rect 1111 24 1123 64
rect 1131 24 1143 64
rect 1183 24 1195 104
rect 1211 24 1223 104
rect 1251 24 1263 64
rect 1271 24 1283 64
rect 1316 24 1328 64
rect 1338 24 1350 104
rect 1366 24 1378 104
rect 1411 24 1423 64
rect 1431 24 1443 64
rect 1471 24 1483 64
rect 1491 24 1503 64
rect 1517 24 1529 104
rect 1545 24 1557 104
rect 1611 24 1623 104
rect 1631 24 1643 104
rect 1651 24 1663 92
rect 1671 24 1683 96
rect 1701 24 1713 104
rect 1721 24 1733 64
rect 1755 24 1767 64
rect 1787 24 1799 64
rect 1807 24 1819 64
rect 1833 24 1845 64
rect 1861 24 1873 44
rect 1891 24 1903 44
rect 1911 24 1923 104
rect 1956 24 1968 64
rect 1978 24 1990 104
rect 2006 24 2018 104
rect 2037 24 2049 64
rect 2057 24 2069 64
rect 2097 24 2109 104
rect 2125 24 2137 104
rect 2177 24 2189 104
rect 2205 24 2217 104
rect 2283 24 2295 104
rect 2311 24 2323 104
rect 2337 24 2349 104
rect 2365 24 2377 104
rect 2431 24 2443 64
rect 2451 24 2463 64
rect 2477 24 2489 104
rect 2497 24 2509 44
rect 2527 24 2539 44
rect 2555 24 2567 64
rect 2581 24 2593 64
rect 2601 24 2613 64
rect 2633 24 2645 64
rect 2667 24 2679 64
rect 2687 24 2699 104
rect 2717 24 2729 104
rect 2737 24 2749 44
rect 2767 24 2779 44
rect 2795 24 2807 64
rect 2821 24 2833 64
rect 2841 24 2853 64
rect 2873 24 2885 64
rect 2907 24 2919 64
rect 2927 24 2939 104
rect 2957 24 2969 104
rect 2987 24 3009 104
rect 3027 24 3039 104
rect 3101 24 3113 103
rect 3121 24 3133 103
rect 3151 24 3163 104
rect 3182 24 3194 104
rect 3210 24 3222 104
rect 3232 24 3244 64
rect 3291 24 3303 64
rect 3311 24 3323 64
rect 3337 24 3349 64
rect 3357 24 3369 64
rect 3377 24 3389 64
rect 3431 24 3443 64
rect 3451 24 3463 60
rect 3471 24 3483 64
rect 3491 24 3503 64
rect 3531 24 3543 64
rect 3551 24 3563 64
rect 3591 24 3603 104
rect 3611 24 3623 104
rect 3631 24 3643 92
rect 3651 24 3663 96
rect 3703 24 3715 104
rect 3731 24 3743 104
rect 3757 24 3769 64
rect 3777 24 3789 64
rect 3822 24 3834 104
rect 3850 24 3862 104
rect 3872 24 3884 64
rect 3917 24 3929 104
rect 3945 24 3957 104
rect 4011 24 4023 64
rect 4031 24 4043 60
rect 4051 24 4063 64
rect 4071 24 4083 64
rect 4097 24 4109 64
rect 4117 24 4129 64
rect 4137 24 4149 64
rect 4191 24 4203 64
rect 4211 24 4223 60
rect 4231 24 4243 64
rect 4251 24 4263 64
rect 4291 24 4303 64
rect 4311 24 4323 64
rect 4331 24 4343 64
rect 4371 24 4383 64
rect 4391 24 4403 60
rect 4411 24 4423 64
rect 4431 24 4443 64
rect 4457 24 4469 64
rect 4477 24 4489 64
rect 4497 24 4509 64
rect 4537 24 4549 64
rect 4557 24 4569 64
rect 4577 24 4589 60
rect 4597 24 4609 64
rect 4651 24 4663 104
rect 4671 24 4683 104
rect 4691 24 4703 92
rect 4711 24 4723 96
<< psubstratepcontact >>
rect 4 4564 4776 4576
rect 4 4084 4776 4096
rect 4 3604 4776 3616
rect 4 3124 4776 3136
rect 4 2644 4776 2656
rect 4 2164 4776 2176
rect 4 1684 4776 1696
rect 4 1204 4776 1216
rect 4 724 4776 736
rect 4 244 4776 256
<< nsubstratencontact >>
rect 4 4324 4776 4336
rect 4 3844 4776 3856
rect 4 3364 4776 3376
rect 4 2884 4776 2896
rect 4 2404 4776 2416
rect 4 1924 4776 1936
rect 4 1444 4776 1456
rect 4 964 4776 976
rect 4 484 4776 496
rect 4 4 4776 16
<< polysilicon >>
rect 43 4556 47 4560
rect 65 4556 69 4560
rect 133 4556 137 4560
rect 143 4556 147 4560
rect 205 4556 209 4560
rect 225 4556 229 4560
rect 245 4556 249 4560
rect 291 4556 295 4560
rect 313 4556 317 4560
rect 385 4556 389 4560
rect 405 4556 409 4560
rect 465 4556 469 4560
rect 485 4556 489 4560
rect 531 4556 535 4560
rect 553 4556 557 4560
rect 625 4556 629 4560
rect 671 4556 675 4560
rect 691 4556 695 4560
rect 751 4556 755 4560
rect 811 4556 815 4560
rect 833 4556 837 4560
rect 843 4556 847 4560
rect 863 4556 867 4560
rect 871 4556 875 4560
rect 917 4556 921 4560
rect 939 4556 943 4560
rect 949 4556 953 4560
rect 971 4556 975 4560
rect 981 4556 985 4560
rect 1001 4556 1005 4560
rect 1051 4556 1055 4560
rect 1071 4556 1075 4560
rect 1091 4556 1095 4560
rect 1151 4556 1155 4560
rect 1173 4556 1177 4560
rect 1183 4556 1187 4560
rect 1203 4556 1207 4560
rect 1211 4556 1215 4560
rect 1257 4556 1261 4560
rect 1279 4556 1283 4560
rect 1289 4556 1293 4560
rect 1311 4556 1315 4560
rect 1321 4556 1325 4560
rect 1341 4556 1345 4560
rect 1391 4556 1395 4560
rect 1411 4556 1415 4560
rect 1431 4556 1435 4560
rect 1495 4556 1499 4560
rect 1515 4556 1519 4560
rect 1525 4556 1529 4560
rect 1547 4556 1551 4560
rect 1557 4556 1561 4560
rect 1579 4556 1583 4560
rect 1625 4556 1629 4560
rect 1633 4556 1637 4560
rect 1653 4556 1657 4560
rect 1663 4556 1667 4560
rect 1685 4556 1689 4560
rect 1733 4556 1737 4560
rect 1743 4556 1747 4560
rect 1811 4556 1815 4560
rect 1833 4556 1837 4560
rect 1843 4556 1847 4560
rect 1863 4556 1867 4560
rect 1871 4556 1875 4560
rect 1917 4556 1921 4560
rect 1939 4556 1943 4560
rect 1949 4556 1953 4560
rect 1971 4556 1975 4560
rect 1981 4556 1985 4560
rect 2001 4556 2005 4560
rect 2051 4556 2055 4560
rect 2071 4556 2075 4560
rect 2091 4556 2095 4560
rect 2111 4556 2115 4560
rect 2208 4556 2212 4560
rect 2216 4556 2220 4560
rect 2224 4556 2228 4560
rect 2285 4556 2289 4560
rect 2305 4556 2309 4560
rect 2325 4556 2329 4560
rect 2385 4556 2389 4560
rect 2431 4556 2435 4560
rect 2451 4556 2455 4560
rect 2525 4556 2529 4560
rect 2571 4556 2575 4560
rect 2591 4556 2595 4560
rect 2611 4556 2615 4560
rect 2671 4556 2675 4560
rect 2693 4556 2697 4560
rect 2751 4556 2755 4560
rect 2773 4556 2777 4560
rect 2843 4556 2847 4560
rect 2865 4556 2869 4560
rect 2948 4556 2952 4560
rect 2956 4556 2960 4560
rect 2964 4556 2968 4560
rect 3035 4556 3039 4560
rect 3055 4556 3059 4560
rect 3065 4556 3069 4560
rect 3123 4556 3127 4560
rect 3145 4556 3149 4560
rect 3228 4556 3232 4560
rect 3236 4556 3240 4560
rect 3244 4556 3248 4560
rect 3293 4556 3297 4560
rect 3303 4556 3307 4560
rect 3374 4556 3378 4560
rect 3382 4556 3386 4560
rect 3404 4556 3408 4560
rect 3471 4556 3475 4560
rect 3533 4556 3537 4560
rect 3543 4556 3547 4560
rect 3612 4556 3616 4560
rect 3620 4556 3624 4560
rect 3628 4556 3632 4560
rect 3714 4556 3718 4560
rect 3722 4556 3726 4560
rect 3744 4556 3748 4560
rect 3811 4556 3815 4560
rect 3831 4556 3835 4560
rect 3851 4556 3855 4560
rect 3925 4556 3929 4560
rect 3945 4556 3949 4560
rect 3965 4556 3969 4560
rect 4048 4556 4052 4560
rect 4056 4556 4060 4560
rect 4064 4556 4068 4560
rect 4148 4556 4152 4560
rect 4156 4556 4160 4560
rect 4164 4556 4168 4560
rect 4214 4556 4218 4560
rect 4222 4556 4226 4560
rect 4244 4556 4248 4560
rect 4313 4556 4317 4560
rect 4323 4556 4327 4560
rect 4412 4556 4416 4560
rect 4434 4556 4438 4560
rect 4442 4556 4446 4560
rect 4505 4556 4509 4560
rect 4552 4556 4556 4560
rect 4560 4556 4564 4560
rect 4568 4556 4572 4560
rect 4652 4556 4656 4560
rect 4660 4556 4664 4560
rect 4668 4556 4672 4560
rect 43 4510 47 4516
rect 43 4498 45 4510
rect 65 4459 69 4536
rect 133 4496 137 4516
rect 123 4489 137 4496
rect 143 4496 147 4516
rect 143 4489 151 4496
rect 123 4473 129 4489
rect 126 4461 129 4473
rect 65 4447 74 4459
rect 43 4430 45 4442
rect 43 4424 47 4430
rect 65 4384 69 4447
rect 125 4384 129 4461
rect 145 4473 151 4489
rect 145 4461 154 4473
rect 145 4384 149 4461
rect 205 4439 209 4516
rect 225 4493 229 4516
rect 245 4511 249 4516
rect 245 4504 258 4511
rect 225 4481 234 4493
rect 207 4427 214 4439
rect 210 4384 214 4427
rect 232 4424 236 4481
rect 254 4459 258 4504
rect 291 4459 295 4536
rect 313 4510 317 4516
rect 315 4498 317 4510
rect 385 4459 389 4536
rect 405 4459 409 4536
rect 465 4459 469 4536
rect 485 4459 489 4536
rect 531 4459 535 4536
rect 553 4510 557 4516
rect 555 4498 557 4510
rect 286 4447 295 4459
rect 386 4447 401 4459
rect 254 4436 258 4447
rect 240 4428 258 4436
rect 240 4424 244 4428
rect 291 4384 295 4447
rect 315 4430 317 4442
rect 313 4424 317 4430
rect 397 4424 401 4447
rect 405 4447 414 4459
rect 466 4447 481 4459
rect 405 4424 409 4447
rect 477 4424 481 4447
rect 485 4447 494 4459
rect 526 4447 535 4459
rect 485 4424 489 4447
rect 531 4384 535 4447
rect 625 4479 629 4536
rect 625 4467 634 4479
rect 555 4430 557 4442
rect 553 4424 557 4430
rect 625 4384 629 4467
rect 671 4459 675 4536
rect 691 4459 695 4536
rect 751 4479 755 4536
rect 746 4467 755 4479
rect 666 4447 675 4459
rect 671 4424 675 4447
rect 679 4447 694 4459
rect 679 4424 683 4447
rect 751 4384 755 4467
rect 811 4448 815 4516
rect 833 4487 837 4536
rect 843 4515 847 4536
rect 863 4524 867 4536
rect 871 4532 875 4536
rect 871 4528 905 4532
rect 863 4520 893 4524
rect 863 4519 881 4520
rect 843 4511 867 4515
rect 811 4436 813 4448
rect 811 4424 815 4436
rect 833 4429 837 4475
rect 829 4423 837 4429
rect 829 4394 833 4423
rect 861 4416 867 4511
rect 829 4387 837 4394
rect 833 4364 837 4387
rect 841 4364 845 4404
rect 861 4384 865 4416
rect 901 4402 905 4528
rect 917 4422 921 4536
rect 939 4524 943 4536
rect 941 4512 943 4524
rect 949 4524 953 4536
rect 949 4512 951 4524
rect 869 4390 893 4392
rect 869 4388 905 4390
rect 869 4384 873 4388
rect 915 4384 919 4410
rect 933 4402 937 4512
rect 971 4504 975 4536
rect 942 4500 975 4504
rect 942 4436 946 4500
rect 962 4451 966 4480
rect 981 4478 985 4536
rect 1001 4479 1005 4516
rect 1051 4511 1055 4516
rect 1042 4504 1055 4511
rect 962 4443 971 4451
rect 942 4424 945 4436
rect 935 4384 939 4390
rect 947 4384 951 4424
rect 967 4384 971 4443
rect 981 4384 985 4466
rect 1001 4424 1005 4467
rect 1042 4459 1046 4504
rect 1071 4493 1075 4516
rect 1066 4481 1075 4493
rect 1042 4436 1046 4447
rect 1042 4428 1060 4436
rect 1056 4424 1060 4428
rect 1064 4424 1068 4481
rect 1091 4439 1095 4516
rect 1151 4448 1155 4516
rect 1173 4487 1177 4536
rect 1183 4515 1187 4536
rect 1203 4524 1207 4536
rect 1211 4532 1215 4536
rect 1211 4528 1245 4532
rect 1203 4520 1233 4524
rect 1203 4519 1221 4520
rect 1183 4511 1207 4515
rect 1086 4427 1093 4439
rect 1151 4436 1153 4448
rect 1086 4384 1090 4427
rect 1151 4424 1155 4436
rect 1173 4429 1177 4475
rect 1169 4423 1177 4429
rect 1169 4394 1173 4423
rect 1201 4416 1207 4511
rect 1169 4387 1177 4394
rect 1173 4364 1177 4387
rect 1181 4364 1185 4404
rect 1201 4384 1205 4416
rect 1241 4402 1245 4528
rect 1257 4422 1261 4536
rect 1279 4524 1283 4536
rect 1281 4512 1283 4524
rect 1289 4524 1293 4536
rect 1289 4512 1291 4524
rect 1209 4390 1233 4392
rect 1209 4388 1245 4390
rect 1209 4384 1213 4388
rect 1255 4384 1259 4410
rect 1273 4402 1277 4512
rect 1311 4504 1315 4536
rect 1282 4500 1315 4504
rect 1282 4436 1286 4500
rect 1302 4451 1306 4480
rect 1321 4478 1325 4536
rect 1341 4479 1345 4516
rect 1391 4511 1395 4516
rect 1382 4504 1395 4511
rect 1302 4443 1311 4451
rect 1282 4424 1285 4436
rect 1275 4384 1279 4390
rect 1287 4384 1291 4424
rect 1307 4384 1311 4443
rect 1321 4384 1325 4466
rect 1341 4424 1345 4467
rect 1382 4459 1386 4504
rect 1411 4493 1415 4516
rect 1406 4481 1415 4493
rect 1382 4436 1386 4447
rect 1382 4428 1400 4436
rect 1396 4424 1400 4428
rect 1404 4424 1408 4481
rect 1431 4439 1435 4516
rect 1495 4479 1499 4516
rect 1515 4478 1519 4536
rect 1525 4504 1529 4536
rect 1547 4524 1551 4536
rect 1549 4512 1551 4524
rect 1557 4524 1561 4536
rect 1557 4512 1559 4524
rect 1525 4500 1558 4504
rect 1426 4427 1433 4439
rect 1426 4384 1430 4427
rect 1495 4424 1499 4467
rect 1515 4384 1519 4466
rect 1534 4451 1538 4480
rect 1529 4443 1538 4451
rect 1529 4384 1533 4443
rect 1554 4436 1558 4500
rect 1555 4424 1558 4436
rect 1549 4384 1553 4424
rect 1563 4402 1567 4512
rect 1579 4422 1583 4536
rect 1625 4532 1629 4536
rect 1595 4528 1629 4532
rect 1561 4384 1565 4390
rect 1581 4384 1585 4410
rect 1595 4402 1599 4528
rect 1633 4524 1637 4536
rect 1607 4520 1637 4524
rect 1619 4519 1637 4520
rect 1653 4515 1657 4536
rect 1633 4511 1657 4515
rect 1633 4416 1639 4511
rect 1663 4487 1667 4536
rect 1663 4429 1667 4475
rect 1685 4448 1689 4516
rect 1733 4496 1737 4516
rect 1729 4489 1737 4496
rect 1743 4496 1747 4516
rect 1743 4489 1757 4496
rect 1729 4473 1735 4489
rect 1726 4461 1735 4473
rect 1687 4436 1689 4448
rect 1663 4423 1671 4429
rect 1685 4424 1689 4436
rect 1607 4390 1631 4392
rect 1595 4388 1631 4390
rect 1627 4384 1631 4388
rect 1635 4384 1639 4416
rect 1655 4364 1659 4404
rect 1667 4394 1671 4423
rect 1663 4387 1671 4394
rect 1663 4364 1667 4387
rect 1731 4384 1735 4461
rect 1751 4473 1757 4489
rect 1751 4461 1754 4473
rect 1751 4384 1755 4461
rect 1811 4448 1815 4516
rect 1833 4487 1837 4536
rect 1843 4515 1847 4536
rect 1863 4524 1867 4536
rect 1871 4532 1875 4536
rect 1871 4528 1905 4532
rect 1863 4520 1893 4524
rect 1863 4519 1881 4520
rect 1843 4511 1867 4515
rect 1811 4436 1813 4448
rect 1811 4424 1815 4436
rect 1833 4429 1837 4475
rect 1829 4423 1837 4429
rect 1829 4394 1833 4423
rect 1861 4416 1867 4511
rect 1829 4387 1837 4394
rect 1833 4364 1837 4387
rect 1841 4364 1845 4404
rect 1861 4384 1865 4416
rect 1901 4402 1905 4528
rect 1917 4422 1921 4536
rect 1939 4524 1943 4536
rect 1941 4512 1943 4524
rect 1949 4524 1953 4536
rect 1949 4512 1951 4524
rect 1869 4390 1893 4392
rect 1869 4388 1905 4390
rect 1869 4384 1873 4388
rect 1915 4384 1919 4410
rect 1933 4402 1937 4512
rect 1971 4504 1975 4536
rect 1942 4500 1975 4504
rect 1942 4436 1946 4500
rect 1962 4451 1966 4480
rect 1981 4478 1985 4536
rect 2001 4479 2005 4516
rect 2051 4509 2055 4516
rect 2040 4505 2055 4509
rect 1962 4443 1971 4451
rect 1942 4424 1945 4436
rect 1935 4384 1939 4390
rect 1947 4384 1951 4424
rect 1967 4384 1971 4443
rect 1981 4384 1985 4466
rect 2001 4424 2005 4467
rect 2040 4459 2046 4505
rect 2071 4493 2075 4516
rect 2091 4493 2095 4516
rect 2066 4481 2075 4493
rect 2041 4432 2046 4447
rect 2069 4432 2075 4481
rect 2041 4428 2055 4432
rect 2051 4424 2055 4428
rect 2061 4428 2075 4432
rect 2061 4424 2065 4428
rect 2091 4424 2095 4481
rect 2111 4459 2115 4516
rect 2111 4447 2113 4459
rect 2111 4432 2115 4447
rect 2208 4439 2212 4496
rect 2101 4428 2115 4432
rect 2101 4424 2105 4428
rect 2185 4427 2193 4439
rect 2205 4427 2212 4439
rect 2185 4384 2189 4427
rect 2216 4419 2220 4496
rect 2224 4439 2228 4496
rect 2285 4439 2289 4516
rect 2305 4493 2309 4516
rect 2325 4511 2329 4516
rect 2325 4504 2338 4511
rect 2305 4481 2314 4493
rect 2224 4427 2234 4439
rect 2287 4427 2294 4439
rect 2214 4400 2220 4407
rect 2205 4396 2220 4400
rect 2234 4396 2240 4427
rect 2205 4384 2209 4396
rect 2225 4392 2240 4396
rect 2225 4384 2229 4392
rect 2290 4384 2294 4427
rect 2312 4424 2316 4481
rect 2334 4459 2338 4504
rect 2385 4479 2389 4536
rect 2385 4467 2394 4479
rect 2334 4436 2338 4447
rect 2320 4428 2338 4436
rect 2320 4424 2324 4428
rect 2385 4384 2389 4467
rect 2431 4459 2435 4536
rect 2451 4459 2455 4536
rect 2525 4479 2529 4536
rect 2571 4511 2575 4516
rect 2562 4504 2575 4511
rect 2525 4467 2534 4479
rect 2426 4447 2435 4459
rect 2431 4424 2435 4447
rect 2439 4447 2454 4459
rect 2439 4424 2443 4447
rect 2525 4384 2529 4467
rect 2562 4459 2566 4504
rect 2591 4493 2595 4516
rect 2586 4481 2595 4493
rect 2562 4436 2566 4447
rect 2562 4428 2580 4436
rect 2576 4424 2580 4428
rect 2584 4424 2588 4481
rect 2611 4439 2615 4516
rect 2671 4459 2675 4536
rect 2693 4510 2697 4516
rect 2695 4498 2697 4510
rect 2751 4459 2755 4536
rect 2773 4510 2777 4516
rect 2775 4498 2777 4510
rect 2843 4510 2847 4516
rect 2843 4498 2845 4510
rect 2666 4447 2675 4459
rect 2746 4447 2755 4459
rect 2606 4427 2613 4439
rect 2606 4384 2610 4427
rect 2671 4384 2675 4447
rect 2695 4430 2697 4442
rect 2693 4424 2697 4430
rect 2751 4384 2755 4447
rect 2865 4459 2869 4536
rect 3035 4510 3039 4516
rect 3021 4498 3033 4510
rect 2865 4447 2874 4459
rect 2775 4430 2777 4442
rect 2773 4424 2777 4430
rect 2843 4430 2845 4442
rect 2843 4424 2847 4430
rect 2865 4384 2869 4447
rect 2948 4439 2952 4496
rect 2925 4427 2933 4439
rect 2945 4427 2952 4439
rect 2925 4384 2929 4427
rect 2956 4419 2960 4496
rect 2964 4439 2968 4496
rect 2964 4427 2974 4439
rect 2954 4400 2960 4407
rect 2945 4396 2960 4400
rect 2974 4396 2980 4427
rect 3021 4424 3025 4498
rect 3055 4473 3059 4516
rect 3046 4461 3059 4473
rect 2945 4384 2949 4396
rect 2965 4392 2980 4396
rect 2965 4384 2969 4392
rect 3043 4384 3047 4461
rect 3065 4459 3069 4516
rect 3123 4510 3127 4516
rect 3123 4498 3125 4510
rect 3145 4459 3149 4536
rect 3293 4496 3297 4516
rect 3065 4447 3074 4459
rect 3145 4447 3154 4459
rect 3065 4384 3069 4447
rect 3123 4430 3125 4442
rect 3123 4424 3127 4430
rect 3145 4384 3149 4447
rect 3228 4439 3232 4496
rect 3205 4427 3213 4439
rect 3225 4427 3232 4439
rect 3205 4384 3209 4427
rect 3236 4419 3240 4496
rect 3244 4439 3248 4496
rect 3289 4489 3297 4496
rect 3303 4496 3307 4516
rect 3374 4512 3378 4516
rect 3359 4506 3378 4512
rect 3303 4489 3317 4496
rect 3359 4493 3366 4506
rect 3289 4473 3295 4489
rect 3286 4461 3295 4473
rect 3244 4427 3254 4439
rect 3234 4400 3240 4407
rect 3225 4396 3240 4400
rect 3254 4396 3260 4427
rect 3225 4384 3229 4396
rect 3245 4392 3260 4396
rect 3245 4384 3249 4392
rect 3291 4384 3295 4461
rect 3311 4473 3317 4489
rect 3311 4461 3314 4473
rect 3311 4384 3315 4461
rect 3359 4444 3366 4481
rect 3382 4479 3386 4516
rect 3404 4493 3408 4536
rect 3406 4481 3415 4493
rect 3380 4444 3386 4467
rect 3359 4438 3375 4444
rect 3380 4438 3395 4444
rect 3371 4424 3375 4438
rect 3391 4424 3395 4438
rect 3411 4424 3415 4481
rect 3471 4479 3475 4536
rect 3533 4496 3537 4516
rect 3466 4467 3475 4479
rect 3529 4489 3537 4496
rect 3543 4496 3547 4516
rect 3714 4512 3718 4516
rect 3699 4506 3718 4512
rect 3543 4489 3557 4496
rect 3529 4473 3535 4489
rect 3471 4384 3475 4467
rect 3526 4461 3535 4473
rect 3531 4384 3535 4461
rect 3551 4473 3557 4489
rect 3551 4461 3554 4473
rect 3551 4384 3555 4461
rect 3612 4439 3616 4496
rect 3606 4427 3616 4439
rect 3600 4396 3606 4427
rect 3620 4419 3624 4496
rect 3628 4439 3632 4496
rect 3699 4493 3706 4506
rect 3699 4444 3706 4481
rect 3722 4479 3726 4516
rect 3744 4493 3748 4536
rect 3811 4511 3815 4516
rect 3802 4504 3815 4511
rect 3746 4481 3755 4493
rect 3720 4444 3726 4467
rect 3628 4427 3635 4439
rect 3647 4427 3655 4439
rect 3699 4438 3715 4444
rect 3720 4438 3735 4444
rect 3620 4400 3626 4407
rect 3620 4396 3635 4400
rect 3600 4392 3615 4396
rect 3611 4384 3615 4392
rect 3631 4384 3635 4396
rect 3651 4384 3655 4427
rect 3711 4424 3715 4438
rect 3731 4424 3735 4438
rect 3751 4424 3755 4481
rect 3802 4459 3806 4504
rect 3831 4493 3835 4516
rect 3826 4481 3835 4493
rect 3802 4436 3806 4447
rect 3802 4428 3820 4436
rect 3816 4424 3820 4428
rect 3824 4424 3828 4481
rect 3851 4439 3855 4516
rect 3925 4439 3929 4516
rect 3945 4493 3949 4516
rect 3965 4511 3969 4516
rect 3965 4504 3978 4511
rect 3945 4481 3954 4493
rect 3846 4427 3853 4439
rect 3927 4427 3934 4439
rect 3846 4384 3850 4427
rect 3930 4384 3934 4427
rect 3952 4424 3956 4481
rect 3974 4459 3978 4504
rect 4214 4512 4218 4516
rect 4199 4506 4218 4512
rect 3974 4436 3978 4447
rect 4048 4439 4052 4496
rect 3960 4428 3978 4436
rect 3960 4424 3964 4428
rect 4025 4427 4033 4439
rect 4045 4427 4052 4439
rect 4025 4384 4029 4427
rect 4056 4419 4060 4496
rect 4064 4439 4068 4496
rect 4148 4439 4152 4496
rect 4064 4427 4074 4439
rect 4125 4427 4133 4439
rect 4145 4427 4152 4439
rect 4054 4400 4060 4407
rect 4045 4396 4060 4400
rect 4074 4396 4080 4427
rect 4045 4384 4049 4396
rect 4065 4392 4080 4396
rect 4065 4384 4069 4392
rect 4125 4384 4129 4427
rect 4156 4419 4160 4496
rect 4164 4439 4168 4496
rect 4199 4493 4206 4506
rect 4199 4444 4206 4481
rect 4222 4479 4226 4516
rect 4244 4493 4248 4536
rect 4313 4496 4317 4516
rect 4246 4481 4255 4493
rect 4220 4444 4226 4467
rect 4164 4427 4174 4439
rect 4199 4438 4215 4444
rect 4220 4438 4235 4444
rect 4154 4400 4160 4407
rect 4145 4396 4160 4400
rect 4174 4396 4180 4427
rect 4211 4424 4215 4438
rect 4231 4424 4235 4438
rect 4251 4424 4255 4481
rect 4309 4489 4317 4496
rect 4323 4496 4327 4516
rect 4323 4489 4337 4496
rect 4412 4493 4416 4536
rect 4309 4473 4315 4489
rect 4306 4461 4315 4473
rect 4145 4384 4149 4396
rect 4165 4392 4180 4396
rect 4165 4384 4169 4392
rect 4311 4384 4315 4461
rect 4331 4473 4337 4489
rect 4405 4481 4414 4493
rect 4331 4461 4334 4473
rect 4331 4384 4335 4461
rect 4405 4424 4409 4481
rect 4434 4479 4438 4516
rect 4442 4512 4446 4516
rect 4442 4506 4461 4512
rect 4454 4493 4461 4506
rect 4434 4444 4440 4467
rect 4454 4444 4461 4481
rect 4425 4438 4440 4444
rect 4445 4438 4461 4444
rect 4505 4479 4509 4536
rect 4505 4467 4514 4479
rect 4425 4424 4429 4438
rect 4445 4424 4449 4438
rect 4505 4384 4509 4467
rect 4552 4439 4556 4496
rect 4546 4427 4556 4439
rect 4540 4396 4546 4427
rect 4560 4419 4564 4496
rect 4568 4439 4572 4496
rect 4652 4439 4656 4496
rect 4568 4427 4575 4439
rect 4587 4427 4595 4439
rect 4646 4427 4656 4439
rect 4560 4400 4566 4407
rect 4560 4396 4575 4400
rect 4540 4392 4555 4396
rect 4551 4384 4555 4392
rect 4571 4384 4575 4396
rect 4591 4384 4595 4427
rect 4640 4396 4646 4427
rect 4660 4419 4664 4496
rect 4668 4439 4672 4496
rect 4668 4427 4675 4439
rect 4687 4427 4695 4439
rect 4660 4400 4666 4407
rect 4660 4396 4675 4400
rect 4640 4392 4655 4396
rect 4651 4384 4655 4392
rect 4671 4384 4675 4396
rect 4691 4384 4695 4427
rect 43 4340 47 4344
rect 65 4340 69 4344
rect 125 4340 129 4344
rect 145 4340 149 4344
rect 210 4340 214 4344
rect 232 4340 236 4344
rect 240 4340 244 4344
rect 291 4340 295 4344
rect 313 4340 317 4344
rect 397 4340 401 4344
rect 405 4340 409 4344
rect 477 4340 481 4344
rect 485 4340 489 4344
rect 531 4340 535 4344
rect 553 4340 557 4344
rect 625 4340 629 4344
rect 671 4340 675 4344
rect 679 4340 683 4344
rect 751 4340 755 4344
rect 811 4340 815 4344
rect 833 4340 837 4344
rect 841 4340 845 4344
rect 861 4340 865 4344
rect 869 4340 873 4344
rect 915 4340 919 4344
rect 935 4340 939 4344
rect 947 4340 951 4344
rect 967 4340 971 4344
rect 981 4340 985 4344
rect 1001 4340 1005 4344
rect 1056 4340 1060 4344
rect 1064 4340 1068 4344
rect 1086 4340 1090 4344
rect 1151 4340 1155 4344
rect 1173 4340 1177 4344
rect 1181 4340 1185 4344
rect 1201 4340 1205 4344
rect 1209 4340 1213 4344
rect 1255 4340 1259 4344
rect 1275 4340 1279 4344
rect 1287 4340 1291 4344
rect 1307 4340 1311 4344
rect 1321 4340 1325 4344
rect 1341 4340 1345 4344
rect 1396 4340 1400 4344
rect 1404 4340 1408 4344
rect 1426 4340 1430 4344
rect 1495 4340 1499 4344
rect 1515 4340 1519 4344
rect 1529 4340 1533 4344
rect 1549 4340 1553 4344
rect 1561 4340 1565 4344
rect 1581 4340 1585 4344
rect 1627 4340 1631 4344
rect 1635 4340 1639 4344
rect 1655 4340 1659 4344
rect 1663 4340 1667 4344
rect 1685 4340 1689 4344
rect 1731 4340 1735 4344
rect 1751 4340 1755 4344
rect 1811 4340 1815 4344
rect 1833 4340 1837 4344
rect 1841 4340 1845 4344
rect 1861 4340 1865 4344
rect 1869 4340 1873 4344
rect 1915 4340 1919 4344
rect 1935 4340 1939 4344
rect 1947 4340 1951 4344
rect 1967 4340 1971 4344
rect 1981 4340 1985 4344
rect 2001 4340 2005 4344
rect 2051 4340 2055 4344
rect 2061 4340 2065 4344
rect 2091 4340 2095 4344
rect 2101 4340 2105 4344
rect 2185 4340 2189 4344
rect 2205 4340 2209 4344
rect 2225 4340 2229 4344
rect 2290 4340 2294 4344
rect 2312 4340 2316 4344
rect 2320 4340 2324 4344
rect 2385 4340 2389 4344
rect 2431 4340 2435 4344
rect 2439 4340 2443 4344
rect 2525 4340 2529 4344
rect 2576 4340 2580 4344
rect 2584 4340 2588 4344
rect 2606 4340 2610 4344
rect 2671 4340 2675 4344
rect 2693 4340 2697 4344
rect 2751 4340 2755 4344
rect 2773 4340 2777 4344
rect 2843 4340 2847 4344
rect 2865 4340 2869 4344
rect 2925 4340 2929 4344
rect 2945 4340 2949 4344
rect 2965 4340 2969 4344
rect 3021 4340 3025 4344
rect 3043 4340 3047 4344
rect 3065 4340 3069 4344
rect 3123 4340 3127 4344
rect 3145 4340 3149 4344
rect 3205 4340 3209 4344
rect 3225 4340 3229 4344
rect 3245 4340 3249 4344
rect 3291 4340 3295 4344
rect 3311 4340 3315 4344
rect 3371 4340 3375 4344
rect 3391 4340 3395 4344
rect 3411 4340 3415 4344
rect 3471 4340 3475 4344
rect 3531 4340 3535 4344
rect 3551 4340 3555 4344
rect 3611 4340 3615 4344
rect 3631 4340 3635 4344
rect 3651 4340 3655 4344
rect 3711 4340 3715 4344
rect 3731 4340 3735 4344
rect 3751 4340 3755 4344
rect 3816 4340 3820 4344
rect 3824 4340 3828 4344
rect 3846 4340 3850 4344
rect 3930 4340 3934 4344
rect 3952 4340 3956 4344
rect 3960 4340 3964 4344
rect 4025 4340 4029 4344
rect 4045 4340 4049 4344
rect 4065 4340 4069 4344
rect 4125 4340 4129 4344
rect 4145 4340 4149 4344
rect 4165 4340 4169 4344
rect 4211 4340 4215 4344
rect 4231 4340 4235 4344
rect 4251 4340 4255 4344
rect 4311 4340 4315 4344
rect 4331 4340 4335 4344
rect 4405 4340 4409 4344
rect 4425 4340 4429 4344
rect 4445 4340 4449 4344
rect 4505 4340 4509 4344
rect 4551 4340 4555 4344
rect 4571 4340 4575 4344
rect 4591 4340 4595 4344
rect 4651 4340 4655 4344
rect 4671 4340 4675 4344
rect 4691 4340 4695 4344
rect 50 4316 54 4320
rect 72 4316 76 4320
rect 80 4316 84 4320
rect 141 4316 145 4320
rect 163 4316 167 4320
rect 185 4316 189 4320
rect 231 4316 235 4320
rect 239 4316 243 4320
rect 325 4316 329 4320
rect 345 4316 349 4320
rect 365 4316 369 4320
rect 411 4316 415 4320
rect 433 4316 437 4320
rect 455 4316 459 4320
rect 525 4316 529 4320
rect 545 4316 549 4320
rect 565 4316 569 4320
rect 611 4316 615 4320
rect 631 4316 635 4320
rect 651 4316 655 4320
rect 711 4316 715 4320
rect 731 4316 735 4320
rect 751 4316 755 4320
rect 811 4316 815 4320
rect 833 4316 837 4320
rect 855 4316 859 4320
rect 930 4316 934 4320
rect 952 4316 956 4320
rect 960 4316 964 4320
rect 1025 4316 1029 4320
rect 1071 4316 1075 4320
rect 1079 4316 1083 4320
rect 1151 4316 1155 4320
rect 1159 4316 1163 4320
rect 1231 4316 1235 4320
rect 1239 4316 1243 4320
rect 1311 4316 1315 4320
rect 1371 4316 1375 4320
rect 1393 4316 1397 4320
rect 1401 4316 1405 4320
rect 1421 4316 1425 4320
rect 1429 4316 1433 4320
rect 1475 4316 1479 4320
rect 1495 4316 1499 4320
rect 1507 4316 1511 4320
rect 1527 4316 1531 4320
rect 1541 4316 1545 4320
rect 1561 4316 1565 4320
rect 1616 4316 1620 4320
rect 1624 4316 1628 4320
rect 1646 4316 1650 4320
rect 1711 4316 1715 4320
rect 1719 4316 1723 4320
rect 1805 4316 1809 4320
rect 1851 4316 1855 4320
rect 1873 4316 1877 4320
rect 1881 4316 1885 4320
rect 1901 4316 1905 4320
rect 1909 4316 1913 4320
rect 1955 4316 1959 4320
rect 1975 4316 1979 4320
rect 1987 4316 1991 4320
rect 2007 4316 2011 4320
rect 2021 4316 2025 4320
rect 2041 4316 2045 4320
rect 2105 4316 2109 4320
rect 2125 4316 2129 4320
rect 2171 4316 2175 4320
rect 2181 4316 2185 4320
rect 2201 4316 2205 4320
rect 2285 4316 2289 4320
rect 2305 4316 2309 4320
rect 2325 4316 2329 4320
rect 2345 4316 2349 4320
rect 2391 4316 2395 4320
rect 2411 4316 2415 4320
rect 2490 4316 2494 4320
rect 2512 4316 2516 4320
rect 2520 4316 2524 4320
rect 2597 4316 2601 4320
rect 2605 4316 2609 4320
rect 2651 4316 2655 4320
rect 2671 4316 2675 4320
rect 2691 4316 2695 4320
rect 2765 4316 2769 4320
rect 2785 4316 2789 4320
rect 2805 4316 2809 4320
rect 2851 4316 2855 4320
rect 2873 4316 2877 4320
rect 2945 4316 2949 4320
rect 2965 4316 2969 4320
rect 2985 4316 2989 4320
rect 3045 4316 3049 4320
rect 3065 4316 3069 4320
rect 3085 4316 3089 4320
rect 3131 4316 3135 4320
rect 3151 4316 3155 4320
rect 3225 4316 3229 4320
rect 3285 4316 3289 4320
rect 3305 4316 3309 4320
rect 3325 4316 3329 4320
rect 3385 4316 3389 4320
rect 3405 4316 3409 4320
rect 3425 4316 3429 4320
rect 3485 4316 3489 4320
rect 3505 4316 3509 4320
rect 3525 4316 3529 4320
rect 3585 4316 3589 4320
rect 3605 4316 3609 4320
rect 3625 4316 3629 4320
rect 3671 4316 3675 4320
rect 3691 4316 3695 4320
rect 3711 4316 3715 4320
rect 3771 4316 3775 4320
rect 3791 4316 3795 4320
rect 3811 4316 3815 4320
rect 3876 4316 3880 4320
rect 3884 4316 3888 4320
rect 3906 4316 3910 4320
rect 3971 4316 3975 4320
rect 4031 4316 4035 4320
rect 4051 4316 4055 4320
rect 4071 4316 4075 4320
rect 4145 4316 4149 4320
rect 4165 4316 4169 4320
rect 4185 4316 4189 4320
rect 4231 4316 4235 4320
rect 4251 4316 4255 4320
rect 4271 4316 4275 4320
rect 4331 4316 4335 4320
rect 4351 4316 4355 4320
rect 4371 4316 4375 4320
rect 4436 4316 4440 4320
rect 4444 4316 4448 4320
rect 4466 4316 4470 4320
rect 4531 4316 4535 4320
rect 4551 4316 4555 4320
rect 4571 4316 4575 4320
rect 4591 4316 4595 4320
rect 4677 4316 4681 4320
rect 4685 4316 4689 4320
rect 50 4233 54 4276
rect 47 4221 54 4233
rect 45 4144 49 4221
rect 72 4179 76 4236
rect 80 4232 84 4236
rect 80 4224 98 4232
rect 94 4213 98 4224
rect 65 4167 74 4179
rect 65 4144 69 4167
rect 94 4156 98 4201
rect 85 4149 98 4156
rect 141 4162 145 4236
rect 163 4199 167 4276
rect 185 4213 189 4276
rect 231 4213 235 4236
rect 185 4201 194 4213
rect 226 4201 235 4213
rect 239 4213 243 4236
rect 239 4201 254 4213
rect 166 4187 179 4199
rect 141 4150 153 4162
rect 85 4144 89 4149
rect 155 4144 159 4150
rect 175 4144 179 4187
rect 185 4144 189 4201
rect 231 4124 235 4201
rect 251 4124 255 4201
rect 325 4179 329 4236
rect 345 4222 349 4236
rect 365 4222 369 4236
rect 345 4216 360 4222
rect 365 4216 381 4222
rect 354 4193 360 4216
rect 325 4167 334 4179
rect 332 4124 336 4167
rect 354 4144 358 4181
rect 374 4179 381 4216
rect 411 4213 415 4276
rect 406 4201 415 4213
rect 374 4154 381 4167
rect 362 4148 381 4154
rect 362 4144 366 4148
rect 411 4144 415 4201
rect 433 4199 437 4276
rect 611 4268 615 4276
rect 600 4264 615 4268
rect 631 4264 635 4276
rect 421 4187 434 4199
rect 421 4144 425 4187
rect 455 4162 459 4236
rect 525 4179 529 4236
rect 545 4222 549 4236
rect 565 4222 569 4236
rect 600 4233 606 4264
rect 620 4260 635 4264
rect 620 4253 626 4260
rect 545 4216 560 4222
rect 565 4216 581 4222
rect 606 4221 616 4233
rect 554 4193 560 4216
rect 525 4167 534 4179
rect 447 4150 459 4162
rect 441 4144 445 4150
rect 532 4124 536 4167
rect 554 4144 558 4181
rect 574 4179 581 4216
rect 574 4154 581 4167
rect 612 4164 616 4221
rect 620 4164 624 4241
rect 651 4233 655 4276
rect 628 4221 635 4233
rect 647 4221 655 4233
rect 711 4222 715 4236
rect 731 4222 735 4236
rect 628 4164 632 4221
rect 699 4216 715 4222
rect 720 4216 735 4222
rect 699 4179 706 4216
rect 720 4193 726 4216
rect 562 4148 581 4154
rect 562 4144 566 4148
rect 699 4154 706 4167
rect 699 4148 718 4154
rect 714 4144 718 4148
rect 722 4144 726 4181
rect 751 4179 755 4236
rect 811 4213 815 4276
rect 806 4201 815 4213
rect 746 4167 755 4179
rect 744 4124 748 4167
rect 811 4144 815 4201
rect 833 4199 837 4276
rect 821 4187 834 4199
rect 821 4144 825 4187
rect 855 4162 859 4236
rect 930 4233 934 4276
rect 927 4221 934 4233
rect 847 4150 859 4162
rect 841 4144 845 4150
rect 925 4144 929 4221
rect 952 4179 956 4236
rect 960 4232 964 4236
rect 960 4224 978 4232
rect 974 4213 978 4224
rect 945 4167 954 4179
rect 945 4144 949 4167
rect 974 4156 978 4201
rect 965 4149 978 4156
rect 1025 4193 1029 4276
rect 1071 4213 1075 4236
rect 1066 4201 1075 4213
rect 1079 4213 1083 4236
rect 1151 4213 1155 4236
rect 1079 4201 1094 4213
rect 1146 4201 1155 4213
rect 1159 4213 1163 4236
rect 1231 4213 1235 4236
rect 1159 4201 1174 4213
rect 1226 4201 1235 4213
rect 1239 4213 1243 4236
rect 1239 4201 1254 4213
rect 1025 4181 1034 4193
rect 965 4144 969 4149
rect 1025 4124 1029 4181
rect 1071 4124 1075 4201
rect 1091 4124 1095 4201
rect 1151 4124 1155 4201
rect 1171 4124 1175 4201
rect 1231 4124 1235 4201
rect 1251 4124 1255 4201
rect 1311 4193 1315 4276
rect 1393 4273 1397 4296
rect 1389 4266 1397 4273
rect 1389 4237 1393 4266
rect 1401 4256 1405 4296
rect 1421 4244 1425 4276
rect 1429 4272 1433 4276
rect 1429 4270 1465 4272
rect 1429 4268 1453 4270
rect 1306 4181 1315 4193
rect 1311 4124 1315 4181
rect 1371 4224 1375 4236
rect 1389 4231 1397 4237
rect 1371 4212 1373 4224
rect 1371 4144 1375 4212
rect 1393 4185 1397 4231
rect 1393 4124 1397 4173
rect 1421 4149 1427 4244
rect 1403 4145 1427 4149
rect 1403 4124 1407 4145
rect 1423 4140 1441 4141
rect 1423 4136 1453 4140
rect 1423 4124 1427 4136
rect 1461 4132 1465 4258
rect 1475 4250 1479 4276
rect 1495 4270 1499 4276
rect 1431 4128 1465 4132
rect 1431 4124 1435 4128
rect 1477 4124 1481 4238
rect 1493 4148 1497 4258
rect 1507 4236 1511 4276
rect 1502 4224 1505 4236
rect 1502 4160 1506 4224
rect 1527 4217 1531 4276
rect 1522 4209 1531 4217
rect 1522 4180 1526 4209
rect 1541 4194 1545 4276
rect 1561 4193 1565 4236
rect 1616 4232 1620 4236
rect 1602 4224 1620 4232
rect 1602 4213 1606 4224
rect 1502 4156 1535 4160
rect 1501 4136 1503 4148
rect 1499 4124 1503 4136
rect 1509 4136 1511 4148
rect 1509 4124 1513 4136
rect 1531 4124 1535 4156
rect 1541 4124 1545 4182
rect 1561 4144 1565 4181
rect 1602 4156 1606 4201
rect 1624 4179 1628 4236
rect 1646 4233 1650 4276
rect 1646 4221 1653 4233
rect 1626 4167 1635 4179
rect 1602 4149 1615 4156
rect 1611 4144 1615 4149
rect 1631 4144 1635 4167
rect 1651 4144 1655 4221
rect 1711 4213 1715 4236
rect 1706 4201 1715 4213
rect 1719 4213 1723 4236
rect 1719 4201 1734 4213
rect 1711 4124 1715 4201
rect 1731 4124 1735 4201
rect 1805 4193 1809 4276
rect 1873 4273 1877 4296
rect 1869 4266 1877 4273
rect 1869 4237 1873 4266
rect 1881 4256 1885 4296
rect 1901 4244 1905 4276
rect 1909 4272 1913 4276
rect 1909 4270 1945 4272
rect 1909 4268 1933 4270
rect 1851 4224 1855 4236
rect 1869 4231 1877 4237
rect 1851 4212 1853 4224
rect 1805 4181 1814 4193
rect 1805 4124 1809 4181
rect 1851 4144 1855 4212
rect 1873 4185 1877 4231
rect 1873 4124 1877 4173
rect 1901 4149 1907 4244
rect 1883 4145 1907 4149
rect 1883 4124 1887 4145
rect 1903 4140 1921 4141
rect 1903 4136 1933 4140
rect 1903 4124 1907 4136
rect 1941 4132 1945 4258
rect 1955 4250 1959 4276
rect 1975 4270 1979 4276
rect 1911 4128 1945 4132
rect 1911 4124 1915 4128
rect 1957 4124 1961 4238
rect 1973 4148 1977 4258
rect 1987 4236 1991 4276
rect 1982 4224 1985 4236
rect 1982 4160 1986 4224
rect 2007 4217 2011 4276
rect 2002 4209 2011 4217
rect 2002 4180 2006 4209
rect 2021 4194 2025 4276
rect 2041 4193 2045 4236
rect 2105 4199 2109 4276
rect 1982 4156 2015 4160
rect 1981 4136 1983 4148
rect 1979 4124 1983 4136
rect 1989 4136 1991 4148
rect 1989 4124 1993 4136
rect 2011 4124 2015 4156
rect 2021 4124 2025 4182
rect 2106 4187 2109 4199
rect 2041 4144 2045 4181
rect 2103 4171 2109 4187
rect 2125 4199 2129 4276
rect 2171 4232 2175 4236
rect 2162 4227 2175 4232
rect 2125 4187 2134 4199
rect 2162 4193 2166 4227
rect 2181 4213 2185 4236
rect 2201 4231 2205 4236
rect 2285 4213 2289 4236
rect 2286 4201 2289 4213
rect 2125 4171 2131 4187
rect 2103 4164 2117 4171
rect 2113 4144 2117 4164
rect 2123 4164 2131 4171
rect 2123 4144 2127 4164
rect 2162 4136 2166 4181
rect 2181 4137 2185 4201
rect 2205 4152 2215 4164
rect 2211 4144 2215 4152
rect 2280 4153 2286 4201
rect 2305 4179 2309 4236
rect 2325 4214 2329 4236
rect 2345 4214 2349 4236
rect 2325 4208 2338 4214
rect 2345 4213 2365 4214
rect 2345 4208 2353 4213
rect 2334 4179 2338 4208
rect 2307 4167 2309 4179
rect 2305 4165 2309 4167
rect 2305 4158 2318 4165
rect 2280 4149 2310 4153
rect 2306 4144 2310 4149
rect 2314 4144 2318 4158
rect 2334 4144 2338 4167
rect 2353 4159 2359 4201
rect 2391 4199 2395 4276
rect 2386 4187 2395 4199
rect 2389 4171 2395 4187
rect 2411 4199 2415 4276
rect 2490 4233 2494 4276
rect 2487 4221 2494 4233
rect 2411 4187 2414 4199
rect 2411 4171 2417 4187
rect 2389 4164 2397 4171
rect 2342 4152 2359 4159
rect 2342 4144 2346 4152
rect 2393 4144 2397 4164
rect 2403 4164 2417 4171
rect 2403 4144 2407 4164
rect 2485 4144 2489 4221
rect 2512 4179 2516 4236
rect 2520 4232 2524 4236
rect 2520 4224 2538 4232
rect 2534 4213 2538 4224
rect 2597 4213 2601 4236
rect 2586 4201 2601 4213
rect 2605 4213 2609 4236
rect 2651 4222 2655 4236
rect 2671 4222 2675 4236
rect 2639 4216 2655 4222
rect 2660 4216 2675 4222
rect 2605 4201 2614 4213
rect 2505 4167 2514 4179
rect 2505 4144 2509 4167
rect 2534 4156 2538 4201
rect 2525 4149 2538 4156
rect 2525 4144 2529 4149
rect 2162 4131 2175 4136
rect 2181 4131 2195 4137
rect 2171 4124 2175 4131
rect 2191 4124 2195 4131
rect 2585 4124 2589 4201
rect 2605 4124 2609 4201
rect 2639 4179 2646 4216
rect 2660 4193 2666 4216
rect 2639 4154 2646 4167
rect 2639 4148 2658 4154
rect 2654 4144 2658 4148
rect 2662 4144 2666 4181
rect 2691 4179 2695 4236
rect 2686 4167 2695 4179
rect 2765 4179 2769 4236
rect 2785 4222 2789 4236
rect 2805 4222 2809 4236
rect 2785 4216 2800 4222
rect 2805 4216 2821 4222
rect 2794 4193 2800 4216
rect 2765 4167 2774 4179
rect 2684 4124 2688 4167
rect 2772 4124 2776 4167
rect 2794 4144 2798 4181
rect 2814 4179 2821 4216
rect 2851 4213 2855 4276
rect 2873 4230 2877 4236
rect 2875 4218 2877 4230
rect 2945 4233 2949 4276
rect 2965 4264 2969 4276
rect 2985 4268 2989 4276
rect 2985 4264 3000 4268
rect 2965 4260 2980 4264
rect 2974 4253 2980 4260
rect 2945 4221 2953 4233
rect 2965 4221 2972 4233
rect 2846 4201 2855 4213
rect 2814 4154 2821 4167
rect 2802 4148 2821 4154
rect 2802 4144 2806 4148
rect 2851 4124 2855 4201
rect 2968 4164 2972 4221
rect 2976 4164 2980 4241
rect 2994 4233 3000 4264
rect 3045 4233 3049 4276
rect 3065 4264 3069 4276
rect 3085 4268 3089 4276
rect 3085 4264 3100 4268
rect 3065 4260 3080 4264
rect 3074 4253 3080 4260
rect 2984 4221 2994 4233
rect 3045 4221 3053 4233
rect 3065 4221 3072 4233
rect 2984 4164 2988 4221
rect 3068 4164 3072 4221
rect 3076 4164 3080 4241
rect 3094 4233 3100 4264
rect 3084 4221 3094 4233
rect 3084 4164 3088 4221
rect 3131 4199 3135 4276
rect 3126 4187 3135 4199
rect 3129 4171 3135 4187
rect 3151 4199 3155 4276
rect 3151 4187 3154 4199
rect 3225 4193 3229 4276
rect 3285 4233 3289 4276
rect 3305 4264 3309 4276
rect 3325 4268 3329 4276
rect 3325 4264 3340 4268
rect 3305 4260 3320 4264
rect 3314 4253 3320 4260
rect 3285 4221 3293 4233
rect 3305 4221 3312 4233
rect 3151 4171 3157 4187
rect 3129 4164 3137 4171
rect 2875 4150 2877 4162
rect 2873 4144 2877 4150
rect 3133 4144 3137 4164
rect 3143 4164 3157 4171
rect 3225 4181 3234 4193
rect 3143 4144 3147 4164
rect 3225 4124 3229 4181
rect 3308 4164 3312 4221
rect 3316 4164 3320 4241
rect 3334 4233 3340 4264
rect 3385 4233 3389 4276
rect 3405 4264 3409 4276
rect 3425 4268 3429 4276
rect 3425 4264 3440 4268
rect 3405 4260 3420 4264
rect 3414 4253 3420 4260
rect 3324 4221 3334 4233
rect 3385 4221 3393 4233
rect 3405 4221 3412 4233
rect 3324 4164 3328 4221
rect 3408 4164 3412 4221
rect 3416 4164 3420 4241
rect 3434 4233 3440 4264
rect 3485 4233 3489 4276
rect 3505 4264 3509 4276
rect 3525 4268 3529 4276
rect 3525 4264 3540 4268
rect 3505 4260 3520 4264
rect 3514 4253 3520 4260
rect 3424 4221 3434 4233
rect 3485 4221 3493 4233
rect 3505 4221 3512 4233
rect 3424 4164 3428 4221
rect 3508 4164 3512 4221
rect 3516 4164 3520 4241
rect 3534 4233 3540 4264
rect 3585 4233 3589 4276
rect 3605 4264 3609 4276
rect 3625 4268 3629 4276
rect 3671 4268 3675 4276
rect 3625 4264 3640 4268
rect 3605 4260 3620 4264
rect 3614 4253 3620 4260
rect 3524 4221 3534 4233
rect 3585 4221 3593 4233
rect 3605 4221 3612 4233
rect 3524 4164 3528 4221
rect 3608 4164 3612 4221
rect 3616 4164 3620 4241
rect 3634 4233 3640 4264
rect 3660 4264 3675 4268
rect 3691 4264 3695 4276
rect 3660 4233 3666 4264
rect 3680 4260 3695 4264
rect 3680 4253 3686 4260
rect 3624 4221 3634 4233
rect 3666 4221 3676 4233
rect 3624 4164 3628 4221
rect 3672 4164 3676 4221
rect 3680 4164 3684 4241
rect 3711 4233 3715 4276
rect 3688 4221 3695 4233
rect 3707 4221 3715 4233
rect 3771 4222 3775 4236
rect 3791 4222 3795 4236
rect 3688 4164 3692 4221
rect 3759 4216 3775 4222
rect 3780 4216 3795 4222
rect 3759 4179 3766 4216
rect 3780 4193 3786 4216
rect 3759 4154 3766 4167
rect 3759 4148 3778 4154
rect 3774 4144 3778 4148
rect 3782 4144 3786 4181
rect 3811 4179 3815 4236
rect 3876 4232 3880 4236
rect 3862 4224 3880 4232
rect 3862 4213 3866 4224
rect 3806 4167 3815 4179
rect 3804 4124 3808 4167
rect 3862 4156 3866 4201
rect 3884 4179 3888 4236
rect 3906 4233 3910 4276
rect 3906 4221 3913 4233
rect 3886 4167 3895 4179
rect 3862 4149 3875 4156
rect 3871 4144 3875 4149
rect 3891 4144 3895 4167
rect 3911 4144 3915 4221
rect 3971 4193 3975 4276
rect 4031 4222 4035 4236
rect 4051 4222 4055 4236
rect 3966 4181 3975 4193
rect 3971 4124 3975 4181
rect 4019 4216 4035 4222
rect 4040 4216 4055 4222
rect 4019 4179 4026 4216
rect 4040 4193 4046 4216
rect 4019 4154 4026 4167
rect 4019 4148 4038 4154
rect 4034 4144 4038 4148
rect 4042 4144 4046 4181
rect 4071 4179 4075 4236
rect 4145 4233 4149 4276
rect 4165 4264 4169 4276
rect 4185 4268 4189 4276
rect 4231 4268 4235 4276
rect 4185 4264 4200 4268
rect 4165 4260 4180 4264
rect 4174 4253 4180 4260
rect 4145 4221 4153 4233
rect 4165 4221 4172 4233
rect 4066 4167 4075 4179
rect 4064 4124 4068 4167
rect 4168 4164 4172 4221
rect 4176 4164 4180 4241
rect 4194 4233 4200 4264
rect 4220 4264 4235 4268
rect 4251 4264 4255 4276
rect 4220 4233 4226 4264
rect 4240 4260 4255 4264
rect 4240 4253 4246 4260
rect 4184 4221 4194 4233
rect 4226 4221 4236 4233
rect 4184 4164 4188 4221
rect 4232 4164 4236 4221
rect 4240 4164 4244 4241
rect 4271 4233 4275 4276
rect 4248 4221 4255 4233
rect 4267 4221 4275 4233
rect 4331 4222 4335 4236
rect 4351 4222 4355 4236
rect 4248 4164 4252 4221
rect 4319 4216 4335 4222
rect 4340 4216 4355 4222
rect 4319 4179 4326 4216
rect 4340 4193 4346 4216
rect 4319 4154 4326 4167
rect 4319 4148 4338 4154
rect 4334 4144 4338 4148
rect 4342 4144 4346 4181
rect 4371 4179 4375 4236
rect 4436 4232 4440 4236
rect 4422 4224 4440 4232
rect 4422 4213 4426 4224
rect 4366 4167 4375 4179
rect 4364 4124 4368 4167
rect 4422 4156 4426 4201
rect 4444 4179 4448 4236
rect 4466 4233 4470 4276
rect 4466 4221 4473 4233
rect 4446 4167 4455 4179
rect 4422 4149 4435 4156
rect 4431 4144 4435 4149
rect 4451 4144 4455 4167
rect 4471 4144 4475 4221
rect 4531 4214 4535 4236
rect 4551 4214 4555 4236
rect 4515 4213 4535 4214
rect 4527 4208 4535 4213
rect 4542 4208 4555 4214
rect 4521 4159 4527 4201
rect 4542 4179 4546 4208
rect 4571 4179 4575 4236
rect 4591 4213 4595 4236
rect 4677 4213 4681 4236
rect 4591 4201 4594 4213
rect 4666 4201 4681 4213
rect 4685 4213 4689 4236
rect 4685 4201 4694 4213
rect 4571 4167 4573 4179
rect 4521 4152 4538 4159
rect 4534 4144 4538 4152
rect 4542 4144 4546 4167
rect 4571 4165 4575 4167
rect 4562 4158 4575 4165
rect 4562 4144 4566 4158
rect 4594 4153 4600 4201
rect 4570 4149 4600 4153
rect 4570 4144 4574 4149
rect 4665 4124 4669 4201
rect 4685 4124 4689 4201
rect 45 4100 49 4104
rect 65 4100 69 4104
rect 85 4100 89 4104
rect 155 4100 159 4104
rect 175 4100 179 4104
rect 185 4100 189 4104
rect 231 4100 235 4104
rect 251 4100 255 4104
rect 332 4100 336 4104
rect 354 4100 358 4104
rect 362 4100 366 4104
rect 411 4100 415 4104
rect 421 4100 425 4104
rect 441 4100 445 4104
rect 532 4100 536 4104
rect 554 4100 558 4104
rect 562 4100 566 4104
rect 612 4100 616 4104
rect 620 4100 624 4104
rect 628 4100 632 4104
rect 714 4100 718 4104
rect 722 4100 726 4104
rect 744 4100 748 4104
rect 811 4100 815 4104
rect 821 4100 825 4104
rect 841 4100 845 4104
rect 925 4100 929 4104
rect 945 4100 949 4104
rect 965 4100 969 4104
rect 1025 4100 1029 4104
rect 1071 4100 1075 4104
rect 1091 4100 1095 4104
rect 1151 4100 1155 4104
rect 1171 4100 1175 4104
rect 1231 4100 1235 4104
rect 1251 4100 1255 4104
rect 1311 4100 1315 4104
rect 1371 4100 1375 4104
rect 1393 4100 1397 4104
rect 1403 4100 1407 4104
rect 1423 4100 1427 4104
rect 1431 4100 1435 4104
rect 1477 4100 1481 4104
rect 1499 4100 1503 4104
rect 1509 4100 1513 4104
rect 1531 4100 1535 4104
rect 1541 4100 1545 4104
rect 1561 4100 1565 4104
rect 1611 4100 1615 4104
rect 1631 4100 1635 4104
rect 1651 4100 1655 4104
rect 1711 4100 1715 4104
rect 1731 4100 1735 4104
rect 1805 4100 1809 4104
rect 1851 4100 1855 4104
rect 1873 4100 1877 4104
rect 1883 4100 1887 4104
rect 1903 4100 1907 4104
rect 1911 4100 1915 4104
rect 1957 4100 1961 4104
rect 1979 4100 1983 4104
rect 1989 4100 1993 4104
rect 2011 4100 2015 4104
rect 2021 4100 2025 4104
rect 2041 4100 2045 4104
rect 2113 4100 2117 4104
rect 2123 4100 2127 4104
rect 2171 4100 2175 4104
rect 2191 4100 2195 4104
rect 2211 4100 2215 4104
rect 2306 4100 2310 4104
rect 2314 4100 2318 4104
rect 2334 4100 2338 4104
rect 2342 4100 2346 4104
rect 2393 4100 2397 4104
rect 2403 4100 2407 4104
rect 2485 4100 2489 4104
rect 2505 4100 2509 4104
rect 2525 4100 2529 4104
rect 2585 4100 2589 4104
rect 2605 4100 2609 4104
rect 2654 4100 2658 4104
rect 2662 4100 2666 4104
rect 2684 4100 2688 4104
rect 2772 4100 2776 4104
rect 2794 4100 2798 4104
rect 2802 4100 2806 4104
rect 2851 4100 2855 4104
rect 2873 4100 2877 4104
rect 2968 4100 2972 4104
rect 2976 4100 2980 4104
rect 2984 4100 2988 4104
rect 3068 4100 3072 4104
rect 3076 4100 3080 4104
rect 3084 4100 3088 4104
rect 3133 4100 3137 4104
rect 3143 4100 3147 4104
rect 3225 4100 3229 4104
rect 3308 4100 3312 4104
rect 3316 4100 3320 4104
rect 3324 4100 3328 4104
rect 3408 4100 3412 4104
rect 3416 4100 3420 4104
rect 3424 4100 3428 4104
rect 3508 4100 3512 4104
rect 3516 4100 3520 4104
rect 3524 4100 3528 4104
rect 3608 4100 3612 4104
rect 3616 4100 3620 4104
rect 3624 4100 3628 4104
rect 3672 4100 3676 4104
rect 3680 4100 3684 4104
rect 3688 4100 3692 4104
rect 3774 4100 3778 4104
rect 3782 4100 3786 4104
rect 3804 4100 3808 4104
rect 3871 4100 3875 4104
rect 3891 4100 3895 4104
rect 3911 4100 3915 4104
rect 3971 4100 3975 4104
rect 4034 4100 4038 4104
rect 4042 4100 4046 4104
rect 4064 4100 4068 4104
rect 4168 4100 4172 4104
rect 4176 4100 4180 4104
rect 4184 4100 4188 4104
rect 4232 4100 4236 4104
rect 4240 4100 4244 4104
rect 4248 4100 4252 4104
rect 4334 4100 4338 4104
rect 4342 4100 4346 4104
rect 4364 4100 4368 4104
rect 4431 4100 4435 4104
rect 4451 4100 4455 4104
rect 4471 4100 4475 4104
rect 4534 4100 4538 4104
rect 4542 4100 4546 4104
rect 4562 4100 4566 4104
rect 4570 4100 4574 4104
rect 4665 4100 4669 4104
rect 4685 4100 4689 4104
rect 53 4076 57 4080
rect 63 4076 67 4080
rect 133 4076 137 4080
rect 143 4076 147 4080
rect 205 4076 209 4080
rect 225 4076 229 4080
rect 271 4076 275 4080
rect 291 4076 295 4080
rect 311 4076 315 4080
rect 385 4076 389 4080
rect 445 4076 449 4080
rect 505 4076 509 4080
rect 525 4076 529 4080
rect 571 4076 575 4080
rect 581 4076 585 4080
rect 601 4076 605 4080
rect 671 4076 675 4080
rect 691 4076 695 4080
rect 711 4076 715 4080
rect 771 4076 775 4080
rect 831 4076 835 4080
rect 851 4076 855 4080
rect 871 4076 875 4080
rect 933 4076 937 4080
rect 943 4076 947 4080
rect 1025 4076 1029 4080
rect 1085 4076 1089 4080
rect 1105 4076 1109 4080
rect 1151 4076 1155 4080
rect 1211 4076 1215 4080
rect 1231 4076 1235 4080
rect 1291 4076 1295 4080
rect 1365 4076 1369 4080
rect 1385 4076 1389 4080
rect 1445 4076 1449 4080
rect 1491 4076 1495 4080
rect 1511 4076 1515 4080
rect 1531 4076 1535 4080
rect 1591 4076 1595 4080
rect 1611 4076 1615 4080
rect 1631 4076 1635 4080
rect 1651 4076 1655 4080
rect 1713 4076 1717 4080
rect 1723 4076 1727 4080
rect 1812 4076 1816 4080
rect 1834 4076 1838 4080
rect 1842 4076 1846 4080
rect 1892 4076 1896 4080
rect 1900 4076 1904 4080
rect 1908 4076 1912 4080
rect 2005 4076 2009 4080
rect 2025 4076 2029 4080
rect 2045 4076 2049 4080
rect 2105 4076 2109 4080
rect 2188 4076 2192 4080
rect 2196 4076 2200 4080
rect 2204 4076 2208 4080
rect 2288 4076 2292 4080
rect 2296 4076 2300 4080
rect 2304 4076 2308 4080
rect 2372 4076 2376 4080
rect 2394 4076 2398 4080
rect 2402 4076 2406 4080
rect 2465 4076 2469 4080
rect 2525 4076 2529 4080
rect 2545 4076 2549 4080
rect 2565 4076 2569 4080
rect 2648 4076 2652 4080
rect 2656 4076 2660 4080
rect 2664 4076 2668 4080
rect 2732 4076 2736 4080
rect 2754 4076 2758 4080
rect 2762 4076 2766 4080
rect 2825 4076 2829 4080
rect 2845 4076 2849 4080
rect 2865 4076 2869 4080
rect 2911 4076 2915 4080
rect 2931 4076 2935 4080
rect 2951 4076 2955 4080
rect 3048 4076 3052 4080
rect 3056 4076 3060 4080
rect 3064 4076 3068 4080
rect 3125 4076 3129 4080
rect 3171 4076 3175 4080
rect 3191 4076 3195 4080
rect 3211 4076 3215 4080
rect 3274 4076 3278 4080
rect 3282 4076 3286 4080
rect 3304 4076 3308 4080
rect 3371 4076 3375 4080
rect 3391 4076 3395 4080
rect 3411 4076 3415 4080
rect 3485 4076 3489 4080
rect 3505 4076 3509 4080
rect 3525 4076 3529 4080
rect 3585 4076 3589 4080
rect 3605 4076 3609 4080
rect 3625 4076 3629 4080
rect 3692 4076 3696 4080
rect 3714 4076 3718 4080
rect 3722 4076 3726 4080
rect 3808 4076 3812 4080
rect 3816 4076 3820 4080
rect 3824 4076 3828 4080
rect 3893 4076 3897 4080
rect 3903 4076 3907 4080
rect 3973 4076 3977 4080
rect 3983 4076 3987 4080
rect 4033 4076 4037 4080
rect 4043 4076 4047 4080
rect 4148 4076 4152 4080
rect 4156 4076 4160 4080
rect 4164 4076 4168 4080
rect 4225 4076 4229 4080
rect 4245 4076 4249 4080
rect 4265 4076 4269 4080
rect 4311 4076 4315 4080
rect 4331 4076 4335 4080
rect 4351 4076 4355 4080
rect 4425 4076 4429 4080
rect 4508 4076 4512 4080
rect 4516 4076 4520 4080
rect 4524 4076 4528 4080
rect 4608 4076 4612 4080
rect 4616 4076 4620 4080
rect 4624 4076 4628 4080
rect 4674 4076 4678 4080
rect 4682 4076 4686 4080
rect 4704 4076 4708 4080
rect 53 4016 57 4036
rect 43 4009 57 4016
rect 63 4016 67 4036
rect 133 4016 137 4036
rect 63 4009 71 4016
rect 43 3993 49 4009
rect 46 3981 49 3993
rect 45 3904 49 3981
rect 65 3993 71 4009
rect 123 4009 137 4016
rect 143 4016 147 4036
rect 143 4009 151 4016
rect 123 3993 129 4009
rect 65 3981 74 3993
rect 126 3981 129 3993
rect 65 3904 69 3981
rect 125 3904 129 3981
rect 145 3993 151 4009
rect 145 3981 154 3993
rect 145 3904 149 3981
rect 205 3979 209 4056
rect 225 3979 229 4056
rect 271 4031 275 4036
rect 262 4024 275 4031
rect 262 3979 266 4024
rect 291 4013 295 4036
rect 286 4001 295 4013
rect 206 3967 221 3979
rect 217 3944 221 3967
rect 225 3967 234 3979
rect 225 3944 229 3967
rect 262 3956 266 3967
rect 262 3948 280 3956
rect 276 3944 280 3948
rect 284 3944 288 4001
rect 311 3959 315 4036
rect 385 3999 389 4056
rect 445 3999 449 4056
rect 385 3987 394 3999
rect 445 3987 454 3999
rect 306 3947 313 3959
rect 306 3904 310 3947
rect 385 3904 389 3987
rect 445 3904 449 3987
rect 505 3979 509 4056
rect 525 3979 529 4056
rect 571 3979 575 4036
rect 581 3993 585 4036
rect 601 4030 605 4036
rect 671 4031 675 4036
rect 607 4018 619 4030
rect 581 3981 594 3993
rect 506 3967 521 3979
rect 517 3944 521 3967
rect 525 3967 534 3979
rect 566 3967 575 3979
rect 525 3944 529 3967
rect 571 3904 575 3967
rect 593 3904 597 3981
rect 615 3944 619 4018
rect 662 4024 675 4031
rect 662 3979 666 4024
rect 691 4013 695 4036
rect 686 4001 695 4013
rect 662 3956 666 3967
rect 662 3948 680 3956
rect 676 3944 680 3948
rect 684 3944 688 4001
rect 711 3959 715 4036
rect 771 3999 775 4056
rect 831 4031 835 4036
rect 766 3987 775 3999
rect 706 3947 713 3959
rect 706 3904 710 3947
rect 771 3904 775 3987
rect 822 4024 835 4031
rect 822 3979 826 4024
rect 851 4013 855 4036
rect 846 4001 855 4013
rect 822 3956 826 3967
rect 822 3948 840 3956
rect 836 3944 840 3948
rect 844 3944 848 4001
rect 871 3959 875 4036
rect 933 4016 937 4036
rect 929 4009 937 4016
rect 943 4016 947 4036
rect 943 4009 957 4016
rect 929 3993 935 4009
rect 926 3981 935 3993
rect 866 3947 873 3959
rect 866 3904 870 3947
rect 931 3904 935 3981
rect 951 3993 957 4009
rect 1025 3999 1029 4056
rect 951 3981 954 3993
rect 1025 3987 1034 3999
rect 951 3904 955 3981
rect 1025 3904 1029 3987
rect 1085 3979 1089 4056
rect 1105 3979 1109 4056
rect 1151 3999 1155 4056
rect 1146 3987 1155 3999
rect 1086 3967 1101 3979
rect 1097 3944 1101 3967
rect 1105 3967 1114 3979
rect 1105 3944 1109 3967
rect 1151 3904 1155 3987
rect 1211 3979 1215 4056
rect 1231 3979 1235 4056
rect 1291 3999 1295 4056
rect 1286 3987 1295 3999
rect 1206 3967 1215 3979
rect 1211 3944 1215 3967
rect 1219 3967 1234 3979
rect 1219 3944 1223 3967
rect 1291 3904 1295 3987
rect 1365 3979 1369 4056
rect 1385 3979 1389 4056
rect 1445 3999 1449 4056
rect 1491 4031 1495 4036
rect 1482 4024 1495 4031
rect 1445 3987 1454 3999
rect 1366 3967 1381 3979
rect 1377 3944 1381 3967
rect 1385 3967 1394 3979
rect 1385 3944 1389 3967
rect 1445 3904 1449 3987
rect 1482 3979 1486 4024
rect 1511 4013 1515 4036
rect 1506 4001 1515 4013
rect 1482 3956 1486 3967
rect 1482 3948 1500 3956
rect 1496 3944 1500 3948
rect 1504 3944 1508 4001
rect 1531 3959 1535 4036
rect 1591 4029 1595 4036
rect 1580 4025 1595 4029
rect 1580 3979 1586 4025
rect 1611 4013 1615 4036
rect 1631 4013 1635 4036
rect 1606 4001 1615 4013
rect 1526 3947 1533 3959
rect 1581 3952 1586 3967
rect 1609 3952 1615 4001
rect 1581 3948 1595 3952
rect 1526 3904 1530 3947
rect 1591 3944 1595 3948
rect 1601 3948 1615 3952
rect 1601 3944 1605 3948
rect 1631 3944 1635 4001
rect 1651 3979 1655 4036
rect 1713 4016 1717 4036
rect 1709 4009 1717 4016
rect 1723 4016 1727 4036
rect 1723 4009 1737 4016
rect 1812 4013 1816 4056
rect 1709 3993 1715 4009
rect 1706 3981 1715 3993
rect 1651 3967 1653 3979
rect 1651 3952 1655 3967
rect 1641 3948 1655 3952
rect 1641 3944 1645 3948
rect 1711 3904 1715 3981
rect 1731 3993 1737 4009
rect 1805 4001 1814 4013
rect 1731 3981 1734 3993
rect 1731 3904 1735 3981
rect 1805 3944 1809 4001
rect 1834 3999 1838 4036
rect 1842 4032 1846 4036
rect 1842 4026 1861 4032
rect 1854 4013 1861 4026
rect 1834 3964 1840 3987
rect 1854 3964 1861 4001
rect 1825 3958 1840 3964
rect 1845 3958 1861 3964
rect 1892 3959 1896 4016
rect 1825 3944 1829 3958
rect 1845 3944 1849 3958
rect 1886 3947 1896 3959
rect 1880 3916 1886 3947
rect 1900 3939 1904 4016
rect 1908 3959 1912 4016
rect 2005 3959 2009 4036
rect 2025 4013 2029 4036
rect 2045 4031 2049 4036
rect 2045 4024 2058 4031
rect 2025 4001 2034 4013
rect 1908 3947 1915 3959
rect 1927 3947 1935 3959
rect 2007 3947 2014 3959
rect 1900 3920 1906 3927
rect 1900 3916 1915 3920
rect 1880 3912 1895 3916
rect 1891 3904 1895 3912
rect 1911 3904 1915 3916
rect 1931 3904 1935 3947
rect 2010 3904 2014 3947
rect 2032 3944 2036 4001
rect 2054 3979 2058 4024
rect 2105 3999 2109 4056
rect 2105 3987 2114 3999
rect 2054 3956 2058 3967
rect 2040 3948 2058 3956
rect 2040 3944 2044 3948
rect 2105 3904 2109 3987
rect 2188 3959 2192 4016
rect 2165 3947 2173 3959
rect 2185 3947 2192 3959
rect 2165 3904 2169 3947
rect 2196 3939 2200 4016
rect 2204 3959 2208 4016
rect 2288 3959 2292 4016
rect 2204 3947 2214 3959
rect 2265 3947 2273 3959
rect 2285 3947 2292 3959
rect 2194 3920 2200 3927
rect 2185 3916 2200 3920
rect 2214 3916 2220 3947
rect 2185 3904 2189 3916
rect 2205 3912 2220 3916
rect 2205 3904 2209 3912
rect 2265 3904 2269 3947
rect 2296 3939 2300 4016
rect 2304 3959 2308 4016
rect 2372 4013 2376 4056
rect 2365 4001 2374 4013
rect 2304 3947 2314 3959
rect 2294 3920 2300 3927
rect 2285 3916 2300 3920
rect 2314 3916 2320 3947
rect 2365 3944 2369 4001
rect 2394 3999 2398 4036
rect 2402 4032 2406 4036
rect 2402 4026 2421 4032
rect 2414 4013 2421 4026
rect 2394 3964 2400 3987
rect 2414 3964 2421 4001
rect 2385 3958 2400 3964
rect 2405 3958 2421 3964
rect 2465 3999 2469 4056
rect 2465 3987 2474 3999
rect 2385 3944 2389 3958
rect 2405 3944 2409 3958
rect 2285 3904 2289 3916
rect 2305 3912 2320 3916
rect 2305 3904 2309 3912
rect 2465 3904 2469 3987
rect 2525 3959 2529 4036
rect 2545 4013 2549 4036
rect 2565 4031 2569 4036
rect 2565 4024 2578 4031
rect 2545 4001 2554 4013
rect 2527 3947 2534 3959
rect 2530 3904 2534 3947
rect 2552 3944 2556 4001
rect 2574 3979 2578 4024
rect 2574 3956 2578 3967
rect 2648 3959 2652 4016
rect 2560 3948 2578 3956
rect 2560 3944 2564 3948
rect 2625 3947 2633 3959
rect 2645 3947 2652 3959
rect 2625 3904 2629 3947
rect 2656 3939 2660 4016
rect 2664 3959 2668 4016
rect 2732 4013 2736 4056
rect 2725 4001 2734 4013
rect 2664 3947 2674 3959
rect 2654 3920 2660 3927
rect 2645 3916 2660 3920
rect 2674 3916 2680 3947
rect 2725 3944 2729 4001
rect 2754 3999 2758 4036
rect 2762 4032 2766 4036
rect 2762 4026 2781 4032
rect 2774 4013 2781 4026
rect 2754 3964 2760 3987
rect 2774 3964 2781 4001
rect 2745 3958 2760 3964
rect 2765 3958 2781 3964
rect 2825 3959 2829 4036
rect 2845 4013 2849 4036
rect 2865 4031 2869 4036
rect 2911 4031 2915 4036
rect 2865 4024 2878 4031
rect 2845 4001 2854 4013
rect 2745 3944 2749 3958
rect 2765 3944 2769 3958
rect 2827 3947 2834 3959
rect 2645 3904 2649 3916
rect 2665 3912 2680 3916
rect 2665 3904 2669 3912
rect 2830 3904 2834 3947
rect 2852 3944 2856 4001
rect 2874 3979 2878 4024
rect 2902 4024 2915 4031
rect 2902 3979 2906 4024
rect 2931 4013 2935 4036
rect 2926 4001 2935 4013
rect 2874 3956 2878 3967
rect 2860 3948 2878 3956
rect 2902 3956 2906 3967
rect 2902 3948 2920 3956
rect 2860 3944 2864 3948
rect 2916 3944 2920 3948
rect 2924 3944 2928 4001
rect 2951 3959 2955 4036
rect 3048 3959 3052 4016
rect 2946 3947 2953 3959
rect 3025 3947 3033 3959
rect 3045 3947 3052 3959
rect 2946 3904 2950 3947
rect 3025 3904 3029 3947
rect 3056 3939 3060 4016
rect 3064 3959 3068 4016
rect 3125 3999 3129 4056
rect 3171 4031 3175 4036
rect 3162 4024 3175 4031
rect 3125 3987 3134 3999
rect 3064 3947 3074 3959
rect 3054 3920 3060 3927
rect 3045 3916 3060 3920
rect 3074 3916 3080 3947
rect 3045 3904 3049 3916
rect 3065 3912 3080 3916
rect 3065 3904 3069 3912
rect 3125 3904 3129 3987
rect 3162 3979 3166 4024
rect 3191 4013 3195 4036
rect 3186 4001 3195 4013
rect 3162 3956 3166 3967
rect 3162 3948 3180 3956
rect 3176 3944 3180 3948
rect 3184 3944 3188 4001
rect 3211 3959 3215 4036
rect 3274 4032 3278 4036
rect 3259 4026 3278 4032
rect 3259 4013 3266 4026
rect 3259 3964 3266 4001
rect 3282 3999 3286 4036
rect 3304 4013 3308 4056
rect 3371 4031 3375 4036
rect 3362 4024 3375 4031
rect 3306 4001 3315 4013
rect 3280 3964 3286 3987
rect 3206 3947 3213 3959
rect 3259 3958 3275 3964
rect 3280 3958 3295 3964
rect 3206 3904 3210 3947
rect 3271 3944 3275 3958
rect 3291 3944 3295 3958
rect 3311 3944 3315 4001
rect 3362 3979 3366 4024
rect 3391 4013 3395 4036
rect 3386 4001 3395 4013
rect 3362 3956 3366 3967
rect 3362 3948 3380 3956
rect 3376 3944 3380 3948
rect 3384 3944 3388 4001
rect 3411 3959 3415 4036
rect 3485 3959 3489 4036
rect 3505 4013 3509 4036
rect 3525 4031 3529 4036
rect 3525 4024 3538 4031
rect 3505 4001 3514 4013
rect 3406 3947 3413 3959
rect 3487 3947 3494 3959
rect 3406 3904 3410 3947
rect 3490 3904 3494 3947
rect 3512 3944 3516 4001
rect 3534 3979 3538 4024
rect 3534 3956 3538 3967
rect 3585 3959 3589 4036
rect 3605 4013 3609 4036
rect 3625 4031 3629 4036
rect 3625 4024 3638 4031
rect 3605 4001 3614 4013
rect 3520 3948 3538 3956
rect 3520 3944 3524 3948
rect 3587 3947 3594 3959
rect 3590 3904 3594 3947
rect 3612 3944 3616 4001
rect 3634 3979 3638 4024
rect 3692 4013 3696 4056
rect 3685 4001 3694 4013
rect 3634 3956 3638 3967
rect 3620 3948 3638 3956
rect 3620 3944 3624 3948
rect 3685 3944 3689 4001
rect 3714 3999 3718 4036
rect 3722 4032 3726 4036
rect 3722 4026 3741 4032
rect 3734 4013 3741 4026
rect 3893 4016 3897 4036
rect 3714 3964 3720 3987
rect 3734 3964 3741 4001
rect 3705 3958 3720 3964
rect 3725 3958 3741 3964
rect 3808 3959 3812 4016
rect 3705 3944 3709 3958
rect 3725 3944 3729 3958
rect 3785 3947 3793 3959
rect 3805 3947 3812 3959
rect 3785 3904 3789 3947
rect 3816 3939 3820 4016
rect 3824 3959 3828 4016
rect 3883 4009 3897 4016
rect 3903 4016 3907 4036
rect 3973 4016 3977 4036
rect 3903 4009 3911 4016
rect 3883 3993 3889 4009
rect 3886 3981 3889 3993
rect 3824 3947 3834 3959
rect 3814 3920 3820 3927
rect 3805 3916 3820 3920
rect 3834 3916 3840 3947
rect 3805 3904 3809 3916
rect 3825 3912 3840 3916
rect 3825 3904 3829 3912
rect 3885 3904 3889 3981
rect 3905 3993 3911 4009
rect 3963 4009 3977 4016
rect 3983 4016 3987 4036
rect 4033 4016 4037 4036
rect 3983 4009 3991 4016
rect 3963 3993 3969 4009
rect 3905 3981 3914 3993
rect 3966 3981 3969 3993
rect 3905 3904 3909 3981
rect 3965 3904 3969 3981
rect 3985 3993 3991 4009
rect 4029 4009 4037 4016
rect 4043 4016 4047 4036
rect 4043 4009 4057 4016
rect 4029 3993 4035 4009
rect 3985 3981 3994 3993
rect 4026 3981 4035 3993
rect 3985 3904 3989 3981
rect 4031 3904 4035 3981
rect 4051 3993 4057 4009
rect 4051 3981 4054 3993
rect 4051 3904 4055 3981
rect 4148 3959 4152 4016
rect 4125 3947 4133 3959
rect 4145 3947 4152 3959
rect 4125 3904 4129 3947
rect 4156 3939 4160 4016
rect 4164 3959 4168 4016
rect 4225 3959 4229 4036
rect 4245 4013 4249 4036
rect 4265 4031 4269 4036
rect 4311 4031 4315 4036
rect 4265 4024 4278 4031
rect 4245 4001 4254 4013
rect 4164 3947 4174 3959
rect 4227 3947 4234 3959
rect 4154 3920 4160 3927
rect 4145 3916 4160 3920
rect 4174 3916 4180 3947
rect 4145 3904 4149 3916
rect 4165 3912 4180 3916
rect 4165 3904 4169 3912
rect 4230 3904 4234 3947
rect 4252 3944 4256 4001
rect 4274 3979 4278 4024
rect 4302 4024 4315 4031
rect 4302 3979 4306 4024
rect 4331 4013 4335 4036
rect 4326 4001 4335 4013
rect 4274 3956 4278 3967
rect 4260 3948 4278 3956
rect 4302 3956 4306 3967
rect 4302 3948 4320 3956
rect 4260 3944 4264 3948
rect 4316 3944 4320 3948
rect 4324 3944 4328 4001
rect 4351 3959 4355 4036
rect 4425 3999 4429 4056
rect 4674 4032 4678 4036
rect 4659 4026 4678 4032
rect 4425 3987 4434 3999
rect 4346 3947 4353 3959
rect 4346 3904 4350 3947
rect 4425 3904 4429 3987
rect 4508 3959 4512 4016
rect 4485 3947 4493 3959
rect 4505 3947 4512 3959
rect 4485 3904 4489 3947
rect 4516 3939 4520 4016
rect 4524 3959 4528 4016
rect 4608 3959 4612 4016
rect 4524 3947 4534 3959
rect 4585 3947 4593 3959
rect 4605 3947 4612 3959
rect 4514 3920 4520 3927
rect 4505 3916 4520 3920
rect 4534 3916 4540 3947
rect 4505 3904 4509 3916
rect 4525 3912 4540 3916
rect 4525 3904 4529 3912
rect 4585 3904 4589 3947
rect 4616 3939 4620 4016
rect 4624 3959 4628 4016
rect 4659 4013 4666 4026
rect 4659 3964 4666 4001
rect 4682 3999 4686 4036
rect 4704 4013 4708 4056
rect 4706 4001 4715 4013
rect 4680 3964 4686 3987
rect 4624 3947 4634 3959
rect 4659 3958 4675 3964
rect 4680 3958 4695 3964
rect 4614 3920 4620 3927
rect 4605 3916 4620 3920
rect 4634 3916 4640 3947
rect 4671 3944 4675 3958
rect 4691 3944 4695 3958
rect 4711 3944 4715 4001
rect 4605 3904 4609 3916
rect 4625 3912 4640 3916
rect 4625 3904 4629 3912
rect 45 3860 49 3864
rect 65 3860 69 3864
rect 125 3860 129 3864
rect 145 3860 149 3864
rect 217 3860 221 3864
rect 225 3860 229 3864
rect 276 3860 280 3864
rect 284 3860 288 3864
rect 306 3860 310 3864
rect 385 3860 389 3864
rect 445 3860 449 3864
rect 517 3860 521 3864
rect 525 3860 529 3864
rect 571 3860 575 3864
rect 593 3860 597 3864
rect 615 3860 619 3864
rect 676 3860 680 3864
rect 684 3860 688 3864
rect 706 3860 710 3864
rect 771 3860 775 3864
rect 836 3860 840 3864
rect 844 3860 848 3864
rect 866 3860 870 3864
rect 931 3860 935 3864
rect 951 3860 955 3864
rect 1025 3860 1029 3864
rect 1097 3860 1101 3864
rect 1105 3860 1109 3864
rect 1151 3860 1155 3864
rect 1211 3860 1215 3864
rect 1219 3860 1223 3864
rect 1291 3860 1295 3864
rect 1377 3860 1381 3864
rect 1385 3860 1389 3864
rect 1445 3860 1449 3864
rect 1496 3860 1500 3864
rect 1504 3860 1508 3864
rect 1526 3860 1530 3864
rect 1591 3860 1595 3864
rect 1601 3860 1605 3864
rect 1631 3860 1635 3864
rect 1641 3860 1645 3864
rect 1711 3860 1715 3864
rect 1731 3860 1735 3864
rect 1805 3860 1809 3864
rect 1825 3860 1829 3864
rect 1845 3860 1849 3864
rect 1891 3860 1895 3864
rect 1911 3860 1915 3864
rect 1931 3860 1935 3864
rect 2010 3860 2014 3864
rect 2032 3860 2036 3864
rect 2040 3860 2044 3864
rect 2105 3860 2109 3864
rect 2165 3860 2169 3864
rect 2185 3860 2189 3864
rect 2205 3860 2209 3864
rect 2265 3860 2269 3864
rect 2285 3860 2289 3864
rect 2305 3860 2309 3864
rect 2365 3860 2369 3864
rect 2385 3860 2389 3864
rect 2405 3860 2409 3864
rect 2465 3860 2469 3864
rect 2530 3860 2534 3864
rect 2552 3860 2556 3864
rect 2560 3860 2564 3864
rect 2625 3860 2629 3864
rect 2645 3860 2649 3864
rect 2665 3860 2669 3864
rect 2725 3860 2729 3864
rect 2745 3860 2749 3864
rect 2765 3860 2769 3864
rect 2830 3860 2834 3864
rect 2852 3860 2856 3864
rect 2860 3860 2864 3864
rect 2916 3860 2920 3864
rect 2924 3860 2928 3864
rect 2946 3860 2950 3864
rect 3025 3860 3029 3864
rect 3045 3860 3049 3864
rect 3065 3860 3069 3864
rect 3125 3860 3129 3864
rect 3176 3860 3180 3864
rect 3184 3860 3188 3864
rect 3206 3860 3210 3864
rect 3271 3860 3275 3864
rect 3291 3860 3295 3864
rect 3311 3860 3315 3864
rect 3376 3860 3380 3864
rect 3384 3860 3388 3864
rect 3406 3860 3410 3864
rect 3490 3860 3494 3864
rect 3512 3860 3516 3864
rect 3520 3860 3524 3864
rect 3590 3860 3594 3864
rect 3612 3860 3616 3864
rect 3620 3860 3624 3864
rect 3685 3860 3689 3864
rect 3705 3860 3709 3864
rect 3725 3860 3729 3864
rect 3785 3860 3789 3864
rect 3805 3860 3809 3864
rect 3825 3860 3829 3864
rect 3885 3860 3889 3864
rect 3905 3860 3909 3864
rect 3965 3860 3969 3864
rect 3985 3860 3989 3864
rect 4031 3860 4035 3864
rect 4051 3860 4055 3864
rect 4125 3860 4129 3864
rect 4145 3860 4149 3864
rect 4165 3860 4169 3864
rect 4230 3860 4234 3864
rect 4252 3860 4256 3864
rect 4260 3860 4264 3864
rect 4316 3860 4320 3864
rect 4324 3860 4328 3864
rect 4346 3860 4350 3864
rect 4425 3860 4429 3864
rect 4485 3860 4489 3864
rect 4505 3860 4509 3864
rect 4525 3860 4529 3864
rect 4585 3860 4589 3864
rect 4605 3860 4609 3864
rect 4625 3860 4629 3864
rect 4671 3860 4675 3864
rect 4691 3860 4695 3864
rect 4711 3860 4715 3864
rect 50 3836 54 3840
rect 72 3836 76 3840
rect 80 3836 84 3840
rect 145 3836 149 3840
rect 191 3836 195 3840
rect 213 3836 217 3840
rect 221 3836 225 3840
rect 241 3836 245 3840
rect 249 3836 253 3840
rect 295 3836 299 3840
rect 315 3836 319 3840
rect 327 3836 331 3840
rect 347 3836 351 3840
rect 361 3836 365 3840
rect 381 3836 385 3840
rect 450 3836 454 3840
rect 472 3836 476 3840
rect 480 3836 484 3840
rect 531 3836 535 3840
rect 553 3836 557 3840
rect 575 3836 579 3840
rect 655 3836 659 3840
rect 675 3836 679 3840
rect 685 3836 689 3840
rect 745 3836 749 3840
rect 765 3836 769 3840
rect 815 3836 819 3840
rect 835 3836 839 3840
rect 849 3836 853 3840
rect 869 3836 873 3840
rect 881 3836 885 3840
rect 901 3836 905 3840
rect 947 3836 951 3840
rect 955 3836 959 3840
rect 975 3836 979 3840
rect 983 3836 987 3840
rect 1005 3836 1009 3840
rect 1063 3836 1067 3840
rect 1085 3836 1089 3840
rect 1131 3836 1135 3840
rect 1153 3836 1157 3840
rect 1161 3836 1165 3840
rect 1181 3836 1185 3840
rect 1189 3836 1193 3840
rect 1235 3836 1239 3840
rect 1255 3836 1259 3840
rect 1267 3836 1271 3840
rect 1287 3836 1291 3840
rect 1301 3836 1305 3840
rect 1321 3836 1325 3840
rect 1376 3836 1380 3840
rect 1384 3836 1388 3840
rect 1406 3836 1410 3840
rect 1471 3836 1475 3840
rect 1491 3836 1495 3840
rect 1551 3836 1555 3840
rect 1571 3836 1575 3840
rect 1631 3836 1635 3840
rect 1653 3836 1657 3840
rect 1711 3836 1715 3840
rect 1733 3836 1737 3840
rect 1741 3836 1745 3840
rect 1761 3836 1765 3840
rect 1769 3836 1773 3840
rect 1815 3836 1819 3840
rect 1835 3836 1839 3840
rect 1847 3836 1851 3840
rect 1867 3836 1871 3840
rect 1881 3836 1885 3840
rect 1901 3836 1905 3840
rect 1965 3836 1969 3840
rect 2025 3836 2029 3840
rect 2045 3836 2049 3840
rect 2065 3836 2069 3840
rect 2125 3836 2129 3840
rect 2171 3836 2175 3840
rect 2191 3836 2195 3840
rect 2211 3836 2215 3840
rect 2290 3836 2294 3840
rect 2312 3836 2316 3840
rect 2320 3836 2324 3840
rect 2385 3836 2389 3840
rect 2405 3836 2409 3840
rect 2425 3836 2429 3840
rect 2485 3836 2489 3840
rect 2505 3836 2509 3840
rect 2525 3836 2529 3840
rect 2585 3836 2589 3840
rect 2605 3836 2609 3840
rect 2625 3836 2629 3840
rect 2671 3836 2675 3840
rect 2691 3836 2695 3840
rect 2711 3836 2715 3840
rect 2785 3836 2789 3840
rect 2805 3836 2809 3840
rect 2825 3836 2829 3840
rect 2885 3836 2889 3840
rect 2945 3836 2949 3840
rect 3005 3836 3009 3840
rect 3025 3836 3029 3840
rect 3045 3836 3049 3840
rect 3105 3836 3109 3840
rect 3125 3836 3129 3840
rect 3145 3836 3149 3840
rect 3205 3836 3209 3840
rect 3225 3836 3229 3840
rect 3245 3836 3249 3840
rect 3305 3836 3309 3840
rect 3370 3836 3374 3840
rect 3392 3836 3396 3840
rect 3400 3836 3404 3840
rect 3465 3836 3469 3840
rect 3485 3836 3489 3840
rect 3531 3836 3535 3840
rect 3553 3836 3557 3840
rect 3575 3836 3579 3840
rect 3645 3836 3649 3840
rect 3665 3836 3669 3840
rect 3685 3836 3689 3840
rect 3745 3836 3749 3840
rect 3765 3836 3769 3840
rect 3785 3836 3789 3840
rect 3845 3836 3849 3840
rect 3891 3836 3895 3840
rect 3911 3836 3915 3840
rect 3931 3836 3935 3840
rect 4010 3836 4014 3840
rect 4032 3836 4036 3840
rect 4040 3836 4044 3840
rect 4096 3836 4100 3840
rect 4104 3836 4108 3840
rect 4126 3836 4130 3840
rect 4191 3836 4195 3840
rect 4211 3836 4215 3840
rect 4231 3836 4235 3840
rect 4305 3836 4309 3840
rect 4325 3836 4329 3840
rect 4345 3836 4349 3840
rect 4391 3836 4395 3840
rect 4411 3836 4415 3840
rect 4431 3836 4435 3840
rect 4505 3836 4509 3840
rect 4565 3836 4569 3840
rect 4585 3836 4589 3840
rect 4605 3836 4609 3840
rect 4651 3836 4655 3840
rect 4671 3836 4675 3840
rect 4691 3836 4695 3840
rect 50 3753 54 3796
rect 47 3741 54 3753
rect 45 3664 49 3741
rect 72 3699 76 3756
rect 80 3752 84 3756
rect 80 3744 98 3752
rect 94 3733 98 3744
rect 65 3687 74 3699
rect 65 3664 69 3687
rect 94 3676 98 3721
rect 85 3669 98 3676
rect 145 3713 149 3796
rect 213 3793 217 3816
rect 209 3786 217 3793
rect 209 3757 213 3786
rect 221 3776 225 3816
rect 241 3764 245 3796
rect 249 3792 253 3796
rect 249 3790 285 3792
rect 249 3788 273 3790
rect 191 3744 195 3756
rect 209 3751 217 3757
rect 191 3732 193 3744
rect 145 3701 154 3713
rect 85 3664 89 3669
rect 145 3644 149 3701
rect 191 3664 195 3732
rect 213 3705 217 3751
rect 213 3644 217 3693
rect 241 3669 247 3764
rect 223 3665 247 3669
rect 223 3644 227 3665
rect 243 3660 261 3661
rect 243 3656 273 3660
rect 243 3644 247 3656
rect 281 3652 285 3778
rect 295 3770 299 3796
rect 315 3790 319 3796
rect 251 3648 285 3652
rect 251 3644 255 3648
rect 297 3644 301 3758
rect 313 3668 317 3778
rect 327 3756 331 3796
rect 322 3744 325 3756
rect 322 3680 326 3744
rect 347 3737 351 3796
rect 342 3729 351 3737
rect 342 3700 346 3729
rect 361 3714 365 3796
rect 381 3713 385 3756
rect 450 3753 454 3796
rect 447 3741 454 3753
rect 322 3676 355 3680
rect 321 3656 323 3668
rect 319 3644 323 3656
rect 329 3656 331 3668
rect 329 3644 333 3656
rect 351 3644 355 3676
rect 361 3644 365 3702
rect 381 3664 385 3701
rect 445 3664 449 3741
rect 472 3699 476 3756
rect 480 3752 484 3756
rect 480 3744 498 3752
rect 494 3733 498 3744
rect 531 3733 535 3796
rect 526 3721 535 3733
rect 465 3687 474 3699
rect 465 3664 469 3687
rect 494 3676 498 3721
rect 485 3669 498 3676
rect 485 3664 489 3669
rect 531 3664 535 3721
rect 553 3719 557 3796
rect 541 3707 554 3719
rect 541 3664 545 3707
rect 575 3682 579 3756
rect 655 3751 659 3756
rect 675 3733 679 3756
rect 685 3752 689 3756
rect 685 3747 698 3752
rect 567 3670 579 3682
rect 645 3672 655 3684
rect 561 3664 565 3670
rect 645 3664 649 3672
rect 675 3657 679 3721
rect 665 3651 679 3657
rect 694 3713 698 3747
rect 745 3719 749 3796
rect 746 3707 749 3719
rect 694 3656 698 3701
rect 743 3691 749 3707
rect 765 3719 769 3796
rect 765 3707 774 3719
rect 815 3713 819 3756
rect 835 3714 839 3796
rect 849 3737 853 3796
rect 869 3756 873 3796
rect 881 3790 885 3796
rect 875 3744 878 3756
rect 849 3729 858 3737
rect 765 3691 771 3707
rect 743 3684 757 3691
rect 753 3664 757 3684
rect 763 3684 771 3691
rect 763 3664 767 3684
rect 815 3664 819 3701
rect 685 3651 698 3656
rect 665 3644 669 3651
rect 685 3644 689 3651
rect 835 3644 839 3702
rect 854 3700 858 3729
rect 874 3680 878 3744
rect 845 3676 878 3680
rect 845 3644 849 3676
rect 883 3668 887 3778
rect 901 3770 905 3796
rect 947 3792 951 3796
rect 915 3790 951 3792
rect 927 3788 951 3790
rect 869 3656 871 3668
rect 867 3644 871 3656
rect 877 3656 879 3668
rect 877 3644 881 3656
rect 899 3644 903 3758
rect 915 3652 919 3778
rect 955 3764 959 3796
rect 975 3776 979 3816
rect 983 3793 987 3816
rect 983 3786 991 3793
rect 953 3669 959 3764
rect 987 3757 991 3786
rect 983 3751 991 3757
rect 983 3705 987 3751
rect 1005 3744 1009 3756
rect 1007 3732 1009 3744
rect 1063 3750 1067 3756
rect 1063 3738 1065 3750
rect 953 3665 977 3669
rect 939 3660 957 3661
rect 927 3656 957 3660
rect 915 3648 949 3652
rect 945 3644 949 3648
rect 953 3644 957 3656
rect 973 3644 977 3665
rect 983 3644 987 3693
rect 1005 3664 1009 3732
rect 1085 3733 1089 3796
rect 1153 3793 1157 3816
rect 1149 3786 1157 3793
rect 1149 3757 1153 3786
rect 1161 3776 1165 3816
rect 1181 3764 1185 3796
rect 1189 3792 1193 3796
rect 1189 3790 1225 3792
rect 1189 3788 1213 3790
rect 1131 3744 1135 3756
rect 1149 3751 1157 3757
rect 1085 3721 1094 3733
rect 1131 3732 1133 3744
rect 1063 3670 1065 3682
rect 1063 3664 1067 3670
rect 1085 3644 1089 3721
rect 1131 3664 1135 3732
rect 1153 3705 1157 3751
rect 1153 3644 1157 3693
rect 1181 3669 1187 3764
rect 1163 3665 1187 3669
rect 1163 3644 1167 3665
rect 1183 3660 1201 3661
rect 1183 3656 1213 3660
rect 1183 3644 1187 3656
rect 1221 3652 1225 3778
rect 1235 3770 1239 3796
rect 1255 3790 1259 3796
rect 1191 3648 1225 3652
rect 1191 3644 1195 3648
rect 1237 3644 1241 3758
rect 1253 3668 1257 3778
rect 1267 3756 1271 3796
rect 1262 3744 1265 3756
rect 1262 3680 1266 3744
rect 1287 3737 1291 3796
rect 1282 3729 1291 3737
rect 1282 3700 1286 3729
rect 1301 3714 1305 3796
rect 1321 3713 1325 3756
rect 1376 3752 1380 3756
rect 1362 3744 1380 3752
rect 1362 3733 1366 3744
rect 1262 3676 1295 3680
rect 1261 3656 1263 3668
rect 1259 3644 1263 3656
rect 1269 3656 1271 3668
rect 1269 3644 1273 3656
rect 1291 3644 1295 3676
rect 1301 3644 1305 3702
rect 1321 3664 1325 3701
rect 1362 3676 1366 3721
rect 1384 3699 1388 3756
rect 1406 3753 1410 3796
rect 1406 3741 1413 3753
rect 1386 3687 1395 3699
rect 1362 3669 1375 3676
rect 1371 3664 1375 3669
rect 1391 3664 1395 3687
rect 1411 3664 1415 3741
rect 1471 3719 1475 3796
rect 1466 3707 1475 3719
rect 1469 3691 1475 3707
rect 1491 3719 1495 3796
rect 1551 3719 1555 3796
rect 1491 3707 1494 3719
rect 1546 3707 1555 3719
rect 1491 3691 1497 3707
rect 1469 3684 1477 3691
rect 1473 3664 1477 3684
rect 1483 3684 1497 3691
rect 1549 3691 1555 3707
rect 1571 3719 1575 3796
rect 1631 3733 1635 3796
rect 1733 3793 1737 3816
rect 1729 3786 1737 3793
rect 1729 3757 1733 3786
rect 1741 3776 1745 3816
rect 1761 3764 1765 3796
rect 1769 3792 1773 3796
rect 1769 3790 1805 3792
rect 1769 3788 1793 3790
rect 1653 3750 1657 3756
rect 1655 3738 1657 3750
rect 1711 3744 1715 3756
rect 1729 3751 1737 3757
rect 1626 3721 1635 3733
rect 1571 3707 1574 3719
rect 1571 3691 1577 3707
rect 1549 3684 1557 3691
rect 1483 3664 1487 3684
rect 1553 3664 1557 3684
rect 1563 3684 1577 3691
rect 1563 3664 1567 3684
rect 1631 3644 1635 3721
rect 1711 3732 1713 3744
rect 1655 3670 1657 3682
rect 1653 3664 1657 3670
rect 1711 3664 1715 3732
rect 1733 3705 1737 3751
rect 1733 3644 1737 3693
rect 1761 3669 1767 3764
rect 1743 3665 1767 3669
rect 1743 3644 1747 3665
rect 1763 3660 1781 3661
rect 1763 3656 1793 3660
rect 1763 3644 1767 3656
rect 1801 3652 1805 3778
rect 1815 3770 1819 3796
rect 1835 3790 1839 3796
rect 1771 3648 1805 3652
rect 1771 3644 1775 3648
rect 1817 3644 1821 3758
rect 1833 3668 1837 3778
rect 1847 3756 1851 3796
rect 1842 3744 1845 3756
rect 1842 3680 1846 3744
rect 1867 3737 1871 3796
rect 1862 3729 1871 3737
rect 1862 3700 1866 3729
rect 1881 3714 1885 3796
rect 1901 3713 1905 3756
rect 1965 3713 1969 3796
rect 1842 3676 1875 3680
rect 1841 3656 1843 3668
rect 1839 3644 1843 3656
rect 1849 3656 1851 3668
rect 1849 3644 1853 3656
rect 1871 3644 1875 3676
rect 1881 3644 1885 3702
rect 1965 3701 1974 3713
rect 1901 3664 1905 3701
rect 1965 3644 1969 3701
rect 2025 3699 2029 3756
rect 2045 3742 2049 3756
rect 2065 3742 2069 3756
rect 2045 3736 2060 3742
rect 2065 3736 2081 3742
rect 2054 3713 2060 3736
rect 2025 3687 2034 3699
rect 2032 3644 2036 3687
rect 2054 3664 2058 3701
rect 2074 3699 2081 3736
rect 2125 3713 2129 3796
rect 2171 3788 2175 3796
rect 2160 3784 2175 3788
rect 2191 3784 2195 3796
rect 2160 3753 2166 3784
rect 2180 3780 2195 3784
rect 2180 3773 2186 3780
rect 2166 3741 2176 3753
rect 2125 3701 2134 3713
rect 2074 3674 2081 3687
rect 2062 3668 2081 3674
rect 2062 3664 2066 3668
rect 2125 3644 2129 3701
rect 2172 3684 2176 3741
rect 2180 3684 2184 3761
rect 2211 3753 2215 3796
rect 2290 3753 2294 3796
rect 2188 3741 2195 3753
rect 2207 3741 2215 3753
rect 2287 3741 2294 3753
rect 2188 3684 2192 3741
rect 2285 3664 2289 3741
rect 2312 3699 2316 3756
rect 2320 3752 2324 3756
rect 2385 3753 2389 3796
rect 2405 3784 2409 3796
rect 2425 3788 2429 3796
rect 2425 3784 2440 3788
rect 2405 3780 2420 3784
rect 2414 3773 2420 3780
rect 2320 3744 2338 3752
rect 2334 3733 2338 3744
rect 2385 3741 2393 3753
rect 2405 3741 2412 3753
rect 2305 3687 2314 3699
rect 2305 3664 2309 3687
rect 2334 3676 2338 3721
rect 2408 3684 2412 3741
rect 2416 3684 2420 3761
rect 2434 3753 2440 3784
rect 2424 3741 2434 3753
rect 2424 3684 2428 3741
rect 2485 3699 2489 3756
rect 2505 3742 2509 3756
rect 2525 3742 2529 3756
rect 2585 3753 2589 3796
rect 2605 3784 2609 3796
rect 2625 3788 2629 3796
rect 2625 3784 2640 3788
rect 2605 3780 2620 3784
rect 2614 3773 2620 3780
rect 2505 3736 2520 3742
rect 2525 3736 2541 3742
rect 2585 3741 2593 3753
rect 2605 3741 2612 3753
rect 2514 3713 2520 3736
rect 2485 3687 2494 3699
rect 2325 3669 2338 3676
rect 2325 3664 2329 3669
rect 2492 3644 2496 3687
rect 2514 3664 2518 3701
rect 2534 3699 2541 3736
rect 2534 3674 2541 3687
rect 2608 3684 2612 3741
rect 2616 3684 2620 3761
rect 2634 3753 2640 3784
rect 2624 3741 2634 3753
rect 2671 3742 2675 3756
rect 2691 3742 2695 3756
rect 2624 3684 2628 3741
rect 2659 3736 2675 3742
rect 2680 3736 2695 3742
rect 2659 3699 2666 3736
rect 2680 3713 2686 3736
rect 2522 3668 2541 3674
rect 2522 3664 2526 3668
rect 2659 3674 2666 3687
rect 2659 3668 2678 3674
rect 2674 3664 2678 3668
rect 2682 3664 2686 3701
rect 2711 3699 2715 3756
rect 2706 3687 2715 3699
rect 2785 3699 2789 3756
rect 2805 3742 2809 3756
rect 2825 3742 2829 3756
rect 2805 3736 2820 3742
rect 2825 3736 2841 3742
rect 2814 3713 2820 3736
rect 2785 3687 2794 3699
rect 2704 3644 2708 3687
rect 2792 3644 2796 3687
rect 2814 3664 2818 3701
rect 2834 3699 2841 3736
rect 2885 3713 2889 3796
rect 2945 3713 2949 3796
rect 3005 3753 3009 3796
rect 3025 3784 3029 3796
rect 3045 3788 3049 3796
rect 3045 3784 3060 3788
rect 3025 3780 3040 3784
rect 3034 3773 3040 3780
rect 3005 3741 3013 3753
rect 3025 3741 3032 3753
rect 2885 3701 2894 3713
rect 2945 3701 2954 3713
rect 2834 3674 2841 3687
rect 2822 3668 2841 3674
rect 2822 3664 2826 3668
rect 2885 3644 2889 3701
rect 2945 3644 2949 3701
rect 3028 3684 3032 3741
rect 3036 3684 3040 3761
rect 3054 3753 3060 3784
rect 3044 3741 3054 3753
rect 3044 3684 3048 3741
rect 3105 3699 3109 3756
rect 3125 3742 3129 3756
rect 3145 3742 3149 3756
rect 3205 3753 3209 3796
rect 3225 3784 3229 3796
rect 3245 3788 3249 3796
rect 3245 3784 3260 3788
rect 3225 3780 3240 3784
rect 3234 3773 3240 3780
rect 3125 3736 3140 3742
rect 3145 3736 3161 3742
rect 3205 3741 3213 3753
rect 3225 3741 3232 3753
rect 3134 3713 3140 3736
rect 3105 3687 3114 3699
rect 3112 3644 3116 3687
rect 3134 3664 3138 3701
rect 3154 3699 3161 3736
rect 3154 3674 3161 3687
rect 3228 3684 3232 3741
rect 3236 3684 3240 3761
rect 3254 3753 3260 3784
rect 3244 3741 3254 3753
rect 3244 3684 3248 3741
rect 3305 3713 3309 3796
rect 3370 3753 3374 3796
rect 3367 3741 3374 3753
rect 3305 3701 3314 3713
rect 3142 3668 3161 3674
rect 3142 3664 3146 3668
rect 3305 3644 3309 3701
rect 3365 3664 3369 3741
rect 3392 3699 3396 3756
rect 3400 3752 3404 3756
rect 3400 3744 3418 3752
rect 3414 3733 3418 3744
rect 3385 3687 3394 3699
rect 3385 3664 3389 3687
rect 3414 3676 3418 3721
rect 3465 3719 3469 3796
rect 3466 3707 3469 3719
rect 3463 3691 3469 3707
rect 3485 3719 3489 3796
rect 3531 3733 3535 3796
rect 3526 3721 3535 3733
rect 3485 3707 3494 3719
rect 3485 3691 3491 3707
rect 3463 3684 3477 3691
rect 3405 3669 3418 3676
rect 3405 3664 3409 3669
rect 3473 3664 3477 3684
rect 3483 3684 3491 3691
rect 3483 3664 3487 3684
rect 3531 3664 3535 3721
rect 3553 3719 3557 3796
rect 3541 3707 3554 3719
rect 3541 3664 3545 3707
rect 3575 3682 3579 3756
rect 3645 3699 3649 3756
rect 3665 3742 3669 3756
rect 3685 3742 3689 3756
rect 3745 3753 3749 3796
rect 3765 3784 3769 3796
rect 3785 3788 3789 3796
rect 3785 3784 3800 3788
rect 3765 3780 3780 3784
rect 3774 3773 3780 3780
rect 3665 3736 3680 3742
rect 3685 3736 3701 3742
rect 3745 3741 3753 3753
rect 3765 3741 3772 3753
rect 3674 3713 3680 3736
rect 3645 3687 3654 3699
rect 3567 3670 3579 3682
rect 3561 3664 3565 3670
rect 3652 3644 3656 3687
rect 3674 3664 3678 3701
rect 3694 3699 3701 3736
rect 3694 3674 3701 3687
rect 3768 3684 3772 3741
rect 3776 3684 3780 3761
rect 3794 3753 3800 3784
rect 3784 3741 3794 3753
rect 3784 3684 3788 3741
rect 3845 3713 3849 3796
rect 3891 3742 3895 3756
rect 3911 3742 3915 3756
rect 3879 3736 3895 3742
rect 3900 3736 3915 3742
rect 3845 3701 3854 3713
rect 3682 3668 3701 3674
rect 3682 3664 3686 3668
rect 3845 3644 3849 3701
rect 3879 3699 3886 3736
rect 3900 3713 3906 3736
rect 3879 3674 3886 3687
rect 3879 3668 3898 3674
rect 3894 3664 3898 3668
rect 3902 3664 3906 3701
rect 3931 3699 3935 3756
rect 4010 3753 4014 3796
rect 4007 3741 4014 3753
rect 3926 3687 3935 3699
rect 3924 3644 3928 3687
rect 4005 3664 4009 3741
rect 4032 3699 4036 3756
rect 4040 3752 4044 3756
rect 4096 3752 4100 3756
rect 4040 3744 4058 3752
rect 4054 3733 4058 3744
rect 4082 3744 4100 3752
rect 4082 3733 4086 3744
rect 4025 3687 4034 3699
rect 4025 3664 4029 3687
rect 4054 3676 4058 3721
rect 4045 3669 4058 3676
rect 4082 3676 4086 3721
rect 4104 3699 4108 3756
rect 4126 3753 4130 3796
rect 4391 3788 4395 3796
rect 4380 3784 4395 3788
rect 4411 3784 4415 3796
rect 4126 3741 4133 3753
rect 4191 3742 4195 3756
rect 4211 3742 4215 3756
rect 4106 3687 4115 3699
rect 4082 3669 4095 3676
rect 4045 3664 4049 3669
rect 4091 3664 4095 3669
rect 4111 3664 4115 3687
rect 4131 3664 4135 3741
rect 4179 3736 4195 3742
rect 4200 3736 4215 3742
rect 4179 3699 4186 3736
rect 4200 3713 4206 3736
rect 4179 3674 4186 3687
rect 4179 3668 4198 3674
rect 4194 3664 4198 3668
rect 4202 3664 4206 3701
rect 4231 3699 4235 3756
rect 4226 3687 4235 3699
rect 4305 3699 4309 3756
rect 4325 3742 4329 3756
rect 4345 3742 4349 3756
rect 4380 3753 4386 3784
rect 4400 3780 4415 3784
rect 4400 3773 4406 3780
rect 4325 3736 4340 3742
rect 4345 3736 4361 3742
rect 4386 3741 4396 3753
rect 4334 3713 4340 3736
rect 4305 3687 4314 3699
rect 4224 3644 4228 3687
rect 4312 3644 4316 3687
rect 4334 3664 4338 3701
rect 4354 3699 4361 3736
rect 4354 3674 4361 3687
rect 4392 3684 4396 3741
rect 4400 3684 4404 3761
rect 4431 3753 4435 3796
rect 4408 3741 4415 3753
rect 4427 3741 4435 3753
rect 4408 3684 4412 3741
rect 4505 3713 4509 3796
rect 4565 3753 4569 3796
rect 4585 3784 4589 3796
rect 4605 3788 4609 3796
rect 4651 3788 4655 3796
rect 4605 3784 4620 3788
rect 4585 3780 4600 3784
rect 4594 3773 4600 3780
rect 4565 3741 4573 3753
rect 4585 3741 4592 3753
rect 4505 3701 4514 3713
rect 4342 3668 4361 3674
rect 4342 3664 4346 3668
rect 4505 3644 4509 3701
rect 4588 3684 4592 3741
rect 4596 3684 4600 3761
rect 4614 3753 4620 3784
rect 4640 3784 4655 3788
rect 4671 3784 4675 3796
rect 4640 3753 4646 3784
rect 4660 3780 4675 3784
rect 4660 3773 4666 3780
rect 4604 3741 4614 3753
rect 4646 3741 4656 3753
rect 4604 3684 4608 3741
rect 4652 3684 4656 3741
rect 4660 3684 4664 3761
rect 4691 3753 4695 3796
rect 4668 3741 4675 3753
rect 4687 3741 4695 3753
rect 4668 3684 4672 3741
rect 45 3620 49 3624
rect 65 3620 69 3624
rect 85 3620 89 3624
rect 145 3620 149 3624
rect 191 3620 195 3624
rect 213 3620 217 3624
rect 223 3620 227 3624
rect 243 3620 247 3624
rect 251 3620 255 3624
rect 297 3620 301 3624
rect 319 3620 323 3624
rect 329 3620 333 3624
rect 351 3620 355 3624
rect 361 3620 365 3624
rect 381 3620 385 3624
rect 445 3620 449 3624
rect 465 3620 469 3624
rect 485 3620 489 3624
rect 531 3620 535 3624
rect 541 3620 545 3624
rect 561 3620 565 3624
rect 645 3620 649 3624
rect 665 3620 669 3624
rect 685 3620 689 3624
rect 753 3620 757 3624
rect 763 3620 767 3624
rect 815 3620 819 3624
rect 835 3620 839 3624
rect 845 3620 849 3624
rect 867 3620 871 3624
rect 877 3620 881 3624
rect 899 3620 903 3624
rect 945 3620 949 3624
rect 953 3620 957 3624
rect 973 3620 977 3624
rect 983 3620 987 3624
rect 1005 3620 1009 3624
rect 1063 3620 1067 3624
rect 1085 3620 1089 3624
rect 1131 3620 1135 3624
rect 1153 3620 1157 3624
rect 1163 3620 1167 3624
rect 1183 3620 1187 3624
rect 1191 3620 1195 3624
rect 1237 3620 1241 3624
rect 1259 3620 1263 3624
rect 1269 3620 1273 3624
rect 1291 3620 1295 3624
rect 1301 3620 1305 3624
rect 1321 3620 1325 3624
rect 1371 3620 1375 3624
rect 1391 3620 1395 3624
rect 1411 3620 1415 3624
rect 1473 3620 1477 3624
rect 1483 3620 1487 3624
rect 1553 3620 1557 3624
rect 1563 3620 1567 3624
rect 1631 3620 1635 3624
rect 1653 3620 1657 3624
rect 1711 3620 1715 3624
rect 1733 3620 1737 3624
rect 1743 3620 1747 3624
rect 1763 3620 1767 3624
rect 1771 3620 1775 3624
rect 1817 3620 1821 3624
rect 1839 3620 1843 3624
rect 1849 3620 1853 3624
rect 1871 3620 1875 3624
rect 1881 3620 1885 3624
rect 1901 3620 1905 3624
rect 1965 3620 1969 3624
rect 2032 3620 2036 3624
rect 2054 3620 2058 3624
rect 2062 3620 2066 3624
rect 2125 3620 2129 3624
rect 2172 3620 2176 3624
rect 2180 3620 2184 3624
rect 2188 3620 2192 3624
rect 2285 3620 2289 3624
rect 2305 3620 2309 3624
rect 2325 3620 2329 3624
rect 2408 3620 2412 3624
rect 2416 3620 2420 3624
rect 2424 3620 2428 3624
rect 2492 3620 2496 3624
rect 2514 3620 2518 3624
rect 2522 3620 2526 3624
rect 2608 3620 2612 3624
rect 2616 3620 2620 3624
rect 2624 3620 2628 3624
rect 2674 3620 2678 3624
rect 2682 3620 2686 3624
rect 2704 3620 2708 3624
rect 2792 3620 2796 3624
rect 2814 3620 2818 3624
rect 2822 3620 2826 3624
rect 2885 3620 2889 3624
rect 2945 3620 2949 3624
rect 3028 3620 3032 3624
rect 3036 3620 3040 3624
rect 3044 3620 3048 3624
rect 3112 3620 3116 3624
rect 3134 3620 3138 3624
rect 3142 3620 3146 3624
rect 3228 3620 3232 3624
rect 3236 3620 3240 3624
rect 3244 3620 3248 3624
rect 3305 3620 3309 3624
rect 3365 3620 3369 3624
rect 3385 3620 3389 3624
rect 3405 3620 3409 3624
rect 3473 3620 3477 3624
rect 3483 3620 3487 3624
rect 3531 3620 3535 3624
rect 3541 3620 3545 3624
rect 3561 3620 3565 3624
rect 3652 3620 3656 3624
rect 3674 3620 3678 3624
rect 3682 3620 3686 3624
rect 3768 3620 3772 3624
rect 3776 3620 3780 3624
rect 3784 3620 3788 3624
rect 3845 3620 3849 3624
rect 3894 3620 3898 3624
rect 3902 3620 3906 3624
rect 3924 3620 3928 3624
rect 4005 3620 4009 3624
rect 4025 3620 4029 3624
rect 4045 3620 4049 3624
rect 4091 3620 4095 3624
rect 4111 3620 4115 3624
rect 4131 3620 4135 3624
rect 4194 3620 4198 3624
rect 4202 3620 4206 3624
rect 4224 3620 4228 3624
rect 4312 3620 4316 3624
rect 4334 3620 4338 3624
rect 4342 3620 4346 3624
rect 4392 3620 4396 3624
rect 4400 3620 4404 3624
rect 4408 3620 4412 3624
rect 4505 3620 4509 3624
rect 4588 3620 4592 3624
rect 4596 3620 4600 3624
rect 4604 3620 4608 3624
rect 4652 3620 4656 3624
rect 4660 3620 4664 3624
rect 4668 3620 4672 3624
rect 35 3596 39 3600
rect 55 3596 59 3600
rect 65 3596 69 3600
rect 87 3596 91 3600
rect 97 3596 101 3600
rect 119 3596 123 3600
rect 165 3596 169 3600
rect 173 3596 177 3600
rect 193 3596 197 3600
rect 203 3596 207 3600
rect 225 3596 229 3600
rect 293 3596 297 3600
rect 303 3596 307 3600
rect 365 3596 369 3600
rect 385 3596 389 3600
rect 405 3596 409 3600
rect 473 3596 477 3600
rect 483 3596 487 3600
rect 568 3596 572 3600
rect 576 3596 580 3600
rect 584 3596 588 3600
rect 645 3596 649 3600
rect 705 3596 709 3600
rect 725 3596 729 3600
rect 745 3596 749 3600
rect 805 3596 809 3600
rect 825 3596 829 3600
rect 845 3596 849 3600
rect 891 3596 895 3600
rect 965 3596 969 3600
rect 985 3596 989 3600
rect 1031 3596 1035 3600
rect 1053 3596 1057 3600
rect 1063 3596 1067 3600
rect 1083 3596 1087 3600
rect 1091 3596 1095 3600
rect 1137 3596 1141 3600
rect 1159 3596 1163 3600
rect 1169 3596 1173 3600
rect 1191 3596 1195 3600
rect 1201 3596 1205 3600
rect 1221 3596 1225 3600
rect 1271 3596 1275 3600
rect 1331 3596 1335 3600
rect 1351 3596 1355 3600
rect 1411 3596 1415 3600
rect 1431 3596 1435 3600
rect 1451 3596 1455 3600
rect 1513 3596 1517 3600
rect 1523 3596 1527 3600
rect 1603 3596 1607 3600
rect 1625 3596 1629 3600
rect 1685 3596 1689 3600
rect 1731 3596 1735 3600
rect 1753 3596 1757 3600
rect 1763 3596 1767 3600
rect 1783 3596 1787 3600
rect 1791 3596 1795 3600
rect 1837 3596 1841 3600
rect 1859 3596 1863 3600
rect 1869 3596 1873 3600
rect 1891 3596 1895 3600
rect 1901 3596 1905 3600
rect 1921 3596 1925 3600
rect 1971 3596 1975 3600
rect 1991 3596 1995 3600
rect 2011 3596 2015 3600
rect 2031 3596 2035 3600
rect 2093 3596 2097 3600
rect 2103 3596 2107 3600
rect 2192 3596 2196 3600
rect 2214 3596 2218 3600
rect 2222 3596 2226 3600
rect 2308 3596 2312 3600
rect 2316 3596 2320 3600
rect 2324 3596 2328 3600
rect 2385 3596 2389 3600
rect 2468 3596 2472 3600
rect 2476 3596 2480 3600
rect 2484 3596 2488 3600
rect 2568 3596 2572 3600
rect 2576 3596 2580 3600
rect 2584 3596 2588 3600
rect 2645 3596 2649 3600
rect 2665 3596 2669 3600
rect 2685 3596 2689 3600
rect 2731 3596 2735 3600
rect 2751 3596 2755 3600
rect 2771 3596 2775 3600
rect 2833 3596 2837 3600
rect 2843 3596 2847 3600
rect 2911 3596 2915 3600
rect 2931 3596 2935 3600
rect 2951 3596 2955 3600
rect 3011 3596 3015 3600
rect 3031 3596 3035 3600
rect 3105 3596 3109 3600
rect 3125 3596 3129 3600
rect 3145 3596 3149 3600
rect 3194 3596 3198 3600
rect 3202 3596 3206 3600
rect 3222 3596 3226 3600
rect 3230 3596 3234 3600
rect 3313 3596 3317 3600
rect 3323 3596 3327 3600
rect 3393 3596 3397 3600
rect 3403 3596 3407 3600
rect 3473 3596 3477 3600
rect 3483 3596 3487 3600
rect 3551 3596 3555 3600
rect 3571 3596 3575 3600
rect 3633 3596 3637 3600
rect 3643 3596 3647 3600
rect 3713 3596 3717 3600
rect 3723 3596 3727 3600
rect 3813 3596 3817 3600
rect 3823 3596 3827 3600
rect 3885 3596 3889 3600
rect 3905 3596 3909 3600
rect 3953 3596 3957 3600
rect 3963 3596 3967 3600
rect 4033 3596 4037 3600
rect 4043 3596 4047 3600
rect 4111 3596 4115 3600
rect 4131 3596 4135 3600
rect 4151 3596 4155 3600
rect 4248 3596 4252 3600
rect 4256 3596 4260 3600
rect 4264 3596 4268 3600
rect 4312 3596 4316 3600
rect 4320 3596 4324 3600
rect 4328 3596 4332 3600
rect 4414 3596 4418 3600
rect 4422 3596 4426 3600
rect 4444 3596 4448 3600
rect 4511 3596 4515 3600
rect 4608 3596 4612 3600
rect 4616 3596 4620 3600
rect 4624 3596 4628 3600
rect 4672 3596 4676 3600
rect 4680 3596 4684 3600
rect 4688 3596 4692 3600
rect 35 3519 39 3556
rect 55 3518 59 3576
rect 65 3544 69 3576
rect 87 3564 91 3576
rect 89 3552 91 3564
rect 97 3564 101 3576
rect 97 3552 99 3564
rect 65 3540 98 3544
rect 35 3464 39 3507
rect 55 3424 59 3506
rect 74 3491 78 3520
rect 69 3483 78 3491
rect 69 3424 73 3483
rect 94 3476 98 3540
rect 95 3464 98 3476
rect 89 3424 93 3464
rect 103 3442 107 3552
rect 119 3462 123 3576
rect 165 3572 169 3576
rect 135 3568 169 3572
rect 101 3424 105 3430
rect 121 3424 125 3450
rect 135 3442 139 3568
rect 173 3564 177 3576
rect 147 3560 177 3564
rect 159 3559 177 3560
rect 193 3555 197 3576
rect 173 3551 197 3555
rect 173 3456 179 3551
rect 203 3527 207 3576
rect 203 3469 207 3515
rect 225 3488 229 3556
rect 293 3536 297 3556
rect 283 3529 297 3536
rect 303 3536 307 3556
rect 303 3529 311 3536
rect 283 3513 289 3529
rect 286 3501 289 3513
rect 227 3476 229 3488
rect 203 3463 211 3469
rect 225 3464 229 3476
rect 147 3430 171 3432
rect 135 3428 171 3430
rect 167 3424 171 3428
rect 175 3424 179 3456
rect 195 3404 199 3444
rect 207 3434 211 3463
rect 203 3427 211 3434
rect 203 3404 207 3427
rect 285 3424 289 3501
rect 305 3513 311 3529
rect 305 3501 314 3513
rect 305 3424 309 3501
rect 365 3479 369 3556
rect 385 3533 389 3556
rect 405 3551 409 3556
rect 405 3544 418 3551
rect 385 3521 394 3533
rect 367 3467 374 3479
rect 370 3424 374 3467
rect 392 3464 396 3521
rect 414 3499 418 3544
rect 473 3536 477 3556
rect 463 3529 477 3536
rect 483 3536 487 3556
rect 483 3529 491 3536
rect 463 3513 469 3529
rect 466 3501 469 3513
rect 414 3476 418 3487
rect 400 3468 418 3476
rect 400 3464 404 3468
rect 465 3424 469 3501
rect 485 3513 491 3529
rect 485 3501 494 3513
rect 485 3424 489 3501
rect 568 3479 572 3536
rect 545 3467 553 3479
rect 565 3467 572 3479
rect 545 3424 549 3467
rect 576 3459 580 3536
rect 584 3479 588 3536
rect 645 3519 649 3576
rect 645 3507 654 3519
rect 584 3467 594 3479
rect 574 3440 580 3447
rect 565 3436 580 3440
rect 594 3436 600 3467
rect 565 3424 569 3436
rect 585 3432 600 3436
rect 585 3424 589 3432
rect 645 3424 649 3507
rect 705 3479 709 3556
rect 725 3533 729 3556
rect 745 3551 749 3556
rect 745 3544 758 3551
rect 725 3521 734 3533
rect 707 3467 714 3479
rect 710 3424 714 3467
rect 732 3464 736 3521
rect 754 3499 758 3544
rect 754 3476 758 3487
rect 805 3479 809 3556
rect 825 3533 829 3556
rect 845 3551 849 3556
rect 845 3544 858 3551
rect 825 3521 834 3533
rect 740 3468 758 3476
rect 740 3464 744 3468
rect 807 3467 814 3479
rect 810 3424 814 3467
rect 832 3464 836 3521
rect 854 3499 858 3544
rect 891 3519 895 3576
rect 886 3507 895 3519
rect 854 3476 858 3487
rect 840 3468 858 3476
rect 840 3464 844 3468
rect 891 3424 895 3507
rect 965 3499 969 3576
rect 985 3499 989 3576
rect 966 3487 981 3499
rect 977 3464 981 3487
rect 985 3487 994 3499
rect 1031 3488 1035 3556
rect 1053 3527 1057 3576
rect 1063 3555 1067 3576
rect 1083 3564 1087 3576
rect 1091 3572 1095 3576
rect 1091 3568 1125 3572
rect 1083 3560 1113 3564
rect 1083 3559 1101 3560
rect 1063 3551 1087 3555
rect 985 3464 989 3487
rect 1031 3476 1033 3488
rect 1031 3464 1035 3476
rect 1053 3469 1057 3515
rect 1049 3463 1057 3469
rect 1049 3434 1053 3463
rect 1081 3456 1087 3551
rect 1049 3427 1057 3434
rect 1053 3404 1057 3427
rect 1061 3404 1065 3444
rect 1081 3424 1085 3456
rect 1121 3442 1125 3568
rect 1137 3462 1141 3576
rect 1159 3564 1163 3576
rect 1161 3552 1163 3564
rect 1169 3564 1173 3576
rect 1169 3552 1171 3564
rect 1089 3430 1113 3432
rect 1089 3428 1125 3430
rect 1089 3424 1093 3428
rect 1135 3424 1139 3450
rect 1153 3442 1157 3552
rect 1191 3544 1195 3576
rect 1162 3540 1195 3544
rect 1162 3476 1166 3540
rect 1182 3491 1186 3520
rect 1201 3518 1205 3576
rect 1221 3519 1225 3556
rect 1271 3519 1275 3576
rect 1266 3507 1275 3519
rect 1182 3483 1191 3491
rect 1162 3464 1165 3476
rect 1155 3424 1159 3430
rect 1167 3424 1171 3464
rect 1187 3424 1191 3483
rect 1201 3424 1205 3506
rect 1221 3464 1225 3507
rect 1271 3424 1275 3507
rect 1331 3499 1335 3576
rect 1351 3499 1355 3576
rect 1411 3551 1415 3556
rect 1402 3544 1415 3551
rect 1402 3499 1406 3544
rect 1431 3533 1435 3556
rect 1426 3521 1435 3533
rect 1326 3487 1335 3499
rect 1331 3464 1335 3487
rect 1339 3487 1354 3499
rect 1339 3464 1343 3487
rect 1402 3476 1406 3487
rect 1402 3468 1420 3476
rect 1416 3464 1420 3468
rect 1424 3464 1428 3521
rect 1451 3479 1455 3556
rect 1513 3536 1517 3556
rect 1509 3529 1517 3536
rect 1523 3536 1527 3556
rect 1603 3550 1607 3556
rect 1603 3538 1605 3550
rect 1523 3529 1537 3536
rect 1509 3513 1515 3529
rect 1506 3501 1515 3513
rect 1446 3467 1453 3479
rect 1446 3424 1450 3467
rect 1511 3424 1515 3501
rect 1531 3513 1537 3529
rect 1531 3501 1534 3513
rect 1531 3424 1535 3501
rect 1625 3499 1629 3576
rect 1685 3519 1689 3576
rect 1685 3507 1694 3519
rect 1625 3487 1634 3499
rect 1603 3470 1605 3482
rect 1603 3464 1607 3470
rect 1625 3424 1629 3487
rect 1685 3424 1689 3507
rect 1731 3488 1735 3556
rect 1753 3527 1757 3576
rect 1763 3555 1767 3576
rect 1783 3564 1787 3576
rect 1791 3572 1795 3576
rect 1791 3568 1825 3572
rect 1783 3560 1813 3564
rect 1783 3559 1801 3560
rect 1763 3551 1787 3555
rect 1731 3476 1733 3488
rect 1731 3464 1735 3476
rect 1753 3469 1757 3515
rect 1749 3463 1757 3469
rect 1749 3434 1753 3463
rect 1781 3456 1787 3551
rect 1749 3427 1757 3434
rect 1753 3404 1757 3427
rect 1761 3404 1765 3444
rect 1781 3424 1785 3456
rect 1821 3442 1825 3568
rect 1837 3462 1841 3576
rect 1859 3564 1863 3576
rect 1861 3552 1863 3564
rect 1869 3564 1873 3576
rect 1869 3552 1871 3564
rect 1789 3430 1813 3432
rect 1789 3428 1825 3430
rect 1789 3424 1793 3428
rect 1835 3424 1839 3450
rect 1853 3442 1857 3552
rect 1891 3544 1895 3576
rect 1862 3540 1895 3544
rect 1862 3476 1866 3540
rect 1882 3491 1886 3520
rect 1901 3518 1905 3576
rect 1921 3519 1925 3556
rect 1971 3549 1975 3556
rect 1960 3545 1975 3549
rect 1882 3483 1891 3491
rect 1862 3464 1865 3476
rect 1855 3424 1859 3430
rect 1867 3424 1871 3464
rect 1887 3424 1891 3483
rect 1901 3424 1905 3506
rect 1921 3464 1925 3507
rect 1960 3499 1966 3545
rect 1991 3533 1995 3556
rect 2011 3533 2015 3556
rect 1986 3521 1995 3533
rect 1961 3472 1966 3487
rect 1989 3472 1995 3521
rect 1961 3468 1975 3472
rect 1971 3464 1975 3468
rect 1981 3468 1995 3472
rect 1981 3464 1985 3468
rect 2011 3464 2015 3521
rect 2031 3499 2035 3556
rect 2093 3536 2097 3556
rect 2089 3529 2097 3536
rect 2103 3536 2107 3556
rect 2103 3529 2117 3536
rect 2192 3533 2196 3576
rect 2089 3513 2095 3529
rect 2086 3501 2095 3513
rect 2031 3487 2033 3499
rect 2031 3472 2035 3487
rect 2021 3468 2035 3472
rect 2021 3464 2025 3468
rect 2091 3424 2095 3501
rect 2111 3513 2117 3529
rect 2185 3521 2194 3533
rect 2111 3501 2114 3513
rect 2111 3424 2115 3501
rect 2185 3464 2189 3521
rect 2214 3519 2218 3556
rect 2222 3552 2226 3556
rect 2222 3546 2241 3552
rect 2234 3533 2241 3546
rect 2214 3484 2220 3507
rect 2234 3484 2241 3521
rect 2205 3478 2220 3484
rect 2225 3478 2241 3484
rect 2308 3479 2312 3536
rect 2205 3464 2209 3478
rect 2225 3464 2229 3478
rect 2285 3467 2293 3479
rect 2305 3467 2312 3479
rect 2285 3424 2289 3467
rect 2316 3459 2320 3536
rect 2324 3479 2328 3536
rect 2385 3519 2389 3576
rect 2385 3507 2394 3519
rect 2324 3467 2334 3479
rect 2314 3440 2320 3447
rect 2305 3436 2320 3440
rect 2334 3436 2340 3467
rect 2305 3424 2309 3436
rect 2325 3432 2340 3436
rect 2325 3424 2329 3432
rect 2385 3424 2389 3507
rect 2468 3479 2472 3536
rect 2445 3467 2453 3479
rect 2465 3467 2472 3479
rect 2445 3424 2449 3467
rect 2476 3459 2480 3536
rect 2484 3479 2488 3536
rect 2568 3479 2572 3536
rect 2484 3467 2494 3479
rect 2545 3467 2553 3479
rect 2565 3467 2572 3479
rect 2474 3440 2480 3447
rect 2465 3436 2480 3440
rect 2494 3436 2500 3467
rect 2465 3424 2469 3436
rect 2485 3432 2500 3436
rect 2485 3424 2489 3432
rect 2545 3424 2549 3467
rect 2576 3459 2580 3536
rect 2584 3479 2588 3536
rect 2645 3479 2649 3556
rect 2665 3533 2669 3556
rect 2685 3551 2689 3556
rect 2731 3551 2735 3556
rect 2685 3544 2698 3551
rect 2665 3521 2674 3533
rect 2584 3467 2594 3479
rect 2647 3467 2654 3479
rect 2574 3440 2580 3447
rect 2565 3436 2580 3440
rect 2594 3436 2600 3467
rect 2565 3424 2569 3436
rect 2585 3432 2600 3436
rect 2585 3424 2589 3432
rect 2650 3424 2654 3467
rect 2672 3464 2676 3521
rect 2694 3499 2698 3544
rect 2722 3544 2735 3551
rect 2722 3499 2726 3544
rect 2751 3533 2755 3556
rect 2746 3521 2755 3533
rect 2694 3476 2698 3487
rect 2680 3468 2698 3476
rect 2722 3476 2726 3487
rect 2722 3468 2740 3476
rect 2680 3464 2684 3468
rect 2736 3464 2740 3468
rect 2744 3464 2748 3521
rect 2771 3479 2775 3556
rect 2833 3536 2837 3556
rect 2829 3529 2837 3536
rect 2843 3536 2847 3556
rect 2911 3551 2915 3556
rect 2902 3544 2915 3551
rect 2843 3529 2857 3536
rect 2829 3513 2835 3529
rect 2826 3501 2835 3513
rect 2766 3467 2773 3479
rect 2766 3424 2770 3467
rect 2831 3424 2835 3501
rect 2851 3513 2857 3529
rect 2851 3501 2854 3513
rect 2851 3424 2855 3501
rect 2902 3499 2906 3544
rect 2931 3533 2935 3556
rect 2926 3521 2935 3533
rect 2902 3476 2906 3487
rect 2902 3468 2920 3476
rect 2916 3464 2920 3468
rect 2924 3464 2928 3521
rect 2951 3479 2955 3556
rect 3011 3499 3015 3576
rect 3031 3499 3035 3576
rect 3006 3487 3015 3499
rect 2946 3467 2953 3479
rect 2946 3424 2950 3467
rect 3011 3464 3015 3487
rect 3019 3487 3034 3499
rect 3019 3464 3023 3487
rect 3105 3479 3109 3556
rect 3125 3533 3129 3556
rect 3145 3551 3149 3556
rect 3145 3544 3158 3551
rect 3194 3548 3198 3556
rect 3125 3521 3134 3533
rect 3107 3467 3114 3479
rect 3110 3424 3114 3467
rect 3132 3464 3136 3521
rect 3154 3499 3158 3544
rect 3181 3541 3198 3548
rect 3181 3499 3187 3541
rect 3202 3533 3206 3556
rect 3222 3542 3226 3556
rect 3230 3551 3234 3556
rect 3230 3547 3260 3551
rect 3222 3535 3235 3542
rect 3231 3533 3235 3535
rect 3231 3521 3233 3533
rect 3202 3492 3206 3521
rect 3187 3487 3195 3492
rect 3154 3476 3158 3487
rect 3175 3486 3195 3487
rect 3202 3486 3215 3492
rect 3140 3468 3158 3476
rect 3140 3464 3144 3468
rect 3191 3464 3195 3486
rect 3211 3464 3215 3486
rect 3231 3464 3235 3521
rect 3254 3499 3260 3547
rect 3313 3536 3317 3556
rect 3309 3529 3317 3536
rect 3323 3536 3327 3556
rect 3393 3536 3397 3556
rect 3323 3529 3337 3536
rect 3309 3513 3315 3529
rect 3306 3501 3315 3513
rect 3251 3487 3254 3499
rect 3251 3464 3255 3487
rect 3311 3424 3315 3501
rect 3331 3513 3337 3529
rect 3389 3529 3397 3536
rect 3403 3536 3407 3556
rect 3473 3536 3477 3556
rect 3403 3529 3417 3536
rect 3389 3513 3395 3529
rect 3331 3501 3334 3513
rect 3386 3501 3395 3513
rect 3331 3424 3335 3501
rect 3391 3424 3395 3501
rect 3411 3513 3417 3529
rect 3469 3529 3477 3536
rect 3483 3536 3487 3556
rect 3483 3529 3497 3536
rect 3469 3513 3475 3529
rect 3411 3501 3414 3513
rect 3466 3501 3475 3513
rect 3411 3424 3415 3501
rect 3471 3424 3475 3501
rect 3491 3513 3497 3529
rect 3491 3501 3494 3513
rect 3491 3424 3495 3501
rect 3551 3499 3555 3576
rect 3571 3499 3575 3576
rect 3633 3536 3637 3556
rect 3629 3529 3637 3536
rect 3643 3536 3647 3556
rect 3713 3536 3717 3556
rect 3643 3529 3657 3536
rect 3629 3513 3635 3529
rect 3626 3501 3635 3513
rect 3546 3487 3555 3499
rect 3551 3464 3555 3487
rect 3559 3487 3574 3499
rect 3559 3464 3563 3487
rect 3631 3424 3635 3501
rect 3651 3513 3657 3529
rect 3709 3529 3717 3536
rect 3723 3536 3727 3556
rect 3813 3536 3817 3556
rect 3723 3529 3737 3536
rect 3709 3513 3715 3529
rect 3651 3501 3654 3513
rect 3706 3501 3715 3513
rect 3651 3424 3655 3501
rect 3711 3424 3715 3501
rect 3731 3513 3737 3529
rect 3803 3529 3817 3536
rect 3823 3536 3827 3556
rect 3823 3529 3831 3536
rect 3803 3513 3809 3529
rect 3731 3501 3734 3513
rect 3806 3501 3809 3513
rect 3731 3424 3735 3501
rect 3805 3424 3809 3501
rect 3825 3513 3831 3529
rect 3825 3501 3834 3513
rect 3825 3424 3829 3501
rect 3885 3499 3889 3576
rect 3905 3499 3909 3576
rect 3953 3536 3957 3556
rect 3949 3529 3957 3536
rect 3963 3536 3967 3556
rect 4033 3536 4037 3556
rect 3963 3529 3977 3536
rect 3949 3513 3955 3529
rect 3946 3501 3955 3513
rect 3886 3487 3901 3499
rect 3897 3464 3901 3487
rect 3905 3487 3914 3499
rect 3905 3464 3909 3487
rect 3951 3424 3955 3501
rect 3971 3513 3977 3529
rect 4029 3529 4037 3536
rect 4043 3536 4047 3556
rect 4111 3551 4115 3556
rect 4102 3544 4115 3551
rect 4043 3529 4057 3536
rect 4029 3513 4035 3529
rect 3971 3501 3974 3513
rect 4026 3501 4035 3513
rect 3971 3424 3975 3501
rect 4031 3424 4035 3501
rect 4051 3513 4057 3529
rect 4051 3501 4054 3513
rect 4051 3424 4055 3501
rect 4102 3499 4106 3544
rect 4131 3533 4135 3556
rect 4126 3521 4135 3533
rect 4102 3476 4106 3487
rect 4102 3468 4120 3476
rect 4116 3464 4120 3468
rect 4124 3464 4128 3521
rect 4151 3479 4155 3556
rect 4414 3552 4418 3556
rect 4399 3546 4418 3552
rect 4248 3479 4252 3536
rect 4146 3467 4153 3479
rect 4225 3467 4233 3479
rect 4245 3467 4252 3479
rect 4146 3424 4150 3467
rect 4225 3424 4229 3467
rect 4256 3459 4260 3536
rect 4264 3479 4268 3536
rect 4312 3479 4316 3536
rect 4264 3467 4274 3479
rect 4306 3467 4316 3479
rect 4254 3440 4260 3447
rect 4245 3436 4260 3440
rect 4274 3436 4280 3467
rect 4245 3424 4249 3436
rect 4265 3432 4280 3436
rect 4300 3436 4306 3467
rect 4320 3459 4324 3536
rect 4328 3479 4332 3536
rect 4399 3533 4406 3546
rect 4399 3484 4406 3521
rect 4422 3519 4426 3556
rect 4444 3533 4448 3576
rect 4446 3521 4455 3533
rect 4420 3484 4426 3507
rect 4328 3467 4335 3479
rect 4347 3467 4355 3479
rect 4399 3478 4415 3484
rect 4420 3478 4435 3484
rect 4320 3440 4326 3447
rect 4320 3436 4335 3440
rect 4300 3432 4315 3436
rect 4265 3424 4269 3432
rect 4311 3424 4315 3432
rect 4331 3424 4335 3436
rect 4351 3424 4355 3467
rect 4411 3464 4415 3478
rect 4431 3464 4435 3478
rect 4451 3464 4455 3521
rect 4511 3519 4515 3576
rect 4506 3507 4515 3519
rect 4511 3424 4515 3507
rect 4608 3479 4612 3536
rect 4585 3467 4593 3479
rect 4605 3467 4612 3479
rect 4585 3424 4589 3467
rect 4616 3459 4620 3536
rect 4624 3479 4628 3536
rect 4672 3479 4676 3536
rect 4624 3467 4634 3479
rect 4666 3467 4676 3479
rect 4614 3440 4620 3447
rect 4605 3436 4620 3440
rect 4634 3436 4640 3467
rect 4605 3424 4609 3436
rect 4625 3432 4640 3436
rect 4660 3436 4666 3467
rect 4680 3459 4684 3536
rect 4688 3479 4692 3536
rect 4688 3467 4695 3479
rect 4707 3467 4715 3479
rect 4680 3440 4686 3447
rect 4680 3436 4695 3440
rect 4660 3432 4675 3436
rect 4625 3424 4629 3432
rect 4671 3424 4675 3432
rect 4691 3424 4695 3436
rect 4711 3424 4715 3467
rect 35 3380 39 3384
rect 55 3380 59 3384
rect 69 3380 73 3384
rect 89 3380 93 3384
rect 101 3380 105 3384
rect 121 3380 125 3384
rect 167 3380 171 3384
rect 175 3380 179 3384
rect 195 3380 199 3384
rect 203 3380 207 3384
rect 225 3380 229 3384
rect 285 3380 289 3384
rect 305 3380 309 3384
rect 370 3380 374 3384
rect 392 3380 396 3384
rect 400 3380 404 3384
rect 465 3380 469 3384
rect 485 3380 489 3384
rect 545 3380 549 3384
rect 565 3380 569 3384
rect 585 3380 589 3384
rect 645 3380 649 3384
rect 710 3380 714 3384
rect 732 3380 736 3384
rect 740 3380 744 3384
rect 810 3380 814 3384
rect 832 3380 836 3384
rect 840 3380 844 3384
rect 891 3380 895 3384
rect 977 3380 981 3384
rect 985 3380 989 3384
rect 1031 3380 1035 3384
rect 1053 3380 1057 3384
rect 1061 3380 1065 3384
rect 1081 3380 1085 3384
rect 1089 3380 1093 3384
rect 1135 3380 1139 3384
rect 1155 3380 1159 3384
rect 1167 3380 1171 3384
rect 1187 3380 1191 3384
rect 1201 3380 1205 3384
rect 1221 3380 1225 3384
rect 1271 3380 1275 3384
rect 1331 3380 1335 3384
rect 1339 3380 1343 3384
rect 1416 3380 1420 3384
rect 1424 3380 1428 3384
rect 1446 3380 1450 3384
rect 1511 3380 1515 3384
rect 1531 3380 1535 3384
rect 1603 3380 1607 3384
rect 1625 3380 1629 3384
rect 1685 3380 1689 3384
rect 1731 3380 1735 3384
rect 1753 3380 1757 3384
rect 1761 3380 1765 3384
rect 1781 3380 1785 3384
rect 1789 3380 1793 3384
rect 1835 3380 1839 3384
rect 1855 3380 1859 3384
rect 1867 3380 1871 3384
rect 1887 3380 1891 3384
rect 1901 3380 1905 3384
rect 1921 3380 1925 3384
rect 1971 3380 1975 3384
rect 1981 3380 1985 3384
rect 2011 3380 2015 3384
rect 2021 3380 2025 3384
rect 2091 3380 2095 3384
rect 2111 3380 2115 3384
rect 2185 3380 2189 3384
rect 2205 3380 2209 3384
rect 2225 3380 2229 3384
rect 2285 3380 2289 3384
rect 2305 3380 2309 3384
rect 2325 3380 2329 3384
rect 2385 3380 2389 3384
rect 2445 3380 2449 3384
rect 2465 3380 2469 3384
rect 2485 3380 2489 3384
rect 2545 3380 2549 3384
rect 2565 3380 2569 3384
rect 2585 3380 2589 3384
rect 2650 3380 2654 3384
rect 2672 3380 2676 3384
rect 2680 3380 2684 3384
rect 2736 3380 2740 3384
rect 2744 3380 2748 3384
rect 2766 3380 2770 3384
rect 2831 3380 2835 3384
rect 2851 3380 2855 3384
rect 2916 3380 2920 3384
rect 2924 3380 2928 3384
rect 2946 3380 2950 3384
rect 3011 3380 3015 3384
rect 3019 3380 3023 3384
rect 3110 3380 3114 3384
rect 3132 3380 3136 3384
rect 3140 3380 3144 3384
rect 3191 3380 3195 3384
rect 3211 3380 3215 3384
rect 3231 3380 3235 3384
rect 3251 3380 3255 3384
rect 3311 3380 3315 3384
rect 3331 3380 3335 3384
rect 3391 3380 3395 3384
rect 3411 3380 3415 3384
rect 3471 3380 3475 3384
rect 3491 3380 3495 3384
rect 3551 3380 3555 3384
rect 3559 3380 3563 3384
rect 3631 3380 3635 3384
rect 3651 3380 3655 3384
rect 3711 3380 3715 3384
rect 3731 3380 3735 3384
rect 3805 3380 3809 3384
rect 3825 3380 3829 3384
rect 3897 3380 3901 3384
rect 3905 3380 3909 3384
rect 3951 3380 3955 3384
rect 3971 3380 3975 3384
rect 4031 3380 4035 3384
rect 4051 3380 4055 3384
rect 4116 3380 4120 3384
rect 4124 3380 4128 3384
rect 4146 3380 4150 3384
rect 4225 3380 4229 3384
rect 4245 3380 4249 3384
rect 4265 3380 4269 3384
rect 4311 3380 4315 3384
rect 4331 3380 4335 3384
rect 4351 3380 4355 3384
rect 4411 3380 4415 3384
rect 4431 3380 4435 3384
rect 4451 3380 4455 3384
rect 4511 3380 4515 3384
rect 4585 3380 4589 3384
rect 4605 3380 4609 3384
rect 4625 3380 4629 3384
rect 4671 3380 4675 3384
rect 4691 3380 4695 3384
rect 4711 3380 4715 3384
rect 35 3356 39 3360
rect 55 3356 59 3360
rect 69 3356 73 3360
rect 89 3356 93 3360
rect 101 3356 105 3360
rect 121 3356 125 3360
rect 167 3356 171 3360
rect 175 3356 179 3360
rect 195 3356 199 3360
rect 203 3356 207 3360
rect 225 3356 229 3360
rect 285 3356 289 3360
rect 305 3356 309 3360
rect 325 3356 329 3360
rect 345 3356 349 3360
rect 391 3356 395 3360
rect 411 3356 415 3360
rect 476 3356 480 3360
rect 484 3356 488 3360
rect 506 3356 510 3360
rect 576 3356 580 3360
rect 584 3356 588 3360
rect 606 3356 610 3360
rect 685 3356 689 3360
rect 705 3356 709 3360
rect 751 3356 755 3360
rect 825 3356 829 3360
rect 845 3356 849 3360
rect 865 3356 869 3360
rect 885 3356 889 3360
rect 905 3356 909 3360
rect 925 3356 929 3360
rect 945 3356 949 3360
rect 965 3356 969 3360
rect 1011 3356 1015 3360
rect 1031 3356 1035 3360
rect 1051 3356 1055 3360
rect 1071 3356 1075 3360
rect 1091 3356 1095 3360
rect 1111 3356 1115 3360
rect 1131 3356 1135 3360
rect 1151 3356 1155 3360
rect 1225 3356 1229 3360
rect 1271 3356 1275 3360
rect 1293 3356 1297 3360
rect 1301 3356 1305 3360
rect 1321 3356 1325 3360
rect 1329 3356 1333 3360
rect 1375 3356 1379 3360
rect 1395 3356 1399 3360
rect 1407 3356 1411 3360
rect 1427 3356 1431 3360
rect 1441 3356 1445 3360
rect 1461 3356 1465 3360
rect 1516 3356 1520 3360
rect 1524 3356 1528 3360
rect 1546 3356 1550 3360
rect 1630 3356 1634 3360
rect 1652 3356 1656 3360
rect 1660 3356 1664 3360
rect 1730 3356 1734 3360
rect 1752 3356 1756 3360
rect 1760 3356 1764 3360
rect 1825 3356 1829 3360
rect 1890 3356 1894 3360
rect 1912 3356 1916 3360
rect 1920 3356 1924 3360
rect 1990 3356 1994 3360
rect 2012 3356 2016 3360
rect 2020 3356 2024 3360
rect 2071 3356 2075 3360
rect 2093 3356 2097 3360
rect 2101 3356 2105 3360
rect 2121 3356 2125 3360
rect 2129 3356 2133 3360
rect 2175 3356 2179 3360
rect 2195 3356 2199 3360
rect 2207 3356 2211 3360
rect 2227 3356 2231 3360
rect 2241 3356 2245 3360
rect 2261 3356 2265 3360
rect 2325 3356 2329 3360
rect 2385 3356 2389 3360
rect 2445 3356 2449 3360
rect 2465 3356 2469 3360
rect 2485 3356 2489 3360
rect 2531 3356 2535 3360
rect 2551 3356 2555 3360
rect 2571 3356 2575 3360
rect 2645 3356 2649 3360
rect 2710 3356 2714 3360
rect 2732 3356 2736 3360
rect 2740 3356 2744 3360
rect 2791 3356 2795 3360
rect 2799 3356 2803 3360
rect 2876 3356 2880 3360
rect 2884 3356 2888 3360
rect 2906 3356 2910 3360
rect 2971 3356 2975 3360
rect 2991 3356 2995 3360
rect 3051 3356 3055 3360
rect 3071 3356 3075 3360
rect 3145 3356 3149 3360
rect 3165 3356 3169 3360
rect 3185 3356 3189 3360
rect 3245 3356 3249 3360
rect 3265 3356 3269 3360
rect 3285 3356 3289 3360
rect 3350 3356 3354 3360
rect 3372 3356 3376 3360
rect 3380 3356 3384 3360
rect 3441 3356 3445 3360
rect 3463 3356 3467 3360
rect 3485 3356 3489 3360
rect 3531 3356 3535 3360
rect 3551 3356 3555 3360
rect 3621 3356 3625 3360
rect 3643 3356 3647 3360
rect 3665 3356 3669 3360
rect 3725 3356 3729 3360
rect 3745 3356 3749 3360
rect 3765 3356 3769 3360
rect 3785 3356 3789 3360
rect 3845 3356 3849 3360
rect 3865 3356 3869 3360
rect 3916 3356 3920 3360
rect 3924 3356 3928 3360
rect 3946 3356 3950 3360
rect 4011 3356 4015 3360
rect 4031 3356 4035 3360
rect 4101 3356 4105 3360
rect 4123 3356 4127 3360
rect 4145 3356 4149 3360
rect 4191 3356 4195 3360
rect 4211 3356 4215 3360
rect 4271 3356 4275 3360
rect 4293 3356 4297 3360
rect 4315 3356 4319 3360
rect 4371 3356 4375 3360
rect 4391 3356 4395 3360
rect 4411 3356 4415 3360
rect 4476 3356 4480 3360
rect 4484 3356 4488 3360
rect 4506 3356 4510 3360
rect 4576 3356 4580 3360
rect 4584 3356 4588 3360
rect 4606 3356 4610 3360
rect 4685 3356 4689 3360
rect 4705 3356 4709 3360
rect 4725 3356 4729 3360
rect 35 3233 39 3276
rect 55 3234 59 3316
rect 69 3257 73 3316
rect 89 3276 93 3316
rect 101 3310 105 3316
rect 95 3264 98 3276
rect 69 3249 78 3257
rect 35 3184 39 3221
rect 55 3164 59 3222
rect 74 3220 78 3249
rect 94 3200 98 3264
rect 65 3196 98 3200
rect 65 3164 69 3196
rect 103 3188 107 3298
rect 121 3290 125 3316
rect 167 3312 171 3316
rect 135 3310 171 3312
rect 147 3308 171 3310
rect 89 3176 91 3188
rect 87 3164 91 3176
rect 97 3176 99 3188
rect 97 3164 101 3176
rect 119 3164 123 3278
rect 135 3172 139 3298
rect 175 3284 179 3316
rect 195 3296 199 3336
rect 203 3313 207 3336
rect 203 3306 211 3313
rect 173 3189 179 3284
rect 207 3277 211 3306
rect 203 3271 211 3277
rect 203 3225 207 3271
rect 225 3264 229 3276
rect 227 3252 229 3264
rect 285 3253 289 3276
rect 173 3185 197 3189
rect 159 3180 177 3181
rect 147 3176 177 3180
rect 135 3168 169 3172
rect 165 3164 169 3168
rect 173 3164 177 3176
rect 193 3164 197 3185
rect 203 3164 207 3213
rect 225 3184 229 3252
rect 286 3241 289 3253
rect 280 3193 286 3241
rect 305 3219 309 3276
rect 325 3254 329 3276
rect 345 3254 349 3276
rect 325 3248 338 3254
rect 345 3253 365 3254
rect 345 3248 353 3253
rect 334 3219 338 3248
rect 307 3207 309 3219
rect 305 3205 309 3207
rect 305 3198 318 3205
rect 280 3189 310 3193
rect 306 3184 310 3189
rect 314 3184 318 3198
rect 334 3184 338 3207
rect 353 3199 359 3241
rect 391 3239 395 3316
rect 386 3227 395 3239
rect 389 3211 395 3227
rect 411 3239 415 3316
rect 476 3272 480 3276
rect 462 3264 480 3272
rect 462 3253 466 3264
rect 411 3227 414 3239
rect 411 3211 417 3227
rect 389 3204 397 3211
rect 342 3192 359 3199
rect 342 3184 346 3192
rect 393 3184 397 3204
rect 403 3204 417 3211
rect 403 3184 407 3204
rect 462 3196 466 3241
rect 484 3219 488 3276
rect 506 3273 510 3316
rect 506 3261 513 3273
rect 576 3272 580 3276
rect 562 3264 580 3272
rect 486 3207 495 3219
rect 462 3189 475 3196
rect 471 3184 475 3189
rect 491 3184 495 3207
rect 511 3184 515 3261
rect 562 3253 566 3264
rect 562 3196 566 3241
rect 584 3219 588 3276
rect 606 3273 610 3316
rect 606 3261 613 3273
rect 586 3207 595 3219
rect 562 3189 575 3196
rect 571 3184 575 3189
rect 591 3184 595 3207
rect 611 3184 615 3261
rect 685 3239 689 3316
rect 686 3227 689 3239
rect 683 3211 689 3227
rect 705 3239 709 3316
rect 705 3227 714 3239
rect 751 3233 755 3316
rect 705 3211 711 3227
rect 746 3221 755 3233
rect 683 3204 697 3211
rect 693 3184 697 3204
rect 703 3204 711 3211
rect 703 3184 707 3204
rect 751 3164 755 3221
rect 825 3216 829 3276
rect 845 3216 849 3276
rect 865 3216 869 3276
rect 885 3216 889 3276
rect 905 3216 909 3276
rect 925 3216 929 3276
rect 945 3219 949 3276
rect 965 3219 969 3276
rect 825 3204 838 3216
rect 865 3204 878 3216
rect 905 3204 918 3216
rect 945 3207 954 3219
rect 966 3207 969 3219
rect 825 3184 829 3204
rect 845 3184 849 3204
rect 865 3184 869 3204
rect 885 3184 889 3204
rect 905 3184 909 3204
rect 925 3184 929 3204
rect 945 3184 949 3207
rect 965 3184 969 3207
rect 1011 3219 1015 3276
rect 1031 3219 1035 3276
rect 1011 3207 1014 3219
rect 1026 3207 1035 3219
rect 1051 3216 1055 3276
rect 1071 3216 1075 3276
rect 1091 3216 1095 3276
rect 1111 3216 1115 3276
rect 1131 3216 1135 3276
rect 1151 3216 1155 3276
rect 1011 3184 1015 3207
rect 1031 3184 1035 3207
rect 1062 3204 1075 3216
rect 1102 3204 1115 3216
rect 1142 3204 1155 3216
rect 1051 3184 1055 3204
rect 1071 3184 1075 3204
rect 1091 3184 1095 3204
rect 1111 3184 1115 3204
rect 1131 3184 1135 3204
rect 1151 3184 1155 3204
rect 1225 3233 1229 3316
rect 1293 3313 1297 3336
rect 1289 3306 1297 3313
rect 1289 3277 1293 3306
rect 1301 3296 1305 3336
rect 1321 3284 1325 3316
rect 1329 3312 1333 3316
rect 1329 3310 1365 3312
rect 1329 3308 1353 3310
rect 1271 3264 1275 3276
rect 1289 3271 1297 3277
rect 1271 3252 1273 3264
rect 1225 3221 1234 3233
rect 1225 3164 1229 3221
rect 1271 3184 1275 3252
rect 1293 3225 1297 3271
rect 1293 3164 1297 3213
rect 1321 3189 1327 3284
rect 1303 3185 1327 3189
rect 1303 3164 1307 3185
rect 1323 3180 1341 3181
rect 1323 3176 1353 3180
rect 1323 3164 1327 3176
rect 1361 3172 1365 3298
rect 1375 3290 1379 3316
rect 1395 3310 1399 3316
rect 1331 3168 1365 3172
rect 1331 3164 1335 3168
rect 1377 3164 1381 3278
rect 1393 3188 1397 3298
rect 1407 3276 1411 3316
rect 1402 3264 1405 3276
rect 1402 3200 1406 3264
rect 1427 3257 1431 3316
rect 1422 3249 1431 3257
rect 1422 3220 1426 3249
rect 1441 3234 1445 3316
rect 1461 3233 1465 3276
rect 1516 3272 1520 3276
rect 1502 3264 1520 3272
rect 1502 3253 1506 3264
rect 1402 3196 1435 3200
rect 1401 3176 1403 3188
rect 1399 3164 1403 3176
rect 1409 3176 1411 3188
rect 1409 3164 1413 3176
rect 1431 3164 1435 3196
rect 1441 3164 1445 3222
rect 1461 3184 1465 3221
rect 1502 3196 1506 3241
rect 1524 3219 1528 3276
rect 1546 3273 1550 3316
rect 1630 3273 1634 3316
rect 1546 3261 1553 3273
rect 1627 3261 1634 3273
rect 1526 3207 1535 3219
rect 1502 3189 1515 3196
rect 1511 3184 1515 3189
rect 1531 3184 1535 3207
rect 1551 3184 1555 3261
rect 1625 3184 1629 3261
rect 1652 3219 1656 3276
rect 1660 3272 1664 3276
rect 1730 3273 1734 3316
rect 1660 3264 1678 3272
rect 1674 3253 1678 3264
rect 1727 3261 1734 3273
rect 1645 3207 1654 3219
rect 1645 3184 1649 3207
rect 1674 3196 1678 3241
rect 1665 3189 1678 3196
rect 1665 3184 1669 3189
rect 1725 3184 1729 3261
rect 1752 3219 1756 3276
rect 1760 3272 1764 3276
rect 1760 3264 1778 3272
rect 1774 3253 1778 3264
rect 1745 3207 1754 3219
rect 1745 3184 1749 3207
rect 1774 3196 1778 3241
rect 1765 3189 1778 3196
rect 1825 3233 1829 3316
rect 1890 3273 1894 3316
rect 1887 3261 1894 3273
rect 1825 3221 1834 3233
rect 1765 3184 1769 3189
rect 1825 3164 1829 3221
rect 1885 3184 1889 3261
rect 1912 3219 1916 3276
rect 1920 3272 1924 3276
rect 1990 3273 1994 3316
rect 2093 3313 2097 3336
rect 2089 3306 2097 3313
rect 2089 3277 2093 3306
rect 2101 3296 2105 3336
rect 2121 3284 2125 3316
rect 2129 3312 2133 3316
rect 2129 3310 2165 3312
rect 2129 3308 2153 3310
rect 1920 3264 1938 3272
rect 1934 3253 1938 3264
rect 1987 3261 1994 3273
rect 1905 3207 1914 3219
rect 1905 3184 1909 3207
rect 1934 3196 1938 3241
rect 1925 3189 1938 3196
rect 1925 3184 1929 3189
rect 1985 3184 1989 3261
rect 2012 3219 2016 3276
rect 2020 3272 2024 3276
rect 2020 3264 2038 3272
rect 2034 3253 2038 3264
rect 2071 3264 2075 3276
rect 2089 3271 2097 3277
rect 2071 3252 2073 3264
rect 2005 3207 2014 3219
rect 2005 3184 2009 3207
rect 2034 3196 2038 3241
rect 2025 3189 2038 3196
rect 2025 3184 2029 3189
rect 2071 3184 2075 3252
rect 2093 3225 2097 3271
rect 2093 3164 2097 3213
rect 2121 3189 2127 3284
rect 2103 3185 2127 3189
rect 2103 3164 2107 3185
rect 2123 3180 2141 3181
rect 2123 3176 2153 3180
rect 2123 3164 2127 3176
rect 2161 3172 2165 3298
rect 2175 3290 2179 3316
rect 2195 3310 2199 3316
rect 2131 3168 2165 3172
rect 2131 3164 2135 3168
rect 2177 3164 2181 3278
rect 2193 3188 2197 3298
rect 2207 3276 2211 3316
rect 2202 3264 2205 3276
rect 2202 3200 2206 3264
rect 2227 3257 2231 3316
rect 2222 3249 2231 3257
rect 2222 3220 2226 3249
rect 2241 3234 2245 3316
rect 2261 3233 2265 3276
rect 2325 3233 2329 3316
rect 2385 3233 2389 3316
rect 2445 3273 2449 3316
rect 2465 3304 2469 3316
rect 2485 3308 2489 3316
rect 2485 3304 2500 3308
rect 2465 3300 2480 3304
rect 2474 3293 2480 3300
rect 2445 3261 2453 3273
rect 2465 3261 2472 3273
rect 2202 3196 2235 3200
rect 2201 3176 2203 3188
rect 2199 3164 2203 3176
rect 2209 3176 2211 3188
rect 2209 3164 2213 3176
rect 2231 3164 2235 3196
rect 2241 3164 2245 3222
rect 2325 3221 2334 3233
rect 2385 3221 2394 3233
rect 2261 3184 2265 3221
rect 2325 3164 2329 3221
rect 2385 3164 2389 3221
rect 2468 3204 2472 3261
rect 2476 3204 2480 3281
rect 2494 3273 2500 3304
rect 2484 3261 2494 3273
rect 2531 3262 2535 3276
rect 2551 3262 2555 3276
rect 2484 3204 2488 3261
rect 2519 3256 2535 3262
rect 2540 3256 2555 3262
rect 2519 3219 2526 3256
rect 2540 3233 2546 3256
rect 2519 3194 2526 3207
rect 2519 3188 2538 3194
rect 2534 3184 2538 3188
rect 2542 3184 2546 3221
rect 2571 3219 2575 3276
rect 2566 3207 2575 3219
rect 2645 3233 2649 3316
rect 2710 3273 2714 3316
rect 2707 3261 2714 3273
rect 2645 3221 2654 3233
rect 2564 3164 2568 3207
rect 2645 3164 2649 3221
rect 2705 3184 2709 3261
rect 2732 3219 2736 3276
rect 2740 3272 2744 3276
rect 2740 3264 2758 3272
rect 2754 3253 2758 3264
rect 2791 3253 2795 3276
rect 2786 3241 2795 3253
rect 2799 3253 2803 3276
rect 2876 3272 2880 3276
rect 2862 3264 2880 3272
rect 2862 3253 2866 3264
rect 2799 3241 2814 3253
rect 2725 3207 2734 3219
rect 2725 3184 2729 3207
rect 2754 3196 2758 3241
rect 2745 3189 2758 3196
rect 2745 3184 2749 3189
rect 2791 3164 2795 3241
rect 2811 3164 2815 3241
rect 2862 3196 2866 3241
rect 2884 3219 2888 3276
rect 2906 3273 2910 3316
rect 2906 3261 2913 3273
rect 2886 3207 2895 3219
rect 2862 3189 2875 3196
rect 2871 3184 2875 3189
rect 2891 3184 2895 3207
rect 2911 3184 2915 3261
rect 2971 3239 2975 3316
rect 2966 3227 2975 3239
rect 2969 3211 2975 3227
rect 2991 3239 2995 3316
rect 3051 3239 3055 3316
rect 2991 3227 2994 3239
rect 3046 3227 3055 3239
rect 2991 3211 2997 3227
rect 2969 3204 2977 3211
rect 2973 3184 2977 3204
rect 2983 3204 2997 3211
rect 3049 3211 3055 3227
rect 3071 3239 3075 3316
rect 3071 3227 3074 3239
rect 3071 3211 3077 3227
rect 3049 3204 3057 3211
rect 2983 3184 2987 3204
rect 3053 3184 3057 3204
rect 3063 3204 3077 3211
rect 3145 3219 3149 3276
rect 3165 3262 3169 3276
rect 3185 3262 3189 3276
rect 3245 3273 3249 3316
rect 3265 3304 3269 3316
rect 3285 3308 3289 3316
rect 3285 3304 3300 3308
rect 3265 3300 3280 3304
rect 3274 3293 3280 3300
rect 3165 3256 3180 3262
rect 3185 3256 3201 3262
rect 3245 3261 3253 3273
rect 3265 3261 3272 3273
rect 3174 3233 3180 3256
rect 3145 3207 3154 3219
rect 3063 3184 3067 3204
rect 3152 3164 3156 3207
rect 3174 3184 3178 3221
rect 3194 3219 3201 3256
rect 3194 3194 3201 3207
rect 3268 3204 3272 3261
rect 3276 3204 3280 3281
rect 3294 3273 3300 3304
rect 3350 3273 3354 3316
rect 3284 3261 3294 3273
rect 3347 3261 3354 3273
rect 3284 3204 3288 3261
rect 3182 3188 3201 3194
rect 3182 3184 3186 3188
rect 3345 3184 3349 3261
rect 3372 3219 3376 3276
rect 3380 3272 3384 3276
rect 3380 3264 3398 3272
rect 3394 3253 3398 3264
rect 3365 3207 3374 3219
rect 3365 3184 3369 3207
rect 3394 3196 3398 3241
rect 3385 3189 3398 3196
rect 3441 3202 3445 3276
rect 3463 3239 3467 3316
rect 3485 3253 3489 3316
rect 3485 3241 3494 3253
rect 3466 3227 3479 3239
rect 3441 3190 3453 3202
rect 3385 3184 3389 3189
rect 3455 3184 3459 3190
rect 3475 3184 3479 3227
rect 3485 3184 3489 3241
rect 3531 3239 3535 3316
rect 3526 3227 3535 3239
rect 3529 3211 3535 3227
rect 3551 3239 3555 3316
rect 3551 3227 3554 3239
rect 3551 3211 3557 3227
rect 3529 3204 3537 3211
rect 3533 3184 3537 3204
rect 3543 3204 3557 3211
rect 3543 3184 3547 3204
rect 3621 3202 3625 3276
rect 3643 3239 3647 3316
rect 3665 3253 3669 3316
rect 3725 3253 3729 3276
rect 3665 3241 3674 3253
rect 3726 3241 3729 3253
rect 3646 3227 3659 3239
rect 3621 3190 3633 3202
rect 3635 3184 3639 3190
rect 3655 3184 3659 3227
rect 3665 3184 3669 3241
rect 3720 3193 3726 3241
rect 3745 3219 3749 3276
rect 3765 3254 3769 3276
rect 3785 3254 3789 3276
rect 3765 3248 3778 3254
rect 3785 3253 3805 3254
rect 3785 3248 3793 3253
rect 3774 3219 3778 3248
rect 3747 3207 3749 3219
rect 3745 3205 3749 3207
rect 3745 3198 3758 3205
rect 3720 3189 3750 3193
rect 3746 3184 3750 3189
rect 3754 3184 3758 3198
rect 3774 3184 3778 3207
rect 3793 3199 3799 3241
rect 3845 3239 3849 3316
rect 3846 3227 3849 3239
rect 3843 3211 3849 3227
rect 3865 3239 3869 3316
rect 3916 3272 3920 3276
rect 3902 3264 3920 3272
rect 3902 3253 3906 3264
rect 3865 3227 3874 3239
rect 3865 3211 3871 3227
rect 3843 3204 3857 3211
rect 3782 3192 3799 3199
rect 3782 3184 3786 3192
rect 3853 3184 3857 3204
rect 3863 3204 3871 3211
rect 3863 3184 3867 3204
rect 3902 3196 3906 3241
rect 3924 3219 3928 3276
rect 3946 3273 3950 3316
rect 3946 3261 3953 3273
rect 3926 3207 3935 3219
rect 3902 3189 3915 3196
rect 3911 3184 3915 3189
rect 3931 3184 3935 3207
rect 3951 3184 3955 3261
rect 4011 3239 4015 3316
rect 4006 3227 4015 3239
rect 4009 3211 4015 3227
rect 4031 3239 4035 3316
rect 4031 3227 4034 3239
rect 4031 3211 4037 3227
rect 4009 3204 4017 3211
rect 4013 3184 4017 3204
rect 4023 3204 4037 3211
rect 4023 3184 4027 3204
rect 4101 3202 4105 3276
rect 4123 3239 4127 3316
rect 4145 3253 4149 3316
rect 4145 3241 4154 3253
rect 4126 3227 4139 3239
rect 4101 3190 4113 3202
rect 4115 3184 4119 3190
rect 4135 3184 4139 3227
rect 4145 3184 4149 3241
rect 4191 3239 4195 3316
rect 4186 3227 4195 3239
rect 4189 3211 4195 3227
rect 4211 3239 4215 3316
rect 4271 3253 4275 3316
rect 4266 3241 4275 3253
rect 4211 3227 4214 3239
rect 4211 3211 4217 3227
rect 4189 3204 4197 3211
rect 4193 3184 4197 3204
rect 4203 3204 4217 3211
rect 4203 3184 4207 3204
rect 4271 3184 4275 3241
rect 4293 3239 4297 3316
rect 4281 3227 4294 3239
rect 4281 3184 4285 3227
rect 4315 3202 4319 3276
rect 4371 3262 4375 3276
rect 4391 3262 4395 3276
rect 4359 3256 4375 3262
rect 4380 3256 4395 3262
rect 4359 3219 4366 3256
rect 4380 3233 4386 3256
rect 4307 3190 4319 3202
rect 4359 3194 4366 3207
rect 4301 3184 4305 3190
rect 4359 3188 4378 3194
rect 4374 3184 4378 3188
rect 4382 3184 4386 3221
rect 4411 3219 4415 3276
rect 4476 3272 4480 3276
rect 4462 3264 4480 3272
rect 4462 3253 4466 3264
rect 4406 3207 4415 3219
rect 4404 3164 4408 3207
rect 4462 3196 4466 3241
rect 4484 3219 4488 3276
rect 4506 3273 4510 3316
rect 4506 3261 4513 3273
rect 4576 3272 4580 3276
rect 4562 3264 4580 3272
rect 4486 3207 4495 3219
rect 4462 3189 4475 3196
rect 4471 3184 4475 3189
rect 4491 3184 4495 3207
rect 4511 3184 4515 3261
rect 4562 3253 4566 3264
rect 4562 3196 4566 3241
rect 4584 3219 4588 3276
rect 4606 3273 4610 3316
rect 4685 3273 4689 3316
rect 4705 3304 4709 3316
rect 4725 3308 4729 3316
rect 4725 3304 4740 3308
rect 4705 3300 4720 3304
rect 4714 3293 4720 3300
rect 4606 3261 4613 3273
rect 4685 3261 4693 3273
rect 4705 3261 4712 3273
rect 4586 3207 4595 3219
rect 4562 3189 4575 3196
rect 4571 3184 4575 3189
rect 4591 3184 4595 3207
rect 4611 3184 4615 3261
rect 4708 3204 4712 3261
rect 4716 3204 4720 3281
rect 4734 3273 4740 3304
rect 4724 3261 4734 3273
rect 4724 3204 4728 3261
rect 35 3140 39 3144
rect 55 3140 59 3144
rect 65 3140 69 3144
rect 87 3140 91 3144
rect 97 3140 101 3144
rect 119 3140 123 3144
rect 165 3140 169 3144
rect 173 3140 177 3144
rect 193 3140 197 3144
rect 203 3140 207 3144
rect 225 3140 229 3144
rect 306 3140 310 3144
rect 314 3140 318 3144
rect 334 3140 338 3144
rect 342 3140 346 3144
rect 393 3140 397 3144
rect 403 3140 407 3144
rect 471 3140 475 3144
rect 491 3140 495 3144
rect 511 3140 515 3144
rect 571 3140 575 3144
rect 591 3140 595 3144
rect 611 3140 615 3144
rect 693 3140 697 3144
rect 703 3140 707 3144
rect 751 3140 755 3144
rect 825 3140 829 3144
rect 845 3140 849 3144
rect 865 3140 869 3144
rect 885 3140 889 3144
rect 905 3140 909 3144
rect 925 3140 929 3144
rect 945 3140 949 3144
rect 965 3140 969 3144
rect 1011 3140 1015 3144
rect 1031 3140 1035 3144
rect 1051 3140 1055 3144
rect 1071 3140 1075 3144
rect 1091 3140 1095 3144
rect 1111 3140 1115 3144
rect 1131 3140 1135 3144
rect 1151 3140 1155 3144
rect 1225 3140 1229 3144
rect 1271 3140 1275 3144
rect 1293 3140 1297 3144
rect 1303 3140 1307 3144
rect 1323 3140 1327 3144
rect 1331 3140 1335 3144
rect 1377 3140 1381 3144
rect 1399 3140 1403 3144
rect 1409 3140 1413 3144
rect 1431 3140 1435 3144
rect 1441 3140 1445 3144
rect 1461 3140 1465 3144
rect 1511 3140 1515 3144
rect 1531 3140 1535 3144
rect 1551 3140 1555 3144
rect 1625 3140 1629 3144
rect 1645 3140 1649 3144
rect 1665 3140 1669 3144
rect 1725 3140 1729 3144
rect 1745 3140 1749 3144
rect 1765 3140 1769 3144
rect 1825 3140 1829 3144
rect 1885 3140 1889 3144
rect 1905 3140 1909 3144
rect 1925 3140 1929 3144
rect 1985 3140 1989 3144
rect 2005 3140 2009 3144
rect 2025 3140 2029 3144
rect 2071 3140 2075 3144
rect 2093 3140 2097 3144
rect 2103 3140 2107 3144
rect 2123 3140 2127 3144
rect 2131 3140 2135 3144
rect 2177 3140 2181 3144
rect 2199 3140 2203 3144
rect 2209 3140 2213 3144
rect 2231 3140 2235 3144
rect 2241 3140 2245 3144
rect 2261 3140 2265 3144
rect 2325 3140 2329 3144
rect 2385 3140 2389 3144
rect 2468 3140 2472 3144
rect 2476 3140 2480 3144
rect 2484 3140 2488 3144
rect 2534 3140 2538 3144
rect 2542 3140 2546 3144
rect 2564 3140 2568 3144
rect 2645 3140 2649 3144
rect 2705 3140 2709 3144
rect 2725 3140 2729 3144
rect 2745 3140 2749 3144
rect 2791 3140 2795 3144
rect 2811 3140 2815 3144
rect 2871 3140 2875 3144
rect 2891 3140 2895 3144
rect 2911 3140 2915 3144
rect 2973 3140 2977 3144
rect 2983 3140 2987 3144
rect 3053 3140 3057 3144
rect 3063 3140 3067 3144
rect 3152 3140 3156 3144
rect 3174 3140 3178 3144
rect 3182 3140 3186 3144
rect 3268 3140 3272 3144
rect 3276 3140 3280 3144
rect 3284 3140 3288 3144
rect 3345 3140 3349 3144
rect 3365 3140 3369 3144
rect 3385 3140 3389 3144
rect 3455 3140 3459 3144
rect 3475 3140 3479 3144
rect 3485 3140 3489 3144
rect 3533 3140 3537 3144
rect 3543 3140 3547 3144
rect 3635 3140 3639 3144
rect 3655 3140 3659 3144
rect 3665 3140 3669 3144
rect 3746 3140 3750 3144
rect 3754 3140 3758 3144
rect 3774 3140 3778 3144
rect 3782 3140 3786 3144
rect 3853 3140 3857 3144
rect 3863 3140 3867 3144
rect 3911 3140 3915 3144
rect 3931 3140 3935 3144
rect 3951 3140 3955 3144
rect 4013 3140 4017 3144
rect 4023 3140 4027 3144
rect 4115 3140 4119 3144
rect 4135 3140 4139 3144
rect 4145 3140 4149 3144
rect 4193 3140 4197 3144
rect 4203 3140 4207 3144
rect 4271 3140 4275 3144
rect 4281 3140 4285 3144
rect 4301 3140 4305 3144
rect 4374 3140 4378 3144
rect 4382 3140 4386 3144
rect 4404 3140 4408 3144
rect 4471 3140 4475 3144
rect 4491 3140 4495 3144
rect 4511 3140 4515 3144
rect 4571 3140 4575 3144
rect 4591 3140 4595 3144
rect 4611 3140 4615 3144
rect 4708 3140 4712 3144
rect 4716 3140 4720 3144
rect 4724 3140 4728 3144
rect 35 3116 39 3120
rect 55 3116 59 3120
rect 65 3116 69 3120
rect 87 3116 91 3120
rect 97 3116 101 3120
rect 119 3116 123 3120
rect 165 3116 169 3120
rect 173 3116 177 3120
rect 193 3116 197 3120
rect 203 3116 207 3120
rect 225 3116 229 3120
rect 285 3116 289 3120
rect 305 3116 309 3120
rect 325 3116 329 3120
rect 393 3116 397 3120
rect 403 3116 407 3120
rect 451 3116 455 3120
rect 473 3116 477 3120
rect 483 3116 487 3120
rect 503 3116 507 3120
rect 511 3116 515 3120
rect 557 3116 561 3120
rect 579 3116 583 3120
rect 589 3116 593 3120
rect 611 3116 615 3120
rect 621 3116 625 3120
rect 641 3116 645 3120
rect 695 3116 699 3120
rect 715 3116 719 3120
rect 725 3116 729 3120
rect 747 3116 751 3120
rect 757 3116 761 3120
rect 779 3116 783 3120
rect 825 3116 829 3120
rect 833 3116 837 3120
rect 853 3116 857 3120
rect 863 3116 867 3120
rect 885 3116 889 3120
rect 931 3116 935 3120
rect 1005 3116 1009 3120
rect 1025 3116 1029 3120
rect 1093 3116 1097 3120
rect 1103 3116 1107 3120
rect 1151 3116 1155 3120
rect 1171 3116 1175 3120
rect 1191 3116 1195 3120
rect 1254 3116 1258 3120
rect 1262 3116 1266 3120
rect 1284 3116 1288 3120
rect 1355 3116 1359 3120
rect 1375 3116 1379 3120
rect 1385 3116 1389 3120
rect 1407 3116 1411 3120
rect 1417 3116 1421 3120
rect 1439 3116 1443 3120
rect 1485 3116 1489 3120
rect 1493 3116 1497 3120
rect 1513 3116 1517 3120
rect 1523 3116 1527 3120
rect 1545 3116 1549 3120
rect 1605 3116 1609 3120
rect 1625 3116 1629 3120
rect 1693 3116 1697 3120
rect 1703 3116 1707 3120
rect 1751 3116 1755 3120
rect 1771 3116 1775 3120
rect 1791 3116 1795 3120
rect 1865 3116 1869 3120
rect 1885 3116 1889 3120
rect 1905 3116 1909 3120
rect 1951 3116 1955 3120
rect 1973 3116 1977 3120
rect 1983 3116 1987 3120
rect 2003 3116 2007 3120
rect 2011 3116 2015 3120
rect 2057 3116 2061 3120
rect 2079 3116 2083 3120
rect 2089 3116 2093 3120
rect 2111 3116 2115 3120
rect 2121 3116 2125 3120
rect 2141 3116 2145 3120
rect 2205 3116 2209 3120
rect 2225 3116 2229 3120
rect 2285 3116 2289 3120
rect 2368 3116 2372 3120
rect 2376 3116 2380 3120
rect 2384 3116 2388 3120
rect 2452 3116 2456 3120
rect 2474 3116 2478 3120
rect 2482 3116 2486 3120
rect 2568 3116 2572 3120
rect 2576 3116 2580 3120
rect 2584 3116 2588 3120
rect 2645 3116 2649 3120
rect 2665 3116 2669 3120
rect 2685 3116 2689 3120
rect 2745 3116 2749 3120
rect 2765 3116 2769 3120
rect 2813 3116 2817 3120
rect 2823 3116 2827 3120
rect 2893 3116 2897 3120
rect 2903 3116 2907 3120
rect 2974 3116 2978 3120
rect 2982 3116 2986 3120
rect 3002 3116 3006 3120
rect 3010 3116 3014 3120
rect 3093 3116 3097 3120
rect 3103 3116 3107 3120
rect 3171 3116 3175 3120
rect 3191 3116 3195 3120
rect 3211 3116 3215 3120
rect 3271 3116 3275 3120
rect 3331 3116 3335 3120
rect 3341 3116 3345 3120
rect 3361 3116 3365 3120
rect 3443 3116 3447 3120
rect 3465 3116 3469 3120
rect 3523 3116 3527 3120
rect 3545 3116 3549 3120
rect 3593 3116 3597 3120
rect 3603 3116 3607 3120
rect 3671 3116 3675 3120
rect 3691 3116 3695 3120
rect 3711 3116 3715 3120
rect 3783 3116 3787 3120
rect 3805 3116 3809 3120
rect 3851 3116 3855 3120
rect 3871 3116 3875 3120
rect 3891 3116 3895 3120
rect 3952 3116 3956 3120
rect 3960 3116 3964 3120
rect 3968 3116 3972 3120
rect 4051 3116 4055 3120
rect 4073 3116 4077 3120
rect 4152 3116 4156 3120
rect 4174 3116 4178 3120
rect 4182 3116 4186 3120
rect 4232 3116 4236 3120
rect 4240 3116 4244 3120
rect 4248 3116 4252 3120
rect 4352 3116 4356 3120
rect 4374 3116 4378 3120
rect 4382 3116 4386 3120
rect 4468 3116 4472 3120
rect 4476 3116 4480 3120
rect 4484 3116 4488 3120
rect 4545 3116 4549 3120
rect 4605 3116 4609 3120
rect 4625 3116 4629 3120
rect 4645 3116 4649 3120
rect 4691 3116 4695 3120
rect 4711 3116 4715 3120
rect 4731 3116 4735 3120
rect 35 3039 39 3076
rect 55 3038 59 3096
rect 65 3064 69 3096
rect 87 3084 91 3096
rect 89 3072 91 3084
rect 97 3084 101 3096
rect 97 3072 99 3084
rect 65 3060 98 3064
rect 35 2984 39 3027
rect 55 2944 59 3026
rect 74 3011 78 3040
rect 69 3003 78 3011
rect 69 2944 73 3003
rect 94 2996 98 3060
rect 95 2984 98 2996
rect 89 2944 93 2984
rect 103 2962 107 3072
rect 119 2982 123 3096
rect 165 3092 169 3096
rect 135 3088 169 3092
rect 101 2944 105 2950
rect 121 2944 125 2970
rect 135 2962 139 3088
rect 173 3084 177 3096
rect 147 3080 177 3084
rect 159 3079 177 3080
rect 193 3075 197 3096
rect 173 3071 197 3075
rect 173 2976 179 3071
rect 203 3047 207 3096
rect 203 2989 207 3035
rect 225 3008 229 3076
rect 227 2996 229 3008
rect 285 2999 289 3076
rect 305 3053 309 3076
rect 325 3071 329 3076
rect 325 3064 338 3071
rect 305 3041 314 3053
rect 203 2983 211 2989
rect 225 2984 229 2996
rect 287 2987 294 2999
rect 147 2950 171 2952
rect 135 2948 171 2950
rect 167 2944 171 2948
rect 175 2944 179 2976
rect 195 2924 199 2964
rect 207 2954 211 2983
rect 203 2947 211 2954
rect 203 2924 207 2947
rect 290 2944 294 2987
rect 312 2984 316 3041
rect 334 3019 338 3064
rect 393 3056 397 3076
rect 383 3049 397 3056
rect 403 3056 407 3076
rect 403 3049 411 3056
rect 383 3033 389 3049
rect 386 3021 389 3033
rect 334 2996 338 3007
rect 320 2988 338 2996
rect 320 2984 324 2988
rect 385 2944 389 3021
rect 405 3033 411 3049
rect 405 3021 414 3033
rect 405 2944 409 3021
rect 451 3008 455 3076
rect 473 3047 477 3096
rect 483 3075 487 3096
rect 503 3084 507 3096
rect 511 3092 515 3096
rect 511 3088 545 3092
rect 503 3080 533 3084
rect 503 3079 521 3080
rect 483 3071 507 3075
rect 451 2996 453 3008
rect 451 2984 455 2996
rect 473 2989 477 3035
rect 469 2983 477 2989
rect 469 2954 473 2983
rect 501 2976 507 3071
rect 469 2947 477 2954
rect 473 2924 477 2947
rect 481 2924 485 2964
rect 501 2944 505 2976
rect 541 2962 545 3088
rect 557 2982 561 3096
rect 579 3084 583 3096
rect 581 3072 583 3084
rect 589 3084 593 3096
rect 589 3072 591 3084
rect 509 2950 533 2952
rect 509 2948 545 2950
rect 509 2944 513 2948
rect 555 2944 559 2970
rect 573 2962 577 3072
rect 611 3064 615 3096
rect 582 3060 615 3064
rect 582 2996 586 3060
rect 602 3011 606 3040
rect 621 3038 625 3096
rect 641 3039 645 3076
rect 695 3039 699 3076
rect 715 3038 719 3096
rect 725 3064 729 3096
rect 747 3084 751 3096
rect 749 3072 751 3084
rect 757 3084 761 3096
rect 757 3072 759 3084
rect 725 3060 758 3064
rect 602 3003 611 3011
rect 582 2984 585 2996
rect 575 2944 579 2950
rect 587 2944 591 2984
rect 607 2944 611 3003
rect 621 2944 625 3026
rect 641 2984 645 3027
rect 695 2984 699 3027
rect 715 2944 719 3026
rect 734 3011 738 3040
rect 729 3003 738 3011
rect 729 2944 733 3003
rect 754 2996 758 3060
rect 755 2984 758 2996
rect 749 2944 753 2984
rect 763 2962 767 3072
rect 779 2982 783 3096
rect 825 3092 829 3096
rect 795 3088 829 3092
rect 761 2944 765 2950
rect 781 2944 785 2970
rect 795 2962 799 3088
rect 833 3084 837 3096
rect 807 3080 837 3084
rect 819 3079 837 3080
rect 853 3075 857 3096
rect 833 3071 857 3075
rect 833 2976 839 3071
rect 863 3047 867 3096
rect 863 2989 867 3035
rect 885 3008 889 3076
rect 931 3039 935 3096
rect 926 3027 935 3039
rect 887 2996 889 3008
rect 863 2983 871 2989
rect 885 2984 889 2996
rect 807 2950 831 2952
rect 795 2948 831 2950
rect 827 2944 831 2948
rect 835 2944 839 2976
rect 855 2924 859 2964
rect 867 2954 871 2983
rect 863 2947 871 2954
rect 863 2924 867 2947
rect 931 2944 935 3027
rect 1005 3019 1009 3096
rect 1025 3019 1029 3096
rect 1093 3056 1097 3076
rect 1083 3049 1097 3056
rect 1103 3056 1107 3076
rect 1151 3071 1155 3076
rect 1142 3064 1155 3071
rect 1103 3049 1111 3056
rect 1083 3033 1089 3049
rect 1086 3021 1089 3033
rect 1006 3007 1021 3019
rect 1017 2984 1021 3007
rect 1025 3007 1034 3019
rect 1025 2984 1029 3007
rect 1085 2944 1089 3021
rect 1105 3033 1111 3049
rect 1105 3021 1114 3033
rect 1105 2944 1109 3021
rect 1142 3019 1146 3064
rect 1171 3053 1175 3076
rect 1166 3041 1175 3053
rect 1142 2996 1146 3007
rect 1142 2988 1160 2996
rect 1156 2984 1160 2988
rect 1164 2984 1168 3041
rect 1191 2999 1195 3076
rect 1254 3072 1258 3076
rect 1239 3066 1258 3072
rect 1239 3053 1246 3066
rect 1239 3004 1246 3041
rect 1262 3039 1266 3076
rect 1284 3053 1288 3096
rect 1286 3041 1295 3053
rect 1260 3004 1266 3027
rect 1186 2987 1193 2999
rect 1239 2998 1255 3004
rect 1260 2998 1275 3004
rect 1186 2944 1190 2987
rect 1251 2984 1255 2998
rect 1271 2984 1275 2998
rect 1291 2984 1295 3041
rect 1355 3039 1359 3076
rect 1375 3038 1379 3096
rect 1385 3064 1389 3096
rect 1407 3084 1411 3096
rect 1409 3072 1411 3084
rect 1417 3084 1421 3096
rect 1417 3072 1419 3084
rect 1385 3060 1418 3064
rect 1355 2984 1359 3027
rect 1375 2944 1379 3026
rect 1394 3011 1398 3040
rect 1389 3003 1398 3011
rect 1389 2944 1393 3003
rect 1414 2996 1418 3060
rect 1415 2984 1418 2996
rect 1409 2944 1413 2984
rect 1423 2962 1427 3072
rect 1439 2982 1443 3096
rect 1485 3092 1489 3096
rect 1455 3088 1489 3092
rect 1421 2944 1425 2950
rect 1441 2944 1445 2970
rect 1455 2962 1459 3088
rect 1493 3084 1497 3096
rect 1467 3080 1497 3084
rect 1479 3079 1497 3080
rect 1513 3075 1517 3096
rect 1493 3071 1517 3075
rect 1493 2976 1499 3071
rect 1523 3047 1527 3096
rect 1523 2989 1527 3035
rect 1545 3008 1549 3076
rect 1605 3019 1609 3096
rect 1625 3019 1629 3096
rect 1693 3056 1697 3076
rect 1683 3049 1697 3056
rect 1703 3056 1707 3076
rect 1751 3071 1755 3076
rect 1742 3064 1755 3071
rect 1703 3049 1711 3056
rect 1683 3033 1689 3049
rect 1686 3021 1689 3033
rect 1547 2996 1549 3008
rect 1606 3007 1621 3019
rect 1523 2983 1531 2989
rect 1545 2984 1549 2996
rect 1617 2984 1621 3007
rect 1625 3007 1634 3019
rect 1625 2984 1629 3007
rect 1467 2950 1491 2952
rect 1455 2948 1491 2950
rect 1487 2944 1491 2948
rect 1495 2944 1499 2976
rect 1515 2924 1519 2964
rect 1527 2954 1531 2983
rect 1523 2947 1531 2954
rect 1523 2924 1527 2947
rect 1685 2944 1689 3021
rect 1705 3033 1711 3049
rect 1705 3021 1714 3033
rect 1705 2944 1709 3021
rect 1742 3019 1746 3064
rect 1771 3053 1775 3076
rect 1766 3041 1775 3053
rect 1742 2996 1746 3007
rect 1742 2988 1760 2996
rect 1756 2984 1760 2988
rect 1764 2984 1768 3041
rect 1791 2999 1795 3076
rect 1865 2999 1869 3076
rect 1885 3053 1889 3076
rect 1905 3071 1909 3076
rect 1905 3064 1918 3071
rect 1885 3041 1894 3053
rect 1786 2987 1793 2999
rect 1867 2987 1874 2999
rect 1786 2944 1790 2987
rect 1870 2944 1874 2987
rect 1892 2984 1896 3041
rect 1914 3019 1918 3064
rect 1951 3008 1955 3076
rect 1973 3047 1977 3096
rect 1983 3075 1987 3096
rect 2003 3084 2007 3096
rect 2011 3092 2015 3096
rect 2011 3088 2045 3092
rect 2003 3080 2033 3084
rect 2003 3079 2021 3080
rect 1983 3071 2007 3075
rect 1914 2996 1918 3007
rect 1900 2988 1918 2996
rect 1951 2996 1953 3008
rect 1900 2984 1904 2988
rect 1951 2984 1955 2996
rect 1973 2989 1977 3035
rect 1969 2983 1977 2989
rect 1969 2954 1973 2983
rect 2001 2976 2007 3071
rect 1969 2947 1977 2954
rect 1973 2924 1977 2947
rect 1981 2924 1985 2964
rect 2001 2944 2005 2976
rect 2041 2962 2045 3088
rect 2057 2982 2061 3096
rect 2079 3084 2083 3096
rect 2081 3072 2083 3084
rect 2089 3084 2093 3096
rect 2089 3072 2091 3084
rect 2009 2950 2033 2952
rect 2009 2948 2045 2950
rect 2009 2944 2013 2948
rect 2055 2944 2059 2970
rect 2073 2962 2077 3072
rect 2111 3064 2115 3096
rect 2082 3060 2115 3064
rect 2082 2996 2086 3060
rect 2102 3011 2106 3040
rect 2121 3038 2125 3096
rect 2141 3039 2145 3076
rect 2102 3003 2111 3011
rect 2082 2984 2085 2996
rect 2075 2944 2079 2950
rect 2087 2944 2091 2984
rect 2107 2944 2111 3003
rect 2121 2944 2125 3026
rect 2141 2984 2145 3027
rect 2205 3019 2209 3096
rect 2225 3019 2229 3096
rect 2285 3039 2289 3096
rect 2285 3027 2294 3039
rect 2206 3007 2221 3019
rect 2217 2984 2221 3007
rect 2225 3007 2234 3019
rect 2225 2984 2229 3007
rect 2285 2944 2289 3027
rect 2368 2999 2372 3056
rect 2345 2987 2353 2999
rect 2365 2987 2372 2999
rect 2345 2944 2349 2987
rect 2376 2979 2380 3056
rect 2384 2999 2388 3056
rect 2452 3053 2456 3096
rect 2445 3041 2454 3053
rect 2384 2987 2394 2999
rect 2374 2960 2380 2967
rect 2365 2956 2380 2960
rect 2394 2956 2400 2987
rect 2445 2984 2449 3041
rect 2474 3039 2478 3076
rect 2482 3072 2486 3076
rect 2482 3066 2501 3072
rect 2494 3053 2501 3066
rect 2474 3004 2480 3027
rect 2494 3004 2501 3041
rect 2465 2998 2480 3004
rect 2485 2998 2501 3004
rect 2568 2999 2572 3056
rect 2465 2984 2469 2998
rect 2485 2984 2489 2998
rect 2545 2987 2553 2999
rect 2565 2987 2572 2999
rect 2365 2944 2369 2956
rect 2385 2952 2400 2956
rect 2385 2944 2389 2952
rect 2545 2944 2549 2987
rect 2576 2979 2580 3056
rect 2584 2999 2588 3056
rect 2645 2999 2649 3076
rect 2665 3053 2669 3076
rect 2685 3071 2689 3076
rect 2685 3064 2698 3071
rect 2665 3041 2674 3053
rect 2584 2987 2594 2999
rect 2647 2987 2654 2999
rect 2574 2960 2580 2967
rect 2565 2956 2580 2960
rect 2594 2956 2600 2987
rect 2565 2944 2569 2956
rect 2585 2952 2600 2956
rect 2585 2944 2589 2952
rect 2650 2944 2654 2987
rect 2672 2984 2676 3041
rect 2694 3019 2698 3064
rect 2745 3019 2749 3096
rect 2765 3019 2769 3096
rect 2813 3056 2817 3076
rect 2809 3049 2817 3056
rect 2823 3056 2827 3076
rect 2893 3056 2897 3076
rect 2823 3049 2837 3056
rect 2809 3033 2815 3049
rect 2806 3021 2815 3033
rect 2746 3007 2761 3019
rect 2694 2996 2698 3007
rect 2680 2988 2698 2996
rect 2680 2984 2684 2988
rect 2757 2984 2761 3007
rect 2765 3007 2774 3019
rect 2765 2984 2769 3007
rect 2811 2944 2815 3021
rect 2831 3033 2837 3049
rect 2889 3049 2897 3056
rect 2903 3056 2907 3076
rect 2974 3068 2978 3076
rect 2961 3061 2978 3068
rect 2903 3049 2917 3056
rect 2889 3033 2895 3049
rect 2831 3021 2834 3033
rect 2886 3021 2895 3033
rect 2831 2944 2835 3021
rect 2891 2944 2895 3021
rect 2911 3033 2917 3049
rect 2911 3021 2914 3033
rect 2911 2944 2915 3021
rect 2961 3019 2967 3061
rect 2982 3053 2986 3076
rect 3002 3062 3006 3076
rect 3010 3071 3014 3076
rect 3010 3067 3040 3071
rect 3002 3055 3015 3062
rect 3011 3053 3015 3055
rect 3011 3041 3013 3053
rect 2982 3012 2986 3041
rect 2967 3007 2975 3012
rect 2955 3006 2975 3007
rect 2982 3006 2995 3012
rect 2971 2984 2975 3006
rect 2991 2984 2995 3006
rect 3011 2984 3015 3041
rect 3034 3019 3040 3067
rect 3093 3056 3097 3076
rect 3089 3049 3097 3056
rect 3103 3056 3107 3076
rect 3171 3071 3175 3076
rect 3162 3064 3175 3071
rect 3103 3049 3117 3056
rect 3089 3033 3095 3049
rect 3086 3021 3095 3033
rect 3031 3007 3034 3019
rect 3031 2984 3035 3007
rect 3091 2944 3095 3021
rect 3111 3033 3117 3049
rect 3111 3021 3114 3033
rect 3111 2944 3115 3021
rect 3162 3019 3166 3064
rect 3191 3053 3195 3076
rect 3186 3041 3195 3053
rect 3162 2996 3166 3007
rect 3162 2988 3180 2996
rect 3176 2984 3180 2988
rect 3184 2984 3188 3041
rect 3211 2999 3215 3076
rect 3271 3053 3275 3076
rect 3266 3041 3275 3053
rect 3206 2987 3213 2999
rect 3206 2944 3210 2987
rect 3271 2984 3275 3041
rect 3331 3019 3335 3076
rect 3341 3033 3345 3076
rect 3361 3070 3365 3076
rect 3443 3070 3447 3076
rect 3367 3058 3379 3070
rect 3443 3058 3445 3070
rect 3341 3021 3354 3033
rect 3326 3007 3335 3019
rect 3331 2944 3335 3007
rect 3353 2944 3357 3021
rect 3375 2984 3379 3058
rect 3465 3019 3469 3096
rect 3523 3070 3527 3076
rect 3523 3058 3525 3070
rect 3545 3019 3549 3096
rect 3593 3056 3597 3076
rect 3589 3049 3597 3056
rect 3603 3056 3607 3076
rect 3671 3071 3675 3076
rect 3662 3064 3675 3071
rect 3603 3049 3617 3056
rect 3589 3033 3595 3049
rect 3586 3021 3595 3033
rect 3465 3007 3474 3019
rect 3545 3007 3554 3019
rect 3443 2990 3445 3002
rect 3443 2984 3447 2990
rect 3465 2944 3469 3007
rect 3523 2990 3525 3002
rect 3523 2984 3527 2990
rect 3545 2944 3549 3007
rect 3591 2944 3595 3021
rect 3611 3033 3617 3049
rect 3611 3021 3614 3033
rect 3611 2944 3615 3021
rect 3662 3019 3666 3064
rect 3691 3053 3695 3076
rect 3686 3041 3695 3053
rect 3662 2996 3666 3007
rect 3662 2988 3680 2996
rect 3676 2984 3680 2988
rect 3684 2984 3688 3041
rect 3711 2999 3715 3076
rect 3783 3070 3787 3076
rect 3783 3058 3785 3070
rect 3805 3019 3809 3096
rect 3851 3071 3855 3076
rect 3842 3064 3855 3071
rect 3842 3019 3846 3064
rect 3871 3053 3875 3076
rect 3866 3041 3875 3053
rect 3805 3007 3814 3019
rect 3706 2987 3713 2999
rect 3783 2990 3785 3002
rect 3706 2944 3710 2987
rect 3783 2984 3787 2990
rect 3805 2944 3809 3007
rect 3842 2996 3846 3007
rect 3842 2988 3860 2996
rect 3856 2984 3860 2988
rect 3864 2984 3868 3041
rect 3891 2999 3895 3076
rect 3952 2999 3956 3056
rect 3886 2987 3893 2999
rect 3946 2987 3956 2999
rect 3886 2944 3890 2987
rect 3940 2956 3946 2987
rect 3960 2979 3964 3056
rect 3968 2999 3972 3056
rect 4051 3019 4055 3096
rect 4073 3070 4077 3076
rect 4075 3058 4077 3070
rect 4152 3053 4156 3096
rect 4046 3007 4055 3019
rect 3968 2987 3975 2999
rect 3987 2987 3995 2999
rect 3960 2960 3966 2967
rect 3960 2956 3975 2960
rect 3940 2952 3955 2956
rect 3951 2944 3955 2952
rect 3971 2944 3975 2956
rect 3991 2944 3995 2987
rect 4051 2944 4055 3007
rect 4145 3041 4154 3053
rect 4075 2990 4077 3002
rect 4073 2984 4077 2990
rect 4145 2984 4149 3041
rect 4174 3039 4178 3076
rect 4182 3072 4186 3076
rect 4182 3066 4201 3072
rect 4194 3053 4201 3066
rect 4174 3004 4180 3027
rect 4194 3004 4201 3041
rect 4165 2998 4180 3004
rect 4185 2998 4201 3004
rect 4232 2999 4236 3056
rect 4165 2984 4169 2998
rect 4185 2984 4189 2998
rect 4226 2987 4236 2999
rect 4220 2956 4226 2987
rect 4240 2979 4244 3056
rect 4248 2999 4252 3056
rect 4352 3053 4356 3096
rect 4345 3041 4354 3053
rect 4248 2987 4255 2999
rect 4267 2987 4275 2999
rect 4240 2960 4246 2967
rect 4240 2956 4255 2960
rect 4220 2952 4235 2956
rect 4231 2944 4235 2952
rect 4251 2944 4255 2956
rect 4271 2944 4275 2987
rect 4345 2984 4349 3041
rect 4374 3039 4378 3076
rect 4382 3072 4386 3076
rect 4382 3066 4401 3072
rect 4394 3053 4401 3066
rect 4374 3004 4380 3027
rect 4394 3004 4401 3041
rect 4365 2998 4380 3004
rect 4385 2998 4401 3004
rect 4468 2999 4472 3056
rect 4365 2984 4369 2998
rect 4385 2984 4389 2998
rect 4445 2987 4453 2999
rect 4465 2987 4472 2999
rect 4445 2944 4449 2987
rect 4476 2979 4480 3056
rect 4484 2999 4488 3056
rect 4545 3039 4549 3096
rect 4545 3027 4554 3039
rect 4484 2987 4494 2999
rect 4474 2960 4480 2967
rect 4465 2956 4480 2960
rect 4494 2956 4500 2987
rect 4465 2944 4469 2956
rect 4485 2952 4500 2956
rect 4485 2944 4489 2952
rect 4545 2944 4549 3027
rect 4605 2999 4609 3076
rect 4625 3053 4629 3076
rect 4645 3071 4649 3076
rect 4691 3071 4695 3076
rect 4645 3064 4658 3071
rect 4625 3041 4634 3053
rect 4607 2987 4614 2999
rect 4610 2944 4614 2987
rect 4632 2984 4636 3041
rect 4654 3019 4658 3064
rect 4682 3064 4695 3071
rect 4682 3019 4686 3064
rect 4711 3053 4715 3076
rect 4706 3041 4715 3053
rect 4654 2996 4658 3007
rect 4640 2988 4658 2996
rect 4682 2996 4686 3007
rect 4682 2988 4700 2996
rect 4640 2984 4644 2988
rect 4696 2984 4700 2988
rect 4704 2984 4708 3041
rect 4731 2999 4735 3076
rect 4726 2987 4733 2999
rect 4726 2944 4730 2987
rect 35 2900 39 2904
rect 55 2900 59 2904
rect 69 2900 73 2904
rect 89 2900 93 2904
rect 101 2900 105 2904
rect 121 2900 125 2904
rect 167 2900 171 2904
rect 175 2900 179 2904
rect 195 2900 199 2904
rect 203 2900 207 2904
rect 225 2900 229 2904
rect 290 2900 294 2904
rect 312 2900 316 2904
rect 320 2900 324 2904
rect 385 2900 389 2904
rect 405 2900 409 2904
rect 451 2900 455 2904
rect 473 2900 477 2904
rect 481 2900 485 2904
rect 501 2900 505 2904
rect 509 2900 513 2904
rect 555 2900 559 2904
rect 575 2900 579 2904
rect 587 2900 591 2904
rect 607 2900 611 2904
rect 621 2900 625 2904
rect 641 2900 645 2904
rect 695 2900 699 2904
rect 715 2900 719 2904
rect 729 2900 733 2904
rect 749 2900 753 2904
rect 761 2900 765 2904
rect 781 2900 785 2904
rect 827 2900 831 2904
rect 835 2900 839 2904
rect 855 2900 859 2904
rect 863 2900 867 2904
rect 885 2900 889 2904
rect 931 2900 935 2904
rect 1017 2900 1021 2904
rect 1025 2900 1029 2904
rect 1085 2900 1089 2904
rect 1105 2900 1109 2904
rect 1156 2900 1160 2904
rect 1164 2900 1168 2904
rect 1186 2900 1190 2904
rect 1251 2900 1255 2904
rect 1271 2900 1275 2904
rect 1291 2900 1295 2904
rect 1355 2900 1359 2904
rect 1375 2900 1379 2904
rect 1389 2900 1393 2904
rect 1409 2900 1413 2904
rect 1421 2900 1425 2904
rect 1441 2900 1445 2904
rect 1487 2900 1491 2904
rect 1495 2900 1499 2904
rect 1515 2900 1519 2904
rect 1523 2900 1527 2904
rect 1545 2900 1549 2904
rect 1617 2900 1621 2904
rect 1625 2900 1629 2904
rect 1685 2900 1689 2904
rect 1705 2900 1709 2904
rect 1756 2900 1760 2904
rect 1764 2900 1768 2904
rect 1786 2900 1790 2904
rect 1870 2900 1874 2904
rect 1892 2900 1896 2904
rect 1900 2900 1904 2904
rect 1951 2900 1955 2904
rect 1973 2900 1977 2904
rect 1981 2900 1985 2904
rect 2001 2900 2005 2904
rect 2009 2900 2013 2904
rect 2055 2900 2059 2904
rect 2075 2900 2079 2904
rect 2087 2900 2091 2904
rect 2107 2900 2111 2904
rect 2121 2900 2125 2904
rect 2141 2900 2145 2904
rect 2217 2900 2221 2904
rect 2225 2900 2229 2904
rect 2285 2900 2289 2904
rect 2345 2900 2349 2904
rect 2365 2900 2369 2904
rect 2385 2900 2389 2904
rect 2445 2900 2449 2904
rect 2465 2900 2469 2904
rect 2485 2900 2489 2904
rect 2545 2900 2549 2904
rect 2565 2900 2569 2904
rect 2585 2900 2589 2904
rect 2650 2900 2654 2904
rect 2672 2900 2676 2904
rect 2680 2900 2684 2904
rect 2757 2900 2761 2904
rect 2765 2900 2769 2904
rect 2811 2900 2815 2904
rect 2831 2900 2835 2904
rect 2891 2900 2895 2904
rect 2911 2900 2915 2904
rect 2971 2900 2975 2904
rect 2991 2900 2995 2904
rect 3011 2900 3015 2904
rect 3031 2900 3035 2904
rect 3091 2900 3095 2904
rect 3111 2900 3115 2904
rect 3176 2900 3180 2904
rect 3184 2900 3188 2904
rect 3206 2900 3210 2904
rect 3271 2900 3275 2904
rect 3331 2900 3335 2904
rect 3353 2900 3357 2904
rect 3375 2900 3379 2904
rect 3443 2900 3447 2904
rect 3465 2900 3469 2904
rect 3523 2900 3527 2904
rect 3545 2900 3549 2904
rect 3591 2900 3595 2904
rect 3611 2900 3615 2904
rect 3676 2900 3680 2904
rect 3684 2900 3688 2904
rect 3706 2900 3710 2904
rect 3783 2900 3787 2904
rect 3805 2900 3809 2904
rect 3856 2900 3860 2904
rect 3864 2900 3868 2904
rect 3886 2900 3890 2904
rect 3951 2900 3955 2904
rect 3971 2900 3975 2904
rect 3991 2900 3995 2904
rect 4051 2900 4055 2904
rect 4073 2900 4077 2904
rect 4145 2900 4149 2904
rect 4165 2900 4169 2904
rect 4185 2900 4189 2904
rect 4231 2900 4235 2904
rect 4251 2900 4255 2904
rect 4271 2900 4275 2904
rect 4345 2900 4349 2904
rect 4365 2900 4369 2904
rect 4385 2900 4389 2904
rect 4445 2900 4449 2904
rect 4465 2900 4469 2904
rect 4485 2900 4489 2904
rect 4545 2900 4549 2904
rect 4610 2900 4614 2904
rect 4632 2900 4636 2904
rect 4640 2900 4644 2904
rect 4696 2900 4700 2904
rect 4704 2900 4708 2904
rect 4726 2900 4730 2904
rect 35 2876 39 2880
rect 55 2876 59 2880
rect 69 2876 73 2880
rect 89 2876 93 2880
rect 101 2876 105 2880
rect 121 2876 125 2880
rect 167 2876 171 2880
rect 175 2876 179 2880
rect 195 2876 199 2880
rect 203 2876 207 2880
rect 225 2876 229 2880
rect 285 2876 289 2880
rect 305 2876 309 2880
rect 325 2876 329 2880
rect 345 2876 349 2880
rect 391 2876 395 2880
rect 411 2876 415 2880
rect 490 2876 494 2880
rect 512 2876 516 2880
rect 520 2876 524 2880
rect 583 2876 587 2880
rect 605 2876 609 2880
rect 651 2876 655 2880
rect 671 2876 675 2880
rect 750 2876 754 2880
rect 772 2876 776 2880
rect 780 2876 784 2880
rect 857 2876 861 2880
rect 865 2876 869 2880
rect 925 2876 929 2880
rect 945 2876 949 2880
rect 991 2876 995 2880
rect 1065 2876 1069 2880
rect 1085 2876 1089 2880
rect 1131 2876 1135 2880
rect 1139 2876 1143 2880
rect 1223 2876 1227 2880
rect 1245 2876 1249 2880
rect 1295 2876 1299 2880
rect 1315 2876 1319 2880
rect 1329 2876 1333 2880
rect 1349 2876 1353 2880
rect 1361 2876 1365 2880
rect 1381 2876 1385 2880
rect 1427 2876 1431 2880
rect 1435 2876 1439 2880
rect 1455 2876 1459 2880
rect 1463 2876 1467 2880
rect 1485 2876 1489 2880
rect 1531 2876 1535 2880
rect 1551 2876 1555 2880
rect 1630 2876 1634 2880
rect 1652 2876 1656 2880
rect 1660 2876 1664 2880
rect 1730 2876 1734 2880
rect 1752 2876 1756 2880
rect 1760 2876 1764 2880
rect 1837 2876 1841 2880
rect 1845 2876 1849 2880
rect 1905 2876 1909 2880
rect 1925 2876 1929 2880
rect 1945 2876 1949 2880
rect 2003 2876 2007 2880
rect 2025 2876 2029 2880
rect 2085 2876 2089 2880
rect 2105 2876 2109 2880
rect 2125 2876 2129 2880
rect 2171 2876 2175 2880
rect 2193 2876 2197 2880
rect 2255 2876 2259 2880
rect 2275 2876 2279 2880
rect 2289 2876 2293 2880
rect 2309 2876 2313 2880
rect 2321 2876 2325 2880
rect 2341 2876 2345 2880
rect 2387 2876 2391 2880
rect 2395 2876 2399 2880
rect 2415 2876 2419 2880
rect 2423 2876 2427 2880
rect 2445 2876 2449 2880
rect 2510 2876 2514 2880
rect 2532 2876 2536 2880
rect 2540 2876 2544 2880
rect 2610 2876 2614 2880
rect 2632 2876 2636 2880
rect 2640 2876 2644 2880
rect 2696 2876 2700 2880
rect 2704 2876 2708 2880
rect 2726 2876 2730 2880
rect 2791 2876 2795 2880
rect 2811 2876 2815 2880
rect 2871 2876 2875 2880
rect 2891 2876 2895 2880
rect 2956 2876 2960 2880
rect 2964 2876 2968 2880
rect 2986 2876 2990 2880
rect 3056 2876 3060 2880
rect 3064 2876 3068 2880
rect 3086 2876 3090 2880
rect 3151 2876 3155 2880
rect 3171 2876 3175 2880
rect 3250 2876 3254 2880
rect 3272 2876 3276 2880
rect 3280 2876 3284 2880
rect 3345 2876 3349 2880
rect 3365 2876 3369 2880
rect 3411 2876 3415 2880
rect 3431 2876 3435 2880
rect 3451 2876 3455 2880
rect 3530 2876 3534 2880
rect 3552 2876 3556 2880
rect 3560 2876 3564 2880
rect 3616 2876 3620 2880
rect 3624 2876 3628 2880
rect 3646 2876 3650 2880
rect 3725 2876 3729 2880
rect 3745 2876 3749 2880
rect 3810 2876 3814 2880
rect 3832 2876 3836 2880
rect 3840 2876 3844 2880
rect 3891 2876 3895 2880
rect 3911 2876 3915 2880
rect 3931 2876 3935 2880
rect 3991 2876 3995 2880
rect 4065 2876 4069 2880
rect 4085 2876 4089 2880
rect 4105 2876 4109 2880
rect 4125 2876 4129 2880
rect 4171 2876 4175 2880
rect 4191 2876 4195 2880
rect 4211 2876 4215 2880
rect 4276 2876 4280 2880
rect 4284 2876 4288 2880
rect 4306 2876 4310 2880
rect 4371 2876 4375 2880
rect 4393 2876 4397 2880
rect 4415 2876 4419 2880
rect 4471 2876 4475 2880
rect 4491 2876 4495 2880
rect 4511 2876 4515 2880
rect 4531 2876 4535 2880
rect 4591 2876 4595 2880
rect 4651 2876 4655 2880
rect 4671 2876 4675 2880
rect 4691 2876 4695 2880
rect 35 2753 39 2796
rect 55 2754 59 2836
rect 69 2777 73 2836
rect 89 2796 93 2836
rect 101 2830 105 2836
rect 95 2784 98 2796
rect 69 2769 78 2777
rect 35 2704 39 2741
rect 55 2684 59 2742
rect 74 2740 78 2769
rect 94 2720 98 2784
rect 65 2716 98 2720
rect 65 2684 69 2716
rect 103 2708 107 2818
rect 121 2810 125 2836
rect 167 2832 171 2836
rect 135 2830 171 2832
rect 147 2828 171 2830
rect 89 2696 91 2708
rect 87 2684 91 2696
rect 97 2696 99 2708
rect 97 2684 101 2696
rect 119 2684 123 2798
rect 135 2692 139 2818
rect 175 2804 179 2836
rect 195 2816 199 2856
rect 203 2833 207 2856
rect 203 2826 211 2833
rect 173 2709 179 2804
rect 207 2797 211 2826
rect 203 2791 211 2797
rect 203 2745 207 2791
rect 225 2784 229 2796
rect 227 2772 229 2784
rect 285 2773 289 2796
rect 173 2705 197 2709
rect 159 2700 177 2701
rect 147 2696 177 2700
rect 135 2688 169 2692
rect 165 2684 169 2688
rect 173 2684 177 2696
rect 193 2684 197 2705
rect 203 2684 207 2733
rect 225 2704 229 2772
rect 286 2761 289 2773
rect 280 2713 286 2761
rect 305 2739 309 2796
rect 325 2774 329 2796
rect 345 2774 349 2796
rect 325 2768 338 2774
rect 345 2773 365 2774
rect 345 2768 353 2773
rect 334 2739 338 2768
rect 307 2727 309 2739
rect 305 2725 309 2727
rect 305 2718 318 2725
rect 280 2709 310 2713
rect 306 2704 310 2709
rect 314 2704 318 2718
rect 334 2704 338 2727
rect 353 2719 359 2761
rect 391 2759 395 2836
rect 386 2747 395 2759
rect 389 2731 395 2747
rect 411 2759 415 2836
rect 490 2793 494 2836
rect 487 2781 494 2793
rect 411 2747 414 2759
rect 411 2731 417 2747
rect 389 2724 397 2731
rect 342 2712 359 2719
rect 342 2704 346 2712
rect 393 2704 397 2724
rect 403 2724 417 2731
rect 403 2704 407 2724
rect 485 2704 489 2781
rect 512 2739 516 2796
rect 520 2792 524 2796
rect 520 2784 538 2792
rect 534 2773 538 2784
rect 583 2790 587 2796
rect 583 2778 585 2790
rect 605 2773 609 2836
rect 605 2761 614 2773
rect 505 2727 514 2739
rect 505 2704 509 2727
rect 534 2716 538 2761
rect 525 2709 538 2716
rect 583 2710 585 2722
rect 525 2704 529 2709
rect 583 2704 587 2710
rect 605 2684 609 2761
rect 651 2759 655 2836
rect 646 2747 655 2759
rect 649 2731 655 2747
rect 671 2759 675 2836
rect 750 2793 754 2836
rect 747 2781 754 2793
rect 671 2747 674 2759
rect 671 2731 677 2747
rect 649 2724 657 2731
rect 653 2704 657 2724
rect 663 2724 677 2731
rect 663 2704 667 2724
rect 745 2704 749 2781
rect 772 2739 776 2796
rect 780 2792 784 2796
rect 780 2784 798 2792
rect 794 2773 798 2784
rect 857 2773 861 2796
rect 846 2761 861 2773
rect 865 2773 869 2796
rect 865 2761 874 2773
rect 765 2727 774 2739
rect 765 2704 769 2727
rect 794 2716 798 2761
rect 785 2709 798 2716
rect 785 2704 789 2709
rect 845 2684 849 2761
rect 865 2684 869 2761
rect 925 2759 929 2836
rect 926 2747 929 2759
rect 923 2731 929 2747
rect 945 2759 949 2836
rect 945 2747 954 2759
rect 991 2753 995 2836
rect 1065 2759 1069 2836
rect 945 2731 951 2747
rect 986 2741 995 2753
rect 1066 2747 1069 2759
rect 923 2724 937 2731
rect 933 2704 937 2724
rect 943 2724 951 2731
rect 943 2704 947 2724
rect 991 2684 995 2741
rect 1063 2731 1069 2747
rect 1085 2759 1089 2836
rect 1131 2773 1135 2796
rect 1126 2761 1135 2773
rect 1139 2773 1143 2796
rect 1223 2790 1227 2796
rect 1223 2778 1225 2790
rect 1245 2773 1249 2836
rect 1139 2761 1154 2773
rect 1245 2761 1254 2773
rect 1085 2747 1094 2759
rect 1085 2731 1091 2747
rect 1063 2724 1077 2731
rect 1073 2704 1077 2724
rect 1083 2724 1091 2731
rect 1083 2704 1087 2724
rect 1131 2684 1135 2761
rect 1151 2684 1155 2761
rect 1223 2710 1225 2722
rect 1223 2704 1227 2710
rect 1245 2684 1249 2761
rect 1295 2753 1299 2796
rect 1315 2754 1319 2836
rect 1329 2777 1333 2836
rect 1349 2796 1353 2836
rect 1361 2830 1365 2836
rect 1355 2784 1358 2796
rect 1329 2769 1338 2777
rect 1295 2704 1299 2741
rect 1315 2684 1319 2742
rect 1334 2740 1338 2769
rect 1354 2720 1358 2784
rect 1325 2716 1358 2720
rect 1325 2684 1329 2716
rect 1363 2708 1367 2818
rect 1381 2810 1385 2836
rect 1427 2832 1431 2836
rect 1395 2830 1431 2832
rect 1407 2828 1431 2830
rect 1349 2696 1351 2708
rect 1347 2684 1351 2696
rect 1357 2696 1359 2708
rect 1357 2684 1361 2696
rect 1379 2684 1383 2798
rect 1395 2692 1399 2818
rect 1435 2804 1439 2836
rect 1455 2816 1459 2856
rect 1463 2833 1467 2856
rect 1463 2826 1471 2833
rect 1433 2709 1439 2804
rect 1467 2797 1471 2826
rect 1463 2791 1471 2797
rect 1463 2745 1467 2791
rect 1485 2784 1489 2796
rect 1487 2772 1489 2784
rect 1433 2705 1457 2709
rect 1419 2700 1437 2701
rect 1407 2696 1437 2700
rect 1395 2688 1429 2692
rect 1425 2684 1429 2688
rect 1433 2684 1437 2696
rect 1453 2684 1457 2705
rect 1463 2684 1467 2733
rect 1485 2704 1489 2772
rect 1531 2759 1535 2836
rect 1526 2747 1535 2759
rect 1529 2731 1535 2747
rect 1551 2759 1555 2836
rect 1630 2793 1634 2836
rect 1627 2781 1634 2793
rect 1551 2747 1554 2759
rect 1551 2731 1557 2747
rect 1529 2724 1537 2731
rect 1533 2704 1537 2724
rect 1543 2724 1557 2731
rect 1543 2704 1547 2724
rect 1625 2704 1629 2781
rect 1652 2739 1656 2796
rect 1660 2792 1664 2796
rect 1730 2793 1734 2836
rect 1660 2784 1678 2792
rect 1674 2773 1678 2784
rect 1727 2781 1734 2793
rect 1645 2727 1654 2739
rect 1645 2704 1649 2727
rect 1674 2716 1678 2761
rect 1665 2709 1678 2716
rect 1665 2704 1669 2709
rect 1725 2704 1729 2781
rect 1752 2739 1756 2796
rect 1760 2792 1764 2796
rect 1760 2784 1778 2792
rect 1774 2773 1778 2784
rect 1837 2773 1841 2796
rect 1826 2761 1841 2773
rect 1845 2773 1849 2796
rect 1845 2761 1854 2773
rect 1745 2727 1754 2739
rect 1745 2704 1749 2727
rect 1774 2716 1778 2761
rect 1765 2709 1778 2716
rect 1765 2704 1769 2709
rect 1825 2684 1829 2761
rect 1845 2684 1849 2761
rect 1905 2739 1909 2796
rect 1925 2782 1929 2796
rect 1945 2782 1949 2796
rect 2003 2790 2007 2796
rect 1925 2776 1940 2782
rect 1945 2776 1961 2782
rect 2003 2778 2005 2790
rect 1934 2753 1940 2776
rect 1905 2727 1914 2739
rect 1912 2684 1916 2727
rect 1934 2704 1938 2741
rect 1954 2739 1961 2776
rect 2025 2773 2029 2836
rect 2085 2793 2089 2836
rect 2105 2824 2109 2836
rect 2125 2828 2129 2836
rect 2125 2824 2140 2828
rect 2105 2820 2120 2824
rect 2114 2813 2120 2820
rect 2085 2781 2093 2793
rect 2105 2781 2112 2793
rect 2025 2761 2034 2773
rect 1954 2714 1961 2727
rect 1942 2708 1961 2714
rect 2003 2710 2005 2722
rect 1942 2704 1946 2708
rect 2003 2704 2007 2710
rect 2025 2684 2029 2761
rect 2108 2724 2112 2781
rect 2116 2724 2120 2801
rect 2134 2793 2140 2824
rect 2124 2781 2134 2793
rect 2124 2724 2128 2781
rect 2171 2773 2175 2836
rect 2193 2790 2197 2796
rect 2195 2778 2197 2790
rect 2166 2761 2175 2773
rect 2171 2684 2175 2761
rect 2255 2753 2259 2796
rect 2275 2754 2279 2836
rect 2289 2777 2293 2836
rect 2309 2796 2313 2836
rect 2321 2830 2325 2836
rect 2315 2784 2318 2796
rect 2289 2769 2298 2777
rect 2195 2710 2197 2722
rect 2193 2704 2197 2710
rect 2255 2704 2259 2741
rect 2275 2684 2279 2742
rect 2294 2740 2298 2769
rect 2314 2720 2318 2784
rect 2285 2716 2318 2720
rect 2285 2684 2289 2716
rect 2323 2708 2327 2818
rect 2341 2810 2345 2836
rect 2387 2832 2391 2836
rect 2355 2830 2391 2832
rect 2367 2828 2391 2830
rect 2309 2696 2311 2708
rect 2307 2684 2311 2696
rect 2317 2696 2319 2708
rect 2317 2684 2321 2696
rect 2339 2684 2343 2798
rect 2355 2692 2359 2818
rect 2395 2804 2399 2836
rect 2415 2816 2419 2856
rect 2423 2833 2427 2856
rect 2423 2826 2431 2833
rect 2393 2709 2399 2804
rect 2427 2797 2431 2826
rect 2423 2791 2431 2797
rect 2423 2745 2427 2791
rect 2445 2784 2449 2796
rect 2510 2793 2514 2836
rect 2447 2772 2449 2784
rect 2507 2781 2514 2793
rect 2393 2705 2417 2709
rect 2379 2700 2397 2701
rect 2367 2696 2397 2700
rect 2355 2688 2389 2692
rect 2385 2684 2389 2688
rect 2393 2684 2397 2696
rect 2413 2684 2417 2705
rect 2423 2684 2427 2733
rect 2445 2704 2449 2772
rect 2505 2704 2509 2781
rect 2532 2739 2536 2796
rect 2540 2792 2544 2796
rect 2610 2793 2614 2836
rect 2540 2784 2558 2792
rect 2554 2773 2558 2784
rect 2607 2781 2614 2793
rect 2525 2727 2534 2739
rect 2525 2704 2529 2727
rect 2554 2716 2558 2761
rect 2545 2709 2558 2716
rect 2545 2704 2549 2709
rect 2605 2704 2609 2781
rect 2632 2739 2636 2796
rect 2640 2792 2644 2796
rect 2696 2792 2700 2796
rect 2640 2784 2658 2792
rect 2654 2773 2658 2784
rect 2682 2784 2700 2792
rect 2682 2773 2686 2784
rect 2625 2727 2634 2739
rect 2625 2704 2629 2727
rect 2654 2716 2658 2761
rect 2645 2709 2658 2716
rect 2682 2716 2686 2761
rect 2704 2739 2708 2796
rect 2726 2793 2730 2836
rect 2726 2781 2733 2793
rect 2706 2727 2715 2739
rect 2682 2709 2695 2716
rect 2645 2704 2649 2709
rect 2691 2704 2695 2709
rect 2711 2704 2715 2727
rect 2731 2704 2735 2781
rect 2791 2759 2795 2836
rect 2786 2747 2795 2759
rect 2789 2731 2795 2747
rect 2811 2759 2815 2836
rect 2871 2759 2875 2836
rect 2811 2747 2814 2759
rect 2866 2747 2875 2759
rect 2811 2731 2817 2747
rect 2789 2724 2797 2731
rect 2793 2704 2797 2724
rect 2803 2724 2817 2731
rect 2869 2731 2875 2747
rect 2891 2759 2895 2836
rect 2956 2792 2960 2796
rect 2942 2784 2960 2792
rect 2942 2773 2946 2784
rect 2891 2747 2894 2759
rect 2891 2731 2897 2747
rect 2869 2724 2877 2731
rect 2803 2704 2807 2724
rect 2873 2704 2877 2724
rect 2883 2724 2897 2731
rect 2883 2704 2887 2724
rect 2942 2716 2946 2761
rect 2964 2739 2968 2796
rect 2986 2793 2990 2836
rect 2986 2781 2993 2793
rect 3056 2792 3060 2796
rect 3042 2784 3060 2792
rect 2966 2727 2975 2739
rect 2942 2709 2955 2716
rect 2951 2704 2955 2709
rect 2971 2704 2975 2727
rect 2991 2704 2995 2781
rect 3042 2773 3046 2784
rect 3042 2716 3046 2761
rect 3064 2739 3068 2796
rect 3086 2793 3090 2836
rect 3086 2781 3093 2793
rect 3066 2727 3075 2739
rect 3042 2709 3055 2716
rect 3051 2704 3055 2709
rect 3071 2704 3075 2727
rect 3091 2704 3095 2781
rect 3151 2759 3155 2836
rect 3146 2747 3155 2759
rect 3149 2731 3155 2747
rect 3171 2759 3175 2836
rect 3250 2793 3254 2836
rect 3247 2781 3254 2793
rect 3171 2747 3174 2759
rect 3171 2731 3177 2747
rect 3149 2724 3157 2731
rect 3153 2704 3157 2724
rect 3163 2724 3177 2731
rect 3163 2704 3167 2724
rect 3245 2704 3249 2781
rect 3272 2739 3276 2796
rect 3280 2792 3284 2796
rect 3280 2784 3298 2792
rect 3294 2773 3298 2784
rect 3265 2727 3274 2739
rect 3265 2704 3269 2727
rect 3294 2716 3298 2761
rect 3345 2759 3349 2836
rect 3346 2747 3349 2759
rect 3343 2731 3349 2747
rect 3365 2759 3369 2836
rect 3411 2828 3415 2836
rect 3400 2824 3415 2828
rect 3431 2824 3435 2836
rect 3400 2793 3406 2824
rect 3420 2820 3435 2824
rect 3420 2813 3426 2820
rect 3406 2781 3416 2793
rect 3365 2747 3374 2759
rect 3365 2731 3371 2747
rect 3343 2724 3357 2731
rect 3285 2709 3298 2716
rect 3285 2704 3289 2709
rect 3353 2704 3357 2724
rect 3363 2724 3371 2731
rect 3412 2724 3416 2781
rect 3420 2724 3424 2801
rect 3451 2793 3455 2836
rect 3530 2793 3534 2836
rect 3428 2781 3435 2793
rect 3447 2781 3455 2793
rect 3527 2781 3534 2793
rect 3428 2724 3432 2781
rect 3363 2704 3367 2724
rect 3525 2704 3529 2781
rect 3552 2739 3556 2796
rect 3560 2792 3564 2796
rect 3616 2792 3620 2796
rect 3560 2784 3578 2792
rect 3574 2773 3578 2784
rect 3602 2784 3620 2792
rect 3602 2773 3606 2784
rect 3545 2727 3554 2739
rect 3545 2704 3549 2727
rect 3574 2716 3578 2761
rect 3565 2709 3578 2716
rect 3602 2716 3606 2761
rect 3624 2739 3628 2796
rect 3646 2793 3650 2836
rect 3646 2781 3653 2793
rect 3626 2727 3635 2739
rect 3602 2709 3615 2716
rect 3565 2704 3569 2709
rect 3611 2704 3615 2709
rect 3631 2704 3635 2727
rect 3651 2704 3655 2781
rect 3725 2759 3729 2836
rect 3726 2747 3729 2759
rect 3723 2731 3729 2747
rect 3745 2759 3749 2836
rect 3810 2793 3814 2836
rect 3891 2828 3895 2836
rect 3880 2824 3895 2828
rect 3911 2824 3915 2836
rect 3807 2781 3814 2793
rect 3745 2747 3754 2759
rect 3745 2731 3751 2747
rect 3723 2724 3737 2731
rect 3733 2704 3737 2724
rect 3743 2724 3751 2731
rect 3743 2704 3747 2724
rect 3805 2704 3809 2781
rect 3832 2739 3836 2796
rect 3840 2792 3844 2796
rect 3880 2793 3886 2824
rect 3900 2820 3915 2824
rect 3900 2813 3906 2820
rect 3840 2784 3858 2792
rect 3854 2773 3858 2784
rect 3886 2781 3896 2793
rect 3825 2727 3834 2739
rect 3825 2704 3829 2727
rect 3854 2716 3858 2761
rect 3892 2724 3896 2781
rect 3900 2724 3904 2801
rect 3931 2793 3935 2836
rect 3908 2781 3915 2793
rect 3927 2781 3935 2793
rect 3908 2724 3912 2781
rect 3991 2753 3995 2836
rect 4171 2828 4175 2836
rect 4160 2824 4175 2828
rect 4191 2824 4195 2836
rect 4065 2773 4069 2796
rect 4066 2761 4069 2773
rect 3986 2741 3995 2753
rect 3845 2709 3858 2716
rect 3845 2704 3849 2709
rect 3991 2684 3995 2741
rect 4060 2713 4066 2761
rect 4085 2739 4089 2796
rect 4105 2774 4109 2796
rect 4125 2774 4129 2796
rect 4160 2793 4166 2824
rect 4180 2820 4195 2824
rect 4180 2813 4186 2820
rect 4166 2781 4176 2793
rect 4105 2768 4118 2774
rect 4125 2773 4145 2774
rect 4125 2768 4133 2773
rect 4114 2739 4118 2768
rect 4087 2727 4089 2739
rect 4085 2725 4089 2727
rect 4085 2718 4098 2725
rect 4060 2709 4090 2713
rect 4086 2704 4090 2709
rect 4094 2704 4098 2718
rect 4114 2704 4118 2727
rect 4133 2719 4139 2761
rect 4172 2724 4176 2781
rect 4180 2724 4184 2801
rect 4211 2793 4215 2836
rect 4188 2781 4195 2793
rect 4207 2781 4215 2793
rect 4276 2792 4280 2796
rect 4262 2784 4280 2792
rect 4188 2724 4192 2781
rect 4262 2773 4266 2784
rect 4122 2712 4139 2719
rect 4122 2704 4126 2712
rect 4262 2716 4266 2761
rect 4284 2739 4288 2796
rect 4306 2793 4310 2836
rect 4306 2781 4313 2793
rect 4286 2727 4295 2739
rect 4262 2709 4275 2716
rect 4271 2704 4275 2709
rect 4291 2704 4295 2727
rect 4311 2704 4315 2781
rect 4371 2773 4375 2836
rect 4366 2761 4375 2773
rect 4371 2704 4375 2761
rect 4393 2759 4397 2836
rect 4381 2747 4394 2759
rect 4381 2704 4385 2747
rect 4415 2722 4419 2796
rect 4471 2774 4475 2796
rect 4491 2774 4495 2796
rect 4455 2773 4475 2774
rect 4467 2768 4475 2773
rect 4482 2768 4495 2774
rect 4407 2710 4419 2722
rect 4461 2719 4467 2761
rect 4482 2739 4486 2768
rect 4511 2739 4515 2796
rect 4531 2773 4535 2796
rect 4531 2761 4534 2773
rect 4511 2727 4513 2739
rect 4461 2712 4478 2719
rect 4401 2704 4405 2710
rect 4474 2704 4478 2712
rect 4482 2704 4486 2727
rect 4511 2725 4515 2727
rect 4502 2718 4515 2725
rect 4502 2704 4506 2718
rect 4534 2713 4540 2761
rect 4591 2753 4595 2836
rect 4651 2782 4655 2796
rect 4671 2782 4675 2796
rect 4586 2741 4595 2753
rect 4510 2709 4540 2713
rect 4510 2704 4514 2709
rect 4591 2684 4595 2741
rect 4639 2776 4655 2782
rect 4660 2776 4675 2782
rect 4639 2739 4646 2776
rect 4660 2753 4666 2776
rect 4639 2714 4646 2727
rect 4639 2708 4658 2714
rect 4654 2704 4658 2708
rect 4662 2704 4666 2741
rect 4691 2739 4695 2796
rect 4686 2727 4695 2739
rect 4684 2684 4688 2727
rect 35 2660 39 2664
rect 55 2660 59 2664
rect 65 2660 69 2664
rect 87 2660 91 2664
rect 97 2660 101 2664
rect 119 2660 123 2664
rect 165 2660 169 2664
rect 173 2660 177 2664
rect 193 2660 197 2664
rect 203 2660 207 2664
rect 225 2660 229 2664
rect 306 2660 310 2664
rect 314 2660 318 2664
rect 334 2660 338 2664
rect 342 2660 346 2664
rect 393 2660 397 2664
rect 403 2660 407 2664
rect 485 2660 489 2664
rect 505 2660 509 2664
rect 525 2660 529 2664
rect 583 2660 587 2664
rect 605 2660 609 2664
rect 653 2660 657 2664
rect 663 2660 667 2664
rect 745 2660 749 2664
rect 765 2660 769 2664
rect 785 2660 789 2664
rect 845 2660 849 2664
rect 865 2660 869 2664
rect 933 2660 937 2664
rect 943 2660 947 2664
rect 991 2660 995 2664
rect 1073 2660 1077 2664
rect 1083 2660 1087 2664
rect 1131 2660 1135 2664
rect 1151 2660 1155 2664
rect 1223 2660 1227 2664
rect 1245 2660 1249 2664
rect 1295 2660 1299 2664
rect 1315 2660 1319 2664
rect 1325 2660 1329 2664
rect 1347 2660 1351 2664
rect 1357 2660 1361 2664
rect 1379 2660 1383 2664
rect 1425 2660 1429 2664
rect 1433 2660 1437 2664
rect 1453 2660 1457 2664
rect 1463 2660 1467 2664
rect 1485 2660 1489 2664
rect 1533 2660 1537 2664
rect 1543 2660 1547 2664
rect 1625 2660 1629 2664
rect 1645 2660 1649 2664
rect 1665 2660 1669 2664
rect 1725 2660 1729 2664
rect 1745 2660 1749 2664
rect 1765 2660 1769 2664
rect 1825 2660 1829 2664
rect 1845 2660 1849 2664
rect 1912 2660 1916 2664
rect 1934 2660 1938 2664
rect 1942 2660 1946 2664
rect 2003 2660 2007 2664
rect 2025 2660 2029 2664
rect 2108 2660 2112 2664
rect 2116 2660 2120 2664
rect 2124 2660 2128 2664
rect 2171 2660 2175 2664
rect 2193 2660 2197 2664
rect 2255 2660 2259 2664
rect 2275 2660 2279 2664
rect 2285 2660 2289 2664
rect 2307 2660 2311 2664
rect 2317 2660 2321 2664
rect 2339 2660 2343 2664
rect 2385 2660 2389 2664
rect 2393 2660 2397 2664
rect 2413 2660 2417 2664
rect 2423 2660 2427 2664
rect 2445 2660 2449 2664
rect 2505 2660 2509 2664
rect 2525 2660 2529 2664
rect 2545 2660 2549 2664
rect 2605 2660 2609 2664
rect 2625 2660 2629 2664
rect 2645 2660 2649 2664
rect 2691 2660 2695 2664
rect 2711 2660 2715 2664
rect 2731 2660 2735 2664
rect 2793 2660 2797 2664
rect 2803 2660 2807 2664
rect 2873 2660 2877 2664
rect 2883 2660 2887 2664
rect 2951 2660 2955 2664
rect 2971 2660 2975 2664
rect 2991 2660 2995 2664
rect 3051 2660 3055 2664
rect 3071 2660 3075 2664
rect 3091 2660 3095 2664
rect 3153 2660 3157 2664
rect 3163 2660 3167 2664
rect 3245 2660 3249 2664
rect 3265 2660 3269 2664
rect 3285 2660 3289 2664
rect 3353 2660 3357 2664
rect 3363 2660 3367 2664
rect 3412 2660 3416 2664
rect 3420 2660 3424 2664
rect 3428 2660 3432 2664
rect 3525 2660 3529 2664
rect 3545 2660 3549 2664
rect 3565 2660 3569 2664
rect 3611 2660 3615 2664
rect 3631 2660 3635 2664
rect 3651 2660 3655 2664
rect 3733 2660 3737 2664
rect 3743 2660 3747 2664
rect 3805 2660 3809 2664
rect 3825 2660 3829 2664
rect 3845 2660 3849 2664
rect 3892 2660 3896 2664
rect 3900 2660 3904 2664
rect 3908 2660 3912 2664
rect 3991 2660 3995 2664
rect 4086 2660 4090 2664
rect 4094 2660 4098 2664
rect 4114 2660 4118 2664
rect 4122 2660 4126 2664
rect 4172 2660 4176 2664
rect 4180 2660 4184 2664
rect 4188 2660 4192 2664
rect 4271 2660 4275 2664
rect 4291 2660 4295 2664
rect 4311 2660 4315 2664
rect 4371 2660 4375 2664
rect 4381 2660 4385 2664
rect 4401 2660 4405 2664
rect 4474 2660 4478 2664
rect 4482 2660 4486 2664
rect 4502 2660 4506 2664
rect 4510 2660 4514 2664
rect 4591 2660 4595 2664
rect 4654 2660 4658 2664
rect 4662 2660 4666 2664
rect 4684 2660 4688 2664
rect 35 2636 39 2640
rect 55 2636 59 2640
rect 65 2636 69 2640
rect 87 2636 91 2640
rect 97 2636 101 2640
rect 119 2636 123 2640
rect 165 2636 169 2640
rect 173 2636 177 2640
rect 193 2636 197 2640
rect 203 2636 207 2640
rect 225 2636 229 2640
rect 285 2636 289 2640
rect 305 2636 309 2640
rect 325 2636 329 2640
rect 371 2636 375 2640
rect 393 2636 397 2640
rect 453 2636 457 2640
rect 463 2636 467 2640
rect 545 2636 549 2640
rect 565 2636 569 2640
rect 585 2636 589 2640
rect 631 2636 635 2640
rect 653 2636 657 2640
rect 725 2636 729 2640
rect 745 2636 749 2640
rect 765 2636 769 2640
rect 811 2636 815 2640
rect 831 2636 835 2640
rect 895 2636 899 2640
rect 915 2636 919 2640
rect 925 2636 929 2640
rect 947 2636 951 2640
rect 957 2636 961 2640
rect 979 2636 983 2640
rect 1025 2636 1029 2640
rect 1033 2636 1037 2640
rect 1053 2636 1057 2640
rect 1063 2636 1067 2640
rect 1085 2636 1089 2640
rect 1131 2636 1135 2640
rect 1191 2636 1195 2640
rect 1211 2636 1215 2640
rect 1231 2636 1235 2640
rect 1291 2636 1295 2640
rect 1353 2636 1357 2640
rect 1363 2636 1367 2640
rect 1431 2636 1435 2640
rect 1453 2636 1457 2640
rect 1463 2636 1467 2640
rect 1483 2636 1487 2640
rect 1491 2636 1495 2640
rect 1537 2636 1541 2640
rect 1559 2636 1563 2640
rect 1569 2636 1573 2640
rect 1591 2636 1595 2640
rect 1601 2636 1605 2640
rect 1621 2636 1625 2640
rect 1671 2636 1675 2640
rect 1691 2636 1695 2640
rect 1711 2636 1715 2640
rect 1771 2636 1775 2640
rect 1793 2636 1797 2640
rect 1803 2636 1807 2640
rect 1823 2636 1827 2640
rect 1831 2636 1835 2640
rect 1877 2636 1881 2640
rect 1899 2636 1903 2640
rect 1909 2636 1913 2640
rect 1931 2636 1935 2640
rect 1941 2636 1945 2640
rect 1961 2636 1965 2640
rect 2011 2636 2015 2640
rect 2031 2636 2035 2640
rect 2051 2636 2055 2640
rect 2071 2636 2075 2640
rect 2091 2636 2095 2640
rect 2111 2636 2115 2640
rect 2131 2636 2135 2640
rect 2151 2636 2155 2640
rect 2215 2636 2219 2640
rect 2235 2636 2239 2640
rect 2245 2636 2249 2640
rect 2267 2636 2271 2640
rect 2277 2636 2281 2640
rect 2299 2636 2303 2640
rect 2345 2636 2349 2640
rect 2353 2636 2357 2640
rect 2373 2636 2377 2640
rect 2383 2636 2387 2640
rect 2405 2636 2409 2640
rect 2473 2636 2477 2640
rect 2483 2636 2487 2640
rect 2531 2636 2535 2640
rect 2605 2636 2609 2640
rect 2625 2636 2629 2640
rect 2645 2636 2649 2640
rect 2691 2636 2695 2640
rect 2773 2636 2777 2640
rect 2783 2636 2787 2640
rect 2845 2636 2849 2640
rect 2865 2636 2869 2640
rect 2885 2636 2889 2640
rect 2931 2636 2935 2640
rect 2941 2636 2945 2640
rect 2961 2636 2965 2640
rect 3031 2636 3035 2640
rect 3051 2636 3055 2640
rect 3071 2636 3075 2640
rect 3153 2636 3157 2640
rect 3163 2636 3167 2640
rect 3211 2636 3215 2640
rect 3221 2636 3225 2640
rect 3241 2636 3245 2640
rect 3348 2636 3352 2640
rect 3356 2636 3360 2640
rect 3364 2636 3368 2640
rect 3411 2636 3415 2640
rect 3473 2636 3477 2640
rect 3483 2636 3487 2640
rect 3551 2636 3555 2640
rect 3561 2636 3565 2640
rect 3581 2636 3585 2640
rect 3651 2636 3655 2640
rect 3673 2636 3677 2640
rect 3731 2636 3735 2640
rect 3815 2636 3819 2640
rect 3835 2636 3839 2640
rect 3845 2636 3849 2640
rect 3926 2636 3930 2640
rect 3934 2636 3938 2640
rect 3954 2636 3958 2640
rect 3962 2636 3966 2640
rect 4033 2636 4037 2640
rect 4043 2636 4047 2640
rect 4113 2636 4117 2640
rect 4123 2636 4127 2640
rect 4171 2636 4175 2640
rect 4191 2636 4195 2640
rect 4211 2636 4215 2640
rect 4273 2636 4277 2640
rect 4283 2636 4287 2640
rect 4388 2636 4392 2640
rect 4396 2636 4400 2640
rect 4404 2636 4408 2640
rect 4488 2636 4492 2640
rect 4496 2636 4500 2640
rect 4504 2636 4508 2640
rect 4554 2636 4558 2640
rect 4562 2636 4566 2640
rect 4584 2636 4588 2640
rect 4688 2636 4692 2640
rect 4696 2636 4700 2640
rect 4704 2636 4708 2640
rect 35 2559 39 2596
rect 55 2558 59 2616
rect 65 2584 69 2616
rect 87 2604 91 2616
rect 89 2592 91 2604
rect 97 2604 101 2616
rect 97 2592 99 2604
rect 65 2580 98 2584
rect 35 2504 39 2547
rect 55 2464 59 2546
rect 74 2531 78 2560
rect 69 2523 78 2531
rect 69 2464 73 2523
rect 94 2516 98 2580
rect 95 2504 98 2516
rect 89 2464 93 2504
rect 103 2482 107 2592
rect 119 2502 123 2616
rect 165 2612 169 2616
rect 135 2608 169 2612
rect 101 2464 105 2470
rect 121 2464 125 2490
rect 135 2482 139 2608
rect 173 2604 177 2616
rect 147 2600 177 2604
rect 159 2599 177 2600
rect 193 2595 197 2616
rect 173 2591 197 2595
rect 173 2496 179 2591
rect 203 2567 207 2616
rect 203 2509 207 2555
rect 225 2528 229 2596
rect 227 2516 229 2528
rect 285 2519 289 2596
rect 305 2573 309 2596
rect 325 2591 329 2596
rect 325 2584 338 2591
rect 305 2561 314 2573
rect 203 2503 211 2509
rect 225 2504 229 2516
rect 287 2507 294 2519
rect 147 2470 171 2472
rect 135 2468 171 2470
rect 167 2464 171 2468
rect 175 2464 179 2496
rect 195 2444 199 2484
rect 207 2474 211 2503
rect 203 2467 211 2474
rect 203 2444 207 2467
rect 290 2464 294 2507
rect 312 2504 316 2561
rect 334 2539 338 2584
rect 371 2539 375 2616
rect 393 2590 397 2596
rect 395 2578 397 2590
rect 453 2576 457 2596
rect 449 2569 457 2576
rect 463 2576 467 2596
rect 463 2569 477 2576
rect 449 2553 455 2569
rect 446 2541 455 2553
rect 366 2527 375 2539
rect 334 2516 338 2527
rect 320 2508 338 2516
rect 320 2504 324 2508
rect 371 2464 375 2527
rect 395 2510 397 2522
rect 393 2504 397 2510
rect 451 2464 455 2541
rect 471 2553 477 2569
rect 471 2541 474 2553
rect 471 2464 475 2541
rect 545 2519 549 2596
rect 565 2573 569 2596
rect 585 2591 589 2596
rect 585 2584 598 2591
rect 565 2561 574 2573
rect 547 2507 554 2519
rect 550 2464 554 2507
rect 572 2504 576 2561
rect 594 2539 598 2584
rect 631 2539 635 2616
rect 653 2590 657 2596
rect 655 2578 657 2590
rect 626 2527 635 2539
rect 594 2516 598 2527
rect 580 2508 598 2516
rect 580 2504 584 2508
rect 631 2464 635 2527
rect 655 2510 657 2522
rect 725 2519 729 2596
rect 745 2573 749 2596
rect 765 2591 769 2596
rect 765 2584 778 2591
rect 745 2561 754 2573
rect 653 2504 657 2510
rect 727 2507 734 2519
rect 730 2464 734 2507
rect 752 2504 756 2561
rect 774 2539 778 2584
rect 811 2539 815 2616
rect 831 2539 835 2616
rect 895 2559 899 2596
rect 915 2558 919 2616
rect 925 2584 929 2616
rect 947 2604 951 2616
rect 949 2592 951 2604
rect 957 2604 961 2616
rect 957 2592 959 2604
rect 925 2580 958 2584
rect 806 2527 815 2539
rect 774 2516 778 2527
rect 760 2508 778 2516
rect 760 2504 764 2508
rect 811 2504 815 2527
rect 819 2527 834 2539
rect 819 2504 823 2527
rect 895 2504 899 2547
rect 915 2464 919 2546
rect 934 2531 938 2560
rect 929 2523 938 2531
rect 929 2464 933 2523
rect 954 2516 958 2580
rect 955 2504 958 2516
rect 949 2464 953 2504
rect 963 2482 967 2592
rect 979 2502 983 2616
rect 1025 2612 1029 2616
rect 995 2608 1029 2612
rect 961 2464 965 2470
rect 981 2464 985 2490
rect 995 2482 999 2608
rect 1033 2604 1037 2616
rect 1007 2600 1037 2604
rect 1019 2599 1037 2600
rect 1053 2595 1057 2616
rect 1033 2591 1057 2595
rect 1033 2496 1039 2591
rect 1063 2567 1067 2616
rect 1063 2509 1067 2555
rect 1085 2528 1089 2596
rect 1131 2559 1135 2616
rect 1191 2591 1195 2596
rect 1126 2547 1135 2559
rect 1087 2516 1089 2528
rect 1063 2503 1071 2509
rect 1085 2504 1089 2516
rect 1007 2470 1031 2472
rect 995 2468 1031 2470
rect 1027 2464 1031 2468
rect 1035 2464 1039 2496
rect 1055 2444 1059 2484
rect 1067 2474 1071 2503
rect 1063 2467 1071 2474
rect 1063 2444 1067 2467
rect 1131 2464 1135 2547
rect 1182 2584 1195 2591
rect 1182 2539 1186 2584
rect 1211 2573 1215 2596
rect 1206 2561 1215 2573
rect 1182 2516 1186 2527
rect 1182 2508 1200 2516
rect 1196 2504 1200 2508
rect 1204 2504 1208 2561
rect 1231 2519 1235 2596
rect 1291 2559 1295 2616
rect 1353 2576 1357 2596
rect 1286 2547 1295 2559
rect 1349 2569 1357 2576
rect 1363 2576 1367 2596
rect 1363 2569 1377 2576
rect 1349 2553 1355 2569
rect 1226 2507 1233 2519
rect 1226 2464 1230 2507
rect 1291 2464 1295 2547
rect 1346 2541 1355 2553
rect 1351 2464 1355 2541
rect 1371 2553 1377 2569
rect 1371 2541 1374 2553
rect 1371 2464 1375 2541
rect 1431 2528 1435 2596
rect 1453 2567 1457 2616
rect 1463 2595 1467 2616
rect 1483 2604 1487 2616
rect 1491 2612 1495 2616
rect 1491 2608 1525 2612
rect 1483 2600 1513 2604
rect 1483 2599 1501 2600
rect 1463 2591 1487 2595
rect 1431 2516 1433 2528
rect 1431 2504 1435 2516
rect 1453 2509 1457 2555
rect 1449 2503 1457 2509
rect 1449 2474 1453 2503
rect 1481 2496 1487 2591
rect 1449 2467 1457 2474
rect 1453 2444 1457 2467
rect 1461 2444 1465 2484
rect 1481 2464 1485 2496
rect 1521 2482 1525 2608
rect 1537 2502 1541 2616
rect 1559 2604 1563 2616
rect 1561 2592 1563 2604
rect 1569 2604 1573 2616
rect 1569 2592 1571 2604
rect 1489 2470 1513 2472
rect 1489 2468 1525 2470
rect 1489 2464 1493 2468
rect 1535 2464 1539 2490
rect 1553 2482 1557 2592
rect 1591 2584 1595 2616
rect 1562 2580 1595 2584
rect 1562 2516 1566 2580
rect 1582 2531 1586 2560
rect 1601 2558 1605 2616
rect 1621 2559 1625 2596
rect 1671 2591 1675 2596
rect 1662 2584 1675 2591
rect 1582 2523 1591 2531
rect 1562 2504 1565 2516
rect 1555 2464 1559 2470
rect 1567 2464 1571 2504
rect 1587 2464 1591 2523
rect 1601 2464 1605 2546
rect 1621 2504 1625 2547
rect 1662 2539 1666 2584
rect 1691 2573 1695 2596
rect 1686 2561 1695 2573
rect 1662 2516 1666 2527
rect 1662 2508 1680 2516
rect 1676 2504 1680 2508
rect 1684 2504 1688 2561
rect 1711 2519 1715 2596
rect 1771 2528 1775 2596
rect 1793 2567 1797 2616
rect 1803 2595 1807 2616
rect 1823 2604 1827 2616
rect 1831 2612 1835 2616
rect 1831 2608 1865 2612
rect 1823 2600 1853 2604
rect 1823 2599 1841 2600
rect 1803 2591 1827 2595
rect 1706 2507 1713 2519
rect 1771 2516 1773 2528
rect 1706 2464 1710 2507
rect 1771 2504 1775 2516
rect 1793 2509 1797 2555
rect 1789 2503 1797 2509
rect 1789 2474 1793 2503
rect 1821 2496 1827 2591
rect 1789 2467 1797 2474
rect 1793 2444 1797 2467
rect 1801 2444 1805 2484
rect 1821 2464 1825 2496
rect 1861 2482 1865 2608
rect 1877 2502 1881 2616
rect 1899 2604 1903 2616
rect 1901 2592 1903 2604
rect 1909 2604 1913 2616
rect 1909 2592 1911 2604
rect 1829 2470 1853 2472
rect 1829 2468 1865 2470
rect 1829 2464 1833 2468
rect 1875 2464 1879 2490
rect 1893 2482 1897 2592
rect 1931 2584 1935 2616
rect 1902 2580 1935 2584
rect 1902 2516 1906 2580
rect 1922 2531 1926 2560
rect 1941 2558 1945 2616
rect 1961 2559 1965 2596
rect 2011 2573 2015 2596
rect 2031 2573 2035 2596
rect 2051 2576 2055 2596
rect 2071 2576 2075 2596
rect 2091 2576 2095 2596
rect 2111 2576 2115 2596
rect 2131 2576 2135 2596
rect 2151 2576 2155 2596
rect 2011 2561 2014 2573
rect 2026 2561 2035 2573
rect 2062 2564 2075 2576
rect 2102 2564 2115 2576
rect 2142 2564 2155 2576
rect 1922 2523 1931 2531
rect 1902 2504 1905 2516
rect 1895 2464 1899 2470
rect 1907 2464 1911 2504
rect 1927 2464 1931 2523
rect 1941 2464 1945 2546
rect 1961 2504 1965 2547
rect 2011 2504 2015 2561
rect 2031 2504 2035 2561
rect 2051 2504 2055 2564
rect 2071 2504 2075 2564
rect 2091 2504 2095 2564
rect 2111 2504 2115 2564
rect 2131 2504 2135 2564
rect 2151 2504 2155 2564
rect 2215 2559 2219 2596
rect 2235 2558 2239 2616
rect 2245 2584 2249 2616
rect 2267 2604 2271 2616
rect 2269 2592 2271 2604
rect 2277 2604 2281 2616
rect 2277 2592 2279 2604
rect 2245 2580 2278 2584
rect 2215 2504 2219 2547
rect 2235 2464 2239 2546
rect 2254 2531 2258 2560
rect 2249 2523 2258 2531
rect 2249 2464 2253 2523
rect 2274 2516 2278 2580
rect 2275 2504 2278 2516
rect 2269 2464 2273 2504
rect 2283 2482 2287 2592
rect 2299 2502 2303 2616
rect 2345 2612 2349 2616
rect 2315 2608 2349 2612
rect 2281 2464 2285 2470
rect 2301 2464 2305 2490
rect 2315 2482 2319 2608
rect 2353 2604 2357 2616
rect 2327 2600 2357 2604
rect 2339 2599 2357 2600
rect 2373 2595 2377 2616
rect 2353 2591 2377 2595
rect 2353 2496 2359 2591
rect 2383 2567 2387 2616
rect 2383 2509 2387 2555
rect 2405 2528 2409 2596
rect 2473 2576 2477 2596
rect 2463 2569 2477 2576
rect 2483 2576 2487 2596
rect 2483 2569 2491 2576
rect 2463 2553 2469 2569
rect 2466 2541 2469 2553
rect 2407 2516 2409 2528
rect 2383 2503 2391 2509
rect 2405 2504 2409 2516
rect 2327 2470 2351 2472
rect 2315 2468 2351 2470
rect 2347 2464 2351 2468
rect 2355 2464 2359 2496
rect 2375 2444 2379 2484
rect 2387 2474 2391 2503
rect 2383 2467 2391 2474
rect 2383 2444 2387 2467
rect 2465 2464 2469 2541
rect 2485 2553 2491 2569
rect 2531 2559 2535 2616
rect 2485 2541 2494 2553
rect 2526 2547 2535 2559
rect 2485 2464 2489 2541
rect 2531 2464 2535 2547
rect 2605 2519 2609 2596
rect 2625 2573 2629 2596
rect 2645 2591 2649 2596
rect 2645 2584 2658 2591
rect 2625 2561 2634 2573
rect 2607 2507 2614 2519
rect 2610 2464 2614 2507
rect 2632 2504 2636 2561
rect 2654 2539 2658 2584
rect 2691 2559 2695 2616
rect 2773 2576 2777 2596
rect 2686 2547 2695 2559
rect 2763 2569 2777 2576
rect 2783 2576 2787 2596
rect 2783 2569 2791 2576
rect 2763 2553 2769 2569
rect 2654 2516 2658 2527
rect 2640 2508 2658 2516
rect 2640 2504 2644 2508
rect 2691 2464 2695 2547
rect 2766 2541 2769 2553
rect 2765 2464 2769 2541
rect 2785 2553 2791 2569
rect 2785 2541 2794 2553
rect 2785 2464 2789 2541
rect 2845 2519 2849 2596
rect 2865 2573 2869 2596
rect 2885 2591 2889 2596
rect 2885 2584 2898 2591
rect 2865 2561 2874 2573
rect 2847 2507 2854 2519
rect 2850 2464 2854 2507
rect 2872 2504 2876 2561
rect 2894 2539 2898 2584
rect 2931 2539 2935 2596
rect 2941 2553 2945 2596
rect 2961 2590 2965 2596
rect 3031 2591 3035 2596
rect 2967 2578 2979 2590
rect 2941 2541 2954 2553
rect 2926 2527 2935 2539
rect 2894 2516 2898 2527
rect 2880 2508 2898 2516
rect 2880 2504 2884 2508
rect 2931 2464 2935 2527
rect 2953 2464 2957 2541
rect 2975 2504 2979 2578
rect 3022 2584 3035 2591
rect 3022 2539 3026 2584
rect 3051 2573 3055 2596
rect 3046 2561 3055 2573
rect 3022 2516 3026 2527
rect 3022 2508 3040 2516
rect 3036 2504 3040 2508
rect 3044 2504 3048 2561
rect 3071 2519 3075 2596
rect 3153 2576 3157 2596
rect 3143 2569 3157 2576
rect 3163 2576 3167 2596
rect 3163 2569 3171 2576
rect 3143 2553 3149 2569
rect 3146 2541 3149 2553
rect 3066 2507 3073 2519
rect 3066 2464 3070 2507
rect 3145 2464 3149 2541
rect 3165 2553 3171 2569
rect 3165 2541 3174 2553
rect 3165 2464 3169 2541
rect 3211 2539 3215 2596
rect 3221 2553 3225 2596
rect 3241 2590 3245 2596
rect 3247 2578 3259 2590
rect 3221 2541 3234 2553
rect 3206 2527 3215 2539
rect 3211 2464 3215 2527
rect 3233 2464 3237 2541
rect 3255 2504 3259 2578
rect 3348 2519 3352 2576
rect 3325 2507 3333 2519
rect 3345 2507 3352 2519
rect 3325 2464 3329 2507
rect 3356 2499 3360 2576
rect 3364 2519 3368 2576
rect 3411 2559 3415 2616
rect 3473 2576 3477 2596
rect 3406 2547 3415 2559
rect 3469 2569 3477 2576
rect 3483 2576 3487 2596
rect 3483 2569 3497 2576
rect 3469 2553 3475 2569
rect 3364 2507 3374 2519
rect 3354 2480 3360 2487
rect 3345 2476 3360 2480
rect 3374 2476 3380 2507
rect 3345 2464 3349 2476
rect 3365 2472 3380 2476
rect 3365 2464 3369 2472
rect 3411 2464 3415 2547
rect 3466 2541 3475 2553
rect 3471 2464 3475 2541
rect 3491 2553 3497 2569
rect 3491 2541 3494 2553
rect 3491 2464 3495 2541
rect 3551 2539 3555 2596
rect 3561 2553 3565 2596
rect 3581 2590 3585 2596
rect 3587 2578 3599 2590
rect 3561 2541 3574 2553
rect 3546 2527 3555 2539
rect 3551 2464 3555 2527
rect 3573 2464 3577 2541
rect 3595 2504 3599 2578
rect 3651 2539 3655 2616
rect 3673 2590 3677 2596
rect 3675 2578 3677 2590
rect 3731 2559 3735 2616
rect 3815 2590 3819 2596
rect 3726 2547 3735 2559
rect 3646 2527 3655 2539
rect 3651 2464 3655 2527
rect 3675 2510 3677 2522
rect 3673 2504 3677 2510
rect 3731 2464 3735 2547
rect 3801 2578 3813 2590
rect 3801 2504 3805 2578
rect 3835 2553 3839 2596
rect 3826 2541 3839 2553
rect 3823 2464 3827 2541
rect 3845 2539 3849 2596
rect 3926 2591 3930 2596
rect 3900 2587 3930 2591
rect 3900 2539 3906 2587
rect 3934 2582 3938 2596
rect 3925 2575 3938 2582
rect 3925 2573 3929 2575
rect 3954 2573 3958 2596
rect 3962 2588 3966 2596
rect 3962 2581 3979 2588
rect 3927 2561 3929 2573
rect 3845 2527 3854 2539
rect 3906 2527 3909 2539
rect 3845 2464 3849 2527
rect 3905 2504 3909 2527
rect 3925 2504 3929 2561
rect 3954 2532 3958 2561
rect 3973 2539 3979 2581
rect 4033 2576 4037 2596
rect 4023 2569 4037 2576
rect 4043 2576 4047 2596
rect 4113 2576 4117 2596
rect 4043 2569 4051 2576
rect 4023 2553 4029 2569
rect 4026 2541 4029 2553
rect 3945 2526 3958 2532
rect 3965 2527 3973 2532
rect 3965 2526 3985 2527
rect 3945 2504 3949 2526
rect 3965 2504 3969 2526
rect 4025 2464 4029 2541
rect 4045 2553 4051 2569
rect 4103 2569 4117 2576
rect 4123 2576 4127 2596
rect 4171 2591 4175 2596
rect 4162 2584 4175 2591
rect 4123 2569 4131 2576
rect 4103 2553 4109 2569
rect 4045 2541 4054 2553
rect 4106 2541 4109 2553
rect 4045 2464 4049 2541
rect 4105 2464 4109 2541
rect 4125 2553 4131 2569
rect 4125 2541 4134 2553
rect 4125 2464 4129 2541
rect 4162 2539 4166 2584
rect 4191 2573 4195 2596
rect 4186 2561 4195 2573
rect 4162 2516 4166 2527
rect 4162 2508 4180 2516
rect 4176 2504 4180 2508
rect 4184 2504 4188 2561
rect 4211 2519 4215 2596
rect 4273 2576 4277 2596
rect 4269 2569 4277 2576
rect 4283 2576 4287 2596
rect 4554 2592 4558 2596
rect 4539 2586 4558 2592
rect 4283 2569 4297 2576
rect 4269 2553 4275 2569
rect 4266 2541 4275 2553
rect 4206 2507 4213 2519
rect 4206 2464 4210 2507
rect 4271 2464 4275 2541
rect 4291 2553 4297 2569
rect 4291 2541 4294 2553
rect 4291 2464 4295 2541
rect 4388 2519 4392 2576
rect 4365 2507 4373 2519
rect 4385 2507 4392 2519
rect 4365 2464 4369 2507
rect 4396 2499 4400 2576
rect 4404 2519 4408 2576
rect 4488 2519 4492 2576
rect 4404 2507 4414 2519
rect 4465 2507 4473 2519
rect 4485 2507 4492 2519
rect 4394 2480 4400 2487
rect 4385 2476 4400 2480
rect 4414 2476 4420 2507
rect 4385 2464 4389 2476
rect 4405 2472 4420 2476
rect 4405 2464 4409 2472
rect 4465 2464 4469 2507
rect 4496 2499 4500 2576
rect 4504 2519 4508 2576
rect 4539 2573 4546 2586
rect 4539 2524 4546 2561
rect 4562 2559 4566 2596
rect 4584 2573 4588 2616
rect 4586 2561 4595 2573
rect 4560 2524 4566 2547
rect 4504 2507 4514 2519
rect 4539 2518 4555 2524
rect 4560 2518 4575 2524
rect 4494 2480 4500 2487
rect 4485 2476 4500 2480
rect 4514 2476 4520 2507
rect 4551 2504 4555 2518
rect 4571 2504 4575 2518
rect 4591 2504 4595 2561
rect 4688 2519 4692 2576
rect 4665 2507 4673 2519
rect 4685 2507 4692 2519
rect 4485 2464 4489 2476
rect 4505 2472 4520 2476
rect 4505 2464 4509 2472
rect 4665 2464 4669 2507
rect 4696 2499 4700 2576
rect 4704 2519 4708 2576
rect 4704 2507 4714 2519
rect 4694 2480 4700 2487
rect 4685 2476 4700 2480
rect 4714 2476 4720 2507
rect 4685 2464 4689 2476
rect 4705 2472 4720 2476
rect 4705 2464 4709 2472
rect 35 2420 39 2424
rect 55 2420 59 2424
rect 69 2420 73 2424
rect 89 2420 93 2424
rect 101 2420 105 2424
rect 121 2420 125 2424
rect 167 2420 171 2424
rect 175 2420 179 2424
rect 195 2420 199 2424
rect 203 2420 207 2424
rect 225 2420 229 2424
rect 290 2420 294 2424
rect 312 2420 316 2424
rect 320 2420 324 2424
rect 371 2420 375 2424
rect 393 2420 397 2424
rect 451 2420 455 2424
rect 471 2420 475 2424
rect 550 2420 554 2424
rect 572 2420 576 2424
rect 580 2420 584 2424
rect 631 2420 635 2424
rect 653 2420 657 2424
rect 730 2420 734 2424
rect 752 2420 756 2424
rect 760 2420 764 2424
rect 811 2420 815 2424
rect 819 2420 823 2424
rect 895 2420 899 2424
rect 915 2420 919 2424
rect 929 2420 933 2424
rect 949 2420 953 2424
rect 961 2420 965 2424
rect 981 2420 985 2424
rect 1027 2420 1031 2424
rect 1035 2420 1039 2424
rect 1055 2420 1059 2424
rect 1063 2420 1067 2424
rect 1085 2420 1089 2424
rect 1131 2420 1135 2424
rect 1196 2420 1200 2424
rect 1204 2420 1208 2424
rect 1226 2420 1230 2424
rect 1291 2420 1295 2424
rect 1351 2420 1355 2424
rect 1371 2420 1375 2424
rect 1431 2420 1435 2424
rect 1453 2420 1457 2424
rect 1461 2420 1465 2424
rect 1481 2420 1485 2424
rect 1489 2420 1493 2424
rect 1535 2420 1539 2424
rect 1555 2420 1559 2424
rect 1567 2420 1571 2424
rect 1587 2420 1591 2424
rect 1601 2420 1605 2424
rect 1621 2420 1625 2424
rect 1676 2420 1680 2424
rect 1684 2420 1688 2424
rect 1706 2420 1710 2424
rect 1771 2420 1775 2424
rect 1793 2420 1797 2424
rect 1801 2420 1805 2424
rect 1821 2420 1825 2424
rect 1829 2420 1833 2424
rect 1875 2420 1879 2424
rect 1895 2420 1899 2424
rect 1907 2420 1911 2424
rect 1927 2420 1931 2424
rect 1941 2420 1945 2424
rect 1961 2420 1965 2424
rect 2011 2420 2015 2424
rect 2031 2420 2035 2424
rect 2051 2420 2055 2424
rect 2071 2420 2075 2424
rect 2091 2420 2095 2424
rect 2111 2420 2115 2424
rect 2131 2420 2135 2424
rect 2151 2420 2155 2424
rect 2215 2420 2219 2424
rect 2235 2420 2239 2424
rect 2249 2420 2253 2424
rect 2269 2420 2273 2424
rect 2281 2420 2285 2424
rect 2301 2420 2305 2424
rect 2347 2420 2351 2424
rect 2355 2420 2359 2424
rect 2375 2420 2379 2424
rect 2383 2420 2387 2424
rect 2405 2420 2409 2424
rect 2465 2420 2469 2424
rect 2485 2420 2489 2424
rect 2531 2420 2535 2424
rect 2610 2420 2614 2424
rect 2632 2420 2636 2424
rect 2640 2420 2644 2424
rect 2691 2420 2695 2424
rect 2765 2420 2769 2424
rect 2785 2420 2789 2424
rect 2850 2420 2854 2424
rect 2872 2420 2876 2424
rect 2880 2420 2884 2424
rect 2931 2420 2935 2424
rect 2953 2420 2957 2424
rect 2975 2420 2979 2424
rect 3036 2420 3040 2424
rect 3044 2420 3048 2424
rect 3066 2420 3070 2424
rect 3145 2420 3149 2424
rect 3165 2420 3169 2424
rect 3211 2420 3215 2424
rect 3233 2420 3237 2424
rect 3255 2420 3259 2424
rect 3325 2420 3329 2424
rect 3345 2420 3349 2424
rect 3365 2420 3369 2424
rect 3411 2420 3415 2424
rect 3471 2420 3475 2424
rect 3491 2420 3495 2424
rect 3551 2420 3555 2424
rect 3573 2420 3577 2424
rect 3595 2420 3599 2424
rect 3651 2420 3655 2424
rect 3673 2420 3677 2424
rect 3731 2420 3735 2424
rect 3801 2420 3805 2424
rect 3823 2420 3827 2424
rect 3845 2420 3849 2424
rect 3905 2420 3909 2424
rect 3925 2420 3929 2424
rect 3945 2420 3949 2424
rect 3965 2420 3969 2424
rect 4025 2420 4029 2424
rect 4045 2420 4049 2424
rect 4105 2420 4109 2424
rect 4125 2420 4129 2424
rect 4176 2420 4180 2424
rect 4184 2420 4188 2424
rect 4206 2420 4210 2424
rect 4271 2420 4275 2424
rect 4291 2420 4295 2424
rect 4365 2420 4369 2424
rect 4385 2420 4389 2424
rect 4405 2420 4409 2424
rect 4465 2420 4469 2424
rect 4485 2420 4489 2424
rect 4505 2420 4509 2424
rect 4551 2420 4555 2424
rect 4571 2420 4575 2424
rect 4591 2420 4595 2424
rect 4665 2420 4669 2424
rect 4685 2420 4689 2424
rect 4705 2420 4709 2424
rect 35 2396 39 2400
rect 55 2396 59 2400
rect 69 2396 73 2400
rect 89 2396 93 2400
rect 101 2396 105 2400
rect 121 2396 125 2400
rect 167 2396 171 2400
rect 175 2396 179 2400
rect 195 2396 199 2400
rect 203 2396 207 2400
rect 225 2396 229 2400
rect 276 2396 280 2400
rect 284 2396 288 2400
rect 306 2396 310 2400
rect 371 2396 375 2400
rect 391 2396 395 2400
rect 411 2396 415 2400
rect 431 2396 435 2400
rect 491 2396 495 2400
rect 513 2396 517 2400
rect 571 2396 575 2400
rect 591 2396 595 2400
rect 665 2396 669 2400
rect 711 2396 715 2400
rect 719 2396 723 2400
rect 805 2396 809 2400
rect 825 2396 829 2400
rect 845 2396 849 2400
rect 891 2396 895 2400
rect 899 2396 903 2400
rect 971 2396 975 2400
rect 979 2396 983 2400
rect 1051 2396 1055 2400
rect 1111 2396 1115 2400
rect 1133 2396 1137 2400
rect 1141 2396 1145 2400
rect 1161 2396 1165 2400
rect 1169 2396 1173 2400
rect 1215 2396 1219 2400
rect 1235 2396 1239 2400
rect 1247 2396 1251 2400
rect 1267 2396 1271 2400
rect 1281 2396 1285 2400
rect 1301 2396 1305 2400
rect 1356 2396 1360 2400
rect 1364 2396 1368 2400
rect 1386 2396 1390 2400
rect 1451 2396 1455 2400
rect 1473 2396 1477 2400
rect 1481 2396 1485 2400
rect 1501 2396 1505 2400
rect 1509 2396 1513 2400
rect 1555 2396 1559 2400
rect 1575 2396 1579 2400
rect 1587 2396 1591 2400
rect 1607 2396 1611 2400
rect 1621 2396 1625 2400
rect 1641 2396 1645 2400
rect 1717 2396 1721 2400
rect 1725 2396 1729 2400
rect 1785 2396 1789 2400
rect 1805 2396 1809 2400
rect 1825 2396 1829 2400
rect 1871 2396 1875 2400
rect 1957 2396 1961 2400
rect 1965 2396 1969 2400
rect 2011 2396 2015 2400
rect 2031 2396 2035 2400
rect 2051 2396 2055 2400
rect 2071 2396 2075 2400
rect 2091 2396 2095 2400
rect 2111 2396 2115 2400
rect 2131 2396 2135 2400
rect 2151 2396 2155 2400
rect 2216 2396 2220 2400
rect 2224 2396 2228 2400
rect 2246 2396 2250 2400
rect 2315 2396 2319 2400
rect 2335 2396 2339 2400
rect 2349 2396 2353 2400
rect 2369 2396 2373 2400
rect 2381 2396 2385 2400
rect 2401 2396 2405 2400
rect 2447 2396 2451 2400
rect 2455 2396 2459 2400
rect 2475 2396 2479 2400
rect 2483 2396 2487 2400
rect 2505 2396 2509 2400
rect 2565 2396 2569 2400
rect 2585 2396 2589 2400
rect 2631 2396 2635 2400
rect 2651 2396 2655 2400
rect 2711 2396 2715 2400
rect 2731 2396 2735 2400
rect 2810 2396 2814 2400
rect 2832 2396 2836 2400
rect 2840 2396 2844 2400
rect 2910 2396 2914 2400
rect 2932 2396 2936 2400
rect 2940 2396 2944 2400
rect 2995 2396 2999 2400
rect 3015 2396 3019 2400
rect 3029 2396 3033 2400
rect 3049 2396 3053 2400
rect 3061 2396 3065 2400
rect 3081 2396 3085 2400
rect 3127 2396 3131 2400
rect 3135 2396 3139 2400
rect 3155 2396 3159 2400
rect 3163 2396 3167 2400
rect 3185 2396 3189 2400
rect 3236 2396 3240 2400
rect 3244 2396 3248 2400
rect 3266 2396 3270 2400
rect 3331 2396 3335 2400
rect 3351 2396 3355 2400
rect 3411 2396 3415 2400
rect 3431 2396 3435 2400
rect 3505 2396 3509 2400
rect 3525 2396 3529 2400
rect 3585 2396 3589 2400
rect 3645 2396 3649 2400
rect 3705 2396 3709 2400
rect 3756 2396 3760 2400
rect 3764 2396 3768 2400
rect 3786 2396 3790 2400
rect 3863 2396 3867 2400
rect 3885 2396 3889 2400
rect 3931 2396 3935 2400
rect 3991 2396 3995 2400
rect 4013 2396 4017 2400
rect 4035 2396 4039 2400
rect 4110 2396 4114 2400
rect 4132 2396 4136 2400
rect 4140 2396 4144 2400
rect 4205 2396 4209 2400
rect 4225 2396 4229 2400
rect 4245 2396 4249 2400
rect 4291 2396 4295 2400
rect 4311 2396 4315 2400
rect 4331 2396 4335 2400
rect 4410 2396 4414 2400
rect 4432 2396 4436 2400
rect 4440 2396 4444 2400
rect 4496 2396 4500 2400
rect 4504 2396 4508 2400
rect 4526 2396 4530 2400
rect 4610 2396 4614 2400
rect 4632 2396 4636 2400
rect 4640 2396 4644 2400
rect 4691 2396 4695 2400
rect 4711 2396 4715 2400
rect 4731 2396 4735 2400
rect 35 2273 39 2316
rect 55 2274 59 2356
rect 69 2297 73 2356
rect 89 2316 93 2356
rect 101 2350 105 2356
rect 95 2304 98 2316
rect 69 2289 78 2297
rect 35 2224 39 2261
rect 55 2204 59 2262
rect 74 2260 78 2289
rect 94 2240 98 2304
rect 65 2236 98 2240
rect 65 2204 69 2236
rect 103 2228 107 2338
rect 121 2330 125 2356
rect 167 2352 171 2356
rect 135 2350 171 2352
rect 147 2348 171 2350
rect 89 2216 91 2228
rect 87 2204 91 2216
rect 97 2216 99 2228
rect 97 2204 101 2216
rect 119 2204 123 2318
rect 135 2212 139 2338
rect 175 2324 179 2356
rect 195 2336 199 2376
rect 203 2353 207 2376
rect 203 2346 211 2353
rect 173 2229 179 2324
rect 207 2317 211 2346
rect 203 2311 211 2317
rect 203 2265 207 2311
rect 225 2304 229 2316
rect 276 2312 280 2316
rect 227 2292 229 2304
rect 262 2304 280 2312
rect 262 2293 266 2304
rect 173 2225 197 2229
rect 159 2220 177 2221
rect 147 2216 177 2220
rect 135 2208 169 2212
rect 165 2204 169 2208
rect 173 2204 177 2216
rect 193 2204 197 2225
rect 203 2204 207 2253
rect 225 2224 229 2292
rect 262 2236 266 2281
rect 284 2259 288 2316
rect 306 2313 310 2356
rect 306 2301 313 2313
rect 286 2247 295 2259
rect 262 2229 275 2236
rect 271 2224 275 2229
rect 291 2224 295 2247
rect 311 2224 315 2301
rect 371 2294 375 2316
rect 391 2294 395 2316
rect 355 2293 375 2294
rect 367 2288 375 2293
rect 382 2288 395 2294
rect 361 2239 367 2281
rect 382 2259 386 2288
rect 411 2259 415 2316
rect 431 2293 435 2316
rect 491 2293 495 2356
rect 513 2310 517 2316
rect 515 2298 517 2310
rect 431 2281 434 2293
rect 486 2281 495 2293
rect 411 2247 413 2259
rect 361 2232 378 2239
rect 374 2224 378 2232
rect 382 2224 386 2247
rect 411 2245 415 2247
rect 402 2238 415 2245
rect 402 2224 406 2238
rect 434 2233 440 2281
rect 410 2229 440 2233
rect 410 2224 414 2229
rect 491 2204 495 2281
rect 571 2279 575 2356
rect 566 2267 575 2279
rect 569 2251 575 2267
rect 591 2279 595 2356
rect 591 2267 594 2279
rect 665 2273 669 2356
rect 711 2293 715 2316
rect 706 2281 715 2293
rect 719 2293 723 2316
rect 719 2281 734 2293
rect 591 2251 597 2267
rect 569 2244 577 2251
rect 515 2230 517 2242
rect 513 2224 517 2230
rect 573 2224 577 2244
rect 583 2244 597 2251
rect 665 2261 674 2273
rect 583 2224 587 2244
rect 665 2204 669 2261
rect 711 2204 715 2281
rect 731 2204 735 2281
rect 805 2259 809 2316
rect 825 2302 829 2316
rect 845 2302 849 2316
rect 825 2296 840 2302
rect 845 2296 861 2302
rect 834 2273 840 2296
rect 805 2247 814 2259
rect 812 2204 816 2247
rect 834 2224 838 2261
rect 854 2259 861 2296
rect 891 2293 895 2316
rect 886 2281 895 2293
rect 899 2293 903 2316
rect 971 2293 975 2316
rect 899 2281 914 2293
rect 966 2281 975 2293
rect 979 2293 983 2316
rect 979 2281 994 2293
rect 854 2234 861 2247
rect 842 2228 861 2234
rect 842 2224 846 2228
rect 891 2204 895 2281
rect 911 2204 915 2281
rect 971 2204 975 2281
rect 991 2204 995 2281
rect 1051 2273 1055 2356
rect 1133 2353 1137 2376
rect 1129 2346 1137 2353
rect 1129 2317 1133 2346
rect 1141 2336 1145 2376
rect 1161 2324 1165 2356
rect 1169 2352 1173 2356
rect 1169 2350 1205 2352
rect 1169 2348 1193 2350
rect 1046 2261 1055 2273
rect 1051 2204 1055 2261
rect 1111 2304 1115 2316
rect 1129 2311 1137 2317
rect 1111 2292 1113 2304
rect 1111 2224 1115 2292
rect 1133 2265 1137 2311
rect 1133 2204 1137 2253
rect 1161 2229 1167 2324
rect 1143 2225 1167 2229
rect 1143 2204 1147 2225
rect 1163 2220 1181 2221
rect 1163 2216 1193 2220
rect 1163 2204 1167 2216
rect 1201 2212 1205 2338
rect 1215 2330 1219 2356
rect 1235 2350 1239 2356
rect 1171 2208 1205 2212
rect 1171 2204 1175 2208
rect 1217 2204 1221 2318
rect 1233 2228 1237 2338
rect 1247 2316 1251 2356
rect 1242 2304 1245 2316
rect 1242 2240 1246 2304
rect 1267 2297 1271 2356
rect 1262 2289 1271 2297
rect 1262 2260 1266 2289
rect 1281 2274 1285 2356
rect 1301 2273 1305 2316
rect 1356 2312 1360 2316
rect 1342 2304 1360 2312
rect 1342 2293 1346 2304
rect 1242 2236 1275 2240
rect 1241 2216 1243 2228
rect 1239 2204 1243 2216
rect 1249 2216 1251 2228
rect 1249 2204 1253 2216
rect 1271 2204 1275 2236
rect 1281 2204 1285 2262
rect 1301 2224 1305 2261
rect 1342 2236 1346 2281
rect 1364 2259 1368 2316
rect 1386 2313 1390 2356
rect 1473 2353 1477 2376
rect 1469 2346 1477 2353
rect 1469 2317 1473 2346
rect 1481 2336 1485 2376
rect 1501 2324 1505 2356
rect 1509 2352 1513 2356
rect 1509 2350 1545 2352
rect 1509 2348 1533 2350
rect 1386 2301 1393 2313
rect 1451 2304 1455 2316
rect 1469 2311 1477 2317
rect 1366 2247 1375 2259
rect 1342 2229 1355 2236
rect 1351 2224 1355 2229
rect 1371 2224 1375 2247
rect 1391 2224 1395 2301
rect 1451 2292 1453 2304
rect 1451 2224 1455 2292
rect 1473 2265 1477 2311
rect 1473 2204 1477 2253
rect 1501 2229 1507 2324
rect 1483 2225 1507 2229
rect 1483 2204 1487 2225
rect 1503 2220 1521 2221
rect 1503 2216 1533 2220
rect 1503 2204 1507 2216
rect 1541 2212 1545 2338
rect 1555 2330 1559 2356
rect 1575 2350 1579 2356
rect 1511 2208 1545 2212
rect 1511 2204 1515 2208
rect 1557 2204 1561 2318
rect 1573 2228 1577 2338
rect 1587 2316 1591 2356
rect 1582 2304 1585 2316
rect 1582 2240 1586 2304
rect 1607 2297 1611 2356
rect 1602 2289 1611 2297
rect 1602 2260 1606 2289
rect 1621 2274 1625 2356
rect 1641 2273 1645 2316
rect 1717 2293 1721 2316
rect 1706 2281 1721 2293
rect 1725 2293 1729 2316
rect 1725 2281 1734 2293
rect 1582 2236 1615 2240
rect 1581 2216 1583 2228
rect 1579 2204 1583 2216
rect 1589 2216 1591 2228
rect 1589 2204 1593 2216
rect 1611 2204 1615 2236
rect 1621 2204 1625 2262
rect 1641 2224 1645 2261
rect 1705 2204 1709 2281
rect 1725 2204 1729 2281
rect 1785 2259 1789 2316
rect 1805 2302 1809 2316
rect 1825 2302 1829 2316
rect 1805 2296 1820 2302
rect 1825 2296 1841 2302
rect 1814 2273 1820 2296
rect 1785 2247 1794 2259
rect 1792 2204 1796 2247
rect 1814 2224 1818 2261
rect 1834 2259 1841 2296
rect 1871 2259 1875 2316
rect 1957 2293 1961 2316
rect 1946 2281 1961 2293
rect 1965 2293 1969 2316
rect 1965 2281 1974 2293
rect 1866 2247 1875 2259
rect 1834 2234 1841 2247
rect 1822 2228 1841 2234
rect 1822 2224 1826 2228
rect 1871 2224 1875 2247
rect 1945 2204 1949 2281
rect 1965 2204 1969 2281
rect 2011 2259 2015 2316
rect 2031 2259 2035 2316
rect 2011 2247 2014 2259
rect 2026 2247 2035 2259
rect 2051 2256 2055 2316
rect 2071 2256 2075 2316
rect 2091 2256 2095 2316
rect 2111 2256 2115 2316
rect 2131 2256 2135 2316
rect 2151 2256 2155 2316
rect 2216 2312 2220 2316
rect 2202 2304 2220 2312
rect 2202 2293 2206 2304
rect 2011 2224 2015 2247
rect 2031 2224 2035 2247
rect 2062 2244 2075 2256
rect 2102 2244 2115 2256
rect 2142 2244 2155 2256
rect 2051 2224 2055 2244
rect 2071 2224 2075 2244
rect 2091 2224 2095 2244
rect 2111 2224 2115 2244
rect 2131 2224 2135 2244
rect 2151 2224 2155 2244
rect 2202 2236 2206 2281
rect 2224 2259 2228 2316
rect 2246 2313 2250 2356
rect 2246 2301 2253 2313
rect 2226 2247 2235 2259
rect 2202 2229 2215 2236
rect 2211 2224 2215 2229
rect 2231 2224 2235 2247
rect 2251 2224 2255 2301
rect 2315 2273 2319 2316
rect 2335 2274 2339 2356
rect 2349 2297 2353 2356
rect 2369 2316 2373 2356
rect 2381 2350 2385 2356
rect 2375 2304 2378 2316
rect 2349 2289 2358 2297
rect 2315 2224 2319 2261
rect 2335 2204 2339 2262
rect 2354 2260 2358 2289
rect 2374 2240 2378 2304
rect 2345 2236 2378 2240
rect 2345 2204 2349 2236
rect 2383 2228 2387 2338
rect 2401 2330 2405 2356
rect 2447 2352 2451 2356
rect 2415 2350 2451 2352
rect 2427 2348 2451 2350
rect 2369 2216 2371 2228
rect 2367 2204 2371 2216
rect 2377 2216 2379 2228
rect 2377 2204 2381 2216
rect 2399 2204 2403 2318
rect 2415 2212 2419 2338
rect 2455 2324 2459 2356
rect 2475 2336 2479 2376
rect 2483 2353 2487 2376
rect 2483 2346 2491 2353
rect 2453 2229 2459 2324
rect 2487 2317 2491 2346
rect 2483 2311 2491 2317
rect 2483 2265 2487 2311
rect 2505 2304 2509 2316
rect 2507 2292 2509 2304
rect 2453 2225 2477 2229
rect 2439 2220 2457 2221
rect 2427 2216 2457 2220
rect 2415 2208 2449 2212
rect 2445 2204 2449 2208
rect 2453 2204 2457 2216
rect 2473 2204 2477 2225
rect 2483 2204 2487 2253
rect 2505 2224 2509 2292
rect 2565 2279 2569 2356
rect 2566 2267 2569 2279
rect 2563 2251 2569 2267
rect 2585 2279 2589 2356
rect 2631 2279 2635 2356
rect 2585 2267 2594 2279
rect 2626 2267 2635 2279
rect 2585 2251 2591 2267
rect 2563 2244 2577 2251
rect 2573 2224 2577 2244
rect 2583 2244 2591 2251
rect 2629 2251 2635 2267
rect 2651 2279 2655 2356
rect 2711 2279 2715 2356
rect 2651 2267 2654 2279
rect 2706 2267 2715 2279
rect 2651 2251 2657 2267
rect 2629 2244 2637 2251
rect 2583 2224 2587 2244
rect 2633 2224 2637 2244
rect 2643 2244 2657 2251
rect 2709 2251 2715 2267
rect 2731 2279 2735 2356
rect 2810 2313 2814 2356
rect 2807 2301 2814 2313
rect 2731 2267 2734 2279
rect 2731 2251 2737 2267
rect 2709 2244 2717 2251
rect 2643 2224 2647 2244
rect 2713 2224 2717 2244
rect 2723 2244 2737 2251
rect 2723 2224 2727 2244
rect 2805 2224 2809 2301
rect 2832 2259 2836 2316
rect 2840 2312 2844 2316
rect 2910 2313 2914 2356
rect 2840 2304 2858 2312
rect 2854 2293 2858 2304
rect 2907 2301 2914 2313
rect 2825 2247 2834 2259
rect 2825 2224 2829 2247
rect 2854 2236 2858 2281
rect 2845 2229 2858 2236
rect 2845 2224 2849 2229
rect 2905 2224 2909 2301
rect 2932 2259 2936 2316
rect 2940 2312 2944 2316
rect 2940 2304 2958 2312
rect 2954 2293 2958 2304
rect 2925 2247 2934 2259
rect 2925 2224 2929 2247
rect 2954 2236 2958 2281
rect 2995 2273 2999 2316
rect 3015 2274 3019 2356
rect 3029 2297 3033 2356
rect 3049 2316 3053 2356
rect 3061 2350 3065 2356
rect 3055 2304 3058 2316
rect 3029 2289 3038 2297
rect 2945 2229 2958 2236
rect 2945 2224 2949 2229
rect 2995 2224 2999 2261
rect 3015 2204 3019 2262
rect 3034 2260 3038 2289
rect 3054 2240 3058 2304
rect 3025 2236 3058 2240
rect 3025 2204 3029 2236
rect 3063 2228 3067 2338
rect 3081 2330 3085 2356
rect 3127 2352 3131 2356
rect 3095 2350 3131 2352
rect 3107 2348 3131 2350
rect 3049 2216 3051 2228
rect 3047 2204 3051 2216
rect 3057 2216 3059 2228
rect 3057 2204 3061 2216
rect 3079 2204 3083 2318
rect 3095 2212 3099 2338
rect 3135 2324 3139 2356
rect 3155 2336 3159 2376
rect 3163 2353 3167 2376
rect 3163 2346 3171 2353
rect 3133 2229 3139 2324
rect 3167 2317 3171 2346
rect 3163 2311 3171 2317
rect 3163 2265 3167 2311
rect 3185 2304 3189 2316
rect 3236 2312 3240 2316
rect 3187 2292 3189 2304
rect 3222 2304 3240 2312
rect 3222 2293 3226 2304
rect 3133 2225 3157 2229
rect 3119 2220 3137 2221
rect 3107 2216 3137 2220
rect 3095 2208 3129 2212
rect 3125 2204 3129 2208
rect 3133 2204 3137 2216
rect 3153 2204 3157 2225
rect 3163 2204 3167 2253
rect 3185 2224 3189 2292
rect 3222 2236 3226 2281
rect 3244 2259 3248 2316
rect 3266 2313 3270 2356
rect 3266 2301 3273 2313
rect 3246 2247 3255 2259
rect 3222 2229 3235 2236
rect 3231 2224 3235 2229
rect 3251 2224 3255 2247
rect 3271 2224 3275 2301
rect 3331 2279 3335 2356
rect 3326 2267 3335 2279
rect 3329 2251 3335 2267
rect 3351 2279 3355 2356
rect 3411 2279 3415 2356
rect 3351 2267 3354 2279
rect 3406 2267 3415 2279
rect 3351 2251 3357 2267
rect 3329 2244 3337 2251
rect 3333 2224 3337 2244
rect 3343 2244 3357 2251
rect 3409 2251 3415 2267
rect 3431 2279 3435 2356
rect 3505 2279 3509 2356
rect 3431 2267 3434 2279
rect 3506 2267 3509 2279
rect 3431 2251 3437 2267
rect 3409 2244 3417 2251
rect 3343 2224 3347 2244
rect 3413 2224 3417 2244
rect 3423 2244 3437 2251
rect 3503 2251 3509 2267
rect 3525 2279 3529 2356
rect 3525 2267 3534 2279
rect 3525 2251 3531 2267
rect 3503 2244 3517 2251
rect 3423 2224 3427 2244
rect 3513 2224 3517 2244
rect 3523 2244 3531 2251
rect 3585 2259 3589 2316
rect 3645 2259 3649 2316
rect 3705 2273 3709 2356
rect 3756 2312 3760 2316
rect 3742 2304 3760 2312
rect 3742 2293 3746 2304
rect 3705 2261 3714 2273
rect 3585 2247 3594 2259
rect 3645 2247 3654 2259
rect 3523 2224 3527 2244
rect 3585 2224 3589 2247
rect 3645 2224 3649 2247
rect 3705 2204 3709 2261
rect 3742 2236 3746 2281
rect 3764 2259 3768 2316
rect 3786 2313 3790 2356
rect 3786 2301 3793 2313
rect 3863 2310 3867 2316
rect 3766 2247 3775 2259
rect 3742 2229 3755 2236
rect 3751 2224 3755 2229
rect 3771 2224 3775 2247
rect 3791 2224 3795 2301
rect 3863 2298 3865 2310
rect 3885 2293 3889 2356
rect 3885 2281 3894 2293
rect 3863 2230 3865 2242
rect 3863 2224 3867 2230
rect 3885 2204 3889 2281
rect 3931 2259 3935 2316
rect 3991 2293 3995 2356
rect 3986 2281 3995 2293
rect 3926 2247 3935 2259
rect 3931 2224 3935 2247
rect 3991 2224 3995 2281
rect 4013 2279 4017 2356
rect 4001 2267 4014 2279
rect 4001 2224 4005 2267
rect 4035 2242 4039 2316
rect 4110 2313 4114 2356
rect 4107 2301 4114 2313
rect 4027 2230 4039 2242
rect 4021 2224 4025 2230
rect 4105 2224 4109 2301
rect 4132 2259 4136 2316
rect 4140 2312 4144 2316
rect 4205 2313 4209 2356
rect 4225 2344 4229 2356
rect 4245 2348 4249 2356
rect 4245 2344 4260 2348
rect 4225 2340 4240 2344
rect 4234 2333 4240 2340
rect 4140 2304 4158 2312
rect 4154 2293 4158 2304
rect 4205 2301 4213 2313
rect 4225 2301 4232 2313
rect 4125 2247 4134 2259
rect 4125 2224 4129 2247
rect 4154 2236 4158 2281
rect 4228 2244 4232 2301
rect 4236 2244 4240 2321
rect 4254 2313 4260 2344
rect 4244 2301 4254 2313
rect 4291 2302 4295 2316
rect 4311 2302 4315 2316
rect 4244 2244 4248 2301
rect 4279 2296 4295 2302
rect 4300 2296 4315 2302
rect 4279 2259 4286 2296
rect 4300 2273 4306 2296
rect 4145 2229 4158 2236
rect 4145 2224 4149 2229
rect 4279 2234 4286 2247
rect 4279 2228 4298 2234
rect 4294 2224 4298 2228
rect 4302 2224 4306 2261
rect 4331 2259 4335 2316
rect 4410 2313 4414 2356
rect 4407 2301 4414 2313
rect 4326 2247 4335 2259
rect 4324 2204 4328 2247
rect 4405 2224 4409 2301
rect 4432 2259 4436 2316
rect 4440 2312 4444 2316
rect 4496 2312 4500 2316
rect 4440 2304 4458 2312
rect 4454 2293 4458 2304
rect 4482 2304 4500 2312
rect 4482 2293 4486 2304
rect 4425 2247 4434 2259
rect 4425 2224 4429 2247
rect 4454 2236 4458 2281
rect 4445 2229 4458 2236
rect 4482 2236 4486 2281
rect 4504 2259 4508 2316
rect 4526 2313 4530 2356
rect 4610 2313 4614 2356
rect 4526 2301 4533 2313
rect 4607 2301 4614 2313
rect 4506 2247 4515 2259
rect 4482 2229 4495 2236
rect 4445 2224 4449 2229
rect 4491 2224 4495 2229
rect 4511 2224 4515 2247
rect 4531 2224 4535 2301
rect 4605 2224 4609 2301
rect 4632 2259 4636 2316
rect 4640 2312 4644 2316
rect 4640 2304 4658 2312
rect 4654 2293 4658 2304
rect 4691 2302 4695 2316
rect 4711 2302 4715 2316
rect 4679 2296 4695 2302
rect 4700 2296 4715 2302
rect 4625 2247 4634 2259
rect 4625 2224 4629 2247
rect 4654 2236 4658 2281
rect 4679 2259 4686 2296
rect 4700 2273 4706 2296
rect 4645 2229 4658 2236
rect 4679 2234 4686 2247
rect 4645 2224 4649 2229
rect 4679 2228 4698 2234
rect 4694 2224 4698 2228
rect 4702 2224 4706 2261
rect 4731 2259 4735 2316
rect 4726 2247 4735 2259
rect 4724 2204 4728 2247
rect 35 2180 39 2184
rect 55 2180 59 2184
rect 65 2180 69 2184
rect 87 2180 91 2184
rect 97 2180 101 2184
rect 119 2180 123 2184
rect 165 2180 169 2184
rect 173 2180 177 2184
rect 193 2180 197 2184
rect 203 2180 207 2184
rect 225 2180 229 2184
rect 271 2180 275 2184
rect 291 2180 295 2184
rect 311 2180 315 2184
rect 374 2180 378 2184
rect 382 2180 386 2184
rect 402 2180 406 2184
rect 410 2180 414 2184
rect 491 2180 495 2184
rect 513 2180 517 2184
rect 573 2180 577 2184
rect 583 2180 587 2184
rect 665 2180 669 2184
rect 711 2180 715 2184
rect 731 2180 735 2184
rect 812 2180 816 2184
rect 834 2180 838 2184
rect 842 2180 846 2184
rect 891 2180 895 2184
rect 911 2180 915 2184
rect 971 2180 975 2184
rect 991 2180 995 2184
rect 1051 2180 1055 2184
rect 1111 2180 1115 2184
rect 1133 2180 1137 2184
rect 1143 2180 1147 2184
rect 1163 2180 1167 2184
rect 1171 2180 1175 2184
rect 1217 2180 1221 2184
rect 1239 2180 1243 2184
rect 1249 2180 1253 2184
rect 1271 2180 1275 2184
rect 1281 2180 1285 2184
rect 1301 2180 1305 2184
rect 1351 2180 1355 2184
rect 1371 2180 1375 2184
rect 1391 2180 1395 2184
rect 1451 2180 1455 2184
rect 1473 2180 1477 2184
rect 1483 2180 1487 2184
rect 1503 2180 1507 2184
rect 1511 2180 1515 2184
rect 1557 2180 1561 2184
rect 1579 2180 1583 2184
rect 1589 2180 1593 2184
rect 1611 2180 1615 2184
rect 1621 2180 1625 2184
rect 1641 2180 1645 2184
rect 1705 2180 1709 2184
rect 1725 2180 1729 2184
rect 1792 2180 1796 2184
rect 1814 2180 1818 2184
rect 1822 2180 1826 2184
rect 1871 2180 1875 2184
rect 1945 2180 1949 2184
rect 1965 2180 1969 2184
rect 2011 2180 2015 2184
rect 2031 2180 2035 2184
rect 2051 2180 2055 2184
rect 2071 2180 2075 2184
rect 2091 2180 2095 2184
rect 2111 2180 2115 2184
rect 2131 2180 2135 2184
rect 2151 2180 2155 2184
rect 2211 2180 2215 2184
rect 2231 2180 2235 2184
rect 2251 2180 2255 2184
rect 2315 2180 2319 2184
rect 2335 2180 2339 2184
rect 2345 2180 2349 2184
rect 2367 2180 2371 2184
rect 2377 2180 2381 2184
rect 2399 2180 2403 2184
rect 2445 2180 2449 2184
rect 2453 2180 2457 2184
rect 2473 2180 2477 2184
rect 2483 2180 2487 2184
rect 2505 2180 2509 2184
rect 2573 2180 2577 2184
rect 2583 2180 2587 2184
rect 2633 2180 2637 2184
rect 2643 2180 2647 2184
rect 2713 2180 2717 2184
rect 2723 2180 2727 2184
rect 2805 2180 2809 2184
rect 2825 2180 2829 2184
rect 2845 2180 2849 2184
rect 2905 2180 2909 2184
rect 2925 2180 2929 2184
rect 2945 2180 2949 2184
rect 2995 2180 2999 2184
rect 3015 2180 3019 2184
rect 3025 2180 3029 2184
rect 3047 2180 3051 2184
rect 3057 2180 3061 2184
rect 3079 2180 3083 2184
rect 3125 2180 3129 2184
rect 3133 2180 3137 2184
rect 3153 2180 3157 2184
rect 3163 2180 3167 2184
rect 3185 2180 3189 2184
rect 3231 2180 3235 2184
rect 3251 2180 3255 2184
rect 3271 2180 3275 2184
rect 3333 2180 3337 2184
rect 3343 2180 3347 2184
rect 3413 2180 3417 2184
rect 3423 2180 3427 2184
rect 3513 2180 3517 2184
rect 3523 2180 3527 2184
rect 3585 2180 3589 2184
rect 3645 2180 3649 2184
rect 3705 2180 3709 2184
rect 3751 2180 3755 2184
rect 3771 2180 3775 2184
rect 3791 2180 3795 2184
rect 3863 2180 3867 2184
rect 3885 2180 3889 2184
rect 3931 2180 3935 2184
rect 3991 2180 3995 2184
rect 4001 2180 4005 2184
rect 4021 2180 4025 2184
rect 4105 2180 4109 2184
rect 4125 2180 4129 2184
rect 4145 2180 4149 2184
rect 4228 2180 4232 2184
rect 4236 2180 4240 2184
rect 4244 2180 4248 2184
rect 4294 2180 4298 2184
rect 4302 2180 4306 2184
rect 4324 2180 4328 2184
rect 4405 2180 4409 2184
rect 4425 2180 4429 2184
rect 4445 2180 4449 2184
rect 4491 2180 4495 2184
rect 4511 2180 4515 2184
rect 4531 2180 4535 2184
rect 4605 2180 4609 2184
rect 4625 2180 4629 2184
rect 4645 2180 4649 2184
rect 4694 2180 4698 2184
rect 4702 2180 4706 2184
rect 4724 2180 4728 2184
rect 31 2156 35 2160
rect 51 2156 55 2160
rect 71 2156 75 2160
rect 91 2156 95 2160
rect 111 2156 115 2160
rect 131 2156 135 2160
rect 151 2156 155 2160
rect 171 2156 175 2160
rect 253 2156 257 2160
rect 263 2156 267 2160
rect 325 2156 329 2160
rect 345 2156 349 2160
rect 365 2156 369 2160
rect 414 2156 418 2160
rect 422 2156 426 2160
rect 442 2156 446 2160
rect 450 2156 454 2160
rect 535 2156 539 2160
rect 555 2156 559 2160
rect 565 2156 569 2160
rect 587 2156 591 2160
rect 597 2156 601 2160
rect 619 2156 623 2160
rect 665 2156 669 2160
rect 673 2156 677 2160
rect 693 2156 697 2160
rect 703 2156 707 2160
rect 725 2156 729 2160
rect 793 2156 797 2160
rect 803 2156 807 2160
rect 865 2156 869 2160
rect 885 2156 889 2160
rect 905 2156 909 2160
rect 953 2156 957 2160
rect 963 2156 967 2160
rect 1031 2156 1035 2160
rect 1051 2156 1055 2160
rect 1111 2156 1115 2160
rect 1131 2156 1135 2160
rect 1151 2156 1155 2160
rect 1213 2156 1217 2160
rect 1223 2156 1227 2160
rect 1291 2156 1295 2160
rect 1311 2156 1315 2160
rect 1371 2156 1375 2160
rect 1393 2156 1397 2160
rect 1403 2156 1407 2160
rect 1423 2156 1427 2160
rect 1431 2156 1435 2160
rect 1477 2156 1481 2160
rect 1499 2156 1503 2160
rect 1509 2156 1513 2160
rect 1531 2156 1535 2160
rect 1541 2156 1545 2160
rect 1561 2156 1565 2160
rect 1632 2156 1636 2160
rect 1654 2156 1658 2160
rect 1662 2156 1666 2160
rect 1723 2156 1727 2160
rect 1745 2156 1749 2160
rect 1791 2156 1795 2160
rect 1813 2156 1817 2160
rect 1823 2156 1827 2160
rect 1843 2156 1847 2160
rect 1851 2156 1855 2160
rect 1897 2156 1901 2160
rect 1919 2156 1923 2160
rect 1929 2156 1933 2160
rect 1951 2156 1955 2160
rect 1961 2156 1965 2160
rect 1981 2156 1985 2160
rect 2045 2156 2049 2160
rect 2113 2156 2117 2160
rect 2123 2156 2127 2160
rect 2171 2156 2175 2160
rect 2193 2156 2197 2160
rect 2253 2156 2257 2160
rect 2263 2156 2267 2160
rect 2345 2156 2349 2160
rect 2365 2156 2369 2160
rect 2385 2156 2389 2160
rect 2453 2156 2457 2160
rect 2463 2156 2467 2160
rect 2533 2156 2537 2160
rect 2543 2156 2547 2160
rect 2605 2156 2609 2160
rect 2625 2156 2629 2160
rect 2645 2156 2649 2160
rect 2705 2156 2709 2160
rect 2725 2156 2729 2160
rect 2745 2156 2749 2160
rect 2795 2156 2799 2160
rect 2815 2156 2819 2160
rect 2825 2156 2829 2160
rect 2847 2156 2851 2160
rect 2857 2156 2861 2160
rect 2879 2156 2883 2160
rect 2925 2156 2929 2160
rect 2933 2156 2937 2160
rect 2953 2156 2957 2160
rect 2963 2156 2967 2160
rect 2985 2156 2989 2160
rect 3031 2156 3035 2160
rect 3041 2156 3045 2160
rect 3061 2156 3065 2160
rect 3145 2156 3149 2160
rect 3165 2156 3169 2160
rect 3185 2156 3189 2160
rect 3245 2156 3249 2160
rect 3265 2156 3269 2160
rect 3285 2156 3289 2160
rect 3333 2156 3337 2160
rect 3343 2156 3347 2160
rect 3425 2156 3429 2160
rect 3445 2156 3449 2160
rect 3465 2156 3469 2160
rect 3512 2156 3516 2160
rect 3520 2156 3524 2160
rect 3528 2156 3532 2160
rect 3611 2156 3615 2160
rect 3672 2156 3676 2160
rect 3680 2156 3684 2160
rect 3688 2156 3692 2160
rect 3773 2156 3777 2160
rect 3783 2156 3787 2160
rect 3851 2156 3855 2160
rect 3873 2156 3877 2160
rect 3931 2156 3935 2160
rect 3951 2156 3955 2160
rect 3971 2156 3975 2160
rect 4053 2156 4057 2160
rect 4063 2156 4067 2160
rect 4133 2156 4137 2160
rect 4143 2156 4147 2160
rect 4213 2156 4217 2160
rect 4223 2156 4227 2160
rect 4271 2156 4275 2160
rect 4281 2156 4285 2160
rect 4301 2156 4305 2160
rect 4374 2156 4378 2160
rect 4382 2156 4386 2160
rect 4404 2156 4408 2160
rect 4492 2156 4496 2160
rect 4514 2156 4518 2160
rect 4522 2156 4526 2160
rect 4572 2156 4576 2160
rect 4580 2156 4584 2160
rect 4588 2156 4592 2160
rect 4672 2156 4676 2160
rect 4680 2156 4684 2160
rect 4688 2156 4692 2160
rect 31 2093 35 2116
rect 51 2093 55 2116
rect 71 2096 75 2116
rect 91 2096 95 2116
rect 111 2096 115 2116
rect 131 2096 135 2116
rect 151 2096 155 2116
rect 171 2096 175 2116
rect 253 2096 257 2116
rect 31 2081 34 2093
rect 46 2081 55 2093
rect 82 2084 95 2096
rect 122 2084 135 2096
rect 162 2084 175 2096
rect 31 2024 35 2081
rect 51 2024 55 2081
rect 71 2024 75 2084
rect 91 2024 95 2084
rect 111 2024 115 2084
rect 131 2024 135 2084
rect 151 2024 155 2084
rect 171 2024 175 2084
rect 243 2089 257 2096
rect 263 2096 267 2116
rect 263 2089 271 2096
rect 243 2073 249 2089
rect 246 2061 249 2073
rect 245 1984 249 2061
rect 265 2073 271 2089
rect 265 2061 274 2073
rect 265 1984 269 2061
rect 325 2039 329 2116
rect 345 2093 349 2116
rect 365 2111 369 2116
rect 365 2104 378 2111
rect 414 2108 418 2116
rect 345 2081 354 2093
rect 327 2027 334 2039
rect 330 1984 334 2027
rect 352 2024 356 2081
rect 374 2059 378 2104
rect 401 2101 418 2108
rect 401 2059 407 2101
rect 422 2093 426 2116
rect 442 2102 446 2116
rect 450 2111 454 2116
rect 450 2107 480 2111
rect 442 2095 455 2102
rect 451 2093 455 2095
rect 451 2081 453 2093
rect 422 2052 426 2081
rect 407 2047 415 2052
rect 374 2036 378 2047
rect 395 2046 415 2047
rect 422 2046 435 2052
rect 360 2028 378 2036
rect 360 2024 364 2028
rect 411 2024 415 2046
rect 431 2024 435 2046
rect 451 2024 455 2081
rect 474 2059 480 2107
rect 535 2079 539 2116
rect 555 2078 559 2136
rect 565 2104 569 2136
rect 587 2124 591 2136
rect 589 2112 591 2124
rect 597 2124 601 2136
rect 597 2112 599 2124
rect 565 2100 598 2104
rect 471 2047 474 2059
rect 471 2024 475 2047
rect 535 2024 539 2067
rect 555 1984 559 2066
rect 574 2051 578 2080
rect 569 2043 578 2051
rect 569 1984 573 2043
rect 594 2036 598 2100
rect 595 2024 598 2036
rect 589 1984 593 2024
rect 603 2002 607 2112
rect 619 2022 623 2136
rect 665 2132 669 2136
rect 635 2128 669 2132
rect 601 1984 605 1990
rect 621 1984 625 2010
rect 635 2002 639 2128
rect 673 2124 677 2136
rect 647 2120 677 2124
rect 659 2119 677 2120
rect 693 2115 697 2136
rect 673 2111 697 2115
rect 673 2016 679 2111
rect 703 2087 707 2136
rect 885 2129 889 2136
rect 905 2129 909 2136
rect 885 2123 899 2129
rect 905 2124 918 2129
rect 703 2029 707 2075
rect 725 2048 729 2116
rect 793 2096 797 2116
rect 783 2089 797 2096
rect 803 2096 807 2116
rect 865 2108 869 2116
rect 865 2096 875 2108
rect 803 2089 811 2096
rect 783 2073 789 2089
rect 786 2061 789 2073
rect 727 2036 729 2048
rect 703 2023 711 2029
rect 725 2024 729 2036
rect 647 1990 671 1992
rect 635 1988 671 1990
rect 667 1984 671 1988
rect 675 1984 679 2016
rect 695 1964 699 2004
rect 707 1994 711 2023
rect 703 1987 711 1994
rect 703 1964 707 1987
rect 785 1984 789 2061
rect 805 2073 811 2089
rect 805 2061 814 2073
rect 805 1984 809 2061
rect 895 2059 899 2123
rect 914 2079 918 2124
rect 953 2096 957 2116
rect 949 2089 957 2096
rect 963 2096 967 2116
rect 963 2089 977 2096
rect 949 2073 955 2089
rect 875 2024 879 2029
rect 895 2024 899 2047
rect 914 2033 918 2067
rect 946 2061 955 2073
rect 905 2028 918 2033
rect 905 2024 909 2028
rect 951 1984 955 2061
rect 971 2073 977 2089
rect 971 2061 974 2073
rect 971 1984 975 2061
rect 1031 2059 1035 2136
rect 1051 2059 1055 2136
rect 1111 2111 1115 2116
rect 1102 2104 1115 2111
rect 1102 2059 1106 2104
rect 1131 2093 1135 2116
rect 1126 2081 1135 2093
rect 1026 2047 1035 2059
rect 1031 2024 1035 2047
rect 1039 2047 1054 2059
rect 1039 2024 1043 2047
rect 1102 2036 1106 2047
rect 1102 2028 1120 2036
rect 1116 2024 1120 2028
rect 1124 2024 1128 2081
rect 1151 2039 1155 2116
rect 1213 2096 1217 2116
rect 1209 2089 1217 2096
rect 1223 2096 1227 2116
rect 1223 2089 1237 2096
rect 1209 2073 1215 2089
rect 1206 2061 1215 2073
rect 1146 2027 1153 2039
rect 1146 1984 1150 2027
rect 1211 1984 1215 2061
rect 1231 2073 1237 2089
rect 1231 2061 1234 2073
rect 1231 1984 1235 2061
rect 1291 2059 1295 2136
rect 1311 2059 1315 2136
rect 1286 2047 1295 2059
rect 1291 2024 1295 2047
rect 1299 2047 1314 2059
rect 1371 2048 1375 2116
rect 1393 2087 1397 2136
rect 1403 2115 1407 2136
rect 1423 2124 1427 2136
rect 1431 2132 1435 2136
rect 1431 2128 1465 2132
rect 1423 2120 1453 2124
rect 1423 2119 1441 2120
rect 1403 2111 1427 2115
rect 1299 2024 1303 2047
rect 1371 2036 1373 2048
rect 1371 2024 1375 2036
rect 1393 2029 1397 2075
rect 1389 2023 1397 2029
rect 1389 1994 1393 2023
rect 1421 2016 1427 2111
rect 1389 1987 1397 1994
rect 1393 1964 1397 1987
rect 1401 1964 1405 2004
rect 1421 1984 1425 2016
rect 1461 2002 1465 2128
rect 1477 2022 1481 2136
rect 1499 2124 1503 2136
rect 1501 2112 1503 2124
rect 1509 2124 1513 2136
rect 1509 2112 1511 2124
rect 1429 1990 1453 1992
rect 1429 1988 1465 1990
rect 1429 1984 1433 1988
rect 1475 1984 1479 2010
rect 1493 2002 1497 2112
rect 1531 2104 1535 2136
rect 1502 2100 1535 2104
rect 1502 2036 1506 2100
rect 1522 2051 1526 2080
rect 1541 2078 1545 2136
rect 1561 2079 1565 2116
rect 1632 2093 1636 2136
rect 1625 2081 1634 2093
rect 1522 2043 1531 2051
rect 1502 2024 1505 2036
rect 1495 1984 1499 1990
rect 1507 1984 1511 2024
rect 1527 1984 1531 2043
rect 1541 1984 1545 2066
rect 1561 2024 1565 2067
rect 1625 2024 1629 2081
rect 1654 2079 1658 2116
rect 1662 2112 1666 2116
rect 1662 2106 1681 2112
rect 1674 2093 1681 2106
rect 1723 2110 1727 2116
rect 1723 2098 1725 2110
rect 1654 2044 1660 2067
rect 1674 2044 1681 2081
rect 1645 2038 1660 2044
rect 1665 2038 1681 2044
rect 1745 2059 1749 2136
rect 1745 2047 1754 2059
rect 1791 2048 1795 2116
rect 1813 2087 1817 2136
rect 1823 2115 1827 2136
rect 1843 2124 1847 2136
rect 1851 2132 1855 2136
rect 1851 2128 1885 2132
rect 1843 2120 1873 2124
rect 1843 2119 1861 2120
rect 1823 2111 1847 2115
rect 1645 2024 1649 2038
rect 1665 2024 1669 2038
rect 1723 2030 1725 2042
rect 1723 2024 1727 2030
rect 1745 1984 1749 2047
rect 1791 2036 1793 2048
rect 1791 2024 1795 2036
rect 1813 2029 1817 2075
rect 1809 2023 1817 2029
rect 1809 1994 1813 2023
rect 1841 2016 1847 2111
rect 1809 1987 1817 1994
rect 1813 1964 1817 1987
rect 1821 1964 1825 2004
rect 1841 1984 1845 2016
rect 1881 2002 1885 2128
rect 1897 2022 1901 2136
rect 1919 2124 1923 2136
rect 1921 2112 1923 2124
rect 1929 2124 1933 2136
rect 1929 2112 1931 2124
rect 1849 1990 1873 1992
rect 1849 1988 1885 1990
rect 1849 1984 1853 1988
rect 1895 1984 1899 2010
rect 1913 2002 1917 2112
rect 1951 2104 1955 2136
rect 1922 2100 1955 2104
rect 1922 2036 1926 2100
rect 1942 2051 1946 2080
rect 1961 2078 1965 2136
rect 1981 2079 1985 2116
rect 2045 2079 2049 2136
rect 2113 2096 2117 2116
rect 2103 2089 2117 2096
rect 2123 2096 2127 2116
rect 2123 2089 2131 2096
rect 2045 2067 2054 2079
rect 2103 2073 2109 2089
rect 1942 2043 1951 2051
rect 1922 2024 1925 2036
rect 1915 1984 1919 1990
rect 1927 1984 1931 2024
rect 1947 1984 1951 2043
rect 1961 1984 1965 2066
rect 1981 2024 1985 2067
rect 2045 1984 2049 2067
rect 2106 2061 2109 2073
rect 2105 1984 2109 2061
rect 2125 2073 2131 2089
rect 2125 2061 2134 2073
rect 2125 1984 2129 2061
rect 2171 2059 2175 2136
rect 2193 2110 2197 2116
rect 2195 2098 2197 2110
rect 2253 2096 2257 2116
rect 2249 2089 2257 2096
rect 2263 2096 2267 2116
rect 2263 2089 2277 2096
rect 2249 2073 2255 2089
rect 2246 2061 2255 2073
rect 2166 2047 2175 2059
rect 2171 1984 2175 2047
rect 2195 2030 2197 2042
rect 2193 2024 2197 2030
rect 2251 1984 2255 2061
rect 2271 2073 2277 2089
rect 2271 2061 2274 2073
rect 2271 1984 2275 2061
rect 2345 2039 2349 2116
rect 2365 2093 2369 2116
rect 2385 2111 2389 2116
rect 2385 2104 2398 2111
rect 2365 2081 2374 2093
rect 2347 2027 2354 2039
rect 2350 1984 2354 2027
rect 2372 2024 2376 2081
rect 2394 2059 2398 2104
rect 2453 2096 2457 2116
rect 2443 2089 2457 2096
rect 2463 2096 2467 2116
rect 2533 2096 2537 2116
rect 2463 2089 2471 2096
rect 2443 2073 2449 2089
rect 2446 2061 2449 2073
rect 2394 2036 2398 2047
rect 2380 2028 2398 2036
rect 2380 2024 2384 2028
rect 2445 1984 2449 2061
rect 2465 2073 2471 2089
rect 2523 2089 2537 2096
rect 2543 2096 2547 2116
rect 2543 2089 2551 2096
rect 2523 2073 2529 2089
rect 2465 2061 2474 2073
rect 2526 2061 2529 2073
rect 2465 1984 2469 2061
rect 2525 1984 2529 2061
rect 2545 2073 2551 2089
rect 2545 2061 2554 2073
rect 2545 1984 2549 2061
rect 2605 2039 2609 2116
rect 2625 2093 2629 2116
rect 2645 2111 2649 2116
rect 2645 2104 2658 2111
rect 2625 2081 2634 2093
rect 2607 2027 2614 2039
rect 2610 1984 2614 2027
rect 2632 2024 2636 2081
rect 2654 2059 2658 2104
rect 2654 2036 2658 2047
rect 2705 2039 2709 2116
rect 2725 2093 2729 2116
rect 2745 2111 2749 2116
rect 2745 2104 2758 2111
rect 2725 2081 2734 2093
rect 2640 2028 2658 2036
rect 2640 2024 2644 2028
rect 2707 2027 2714 2039
rect 2710 1984 2714 2027
rect 2732 2024 2736 2081
rect 2754 2059 2758 2104
rect 2795 2079 2799 2116
rect 2815 2078 2819 2136
rect 2825 2104 2829 2136
rect 2847 2124 2851 2136
rect 2849 2112 2851 2124
rect 2857 2124 2861 2136
rect 2857 2112 2859 2124
rect 2825 2100 2858 2104
rect 2754 2036 2758 2047
rect 2740 2028 2758 2036
rect 2740 2024 2744 2028
rect 2795 2024 2799 2067
rect 2815 1984 2819 2066
rect 2834 2051 2838 2080
rect 2829 2043 2838 2051
rect 2829 1984 2833 2043
rect 2854 2036 2858 2100
rect 2855 2024 2858 2036
rect 2849 1984 2853 2024
rect 2863 2002 2867 2112
rect 2879 2022 2883 2136
rect 2925 2132 2929 2136
rect 2895 2128 2929 2132
rect 2861 1984 2865 1990
rect 2881 1984 2885 2010
rect 2895 2002 2899 2128
rect 2933 2124 2937 2136
rect 2907 2120 2937 2124
rect 2919 2119 2937 2120
rect 2953 2115 2957 2136
rect 2933 2111 2957 2115
rect 2933 2016 2939 2111
rect 2963 2087 2967 2136
rect 2963 2029 2967 2075
rect 2985 2048 2989 2116
rect 3031 2059 3035 2116
rect 3041 2073 3045 2116
rect 3061 2110 3065 2116
rect 3067 2098 3079 2110
rect 3041 2061 3054 2073
rect 2987 2036 2989 2048
rect 3026 2047 3035 2059
rect 2963 2023 2971 2029
rect 2985 2024 2989 2036
rect 2907 1990 2931 1992
rect 2895 1988 2931 1990
rect 2927 1984 2931 1988
rect 2935 1984 2939 2016
rect 2955 1964 2959 2004
rect 2967 1994 2971 2023
rect 2963 1987 2971 1994
rect 2963 1964 2967 1987
rect 3031 1984 3035 2047
rect 3053 1984 3057 2061
rect 3075 2024 3079 2098
rect 3145 2039 3149 2116
rect 3165 2093 3169 2116
rect 3185 2111 3189 2116
rect 3185 2104 3198 2111
rect 3165 2081 3174 2093
rect 3147 2027 3154 2039
rect 3150 1984 3154 2027
rect 3172 2024 3176 2081
rect 3194 2059 3198 2104
rect 3194 2036 3198 2047
rect 3245 2039 3249 2116
rect 3265 2093 3269 2116
rect 3285 2111 3289 2116
rect 3285 2104 3298 2111
rect 3265 2081 3274 2093
rect 3180 2028 3198 2036
rect 3180 2024 3184 2028
rect 3247 2027 3254 2039
rect 3250 1984 3254 2027
rect 3272 2024 3276 2081
rect 3294 2059 3298 2104
rect 3333 2096 3337 2116
rect 3329 2089 3337 2096
rect 3343 2096 3347 2116
rect 3343 2089 3357 2096
rect 3329 2073 3335 2089
rect 3326 2061 3335 2073
rect 3294 2036 3298 2047
rect 3280 2028 3298 2036
rect 3280 2024 3284 2028
rect 3331 1984 3335 2061
rect 3351 2073 3357 2089
rect 3351 2061 3354 2073
rect 3351 1984 3355 2061
rect 3425 2039 3429 2116
rect 3445 2093 3449 2116
rect 3465 2111 3469 2116
rect 3465 2104 3478 2111
rect 3445 2081 3454 2093
rect 3427 2027 3434 2039
rect 3430 1984 3434 2027
rect 3452 2024 3456 2081
rect 3474 2059 3478 2104
rect 3474 2036 3478 2047
rect 3512 2039 3516 2096
rect 3460 2028 3478 2036
rect 3460 2024 3464 2028
rect 3506 2027 3516 2039
rect 3500 1996 3506 2027
rect 3520 2019 3524 2096
rect 3528 2039 3532 2096
rect 3611 2079 3615 2136
rect 3773 2096 3777 2116
rect 3606 2067 3615 2079
rect 3528 2027 3535 2039
rect 3547 2027 3555 2039
rect 3520 2000 3526 2007
rect 3520 1996 3535 2000
rect 3500 1992 3515 1996
rect 3511 1984 3515 1992
rect 3531 1984 3535 1996
rect 3551 1984 3555 2027
rect 3611 1984 3615 2067
rect 3672 2039 3676 2096
rect 3666 2027 3676 2039
rect 3660 1996 3666 2027
rect 3680 2019 3684 2096
rect 3688 2039 3692 2096
rect 3769 2089 3777 2096
rect 3783 2096 3787 2116
rect 3783 2089 3797 2096
rect 3769 2073 3775 2089
rect 3766 2061 3775 2073
rect 3688 2027 3695 2039
rect 3707 2027 3715 2039
rect 3680 2000 3686 2007
rect 3680 1996 3695 2000
rect 3660 1992 3675 1996
rect 3671 1984 3675 1992
rect 3691 1984 3695 1996
rect 3711 1984 3715 2027
rect 3771 1984 3775 2061
rect 3791 2073 3797 2089
rect 3791 2061 3794 2073
rect 3791 1984 3795 2061
rect 3851 2059 3855 2136
rect 3873 2110 3877 2116
rect 3931 2111 3935 2116
rect 3875 2098 3877 2110
rect 3922 2104 3935 2111
rect 3922 2059 3926 2104
rect 3951 2093 3955 2116
rect 3946 2081 3955 2093
rect 3846 2047 3855 2059
rect 3851 1984 3855 2047
rect 3875 2030 3877 2042
rect 3873 2024 3877 2030
rect 3922 2036 3926 2047
rect 3922 2028 3940 2036
rect 3936 2024 3940 2028
rect 3944 2024 3948 2081
rect 3971 2039 3975 2116
rect 4053 2096 4057 2116
rect 4043 2089 4057 2096
rect 4063 2096 4067 2116
rect 4133 2096 4137 2116
rect 4063 2089 4071 2096
rect 4043 2073 4049 2089
rect 4046 2061 4049 2073
rect 3966 2027 3973 2039
rect 3966 1984 3970 2027
rect 4045 1984 4049 2061
rect 4065 2073 4071 2089
rect 4123 2089 4137 2096
rect 4143 2096 4147 2116
rect 4213 2096 4217 2116
rect 4143 2089 4151 2096
rect 4123 2073 4129 2089
rect 4065 2061 4074 2073
rect 4126 2061 4129 2073
rect 4065 1984 4069 2061
rect 4125 1984 4129 2061
rect 4145 2073 4151 2089
rect 4203 2089 4217 2096
rect 4223 2096 4227 2116
rect 4223 2089 4231 2096
rect 4203 2073 4209 2089
rect 4145 2061 4154 2073
rect 4206 2061 4209 2073
rect 4145 1984 4149 2061
rect 4205 1984 4209 2061
rect 4225 2073 4231 2089
rect 4225 2061 4234 2073
rect 4225 1984 4229 2061
rect 4271 2059 4275 2116
rect 4281 2073 4285 2116
rect 4301 2110 4305 2116
rect 4374 2112 4378 2116
rect 4307 2098 4319 2110
rect 4281 2061 4294 2073
rect 4266 2047 4275 2059
rect 4271 1984 4275 2047
rect 4293 1984 4297 2061
rect 4315 2024 4319 2098
rect 4359 2106 4378 2112
rect 4359 2093 4366 2106
rect 4359 2044 4366 2081
rect 4382 2079 4386 2116
rect 4404 2093 4408 2136
rect 4492 2093 4496 2136
rect 4406 2081 4415 2093
rect 4380 2044 4386 2067
rect 4359 2038 4375 2044
rect 4380 2038 4395 2044
rect 4371 2024 4375 2038
rect 4391 2024 4395 2038
rect 4411 2024 4415 2081
rect 4485 2081 4494 2093
rect 4485 2024 4489 2081
rect 4514 2079 4518 2116
rect 4522 2112 4526 2116
rect 4522 2106 4541 2112
rect 4534 2093 4541 2106
rect 4514 2044 4520 2067
rect 4534 2044 4541 2081
rect 4505 2038 4520 2044
rect 4525 2038 4541 2044
rect 4572 2039 4576 2096
rect 4505 2024 4509 2038
rect 4525 2024 4529 2038
rect 4566 2027 4576 2039
rect 4560 1996 4566 2027
rect 4580 2019 4584 2096
rect 4588 2039 4592 2096
rect 4672 2039 4676 2096
rect 4588 2027 4595 2039
rect 4607 2027 4615 2039
rect 4666 2027 4676 2039
rect 4580 2000 4586 2007
rect 4580 1996 4595 2000
rect 4560 1992 4575 1996
rect 4571 1984 4575 1992
rect 4591 1984 4595 1996
rect 4611 1984 4615 2027
rect 4660 1996 4666 2027
rect 4680 2019 4684 2096
rect 4688 2039 4692 2096
rect 4688 2027 4695 2039
rect 4707 2027 4715 2039
rect 4680 2000 4686 2007
rect 4680 1996 4695 2000
rect 4660 1992 4675 1996
rect 4671 1984 4675 1992
rect 4691 1984 4695 1996
rect 4711 1984 4715 2027
rect 31 1940 35 1944
rect 51 1940 55 1944
rect 71 1940 75 1944
rect 91 1940 95 1944
rect 111 1940 115 1944
rect 131 1940 135 1944
rect 151 1940 155 1944
rect 171 1940 175 1944
rect 245 1940 249 1944
rect 265 1940 269 1944
rect 330 1940 334 1944
rect 352 1940 356 1944
rect 360 1940 364 1944
rect 411 1940 415 1944
rect 431 1940 435 1944
rect 451 1940 455 1944
rect 471 1940 475 1944
rect 535 1940 539 1944
rect 555 1940 559 1944
rect 569 1940 573 1944
rect 589 1940 593 1944
rect 601 1940 605 1944
rect 621 1940 625 1944
rect 667 1940 671 1944
rect 675 1940 679 1944
rect 695 1940 699 1944
rect 703 1940 707 1944
rect 725 1940 729 1944
rect 785 1940 789 1944
rect 805 1940 809 1944
rect 875 1940 879 1944
rect 895 1940 899 1944
rect 905 1940 909 1944
rect 951 1940 955 1944
rect 971 1940 975 1944
rect 1031 1940 1035 1944
rect 1039 1940 1043 1944
rect 1116 1940 1120 1944
rect 1124 1940 1128 1944
rect 1146 1940 1150 1944
rect 1211 1940 1215 1944
rect 1231 1940 1235 1944
rect 1291 1940 1295 1944
rect 1299 1940 1303 1944
rect 1371 1940 1375 1944
rect 1393 1940 1397 1944
rect 1401 1940 1405 1944
rect 1421 1940 1425 1944
rect 1429 1940 1433 1944
rect 1475 1940 1479 1944
rect 1495 1940 1499 1944
rect 1507 1940 1511 1944
rect 1527 1940 1531 1944
rect 1541 1940 1545 1944
rect 1561 1940 1565 1944
rect 1625 1940 1629 1944
rect 1645 1940 1649 1944
rect 1665 1940 1669 1944
rect 1723 1940 1727 1944
rect 1745 1940 1749 1944
rect 1791 1940 1795 1944
rect 1813 1940 1817 1944
rect 1821 1940 1825 1944
rect 1841 1940 1845 1944
rect 1849 1940 1853 1944
rect 1895 1940 1899 1944
rect 1915 1940 1919 1944
rect 1927 1940 1931 1944
rect 1947 1940 1951 1944
rect 1961 1940 1965 1944
rect 1981 1940 1985 1944
rect 2045 1940 2049 1944
rect 2105 1940 2109 1944
rect 2125 1940 2129 1944
rect 2171 1940 2175 1944
rect 2193 1940 2197 1944
rect 2251 1940 2255 1944
rect 2271 1940 2275 1944
rect 2350 1940 2354 1944
rect 2372 1940 2376 1944
rect 2380 1940 2384 1944
rect 2445 1940 2449 1944
rect 2465 1940 2469 1944
rect 2525 1940 2529 1944
rect 2545 1940 2549 1944
rect 2610 1940 2614 1944
rect 2632 1940 2636 1944
rect 2640 1940 2644 1944
rect 2710 1940 2714 1944
rect 2732 1940 2736 1944
rect 2740 1940 2744 1944
rect 2795 1940 2799 1944
rect 2815 1940 2819 1944
rect 2829 1940 2833 1944
rect 2849 1940 2853 1944
rect 2861 1940 2865 1944
rect 2881 1940 2885 1944
rect 2927 1940 2931 1944
rect 2935 1940 2939 1944
rect 2955 1940 2959 1944
rect 2963 1940 2967 1944
rect 2985 1940 2989 1944
rect 3031 1940 3035 1944
rect 3053 1940 3057 1944
rect 3075 1940 3079 1944
rect 3150 1940 3154 1944
rect 3172 1940 3176 1944
rect 3180 1940 3184 1944
rect 3250 1940 3254 1944
rect 3272 1940 3276 1944
rect 3280 1940 3284 1944
rect 3331 1940 3335 1944
rect 3351 1940 3355 1944
rect 3430 1940 3434 1944
rect 3452 1940 3456 1944
rect 3460 1940 3464 1944
rect 3511 1940 3515 1944
rect 3531 1940 3535 1944
rect 3551 1940 3555 1944
rect 3611 1940 3615 1944
rect 3671 1940 3675 1944
rect 3691 1940 3695 1944
rect 3711 1940 3715 1944
rect 3771 1940 3775 1944
rect 3791 1940 3795 1944
rect 3851 1940 3855 1944
rect 3873 1940 3877 1944
rect 3936 1940 3940 1944
rect 3944 1940 3948 1944
rect 3966 1940 3970 1944
rect 4045 1940 4049 1944
rect 4065 1940 4069 1944
rect 4125 1940 4129 1944
rect 4145 1940 4149 1944
rect 4205 1940 4209 1944
rect 4225 1940 4229 1944
rect 4271 1940 4275 1944
rect 4293 1940 4297 1944
rect 4315 1940 4319 1944
rect 4371 1940 4375 1944
rect 4391 1940 4395 1944
rect 4411 1940 4415 1944
rect 4485 1940 4489 1944
rect 4505 1940 4509 1944
rect 4525 1940 4529 1944
rect 4571 1940 4575 1944
rect 4591 1940 4595 1944
rect 4611 1940 4615 1944
rect 4671 1940 4675 1944
rect 4691 1940 4695 1944
rect 4711 1940 4715 1944
rect 35 1916 39 1920
rect 55 1916 59 1920
rect 69 1916 73 1920
rect 89 1916 93 1920
rect 101 1916 105 1920
rect 121 1916 125 1920
rect 167 1916 171 1920
rect 175 1916 179 1920
rect 195 1916 199 1920
rect 203 1916 207 1920
rect 225 1916 229 1920
rect 276 1916 280 1920
rect 284 1916 288 1920
rect 306 1916 310 1920
rect 390 1916 394 1920
rect 412 1916 416 1920
rect 420 1916 424 1920
rect 490 1916 494 1920
rect 512 1916 516 1920
rect 520 1916 524 1920
rect 590 1916 594 1920
rect 612 1916 616 1920
rect 620 1916 624 1920
rect 671 1916 675 1920
rect 731 1916 735 1920
rect 817 1916 821 1920
rect 825 1916 829 1920
rect 871 1916 875 1920
rect 891 1916 895 1920
rect 911 1916 915 1920
rect 975 1916 979 1920
rect 995 1916 999 1920
rect 1009 1916 1013 1920
rect 1029 1916 1033 1920
rect 1041 1916 1045 1920
rect 1061 1916 1065 1920
rect 1107 1916 1111 1920
rect 1115 1916 1119 1920
rect 1135 1916 1139 1920
rect 1143 1916 1147 1920
rect 1165 1916 1169 1920
rect 1211 1916 1215 1920
rect 1231 1916 1235 1920
rect 1310 1916 1314 1920
rect 1332 1916 1336 1920
rect 1340 1916 1344 1920
rect 1405 1916 1409 1920
rect 1425 1916 1429 1920
rect 1445 1916 1449 1920
rect 1465 1916 1469 1920
rect 1485 1916 1489 1920
rect 1505 1916 1509 1920
rect 1525 1916 1529 1920
rect 1545 1916 1549 1920
rect 1595 1916 1599 1920
rect 1615 1916 1619 1920
rect 1629 1916 1633 1920
rect 1649 1916 1653 1920
rect 1661 1916 1665 1920
rect 1681 1916 1685 1920
rect 1727 1916 1731 1920
rect 1735 1916 1739 1920
rect 1755 1916 1759 1920
rect 1763 1916 1767 1920
rect 1785 1916 1789 1920
rect 1845 1916 1849 1920
rect 1865 1916 1869 1920
rect 1885 1916 1889 1920
rect 1931 1916 1935 1920
rect 1939 1916 1943 1920
rect 2025 1916 2029 1920
rect 2045 1916 2049 1920
rect 2065 1916 2069 1920
rect 2137 1916 2141 1920
rect 2145 1916 2149 1920
rect 2191 1916 2195 1920
rect 2211 1916 2215 1920
rect 2231 1916 2235 1920
rect 2291 1916 2295 1920
rect 2313 1916 2317 1920
rect 2321 1916 2325 1920
rect 2341 1916 2345 1920
rect 2349 1916 2353 1920
rect 2395 1916 2399 1920
rect 2415 1916 2419 1920
rect 2427 1916 2431 1920
rect 2447 1916 2451 1920
rect 2461 1916 2465 1920
rect 2481 1916 2485 1920
rect 2535 1916 2539 1920
rect 2555 1916 2559 1920
rect 2569 1916 2573 1920
rect 2589 1916 2593 1920
rect 2601 1916 2605 1920
rect 2621 1916 2625 1920
rect 2667 1916 2671 1920
rect 2675 1916 2679 1920
rect 2695 1916 2699 1920
rect 2703 1916 2707 1920
rect 2725 1916 2729 1920
rect 2775 1916 2779 1920
rect 2795 1916 2799 1920
rect 2809 1916 2813 1920
rect 2829 1916 2833 1920
rect 2841 1916 2845 1920
rect 2861 1916 2865 1920
rect 2907 1916 2911 1920
rect 2915 1916 2919 1920
rect 2935 1916 2939 1920
rect 2943 1916 2947 1920
rect 2965 1916 2969 1920
rect 3025 1916 3029 1920
rect 3085 1916 3089 1920
rect 3105 1916 3109 1920
rect 3165 1916 3169 1920
rect 3211 1916 3215 1920
rect 3231 1916 3235 1920
rect 3251 1916 3255 1920
rect 3311 1916 3315 1920
rect 3319 1916 3323 1920
rect 3401 1916 3405 1920
rect 3423 1916 3427 1920
rect 3445 1916 3449 1920
rect 3491 1916 3495 1920
rect 3565 1916 3569 1920
rect 3585 1916 3589 1920
rect 3605 1916 3609 1920
rect 3625 1916 3629 1920
rect 3685 1916 3689 1920
rect 3757 1916 3761 1920
rect 3765 1916 3769 1920
rect 3811 1916 3815 1920
rect 3833 1916 3837 1920
rect 3891 1916 3895 1920
rect 3913 1916 3917 1920
rect 3935 1916 3939 1920
rect 4005 1916 4009 1920
rect 4025 1916 4029 1920
rect 4045 1916 4049 1920
rect 4065 1916 4069 1920
rect 4111 1916 4115 1920
rect 4131 1916 4135 1920
rect 4151 1916 4155 1920
rect 4171 1916 4175 1920
rect 4231 1916 4235 1920
rect 4251 1916 4255 1920
rect 4311 1916 4315 1920
rect 4333 1916 4337 1920
rect 4355 1916 4359 1920
rect 4411 1916 4415 1920
rect 4431 1916 4435 1920
rect 4451 1916 4455 1920
rect 4471 1916 4475 1920
rect 4545 1916 4549 1920
rect 4596 1916 4600 1920
rect 4604 1916 4608 1920
rect 4626 1916 4630 1920
rect 4691 1916 4695 1920
rect 35 1793 39 1836
rect 55 1794 59 1876
rect 69 1817 73 1876
rect 89 1836 93 1876
rect 101 1870 105 1876
rect 95 1824 98 1836
rect 69 1809 78 1817
rect 35 1744 39 1781
rect 55 1724 59 1782
rect 74 1780 78 1809
rect 94 1760 98 1824
rect 65 1756 98 1760
rect 65 1724 69 1756
rect 103 1748 107 1858
rect 121 1850 125 1876
rect 167 1872 171 1876
rect 135 1870 171 1872
rect 147 1868 171 1870
rect 89 1736 91 1748
rect 87 1724 91 1736
rect 97 1736 99 1748
rect 97 1724 101 1736
rect 119 1724 123 1838
rect 135 1732 139 1858
rect 175 1844 179 1876
rect 195 1856 199 1896
rect 203 1873 207 1896
rect 203 1866 211 1873
rect 173 1749 179 1844
rect 207 1837 211 1866
rect 203 1831 211 1837
rect 203 1785 207 1831
rect 225 1824 229 1836
rect 276 1832 280 1836
rect 227 1812 229 1824
rect 262 1824 280 1832
rect 262 1813 266 1824
rect 173 1745 197 1749
rect 159 1740 177 1741
rect 147 1736 177 1740
rect 135 1728 169 1732
rect 165 1724 169 1728
rect 173 1724 177 1736
rect 193 1724 197 1745
rect 203 1724 207 1773
rect 225 1744 229 1812
rect 262 1756 266 1801
rect 284 1779 288 1836
rect 306 1833 310 1876
rect 390 1833 394 1876
rect 306 1821 313 1833
rect 387 1821 394 1833
rect 286 1767 295 1779
rect 262 1749 275 1756
rect 271 1744 275 1749
rect 291 1744 295 1767
rect 311 1744 315 1821
rect 385 1744 389 1821
rect 412 1779 416 1836
rect 420 1832 424 1836
rect 490 1833 494 1876
rect 420 1824 438 1832
rect 434 1813 438 1824
rect 487 1821 494 1833
rect 405 1767 414 1779
rect 405 1744 409 1767
rect 434 1756 438 1801
rect 425 1749 438 1756
rect 425 1744 429 1749
rect 485 1744 489 1821
rect 512 1779 516 1836
rect 520 1832 524 1836
rect 590 1833 594 1876
rect 520 1824 538 1832
rect 534 1813 538 1824
rect 587 1821 594 1833
rect 505 1767 514 1779
rect 505 1744 509 1767
rect 534 1756 538 1801
rect 525 1749 538 1756
rect 525 1744 529 1749
rect 585 1744 589 1821
rect 612 1779 616 1836
rect 620 1832 624 1836
rect 620 1824 638 1832
rect 634 1813 638 1824
rect 605 1767 614 1779
rect 605 1744 609 1767
rect 634 1756 638 1801
rect 671 1793 675 1876
rect 731 1793 735 1876
rect 871 1868 875 1876
rect 860 1864 875 1868
rect 891 1864 895 1876
rect 817 1813 821 1836
rect 806 1801 821 1813
rect 825 1813 829 1836
rect 860 1833 866 1864
rect 880 1860 895 1864
rect 880 1853 886 1860
rect 866 1821 876 1833
rect 825 1801 834 1813
rect 666 1781 675 1793
rect 726 1781 735 1793
rect 625 1749 638 1756
rect 625 1744 629 1749
rect 671 1724 675 1781
rect 731 1724 735 1781
rect 805 1724 809 1801
rect 825 1724 829 1801
rect 872 1764 876 1821
rect 880 1764 884 1841
rect 911 1833 915 1876
rect 888 1821 895 1833
rect 907 1821 915 1833
rect 888 1764 892 1821
rect 975 1793 979 1836
rect 995 1794 999 1876
rect 1009 1817 1013 1876
rect 1029 1836 1033 1876
rect 1041 1870 1045 1876
rect 1035 1824 1038 1836
rect 1009 1809 1018 1817
rect 975 1744 979 1781
rect 995 1724 999 1782
rect 1014 1780 1018 1809
rect 1034 1760 1038 1824
rect 1005 1756 1038 1760
rect 1005 1724 1009 1756
rect 1043 1748 1047 1858
rect 1061 1850 1065 1876
rect 1107 1872 1111 1876
rect 1075 1870 1111 1872
rect 1087 1868 1111 1870
rect 1029 1736 1031 1748
rect 1027 1724 1031 1736
rect 1037 1736 1039 1748
rect 1037 1724 1041 1736
rect 1059 1724 1063 1838
rect 1075 1732 1079 1858
rect 1115 1844 1119 1876
rect 1135 1856 1139 1896
rect 1143 1873 1147 1896
rect 1143 1866 1151 1873
rect 1113 1749 1119 1844
rect 1147 1837 1151 1866
rect 1143 1831 1151 1837
rect 1143 1785 1147 1831
rect 1165 1824 1169 1836
rect 1167 1812 1169 1824
rect 1113 1745 1137 1749
rect 1099 1740 1117 1741
rect 1087 1736 1117 1740
rect 1075 1728 1109 1732
rect 1105 1724 1109 1728
rect 1113 1724 1117 1736
rect 1133 1724 1137 1745
rect 1143 1724 1147 1773
rect 1165 1744 1169 1812
rect 1211 1799 1215 1876
rect 1206 1787 1215 1799
rect 1209 1771 1215 1787
rect 1231 1799 1235 1876
rect 1310 1833 1314 1876
rect 1307 1821 1314 1833
rect 1231 1787 1234 1799
rect 1231 1771 1237 1787
rect 1209 1764 1217 1771
rect 1213 1744 1217 1764
rect 1223 1764 1237 1771
rect 1223 1744 1227 1764
rect 1305 1744 1309 1821
rect 1332 1779 1336 1836
rect 1340 1832 1344 1836
rect 1340 1824 1358 1832
rect 1354 1813 1358 1824
rect 1325 1767 1334 1779
rect 1325 1744 1329 1767
rect 1354 1756 1358 1801
rect 1345 1749 1358 1756
rect 1405 1776 1409 1836
rect 1425 1776 1429 1836
rect 1445 1776 1449 1836
rect 1465 1776 1469 1836
rect 1485 1776 1489 1836
rect 1505 1776 1509 1836
rect 1525 1779 1529 1836
rect 1545 1779 1549 1836
rect 1595 1793 1599 1836
rect 1615 1794 1619 1876
rect 1629 1817 1633 1876
rect 1649 1836 1653 1876
rect 1661 1870 1665 1876
rect 1655 1824 1658 1836
rect 1629 1809 1638 1817
rect 1405 1764 1418 1776
rect 1445 1764 1458 1776
rect 1485 1764 1498 1776
rect 1525 1767 1534 1779
rect 1546 1767 1549 1779
rect 1345 1744 1349 1749
rect 1405 1744 1409 1764
rect 1425 1744 1429 1764
rect 1445 1744 1449 1764
rect 1465 1744 1469 1764
rect 1485 1744 1489 1764
rect 1505 1744 1509 1764
rect 1525 1744 1529 1767
rect 1545 1744 1549 1767
rect 1595 1744 1599 1781
rect 1615 1724 1619 1782
rect 1634 1780 1638 1809
rect 1654 1760 1658 1824
rect 1625 1756 1658 1760
rect 1625 1724 1629 1756
rect 1663 1748 1667 1858
rect 1681 1850 1685 1876
rect 1727 1872 1731 1876
rect 1695 1870 1731 1872
rect 1707 1868 1731 1870
rect 1649 1736 1651 1748
rect 1647 1724 1651 1736
rect 1657 1736 1659 1748
rect 1657 1724 1661 1736
rect 1679 1724 1683 1838
rect 1695 1732 1699 1858
rect 1735 1844 1739 1876
rect 1755 1856 1759 1896
rect 1763 1873 1767 1896
rect 1763 1866 1771 1873
rect 1733 1749 1739 1844
rect 1767 1837 1771 1866
rect 1763 1831 1771 1837
rect 2313 1873 2317 1896
rect 2309 1866 2317 1873
rect 2309 1837 2313 1866
rect 2321 1856 2325 1896
rect 2341 1844 2345 1876
rect 2349 1872 2353 1876
rect 2349 1870 2385 1872
rect 2349 1868 2373 1870
rect 1763 1785 1767 1831
rect 1785 1824 1789 1836
rect 1787 1812 1789 1824
rect 1733 1745 1757 1749
rect 1719 1740 1737 1741
rect 1707 1736 1737 1740
rect 1695 1728 1729 1732
rect 1725 1724 1729 1728
rect 1733 1724 1737 1736
rect 1753 1724 1757 1745
rect 1763 1724 1767 1773
rect 1785 1744 1789 1812
rect 1845 1779 1849 1836
rect 1865 1822 1869 1836
rect 1885 1822 1889 1836
rect 1865 1816 1880 1822
rect 1885 1816 1901 1822
rect 1874 1793 1880 1816
rect 1845 1767 1854 1779
rect 1852 1724 1856 1767
rect 1874 1744 1878 1781
rect 1894 1779 1901 1816
rect 1931 1813 1935 1836
rect 1926 1801 1935 1813
rect 1939 1813 1943 1836
rect 1939 1801 1954 1813
rect 1894 1754 1901 1767
rect 1882 1748 1901 1754
rect 1882 1744 1886 1748
rect 1931 1724 1935 1801
rect 1951 1724 1955 1801
rect 2025 1779 2029 1836
rect 2045 1822 2049 1836
rect 2065 1822 2069 1836
rect 2045 1816 2060 1822
rect 2065 1816 2081 1822
rect 2054 1793 2060 1816
rect 2025 1767 2034 1779
rect 2032 1724 2036 1767
rect 2054 1744 2058 1781
rect 2074 1779 2081 1816
rect 2137 1813 2141 1836
rect 2126 1801 2141 1813
rect 2145 1813 2149 1836
rect 2191 1822 2195 1836
rect 2211 1822 2215 1836
rect 2179 1816 2195 1822
rect 2200 1816 2215 1822
rect 2145 1801 2154 1813
rect 2074 1754 2081 1767
rect 2062 1748 2081 1754
rect 2062 1744 2066 1748
rect 2125 1724 2129 1801
rect 2145 1724 2149 1801
rect 2179 1779 2186 1816
rect 2200 1793 2206 1816
rect 2179 1754 2186 1767
rect 2179 1748 2198 1754
rect 2194 1744 2198 1748
rect 2202 1744 2206 1781
rect 2231 1779 2235 1836
rect 2226 1767 2235 1779
rect 2291 1824 2295 1836
rect 2309 1831 2317 1837
rect 2291 1812 2293 1824
rect 2224 1724 2228 1767
rect 2291 1744 2295 1812
rect 2313 1785 2317 1831
rect 2313 1724 2317 1773
rect 2341 1749 2347 1844
rect 2323 1745 2347 1749
rect 2323 1724 2327 1745
rect 2343 1740 2361 1741
rect 2343 1736 2373 1740
rect 2343 1724 2347 1736
rect 2381 1732 2385 1858
rect 2395 1850 2399 1876
rect 2415 1870 2419 1876
rect 2351 1728 2385 1732
rect 2351 1724 2355 1728
rect 2397 1724 2401 1838
rect 2413 1748 2417 1858
rect 2427 1836 2431 1876
rect 2422 1824 2425 1836
rect 2422 1760 2426 1824
rect 2447 1817 2451 1876
rect 2442 1809 2451 1817
rect 2442 1780 2446 1809
rect 2461 1794 2465 1876
rect 2481 1793 2485 1836
rect 2535 1793 2539 1836
rect 2555 1794 2559 1876
rect 2569 1817 2573 1876
rect 2589 1836 2593 1876
rect 2601 1870 2605 1876
rect 2595 1824 2598 1836
rect 2569 1809 2578 1817
rect 2422 1756 2455 1760
rect 2421 1736 2423 1748
rect 2419 1724 2423 1736
rect 2429 1736 2431 1748
rect 2429 1724 2433 1736
rect 2451 1724 2455 1756
rect 2461 1724 2465 1782
rect 2481 1744 2485 1781
rect 2535 1744 2539 1781
rect 2555 1724 2559 1782
rect 2574 1780 2578 1809
rect 2594 1760 2598 1824
rect 2565 1756 2598 1760
rect 2565 1724 2569 1756
rect 2603 1748 2607 1858
rect 2621 1850 2625 1876
rect 2667 1872 2671 1876
rect 2635 1870 2671 1872
rect 2647 1868 2671 1870
rect 2589 1736 2591 1748
rect 2587 1724 2591 1736
rect 2597 1736 2599 1748
rect 2597 1724 2601 1736
rect 2619 1724 2623 1838
rect 2635 1732 2639 1858
rect 2675 1844 2679 1876
rect 2695 1856 2699 1896
rect 2703 1873 2707 1896
rect 2703 1866 2711 1873
rect 2673 1749 2679 1844
rect 2707 1837 2711 1866
rect 2703 1831 2711 1837
rect 2703 1785 2707 1831
rect 2725 1824 2729 1836
rect 2727 1812 2729 1824
rect 2673 1745 2697 1749
rect 2659 1740 2677 1741
rect 2647 1736 2677 1740
rect 2635 1728 2669 1732
rect 2665 1724 2669 1728
rect 2673 1724 2677 1736
rect 2693 1724 2697 1745
rect 2703 1724 2707 1773
rect 2725 1744 2729 1812
rect 2775 1793 2779 1836
rect 2795 1794 2799 1876
rect 2809 1817 2813 1876
rect 2829 1836 2833 1876
rect 2841 1870 2845 1876
rect 2835 1824 2838 1836
rect 2809 1809 2818 1817
rect 2775 1744 2779 1781
rect 2795 1724 2799 1782
rect 2814 1780 2818 1809
rect 2834 1760 2838 1824
rect 2805 1756 2838 1760
rect 2805 1724 2809 1756
rect 2843 1748 2847 1858
rect 2861 1850 2865 1876
rect 2907 1872 2911 1876
rect 2875 1870 2911 1872
rect 2887 1868 2911 1870
rect 2829 1736 2831 1748
rect 2827 1724 2831 1736
rect 2837 1736 2839 1748
rect 2837 1724 2841 1736
rect 2859 1724 2863 1838
rect 2875 1732 2879 1858
rect 2915 1844 2919 1876
rect 2935 1856 2939 1896
rect 2943 1873 2947 1896
rect 2943 1866 2951 1873
rect 2913 1749 2919 1844
rect 2947 1837 2951 1866
rect 2943 1831 2951 1837
rect 2943 1785 2947 1831
rect 2965 1824 2969 1836
rect 2967 1812 2969 1824
rect 2913 1745 2937 1749
rect 2899 1740 2917 1741
rect 2887 1736 2917 1740
rect 2875 1728 2909 1732
rect 2905 1724 2909 1728
rect 2913 1724 2917 1736
rect 2933 1724 2937 1745
rect 2943 1724 2947 1773
rect 2965 1744 2969 1812
rect 3025 1779 3029 1836
rect 3085 1799 3089 1876
rect 3086 1787 3089 1799
rect 3025 1767 3034 1779
rect 3083 1771 3089 1787
rect 3105 1799 3109 1876
rect 3105 1787 3114 1799
rect 3105 1771 3111 1787
rect 3025 1744 3029 1767
rect 3083 1764 3097 1771
rect 3093 1744 3097 1764
rect 3103 1764 3111 1771
rect 3165 1779 3169 1836
rect 3211 1822 3215 1836
rect 3231 1822 3235 1836
rect 3199 1816 3215 1822
rect 3220 1816 3235 1822
rect 3199 1779 3206 1816
rect 3220 1793 3226 1816
rect 3165 1767 3174 1779
rect 3103 1744 3107 1764
rect 3165 1744 3169 1767
rect 3199 1754 3206 1767
rect 3199 1748 3218 1754
rect 3214 1744 3218 1748
rect 3222 1744 3226 1781
rect 3251 1779 3255 1836
rect 3311 1813 3315 1836
rect 3306 1801 3315 1813
rect 3319 1813 3323 1836
rect 3319 1801 3334 1813
rect 3246 1767 3255 1779
rect 3244 1724 3248 1767
rect 3311 1724 3315 1801
rect 3331 1724 3335 1801
rect 3401 1762 3405 1836
rect 3423 1799 3427 1876
rect 3445 1813 3449 1876
rect 3445 1801 3454 1813
rect 3426 1787 3439 1799
rect 3401 1750 3413 1762
rect 3415 1744 3419 1750
rect 3435 1744 3439 1787
rect 3445 1744 3449 1801
rect 3491 1779 3495 1836
rect 3565 1813 3569 1836
rect 3566 1801 3569 1813
rect 3486 1767 3495 1779
rect 3491 1744 3495 1767
rect 3560 1753 3566 1801
rect 3585 1779 3589 1836
rect 3605 1814 3609 1836
rect 3625 1814 3629 1836
rect 3605 1808 3618 1814
rect 3625 1813 3645 1814
rect 3625 1808 3633 1813
rect 3614 1779 3618 1808
rect 3587 1767 3589 1779
rect 3585 1765 3589 1767
rect 3585 1758 3598 1765
rect 3560 1749 3590 1753
rect 3586 1744 3590 1749
rect 3594 1744 3598 1758
rect 3614 1744 3618 1767
rect 3633 1759 3639 1801
rect 3622 1752 3639 1759
rect 3685 1779 3689 1836
rect 3757 1813 3761 1836
rect 3746 1801 3761 1813
rect 3765 1813 3769 1836
rect 3811 1813 3815 1876
rect 3833 1830 3837 1836
rect 3835 1818 3837 1830
rect 3891 1813 3895 1876
rect 3765 1801 3774 1813
rect 3806 1801 3815 1813
rect 3886 1801 3895 1813
rect 3685 1767 3694 1779
rect 3622 1744 3626 1752
rect 3685 1744 3689 1767
rect 3745 1724 3749 1801
rect 3765 1724 3769 1801
rect 3811 1724 3815 1801
rect 3835 1750 3837 1762
rect 3833 1744 3837 1750
rect 3891 1744 3895 1801
rect 3913 1799 3917 1876
rect 3901 1787 3914 1799
rect 3901 1744 3905 1787
rect 3935 1762 3939 1836
rect 4005 1813 4009 1836
rect 4006 1801 4009 1813
rect 3927 1750 3939 1762
rect 4000 1753 4006 1801
rect 4025 1779 4029 1836
rect 4045 1814 4049 1836
rect 4065 1814 4069 1836
rect 4111 1814 4115 1836
rect 4131 1814 4135 1836
rect 4045 1808 4058 1814
rect 4065 1813 4085 1814
rect 4065 1808 4073 1813
rect 4054 1779 4058 1808
rect 4095 1813 4115 1814
rect 4107 1808 4115 1813
rect 4122 1808 4135 1814
rect 4027 1767 4029 1779
rect 4025 1765 4029 1767
rect 4025 1758 4038 1765
rect 3921 1744 3925 1750
rect 4000 1749 4030 1753
rect 4026 1744 4030 1749
rect 4034 1744 4038 1758
rect 4054 1744 4058 1767
rect 4073 1759 4079 1801
rect 4062 1752 4079 1759
rect 4101 1759 4107 1801
rect 4122 1779 4126 1808
rect 4151 1779 4155 1836
rect 4171 1813 4175 1836
rect 4171 1801 4174 1813
rect 4151 1767 4153 1779
rect 4101 1752 4118 1759
rect 4062 1744 4066 1752
rect 4114 1744 4118 1752
rect 4122 1744 4126 1767
rect 4151 1765 4155 1767
rect 4142 1758 4155 1765
rect 4142 1744 4146 1758
rect 4174 1753 4180 1801
rect 4231 1799 4235 1876
rect 4226 1787 4235 1799
rect 4229 1771 4235 1787
rect 4251 1799 4255 1876
rect 4311 1813 4315 1876
rect 4306 1801 4315 1813
rect 4251 1787 4254 1799
rect 4251 1771 4257 1787
rect 4229 1764 4237 1771
rect 4150 1749 4180 1753
rect 4150 1744 4154 1749
rect 4233 1744 4237 1764
rect 4243 1764 4257 1771
rect 4243 1744 4247 1764
rect 4311 1744 4315 1801
rect 4333 1799 4337 1876
rect 4321 1787 4334 1799
rect 4321 1744 4325 1787
rect 4355 1762 4359 1836
rect 4411 1814 4415 1836
rect 4431 1814 4435 1836
rect 4395 1813 4415 1814
rect 4407 1808 4415 1813
rect 4422 1808 4435 1814
rect 4347 1750 4359 1762
rect 4401 1759 4407 1801
rect 4422 1779 4426 1808
rect 4451 1779 4455 1836
rect 4471 1813 4475 1836
rect 4471 1801 4474 1813
rect 4451 1767 4453 1779
rect 4401 1752 4418 1759
rect 4341 1744 4345 1750
rect 4414 1744 4418 1752
rect 4422 1744 4426 1767
rect 4451 1765 4455 1767
rect 4442 1758 4455 1765
rect 4442 1744 4446 1758
rect 4474 1753 4480 1801
rect 4450 1749 4480 1753
rect 4545 1793 4549 1876
rect 4596 1832 4600 1836
rect 4582 1824 4600 1832
rect 4582 1813 4586 1824
rect 4545 1781 4554 1793
rect 4450 1744 4454 1749
rect 4545 1724 4549 1781
rect 4582 1756 4586 1801
rect 4604 1779 4608 1836
rect 4626 1833 4630 1876
rect 4626 1821 4633 1833
rect 4606 1767 4615 1779
rect 4582 1749 4595 1756
rect 4591 1744 4595 1749
rect 4611 1744 4615 1767
rect 4631 1744 4635 1821
rect 4691 1793 4695 1876
rect 4686 1781 4695 1793
rect 4691 1724 4695 1781
rect 35 1700 39 1704
rect 55 1700 59 1704
rect 65 1700 69 1704
rect 87 1700 91 1704
rect 97 1700 101 1704
rect 119 1700 123 1704
rect 165 1700 169 1704
rect 173 1700 177 1704
rect 193 1700 197 1704
rect 203 1700 207 1704
rect 225 1700 229 1704
rect 271 1700 275 1704
rect 291 1700 295 1704
rect 311 1700 315 1704
rect 385 1700 389 1704
rect 405 1700 409 1704
rect 425 1700 429 1704
rect 485 1700 489 1704
rect 505 1700 509 1704
rect 525 1700 529 1704
rect 585 1700 589 1704
rect 605 1700 609 1704
rect 625 1700 629 1704
rect 671 1700 675 1704
rect 731 1700 735 1704
rect 805 1700 809 1704
rect 825 1700 829 1704
rect 872 1700 876 1704
rect 880 1700 884 1704
rect 888 1700 892 1704
rect 975 1700 979 1704
rect 995 1700 999 1704
rect 1005 1700 1009 1704
rect 1027 1700 1031 1704
rect 1037 1700 1041 1704
rect 1059 1700 1063 1704
rect 1105 1700 1109 1704
rect 1113 1700 1117 1704
rect 1133 1700 1137 1704
rect 1143 1700 1147 1704
rect 1165 1700 1169 1704
rect 1213 1700 1217 1704
rect 1223 1700 1227 1704
rect 1305 1700 1309 1704
rect 1325 1700 1329 1704
rect 1345 1700 1349 1704
rect 1405 1700 1409 1704
rect 1425 1700 1429 1704
rect 1445 1700 1449 1704
rect 1465 1700 1469 1704
rect 1485 1700 1489 1704
rect 1505 1700 1509 1704
rect 1525 1700 1529 1704
rect 1545 1700 1549 1704
rect 1595 1700 1599 1704
rect 1615 1700 1619 1704
rect 1625 1700 1629 1704
rect 1647 1700 1651 1704
rect 1657 1700 1661 1704
rect 1679 1700 1683 1704
rect 1725 1700 1729 1704
rect 1733 1700 1737 1704
rect 1753 1700 1757 1704
rect 1763 1700 1767 1704
rect 1785 1700 1789 1704
rect 1852 1700 1856 1704
rect 1874 1700 1878 1704
rect 1882 1700 1886 1704
rect 1931 1700 1935 1704
rect 1951 1700 1955 1704
rect 2032 1700 2036 1704
rect 2054 1700 2058 1704
rect 2062 1700 2066 1704
rect 2125 1700 2129 1704
rect 2145 1700 2149 1704
rect 2194 1700 2198 1704
rect 2202 1700 2206 1704
rect 2224 1700 2228 1704
rect 2291 1700 2295 1704
rect 2313 1700 2317 1704
rect 2323 1700 2327 1704
rect 2343 1700 2347 1704
rect 2351 1700 2355 1704
rect 2397 1700 2401 1704
rect 2419 1700 2423 1704
rect 2429 1700 2433 1704
rect 2451 1700 2455 1704
rect 2461 1700 2465 1704
rect 2481 1700 2485 1704
rect 2535 1700 2539 1704
rect 2555 1700 2559 1704
rect 2565 1700 2569 1704
rect 2587 1700 2591 1704
rect 2597 1700 2601 1704
rect 2619 1700 2623 1704
rect 2665 1700 2669 1704
rect 2673 1700 2677 1704
rect 2693 1700 2697 1704
rect 2703 1700 2707 1704
rect 2725 1700 2729 1704
rect 2775 1700 2779 1704
rect 2795 1700 2799 1704
rect 2805 1700 2809 1704
rect 2827 1700 2831 1704
rect 2837 1700 2841 1704
rect 2859 1700 2863 1704
rect 2905 1700 2909 1704
rect 2913 1700 2917 1704
rect 2933 1700 2937 1704
rect 2943 1700 2947 1704
rect 2965 1700 2969 1704
rect 3025 1700 3029 1704
rect 3093 1700 3097 1704
rect 3103 1700 3107 1704
rect 3165 1700 3169 1704
rect 3214 1700 3218 1704
rect 3222 1700 3226 1704
rect 3244 1700 3248 1704
rect 3311 1700 3315 1704
rect 3331 1700 3335 1704
rect 3415 1700 3419 1704
rect 3435 1700 3439 1704
rect 3445 1700 3449 1704
rect 3491 1700 3495 1704
rect 3586 1700 3590 1704
rect 3594 1700 3598 1704
rect 3614 1700 3618 1704
rect 3622 1700 3626 1704
rect 3685 1700 3689 1704
rect 3745 1700 3749 1704
rect 3765 1700 3769 1704
rect 3811 1700 3815 1704
rect 3833 1700 3837 1704
rect 3891 1700 3895 1704
rect 3901 1700 3905 1704
rect 3921 1700 3925 1704
rect 4026 1700 4030 1704
rect 4034 1700 4038 1704
rect 4054 1700 4058 1704
rect 4062 1700 4066 1704
rect 4114 1700 4118 1704
rect 4122 1700 4126 1704
rect 4142 1700 4146 1704
rect 4150 1700 4154 1704
rect 4233 1700 4237 1704
rect 4243 1700 4247 1704
rect 4311 1700 4315 1704
rect 4321 1700 4325 1704
rect 4341 1700 4345 1704
rect 4414 1700 4418 1704
rect 4422 1700 4426 1704
rect 4442 1700 4446 1704
rect 4450 1700 4454 1704
rect 4545 1700 4549 1704
rect 4591 1700 4595 1704
rect 4611 1700 4615 1704
rect 4631 1700 4635 1704
rect 4691 1700 4695 1704
rect 31 1676 35 1680
rect 51 1676 55 1680
rect 71 1676 75 1680
rect 91 1676 95 1680
rect 111 1676 115 1680
rect 131 1676 135 1680
rect 151 1676 155 1680
rect 171 1676 175 1680
rect 245 1676 249 1680
rect 265 1676 269 1680
rect 323 1676 327 1680
rect 345 1676 349 1680
rect 395 1676 399 1680
rect 415 1676 419 1680
rect 425 1676 429 1680
rect 447 1676 451 1680
rect 457 1676 461 1680
rect 479 1676 483 1680
rect 525 1676 529 1680
rect 533 1676 537 1680
rect 553 1676 557 1680
rect 563 1676 567 1680
rect 585 1676 589 1680
rect 635 1676 639 1680
rect 655 1676 659 1680
rect 665 1676 669 1680
rect 687 1676 691 1680
rect 697 1676 701 1680
rect 719 1676 723 1680
rect 765 1676 769 1680
rect 773 1676 777 1680
rect 793 1676 797 1680
rect 803 1676 807 1680
rect 825 1676 829 1680
rect 871 1676 875 1680
rect 893 1676 897 1680
rect 903 1676 907 1680
rect 923 1676 927 1680
rect 931 1676 935 1680
rect 977 1676 981 1680
rect 999 1676 1003 1680
rect 1009 1676 1013 1680
rect 1031 1676 1035 1680
rect 1041 1676 1045 1680
rect 1061 1676 1065 1680
rect 1133 1676 1137 1680
rect 1143 1676 1147 1680
rect 1205 1676 1209 1680
rect 1225 1676 1229 1680
rect 1245 1676 1249 1680
rect 1291 1676 1295 1680
rect 1313 1676 1317 1680
rect 1323 1676 1327 1680
rect 1343 1676 1347 1680
rect 1351 1676 1355 1680
rect 1397 1676 1401 1680
rect 1419 1676 1423 1680
rect 1429 1676 1433 1680
rect 1451 1676 1455 1680
rect 1461 1676 1465 1680
rect 1481 1676 1485 1680
rect 1535 1676 1539 1680
rect 1555 1676 1559 1680
rect 1565 1676 1569 1680
rect 1587 1676 1591 1680
rect 1597 1676 1601 1680
rect 1619 1676 1623 1680
rect 1665 1676 1669 1680
rect 1673 1676 1677 1680
rect 1693 1676 1697 1680
rect 1703 1676 1707 1680
rect 1725 1676 1729 1680
rect 1792 1676 1796 1680
rect 1814 1676 1818 1680
rect 1822 1676 1826 1680
rect 1871 1676 1875 1680
rect 1891 1676 1895 1680
rect 1955 1676 1959 1680
rect 1975 1676 1979 1680
rect 1985 1676 1989 1680
rect 2007 1676 2011 1680
rect 2017 1676 2021 1680
rect 2039 1676 2043 1680
rect 2085 1676 2089 1680
rect 2093 1676 2097 1680
rect 2113 1676 2117 1680
rect 2123 1676 2127 1680
rect 2145 1676 2149 1680
rect 2205 1676 2209 1680
rect 2225 1676 2229 1680
rect 2293 1676 2297 1680
rect 2303 1676 2307 1680
rect 2351 1676 2355 1680
rect 2371 1676 2375 1680
rect 2391 1676 2395 1680
rect 2451 1676 2455 1680
rect 2473 1676 2477 1680
rect 2483 1676 2487 1680
rect 2503 1676 2507 1680
rect 2511 1676 2515 1680
rect 2557 1676 2561 1680
rect 2579 1676 2583 1680
rect 2589 1676 2593 1680
rect 2611 1676 2615 1680
rect 2621 1676 2625 1680
rect 2641 1676 2645 1680
rect 2695 1676 2699 1680
rect 2715 1676 2719 1680
rect 2725 1676 2729 1680
rect 2747 1676 2751 1680
rect 2757 1676 2761 1680
rect 2779 1676 2783 1680
rect 2825 1676 2829 1680
rect 2833 1676 2837 1680
rect 2853 1676 2857 1680
rect 2863 1676 2867 1680
rect 2885 1676 2889 1680
rect 2931 1676 2935 1680
rect 2993 1676 2997 1680
rect 3003 1676 3007 1680
rect 3093 1676 3097 1680
rect 3103 1676 3107 1680
rect 3151 1676 3155 1680
rect 3171 1676 3175 1680
rect 3191 1676 3195 1680
rect 3253 1676 3257 1680
rect 3263 1676 3267 1680
rect 3353 1676 3357 1680
rect 3363 1676 3367 1680
rect 3425 1676 3429 1680
rect 3445 1676 3449 1680
rect 3465 1676 3469 1680
rect 3512 1676 3516 1680
rect 3520 1676 3524 1680
rect 3528 1676 3532 1680
rect 3625 1676 3629 1680
rect 3645 1676 3649 1680
rect 3665 1676 3669 1680
rect 3685 1676 3689 1680
rect 3731 1676 3735 1680
rect 3792 1676 3796 1680
rect 3800 1676 3804 1680
rect 3808 1676 3812 1680
rect 3894 1676 3898 1680
rect 3902 1676 3906 1680
rect 3924 1676 3928 1680
rect 3991 1676 3995 1680
rect 4011 1676 4015 1680
rect 4031 1676 4035 1680
rect 4113 1676 4117 1680
rect 4123 1676 4127 1680
rect 4174 1676 4178 1680
rect 4182 1676 4186 1680
rect 4204 1676 4208 1680
rect 4271 1676 4275 1680
rect 4291 1676 4295 1680
rect 4311 1676 4315 1680
rect 4371 1676 4375 1680
rect 4431 1676 4435 1680
rect 4451 1676 4455 1680
rect 4513 1676 4517 1680
rect 4523 1676 4527 1680
rect 4593 1676 4597 1680
rect 4603 1676 4607 1680
rect 4673 1676 4677 1680
rect 4683 1676 4687 1680
rect 31 1613 35 1636
rect 51 1613 55 1636
rect 71 1616 75 1636
rect 91 1616 95 1636
rect 111 1616 115 1636
rect 131 1616 135 1636
rect 151 1616 155 1636
rect 171 1616 175 1636
rect 31 1601 34 1613
rect 46 1601 55 1613
rect 82 1604 95 1616
rect 122 1604 135 1616
rect 162 1604 175 1616
rect 31 1544 35 1601
rect 51 1544 55 1601
rect 71 1544 75 1604
rect 91 1544 95 1604
rect 111 1544 115 1604
rect 131 1544 135 1604
rect 151 1544 155 1604
rect 171 1544 175 1604
rect 245 1579 249 1656
rect 265 1579 269 1656
rect 323 1630 327 1636
rect 323 1618 325 1630
rect 345 1579 349 1656
rect 395 1599 399 1636
rect 415 1598 419 1656
rect 425 1624 429 1656
rect 447 1644 451 1656
rect 449 1632 451 1644
rect 457 1644 461 1656
rect 457 1632 459 1644
rect 425 1620 458 1624
rect 246 1567 261 1579
rect 257 1544 261 1567
rect 265 1567 274 1579
rect 345 1567 354 1579
rect 265 1544 269 1567
rect 323 1550 325 1562
rect 323 1544 327 1550
rect 345 1504 349 1567
rect 395 1544 399 1587
rect 415 1504 419 1586
rect 434 1571 438 1600
rect 429 1563 438 1571
rect 429 1504 433 1563
rect 454 1556 458 1620
rect 455 1544 458 1556
rect 449 1504 453 1544
rect 463 1522 467 1632
rect 479 1542 483 1656
rect 525 1652 529 1656
rect 495 1648 529 1652
rect 461 1504 465 1510
rect 481 1504 485 1530
rect 495 1522 499 1648
rect 533 1644 537 1656
rect 507 1640 537 1644
rect 519 1639 537 1640
rect 553 1635 557 1656
rect 533 1631 557 1635
rect 533 1536 539 1631
rect 563 1607 567 1656
rect 563 1549 567 1595
rect 585 1568 589 1636
rect 635 1599 639 1636
rect 655 1598 659 1656
rect 665 1624 669 1656
rect 687 1644 691 1656
rect 689 1632 691 1644
rect 697 1644 701 1656
rect 697 1632 699 1644
rect 665 1620 698 1624
rect 587 1556 589 1568
rect 563 1543 571 1549
rect 585 1544 589 1556
rect 635 1544 639 1587
rect 507 1510 531 1512
rect 495 1508 531 1510
rect 527 1504 531 1508
rect 535 1504 539 1536
rect 555 1484 559 1524
rect 567 1514 571 1543
rect 563 1507 571 1514
rect 563 1484 567 1507
rect 655 1504 659 1586
rect 674 1571 678 1600
rect 669 1563 678 1571
rect 669 1504 673 1563
rect 694 1556 698 1620
rect 695 1544 698 1556
rect 689 1504 693 1544
rect 703 1522 707 1632
rect 719 1542 723 1656
rect 765 1652 769 1656
rect 735 1648 769 1652
rect 701 1504 705 1510
rect 721 1504 725 1530
rect 735 1522 739 1648
rect 773 1644 777 1656
rect 747 1640 777 1644
rect 759 1639 777 1640
rect 793 1635 797 1656
rect 773 1631 797 1635
rect 773 1536 779 1631
rect 803 1607 807 1656
rect 803 1549 807 1595
rect 825 1568 829 1636
rect 827 1556 829 1568
rect 803 1543 811 1549
rect 825 1544 829 1556
rect 871 1568 875 1636
rect 893 1607 897 1656
rect 903 1635 907 1656
rect 923 1644 927 1656
rect 931 1652 935 1656
rect 931 1648 965 1652
rect 923 1640 953 1644
rect 923 1639 941 1640
rect 903 1631 927 1635
rect 871 1556 873 1568
rect 871 1544 875 1556
rect 893 1549 897 1595
rect 747 1510 771 1512
rect 735 1508 771 1510
rect 767 1504 771 1508
rect 775 1504 779 1536
rect 795 1484 799 1524
rect 807 1514 811 1543
rect 803 1507 811 1514
rect 803 1484 807 1507
rect 889 1543 897 1549
rect 889 1514 893 1543
rect 921 1536 927 1631
rect 889 1507 897 1514
rect 893 1484 897 1507
rect 901 1484 905 1524
rect 921 1504 925 1536
rect 961 1522 965 1648
rect 977 1542 981 1656
rect 999 1644 1003 1656
rect 1001 1632 1003 1644
rect 1009 1644 1013 1656
rect 1009 1632 1011 1644
rect 929 1510 953 1512
rect 929 1508 965 1510
rect 929 1504 933 1508
rect 975 1504 979 1530
rect 993 1522 997 1632
rect 1031 1624 1035 1656
rect 1002 1620 1035 1624
rect 1002 1556 1006 1620
rect 1022 1571 1026 1600
rect 1041 1598 1045 1656
rect 1061 1599 1065 1636
rect 1133 1616 1137 1636
rect 1123 1609 1137 1616
rect 1143 1616 1147 1636
rect 1143 1609 1151 1616
rect 1123 1593 1129 1609
rect 1022 1563 1031 1571
rect 1002 1544 1005 1556
rect 995 1504 999 1510
rect 1007 1504 1011 1544
rect 1027 1504 1031 1563
rect 1041 1504 1045 1586
rect 1061 1544 1065 1587
rect 1126 1581 1129 1593
rect 1125 1504 1129 1581
rect 1145 1593 1151 1609
rect 1145 1581 1154 1593
rect 1145 1504 1149 1581
rect 1205 1559 1209 1636
rect 1225 1613 1229 1636
rect 1245 1631 1249 1636
rect 1245 1624 1258 1631
rect 1225 1601 1234 1613
rect 1207 1547 1214 1559
rect 1210 1504 1214 1547
rect 1232 1544 1236 1601
rect 1254 1579 1258 1624
rect 1291 1568 1295 1636
rect 1313 1607 1317 1656
rect 1323 1635 1327 1656
rect 1343 1644 1347 1656
rect 1351 1652 1355 1656
rect 1351 1648 1385 1652
rect 1343 1640 1373 1644
rect 1343 1639 1361 1640
rect 1323 1631 1347 1635
rect 1254 1556 1258 1567
rect 1240 1548 1258 1556
rect 1291 1556 1293 1568
rect 1240 1544 1244 1548
rect 1291 1544 1295 1556
rect 1313 1549 1317 1595
rect 1309 1543 1317 1549
rect 1309 1514 1313 1543
rect 1341 1536 1347 1631
rect 1309 1507 1317 1514
rect 1313 1484 1317 1507
rect 1321 1484 1325 1524
rect 1341 1504 1345 1536
rect 1381 1522 1385 1648
rect 1397 1542 1401 1656
rect 1419 1644 1423 1656
rect 1421 1632 1423 1644
rect 1429 1644 1433 1656
rect 1429 1632 1431 1644
rect 1349 1510 1373 1512
rect 1349 1508 1385 1510
rect 1349 1504 1353 1508
rect 1395 1504 1399 1530
rect 1413 1522 1417 1632
rect 1451 1624 1455 1656
rect 1422 1620 1455 1624
rect 1422 1556 1426 1620
rect 1442 1571 1446 1600
rect 1461 1598 1465 1656
rect 1481 1599 1485 1636
rect 1535 1599 1539 1636
rect 1555 1598 1559 1656
rect 1565 1624 1569 1656
rect 1587 1644 1591 1656
rect 1589 1632 1591 1644
rect 1597 1644 1601 1656
rect 1597 1632 1599 1644
rect 1565 1620 1598 1624
rect 1442 1563 1451 1571
rect 1422 1544 1425 1556
rect 1415 1504 1419 1510
rect 1427 1504 1431 1544
rect 1447 1504 1451 1563
rect 1461 1504 1465 1586
rect 1481 1544 1485 1587
rect 1535 1544 1539 1587
rect 1555 1504 1559 1586
rect 1574 1571 1578 1600
rect 1569 1563 1578 1571
rect 1569 1504 1573 1563
rect 1594 1556 1598 1620
rect 1595 1544 1598 1556
rect 1589 1504 1593 1544
rect 1603 1522 1607 1632
rect 1619 1542 1623 1656
rect 1665 1652 1669 1656
rect 1635 1648 1669 1652
rect 1601 1504 1605 1510
rect 1621 1504 1625 1530
rect 1635 1522 1639 1648
rect 1673 1644 1677 1656
rect 1647 1640 1677 1644
rect 1659 1639 1677 1640
rect 1693 1635 1697 1656
rect 1673 1631 1697 1635
rect 1673 1536 1679 1631
rect 1703 1607 1707 1656
rect 1703 1549 1707 1595
rect 1725 1568 1729 1636
rect 1792 1613 1796 1656
rect 1727 1556 1729 1568
rect 1703 1543 1711 1549
rect 1725 1544 1729 1556
rect 1785 1601 1794 1613
rect 1785 1544 1789 1601
rect 1814 1599 1818 1636
rect 1822 1632 1826 1636
rect 1822 1626 1841 1632
rect 1834 1613 1841 1626
rect 1814 1564 1820 1587
rect 1834 1564 1841 1601
rect 1871 1579 1875 1656
rect 1891 1579 1895 1656
rect 1955 1599 1959 1636
rect 1975 1598 1979 1656
rect 1985 1624 1989 1656
rect 2007 1644 2011 1656
rect 2009 1632 2011 1644
rect 2017 1644 2021 1656
rect 2017 1632 2019 1644
rect 1985 1620 2018 1624
rect 1866 1567 1875 1579
rect 1805 1558 1820 1564
rect 1825 1558 1841 1564
rect 1805 1544 1809 1558
rect 1825 1544 1829 1558
rect 1871 1544 1875 1567
rect 1879 1567 1894 1579
rect 1879 1544 1883 1567
rect 1955 1544 1959 1587
rect 1647 1510 1671 1512
rect 1635 1508 1671 1510
rect 1667 1504 1671 1508
rect 1675 1504 1679 1536
rect 1695 1484 1699 1524
rect 1707 1514 1711 1543
rect 1703 1507 1711 1514
rect 1703 1484 1707 1507
rect 1975 1504 1979 1586
rect 1994 1571 1998 1600
rect 1989 1563 1998 1571
rect 1989 1504 1993 1563
rect 2014 1556 2018 1620
rect 2015 1544 2018 1556
rect 2009 1504 2013 1544
rect 2023 1522 2027 1632
rect 2039 1542 2043 1656
rect 2085 1652 2089 1656
rect 2055 1648 2089 1652
rect 2021 1504 2025 1510
rect 2041 1504 2045 1530
rect 2055 1522 2059 1648
rect 2093 1644 2097 1656
rect 2067 1640 2097 1644
rect 2079 1639 2097 1640
rect 2113 1635 2117 1656
rect 2093 1631 2117 1635
rect 2093 1536 2099 1631
rect 2123 1607 2127 1656
rect 2123 1549 2127 1595
rect 2145 1568 2149 1636
rect 2205 1579 2209 1656
rect 2225 1579 2229 1656
rect 2293 1616 2297 1636
rect 2283 1609 2297 1616
rect 2303 1616 2307 1636
rect 2351 1631 2355 1636
rect 2342 1624 2355 1631
rect 2303 1609 2311 1616
rect 2283 1593 2289 1609
rect 2286 1581 2289 1593
rect 2147 1556 2149 1568
rect 2206 1567 2221 1579
rect 2123 1543 2131 1549
rect 2145 1544 2149 1556
rect 2217 1544 2221 1567
rect 2225 1567 2234 1579
rect 2225 1544 2229 1567
rect 2067 1510 2091 1512
rect 2055 1508 2091 1510
rect 2087 1504 2091 1508
rect 2095 1504 2099 1536
rect 2115 1484 2119 1524
rect 2127 1514 2131 1543
rect 2123 1507 2131 1514
rect 2123 1484 2127 1507
rect 2285 1504 2289 1581
rect 2305 1593 2311 1609
rect 2305 1581 2314 1593
rect 2305 1504 2309 1581
rect 2342 1579 2346 1624
rect 2371 1613 2375 1636
rect 2366 1601 2375 1613
rect 2342 1556 2346 1567
rect 2342 1548 2360 1556
rect 2356 1544 2360 1548
rect 2364 1544 2368 1601
rect 2391 1559 2395 1636
rect 2451 1568 2455 1636
rect 2473 1607 2477 1656
rect 2483 1635 2487 1656
rect 2503 1644 2507 1656
rect 2511 1652 2515 1656
rect 2511 1648 2545 1652
rect 2503 1640 2533 1644
rect 2503 1639 2521 1640
rect 2483 1631 2507 1635
rect 2386 1547 2393 1559
rect 2451 1556 2453 1568
rect 2386 1504 2390 1547
rect 2451 1544 2455 1556
rect 2473 1549 2477 1595
rect 2469 1543 2477 1549
rect 2469 1514 2473 1543
rect 2501 1536 2507 1631
rect 2469 1507 2477 1514
rect 2473 1484 2477 1507
rect 2481 1484 2485 1524
rect 2501 1504 2505 1536
rect 2541 1522 2545 1648
rect 2557 1542 2561 1656
rect 2579 1644 2583 1656
rect 2581 1632 2583 1644
rect 2589 1644 2593 1656
rect 2589 1632 2591 1644
rect 2509 1510 2533 1512
rect 2509 1508 2545 1510
rect 2509 1504 2513 1508
rect 2555 1504 2559 1530
rect 2573 1522 2577 1632
rect 2611 1624 2615 1656
rect 2582 1620 2615 1624
rect 2582 1556 2586 1620
rect 2602 1571 2606 1600
rect 2621 1598 2625 1656
rect 2641 1599 2645 1636
rect 2695 1599 2699 1636
rect 2715 1598 2719 1656
rect 2725 1624 2729 1656
rect 2747 1644 2751 1656
rect 2749 1632 2751 1644
rect 2757 1644 2761 1656
rect 2757 1632 2759 1644
rect 2725 1620 2758 1624
rect 2602 1563 2611 1571
rect 2582 1544 2585 1556
rect 2575 1504 2579 1510
rect 2587 1504 2591 1544
rect 2607 1504 2611 1563
rect 2621 1504 2625 1586
rect 2641 1544 2645 1587
rect 2695 1544 2699 1587
rect 2715 1504 2719 1586
rect 2734 1571 2738 1600
rect 2729 1563 2738 1571
rect 2729 1504 2733 1563
rect 2754 1556 2758 1620
rect 2755 1544 2758 1556
rect 2749 1504 2753 1544
rect 2763 1522 2767 1632
rect 2779 1542 2783 1656
rect 2825 1652 2829 1656
rect 2795 1648 2829 1652
rect 2761 1504 2765 1510
rect 2781 1504 2785 1530
rect 2795 1522 2799 1648
rect 2833 1644 2837 1656
rect 2807 1640 2837 1644
rect 2819 1639 2837 1640
rect 2853 1635 2857 1656
rect 2833 1631 2857 1635
rect 2833 1536 2839 1631
rect 2863 1607 2867 1656
rect 2863 1549 2867 1595
rect 2885 1568 2889 1636
rect 2931 1613 2935 1636
rect 2993 1616 2997 1636
rect 2926 1601 2935 1613
rect 2887 1556 2889 1568
rect 2863 1543 2871 1549
rect 2885 1544 2889 1556
rect 2931 1544 2935 1601
rect 2989 1609 2997 1616
rect 3003 1616 3007 1636
rect 3093 1616 3097 1636
rect 3003 1609 3017 1616
rect 2989 1593 2995 1609
rect 2986 1581 2995 1593
rect 2807 1510 2831 1512
rect 2795 1508 2831 1510
rect 2827 1504 2831 1508
rect 2835 1504 2839 1536
rect 2855 1484 2859 1524
rect 2867 1514 2871 1543
rect 2863 1507 2871 1514
rect 2863 1484 2867 1507
rect 2991 1504 2995 1581
rect 3011 1593 3017 1609
rect 3083 1609 3097 1616
rect 3103 1616 3107 1636
rect 3151 1631 3155 1636
rect 3142 1624 3155 1631
rect 3103 1609 3111 1616
rect 3083 1593 3089 1609
rect 3011 1581 3014 1593
rect 3086 1581 3089 1593
rect 3011 1504 3015 1581
rect 3085 1504 3089 1581
rect 3105 1593 3111 1609
rect 3105 1581 3114 1593
rect 3105 1504 3109 1581
rect 3142 1579 3146 1624
rect 3171 1613 3175 1636
rect 3166 1601 3175 1613
rect 3142 1556 3146 1567
rect 3142 1548 3160 1556
rect 3156 1544 3160 1548
rect 3164 1544 3168 1601
rect 3191 1559 3195 1636
rect 3253 1616 3257 1636
rect 3249 1609 3257 1616
rect 3263 1616 3267 1636
rect 3353 1616 3357 1636
rect 3263 1609 3277 1616
rect 3249 1593 3255 1609
rect 3246 1581 3255 1593
rect 3186 1547 3193 1559
rect 3186 1504 3190 1547
rect 3251 1504 3255 1581
rect 3271 1593 3277 1609
rect 3343 1609 3357 1616
rect 3363 1616 3367 1636
rect 3363 1609 3371 1616
rect 3343 1593 3349 1609
rect 3271 1581 3274 1593
rect 3346 1581 3349 1593
rect 3271 1504 3275 1581
rect 3345 1504 3349 1581
rect 3365 1593 3371 1609
rect 3365 1581 3374 1593
rect 3365 1504 3369 1581
rect 3425 1559 3429 1636
rect 3445 1613 3449 1636
rect 3465 1631 3469 1636
rect 3465 1624 3478 1631
rect 3445 1601 3454 1613
rect 3427 1547 3434 1559
rect 3430 1504 3434 1547
rect 3452 1544 3456 1601
rect 3474 1579 3478 1624
rect 3474 1556 3478 1567
rect 3512 1559 3516 1616
rect 3460 1548 3478 1556
rect 3460 1544 3464 1548
rect 3506 1547 3516 1559
rect 3500 1516 3506 1547
rect 3520 1539 3524 1616
rect 3528 1559 3532 1616
rect 3625 1579 3629 1636
rect 3645 1613 3649 1636
rect 3665 1613 3669 1636
rect 3685 1629 3689 1636
rect 3685 1625 3700 1629
rect 3665 1601 3674 1613
rect 3627 1567 3629 1579
rect 3528 1547 3535 1559
rect 3547 1547 3555 1559
rect 3625 1552 3629 1567
rect 3625 1548 3639 1552
rect 3520 1520 3526 1527
rect 3520 1516 3535 1520
rect 3500 1512 3515 1516
rect 3511 1504 3515 1512
rect 3531 1504 3535 1516
rect 3551 1504 3555 1547
rect 3635 1544 3639 1548
rect 3645 1544 3649 1601
rect 3665 1552 3671 1601
rect 3694 1579 3700 1625
rect 3731 1599 3735 1656
rect 3894 1632 3898 1636
rect 3879 1626 3898 1632
rect 3726 1587 3735 1599
rect 3694 1552 3699 1567
rect 3665 1548 3679 1552
rect 3675 1544 3679 1548
rect 3685 1548 3699 1552
rect 3685 1544 3689 1548
rect 3731 1504 3735 1587
rect 3792 1559 3796 1616
rect 3786 1547 3796 1559
rect 3780 1516 3786 1547
rect 3800 1539 3804 1616
rect 3808 1559 3812 1616
rect 3879 1613 3886 1626
rect 3879 1564 3886 1601
rect 3902 1599 3906 1636
rect 3924 1613 3928 1656
rect 3991 1631 3995 1636
rect 3982 1624 3995 1631
rect 3926 1601 3935 1613
rect 3900 1564 3906 1587
rect 3808 1547 3815 1559
rect 3827 1547 3835 1559
rect 3879 1558 3895 1564
rect 3900 1558 3915 1564
rect 3800 1520 3806 1527
rect 3800 1516 3815 1520
rect 3780 1512 3795 1516
rect 3791 1504 3795 1512
rect 3811 1504 3815 1516
rect 3831 1504 3835 1547
rect 3891 1544 3895 1558
rect 3911 1544 3915 1558
rect 3931 1544 3935 1601
rect 3982 1579 3986 1624
rect 4011 1613 4015 1636
rect 4006 1601 4015 1613
rect 3982 1556 3986 1567
rect 3982 1548 4000 1556
rect 3996 1544 4000 1548
rect 4004 1544 4008 1601
rect 4031 1559 4035 1636
rect 4113 1616 4117 1636
rect 4103 1609 4117 1616
rect 4123 1616 4127 1636
rect 4174 1632 4178 1636
rect 4159 1626 4178 1632
rect 4123 1609 4131 1616
rect 4159 1613 4166 1626
rect 4103 1593 4109 1609
rect 4106 1581 4109 1593
rect 4026 1547 4033 1559
rect 4026 1504 4030 1547
rect 4105 1504 4109 1581
rect 4125 1593 4131 1609
rect 4125 1581 4134 1593
rect 4125 1504 4129 1581
rect 4159 1564 4166 1601
rect 4182 1599 4186 1636
rect 4204 1613 4208 1656
rect 4271 1631 4275 1636
rect 4262 1624 4275 1631
rect 4206 1601 4215 1613
rect 4180 1564 4186 1587
rect 4159 1558 4175 1564
rect 4180 1558 4195 1564
rect 4171 1544 4175 1558
rect 4191 1544 4195 1558
rect 4211 1544 4215 1601
rect 4262 1579 4266 1624
rect 4291 1613 4295 1636
rect 4286 1601 4295 1613
rect 4262 1556 4266 1567
rect 4262 1548 4280 1556
rect 4276 1544 4280 1548
rect 4284 1544 4288 1601
rect 4311 1559 4315 1636
rect 4371 1599 4375 1656
rect 4366 1587 4375 1599
rect 4306 1547 4313 1559
rect 4306 1504 4310 1547
rect 4371 1504 4375 1587
rect 4431 1579 4435 1656
rect 4451 1579 4455 1656
rect 4513 1616 4517 1636
rect 4509 1609 4517 1616
rect 4523 1616 4527 1636
rect 4593 1616 4597 1636
rect 4523 1609 4537 1616
rect 4509 1593 4515 1609
rect 4506 1581 4515 1593
rect 4426 1567 4435 1579
rect 4431 1544 4435 1567
rect 4439 1567 4454 1579
rect 4439 1544 4443 1567
rect 4511 1504 4515 1581
rect 4531 1593 4537 1609
rect 4589 1609 4597 1616
rect 4603 1616 4607 1636
rect 4673 1616 4677 1636
rect 4603 1609 4617 1616
rect 4589 1593 4595 1609
rect 4531 1581 4534 1593
rect 4586 1581 4595 1593
rect 4531 1504 4535 1581
rect 4591 1504 4595 1581
rect 4611 1593 4617 1609
rect 4669 1609 4677 1616
rect 4683 1616 4687 1636
rect 4683 1609 4697 1616
rect 4669 1593 4675 1609
rect 4611 1581 4614 1593
rect 4666 1581 4675 1593
rect 4611 1504 4615 1581
rect 4671 1504 4675 1581
rect 4691 1593 4697 1609
rect 4691 1581 4694 1593
rect 4691 1504 4695 1581
rect 31 1460 35 1464
rect 51 1460 55 1464
rect 71 1460 75 1464
rect 91 1460 95 1464
rect 111 1460 115 1464
rect 131 1460 135 1464
rect 151 1460 155 1464
rect 171 1460 175 1464
rect 257 1460 261 1464
rect 265 1460 269 1464
rect 323 1460 327 1464
rect 345 1460 349 1464
rect 395 1460 399 1464
rect 415 1460 419 1464
rect 429 1460 433 1464
rect 449 1460 453 1464
rect 461 1460 465 1464
rect 481 1460 485 1464
rect 527 1460 531 1464
rect 535 1460 539 1464
rect 555 1460 559 1464
rect 563 1460 567 1464
rect 585 1460 589 1464
rect 635 1460 639 1464
rect 655 1460 659 1464
rect 669 1460 673 1464
rect 689 1460 693 1464
rect 701 1460 705 1464
rect 721 1460 725 1464
rect 767 1460 771 1464
rect 775 1460 779 1464
rect 795 1460 799 1464
rect 803 1460 807 1464
rect 825 1460 829 1464
rect 871 1460 875 1464
rect 893 1460 897 1464
rect 901 1460 905 1464
rect 921 1460 925 1464
rect 929 1460 933 1464
rect 975 1460 979 1464
rect 995 1460 999 1464
rect 1007 1460 1011 1464
rect 1027 1460 1031 1464
rect 1041 1460 1045 1464
rect 1061 1460 1065 1464
rect 1125 1460 1129 1464
rect 1145 1460 1149 1464
rect 1210 1460 1214 1464
rect 1232 1460 1236 1464
rect 1240 1460 1244 1464
rect 1291 1460 1295 1464
rect 1313 1460 1317 1464
rect 1321 1460 1325 1464
rect 1341 1460 1345 1464
rect 1349 1460 1353 1464
rect 1395 1460 1399 1464
rect 1415 1460 1419 1464
rect 1427 1460 1431 1464
rect 1447 1460 1451 1464
rect 1461 1460 1465 1464
rect 1481 1460 1485 1464
rect 1535 1460 1539 1464
rect 1555 1460 1559 1464
rect 1569 1460 1573 1464
rect 1589 1460 1593 1464
rect 1601 1460 1605 1464
rect 1621 1460 1625 1464
rect 1667 1460 1671 1464
rect 1675 1460 1679 1464
rect 1695 1460 1699 1464
rect 1703 1460 1707 1464
rect 1725 1460 1729 1464
rect 1785 1460 1789 1464
rect 1805 1460 1809 1464
rect 1825 1460 1829 1464
rect 1871 1460 1875 1464
rect 1879 1460 1883 1464
rect 1955 1460 1959 1464
rect 1975 1460 1979 1464
rect 1989 1460 1993 1464
rect 2009 1460 2013 1464
rect 2021 1460 2025 1464
rect 2041 1460 2045 1464
rect 2087 1460 2091 1464
rect 2095 1460 2099 1464
rect 2115 1460 2119 1464
rect 2123 1460 2127 1464
rect 2145 1460 2149 1464
rect 2217 1460 2221 1464
rect 2225 1460 2229 1464
rect 2285 1460 2289 1464
rect 2305 1460 2309 1464
rect 2356 1460 2360 1464
rect 2364 1460 2368 1464
rect 2386 1460 2390 1464
rect 2451 1460 2455 1464
rect 2473 1460 2477 1464
rect 2481 1460 2485 1464
rect 2501 1460 2505 1464
rect 2509 1460 2513 1464
rect 2555 1460 2559 1464
rect 2575 1460 2579 1464
rect 2587 1460 2591 1464
rect 2607 1460 2611 1464
rect 2621 1460 2625 1464
rect 2641 1460 2645 1464
rect 2695 1460 2699 1464
rect 2715 1460 2719 1464
rect 2729 1460 2733 1464
rect 2749 1460 2753 1464
rect 2761 1460 2765 1464
rect 2781 1460 2785 1464
rect 2827 1460 2831 1464
rect 2835 1460 2839 1464
rect 2855 1460 2859 1464
rect 2863 1460 2867 1464
rect 2885 1460 2889 1464
rect 2931 1460 2935 1464
rect 2991 1460 2995 1464
rect 3011 1460 3015 1464
rect 3085 1460 3089 1464
rect 3105 1460 3109 1464
rect 3156 1460 3160 1464
rect 3164 1460 3168 1464
rect 3186 1460 3190 1464
rect 3251 1460 3255 1464
rect 3271 1460 3275 1464
rect 3345 1460 3349 1464
rect 3365 1460 3369 1464
rect 3430 1460 3434 1464
rect 3452 1460 3456 1464
rect 3460 1460 3464 1464
rect 3511 1460 3515 1464
rect 3531 1460 3535 1464
rect 3551 1460 3555 1464
rect 3635 1460 3639 1464
rect 3645 1460 3649 1464
rect 3675 1460 3679 1464
rect 3685 1460 3689 1464
rect 3731 1460 3735 1464
rect 3791 1460 3795 1464
rect 3811 1460 3815 1464
rect 3831 1460 3835 1464
rect 3891 1460 3895 1464
rect 3911 1460 3915 1464
rect 3931 1460 3935 1464
rect 3996 1460 4000 1464
rect 4004 1460 4008 1464
rect 4026 1460 4030 1464
rect 4105 1460 4109 1464
rect 4125 1460 4129 1464
rect 4171 1460 4175 1464
rect 4191 1460 4195 1464
rect 4211 1460 4215 1464
rect 4276 1460 4280 1464
rect 4284 1460 4288 1464
rect 4306 1460 4310 1464
rect 4371 1460 4375 1464
rect 4431 1460 4435 1464
rect 4439 1460 4443 1464
rect 4511 1460 4515 1464
rect 4531 1460 4535 1464
rect 4591 1460 4595 1464
rect 4611 1460 4615 1464
rect 4671 1460 4675 1464
rect 4691 1460 4695 1464
rect 31 1436 35 1440
rect 53 1436 57 1440
rect 61 1436 65 1440
rect 81 1436 85 1440
rect 89 1436 93 1440
rect 135 1436 139 1440
rect 155 1436 159 1440
rect 167 1436 171 1440
rect 187 1436 191 1440
rect 201 1436 205 1440
rect 221 1436 225 1440
rect 275 1436 279 1440
rect 295 1436 299 1440
rect 309 1436 313 1440
rect 329 1436 333 1440
rect 341 1436 345 1440
rect 361 1436 365 1440
rect 407 1436 411 1440
rect 415 1436 419 1440
rect 435 1436 439 1440
rect 443 1436 447 1440
rect 465 1436 469 1440
rect 511 1436 515 1440
rect 531 1436 535 1440
rect 610 1436 614 1440
rect 632 1436 636 1440
rect 640 1436 644 1440
rect 710 1436 714 1440
rect 732 1436 736 1440
rect 740 1436 744 1440
rect 803 1436 807 1440
rect 825 1436 829 1440
rect 871 1436 875 1440
rect 891 1436 895 1440
rect 970 1436 974 1440
rect 992 1436 996 1440
rect 1000 1436 1004 1440
rect 1065 1436 1069 1440
rect 1111 1436 1115 1440
rect 1131 1436 1135 1440
rect 1151 1436 1155 1440
rect 1171 1436 1175 1440
rect 1245 1436 1249 1440
rect 1265 1436 1269 1440
rect 1330 1436 1334 1440
rect 1352 1436 1356 1440
rect 1360 1436 1364 1440
rect 1425 1436 1429 1440
rect 1445 1436 1449 1440
rect 1510 1436 1514 1440
rect 1532 1436 1536 1440
rect 1540 1436 1544 1440
rect 1591 1436 1595 1440
rect 1613 1436 1617 1440
rect 1671 1436 1675 1440
rect 1691 1436 1695 1440
rect 1770 1436 1774 1440
rect 1792 1436 1796 1440
rect 1800 1436 1804 1440
rect 1851 1436 1855 1440
rect 1873 1436 1877 1440
rect 1881 1436 1885 1440
rect 1901 1436 1905 1440
rect 1909 1436 1913 1440
rect 1955 1436 1959 1440
rect 1975 1436 1979 1440
rect 1987 1436 1991 1440
rect 2007 1436 2011 1440
rect 2021 1436 2025 1440
rect 2041 1436 2045 1440
rect 2091 1436 2095 1440
rect 2156 1436 2160 1440
rect 2164 1436 2168 1440
rect 2186 1436 2190 1440
rect 2265 1436 2269 1440
rect 2285 1436 2289 1440
rect 2357 1436 2361 1440
rect 2365 1436 2369 1440
rect 2425 1436 2429 1440
rect 2471 1436 2475 1440
rect 2479 1436 2483 1440
rect 2551 1436 2555 1440
rect 2573 1436 2577 1440
rect 2581 1436 2585 1440
rect 2601 1436 2605 1440
rect 2609 1436 2613 1440
rect 2655 1436 2659 1440
rect 2675 1436 2679 1440
rect 2687 1436 2691 1440
rect 2707 1436 2711 1440
rect 2721 1436 2725 1440
rect 2741 1436 2745 1440
rect 2791 1436 2795 1440
rect 2799 1436 2803 1440
rect 2885 1436 2889 1440
rect 2936 1436 2940 1440
rect 2944 1436 2948 1440
rect 2966 1436 2970 1440
rect 3036 1436 3040 1440
rect 3044 1436 3048 1440
rect 3066 1436 3070 1440
rect 3136 1436 3140 1440
rect 3144 1436 3148 1440
rect 3166 1436 3170 1440
rect 3231 1436 3235 1440
rect 3253 1436 3257 1440
rect 3275 1436 3279 1440
rect 3357 1436 3361 1440
rect 3365 1436 3369 1440
rect 3411 1436 3415 1440
rect 3431 1436 3435 1440
rect 3451 1436 3455 1440
rect 3530 1436 3534 1440
rect 3552 1436 3556 1440
rect 3560 1436 3564 1440
rect 3616 1436 3620 1440
rect 3624 1436 3628 1440
rect 3646 1436 3650 1440
rect 3725 1436 3729 1440
rect 3745 1436 3749 1440
rect 3805 1436 3809 1440
rect 3825 1436 3829 1440
rect 3871 1436 3875 1440
rect 3893 1436 3897 1440
rect 3915 1436 3919 1440
rect 3990 1436 3994 1440
rect 4012 1436 4016 1440
rect 4020 1436 4024 1440
rect 4071 1436 4075 1440
rect 4145 1436 4149 1440
rect 4165 1436 4169 1440
rect 4225 1436 4229 1440
rect 4245 1436 4249 1440
rect 4317 1436 4321 1440
rect 4325 1436 4329 1440
rect 4390 1436 4394 1440
rect 4412 1436 4416 1440
rect 4420 1436 4424 1440
rect 4476 1436 4480 1440
rect 4484 1436 4488 1440
rect 4506 1436 4510 1440
rect 4585 1436 4589 1440
rect 4605 1436 4609 1440
rect 4625 1436 4629 1440
rect 4671 1436 4675 1440
rect 4691 1436 4695 1440
rect 53 1393 57 1416
rect 49 1386 57 1393
rect 49 1357 53 1386
rect 61 1376 65 1416
rect 81 1364 85 1396
rect 89 1392 93 1396
rect 89 1390 125 1392
rect 89 1388 113 1390
rect 31 1344 35 1356
rect 49 1351 57 1357
rect 31 1332 33 1344
rect 31 1264 35 1332
rect 53 1305 57 1351
rect 53 1244 57 1293
rect 81 1269 87 1364
rect 63 1265 87 1269
rect 63 1244 67 1265
rect 83 1260 101 1261
rect 83 1256 113 1260
rect 83 1244 87 1256
rect 121 1252 125 1378
rect 135 1370 139 1396
rect 155 1390 159 1396
rect 91 1248 125 1252
rect 91 1244 95 1248
rect 137 1244 141 1358
rect 153 1268 157 1378
rect 167 1356 171 1396
rect 162 1344 165 1356
rect 162 1280 166 1344
rect 187 1337 191 1396
rect 182 1329 191 1337
rect 182 1300 186 1329
rect 201 1314 205 1396
rect 221 1313 225 1356
rect 275 1313 279 1356
rect 295 1314 299 1396
rect 309 1337 313 1396
rect 329 1356 333 1396
rect 341 1390 345 1396
rect 335 1344 338 1356
rect 309 1329 318 1337
rect 162 1276 195 1280
rect 161 1256 163 1268
rect 159 1244 163 1256
rect 169 1256 171 1268
rect 169 1244 173 1256
rect 191 1244 195 1276
rect 201 1244 205 1302
rect 221 1264 225 1301
rect 275 1264 279 1301
rect 295 1244 299 1302
rect 314 1300 318 1329
rect 334 1280 338 1344
rect 305 1276 338 1280
rect 305 1244 309 1276
rect 343 1268 347 1378
rect 361 1370 365 1396
rect 407 1392 411 1396
rect 375 1390 411 1392
rect 387 1388 411 1390
rect 329 1256 331 1268
rect 327 1244 331 1256
rect 337 1256 339 1268
rect 337 1244 341 1256
rect 359 1244 363 1358
rect 375 1252 379 1378
rect 415 1364 419 1396
rect 435 1376 439 1416
rect 443 1393 447 1416
rect 443 1386 451 1393
rect 413 1269 419 1364
rect 447 1357 451 1386
rect 443 1351 451 1357
rect 443 1305 447 1351
rect 465 1344 469 1356
rect 467 1332 469 1344
rect 413 1265 437 1269
rect 399 1260 417 1261
rect 387 1256 417 1260
rect 375 1248 409 1252
rect 405 1244 409 1248
rect 413 1244 417 1256
rect 433 1244 437 1265
rect 443 1244 447 1293
rect 465 1264 469 1332
rect 511 1319 515 1396
rect 506 1307 515 1319
rect 509 1291 515 1307
rect 531 1319 535 1396
rect 610 1353 614 1396
rect 607 1341 614 1353
rect 531 1307 534 1319
rect 531 1291 537 1307
rect 509 1284 517 1291
rect 513 1264 517 1284
rect 523 1284 537 1291
rect 523 1264 527 1284
rect 605 1264 609 1341
rect 632 1299 636 1356
rect 640 1352 644 1356
rect 710 1353 714 1396
rect 640 1344 658 1352
rect 654 1333 658 1344
rect 707 1341 714 1353
rect 625 1287 634 1299
rect 625 1264 629 1287
rect 654 1276 658 1321
rect 645 1269 658 1276
rect 645 1264 649 1269
rect 705 1264 709 1341
rect 732 1299 736 1356
rect 740 1352 744 1356
rect 740 1344 758 1352
rect 754 1333 758 1344
rect 803 1350 807 1356
rect 803 1338 805 1350
rect 825 1333 829 1396
rect 825 1321 834 1333
rect 725 1287 734 1299
rect 725 1264 729 1287
rect 754 1276 758 1321
rect 745 1269 758 1276
rect 803 1270 805 1282
rect 745 1264 749 1269
rect 803 1264 807 1270
rect 825 1244 829 1321
rect 871 1319 875 1396
rect 866 1307 875 1319
rect 869 1291 875 1307
rect 891 1319 895 1396
rect 970 1353 974 1396
rect 967 1341 974 1353
rect 891 1307 894 1319
rect 891 1291 897 1307
rect 869 1284 877 1291
rect 873 1264 877 1284
rect 883 1284 897 1291
rect 883 1264 887 1284
rect 965 1264 969 1341
rect 992 1299 996 1356
rect 1000 1352 1004 1356
rect 1000 1344 1018 1352
rect 1014 1333 1018 1344
rect 985 1287 994 1299
rect 985 1264 989 1287
rect 1014 1276 1018 1321
rect 1005 1269 1018 1276
rect 1065 1313 1069 1396
rect 1111 1352 1115 1356
rect 1131 1352 1135 1356
rect 1151 1352 1155 1356
rect 1171 1352 1175 1356
rect 1111 1348 1175 1352
rect 1111 1333 1117 1348
rect 1111 1321 1114 1333
rect 1065 1301 1074 1313
rect 1005 1264 1009 1269
rect 1065 1244 1069 1301
rect 1111 1272 1117 1321
rect 1245 1319 1249 1396
rect 1246 1307 1249 1319
rect 1243 1291 1249 1307
rect 1265 1319 1269 1396
rect 1330 1353 1334 1396
rect 1327 1341 1334 1353
rect 1265 1307 1274 1319
rect 1265 1291 1271 1307
rect 1243 1284 1257 1291
rect 1111 1268 1175 1272
rect 1111 1264 1115 1268
rect 1131 1264 1135 1268
rect 1151 1264 1155 1268
rect 1171 1264 1175 1268
rect 1253 1264 1257 1284
rect 1263 1284 1271 1291
rect 1263 1264 1267 1284
rect 1325 1264 1329 1341
rect 1352 1299 1356 1356
rect 1360 1352 1364 1356
rect 1360 1344 1378 1352
rect 1374 1333 1378 1344
rect 1345 1287 1354 1299
rect 1345 1264 1349 1287
rect 1374 1276 1378 1321
rect 1425 1319 1429 1396
rect 1426 1307 1429 1319
rect 1423 1291 1429 1307
rect 1445 1319 1449 1396
rect 1510 1353 1514 1396
rect 1507 1341 1514 1353
rect 1445 1307 1454 1319
rect 1445 1291 1451 1307
rect 1423 1284 1437 1291
rect 1365 1269 1378 1276
rect 1365 1264 1369 1269
rect 1433 1264 1437 1284
rect 1443 1284 1451 1291
rect 1443 1264 1447 1284
rect 1505 1264 1509 1341
rect 1532 1299 1536 1356
rect 1540 1352 1544 1356
rect 1540 1344 1558 1352
rect 1554 1333 1558 1344
rect 1591 1333 1595 1396
rect 1613 1350 1617 1356
rect 1615 1338 1617 1350
rect 1586 1321 1595 1333
rect 1525 1287 1534 1299
rect 1525 1264 1529 1287
rect 1554 1276 1558 1321
rect 1545 1269 1558 1276
rect 1545 1264 1549 1269
rect 1591 1244 1595 1321
rect 1671 1319 1675 1396
rect 1666 1307 1675 1319
rect 1669 1291 1675 1307
rect 1691 1319 1695 1396
rect 1770 1353 1774 1396
rect 1873 1393 1877 1416
rect 1869 1386 1877 1393
rect 1869 1357 1873 1386
rect 1881 1376 1885 1416
rect 1901 1364 1905 1396
rect 1909 1392 1913 1396
rect 1909 1390 1945 1392
rect 1909 1388 1933 1390
rect 1767 1341 1774 1353
rect 1691 1307 1694 1319
rect 1691 1291 1697 1307
rect 1669 1284 1677 1291
rect 1615 1270 1617 1282
rect 1613 1264 1617 1270
rect 1673 1264 1677 1284
rect 1683 1284 1697 1291
rect 1683 1264 1687 1284
rect 1765 1264 1769 1341
rect 1792 1299 1796 1356
rect 1800 1352 1804 1356
rect 1800 1344 1818 1352
rect 1814 1333 1818 1344
rect 1851 1344 1855 1356
rect 1869 1351 1877 1357
rect 1851 1332 1853 1344
rect 1785 1287 1794 1299
rect 1785 1264 1789 1287
rect 1814 1276 1818 1321
rect 1805 1269 1818 1276
rect 1805 1264 1809 1269
rect 1851 1264 1855 1332
rect 1873 1305 1877 1351
rect 1873 1244 1877 1293
rect 1901 1269 1907 1364
rect 1883 1265 1907 1269
rect 1883 1244 1887 1265
rect 1903 1260 1921 1261
rect 1903 1256 1933 1260
rect 1903 1244 1907 1256
rect 1941 1252 1945 1378
rect 1955 1370 1959 1396
rect 1975 1390 1979 1396
rect 1911 1248 1945 1252
rect 1911 1244 1915 1248
rect 1957 1244 1961 1358
rect 1973 1268 1977 1378
rect 1987 1356 1991 1396
rect 1982 1344 1985 1356
rect 1982 1280 1986 1344
rect 2007 1337 2011 1396
rect 2002 1329 2011 1337
rect 2002 1300 2006 1329
rect 2021 1314 2025 1396
rect 2041 1313 2045 1356
rect 2091 1313 2095 1396
rect 2156 1352 2160 1356
rect 2142 1344 2160 1352
rect 2142 1333 2146 1344
rect 1982 1276 2015 1280
rect 1981 1256 1983 1268
rect 1979 1244 1983 1256
rect 1989 1256 1991 1268
rect 1989 1244 1993 1256
rect 2011 1244 2015 1276
rect 2021 1244 2025 1302
rect 2086 1301 2095 1313
rect 2041 1264 2045 1301
rect 2091 1244 2095 1301
rect 2142 1276 2146 1321
rect 2164 1299 2168 1356
rect 2186 1353 2190 1396
rect 2186 1341 2193 1353
rect 2166 1287 2175 1299
rect 2142 1269 2155 1276
rect 2151 1264 2155 1269
rect 2171 1264 2175 1287
rect 2191 1264 2195 1341
rect 2265 1319 2269 1396
rect 2266 1307 2269 1319
rect 2263 1291 2269 1307
rect 2285 1319 2289 1396
rect 2357 1333 2361 1356
rect 2346 1321 2361 1333
rect 2365 1333 2369 1356
rect 2365 1321 2374 1333
rect 2285 1307 2294 1319
rect 2285 1291 2291 1307
rect 2263 1284 2277 1291
rect 2273 1264 2277 1284
rect 2283 1284 2291 1291
rect 2283 1264 2287 1284
rect 2345 1244 2349 1321
rect 2365 1244 2369 1321
rect 2425 1313 2429 1396
rect 2573 1393 2577 1416
rect 2569 1386 2577 1393
rect 2569 1357 2573 1386
rect 2581 1376 2585 1416
rect 2601 1364 2605 1396
rect 2609 1392 2613 1396
rect 2609 1390 2645 1392
rect 2609 1388 2633 1390
rect 2471 1333 2475 1356
rect 2466 1321 2475 1333
rect 2479 1333 2483 1356
rect 2551 1344 2555 1356
rect 2569 1351 2577 1357
rect 2479 1321 2494 1333
rect 2551 1332 2553 1344
rect 2425 1301 2434 1313
rect 2425 1244 2429 1301
rect 2471 1244 2475 1321
rect 2491 1244 2495 1321
rect 2551 1264 2555 1332
rect 2573 1305 2577 1351
rect 2573 1244 2577 1293
rect 2601 1269 2607 1364
rect 2583 1265 2607 1269
rect 2583 1244 2587 1265
rect 2603 1260 2621 1261
rect 2603 1256 2633 1260
rect 2603 1244 2607 1256
rect 2641 1252 2645 1378
rect 2655 1370 2659 1396
rect 2675 1390 2679 1396
rect 2611 1248 2645 1252
rect 2611 1244 2615 1248
rect 2657 1244 2661 1358
rect 2673 1268 2677 1378
rect 2687 1356 2691 1396
rect 2682 1344 2685 1356
rect 2682 1280 2686 1344
rect 2707 1337 2711 1396
rect 2702 1329 2711 1337
rect 2702 1300 2706 1329
rect 2721 1314 2725 1396
rect 2741 1313 2745 1356
rect 2791 1333 2795 1356
rect 2786 1321 2795 1333
rect 2799 1333 2803 1356
rect 2799 1321 2814 1333
rect 2682 1276 2715 1280
rect 2681 1256 2683 1268
rect 2679 1244 2683 1256
rect 2689 1256 2691 1268
rect 2689 1244 2693 1256
rect 2711 1244 2715 1276
rect 2721 1244 2725 1302
rect 2741 1264 2745 1301
rect 2791 1244 2795 1321
rect 2811 1244 2815 1321
rect 2885 1299 2889 1356
rect 2936 1352 2940 1356
rect 2922 1344 2940 1352
rect 2922 1333 2926 1344
rect 2885 1287 2894 1299
rect 2885 1264 2889 1287
rect 2922 1276 2926 1321
rect 2944 1299 2948 1356
rect 2966 1353 2970 1396
rect 2966 1341 2973 1353
rect 3036 1352 3040 1356
rect 3022 1344 3040 1352
rect 2946 1287 2955 1299
rect 2922 1269 2935 1276
rect 2931 1264 2935 1269
rect 2951 1264 2955 1287
rect 2971 1264 2975 1341
rect 3022 1333 3026 1344
rect 3022 1276 3026 1321
rect 3044 1299 3048 1356
rect 3066 1353 3070 1396
rect 3066 1341 3073 1353
rect 3136 1352 3140 1356
rect 3122 1344 3140 1352
rect 3046 1287 3055 1299
rect 3022 1269 3035 1276
rect 3031 1264 3035 1269
rect 3051 1264 3055 1287
rect 3071 1264 3075 1341
rect 3122 1333 3126 1344
rect 3122 1276 3126 1321
rect 3144 1299 3148 1356
rect 3166 1353 3170 1396
rect 3166 1341 3173 1353
rect 3146 1287 3155 1299
rect 3122 1269 3135 1276
rect 3131 1264 3135 1269
rect 3151 1264 3155 1287
rect 3171 1264 3175 1341
rect 3231 1333 3235 1396
rect 3226 1321 3235 1333
rect 3231 1264 3235 1321
rect 3253 1319 3257 1396
rect 3411 1388 3415 1396
rect 3400 1384 3415 1388
rect 3431 1384 3435 1396
rect 3241 1307 3254 1319
rect 3241 1264 3245 1307
rect 3275 1282 3279 1356
rect 3357 1333 3361 1356
rect 3346 1321 3361 1333
rect 3365 1333 3369 1356
rect 3400 1353 3406 1384
rect 3420 1380 3435 1384
rect 3420 1373 3426 1380
rect 3406 1341 3416 1353
rect 3365 1321 3374 1333
rect 3267 1270 3279 1282
rect 3261 1264 3265 1270
rect 3345 1244 3349 1321
rect 3365 1244 3369 1321
rect 3412 1284 3416 1341
rect 3420 1284 3424 1361
rect 3451 1353 3455 1396
rect 3530 1353 3534 1396
rect 3428 1341 3435 1353
rect 3447 1341 3455 1353
rect 3527 1341 3534 1353
rect 3428 1284 3432 1341
rect 3525 1264 3529 1341
rect 3552 1299 3556 1356
rect 3560 1352 3564 1356
rect 3616 1352 3620 1356
rect 3560 1344 3578 1352
rect 3574 1333 3578 1344
rect 3602 1344 3620 1352
rect 3602 1333 3606 1344
rect 3545 1287 3554 1299
rect 3545 1264 3549 1287
rect 3574 1276 3578 1321
rect 3565 1269 3578 1276
rect 3602 1276 3606 1321
rect 3624 1299 3628 1356
rect 3646 1353 3650 1396
rect 3646 1341 3653 1353
rect 3626 1287 3635 1299
rect 3602 1269 3615 1276
rect 3565 1264 3569 1269
rect 3611 1264 3615 1269
rect 3631 1264 3635 1287
rect 3651 1264 3655 1341
rect 3725 1319 3729 1396
rect 3726 1307 3729 1319
rect 3723 1291 3729 1307
rect 3745 1319 3749 1396
rect 3805 1319 3809 1396
rect 3745 1307 3754 1319
rect 3806 1307 3809 1319
rect 3745 1291 3751 1307
rect 3723 1284 3737 1291
rect 3733 1264 3737 1284
rect 3743 1284 3751 1291
rect 3803 1291 3809 1307
rect 3825 1319 3829 1396
rect 3871 1333 3875 1396
rect 3866 1321 3875 1333
rect 3825 1307 3834 1319
rect 3825 1291 3831 1307
rect 3803 1284 3817 1291
rect 3743 1264 3747 1284
rect 3813 1264 3817 1284
rect 3823 1284 3831 1291
rect 3823 1264 3827 1284
rect 3871 1264 3875 1321
rect 3893 1319 3897 1396
rect 3881 1307 3894 1319
rect 3881 1264 3885 1307
rect 3915 1282 3919 1356
rect 3990 1353 3994 1396
rect 3987 1341 3994 1353
rect 3907 1270 3919 1282
rect 3901 1264 3905 1270
rect 3985 1264 3989 1341
rect 4012 1299 4016 1356
rect 4020 1352 4024 1356
rect 4020 1344 4038 1352
rect 4034 1333 4038 1344
rect 4005 1287 4014 1299
rect 4005 1264 4009 1287
rect 4034 1276 4038 1321
rect 4071 1313 4075 1396
rect 4145 1319 4149 1396
rect 4066 1301 4075 1313
rect 4146 1307 4149 1319
rect 4025 1269 4038 1276
rect 4025 1264 4029 1269
rect 4071 1244 4075 1301
rect 4143 1291 4149 1307
rect 4165 1319 4169 1396
rect 4225 1319 4229 1396
rect 4165 1307 4174 1319
rect 4226 1307 4229 1319
rect 4165 1291 4171 1307
rect 4143 1284 4157 1291
rect 4153 1264 4157 1284
rect 4163 1284 4171 1291
rect 4223 1291 4229 1307
rect 4245 1319 4249 1396
rect 4317 1333 4321 1356
rect 4306 1321 4321 1333
rect 4325 1333 4329 1356
rect 4390 1353 4394 1396
rect 4387 1341 4394 1353
rect 4325 1321 4334 1333
rect 4245 1307 4254 1319
rect 4245 1291 4251 1307
rect 4223 1284 4237 1291
rect 4163 1264 4167 1284
rect 4233 1264 4237 1284
rect 4243 1284 4251 1291
rect 4243 1264 4247 1284
rect 4305 1244 4309 1321
rect 4325 1244 4329 1321
rect 4385 1264 4389 1341
rect 4412 1299 4416 1356
rect 4420 1352 4424 1356
rect 4476 1352 4480 1356
rect 4420 1344 4438 1352
rect 4434 1333 4438 1344
rect 4462 1344 4480 1352
rect 4462 1333 4466 1344
rect 4405 1287 4414 1299
rect 4405 1264 4409 1287
rect 4434 1276 4438 1321
rect 4425 1269 4438 1276
rect 4462 1276 4466 1321
rect 4484 1299 4488 1356
rect 4506 1353 4510 1396
rect 4506 1341 4513 1353
rect 4486 1287 4495 1299
rect 4462 1269 4475 1276
rect 4425 1264 4429 1269
rect 4471 1264 4475 1269
rect 4491 1264 4495 1287
rect 4511 1264 4515 1341
rect 4585 1299 4589 1356
rect 4605 1342 4609 1356
rect 4625 1342 4629 1356
rect 4605 1336 4620 1342
rect 4625 1336 4641 1342
rect 4614 1313 4620 1336
rect 4585 1287 4594 1299
rect 4592 1244 4596 1287
rect 4614 1264 4618 1301
rect 4634 1299 4641 1336
rect 4671 1319 4675 1396
rect 4666 1307 4675 1319
rect 4669 1291 4675 1307
rect 4691 1319 4695 1396
rect 4691 1307 4694 1319
rect 4691 1291 4697 1307
rect 4634 1274 4641 1287
rect 4669 1284 4677 1291
rect 4622 1268 4641 1274
rect 4622 1264 4626 1268
rect 4673 1264 4677 1284
rect 4683 1284 4697 1291
rect 4683 1264 4687 1284
rect 31 1220 35 1224
rect 53 1220 57 1224
rect 63 1220 67 1224
rect 83 1220 87 1224
rect 91 1220 95 1224
rect 137 1220 141 1224
rect 159 1220 163 1224
rect 169 1220 173 1224
rect 191 1220 195 1224
rect 201 1220 205 1224
rect 221 1220 225 1224
rect 275 1220 279 1224
rect 295 1220 299 1224
rect 305 1220 309 1224
rect 327 1220 331 1224
rect 337 1220 341 1224
rect 359 1220 363 1224
rect 405 1220 409 1224
rect 413 1220 417 1224
rect 433 1220 437 1224
rect 443 1220 447 1224
rect 465 1220 469 1224
rect 513 1220 517 1224
rect 523 1220 527 1224
rect 605 1220 609 1224
rect 625 1220 629 1224
rect 645 1220 649 1224
rect 705 1220 709 1224
rect 725 1220 729 1224
rect 745 1220 749 1224
rect 803 1220 807 1224
rect 825 1220 829 1224
rect 873 1220 877 1224
rect 883 1220 887 1224
rect 965 1220 969 1224
rect 985 1220 989 1224
rect 1005 1220 1009 1224
rect 1065 1220 1069 1224
rect 1111 1220 1115 1224
rect 1131 1220 1135 1224
rect 1151 1220 1155 1224
rect 1171 1220 1175 1224
rect 1253 1220 1257 1224
rect 1263 1220 1267 1224
rect 1325 1220 1329 1224
rect 1345 1220 1349 1224
rect 1365 1220 1369 1224
rect 1433 1220 1437 1224
rect 1443 1220 1447 1224
rect 1505 1220 1509 1224
rect 1525 1220 1529 1224
rect 1545 1220 1549 1224
rect 1591 1220 1595 1224
rect 1613 1220 1617 1224
rect 1673 1220 1677 1224
rect 1683 1220 1687 1224
rect 1765 1220 1769 1224
rect 1785 1220 1789 1224
rect 1805 1220 1809 1224
rect 1851 1220 1855 1224
rect 1873 1220 1877 1224
rect 1883 1220 1887 1224
rect 1903 1220 1907 1224
rect 1911 1220 1915 1224
rect 1957 1220 1961 1224
rect 1979 1220 1983 1224
rect 1989 1220 1993 1224
rect 2011 1220 2015 1224
rect 2021 1220 2025 1224
rect 2041 1220 2045 1224
rect 2091 1220 2095 1224
rect 2151 1220 2155 1224
rect 2171 1220 2175 1224
rect 2191 1220 2195 1224
rect 2273 1220 2277 1224
rect 2283 1220 2287 1224
rect 2345 1220 2349 1224
rect 2365 1220 2369 1224
rect 2425 1220 2429 1224
rect 2471 1220 2475 1224
rect 2491 1220 2495 1224
rect 2551 1220 2555 1224
rect 2573 1220 2577 1224
rect 2583 1220 2587 1224
rect 2603 1220 2607 1224
rect 2611 1220 2615 1224
rect 2657 1220 2661 1224
rect 2679 1220 2683 1224
rect 2689 1220 2693 1224
rect 2711 1220 2715 1224
rect 2721 1220 2725 1224
rect 2741 1220 2745 1224
rect 2791 1220 2795 1224
rect 2811 1220 2815 1224
rect 2885 1220 2889 1224
rect 2931 1220 2935 1224
rect 2951 1220 2955 1224
rect 2971 1220 2975 1224
rect 3031 1220 3035 1224
rect 3051 1220 3055 1224
rect 3071 1220 3075 1224
rect 3131 1220 3135 1224
rect 3151 1220 3155 1224
rect 3171 1220 3175 1224
rect 3231 1220 3235 1224
rect 3241 1220 3245 1224
rect 3261 1220 3265 1224
rect 3345 1220 3349 1224
rect 3365 1220 3369 1224
rect 3412 1220 3416 1224
rect 3420 1220 3424 1224
rect 3428 1220 3432 1224
rect 3525 1220 3529 1224
rect 3545 1220 3549 1224
rect 3565 1220 3569 1224
rect 3611 1220 3615 1224
rect 3631 1220 3635 1224
rect 3651 1220 3655 1224
rect 3733 1220 3737 1224
rect 3743 1220 3747 1224
rect 3813 1220 3817 1224
rect 3823 1220 3827 1224
rect 3871 1220 3875 1224
rect 3881 1220 3885 1224
rect 3901 1220 3905 1224
rect 3985 1220 3989 1224
rect 4005 1220 4009 1224
rect 4025 1220 4029 1224
rect 4071 1220 4075 1224
rect 4153 1220 4157 1224
rect 4163 1220 4167 1224
rect 4233 1220 4237 1224
rect 4243 1220 4247 1224
rect 4305 1220 4309 1224
rect 4325 1220 4329 1224
rect 4385 1220 4389 1224
rect 4405 1220 4409 1224
rect 4425 1220 4429 1224
rect 4471 1220 4475 1224
rect 4491 1220 4495 1224
rect 4511 1220 4515 1224
rect 4592 1220 4596 1224
rect 4614 1220 4618 1224
rect 4622 1220 4626 1224
rect 4673 1220 4677 1224
rect 4683 1220 4687 1224
rect 31 1196 35 1200
rect 113 1196 117 1200
rect 123 1196 127 1200
rect 185 1196 189 1200
rect 205 1196 209 1200
rect 225 1196 229 1200
rect 274 1196 278 1200
rect 282 1196 286 1200
rect 302 1196 306 1200
rect 310 1196 314 1200
rect 412 1196 416 1200
rect 434 1196 438 1200
rect 442 1196 446 1200
rect 505 1196 509 1200
rect 525 1196 529 1200
rect 545 1196 549 1200
rect 591 1196 595 1200
rect 611 1196 615 1200
rect 695 1196 699 1200
rect 715 1196 719 1200
rect 725 1196 729 1200
rect 783 1196 787 1200
rect 805 1196 809 1200
rect 865 1196 869 1200
rect 885 1196 889 1200
rect 945 1196 949 1200
rect 1005 1196 1009 1200
rect 1051 1196 1055 1200
rect 1071 1196 1075 1200
rect 1131 1196 1135 1200
rect 1205 1196 1209 1200
rect 1225 1196 1229 1200
rect 1274 1196 1278 1200
rect 1282 1196 1286 1200
rect 1304 1196 1308 1200
rect 1375 1196 1379 1200
rect 1395 1196 1399 1200
rect 1405 1196 1409 1200
rect 1427 1196 1431 1200
rect 1437 1196 1441 1200
rect 1459 1196 1463 1200
rect 1505 1196 1509 1200
rect 1513 1196 1517 1200
rect 1533 1196 1537 1200
rect 1543 1196 1547 1200
rect 1565 1196 1569 1200
rect 1625 1196 1629 1200
rect 1673 1196 1677 1200
rect 1683 1196 1687 1200
rect 1751 1196 1755 1200
rect 1771 1196 1775 1200
rect 1835 1196 1839 1200
rect 1855 1196 1859 1200
rect 1865 1196 1869 1200
rect 1887 1196 1891 1200
rect 1897 1196 1901 1200
rect 1919 1196 1923 1200
rect 1965 1196 1969 1200
rect 1973 1196 1977 1200
rect 1993 1196 1997 1200
rect 2003 1196 2007 1200
rect 2025 1196 2029 1200
rect 2085 1196 2089 1200
rect 2131 1196 2135 1200
rect 2151 1196 2155 1200
rect 2211 1196 2215 1200
rect 2231 1196 2235 1200
rect 2305 1196 2309 1200
rect 2351 1196 2355 1200
rect 2373 1196 2377 1200
rect 2383 1196 2387 1200
rect 2403 1196 2407 1200
rect 2411 1196 2415 1200
rect 2457 1196 2461 1200
rect 2479 1196 2483 1200
rect 2489 1196 2493 1200
rect 2511 1196 2515 1200
rect 2521 1196 2525 1200
rect 2541 1196 2545 1200
rect 2591 1196 2595 1200
rect 2651 1196 2655 1200
rect 2671 1196 2675 1200
rect 2691 1196 2695 1200
rect 2751 1196 2755 1200
rect 2771 1196 2775 1200
rect 2791 1196 2795 1200
rect 2811 1196 2815 1200
rect 2871 1196 2875 1200
rect 2891 1196 2895 1200
rect 2973 1196 2977 1200
rect 2983 1196 2987 1200
rect 3031 1196 3035 1200
rect 3041 1196 3045 1200
rect 3061 1196 3065 1200
rect 3131 1196 3135 1200
rect 3151 1196 3155 1200
rect 3171 1196 3175 1200
rect 3231 1196 3235 1200
rect 3251 1196 3255 1200
rect 3271 1196 3275 1200
rect 3353 1196 3357 1200
rect 3363 1196 3367 1200
rect 3433 1196 3437 1200
rect 3443 1196 3447 1200
rect 3493 1196 3497 1200
rect 3503 1196 3507 1200
rect 3573 1196 3577 1200
rect 3583 1196 3587 1200
rect 3651 1196 3655 1200
rect 3671 1196 3675 1200
rect 3691 1196 3695 1200
rect 3788 1196 3792 1200
rect 3796 1196 3800 1200
rect 3804 1196 3808 1200
rect 3854 1196 3858 1200
rect 3862 1196 3866 1200
rect 3884 1196 3888 1200
rect 3965 1196 3969 1200
rect 4048 1196 4052 1200
rect 4056 1196 4060 1200
rect 4064 1196 4068 1200
rect 4114 1196 4118 1200
rect 4122 1196 4126 1200
rect 4144 1196 4148 1200
rect 4211 1196 4215 1200
rect 4292 1196 4296 1200
rect 4314 1196 4318 1200
rect 4322 1196 4326 1200
rect 4385 1196 4389 1200
rect 4405 1196 4409 1200
rect 4425 1196 4429 1200
rect 4471 1196 4475 1200
rect 4491 1196 4495 1200
rect 4511 1196 4515 1200
rect 4571 1196 4575 1200
rect 4591 1196 4595 1200
rect 4673 1196 4677 1200
rect 4683 1196 4687 1200
rect 4745 1196 4749 1200
rect 31 1119 35 1176
rect 113 1136 117 1156
rect 26 1107 35 1119
rect 103 1129 117 1136
rect 123 1136 127 1156
rect 123 1129 131 1136
rect 103 1113 109 1129
rect 31 1024 35 1107
rect 106 1101 109 1113
rect 105 1024 109 1101
rect 125 1113 131 1129
rect 125 1101 134 1113
rect 125 1024 129 1101
rect 185 1079 189 1156
rect 205 1133 209 1156
rect 225 1151 229 1156
rect 225 1144 238 1151
rect 274 1148 278 1156
rect 205 1121 214 1133
rect 187 1067 194 1079
rect 190 1024 194 1067
rect 212 1064 216 1121
rect 234 1099 238 1144
rect 261 1141 278 1148
rect 261 1099 267 1141
rect 282 1133 286 1156
rect 302 1142 306 1156
rect 310 1151 314 1156
rect 310 1147 340 1151
rect 302 1135 315 1142
rect 311 1133 315 1135
rect 311 1121 313 1133
rect 282 1092 286 1121
rect 267 1087 275 1092
rect 234 1076 238 1087
rect 255 1086 275 1087
rect 282 1086 295 1092
rect 220 1068 238 1076
rect 220 1064 224 1068
rect 271 1064 275 1086
rect 291 1064 295 1086
rect 311 1064 315 1121
rect 334 1099 340 1147
rect 412 1133 416 1176
rect 525 1169 529 1176
rect 545 1169 549 1176
rect 525 1163 539 1169
rect 545 1164 558 1169
rect 405 1121 414 1133
rect 331 1087 334 1099
rect 331 1064 335 1087
rect 405 1064 409 1121
rect 434 1119 438 1156
rect 442 1152 446 1156
rect 442 1146 461 1152
rect 454 1133 461 1146
rect 505 1148 509 1156
rect 505 1136 515 1148
rect 434 1084 440 1107
rect 454 1084 461 1121
rect 535 1099 539 1163
rect 554 1119 558 1164
rect 425 1078 440 1084
rect 445 1078 461 1084
rect 425 1064 429 1078
rect 445 1064 449 1078
rect 515 1064 519 1069
rect 535 1064 539 1087
rect 554 1073 558 1107
rect 591 1099 595 1176
rect 611 1099 615 1176
rect 695 1150 699 1156
rect 681 1138 693 1150
rect 586 1087 595 1099
rect 545 1068 558 1073
rect 545 1064 549 1068
rect 591 1064 595 1087
rect 599 1087 614 1099
rect 599 1064 603 1087
rect 681 1064 685 1138
rect 715 1113 719 1156
rect 706 1101 719 1113
rect 703 1024 707 1101
rect 725 1099 729 1156
rect 783 1150 787 1156
rect 783 1138 785 1150
rect 805 1099 809 1176
rect 865 1099 869 1176
rect 885 1099 889 1176
rect 945 1119 949 1176
rect 1005 1119 1009 1176
rect 945 1107 954 1119
rect 1005 1107 1014 1119
rect 725 1087 734 1099
rect 805 1087 814 1099
rect 866 1087 881 1099
rect 725 1024 729 1087
rect 783 1070 785 1082
rect 783 1064 787 1070
rect 805 1024 809 1087
rect 877 1064 881 1087
rect 885 1087 894 1099
rect 885 1064 889 1087
rect 945 1024 949 1107
rect 1005 1024 1009 1107
rect 1051 1099 1055 1176
rect 1071 1099 1075 1176
rect 1131 1119 1135 1176
rect 1126 1107 1135 1119
rect 1046 1087 1055 1099
rect 1051 1064 1055 1087
rect 1059 1087 1074 1099
rect 1059 1064 1063 1087
rect 1131 1024 1135 1107
rect 1205 1099 1209 1176
rect 1225 1099 1229 1176
rect 1274 1152 1278 1156
rect 1259 1146 1278 1152
rect 1259 1133 1266 1146
rect 1206 1087 1221 1099
rect 1217 1064 1221 1087
rect 1225 1087 1234 1099
rect 1225 1064 1229 1087
rect 1259 1084 1266 1121
rect 1282 1119 1286 1156
rect 1304 1133 1308 1176
rect 1306 1121 1315 1133
rect 1280 1084 1286 1107
rect 1259 1078 1275 1084
rect 1280 1078 1295 1084
rect 1271 1064 1275 1078
rect 1291 1064 1295 1078
rect 1311 1064 1315 1121
rect 1375 1119 1379 1156
rect 1395 1118 1399 1176
rect 1405 1144 1409 1176
rect 1427 1164 1431 1176
rect 1429 1152 1431 1164
rect 1437 1164 1441 1176
rect 1437 1152 1439 1164
rect 1405 1140 1438 1144
rect 1375 1064 1379 1107
rect 1395 1024 1399 1106
rect 1414 1091 1418 1120
rect 1409 1083 1418 1091
rect 1409 1024 1413 1083
rect 1434 1076 1438 1140
rect 1435 1064 1438 1076
rect 1429 1024 1433 1064
rect 1443 1042 1447 1152
rect 1459 1062 1463 1176
rect 1505 1172 1509 1176
rect 1475 1168 1509 1172
rect 1441 1024 1445 1030
rect 1461 1024 1465 1050
rect 1475 1042 1479 1168
rect 1513 1164 1517 1176
rect 1487 1160 1517 1164
rect 1499 1159 1517 1160
rect 1533 1155 1537 1176
rect 1513 1151 1537 1155
rect 1513 1056 1519 1151
rect 1543 1127 1547 1176
rect 1543 1069 1547 1115
rect 1565 1088 1569 1156
rect 1567 1076 1569 1088
rect 1543 1063 1551 1069
rect 1565 1064 1569 1076
rect 1625 1119 1629 1176
rect 1673 1136 1677 1156
rect 1669 1129 1677 1136
rect 1683 1136 1687 1156
rect 1683 1129 1697 1136
rect 1625 1107 1634 1119
rect 1669 1113 1675 1129
rect 1487 1030 1511 1032
rect 1475 1028 1511 1030
rect 1507 1024 1511 1028
rect 1515 1024 1519 1056
rect 1535 1004 1539 1044
rect 1547 1034 1551 1063
rect 1543 1027 1551 1034
rect 1543 1004 1547 1027
rect 1625 1024 1629 1107
rect 1666 1101 1675 1113
rect 1671 1024 1675 1101
rect 1691 1113 1697 1129
rect 1691 1101 1694 1113
rect 1691 1024 1695 1101
rect 1751 1099 1755 1176
rect 1771 1099 1775 1176
rect 1835 1119 1839 1156
rect 1855 1118 1859 1176
rect 1865 1144 1869 1176
rect 1887 1164 1891 1176
rect 1889 1152 1891 1164
rect 1897 1164 1901 1176
rect 1897 1152 1899 1164
rect 1865 1140 1898 1144
rect 1746 1087 1755 1099
rect 1751 1064 1755 1087
rect 1759 1087 1774 1099
rect 1759 1064 1763 1087
rect 1835 1064 1839 1107
rect 1855 1024 1859 1106
rect 1874 1091 1878 1120
rect 1869 1083 1878 1091
rect 1869 1024 1873 1083
rect 1894 1076 1898 1140
rect 1895 1064 1898 1076
rect 1889 1024 1893 1064
rect 1903 1042 1907 1152
rect 1919 1062 1923 1176
rect 1965 1172 1969 1176
rect 1935 1168 1969 1172
rect 1901 1024 1905 1030
rect 1921 1024 1925 1050
rect 1935 1042 1939 1168
rect 1973 1164 1977 1176
rect 1947 1160 1977 1164
rect 1959 1159 1977 1160
rect 1993 1155 1997 1176
rect 1973 1151 1997 1155
rect 1973 1056 1979 1151
rect 2003 1127 2007 1176
rect 2003 1069 2007 1115
rect 2025 1088 2029 1156
rect 2027 1076 2029 1088
rect 2003 1063 2011 1069
rect 2025 1064 2029 1076
rect 2085 1119 2089 1176
rect 2085 1107 2094 1119
rect 1947 1030 1971 1032
rect 1935 1028 1971 1030
rect 1967 1024 1971 1028
rect 1975 1024 1979 1056
rect 1995 1004 1999 1044
rect 2007 1034 2011 1063
rect 2003 1027 2011 1034
rect 2003 1004 2007 1027
rect 2085 1024 2089 1107
rect 2131 1099 2135 1176
rect 2151 1099 2155 1176
rect 2211 1099 2215 1176
rect 2231 1099 2235 1176
rect 2305 1119 2309 1176
rect 2305 1107 2314 1119
rect 2126 1087 2135 1099
rect 2131 1064 2135 1087
rect 2139 1087 2154 1099
rect 2206 1087 2215 1099
rect 2139 1064 2143 1087
rect 2211 1064 2215 1087
rect 2219 1087 2234 1099
rect 2219 1064 2223 1087
rect 2305 1024 2309 1107
rect 2351 1088 2355 1156
rect 2373 1127 2377 1176
rect 2383 1155 2387 1176
rect 2403 1164 2407 1176
rect 2411 1172 2415 1176
rect 2411 1168 2445 1172
rect 2403 1160 2433 1164
rect 2403 1159 2421 1160
rect 2383 1151 2407 1155
rect 2351 1076 2353 1088
rect 2351 1064 2355 1076
rect 2373 1069 2377 1115
rect 2369 1063 2377 1069
rect 2369 1034 2373 1063
rect 2401 1056 2407 1151
rect 2369 1027 2377 1034
rect 2373 1004 2377 1027
rect 2381 1004 2385 1044
rect 2401 1024 2405 1056
rect 2441 1042 2445 1168
rect 2457 1062 2461 1176
rect 2479 1164 2483 1176
rect 2481 1152 2483 1164
rect 2489 1164 2493 1176
rect 2489 1152 2491 1164
rect 2409 1030 2433 1032
rect 2409 1028 2445 1030
rect 2409 1024 2413 1028
rect 2455 1024 2459 1050
rect 2473 1042 2477 1152
rect 2511 1144 2515 1176
rect 2482 1140 2515 1144
rect 2482 1076 2486 1140
rect 2502 1091 2506 1120
rect 2521 1118 2525 1176
rect 2541 1119 2545 1156
rect 2591 1119 2595 1176
rect 2651 1151 2655 1156
rect 2586 1107 2595 1119
rect 2502 1083 2511 1091
rect 2482 1064 2485 1076
rect 2475 1024 2479 1030
rect 2487 1024 2491 1064
rect 2507 1024 2511 1083
rect 2521 1024 2525 1106
rect 2541 1064 2545 1107
rect 2591 1024 2595 1107
rect 2642 1144 2655 1151
rect 2642 1099 2646 1144
rect 2671 1133 2675 1156
rect 2666 1121 2675 1133
rect 2642 1076 2646 1087
rect 2642 1068 2660 1076
rect 2656 1064 2660 1068
rect 2664 1064 2668 1121
rect 2691 1079 2695 1156
rect 2751 1149 2755 1156
rect 2740 1145 2755 1149
rect 2740 1099 2746 1145
rect 2771 1133 2775 1156
rect 2791 1133 2795 1156
rect 2766 1121 2775 1133
rect 2686 1067 2693 1079
rect 2741 1072 2746 1087
rect 2769 1072 2775 1121
rect 2741 1068 2755 1072
rect 2686 1024 2690 1067
rect 2751 1064 2755 1068
rect 2761 1068 2775 1072
rect 2761 1064 2765 1068
rect 2791 1064 2795 1121
rect 2811 1099 2815 1156
rect 2871 1099 2875 1176
rect 2891 1099 2895 1176
rect 3231 1169 3235 1176
rect 3251 1169 3255 1176
rect 3222 1164 3235 1169
rect 2973 1136 2977 1156
rect 2963 1129 2977 1136
rect 2983 1136 2987 1156
rect 2983 1129 2991 1136
rect 2963 1113 2969 1129
rect 2966 1101 2969 1113
rect 2811 1087 2813 1099
rect 2866 1087 2875 1099
rect 2811 1072 2815 1087
rect 2801 1068 2815 1072
rect 2801 1064 2805 1068
rect 2871 1064 2875 1087
rect 2879 1087 2894 1099
rect 2879 1064 2883 1087
rect 2965 1024 2969 1101
rect 2985 1113 2991 1129
rect 2985 1101 2994 1113
rect 2985 1024 2989 1101
rect 3031 1099 3035 1156
rect 3041 1113 3045 1156
rect 3061 1150 3065 1156
rect 3131 1151 3135 1156
rect 3067 1138 3079 1150
rect 3041 1101 3054 1113
rect 3026 1087 3035 1099
rect 3031 1024 3035 1087
rect 3053 1024 3057 1101
rect 3075 1064 3079 1138
rect 3122 1144 3135 1151
rect 3122 1099 3126 1144
rect 3151 1133 3155 1156
rect 3146 1121 3155 1133
rect 3122 1076 3126 1087
rect 3122 1068 3140 1076
rect 3136 1064 3140 1068
rect 3144 1064 3148 1121
rect 3171 1079 3175 1156
rect 3222 1119 3226 1164
rect 3166 1067 3173 1079
rect 3222 1073 3226 1107
rect 3241 1163 3255 1169
rect 3241 1099 3245 1163
rect 3271 1148 3275 1156
rect 3265 1136 3275 1148
rect 3353 1136 3357 1156
rect 3343 1129 3357 1136
rect 3363 1136 3367 1156
rect 3433 1136 3437 1156
rect 3363 1129 3371 1136
rect 3343 1113 3349 1129
rect 3346 1101 3349 1113
rect 3222 1068 3235 1073
rect 3166 1024 3170 1067
rect 3231 1064 3235 1068
rect 3241 1064 3245 1087
rect 3261 1064 3265 1069
rect 3345 1024 3349 1101
rect 3365 1113 3371 1129
rect 3423 1129 3437 1136
rect 3443 1136 3447 1156
rect 3493 1136 3497 1156
rect 3443 1129 3451 1136
rect 3423 1113 3429 1129
rect 3365 1101 3374 1113
rect 3426 1101 3429 1113
rect 3365 1024 3369 1101
rect 3425 1024 3429 1101
rect 3445 1113 3451 1129
rect 3489 1129 3497 1136
rect 3503 1136 3507 1156
rect 3573 1136 3577 1156
rect 3503 1129 3517 1136
rect 3489 1113 3495 1129
rect 3445 1101 3454 1113
rect 3486 1101 3495 1113
rect 3445 1024 3449 1101
rect 3491 1024 3495 1101
rect 3511 1113 3517 1129
rect 3569 1129 3577 1136
rect 3583 1136 3587 1156
rect 3651 1151 3655 1156
rect 3642 1144 3655 1151
rect 3583 1129 3597 1136
rect 3569 1113 3575 1129
rect 3511 1101 3514 1113
rect 3566 1101 3575 1113
rect 3511 1024 3515 1101
rect 3571 1024 3575 1101
rect 3591 1113 3597 1129
rect 3591 1101 3594 1113
rect 3591 1024 3595 1101
rect 3642 1099 3646 1144
rect 3671 1133 3675 1156
rect 3666 1121 3675 1133
rect 3642 1076 3646 1087
rect 3642 1068 3660 1076
rect 3656 1064 3660 1068
rect 3664 1064 3668 1121
rect 3691 1079 3695 1156
rect 3854 1152 3858 1156
rect 3839 1146 3858 1152
rect 3788 1079 3792 1136
rect 3686 1067 3693 1079
rect 3765 1067 3773 1079
rect 3785 1067 3792 1079
rect 3686 1024 3690 1067
rect 3765 1024 3769 1067
rect 3796 1059 3800 1136
rect 3804 1079 3808 1136
rect 3839 1133 3846 1146
rect 3839 1084 3846 1121
rect 3862 1119 3866 1156
rect 3884 1133 3888 1176
rect 3886 1121 3895 1133
rect 3860 1084 3866 1107
rect 3804 1067 3814 1079
rect 3839 1078 3855 1084
rect 3860 1078 3875 1084
rect 3794 1040 3800 1047
rect 3785 1036 3800 1040
rect 3814 1036 3820 1067
rect 3851 1064 3855 1078
rect 3871 1064 3875 1078
rect 3891 1064 3895 1121
rect 3965 1119 3969 1176
rect 4114 1152 4118 1156
rect 4099 1146 4118 1152
rect 3965 1107 3974 1119
rect 3785 1024 3789 1036
rect 3805 1032 3820 1036
rect 3805 1024 3809 1032
rect 3965 1024 3969 1107
rect 4048 1079 4052 1136
rect 4025 1067 4033 1079
rect 4045 1067 4052 1079
rect 4025 1024 4029 1067
rect 4056 1059 4060 1136
rect 4064 1079 4068 1136
rect 4099 1133 4106 1146
rect 4099 1084 4106 1121
rect 4122 1119 4126 1156
rect 4144 1133 4148 1176
rect 4146 1121 4155 1133
rect 4120 1084 4126 1107
rect 4064 1067 4074 1079
rect 4099 1078 4115 1084
rect 4120 1078 4135 1084
rect 4054 1040 4060 1047
rect 4045 1036 4060 1040
rect 4074 1036 4080 1067
rect 4111 1064 4115 1078
rect 4131 1064 4135 1078
rect 4151 1064 4155 1121
rect 4211 1119 4215 1176
rect 4292 1133 4296 1176
rect 4206 1107 4215 1119
rect 4045 1024 4049 1036
rect 4065 1032 4080 1036
rect 4065 1024 4069 1032
rect 4211 1024 4215 1107
rect 4285 1121 4294 1133
rect 4285 1064 4289 1121
rect 4314 1119 4318 1156
rect 4322 1152 4326 1156
rect 4322 1146 4341 1152
rect 4334 1133 4341 1146
rect 4314 1084 4320 1107
rect 4334 1084 4341 1121
rect 4305 1078 4320 1084
rect 4325 1078 4341 1084
rect 4385 1079 4389 1156
rect 4405 1133 4409 1156
rect 4425 1151 4429 1156
rect 4471 1151 4475 1156
rect 4425 1144 4438 1151
rect 4405 1121 4414 1133
rect 4305 1064 4309 1078
rect 4325 1064 4329 1078
rect 4387 1067 4394 1079
rect 4390 1024 4394 1067
rect 4412 1064 4416 1121
rect 4434 1099 4438 1144
rect 4462 1144 4475 1151
rect 4462 1099 4466 1144
rect 4491 1133 4495 1156
rect 4486 1121 4495 1133
rect 4434 1076 4438 1087
rect 4420 1068 4438 1076
rect 4462 1076 4466 1087
rect 4462 1068 4480 1076
rect 4420 1064 4424 1068
rect 4476 1064 4480 1068
rect 4484 1064 4488 1121
rect 4511 1079 4515 1156
rect 4571 1099 4575 1176
rect 4591 1099 4595 1176
rect 4673 1136 4677 1156
rect 4663 1129 4677 1136
rect 4683 1136 4687 1156
rect 4683 1129 4691 1136
rect 4663 1113 4669 1129
rect 4666 1101 4669 1113
rect 4566 1087 4575 1099
rect 4506 1067 4513 1079
rect 4506 1024 4510 1067
rect 4571 1064 4575 1087
rect 4579 1087 4594 1099
rect 4579 1064 4583 1087
rect 4665 1024 4669 1101
rect 4685 1113 4691 1129
rect 4745 1119 4749 1176
rect 4685 1101 4694 1113
rect 4745 1107 4754 1119
rect 4685 1024 4689 1101
rect 4745 1024 4749 1107
rect 31 980 35 984
rect 105 980 109 984
rect 125 980 129 984
rect 190 980 194 984
rect 212 980 216 984
rect 220 980 224 984
rect 271 980 275 984
rect 291 980 295 984
rect 311 980 315 984
rect 331 980 335 984
rect 405 980 409 984
rect 425 980 429 984
rect 445 980 449 984
rect 515 980 519 984
rect 535 980 539 984
rect 545 980 549 984
rect 591 980 595 984
rect 599 980 603 984
rect 681 980 685 984
rect 703 980 707 984
rect 725 980 729 984
rect 783 980 787 984
rect 805 980 809 984
rect 877 980 881 984
rect 885 980 889 984
rect 945 980 949 984
rect 1005 980 1009 984
rect 1051 980 1055 984
rect 1059 980 1063 984
rect 1131 980 1135 984
rect 1217 980 1221 984
rect 1225 980 1229 984
rect 1271 980 1275 984
rect 1291 980 1295 984
rect 1311 980 1315 984
rect 1375 980 1379 984
rect 1395 980 1399 984
rect 1409 980 1413 984
rect 1429 980 1433 984
rect 1441 980 1445 984
rect 1461 980 1465 984
rect 1507 980 1511 984
rect 1515 980 1519 984
rect 1535 980 1539 984
rect 1543 980 1547 984
rect 1565 980 1569 984
rect 1625 980 1629 984
rect 1671 980 1675 984
rect 1691 980 1695 984
rect 1751 980 1755 984
rect 1759 980 1763 984
rect 1835 980 1839 984
rect 1855 980 1859 984
rect 1869 980 1873 984
rect 1889 980 1893 984
rect 1901 980 1905 984
rect 1921 980 1925 984
rect 1967 980 1971 984
rect 1975 980 1979 984
rect 1995 980 1999 984
rect 2003 980 2007 984
rect 2025 980 2029 984
rect 2085 980 2089 984
rect 2131 980 2135 984
rect 2139 980 2143 984
rect 2211 980 2215 984
rect 2219 980 2223 984
rect 2305 980 2309 984
rect 2351 980 2355 984
rect 2373 980 2377 984
rect 2381 980 2385 984
rect 2401 980 2405 984
rect 2409 980 2413 984
rect 2455 980 2459 984
rect 2475 980 2479 984
rect 2487 980 2491 984
rect 2507 980 2511 984
rect 2521 980 2525 984
rect 2541 980 2545 984
rect 2591 980 2595 984
rect 2656 980 2660 984
rect 2664 980 2668 984
rect 2686 980 2690 984
rect 2751 980 2755 984
rect 2761 980 2765 984
rect 2791 980 2795 984
rect 2801 980 2805 984
rect 2871 980 2875 984
rect 2879 980 2883 984
rect 2965 980 2969 984
rect 2985 980 2989 984
rect 3031 980 3035 984
rect 3053 980 3057 984
rect 3075 980 3079 984
rect 3136 980 3140 984
rect 3144 980 3148 984
rect 3166 980 3170 984
rect 3231 980 3235 984
rect 3241 980 3245 984
rect 3261 980 3265 984
rect 3345 980 3349 984
rect 3365 980 3369 984
rect 3425 980 3429 984
rect 3445 980 3449 984
rect 3491 980 3495 984
rect 3511 980 3515 984
rect 3571 980 3575 984
rect 3591 980 3595 984
rect 3656 980 3660 984
rect 3664 980 3668 984
rect 3686 980 3690 984
rect 3765 980 3769 984
rect 3785 980 3789 984
rect 3805 980 3809 984
rect 3851 980 3855 984
rect 3871 980 3875 984
rect 3891 980 3895 984
rect 3965 980 3969 984
rect 4025 980 4029 984
rect 4045 980 4049 984
rect 4065 980 4069 984
rect 4111 980 4115 984
rect 4131 980 4135 984
rect 4151 980 4155 984
rect 4211 980 4215 984
rect 4285 980 4289 984
rect 4305 980 4309 984
rect 4325 980 4329 984
rect 4390 980 4394 984
rect 4412 980 4416 984
rect 4420 980 4424 984
rect 4476 980 4480 984
rect 4484 980 4488 984
rect 4506 980 4510 984
rect 4571 980 4575 984
rect 4579 980 4583 984
rect 4665 980 4669 984
rect 4685 980 4689 984
rect 4745 980 4749 984
rect 35 956 39 960
rect 55 956 59 960
rect 69 956 73 960
rect 89 956 93 960
rect 101 956 105 960
rect 121 956 125 960
rect 167 956 171 960
rect 175 956 179 960
rect 195 956 199 960
rect 203 956 207 960
rect 225 956 229 960
rect 271 956 275 960
rect 291 956 295 960
rect 370 956 374 960
rect 392 956 396 960
rect 400 956 404 960
rect 455 956 459 960
rect 475 956 479 960
rect 489 956 493 960
rect 509 956 513 960
rect 521 956 525 960
rect 541 956 545 960
rect 587 956 591 960
rect 595 956 599 960
rect 615 956 619 960
rect 623 956 627 960
rect 645 956 649 960
rect 691 956 695 960
rect 711 956 715 960
rect 790 956 794 960
rect 812 956 816 960
rect 820 956 824 960
rect 890 956 894 960
rect 912 956 916 960
rect 920 956 924 960
rect 985 956 989 960
rect 1057 956 1061 960
rect 1065 956 1069 960
rect 1111 956 1115 960
rect 1119 956 1123 960
rect 1205 956 1209 960
rect 1225 956 1229 960
rect 1285 956 1289 960
rect 1305 956 1309 960
rect 1365 956 1369 960
rect 1385 956 1389 960
rect 1445 956 1449 960
rect 1465 956 1469 960
rect 1485 956 1489 960
rect 1541 956 1545 960
rect 1563 956 1567 960
rect 1585 956 1589 960
rect 1631 956 1635 960
rect 1651 956 1655 960
rect 1671 956 1675 960
rect 1731 956 1735 960
rect 1751 956 1755 960
rect 1771 956 1775 960
rect 1791 956 1795 960
rect 1811 956 1815 960
rect 1831 956 1835 960
rect 1851 956 1855 960
rect 1871 956 1875 960
rect 1945 956 1949 960
rect 1965 956 1969 960
rect 2037 956 2041 960
rect 2045 956 2049 960
rect 2096 956 2100 960
rect 2104 956 2108 960
rect 2126 956 2130 960
rect 2196 956 2200 960
rect 2204 956 2208 960
rect 2226 956 2230 960
rect 2296 956 2300 960
rect 2304 956 2308 960
rect 2326 956 2330 960
rect 2391 956 2395 960
rect 2411 956 2415 960
rect 2485 956 2489 960
rect 2531 956 2535 960
rect 2553 956 2557 960
rect 2561 956 2565 960
rect 2581 956 2585 960
rect 2589 956 2593 960
rect 2635 956 2639 960
rect 2655 956 2659 960
rect 2667 956 2671 960
rect 2687 956 2691 960
rect 2701 956 2705 960
rect 2721 956 2725 960
rect 2790 956 2794 960
rect 2812 956 2816 960
rect 2820 956 2824 960
rect 2885 956 2889 960
rect 2931 956 2935 960
rect 2991 956 2995 960
rect 3011 956 3015 960
rect 3031 956 3035 960
rect 3091 956 3095 960
rect 3165 956 3169 960
rect 3185 956 3189 960
rect 3231 956 3235 960
rect 3241 956 3245 960
rect 3261 956 3265 960
rect 3331 956 3335 960
rect 3351 956 3355 960
rect 3411 956 3415 960
rect 3431 956 3435 960
rect 3517 956 3521 960
rect 3525 956 3529 960
rect 3571 956 3575 960
rect 3591 956 3595 960
rect 3665 956 3669 960
rect 3685 956 3689 960
rect 3705 956 3709 960
rect 3765 956 3769 960
rect 3785 956 3789 960
rect 3805 956 3809 960
rect 3851 956 3855 960
rect 3871 956 3875 960
rect 3945 956 3949 960
rect 3965 956 3969 960
rect 3985 956 3989 960
rect 4045 956 4049 960
rect 4110 956 4114 960
rect 4132 956 4136 960
rect 4140 956 4144 960
rect 4210 956 4214 960
rect 4232 956 4236 960
rect 4240 956 4244 960
rect 4305 956 4309 960
rect 4325 956 4329 960
rect 4345 956 4349 960
rect 4391 956 4395 960
rect 4411 956 4415 960
rect 4431 956 4435 960
rect 4505 956 4509 960
rect 4525 956 4529 960
rect 4545 956 4549 960
rect 4605 956 4609 960
rect 4625 956 4629 960
rect 4645 956 4649 960
rect 4691 956 4695 960
rect 4711 956 4715 960
rect 4731 956 4735 960
rect 35 833 39 876
rect 55 834 59 916
rect 69 857 73 916
rect 89 876 93 916
rect 101 910 105 916
rect 95 864 98 876
rect 69 849 78 857
rect 35 784 39 821
rect 55 764 59 822
rect 74 820 78 849
rect 94 800 98 864
rect 65 796 98 800
rect 65 764 69 796
rect 103 788 107 898
rect 121 890 125 916
rect 167 912 171 916
rect 135 910 171 912
rect 147 908 171 910
rect 89 776 91 788
rect 87 764 91 776
rect 97 776 99 788
rect 97 764 101 776
rect 119 764 123 878
rect 135 772 139 898
rect 175 884 179 916
rect 195 896 199 936
rect 203 913 207 936
rect 203 906 211 913
rect 173 789 179 884
rect 207 877 211 906
rect 203 871 211 877
rect 203 825 207 871
rect 225 864 229 876
rect 227 852 229 864
rect 173 785 197 789
rect 159 780 177 781
rect 147 776 177 780
rect 135 768 169 772
rect 165 764 169 768
rect 173 764 177 776
rect 193 764 197 785
rect 203 764 207 813
rect 225 784 229 852
rect 271 839 275 916
rect 266 827 275 839
rect 269 811 275 827
rect 291 839 295 916
rect 370 873 374 916
rect 367 861 374 873
rect 291 827 294 839
rect 291 811 297 827
rect 269 804 277 811
rect 273 784 277 804
rect 283 804 297 811
rect 283 784 287 804
rect 365 784 369 861
rect 392 819 396 876
rect 400 872 404 876
rect 400 864 418 872
rect 414 853 418 864
rect 385 807 394 819
rect 385 784 389 807
rect 414 796 418 841
rect 455 833 459 876
rect 475 834 479 916
rect 489 857 493 916
rect 509 876 513 916
rect 521 910 525 916
rect 515 864 518 876
rect 489 849 498 857
rect 405 789 418 796
rect 405 784 409 789
rect 455 784 459 821
rect 475 764 479 822
rect 494 820 498 849
rect 514 800 518 864
rect 485 796 518 800
rect 485 764 489 796
rect 523 788 527 898
rect 541 890 545 916
rect 587 912 591 916
rect 555 910 591 912
rect 567 908 591 910
rect 509 776 511 788
rect 507 764 511 776
rect 517 776 519 788
rect 517 764 521 776
rect 539 764 543 878
rect 555 772 559 898
rect 595 884 599 916
rect 615 896 619 936
rect 623 913 627 936
rect 623 906 631 913
rect 593 789 599 884
rect 627 877 631 906
rect 623 871 631 877
rect 623 825 627 871
rect 645 864 649 876
rect 647 852 649 864
rect 593 785 617 789
rect 579 780 597 781
rect 567 776 597 780
rect 555 768 589 772
rect 585 764 589 768
rect 593 764 597 776
rect 613 764 617 785
rect 623 764 627 813
rect 645 784 649 852
rect 691 839 695 916
rect 686 827 695 839
rect 689 811 695 827
rect 711 839 715 916
rect 790 873 794 916
rect 787 861 794 873
rect 711 827 714 839
rect 711 811 717 827
rect 689 804 697 811
rect 693 784 697 804
rect 703 804 717 811
rect 703 784 707 804
rect 785 784 789 861
rect 812 819 816 876
rect 820 872 824 876
rect 890 873 894 916
rect 820 864 838 872
rect 834 853 838 864
rect 887 861 894 873
rect 805 807 814 819
rect 805 784 809 807
rect 834 796 838 841
rect 825 789 838 796
rect 825 784 829 789
rect 885 784 889 861
rect 912 819 916 876
rect 920 872 924 876
rect 920 864 938 872
rect 934 853 938 864
rect 905 807 914 819
rect 905 784 909 807
rect 934 796 938 841
rect 925 789 938 796
rect 985 833 989 916
rect 1057 853 1061 876
rect 1046 841 1061 853
rect 1065 853 1069 876
rect 1111 853 1115 876
rect 1065 841 1074 853
rect 1106 841 1115 853
rect 1119 853 1123 876
rect 1119 841 1134 853
rect 985 821 994 833
rect 925 784 929 789
rect 985 764 989 821
rect 1045 764 1049 841
rect 1065 764 1069 841
rect 1111 764 1115 841
rect 1131 764 1135 841
rect 1205 839 1209 916
rect 1206 827 1209 839
rect 1203 811 1209 827
rect 1225 839 1229 916
rect 1285 839 1289 916
rect 1225 827 1234 839
rect 1286 827 1289 839
rect 1225 811 1231 827
rect 1203 804 1217 811
rect 1213 784 1217 804
rect 1223 804 1231 811
rect 1283 811 1289 827
rect 1305 839 1309 916
rect 1365 839 1369 916
rect 1305 827 1314 839
rect 1366 827 1369 839
rect 1305 811 1311 827
rect 1283 804 1297 811
rect 1223 784 1227 804
rect 1293 784 1297 804
rect 1303 804 1311 811
rect 1363 811 1369 827
rect 1385 839 1389 916
rect 1385 827 1394 839
rect 1385 811 1391 827
rect 1363 804 1377 811
rect 1303 784 1307 804
rect 1373 784 1377 804
rect 1383 804 1391 811
rect 1445 819 1449 876
rect 1465 862 1469 876
rect 1485 862 1489 876
rect 1465 856 1480 862
rect 1485 856 1501 862
rect 1474 833 1480 856
rect 1445 807 1454 819
rect 1383 784 1387 804
rect 1452 764 1456 807
rect 1474 784 1478 821
rect 1494 819 1501 856
rect 1494 794 1501 807
rect 1482 788 1501 794
rect 1541 802 1545 876
rect 1563 839 1567 916
rect 1585 853 1589 916
rect 1631 862 1635 876
rect 1651 862 1655 876
rect 1619 856 1635 862
rect 1640 856 1655 862
rect 1585 841 1594 853
rect 1566 827 1579 839
rect 1541 790 1553 802
rect 1482 784 1486 788
rect 1555 784 1559 790
rect 1575 784 1579 827
rect 1585 784 1589 841
rect 1619 819 1626 856
rect 1640 833 1646 856
rect 1619 794 1626 807
rect 1619 788 1638 794
rect 1634 784 1638 788
rect 1642 784 1646 821
rect 1671 819 1675 876
rect 1666 807 1675 819
rect 1731 819 1735 876
rect 1751 819 1755 876
rect 1731 807 1734 819
rect 1746 807 1755 819
rect 1771 816 1775 876
rect 1791 816 1795 876
rect 1811 816 1815 876
rect 1831 816 1835 876
rect 1851 816 1855 876
rect 1871 816 1875 876
rect 1945 839 1949 916
rect 1946 827 1949 839
rect 1664 764 1668 807
rect 1731 784 1735 807
rect 1751 784 1755 807
rect 1782 804 1795 816
rect 1822 804 1835 816
rect 1862 804 1875 816
rect 1943 811 1949 827
rect 1965 839 1969 916
rect 2037 853 2041 876
rect 2026 841 2041 853
rect 2045 853 2049 876
rect 2096 872 2100 876
rect 2082 864 2100 872
rect 2082 853 2086 864
rect 2045 841 2054 853
rect 1965 827 1974 839
rect 1965 811 1971 827
rect 1943 804 1957 811
rect 1771 784 1775 804
rect 1791 784 1795 804
rect 1811 784 1815 804
rect 1831 784 1835 804
rect 1851 784 1855 804
rect 1871 784 1875 804
rect 1953 784 1957 804
rect 1963 804 1971 811
rect 1963 784 1967 804
rect 2025 764 2029 841
rect 2045 764 2049 841
rect 2082 796 2086 841
rect 2104 819 2108 876
rect 2126 873 2130 916
rect 2126 861 2133 873
rect 2196 872 2200 876
rect 2182 864 2200 872
rect 2106 807 2115 819
rect 2082 789 2095 796
rect 2091 784 2095 789
rect 2111 784 2115 807
rect 2131 784 2135 861
rect 2182 853 2186 864
rect 2182 796 2186 841
rect 2204 819 2208 876
rect 2226 873 2230 916
rect 2226 861 2233 873
rect 2296 872 2300 876
rect 2282 864 2300 872
rect 2206 807 2215 819
rect 2182 789 2195 796
rect 2191 784 2195 789
rect 2211 784 2215 807
rect 2231 784 2235 861
rect 2282 853 2286 864
rect 2282 796 2286 841
rect 2304 819 2308 876
rect 2326 873 2330 916
rect 2326 861 2333 873
rect 2306 807 2315 819
rect 2282 789 2295 796
rect 2291 784 2295 789
rect 2311 784 2315 807
rect 2331 784 2335 861
rect 2391 839 2395 916
rect 2386 827 2395 839
rect 2389 811 2395 827
rect 2411 839 2415 916
rect 2411 827 2414 839
rect 2485 833 2489 916
rect 2553 913 2557 936
rect 2549 906 2557 913
rect 2549 877 2553 906
rect 2561 896 2565 936
rect 2581 884 2585 916
rect 2589 912 2593 916
rect 2589 910 2625 912
rect 2589 908 2613 910
rect 2531 864 2535 876
rect 2549 871 2557 877
rect 2531 852 2533 864
rect 2411 811 2417 827
rect 2389 804 2397 811
rect 2393 784 2397 804
rect 2403 804 2417 811
rect 2485 821 2494 833
rect 2403 784 2407 804
rect 2485 764 2489 821
rect 2531 784 2535 852
rect 2553 825 2557 871
rect 2553 764 2557 813
rect 2581 789 2587 884
rect 2563 785 2587 789
rect 2563 764 2567 785
rect 2583 780 2601 781
rect 2583 776 2613 780
rect 2583 764 2587 776
rect 2621 772 2625 898
rect 2635 890 2639 916
rect 2655 910 2659 916
rect 2591 768 2625 772
rect 2591 764 2595 768
rect 2637 764 2641 878
rect 2653 788 2657 898
rect 2667 876 2671 916
rect 2662 864 2665 876
rect 2662 800 2666 864
rect 2687 857 2691 916
rect 2682 849 2691 857
rect 2682 820 2686 849
rect 2701 834 2705 916
rect 2721 833 2725 876
rect 2790 873 2794 916
rect 2787 861 2794 873
rect 2662 796 2695 800
rect 2661 776 2663 788
rect 2659 764 2663 776
rect 2669 776 2671 788
rect 2669 764 2673 776
rect 2691 764 2695 796
rect 2701 764 2705 822
rect 2721 784 2725 821
rect 2785 784 2789 861
rect 2812 819 2816 876
rect 2820 872 2824 876
rect 2820 864 2838 872
rect 2834 853 2838 864
rect 2805 807 2814 819
rect 2805 784 2809 807
rect 2834 796 2838 841
rect 2825 789 2838 796
rect 2885 833 2889 916
rect 2931 833 2935 916
rect 2991 908 2995 916
rect 2980 904 2995 908
rect 3011 904 3015 916
rect 2980 873 2986 904
rect 3000 900 3015 904
rect 3000 893 3006 900
rect 2986 861 2996 873
rect 2885 821 2894 833
rect 2926 821 2935 833
rect 2825 784 2829 789
rect 2885 764 2889 821
rect 2931 764 2935 821
rect 2992 804 2996 861
rect 3000 804 3004 881
rect 3031 873 3035 916
rect 3008 861 3015 873
rect 3027 861 3035 873
rect 3008 804 3012 861
rect 3091 833 3095 916
rect 3165 839 3169 916
rect 3086 821 3095 833
rect 3166 827 3169 839
rect 3091 764 3095 821
rect 3163 811 3169 827
rect 3185 839 3189 916
rect 3231 872 3235 876
rect 3222 867 3235 872
rect 3185 827 3194 839
rect 3222 833 3226 867
rect 3241 853 3245 876
rect 3261 871 3265 876
rect 3185 811 3191 827
rect 3163 804 3177 811
rect 3173 784 3177 804
rect 3183 804 3191 811
rect 3183 784 3187 804
rect 3222 776 3226 821
rect 3241 777 3245 841
rect 3331 839 3335 916
rect 3326 827 3335 839
rect 3329 811 3335 827
rect 3351 839 3355 916
rect 3411 839 3415 916
rect 3351 827 3354 839
rect 3406 827 3415 839
rect 3351 811 3357 827
rect 3329 804 3337 811
rect 3265 792 3275 804
rect 3271 784 3275 792
rect 3333 784 3337 804
rect 3343 804 3357 811
rect 3409 811 3415 827
rect 3431 839 3435 916
rect 3517 853 3521 876
rect 3506 841 3521 853
rect 3525 853 3529 876
rect 3525 841 3534 853
rect 3431 827 3434 839
rect 3431 811 3437 827
rect 3409 804 3417 811
rect 3343 784 3347 804
rect 3413 784 3417 804
rect 3423 804 3437 811
rect 3423 784 3427 804
rect 3222 771 3235 776
rect 3241 771 3255 777
rect 3231 764 3235 771
rect 3251 764 3255 771
rect 3505 764 3509 841
rect 3525 764 3529 841
rect 3571 839 3575 916
rect 3566 827 3575 839
rect 3569 811 3575 827
rect 3591 839 3595 916
rect 3665 873 3669 916
rect 3685 904 3689 916
rect 3705 908 3709 916
rect 3705 904 3720 908
rect 3685 900 3700 904
rect 3694 893 3700 900
rect 3665 861 3673 873
rect 3685 861 3692 873
rect 3591 827 3594 839
rect 3591 811 3597 827
rect 3569 804 3577 811
rect 3573 784 3577 804
rect 3583 804 3597 811
rect 3688 804 3692 861
rect 3696 804 3700 881
rect 3714 873 3720 904
rect 3765 873 3769 916
rect 3785 904 3789 916
rect 3805 908 3809 916
rect 3805 904 3820 908
rect 3785 900 3800 904
rect 3794 893 3800 900
rect 3704 861 3714 873
rect 3765 861 3773 873
rect 3785 861 3792 873
rect 3704 804 3708 861
rect 3788 804 3792 861
rect 3796 804 3800 881
rect 3814 873 3820 904
rect 3804 861 3814 873
rect 3804 804 3808 861
rect 3851 839 3855 916
rect 3846 827 3855 839
rect 3849 811 3855 827
rect 3871 839 3875 916
rect 3945 873 3949 916
rect 3965 904 3969 916
rect 3985 908 3989 916
rect 3985 904 4000 908
rect 3965 900 3980 904
rect 3974 893 3980 900
rect 3945 861 3953 873
rect 3965 861 3972 873
rect 3871 827 3874 839
rect 3871 811 3877 827
rect 3849 804 3857 811
rect 3583 784 3587 804
rect 3853 784 3857 804
rect 3863 804 3877 811
rect 3968 804 3972 861
rect 3976 804 3980 881
rect 3994 873 4000 904
rect 3984 861 3994 873
rect 3984 804 3988 861
rect 4045 833 4049 916
rect 4110 873 4114 916
rect 4107 861 4114 873
rect 4045 821 4054 833
rect 3863 784 3867 804
rect 4045 764 4049 821
rect 4105 784 4109 861
rect 4132 819 4136 876
rect 4140 872 4144 876
rect 4210 873 4214 916
rect 4391 908 4395 916
rect 4380 904 4395 908
rect 4411 904 4415 916
rect 4140 864 4158 872
rect 4154 853 4158 864
rect 4207 861 4214 873
rect 4125 807 4134 819
rect 4125 784 4129 807
rect 4154 796 4158 841
rect 4145 789 4158 796
rect 4145 784 4149 789
rect 4205 784 4209 861
rect 4232 819 4236 876
rect 4240 872 4244 876
rect 4240 864 4258 872
rect 4254 853 4258 864
rect 4225 807 4234 819
rect 4225 784 4229 807
rect 4254 796 4258 841
rect 4305 819 4309 876
rect 4325 862 4329 876
rect 4345 862 4349 876
rect 4380 873 4386 904
rect 4400 900 4415 904
rect 4400 893 4406 900
rect 4325 856 4340 862
rect 4345 856 4361 862
rect 4386 861 4396 873
rect 4334 833 4340 856
rect 4305 807 4314 819
rect 4245 789 4258 796
rect 4245 784 4249 789
rect 4312 764 4316 807
rect 4334 784 4338 821
rect 4354 819 4361 856
rect 4354 794 4361 807
rect 4392 804 4396 861
rect 4400 804 4404 881
rect 4431 873 4435 916
rect 4408 861 4415 873
rect 4427 861 4435 873
rect 4505 873 4509 916
rect 4525 904 4529 916
rect 4545 908 4549 916
rect 4545 904 4560 908
rect 4525 900 4540 904
rect 4534 893 4540 900
rect 4505 861 4513 873
rect 4525 861 4532 873
rect 4408 804 4412 861
rect 4528 804 4532 861
rect 4536 804 4540 881
rect 4554 873 4560 904
rect 4691 908 4695 916
rect 4680 904 4695 908
rect 4711 904 4715 916
rect 4544 861 4554 873
rect 4544 804 4548 861
rect 4605 819 4609 876
rect 4625 862 4629 876
rect 4645 862 4649 876
rect 4680 873 4686 904
rect 4700 900 4715 904
rect 4700 893 4706 900
rect 4625 856 4640 862
rect 4645 856 4661 862
rect 4686 861 4696 873
rect 4634 833 4640 856
rect 4605 807 4614 819
rect 4342 788 4361 794
rect 4342 784 4346 788
rect 4612 764 4616 807
rect 4634 784 4638 821
rect 4654 819 4661 856
rect 4654 794 4661 807
rect 4692 804 4696 861
rect 4700 804 4704 881
rect 4731 873 4735 916
rect 4708 861 4715 873
rect 4727 861 4735 873
rect 4708 804 4712 861
rect 4642 788 4661 794
rect 4642 784 4646 788
rect 35 740 39 744
rect 55 740 59 744
rect 65 740 69 744
rect 87 740 91 744
rect 97 740 101 744
rect 119 740 123 744
rect 165 740 169 744
rect 173 740 177 744
rect 193 740 197 744
rect 203 740 207 744
rect 225 740 229 744
rect 273 740 277 744
rect 283 740 287 744
rect 365 740 369 744
rect 385 740 389 744
rect 405 740 409 744
rect 455 740 459 744
rect 475 740 479 744
rect 485 740 489 744
rect 507 740 511 744
rect 517 740 521 744
rect 539 740 543 744
rect 585 740 589 744
rect 593 740 597 744
rect 613 740 617 744
rect 623 740 627 744
rect 645 740 649 744
rect 693 740 697 744
rect 703 740 707 744
rect 785 740 789 744
rect 805 740 809 744
rect 825 740 829 744
rect 885 740 889 744
rect 905 740 909 744
rect 925 740 929 744
rect 985 740 989 744
rect 1045 740 1049 744
rect 1065 740 1069 744
rect 1111 740 1115 744
rect 1131 740 1135 744
rect 1213 740 1217 744
rect 1223 740 1227 744
rect 1293 740 1297 744
rect 1303 740 1307 744
rect 1373 740 1377 744
rect 1383 740 1387 744
rect 1452 740 1456 744
rect 1474 740 1478 744
rect 1482 740 1486 744
rect 1555 740 1559 744
rect 1575 740 1579 744
rect 1585 740 1589 744
rect 1634 740 1638 744
rect 1642 740 1646 744
rect 1664 740 1668 744
rect 1731 740 1735 744
rect 1751 740 1755 744
rect 1771 740 1775 744
rect 1791 740 1795 744
rect 1811 740 1815 744
rect 1831 740 1835 744
rect 1851 740 1855 744
rect 1871 740 1875 744
rect 1953 740 1957 744
rect 1963 740 1967 744
rect 2025 740 2029 744
rect 2045 740 2049 744
rect 2091 740 2095 744
rect 2111 740 2115 744
rect 2131 740 2135 744
rect 2191 740 2195 744
rect 2211 740 2215 744
rect 2231 740 2235 744
rect 2291 740 2295 744
rect 2311 740 2315 744
rect 2331 740 2335 744
rect 2393 740 2397 744
rect 2403 740 2407 744
rect 2485 740 2489 744
rect 2531 740 2535 744
rect 2553 740 2557 744
rect 2563 740 2567 744
rect 2583 740 2587 744
rect 2591 740 2595 744
rect 2637 740 2641 744
rect 2659 740 2663 744
rect 2669 740 2673 744
rect 2691 740 2695 744
rect 2701 740 2705 744
rect 2721 740 2725 744
rect 2785 740 2789 744
rect 2805 740 2809 744
rect 2825 740 2829 744
rect 2885 740 2889 744
rect 2931 740 2935 744
rect 2992 740 2996 744
rect 3000 740 3004 744
rect 3008 740 3012 744
rect 3091 740 3095 744
rect 3173 740 3177 744
rect 3183 740 3187 744
rect 3231 740 3235 744
rect 3251 740 3255 744
rect 3271 740 3275 744
rect 3333 740 3337 744
rect 3343 740 3347 744
rect 3413 740 3417 744
rect 3423 740 3427 744
rect 3505 740 3509 744
rect 3525 740 3529 744
rect 3573 740 3577 744
rect 3583 740 3587 744
rect 3688 740 3692 744
rect 3696 740 3700 744
rect 3704 740 3708 744
rect 3788 740 3792 744
rect 3796 740 3800 744
rect 3804 740 3808 744
rect 3853 740 3857 744
rect 3863 740 3867 744
rect 3968 740 3972 744
rect 3976 740 3980 744
rect 3984 740 3988 744
rect 4045 740 4049 744
rect 4105 740 4109 744
rect 4125 740 4129 744
rect 4145 740 4149 744
rect 4205 740 4209 744
rect 4225 740 4229 744
rect 4245 740 4249 744
rect 4312 740 4316 744
rect 4334 740 4338 744
rect 4342 740 4346 744
rect 4392 740 4396 744
rect 4400 740 4404 744
rect 4408 740 4412 744
rect 4528 740 4532 744
rect 4536 740 4540 744
rect 4544 740 4548 744
rect 4612 740 4616 744
rect 4634 740 4638 744
rect 4642 740 4646 744
rect 4692 740 4696 744
rect 4700 740 4704 744
rect 4708 740 4712 744
rect 35 716 39 720
rect 55 716 59 720
rect 65 716 69 720
rect 87 716 91 720
rect 97 716 101 720
rect 119 716 123 720
rect 165 716 169 720
rect 173 716 177 720
rect 193 716 197 720
rect 203 716 207 720
rect 225 716 229 720
rect 271 716 275 720
rect 331 716 335 720
rect 351 716 355 720
rect 371 716 375 720
rect 433 716 437 720
rect 443 716 447 720
rect 511 716 515 720
rect 533 716 537 720
rect 605 716 609 720
rect 651 716 655 720
rect 673 716 677 720
rect 683 716 687 720
rect 703 716 707 720
rect 711 716 715 720
rect 757 716 761 720
rect 779 716 783 720
rect 789 716 793 720
rect 811 716 815 720
rect 821 716 825 720
rect 841 716 845 720
rect 891 716 895 720
rect 911 716 915 720
rect 931 716 935 720
rect 1005 716 1009 720
rect 1025 716 1029 720
rect 1071 716 1075 720
rect 1091 716 1095 720
rect 1111 716 1115 720
rect 1185 716 1189 720
rect 1205 716 1209 720
rect 1225 716 1229 720
rect 1295 716 1299 720
rect 1315 716 1319 720
rect 1325 716 1329 720
rect 1371 716 1375 720
rect 1391 716 1395 720
rect 1451 716 1455 720
rect 1473 716 1477 720
rect 1535 716 1539 720
rect 1555 716 1559 720
rect 1565 716 1569 720
rect 1587 716 1591 720
rect 1597 716 1601 720
rect 1619 716 1623 720
rect 1665 716 1669 720
rect 1673 716 1677 720
rect 1693 716 1697 720
rect 1703 716 1707 720
rect 1725 716 1729 720
rect 1771 716 1775 720
rect 1793 716 1797 720
rect 1865 716 1869 720
rect 1885 716 1889 720
rect 1945 716 1949 720
rect 1965 716 1969 720
rect 2025 716 2029 720
rect 2071 716 2075 720
rect 2091 716 2095 720
rect 2151 716 2155 720
rect 2173 716 2177 720
rect 2183 716 2187 720
rect 2203 716 2207 720
rect 2211 716 2215 720
rect 2257 716 2261 720
rect 2279 716 2283 720
rect 2289 716 2293 720
rect 2311 716 2315 720
rect 2321 716 2325 720
rect 2341 716 2345 720
rect 2394 716 2398 720
rect 2402 716 2406 720
rect 2422 716 2426 720
rect 2430 716 2434 720
rect 2525 716 2529 720
rect 2545 716 2549 720
rect 2565 716 2569 720
rect 2632 716 2636 720
rect 2654 716 2658 720
rect 2662 716 2666 720
rect 2732 716 2736 720
rect 2754 716 2758 720
rect 2762 716 2766 720
rect 2811 716 2815 720
rect 2885 716 2889 720
rect 2905 716 2909 720
rect 2925 716 2929 720
rect 2971 716 2975 720
rect 2991 716 2995 720
rect 3011 716 3015 720
rect 3073 716 3077 720
rect 3083 716 3087 720
rect 3165 716 3169 720
rect 3211 716 3215 720
rect 3308 716 3312 720
rect 3316 716 3320 720
rect 3324 716 3328 720
rect 3385 716 3389 720
rect 3405 716 3409 720
rect 3451 716 3455 720
rect 3471 716 3475 720
rect 3491 716 3495 720
rect 3554 716 3558 720
rect 3562 716 3566 720
rect 3584 716 3588 720
rect 3672 716 3676 720
rect 3694 716 3698 720
rect 3702 716 3706 720
rect 3786 716 3790 720
rect 3794 716 3798 720
rect 3814 716 3818 720
rect 3822 716 3826 720
rect 3908 716 3912 720
rect 3916 716 3920 720
rect 3924 716 3928 720
rect 4008 716 4012 720
rect 4016 716 4020 720
rect 4024 716 4028 720
rect 4071 716 4075 720
rect 4132 716 4136 720
rect 4140 716 4144 720
rect 4148 716 4152 720
rect 4232 716 4236 720
rect 4240 716 4244 720
rect 4248 716 4252 720
rect 4368 716 4372 720
rect 4376 716 4380 720
rect 4384 716 4388 720
rect 4468 716 4472 720
rect 4476 716 4480 720
rect 4484 716 4488 720
rect 4531 716 4535 720
rect 4605 716 4609 720
rect 4625 716 4629 720
rect 4645 716 4649 720
rect 4691 716 4695 720
rect 4711 716 4715 720
rect 4731 716 4735 720
rect 35 639 39 676
rect 55 638 59 696
rect 65 664 69 696
rect 87 684 91 696
rect 89 672 91 684
rect 97 684 101 696
rect 97 672 99 684
rect 65 660 98 664
rect 35 584 39 627
rect 55 544 59 626
rect 74 611 78 640
rect 69 603 78 611
rect 69 544 73 603
rect 94 596 98 660
rect 95 584 98 596
rect 89 544 93 584
rect 103 562 107 672
rect 119 582 123 696
rect 165 692 169 696
rect 135 688 169 692
rect 101 544 105 550
rect 121 544 125 570
rect 135 562 139 688
rect 173 684 177 696
rect 147 680 177 684
rect 159 679 177 680
rect 193 675 197 696
rect 173 671 197 675
rect 173 576 179 671
rect 203 647 207 696
rect 203 589 207 635
rect 225 608 229 676
rect 271 639 275 696
rect 331 671 335 676
rect 266 627 275 639
rect 227 596 229 608
rect 203 583 211 589
rect 225 584 229 596
rect 147 550 171 552
rect 135 548 171 550
rect 167 544 171 548
rect 175 544 179 576
rect 195 524 199 564
rect 207 554 211 583
rect 203 547 211 554
rect 203 524 207 547
rect 271 544 275 627
rect 322 664 335 671
rect 322 619 326 664
rect 351 653 355 676
rect 346 641 355 653
rect 322 596 326 607
rect 322 588 340 596
rect 336 584 340 588
rect 344 584 348 641
rect 371 599 375 676
rect 433 656 437 676
rect 429 649 437 656
rect 443 656 447 676
rect 443 649 457 656
rect 429 633 435 649
rect 426 621 435 633
rect 366 587 373 599
rect 366 544 370 587
rect 431 544 435 621
rect 451 633 457 649
rect 451 621 454 633
rect 451 544 455 621
rect 511 619 515 696
rect 533 670 537 676
rect 535 658 537 670
rect 506 607 515 619
rect 511 544 515 607
rect 605 639 609 696
rect 605 627 614 639
rect 535 590 537 602
rect 533 584 537 590
rect 605 544 609 627
rect 651 608 655 676
rect 673 647 677 696
rect 683 675 687 696
rect 703 684 707 696
rect 711 692 715 696
rect 711 688 745 692
rect 703 680 733 684
rect 703 679 721 680
rect 683 671 707 675
rect 651 596 653 608
rect 651 584 655 596
rect 673 589 677 635
rect 669 583 677 589
rect 669 554 673 583
rect 701 576 707 671
rect 669 547 677 554
rect 673 524 677 547
rect 681 524 685 564
rect 701 544 705 576
rect 741 562 745 688
rect 757 582 761 696
rect 779 684 783 696
rect 781 672 783 684
rect 789 684 793 696
rect 789 672 791 684
rect 709 550 733 552
rect 709 548 745 550
rect 709 544 713 548
rect 755 544 759 570
rect 773 562 777 672
rect 811 664 815 696
rect 782 660 815 664
rect 782 596 786 660
rect 802 611 806 640
rect 821 638 825 696
rect 841 639 845 676
rect 891 671 895 676
rect 882 664 895 671
rect 802 603 811 611
rect 782 584 785 596
rect 775 544 779 550
rect 787 544 791 584
rect 807 544 811 603
rect 821 544 825 626
rect 841 584 845 627
rect 882 619 886 664
rect 911 653 915 676
rect 906 641 915 653
rect 882 596 886 607
rect 882 588 900 596
rect 896 584 900 588
rect 904 584 908 641
rect 931 599 935 676
rect 1005 619 1009 696
rect 1025 619 1029 696
rect 1071 689 1075 696
rect 1091 689 1095 696
rect 1062 684 1075 689
rect 1062 639 1066 684
rect 1006 607 1021 619
rect 926 587 933 599
rect 926 544 930 587
rect 1017 584 1021 607
rect 1025 607 1034 619
rect 1025 584 1029 607
rect 1062 593 1066 627
rect 1081 683 1095 689
rect 1081 619 1085 683
rect 1111 668 1115 676
rect 1105 656 1115 668
rect 1062 588 1075 593
rect 1071 584 1075 588
rect 1081 584 1085 607
rect 1185 599 1189 676
rect 1205 653 1209 676
rect 1225 671 1229 676
rect 1225 664 1238 671
rect 1295 670 1299 676
rect 1205 641 1214 653
rect 1101 584 1105 589
rect 1187 587 1194 599
rect 1190 544 1194 587
rect 1212 584 1216 641
rect 1234 619 1238 664
rect 1281 658 1293 670
rect 1234 596 1238 607
rect 1220 588 1238 596
rect 1220 584 1224 588
rect 1281 584 1285 658
rect 1315 633 1319 676
rect 1306 621 1319 633
rect 1303 544 1307 621
rect 1325 619 1329 676
rect 1371 619 1375 696
rect 1391 619 1395 696
rect 1451 619 1455 696
rect 1473 670 1477 676
rect 1475 658 1477 670
rect 1535 639 1539 676
rect 1555 638 1559 696
rect 1565 664 1569 696
rect 1587 684 1591 696
rect 1589 672 1591 684
rect 1597 684 1601 696
rect 1597 672 1599 684
rect 1565 660 1598 664
rect 1325 607 1334 619
rect 1366 607 1375 619
rect 1325 544 1329 607
rect 1371 584 1375 607
rect 1379 607 1394 619
rect 1446 607 1455 619
rect 1379 584 1383 607
rect 1451 544 1455 607
rect 1475 590 1477 602
rect 1473 584 1477 590
rect 1535 584 1539 627
rect 1555 544 1559 626
rect 1574 611 1578 640
rect 1569 603 1578 611
rect 1569 544 1573 603
rect 1594 596 1598 660
rect 1595 584 1598 596
rect 1589 544 1593 584
rect 1603 562 1607 672
rect 1619 582 1623 696
rect 1665 692 1669 696
rect 1635 688 1669 692
rect 1601 544 1605 550
rect 1621 544 1625 570
rect 1635 562 1639 688
rect 1673 684 1677 696
rect 1647 680 1677 684
rect 1659 679 1677 680
rect 1693 675 1697 696
rect 1673 671 1697 675
rect 1673 576 1679 671
rect 1703 647 1707 696
rect 1703 589 1707 635
rect 1725 608 1729 676
rect 1771 619 1775 696
rect 1793 670 1797 676
rect 1795 658 1797 670
rect 1865 619 1869 696
rect 1885 619 1889 696
rect 1945 619 1949 696
rect 1965 619 1969 696
rect 2025 639 2029 696
rect 2025 627 2034 639
rect 1727 596 1729 608
rect 1766 607 1775 619
rect 1866 607 1881 619
rect 1703 583 1711 589
rect 1725 584 1729 596
rect 1647 550 1671 552
rect 1635 548 1671 550
rect 1667 544 1671 548
rect 1675 544 1679 576
rect 1695 524 1699 564
rect 1707 554 1711 583
rect 1703 547 1711 554
rect 1703 524 1707 547
rect 1771 544 1775 607
rect 1795 590 1797 602
rect 1793 584 1797 590
rect 1877 584 1881 607
rect 1885 607 1894 619
rect 1946 607 1961 619
rect 1885 584 1889 607
rect 1957 584 1961 607
rect 1965 607 1974 619
rect 1965 584 1969 607
rect 2025 544 2029 627
rect 2071 619 2075 696
rect 2091 619 2095 696
rect 2066 607 2075 619
rect 2071 584 2075 607
rect 2079 607 2094 619
rect 2151 608 2155 676
rect 2173 647 2177 696
rect 2183 675 2187 696
rect 2203 684 2207 696
rect 2211 692 2215 696
rect 2211 688 2245 692
rect 2203 680 2233 684
rect 2203 679 2221 680
rect 2183 671 2207 675
rect 2079 584 2083 607
rect 2151 596 2153 608
rect 2151 584 2155 596
rect 2173 589 2177 635
rect 2169 583 2177 589
rect 2169 554 2173 583
rect 2201 576 2207 671
rect 2169 547 2177 554
rect 2173 524 2177 547
rect 2181 524 2185 564
rect 2201 544 2205 576
rect 2241 562 2245 688
rect 2257 582 2261 696
rect 2279 684 2283 696
rect 2281 672 2283 684
rect 2289 684 2293 696
rect 2289 672 2291 684
rect 2209 550 2233 552
rect 2209 548 2245 550
rect 2209 544 2213 548
rect 2255 544 2259 570
rect 2273 562 2277 672
rect 2311 664 2315 696
rect 2282 660 2315 664
rect 2282 596 2286 660
rect 2302 611 2306 640
rect 2321 638 2325 696
rect 2545 689 2549 696
rect 2565 689 2569 696
rect 2545 683 2559 689
rect 2565 684 2578 689
rect 2341 639 2345 676
rect 2394 668 2398 676
rect 2381 661 2398 668
rect 2302 603 2311 611
rect 2282 584 2285 596
rect 2275 544 2279 550
rect 2287 544 2291 584
rect 2307 544 2311 603
rect 2321 544 2325 626
rect 2341 584 2345 627
rect 2381 619 2387 661
rect 2402 653 2406 676
rect 2422 662 2426 676
rect 2430 671 2434 676
rect 2430 667 2460 671
rect 2422 655 2435 662
rect 2431 653 2435 655
rect 2431 641 2433 653
rect 2402 612 2406 641
rect 2387 607 2395 612
rect 2375 606 2395 607
rect 2402 606 2415 612
rect 2391 584 2395 606
rect 2411 584 2415 606
rect 2431 584 2435 641
rect 2454 619 2460 667
rect 2525 668 2529 676
rect 2525 656 2535 668
rect 2555 619 2559 683
rect 2574 639 2578 684
rect 2632 653 2636 696
rect 2625 641 2634 653
rect 2451 607 2454 619
rect 2451 584 2455 607
rect 2535 584 2539 589
rect 2555 584 2559 607
rect 2574 593 2578 627
rect 2565 588 2578 593
rect 2565 584 2569 588
rect 2625 584 2629 641
rect 2654 639 2658 676
rect 2662 672 2666 676
rect 2662 666 2681 672
rect 2674 653 2681 666
rect 2732 653 2736 696
rect 2725 641 2734 653
rect 2654 604 2660 627
rect 2674 604 2681 641
rect 2645 598 2660 604
rect 2665 598 2681 604
rect 2645 584 2649 598
rect 2665 584 2669 598
rect 2725 584 2729 641
rect 2754 639 2758 676
rect 2762 672 2766 676
rect 2762 666 2781 672
rect 2774 653 2781 666
rect 2754 604 2760 627
rect 2774 604 2781 641
rect 2811 639 2815 696
rect 2806 627 2815 639
rect 2745 598 2760 604
rect 2765 598 2781 604
rect 2745 584 2749 598
rect 2765 584 2769 598
rect 2811 544 2815 627
rect 2885 599 2889 676
rect 2905 653 2909 676
rect 2925 671 2929 676
rect 2971 671 2975 676
rect 2925 664 2938 671
rect 2905 641 2914 653
rect 2887 587 2894 599
rect 2890 544 2894 587
rect 2912 584 2916 641
rect 2934 619 2938 664
rect 2962 664 2975 671
rect 2962 619 2966 664
rect 2991 653 2995 676
rect 2986 641 2995 653
rect 2934 596 2938 607
rect 2920 588 2938 596
rect 2962 596 2966 607
rect 2962 588 2980 596
rect 2920 584 2924 588
rect 2976 584 2980 588
rect 2984 584 2988 641
rect 3011 599 3015 676
rect 3073 656 3077 676
rect 3069 649 3077 656
rect 3083 656 3087 676
rect 3083 649 3097 656
rect 3069 633 3075 649
rect 3066 621 3075 633
rect 3006 587 3013 599
rect 3006 544 3010 587
rect 3071 544 3075 621
rect 3091 633 3097 649
rect 3165 639 3169 696
rect 3211 639 3215 696
rect 3091 621 3094 633
rect 3165 627 3174 639
rect 3206 627 3215 639
rect 3091 544 3095 621
rect 3165 544 3169 627
rect 3211 544 3215 627
rect 3308 599 3312 656
rect 3285 587 3293 599
rect 3305 587 3312 599
rect 3285 544 3289 587
rect 3316 579 3320 656
rect 3324 599 3328 656
rect 3385 619 3389 696
rect 3405 619 3409 696
rect 3451 671 3455 676
rect 3442 664 3455 671
rect 3442 619 3446 664
rect 3471 653 3475 676
rect 3466 641 3475 653
rect 3386 607 3401 619
rect 3324 587 3334 599
rect 3314 560 3320 567
rect 3305 556 3320 560
rect 3334 556 3340 587
rect 3397 584 3401 607
rect 3405 607 3414 619
rect 3405 584 3409 607
rect 3442 596 3446 607
rect 3442 588 3460 596
rect 3456 584 3460 588
rect 3464 584 3468 641
rect 3491 599 3495 676
rect 3554 672 3558 676
rect 3539 666 3558 672
rect 3539 653 3546 666
rect 3539 604 3546 641
rect 3562 639 3566 676
rect 3584 653 3588 696
rect 3672 653 3676 696
rect 3586 641 3595 653
rect 3560 604 3566 627
rect 3486 587 3493 599
rect 3539 598 3555 604
rect 3560 598 3575 604
rect 3305 544 3309 556
rect 3325 552 3340 556
rect 3325 544 3329 552
rect 3486 544 3490 587
rect 3551 584 3555 598
rect 3571 584 3575 598
rect 3591 584 3595 641
rect 3665 641 3674 653
rect 3665 584 3669 641
rect 3694 639 3698 676
rect 3702 672 3706 676
rect 3702 666 3721 672
rect 3786 671 3790 676
rect 3714 653 3721 666
rect 3760 667 3790 671
rect 3694 604 3700 627
rect 3714 604 3721 641
rect 3760 619 3766 667
rect 3794 662 3798 676
rect 3785 655 3798 662
rect 3785 653 3789 655
rect 3814 653 3818 676
rect 3822 668 3826 676
rect 3822 661 3839 668
rect 3787 641 3789 653
rect 3766 607 3769 619
rect 3685 598 3700 604
rect 3705 598 3721 604
rect 3685 584 3689 598
rect 3705 584 3709 598
rect 3765 584 3769 607
rect 3785 584 3789 641
rect 3814 612 3818 641
rect 3833 619 3839 661
rect 3805 606 3818 612
rect 3825 607 3833 612
rect 3825 606 3845 607
rect 3805 584 3809 606
rect 3825 584 3829 606
rect 3908 599 3912 656
rect 3885 587 3893 599
rect 3905 587 3912 599
rect 3885 544 3889 587
rect 3916 579 3920 656
rect 3924 599 3928 656
rect 4008 599 4012 656
rect 3924 587 3934 599
rect 3985 587 3993 599
rect 4005 587 4012 599
rect 3914 560 3920 567
rect 3905 556 3920 560
rect 3934 556 3940 587
rect 3905 544 3909 556
rect 3925 552 3940 556
rect 3925 544 3929 552
rect 3985 544 3989 587
rect 4016 579 4020 656
rect 4024 599 4028 656
rect 4071 639 4075 696
rect 4066 627 4075 639
rect 4024 587 4034 599
rect 4014 560 4020 567
rect 4005 556 4020 560
rect 4034 556 4040 587
rect 4005 544 4009 556
rect 4025 552 4040 556
rect 4025 544 4029 552
rect 4071 544 4075 627
rect 4132 599 4136 656
rect 4126 587 4136 599
rect 4120 556 4126 587
rect 4140 579 4144 656
rect 4148 599 4152 656
rect 4232 599 4236 656
rect 4148 587 4155 599
rect 4167 587 4175 599
rect 4226 587 4236 599
rect 4140 560 4146 567
rect 4140 556 4155 560
rect 4120 552 4135 556
rect 4131 544 4135 552
rect 4151 544 4155 556
rect 4171 544 4175 587
rect 4220 556 4226 587
rect 4240 579 4244 656
rect 4248 599 4252 656
rect 4368 599 4372 656
rect 4248 587 4255 599
rect 4267 587 4275 599
rect 4240 560 4246 567
rect 4240 556 4255 560
rect 4220 552 4235 556
rect 4231 544 4235 552
rect 4251 544 4255 556
rect 4271 544 4275 587
rect 4345 587 4353 599
rect 4365 587 4372 599
rect 4345 544 4349 587
rect 4376 579 4380 656
rect 4384 599 4388 656
rect 4468 599 4472 656
rect 4384 587 4394 599
rect 4445 587 4453 599
rect 4465 587 4472 599
rect 4374 560 4380 567
rect 4365 556 4380 560
rect 4394 556 4400 587
rect 4365 544 4369 556
rect 4385 552 4400 556
rect 4385 544 4389 552
rect 4445 544 4449 587
rect 4476 579 4480 656
rect 4484 599 4488 656
rect 4531 639 4535 696
rect 4526 627 4535 639
rect 4484 587 4494 599
rect 4474 560 4480 567
rect 4465 556 4480 560
rect 4494 556 4500 587
rect 4465 544 4469 556
rect 4485 552 4500 556
rect 4485 544 4489 552
rect 4531 544 4535 627
rect 4605 599 4609 676
rect 4625 653 4629 676
rect 4645 671 4649 676
rect 4691 671 4695 676
rect 4645 664 4658 671
rect 4625 641 4634 653
rect 4607 587 4614 599
rect 4610 544 4614 587
rect 4632 584 4636 641
rect 4654 619 4658 664
rect 4682 664 4695 671
rect 4682 619 4686 664
rect 4711 653 4715 676
rect 4706 641 4715 653
rect 4654 596 4658 607
rect 4640 588 4658 596
rect 4682 596 4686 607
rect 4682 588 4700 596
rect 4640 584 4644 588
rect 4696 584 4700 588
rect 4704 584 4708 641
rect 4731 599 4735 676
rect 4726 587 4733 599
rect 4726 544 4730 587
rect 35 500 39 504
rect 55 500 59 504
rect 69 500 73 504
rect 89 500 93 504
rect 101 500 105 504
rect 121 500 125 504
rect 167 500 171 504
rect 175 500 179 504
rect 195 500 199 504
rect 203 500 207 504
rect 225 500 229 504
rect 271 500 275 504
rect 336 500 340 504
rect 344 500 348 504
rect 366 500 370 504
rect 431 500 435 504
rect 451 500 455 504
rect 511 500 515 504
rect 533 500 537 504
rect 605 500 609 504
rect 651 500 655 504
rect 673 500 677 504
rect 681 500 685 504
rect 701 500 705 504
rect 709 500 713 504
rect 755 500 759 504
rect 775 500 779 504
rect 787 500 791 504
rect 807 500 811 504
rect 821 500 825 504
rect 841 500 845 504
rect 896 500 900 504
rect 904 500 908 504
rect 926 500 930 504
rect 1017 500 1021 504
rect 1025 500 1029 504
rect 1071 500 1075 504
rect 1081 500 1085 504
rect 1101 500 1105 504
rect 1190 500 1194 504
rect 1212 500 1216 504
rect 1220 500 1224 504
rect 1281 500 1285 504
rect 1303 500 1307 504
rect 1325 500 1329 504
rect 1371 500 1375 504
rect 1379 500 1383 504
rect 1451 500 1455 504
rect 1473 500 1477 504
rect 1535 500 1539 504
rect 1555 500 1559 504
rect 1569 500 1573 504
rect 1589 500 1593 504
rect 1601 500 1605 504
rect 1621 500 1625 504
rect 1667 500 1671 504
rect 1675 500 1679 504
rect 1695 500 1699 504
rect 1703 500 1707 504
rect 1725 500 1729 504
rect 1771 500 1775 504
rect 1793 500 1797 504
rect 1877 500 1881 504
rect 1885 500 1889 504
rect 1957 500 1961 504
rect 1965 500 1969 504
rect 2025 500 2029 504
rect 2071 500 2075 504
rect 2079 500 2083 504
rect 2151 500 2155 504
rect 2173 500 2177 504
rect 2181 500 2185 504
rect 2201 500 2205 504
rect 2209 500 2213 504
rect 2255 500 2259 504
rect 2275 500 2279 504
rect 2287 500 2291 504
rect 2307 500 2311 504
rect 2321 500 2325 504
rect 2341 500 2345 504
rect 2391 500 2395 504
rect 2411 500 2415 504
rect 2431 500 2435 504
rect 2451 500 2455 504
rect 2535 500 2539 504
rect 2555 500 2559 504
rect 2565 500 2569 504
rect 2625 500 2629 504
rect 2645 500 2649 504
rect 2665 500 2669 504
rect 2725 500 2729 504
rect 2745 500 2749 504
rect 2765 500 2769 504
rect 2811 500 2815 504
rect 2890 500 2894 504
rect 2912 500 2916 504
rect 2920 500 2924 504
rect 2976 500 2980 504
rect 2984 500 2988 504
rect 3006 500 3010 504
rect 3071 500 3075 504
rect 3091 500 3095 504
rect 3165 500 3169 504
rect 3211 500 3215 504
rect 3285 500 3289 504
rect 3305 500 3309 504
rect 3325 500 3329 504
rect 3397 500 3401 504
rect 3405 500 3409 504
rect 3456 500 3460 504
rect 3464 500 3468 504
rect 3486 500 3490 504
rect 3551 500 3555 504
rect 3571 500 3575 504
rect 3591 500 3595 504
rect 3665 500 3669 504
rect 3685 500 3689 504
rect 3705 500 3709 504
rect 3765 500 3769 504
rect 3785 500 3789 504
rect 3805 500 3809 504
rect 3825 500 3829 504
rect 3885 500 3889 504
rect 3905 500 3909 504
rect 3925 500 3929 504
rect 3985 500 3989 504
rect 4005 500 4009 504
rect 4025 500 4029 504
rect 4071 500 4075 504
rect 4131 500 4135 504
rect 4151 500 4155 504
rect 4171 500 4175 504
rect 4231 500 4235 504
rect 4251 500 4255 504
rect 4271 500 4275 504
rect 4345 500 4349 504
rect 4365 500 4369 504
rect 4385 500 4389 504
rect 4445 500 4449 504
rect 4465 500 4469 504
rect 4485 500 4489 504
rect 4531 500 4535 504
rect 4610 500 4614 504
rect 4632 500 4636 504
rect 4640 500 4644 504
rect 4696 500 4700 504
rect 4704 500 4708 504
rect 4726 500 4730 504
rect 35 476 39 480
rect 55 476 59 480
rect 69 476 73 480
rect 89 476 93 480
rect 101 476 105 480
rect 121 476 125 480
rect 167 476 171 480
rect 175 476 179 480
rect 195 476 199 480
rect 203 476 207 480
rect 225 476 229 480
rect 271 476 275 480
rect 291 476 295 480
rect 370 476 374 480
rect 392 476 396 480
rect 400 476 404 480
rect 451 476 455 480
rect 511 476 515 480
rect 531 476 535 480
rect 610 476 614 480
rect 632 476 636 480
rect 640 476 644 480
rect 696 476 700 480
rect 704 476 708 480
rect 726 476 730 480
rect 796 476 800 480
rect 804 476 808 480
rect 826 476 830 480
rect 910 476 914 480
rect 932 476 936 480
rect 940 476 944 480
rect 991 476 995 480
rect 1051 476 1055 480
rect 1071 476 1075 480
rect 1145 476 1149 480
rect 1165 476 1169 480
rect 1185 476 1189 480
rect 1245 476 1249 480
rect 1310 476 1314 480
rect 1332 476 1336 480
rect 1340 476 1344 480
rect 1417 476 1421 480
rect 1425 476 1429 480
rect 1476 476 1480 480
rect 1484 476 1488 480
rect 1506 476 1510 480
rect 1571 476 1575 480
rect 1591 476 1595 480
rect 1651 476 1655 480
rect 1673 476 1677 480
rect 1681 476 1685 480
rect 1701 476 1705 480
rect 1709 476 1713 480
rect 1755 476 1759 480
rect 1775 476 1779 480
rect 1787 476 1791 480
rect 1807 476 1811 480
rect 1821 476 1825 480
rect 1841 476 1845 480
rect 1905 476 1909 480
rect 1925 476 1929 480
rect 1990 476 1994 480
rect 2012 476 2016 480
rect 2020 476 2024 480
rect 2075 476 2079 480
rect 2095 476 2099 480
rect 2109 476 2113 480
rect 2129 476 2133 480
rect 2141 476 2145 480
rect 2161 476 2165 480
rect 2207 476 2211 480
rect 2215 476 2219 480
rect 2235 476 2239 480
rect 2243 476 2247 480
rect 2265 476 2269 480
rect 2325 476 2329 480
rect 2371 476 2375 480
rect 2379 476 2383 480
rect 2451 476 2455 480
rect 2525 476 2529 480
rect 2545 476 2549 480
rect 2591 476 2595 480
rect 2613 476 2617 480
rect 2621 476 2625 480
rect 2641 476 2645 480
rect 2649 476 2653 480
rect 2695 476 2699 480
rect 2715 476 2719 480
rect 2727 476 2731 480
rect 2747 476 2751 480
rect 2761 476 2765 480
rect 2781 476 2785 480
rect 2831 476 2835 480
rect 2851 476 2855 480
rect 2911 476 2915 480
rect 2931 476 2935 480
rect 2951 476 2955 480
rect 2971 476 2975 480
rect 3031 476 3035 480
rect 3039 476 3043 480
rect 3111 476 3115 480
rect 3185 476 3189 480
rect 3205 476 3209 480
rect 3225 476 3229 480
rect 3285 476 3289 480
rect 3305 476 3309 480
rect 3325 476 3329 480
rect 3376 476 3380 480
rect 3384 476 3388 480
rect 3406 476 3410 480
rect 3485 476 3489 480
rect 3531 476 3535 480
rect 3551 476 3555 480
rect 3611 476 3615 480
rect 3631 476 3635 480
rect 3696 476 3700 480
rect 3704 476 3708 480
rect 3726 476 3730 480
rect 3817 476 3821 480
rect 3825 476 3829 480
rect 3897 476 3901 480
rect 3905 476 3909 480
rect 3951 476 3955 480
rect 3973 476 3977 480
rect 3995 476 3999 480
rect 4051 476 4055 480
rect 4059 476 4063 480
rect 4145 476 4149 480
rect 4165 476 4169 480
rect 4185 476 4189 480
rect 4245 476 4249 480
rect 4265 476 4269 480
rect 4285 476 4289 480
rect 4331 476 4335 480
rect 4351 476 4355 480
rect 4371 476 4375 480
rect 4431 476 4435 480
rect 4510 476 4514 480
rect 4532 476 4536 480
rect 4540 476 4544 480
rect 4591 476 4595 480
rect 4651 476 4655 480
rect 4711 476 4715 480
rect 35 353 39 396
rect 55 354 59 436
rect 69 377 73 436
rect 89 396 93 436
rect 101 430 105 436
rect 95 384 98 396
rect 69 369 78 377
rect 35 304 39 341
rect 55 284 59 342
rect 74 340 78 369
rect 94 320 98 384
rect 65 316 98 320
rect 65 284 69 316
rect 103 308 107 418
rect 121 410 125 436
rect 167 432 171 436
rect 135 430 171 432
rect 147 428 171 430
rect 89 296 91 308
rect 87 284 91 296
rect 97 296 99 308
rect 97 284 101 296
rect 119 284 123 398
rect 135 292 139 418
rect 175 404 179 436
rect 195 416 199 456
rect 203 433 207 456
rect 203 426 211 433
rect 173 309 179 404
rect 207 397 211 426
rect 203 391 211 397
rect 203 345 207 391
rect 225 384 229 396
rect 227 372 229 384
rect 173 305 197 309
rect 159 300 177 301
rect 147 296 177 300
rect 135 288 169 292
rect 165 284 169 288
rect 173 284 177 296
rect 193 284 197 305
rect 203 284 207 333
rect 225 304 229 372
rect 271 359 275 436
rect 266 347 275 359
rect 269 331 275 347
rect 291 359 295 436
rect 370 393 374 436
rect 367 381 374 393
rect 291 347 294 359
rect 291 331 297 347
rect 269 324 277 331
rect 273 304 277 324
rect 283 324 297 331
rect 283 304 287 324
rect 365 304 369 381
rect 392 339 396 396
rect 400 392 404 396
rect 400 384 418 392
rect 414 373 418 384
rect 385 327 394 339
rect 385 304 389 327
rect 414 316 418 361
rect 451 353 455 436
rect 511 359 515 436
rect 446 341 455 353
rect 506 347 515 359
rect 405 309 418 316
rect 405 304 409 309
rect 451 284 455 341
rect 509 331 515 347
rect 531 359 535 436
rect 610 393 614 436
rect 607 381 614 393
rect 531 347 534 359
rect 531 331 537 347
rect 509 324 517 331
rect 513 304 517 324
rect 523 324 537 331
rect 523 304 527 324
rect 605 304 609 381
rect 632 339 636 396
rect 640 392 644 396
rect 696 392 700 396
rect 640 384 658 392
rect 654 373 658 384
rect 682 384 700 392
rect 682 373 686 384
rect 625 327 634 339
rect 625 304 629 327
rect 654 316 658 361
rect 645 309 658 316
rect 682 316 686 361
rect 704 339 708 396
rect 726 393 730 436
rect 726 381 733 393
rect 796 392 800 396
rect 782 384 800 392
rect 706 327 715 339
rect 682 309 695 316
rect 645 304 649 309
rect 691 304 695 309
rect 711 304 715 327
rect 731 304 735 381
rect 782 373 786 384
rect 782 316 786 361
rect 804 339 808 396
rect 826 393 830 436
rect 910 393 914 436
rect 826 381 833 393
rect 907 381 914 393
rect 806 327 815 339
rect 782 309 795 316
rect 791 304 795 309
rect 811 304 815 327
rect 831 304 835 381
rect 905 304 909 381
rect 932 339 936 396
rect 940 392 944 396
rect 940 384 958 392
rect 954 373 958 384
rect 925 327 934 339
rect 925 304 929 327
rect 954 316 958 361
rect 991 353 995 436
rect 1051 359 1055 436
rect 986 341 995 353
rect 1046 347 1055 359
rect 945 309 958 316
rect 945 304 949 309
rect 991 284 995 341
rect 1049 331 1055 347
rect 1071 359 1075 436
rect 1071 347 1074 359
rect 1071 331 1077 347
rect 1049 324 1057 331
rect 1053 304 1057 324
rect 1063 324 1077 331
rect 1145 339 1149 396
rect 1165 382 1169 396
rect 1185 382 1189 396
rect 1165 376 1180 382
rect 1185 376 1201 382
rect 1174 353 1180 376
rect 1145 327 1154 339
rect 1063 304 1067 324
rect 1152 284 1156 327
rect 1174 304 1178 341
rect 1194 339 1201 376
rect 1245 353 1249 436
rect 1310 393 1314 436
rect 1307 381 1314 393
rect 1245 341 1254 353
rect 1194 314 1201 327
rect 1182 308 1201 314
rect 1182 304 1186 308
rect 1245 284 1249 341
rect 1305 304 1309 381
rect 1332 339 1336 396
rect 1340 392 1344 396
rect 1340 384 1358 392
rect 1354 373 1358 384
rect 1417 373 1421 396
rect 1406 361 1421 373
rect 1425 373 1429 396
rect 1476 392 1480 396
rect 1462 384 1480 392
rect 1462 373 1466 384
rect 1425 361 1434 373
rect 1325 327 1334 339
rect 1325 304 1329 327
rect 1354 316 1358 361
rect 1345 309 1358 316
rect 1345 304 1349 309
rect 1405 284 1409 361
rect 1425 284 1429 361
rect 1462 316 1466 361
rect 1484 339 1488 396
rect 1506 393 1510 436
rect 1506 381 1513 393
rect 1486 327 1495 339
rect 1462 309 1475 316
rect 1471 304 1475 309
rect 1491 304 1495 327
rect 1511 304 1515 381
rect 1571 359 1575 436
rect 1566 347 1575 359
rect 1569 331 1575 347
rect 1591 359 1595 436
rect 1673 433 1677 456
rect 1669 426 1677 433
rect 1669 397 1673 426
rect 1681 416 1685 456
rect 1701 404 1705 436
rect 1709 432 1713 436
rect 1709 430 1745 432
rect 1709 428 1733 430
rect 1651 384 1655 396
rect 1669 391 1677 397
rect 1651 372 1653 384
rect 1591 347 1594 359
rect 1591 331 1597 347
rect 1569 324 1577 331
rect 1573 304 1577 324
rect 1583 324 1597 331
rect 1583 304 1587 324
rect 1651 304 1655 372
rect 1673 345 1677 391
rect 1673 284 1677 333
rect 1701 309 1707 404
rect 1683 305 1707 309
rect 1683 284 1687 305
rect 1703 300 1721 301
rect 1703 296 1733 300
rect 1703 284 1707 296
rect 1741 292 1745 418
rect 1755 410 1759 436
rect 1775 430 1779 436
rect 1711 288 1745 292
rect 1711 284 1715 288
rect 1757 284 1761 398
rect 1773 308 1777 418
rect 1787 396 1791 436
rect 1782 384 1785 396
rect 1782 320 1786 384
rect 1807 377 1811 436
rect 1802 369 1811 377
rect 1802 340 1806 369
rect 1821 354 1825 436
rect 1841 353 1845 396
rect 1905 359 1909 436
rect 1782 316 1815 320
rect 1781 296 1783 308
rect 1779 284 1783 296
rect 1789 296 1791 308
rect 1789 284 1793 296
rect 1811 284 1815 316
rect 1821 284 1825 342
rect 1906 347 1909 359
rect 1841 304 1845 341
rect 1903 331 1909 347
rect 1925 359 1929 436
rect 1990 393 1994 436
rect 1987 381 1994 393
rect 1925 347 1934 359
rect 1925 331 1931 347
rect 1903 324 1917 331
rect 1913 304 1917 324
rect 1923 324 1931 331
rect 1923 304 1927 324
rect 1985 304 1989 381
rect 2012 339 2016 396
rect 2020 392 2024 396
rect 2020 384 2038 392
rect 2034 373 2038 384
rect 2005 327 2014 339
rect 2005 304 2009 327
rect 2034 316 2038 361
rect 2075 353 2079 396
rect 2095 354 2099 436
rect 2109 377 2113 436
rect 2129 396 2133 436
rect 2141 430 2145 436
rect 2135 384 2138 396
rect 2109 369 2118 377
rect 2025 309 2038 316
rect 2025 304 2029 309
rect 2075 304 2079 341
rect 2095 284 2099 342
rect 2114 340 2118 369
rect 2134 320 2138 384
rect 2105 316 2138 320
rect 2105 284 2109 316
rect 2143 308 2147 418
rect 2161 410 2165 436
rect 2207 432 2211 436
rect 2175 430 2211 432
rect 2187 428 2211 430
rect 2129 296 2131 308
rect 2127 284 2131 296
rect 2137 296 2139 308
rect 2137 284 2141 296
rect 2159 284 2163 398
rect 2175 292 2179 418
rect 2215 404 2219 436
rect 2235 416 2239 456
rect 2243 433 2247 456
rect 2243 426 2251 433
rect 2213 309 2219 404
rect 2247 397 2251 426
rect 2243 391 2251 397
rect 2243 345 2247 391
rect 2265 384 2269 396
rect 2267 372 2269 384
rect 2213 305 2237 309
rect 2199 300 2217 301
rect 2187 296 2217 300
rect 2175 288 2209 292
rect 2205 284 2209 288
rect 2213 284 2217 296
rect 2233 284 2237 305
rect 2243 284 2247 333
rect 2265 304 2269 372
rect 2325 353 2329 436
rect 2371 373 2375 396
rect 2366 361 2375 373
rect 2379 373 2383 396
rect 2379 361 2394 373
rect 2325 341 2334 353
rect 2325 284 2329 341
rect 2371 284 2375 361
rect 2391 284 2395 361
rect 2451 353 2455 436
rect 2525 359 2529 436
rect 2446 341 2455 353
rect 2526 347 2529 359
rect 2451 284 2455 341
rect 2523 331 2529 347
rect 2545 359 2549 436
rect 2613 433 2617 456
rect 2609 426 2617 433
rect 2609 397 2613 426
rect 2621 416 2625 456
rect 2641 404 2645 436
rect 2649 432 2653 436
rect 2649 430 2685 432
rect 2649 428 2673 430
rect 2591 384 2595 396
rect 2609 391 2617 397
rect 2591 372 2593 384
rect 2545 347 2554 359
rect 2545 331 2551 347
rect 2523 324 2537 331
rect 2533 304 2537 324
rect 2543 324 2551 331
rect 2543 304 2547 324
rect 2591 304 2595 372
rect 2613 345 2617 391
rect 2613 284 2617 333
rect 2641 309 2647 404
rect 2623 305 2647 309
rect 2623 284 2627 305
rect 2643 300 2661 301
rect 2643 296 2673 300
rect 2643 284 2647 296
rect 2681 292 2685 418
rect 2695 410 2699 436
rect 2715 430 2719 436
rect 2651 288 2685 292
rect 2651 284 2655 288
rect 2697 284 2701 398
rect 2713 308 2717 418
rect 2727 396 2731 436
rect 2722 384 2725 396
rect 2722 320 2726 384
rect 2747 377 2751 436
rect 2742 369 2751 377
rect 2742 340 2746 369
rect 2761 354 2765 436
rect 2781 353 2785 396
rect 2831 359 2835 436
rect 2722 316 2755 320
rect 2721 296 2723 308
rect 2719 284 2723 296
rect 2729 296 2731 308
rect 2729 284 2733 296
rect 2751 284 2755 316
rect 2761 284 2765 342
rect 2826 347 2835 359
rect 2781 304 2785 341
rect 2829 331 2835 347
rect 2851 359 2855 436
rect 2911 374 2915 396
rect 2931 374 2935 396
rect 2895 373 2915 374
rect 2907 368 2915 373
rect 2922 368 2935 374
rect 2851 347 2854 359
rect 2851 331 2857 347
rect 2829 324 2837 331
rect 2833 304 2837 324
rect 2843 324 2857 331
rect 2843 304 2847 324
rect 2901 319 2907 361
rect 2922 339 2926 368
rect 2951 339 2955 396
rect 2971 373 2975 396
rect 3031 373 3035 396
rect 2971 361 2974 373
rect 3026 361 3035 373
rect 3039 373 3043 396
rect 3039 361 3054 373
rect 2951 327 2953 339
rect 2901 312 2918 319
rect 2914 304 2918 312
rect 2922 304 2926 327
rect 2951 325 2955 327
rect 2942 318 2955 325
rect 2942 304 2946 318
rect 2974 313 2980 361
rect 2950 309 2980 313
rect 2950 304 2954 309
rect 3031 284 3035 361
rect 3051 284 3055 361
rect 3111 353 3115 436
rect 3185 393 3189 436
rect 3205 424 3209 436
rect 3225 428 3229 436
rect 3225 424 3240 428
rect 3205 420 3220 424
rect 3214 413 3220 420
rect 3185 381 3193 393
rect 3205 381 3212 393
rect 3106 341 3115 353
rect 3111 284 3115 341
rect 3208 324 3212 381
rect 3216 324 3220 401
rect 3234 393 3240 424
rect 3285 393 3289 436
rect 3305 424 3309 436
rect 3325 428 3329 436
rect 3325 424 3340 428
rect 3305 420 3320 424
rect 3314 413 3320 420
rect 3224 381 3234 393
rect 3285 381 3293 393
rect 3305 381 3312 393
rect 3224 324 3228 381
rect 3308 324 3312 381
rect 3316 324 3320 401
rect 3334 393 3340 424
rect 3324 381 3334 393
rect 3376 392 3380 396
rect 3362 384 3380 392
rect 3324 324 3328 381
rect 3362 373 3366 384
rect 3362 316 3366 361
rect 3384 339 3388 396
rect 3406 393 3410 436
rect 3406 381 3413 393
rect 3386 327 3395 339
rect 3362 309 3375 316
rect 3371 304 3375 309
rect 3391 304 3395 327
rect 3411 304 3415 381
rect 3485 353 3489 436
rect 3531 359 3535 436
rect 3485 341 3494 353
rect 3526 347 3535 359
rect 3485 284 3489 341
rect 3529 331 3535 347
rect 3551 359 3555 436
rect 3611 359 3615 436
rect 3551 347 3554 359
rect 3606 347 3615 359
rect 3551 331 3557 347
rect 3529 324 3537 331
rect 3533 304 3537 324
rect 3543 324 3557 331
rect 3609 331 3615 347
rect 3631 359 3635 436
rect 3696 392 3700 396
rect 3682 384 3700 392
rect 3682 373 3686 384
rect 3631 347 3634 359
rect 3631 331 3637 347
rect 3609 324 3617 331
rect 3543 304 3547 324
rect 3613 304 3617 324
rect 3623 324 3637 331
rect 3623 304 3627 324
rect 3682 316 3686 361
rect 3704 339 3708 396
rect 3726 393 3730 436
rect 3726 381 3733 393
rect 3706 327 3715 339
rect 3682 309 3695 316
rect 3691 304 3695 309
rect 3711 304 3715 327
rect 3731 304 3735 381
rect 3817 373 3821 396
rect 3806 361 3821 373
rect 3825 373 3829 396
rect 3897 373 3901 396
rect 3825 361 3834 373
rect 3886 361 3901 373
rect 3905 373 3909 396
rect 3951 373 3955 436
rect 3905 361 3914 373
rect 3946 361 3955 373
rect 3805 284 3809 361
rect 3825 284 3829 361
rect 3885 284 3889 361
rect 3905 284 3909 361
rect 3951 304 3955 361
rect 3973 359 3977 436
rect 3961 347 3974 359
rect 3961 304 3965 347
rect 3995 322 3999 396
rect 4051 373 4055 396
rect 4046 361 4055 373
rect 4059 373 4063 396
rect 4059 361 4074 373
rect 3987 310 3999 322
rect 3981 304 3985 310
rect 4051 284 4055 361
rect 4071 284 4075 361
rect 4145 339 4149 396
rect 4165 382 4169 396
rect 4185 382 4189 396
rect 4245 393 4249 436
rect 4265 424 4269 436
rect 4285 428 4289 436
rect 4285 424 4300 428
rect 4265 420 4280 424
rect 4274 413 4280 420
rect 4165 376 4180 382
rect 4185 376 4201 382
rect 4245 381 4253 393
rect 4265 381 4272 393
rect 4174 353 4180 376
rect 4145 327 4154 339
rect 4152 284 4156 327
rect 4174 304 4178 341
rect 4194 339 4201 376
rect 4194 314 4201 327
rect 4268 324 4272 381
rect 4276 324 4280 401
rect 4294 393 4300 424
rect 4284 381 4294 393
rect 4331 382 4335 396
rect 4351 382 4355 396
rect 4284 324 4288 381
rect 4319 376 4335 382
rect 4340 376 4355 382
rect 4319 339 4326 376
rect 4340 353 4346 376
rect 4182 308 4201 314
rect 4182 304 4186 308
rect 4319 314 4326 327
rect 4319 308 4338 314
rect 4334 304 4338 308
rect 4342 304 4346 341
rect 4371 339 4375 396
rect 4431 353 4435 436
rect 4510 393 4514 436
rect 4507 381 4514 393
rect 4426 341 4435 353
rect 4366 327 4375 339
rect 4364 284 4368 327
rect 4431 284 4435 341
rect 4505 304 4509 381
rect 4532 339 4536 396
rect 4540 392 4544 396
rect 4540 384 4558 392
rect 4554 373 4558 384
rect 4525 327 4534 339
rect 4525 304 4529 327
rect 4554 316 4558 361
rect 4591 353 4595 436
rect 4651 353 4655 436
rect 4711 353 4715 436
rect 4586 341 4595 353
rect 4646 341 4655 353
rect 4706 341 4715 353
rect 4545 309 4558 316
rect 4545 304 4549 309
rect 4591 284 4595 341
rect 4651 284 4655 341
rect 4711 284 4715 341
rect 35 260 39 264
rect 55 260 59 264
rect 65 260 69 264
rect 87 260 91 264
rect 97 260 101 264
rect 119 260 123 264
rect 165 260 169 264
rect 173 260 177 264
rect 193 260 197 264
rect 203 260 207 264
rect 225 260 229 264
rect 273 260 277 264
rect 283 260 287 264
rect 365 260 369 264
rect 385 260 389 264
rect 405 260 409 264
rect 451 260 455 264
rect 513 260 517 264
rect 523 260 527 264
rect 605 260 609 264
rect 625 260 629 264
rect 645 260 649 264
rect 691 260 695 264
rect 711 260 715 264
rect 731 260 735 264
rect 791 260 795 264
rect 811 260 815 264
rect 831 260 835 264
rect 905 260 909 264
rect 925 260 929 264
rect 945 260 949 264
rect 991 260 995 264
rect 1053 260 1057 264
rect 1063 260 1067 264
rect 1152 260 1156 264
rect 1174 260 1178 264
rect 1182 260 1186 264
rect 1245 260 1249 264
rect 1305 260 1309 264
rect 1325 260 1329 264
rect 1345 260 1349 264
rect 1405 260 1409 264
rect 1425 260 1429 264
rect 1471 260 1475 264
rect 1491 260 1495 264
rect 1511 260 1515 264
rect 1573 260 1577 264
rect 1583 260 1587 264
rect 1651 260 1655 264
rect 1673 260 1677 264
rect 1683 260 1687 264
rect 1703 260 1707 264
rect 1711 260 1715 264
rect 1757 260 1761 264
rect 1779 260 1783 264
rect 1789 260 1793 264
rect 1811 260 1815 264
rect 1821 260 1825 264
rect 1841 260 1845 264
rect 1913 260 1917 264
rect 1923 260 1927 264
rect 1985 260 1989 264
rect 2005 260 2009 264
rect 2025 260 2029 264
rect 2075 260 2079 264
rect 2095 260 2099 264
rect 2105 260 2109 264
rect 2127 260 2131 264
rect 2137 260 2141 264
rect 2159 260 2163 264
rect 2205 260 2209 264
rect 2213 260 2217 264
rect 2233 260 2237 264
rect 2243 260 2247 264
rect 2265 260 2269 264
rect 2325 260 2329 264
rect 2371 260 2375 264
rect 2391 260 2395 264
rect 2451 260 2455 264
rect 2533 260 2537 264
rect 2543 260 2547 264
rect 2591 260 2595 264
rect 2613 260 2617 264
rect 2623 260 2627 264
rect 2643 260 2647 264
rect 2651 260 2655 264
rect 2697 260 2701 264
rect 2719 260 2723 264
rect 2729 260 2733 264
rect 2751 260 2755 264
rect 2761 260 2765 264
rect 2781 260 2785 264
rect 2833 260 2837 264
rect 2843 260 2847 264
rect 2914 260 2918 264
rect 2922 260 2926 264
rect 2942 260 2946 264
rect 2950 260 2954 264
rect 3031 260 3035 264
rect 3051 260 3055 264
rect 3111 260 3115 264
rect 3208 260 3212 264
rect 3216 260 3220 264
rect 3224 260 3228 264
rect 3308 260 3312 264
rect 3316 260 3320 264
rect 3324 260 3328 264
rect 3371 260 3375 264
rect 3391 260 3395 264
rect 3411 260 3415 264
rect 3485 260 3489 264
rect 3533 260 3537 264
rect 3543 260 3547 264
rect 3613 260 3617 264
rect 3623 260 3627 264
rect 3691 260 3695 264
rect 3711 260 3715 264
rect 3731 260 3735 264
rect 3805 260 3809 264
rect 3825 260 3829 264
rect 3885 260 3889 264
rect 3905 260 3909 264
rect 3951 260 3955 264
rect 3961 260 3965 264
rect 3981 260 3985 264
rect 4051 260 4055 264
rect 4071 260 4075 264
rect 4152 260 4156 264
rect 4174 260 4178 264
rect 4182 260 4186 264
rect 4268 260 4272 264
rect 4276 260 4280 264
rect 4284 260 4288 264
rect 4334 260 4338 264
rect 4342 260 4346 264
rect 4364 260 4368 264
rect 4431 260 4435 264
rect 4505 260 4509 264
rect 4525 260 4529 264
rect 4545 260 4549 264
rect 4591 260 4595 264
rect 4651 260 4655 264
rect 4711 260 4715 264
rect 35 236 39 240
rect 55 236 59 240
rect 65 236 69 240
rect 87 236 91 240
rect 97 236 101 240
rect 119 236 123 240
rect 165 236 169 240
rect 173 236 177 240
rect 193 236 197 240
rect 203 236 207 240
rect 225 236 229 240
rect 274 236 278 240
rect 282 236 286 240
rect 302 236 306 240
rect 310 236 314 240
rect 391 236 395 240
rect 411 236 415 240
rect 472 236 476 240
rect 480 236 484 240
rect 488 236 492 240
rect 585 236 589 240
rect 605 236 609 240
rect 625 236 629 240
rect 692 236 696 240
rect 714 236 718 240
rect 722 236 726 240
rect 771 236 775 240
rect 793 236 797 240
rect 803 236 807 240
rect 823 236 827 240
rect 831 236 835 240
rect 877 236 881 240
rect 899 236 903 240
rect 909 236 913 240
rect 931 236 935 240
rect 941 236 945 240
rect 961 236 965 240
rect 1025 236 1029 240
rect 1045 236 1049 240
rect 1065 236 1069 240
rect 1125 236 1129 240
rect 1185 236 1189 240
rect 1205 236 1209 240
rect 1265 236 1269 240
rect 1325 236 1329 240
rect 1345 236 1349 240
rect 1365 236 1369 240
rect 1425 236 1429 240
rect 1485 236 1489 240
rect 1531 236 1535 240
rect 1551 236 1555 240
rect 1632 236 1636 240
rect 1654 236 1658 240
rect 1662 236 1666 240
rect 1715 236 1719 240
rect 1735 236 1739 240
rect 1745 236 1749 240
rect 1767 236 1771 240
rect 1777 236 1781 240
rect 1799 236 1803 240
rect 1845 236 1849 240
rect 1853 236 1857 240
rect 1873 236 1877 240
rect 1883 236 1887 240
rect 1905 236 1909 240
rect 1965 236 1969 240
rect 1985 236 1989 240
rect 2005 236 2009 240
rect 2051 236 2055 240
rect 2111 236 2115 240
rect 2131 236 2135 240
rect 2191 236 2195 240
rect 2211 236 2215 240
rect 2285 236 2289 240
rect 2305 236 2309 240
rect 2351 236 2355 240
rect 2371 236 2375 240
rect 2445 236 2449 240
rect 2491 236 2495 240
rect 2513 236 2517 240
rect 2523 236 2527 240
rect 2543 236 2547 240
rect 2551 236 2555 240
rect 2597 236 2601 240
rect 2619 236 2623 240
rect 2629 236 2633 240
rect 2651 236 2655 240
rect 2661 236 2665 240
rect 2681 236 2685 240
rect 2731 236 2735 240
rect 2753 236 2757 240
rect 2763 236 2767 240
rect 2783 236 2787 240
rect 2791 236 2795 240
rect 2837 236 2841 240
rect 2859 236 2863 240
rect 2869 236 2873 240
rect 2891 236 2895 240
rect 2901 236 2905 240
rect 2921 236 2925 240
rect 2971 236 2975 240
rect 2991 236 2995 240
rect 3011 236 3015 240
rect 3031 236 3035 240
rect 3105 236 3109 240
rect 3125 236 3129 240
rect 3145 236 3149 240
rect 3191 236 3195 240
rect 3211 236 3215 240
rect 3231 236 3235 240
rect 3305 236 3309 240
rect 3353 236 3357 240
rect 3363 236 3367 240
rect 3468 236 3472 240
rect 3476 236 3480 240
rect 3484 236 3488 240
rect 3545 236 3549 240
rect 3612 236 3616 240
rect 3634 236 3638 240
rect 3642 236 3646 240
rect 3705 236 3709 240
rect 3725 236 3729 240
rect 3771 236 3775 240
rect 3831 236 3835 240
rect 3851 236 3855 240
rect 3871 236 3875 240
rect 3931 236 3935 240
rect 3951 236 3955 240
rect 4048 236 4052 240
rect 4056 236 4060 240
rect 4064 236 4068 240
rect 4113 236 4117 240
rect 4123 236 4127 240
rect 4228 236 4232 240
rect 4236 236 4240 240
rect 4244 236 4248 240
rect 4313 236 4317 240
rect 4323 236 4327 240
rect 4408 236 4412 240
rect 4416 236 4420 240
rect 4424 236 4428 240
rect 4473 236 4477 240
rect 4483 236 4487 240
rect 4552 236 4556 240
rect 4560 236 4564 240
rect 4568 236 4572 240
rect 4672 236 4676 240
rect 4694 236 4698 240
rect 4702 236 4706 240
rect 35 159 39 196
rect 55 158 59 216
rect 65 184 69 216
rect 87 204 91 216
rect 89 192 91 204
rect 97 204 101 216
rect 97 192 99 204
rect 65 180 98 184
rect 35 104 39 147
rect 55 64 59 146
rect 74 131 78 160
rect 69 123 78 131
rect 69 64 73 123
rect 94 116 98 180
rect 95 104 98 116
rect 89 64 93 104
rect 103 82 107 192
rect 119 102 123 216
rect 165 212 169 216
rect 135 208 169 212
rect 101 64 105 70
rect 121 64 125 90
rect 135 82 139 208
rect 173 204 177 216
rect 147 200 177 204
rect 159 199 177 200
rect 193 195 197 216
rect 173 191 197 195
rect 173 96 179 191
rect 203 167 207 216
rect 203 109 207 155
rect 225 128 229 196
rect 274 188 278 196
rect 261 181 278 188
rect 261 139 267 181
rect 282 173 286 196
rect 302 182 306 196
rect 310 191 314 196
rect 310 187 340 191
rect 302 175 315 182
rect 311 173 315 175
rect 311 161 313 173
rect 227 116 229 128
rect 282 132 286 161
rect 267 127 275 132
rect 255 126 275 127
rect 282 126 295 132
rect 203 103 211 109
rect 225 104 229 116
rect 271 104 275 126
rect 291 104 295 126
rect 311 104 315 161
rect 334 139 340 187
rect 391 139 395 216
rect 411 139 415 216
rect 605 209 609 216
rect 625 209 629 216
rect 605 203 619 209
rect 625 204 638 209
rect 585 188 589 196
rect 585 176 595 188
rect 331 127 334 139
rect 386 127 395 139
rect 331 104 335 127
rect 391 104 395 127
rect 399 127 414 139
rect 399 104 403 127
rect 472 119 476 176
rect 466 107 476 119
rect 147 70 171 72
rect 135 68 171 70
rect 167 64 171 68
rect 175 64 179 96
rect 195 44 199 84
rect 207 74 211 103
rect 203 67 211 74
rect 203 44 207 67
rect 460 76 466 107
rect 480 99 484 176
rect 488 119 492 176
rect 615 139 619 203
rect 634 159 638 204
rect 692 173 696 216
rect 685 161 694 173
rect 488 107 495 119
rect 507 107 515 119
rect 480 80 486 87
rect 480 76 495 80
rect 460 72 475 76
rect 471 64 475 72
rect 491 64 495 76
rect 511 64 515 107
rect 595 104 599 109
rect 615 104 619 127
rect 634 113 638 147
rect 625 108 638 113
rect 625 104 629 108
rect 685 104 689 161
rect 714 159 718 196
rect 722 192 726 196
rect 722 186 741 192
rect 734 173 741 186
rect 714 124 720 147
rect 734 124 741 161
rect 705 118 720 124
rect 725 118 741 124
rect 771 128 775 196
rect 793 167 797 216
rect 803 195 807 216
rect 823 204 827 216
rect 831 212 835 216
rect 831 208 865 212
rect 823 200 853 204
rect 823 199 841 200
rect 803 191 827 195
rect 705 104 709 118
rect 725 104 729 118
rect 771 116 773 128
rect 771 104 775 116
rect 793 109 797 155
rect 789 103 797 109
rect 789 74 793 103
rect 821 96 827 191
rect 789 67 797 74
rect 793 44 797 67
rect 801 44 805 84
rect 821 64 825 96
rect 861 82 865 208
rect 877 102 881 216
rect 899 204 903 216
rect 901 192 903 204
rect 909 204 913 216
rect 909 192 911 204
rect 829 70 853 72
rect 829 68 865 70
rect 829 64 833 68
rect 875 64 879 90
rect 893 82 897 192
rect 931 184 935 216
rect 902 180 935 184
rect 902 116 906 180
rect 922 131 926 160
rect 941 158 945 216
rect 961 159 965 196
rect 922 123 931 131
rect 902 104 905 116
rect 895 64 899 70
rect 907 64 911 104
rect 927 64 931 123
rect 941 64 945 146
rect 961 104 965 147
rect 1025 119 1029 196
rect 1045 173 1049 196
rect 1065 191 1069 196
rect 1065 184 1078 191
rect 1045 161 1054 173
rect 1027 107 1034 119
rect 1030 64 1034 107
rect 1052 104 1056 161
rect 1074 139 1078 184
rect 1125 159 1129 216
rect 1125 147 1134 159
rect 1074 116 1078 127
rect 1060 108 1078 116
rect 1060 104 1064 108
rect 1125 64 1129 147
rect 1185 139 1189 216
rect 1205 139 1209 216
rect 1265 159 1269 216
rect 1265 147 1274 159
rect 1186 127 1201 139
rect 1197 104 1201 127
rect 1205 127 1214 139
rect 1205 104 1209 127
rect 1265 64 1269 147
rect 1325 119 1329 196
rect 1345 173 1349 196
rect 1365 191 1369 196
rect 1365 184 1378 191
rect 1345 161 1354 173
rect 1327 107 1334 119
rect 1330 64 1334 107
rect 1352 104 1356 161
rect 1374 139 1378 184
rect 1425 159 1429 216
rect 1485 159 1489 216
rect 1425 147 1434 159
rect 1485 147 1494 159
rect 1374 116 1378 127
rect 1360 108 1378 116
rect 1360 104 1364 108
rect 1425 64 1429 147
rect 1485 64 1489 147
rect 1531 139 1535 216
rect 1551 139 1555 216
rect 1632 173 1636 216
rect 1625 161 1634 173
rect 1526 127 1535 139
rect 1531 104 1535 127
rect 1539 127 1554 139
rect 1539 104 1543 127
rect 1625 104 1629 161
rect 1654 159 1658 196
rect 1662 192 1666 196
rect 1662 186 1681 192
rect 1674 173 1681 186
rect 1654 124 1660 147
rect 1674 124 1681 161
rect 1715 159 1719 196
rect 1735 158 1739 216
rect 1745 184 1749 216
rect 1767 204 1771 216
rect 1769 192 1771 204
rect 1777 204 1781 216
rect 1777 192 1779 204
rect 1745 180 1778 184
rect 1645 118 1660 124
rect 1665 118 1681 124
rect 1645 104 1649 118
rect 1665 104 1669 118
rect 1715 104 1719 147
rect 1735 64 1739 146
rect 1754 131 1758 160
rect 1749 123 1758 131
rect 1749 64 1753 123
rect 1774 116 1778 180
rect 1775 104 1778 116
rect 1769 64 1773 104
rect 1783 82 1787 192
rect 1799 102 1803 216
rect 1845 212 1849 216
rect 1815 208 1849 212
rect 1781 64 1785 70
rect 1801 64 1805 90
rect 1815 82 1819 208
rect 1853 204 1857 216
rect 1827 200 1857 204
rect 1839 199 1857 200
rect 1873 195 1877 216
rect 1853 191 1877 195
rect 1853 96 1859 191
rect 1883 167 1887 216
rect 1883 109 1887 155
rect 1905 128 1909 196
rect 1907 116 1909 128
rect 1965 119 1969 196
rect 1985 173 1989 196
rect 2005 191 2009 196
rect 2005 184 2018 191
rect 1985 161 1994 173
rect 1883 103 1891 109
rect 1905 104 1909 116
rect 1967 107 1974 119
rect 1827 70 1851 72
rect 1815 68 1851 70
rect 1847 64 1851 68
rect 1855 64 1859 96
rect 1875 44 1879 84
rect 1887 74 1891 103
rect 1883 67 1891 74
rect 1883 44 1887 67
rect 1970 64 1974 107
rect 1992 104 1996 161
rect 2014 139 2018 184
rect 2051 159 2055 216
rect 2046 147 2055 159
rect 2014 116 2018 127
rect 2000 108 2018 116
rect 2000 104 2004 108
rect 2051 64 2055 147
rect 2111 139 2115 216
rect 2131 139 2135 216
rect 2191 139 2195 216
rect 2211 139 2215 216
rect 2285 139 2289 216
rect 2305 139 2309 216
rect 2351 139 2355 216
rect 2371 139 2375 216
rect 2445 159 2449 216
rect 2445 147 2454 159
rect 2106 127 2115 139
rect 2111 104 2115 127
rect 2119 127 2134 139
rect 2186 127 2195 139
rect 2119 104 2123 127
rect 2191 104 2195 127
rect 2199 127 2214 139
rect 2286 127 2301 139
rect 2199 104 2203 127
rect 2297 104 2301 127
rect 2305 127 2314 139
rect 2346 127 2355 139
rect 2305 104 2309 127
rect 2351 104 2355 127
rect 2359 127 2374 139
rect 2359 104 2363 127
rect 2445 64 2449 147
rect 2491 128 2495 196
rect 2513 167 2517 216
rect 2523 195 2527 216
rect 2543 204 2547 216
rect 2551 212 2555 216
rect 2551 208 2585 212
rect 2543 200 2573 204
rect 2543 199 2561 200
rect 2523 191 2547 195
rect 2491 116 2493 128
rect 2491 104 2495 116
rect 2513 109 2517 155
rect 2509 103 2517 109
rect 2509 74 2513 103
rect 2541 96 2547 191
rect 2509 67 2517 74
rect 2513 44 2517 67
rect 2521 44 2525 84
rect 2541 64 2545 96
rect 2581 82 2585 208
rect 2597 102 2601 216
rect 2619 204 2623 216
rect 2621 192 2623 204
rect 2629 204 2633 216
rect 2629 192 2631 204
rect 2549 70 2573 72
rect 2549 68 2585 70
rect 2549 64 2553 68
rect 2595 64 2599 90
rect 2613 82 2617 192
rect 2651 184 2655 216
rect 2622 180 2655 184
rect 2622 116 2626 180
rect 2642 131 2646 160
rect 2661 158 2665 216
rect 2681 159 2685 196
rect 2642 123 2651 131
rect 2622 104 2625 116
rect 2615 64 2619 70
rect 2627 64 2631 104
rect 2647 64 2651 123
rect 2661 64 2665 146
rect 2681 104 2685 147
rect 2731 128 2735 196
rect 2753 167 2757 216
rect 2763 195 2767 216
rect 2783 204 2787 216
rect 2791 212 2795 216
rect 2791 208 2825 212
rect 2783 200 2813 204
rect 2783 199 2801 200
rect 2763 191 2787 195
rect 2731 116 2733 128
rect 2731 104 2735 116
rect 2753 109 2757 155
rect 2749 103 2757 109
rect 2749 74 2753 103
rect 2781 96 2787 191
rect 2749 67 2757 74
rect 2753 44 2757 67
rect 2761 44 2765 84
rect 2781 64 2785 96
rect 2821 82 2825 208
rect 2837 102 2841 216
rect 2859 204 2863 216
rect 2861 192 2863 204
rect 2869 204 2873 216
rect 2869 192 2871 204
rect 2789 70 2813 72
rect 2789 68 2825 70
rect 2789 64 2793 68
rect 2835 64 2839 90
rect 2853 82 2857 192
rect 2891 184 2895 216
rect 2862 180 2895 184
rect 2862 116 2866 180
rect 2882 131 2886 160
rect 2901 158 2905 216
rect 3125 209 3129 216
rect 3145 209 3149 216
rect 3125 203 3139 209
rect 3145 204 3158 209
rect 2921 159 2925 196
rect 2971 189 2975 196
rect 2960 185 2975 189
rect 2882 123 2891 131
rect 2862 104 2865 116
rect 2855 64 2859 70
rect 2867 64 2871 104
rect 2887 64 2891 123
rect 2901 64 2905 146
rect 2921 104 2925 147
rect 2960 139 2966 185
rect 2991 173 2995 196
rect 3011 173 3015 196
rect 2986 161 2995 173
rect 2961 112 2966 127
rect 2989 112 2995 161
rect 2961 108 2975 112
rect 2971 104 2975 108
rect 2981 108 2995 112
rect 2981 104 2985 108
rect 3011 104 3015 161
rect 3031 139 3035 196
rect 3105 188 3109 196
rect 3105 176 3115 188
rect 3135 139 3139 203
rect 3154 159 3158 204
rect 3191 191 3195 196
rect 3182 184 3195 191
rect 3031 127 3033 139
rect 3031 112 3035 127
rect 3021 108 3035 112
rect 3021 104 3025 108
rect 3115 104 3119 109
rect 3135 104 3139 127
rect 3154 113 3158 147
rect 3182 139 3186 184
rect 3211 173 3215 196
rect 3206 161 3215 173
rect 3145 108 3158 113
rect 3182 116 3186 127
rect 3182 108 3200 116
rect 3145 104 3149 108
rect 3196 104 3200 108
rect 3204 104 3208 161
rect 3231 119 3235 196
rect 3305 159 3309 216
rect 3353 176 3357 196
rect 3349 169 3357 176
rect 3363 176 3367 196
rect 3363 169 3377 176
rect 3305 147 3314 159
rect 3349 153 3355 169
rect 3226 107 3233 119
rect 3226 64 3230 107
rect 3305 64 3309 147
rect 3346 141 3355 153
rect 3351 64 3355 141
rect 3371 153 3377 169
rect 3371 141 3374 153
rect 3371 64 3375 141
rect 3468 119 3472 176
rect 3445 107 3453 119
rect 3465 107 3472 119
rect 3445 64 3449 107
rect 3476 99 3480 176
rect 3484 119 3488 176
rect 3545 159 3549 216
rect 3612 173 3616 216
rect 3605 161 3614 173
rect 3545 147 3554 159
rect 3484 107 3494 119
rect 3474 80 3480 87
rect 3465 76 3480 80
rect 3494 76 3500 107
rect 3465 64 3469 76
rect 3485 72 3500 76
rect 3485 64 3489 72
rect 3545 64 3549 147
rect 3605 104 3609 161
rect 3634 159 3638 196
rect 3642 192 3646 196
rect 3642 186 3661 192
rect 3654 173 3661 186
rect 3634 124 3640 147
rect 3654 124 3661 161
rect 3705 139 3709 216
rect 3725 139 3729 216
rect 3771 159 3775 216
rect 3831 191 3835 196
rect 3766 147 3775 159
rect 3706 127 3721 139
rect 3625 118 3640 124
rect 3645 118 3661 124
rect 3625 104 3629 118
rect 3645 104 3649 118
rect 3717 104 3721 127
rect 3725 127 3734 139
rect 3725 104 3729 127
rect 3771 64 3775 147
rect 3822 184 3835 191
rect 3822 139 3826 184
rect 3851 173 3855 196
rect 3846 161 3855 173
rect 3822 116 3826 127
rect 3822 108 3840 116
rect 3836 104 3840 108
rect 3844 104 3848 161
rect 3871 119 3875 196
rect 3931 139 3935 216
rect 3951 139 3955 216
rect 4113 176 4117 196
rect 3926 127 3935 139
rect 3866 107 3873 119
rect 3866 64 3870 107
rect 3931 104 3935 127
rect 3939 127 3954 139
rect 3939 104 3943 127
rect 4048 119 4052 176
rect 4025 107 4033 119
rect 4045 107 4052 119
rect 4025 64 4029 107
rect 4056 99 4060 176
rect 4064 119 4068 176
rect 4109 169 4117 176
rect 4123 176 4127 196
rect 4313 176 4317 196
rect 4123 169 4137 176
rect 4109 153 4115 169
rect 4106 141 4115 153
rect 4064 107 4074 119
rect 4054 80 4060 87
rect 4045 76 4060 80
rect 4074 76 4080 107
rect 4045 64 4049 76
rect 4065 72 4080 76
rect 4065 64 4069 72
rect 4111 64 4115 141
rect 4131 153 4137 169
rect 4131 141 4134 153
rect 4131 64 4135 141
rect 4228 119 4232 176
rect 4205 107 4213 119
rect 4225 107 4232 119
rect 4205 64 4209 107
rect 4236 99 4240 176
rect 4244 119 4248 176
rect 4303 169 4317 176
rect 4323 176 4327 196
rect 4473 176 4477 196
rect 4323 169 4331 176
rect 4303 153 4309 169
rect 4306 141 4309 153
rect 4244 107 4254 119
rect 4234 80 4240 87
rect 4225 76 4240 80
rect 4254 76 4260 107
rect 4225 64 4229 76
rect 4245 72 4260 76
rect 4245 64 4249 72
rect 4305 64 4309 141
rect 4325 153 4331 169
rect 4325 141 4334 153
rect 4325 64 4329 141
rect 4408 119 4412 176
rect 4385 107 4393 119
rect 4405 107 4412 119
rect 4385 64 4389 107
rect 4416 99 4420 176
rect 4424 119 4428 176
rect 4469 169 4477 176
rect 4483 176 4487 196
rect 4483 169 4497 176
rect 4469 153 4475 169
rect 4466 141 4475 153
rect 4424 107 4434 119
rect 4414 80 4420 87
rect 4405 76 4420 80
rect 4434 76 4440 107
rect 4405 64 4409 76
rect 4425 72 4440 76
rect 4425 64 4429 72
rect 4471 64 4475 141
rect 4491 153 4497 169
rect 4491 141 4494 153
rect 4491 64 4495 141
rect 4552 119 4556 176
rect 4546 107 4556 119
rect 4540 76 4546 107
rect 4560 99 4564 176
rect 4568 119 4572 176
rect 4672 173 4676 216
rect 4665 161 4674 173
rect 4568 107 4575 119
rect 4587 107 4595 119
rect 4560 80 4566 87
rect 4560 76 4575 80
rect 4540 72 4555 76
rect 4551 64 4555 72
rect 4571 64 4575 76
rect 4591 64 4595 107
rect 4665 104 4669 161
rect 4694 159 4698 196
rect 4702 192 4706 196
rect 4702 186 4721 192
rect 4714 173 4721 186
rect 4694 124 4700 147
rect 4714 124 4721 161
rect 4685 118 4700 124
rect 4705 118 4721 124
rect 4685 104 4689 118
rect 4705 104 4709 118
rect 35 20 39 24
rect 55 20 59 24
rect 69 20 73 24
rect 89 20 93 24
rect 101 20 105 24
rect 121 20 125 24
rect 167 20 171 24
rect 175 20 179 24
rect 195 20 199 24
rect 203 20 207 24
rect 225 20 229 24
rect 271 20 275 24
rect 291 20 295 24
rect 311 20 315 24
rect 331 20 335 24
rect 391 20 395 24
rect 399 20 403 24
rect 471 20 475 24
rect 491 20 495 24
rect 511 20 515 24
rect 595 20 599 24
rect 615 20 619 24
rect 625 20 629 24
rect 685 20 689 24
rect 705 20 709 24
rect 725 20 729 24
rect 771 20 775 24
rect 793 20 797 24
rect 801 20 805 24
rect 821 20 825 24
rect 829 20 833 24
rect 875 20 879 24
rect 895 20 899 24
rect 907 20 911 24
rect 927 20 931 24
rect 941 20 945 24
rect 961 20 965 24
rect 1030 20 1034 24
rect 1052 20 1056 24
rect 1060 20 1064 24
rect 1125 20 1129 24
rect 1197 20 1201 24
rect 1205 20 1209 24
rect 1265 20 1269 24
rect 1330 20 1334 24
rect 1352 20 1356 24
rect 1360 20 1364 24
rect 1425 20 1429 24
rect 1485 20 1489 24
rect 1531 20 1535 24
rect 1539 20 1543 24
rect 1625 20 1629 24
rect 1645 20 1649 24
rect 1665 20 1669 24
rect 1715 20 1719 24
rect 1735 20 1739 24
rect 1749 20 1753 24
rect 1769 20 1773 24
rect 1781 20 1785 24
rect 1801 20 1805 24
rect 1847 20 1851 24
rect 1855 20 1859 24
rect 1875 20 1879 24
rect 1883 20 1887 24
rect 1905 20 1909 24
rect 1970 20 1974 24
rect 1992 20 1996 24
rect 2000 20 2004 24
rect 2051 20 2055 24
rect 2111 20 2115 24
rect 2119 20 2123 24
rect 2191 20 2195 24
rect 2199 20 2203 24
rect 2297 20 2301 24
rect 2305 20 2309 24
rect 2351 20 2355 24
rect 2359 20 2363 24
rect 2445 20 2449 24
rect 2491 20 2495 24
rect 2513 20 2517 24
rect 2521 20 2525 24
rect 2541 20 2545 24
rect 2549 20 2553 24
rect 2595 20 2599 24
rect 2615 20 2619 24
rect 2627 20 2631 24
rect 2647 20 2651 24
rect 2661 20 2665 24
rect 2681 20 2685 24
rect 2731 20 2735 24
rect 2753 20 2757 24
rect 2761 20 2765 24
rect 2781 20 2785 24
rect 2789 20 2793 24
rect 2835 20 2839 24
rect 2855 20 2859 24
rect 2867 20 2871 24
rect 2887 20 2891 24
rect 2901 20 2905 24
rect 2921 20 2925 24
rect 2971 20 2975 24
rect 2981 20 2985 24
rect 3011 20 3015 24
rect 3021 20 3025 24
rect 3115 20 3119 24
rect 3135 20 3139 24
rect 3145 20 3149 24
rect 3196 20 3200 24
rect 3204 20 3208 24
rect 3226 20 3230 24
rect 3305 20 3309 24
rect 3351 20 3355 24
rect 3371 20 3375 24
rect 3445 20 3449 24
rect 3465 20 3469 24
rect 3485 20 3489 24
rect 3545 20 3549 24
rect 3605 20 3609 24
rect 3625 20 3629 24
rect 3645 20 3649 24
rect 3717 20 3721 24
rect 3725 20 3729 24
rect 3771 20 3775 24
rect 3836 20 3840 24
rect 3844 20 3848 24
rect 3866 20 3870 24
rect 3931 20 3935 24
rect 3939 20 3943 24
rect 4025 20 4029 24
rect 4045 20 4049 24
rect 4065 20 4069 24
rect 4111 20 4115 24
rect 4131 20 4135 24
rect 4205 20 4209 24
rect 4225 20 4229 24
rect 4245 20 4249 24
rect 4305 20 4309 24
rect 4325 20 4329 24
rect 4385 20 4389 24
rect 4405 20 4409 24
rect 4425 20 4429 24
rect 4471 20 4475 24
rect 4491 20 4495 24
rect 4551 20 4555 24
rect 4571 20 4575 24
rect 4591 20 4595 24
rect 4665 20 4669 24
rect 4685 20 4689 24
rect 4705 20 4709 24
<< polycontact >>
rect 45 4498 57 4510
rect 114 4461 126 4473
rect 74 4447 86 4459
rect 45 4430 57 4442
rect 154 4461 166 4473
rect 234 4481 246 4493
rect 195 4427 207 4439
rect 303 4498 315 4510
rect 543 4498 555 4510
rect 254 4447 266 4459
rect 274 4447 286 4459
rect 374 4447 386 4459
rect 303 4430 315 4442
rect 414 4447 426 4459
rect 454 4447 466 4459
rect 494 4447 506 4459
rect 514 4447 526 4459
rect 634 4467 646 4479
rect 543 4430 555 4442
rect 734 4467 746 4479
rect 654 4447 666 4459
rect 694 4447 706 4459
rect 827 4475 839 4487
rect 813 4436 825 4448
rect 881 4508 893 4520
rect 841 4404 853 4416
rect 865 4404 877 4416
rect 929 4512 941 4524
rect 951 4512 963 4524
rect 913 4410 925 4422
rect 893 4390 905 4402
rect 954 4480 966 4492
rect 974 4466 986 4478
rect 994 4467 1006 4479
rect 945 4424 957 4436
rect 927 4390 939 4402
rect 1054 4481 1066 4493
rect 1034 4447 1046 4459
rect 1167 4475 1179 4487
rect 1093 4427 1105 4439
rect 1153 4436 1165 4448
rect 1221 4508 1233 4520
rect 1181 4404 1193 4416
rect 1205 4404 1217 4416
rect 1269 4512 1281 4524
rect 1291 4512 1303 4524
rect 1253 4410 1265 4422
rect 1233 4390 1245 4402
rect 1294 4480 1306 4492
rect 1314 4466 1326 4478
rect 1334 4467 1346 4479
rect 1285 4424 1297 4436
rect 1267 4390 1279 4402
rect 1394 4481 1406 4493
rect 1374 4447 1386 4459
rect 1494 4467 1506 4479
rect 1537 4512 1549 4524
rect 1559 4512 1571 4524
rect 1534 4480 1546 4492
rect 1433 4427 1445 4439
rect 1514 4466 1526 4478
rect 1543 4424 1555 4436
rect 1575 4410 1587 4422
rect 1561 4390 1573 4402
rect 1607 4508 1619 4520
rect 1661 4475 1673 4487
rect 1714 4461 1726 4473
rect 1675 4436 1687 4448
rect 1623 4404 1635 4416
rect 1595 4390 1607 4402
rect 1647 4404 1659 4416
rect 1754 4461 1766 4473
rect 1827 4475 1839 4487
rect 1813 4436 1825 4448
rect 1881 4508 1893 4520
rect 1841 4404 1853 4416
rect 1865 4404 1877 4416
rect 1929 4512 1941 4524
rect 1951 4512 1963 4524
rect 1913 4410 1925 4422
rect 1893 4390 1905 4402
rect 1954 4480 1966 4492
rect 1974 4466 1986 4478
rect 1994 4467 2006 4479
rect 1945 4424 1957 4436
rect 1927 4390 1939 4402
rect 2054 4481 2066 4493
rect 2090 4481 2102 4493
rect 2034 4447 2046 4459
rect 2113 4447 2125 4459
rect 2193 4427 2205 4439
rect 2314 4481 2326 4493
rect 2234 4427 2246 4439
rect 2275 4427 2287 4439
rect 2214 4407 2226 4419
rect 2394 4467 2406 4479
rect 2334 4447 2346 4459
rect 2534 4467 2546 4479
rect 2414 4447 2426 4459
rect 2454 4447 2466 4459
rect 2574 4481 2586 4493
rect 2554 4447 2566 4459
rect 2683 4498 2695 4510
rect 2763 4498 2775 4510
rect 2845 4498 2857 4510
rect 2654 4447 2666 4459
rect 2734 4447 2746 4459
rect 2613 4427 2625 4439
rect 2683 4430 2695 4442
rect 3033 4498 3045 4510
rect 2874 4447 2886 4459
rect 2763 4430 2775 4442
rect 2845 4430 2857 4442
rect 2933 4427 2945 4439
rect 2974 4427 2986 4439
rect 2954 4407 2966 4419
rect 3034 4461 3046 4473
rect 3125 4498 3137 4510
rect 3074 4447 3086 4459
rect 3154 4447 3166 4459
rect 3125 4430 3137 4442
rect 3213 4427 3225 4439
rect 3274 4461 3286 4473
rect 3254 4427 3266 4439
rect 3234 4407 3246 4419
rect 3354 4481 3366 4493
rect 3314 4461 3326 4473
rect 3394 4481 3406 4493
rect 3374 4467 3386 4479
rect 3454 4467 3466 4479
rect 3514 4461 3526 4473
rect 3554 4461 3566 4473
rect 3594 4427 3606 4439
rect 3694 4481 3706 4493
rect 3734 4481 3746 4493
rect 3714 4467 3726 4479
rect 3635 4427 3647 4439
rect 3614 4407 3626 4419
rect 3814 4481 3826 4493
rect 3794 4447 3806 4459
rect 3954 4481 3966 4493
rect 3853 4427 3865 4439
rect 3915 4427 3927 4439
rect 3974 4447 3986 4459
rect 4033 4427 4045 4439
rect 4074 4427 4086 4439
rect 4133 4427 4145 4439
rect 4054 4407 4066 4419
rect 4194 4481 4206 4493
rect 4234 4481 4246 4493
rect 4214 4467 4226 4479
rect 4174 4427 4186 4439
rect 4154 4407 4166 4419
rect 4294 4461 4306 4473
rect 4414 4481 4426 4493
rect 4334 4461 4346 4473
rect 4454 4481 4466 4493
rect 4434 4467 4446 4479
rect 4514 4467 4526 4479
rect 4534 4427 4546 4439
rect 4575 4427 4587 4439
rect 4634 4427 4646 4439
rect 4554 4407 4566 4419
rect 4675 4427 4687 4439
rect 4654 4407 4666 4419
rect 35 4221 47 4233
rect 94 4201 106 4213
rect 74 4167 86 4179
rect 194 4201 206 4213
rect 214 4201 226 4213
rect 254 4201 266 4213
rect 154 4187 166 4199
rect 153 4150 165 4162
rect 354 4181 366 4193
rect 334 4167 346 4179
rect 394 4201 406 4213
rect 374 4167 386 4179
rect 434 4187 446 4199
rect 614 4241 626 4253
rect 594 4221 606 4233
rect 554 4181 566 4193
rect 534 4167 546 4179
rect 435 4150 447 4162
rect 574 4167 586 4179
rect 635 4221 647 4233
rect 714 4181 726 4193
rect 694 4167 706 4179
rect 794 4201 806 4213
rect 734 4167 746 4179
rect 834 4187 846 4199
rect 915 4221 927 4233
rect 835 4150 847 4162
rect 974 4201 986 4213
rect 954 4167 966 4179
rect 1054 4201 1066 4213
rect 1094 4201 1106 4213
rect 1134 4201 1146 4213
rect 1174 4201 1186 4213
rect 1214 4201 1226 4213
rect 1254 4201 1266 4213
rect 1034 4181 1046 4193
rect 1401 4244 1413 4256
rect 1453 4258 1465 4270
rect 1425 4244 1437 4256
rect 1294 4181 1306 4193
rect 1373 4212 1385 4224
rect 1387 4173 1399 4185
rect 1441 4140 1453 4152
rect 1487 4258 1499 4270
rect 1473 4238 1485 4250
rect 1505 4224 1517 4236
rect 1534 4182 1546 4194
rect 1594 4201 1606 4213
rect 1514 4168 1526 4180
rect 1489 4136 1501 4148
rect 1511 4136 1523 4148
rect 1554 4181 1566 4193
rect 1653 4221 1665 4233
rect 1614 4167 1626 4179
rect 1694 4201 1706 4213
rect 1734 4201 1746 4213
rect 1881 4244 1893 4256
rect 1933 4258 1945 4270
rect 1905 4244 1917 4256
rect 1853 4212 1865 4224
rect 1814 4181 1826 4193
rect 1867 4173 1879 4185
rect 1921 4140 1933 4152
rect 1967 4258 1979 4270
rect 1953 4238 1965 4250
rect 1985 4224 1997 4236
rect 2014 4182 2026 4194
rect 1994 4168 2006 4180
rect 1969 4136 1981 4148
rect 1991 4136 2003 4148
rect 2034 4181 2046 4193
rect 2094 4187 2106 4199
rect 2134 4187 2146 4199
rect 2193 4219 2205 4231
rect 2174 4201 2186 4213
rect 2274 4201 2286 4213
rect 2154 4181 2166 4193
rect 2193 4152 2205 4164
rect 2353 4201 2365 4213
rect 2295 4167 2307 4179
rect 2333 4167 2345 4179
rect 2374 4187 2386 4199
rect 2475 4221 2487 4233
rect 2414 4187 2426 4199
rect 2534 4201 2546 4213
rect 2574 4201 2586 4213
rect 2614 4201 2626 4213
rect 2514 4167 2526 4179
rect 2654 4181 2666 4193
rect 2634 4167 2646 4179
rect 2674 4167 2686 4179
rect 2794 4181 2806 4193
rect 2774 4167 2786 4179
rect 2863 4218 2875 4230
rect 2974 4241 2986 4253
rect 2953 4221 2965 4233
rect 2834 4201 2846 4213
rect 2814 4167 2826 4179
rect 3074 4241 3086 4253
rect 2994 4221 3006 4233
rect 3053 4221 3065 4233
rect 3094 4221 3106 4233
rect 3114 4187 3126 4199
rect 3154 4187 3166 4199
rect 3314 4241 3326 4253
rect 3293 4221 3305 4233
rect 2863 4150 2875 4162
rect 3234 4181 3246 4193
rect 3414 4241 3426 4253
rect 3334 4221 3346 4233
rect 3393 4221 3405 4233
rect 3514 4241 3526 4253
rect 3434 4221 3446 4233
rect 3493 4221 3505 4233
rect 3614 4241 3626 4253
rect 3534 4221 3546 4233
rect 3593 4221 3605 4233
rect 3674 4241 3686 4253
rect 3634 4221 3646 4233
rect 3654 4221 3666 4233
rect 3695 4221 3707 4233
rect 3774 4181 3786 4193
rect 3754 4167 3766 4179
rect 3854 4201 3866 4213
rect 3794 4167 3806 4179
rect 3913 4221 3925 4233
rect 3874 4167 3886 4179
rect 3954 4181 3966 4193
rect 4034 4181 4046 4193
rect 4014 4167 4026 4179
rect 4174 4241 4186 4253
rect 4153 4221 4165 4233
rect 4054 4167 4066 4179
rect 4234 4241 4246 4253
rect 4194 4221 4206 4233
rect 4214 4221 4226 4233
rect 4255 4221 4267 4233
rect 4334 4181 4346 4193
rect 4314 4167 4326 4179
rect 4414 4201 4426 4213
rect 4354 4167 4366 4179
rect 4473 4221 4485 4233
rect 4434 4167 4446 4179
rect 4515 4201 4527 4213
rect 4594 4201 4606 4213
rect 4654 4201 4666 4213
rect 4694 4201 4706 4213
rect 4535 4167 4547 4179
rect 4573 4167 4585 4179
rect 34 3981 46 3993
rect 74 3981 86 3993
rect 114 3981 126 3993
rect 154 3981 166 3993
rect 274 4001 286 4013
rect 194 3967 206 3979
rect 234 3967 246 3979
rect 254 3967 266 3979
rect 394 3987 406 3999
rect 454 3987 466 3999
rect 313 3947 325 3959
rect 595 4018 607 4030
rect 594 3981 606 3993
rect 494 3967 506 3979
rect 534 3967 546 3979
rect 554 3967 566 3979
rect 674 4001 686 4013
rect 654 3967 666 3979
rect 754 3987 766 3999
rect 713 3947 725 3959
rect 834 4001 846 4013
rect 814 3967 826 3979
rect 914 3981 926 3993
rect 873 3947 885 3959
rect 954 3981 966 3993
rect 1034 3987 1046 3999
rect 1134 3987 1146 3999
rect 1074 3967 1086 3979
rect 1114 3967 1126 3979
rect 1274 3987 1286 3999
rect 1194 3967 1206 3979
rect 1234 3967 1246 3979
rect 1454 3987 1466 3999
rect 1354 3967 1366 3979
rect 1394 3967 1406 3979
rect 1494 4001 1506 4013
rect 1474 3967 1486 3979
rect 1594 4001 1606 4013
rect 1630 4001 1642 4013
rect 1574 3967 1586 3979
rect 1533 3947 1545 3959
rect 1694 3981 1706 3993
rect 1653 3967 1665 3979
rect 1814 4001 1826 4013
rect 1734 3981 1746 3993
rect 1854 4001 1866 4013
rect 1834 3987 1846 3999
rect 1874 3947 1886 3959
rect 2034 4001 2046 4013
rect 1915 3947 1927 3959
rect 1995 3947 2007 3959
rect 1894 3927 1906 3939
rect 2114 3987 2126 3999
rect 2054 3967 2066 3979
rect 2173 3947 2185 3959
rect 2214 3947 2226 3959
rect 2273 3947 2285 3959
rect 2194 3927 2206 3939
rect 2374 4001 2386 4013
rect 2314 3947 2326 3959
rect 2294 3927 2306 3939
rect 2414 4001 2426 4013
rect 2394 3987 2406 3999
rect 2474 3987 2486 3999
rect 2554 4001 2566 4013
rect 2515 3947 2527 3959
rect 2574 3967 2586 3979
rect 2633 3947 2645 3959
rect 2734 4001 2746 4013
rect 2674 3947 2686 3959
rect 2654 3927 2666 3939
rect 2774 4001 2786 4013
rect 2754 3987 2766 3999
rect 2854 4001 2866 4013
rect 2815 3947 2827 3959
rect 2914 4001 2926 4013
rect 2874 3967 2886 3979
rect 2894 3967 2906 3979
rect 2953 3947 2965 3959
rect 3033 3947 3045 3959
rect 3134 3987 3146 3999
rect 3074 3947 3086 3959
rect 3054 3927 3066 3939
rect 3174 4001 3186 4013
rect 3154 3967 3166 3979
rect 3254 4001 3266 4013
rect 3294 4001 3306 4013
rect 3274 3987 3286 3999
rect 3213 3947 3225 3959
rect 3374 4001 3386 4013
rect 3354 3967 3366 3979
rect 3514 4001 3526 4013
rect 3413 3947 3425 3959
rect 3475 3947 3487 3959
rect 3534 3967 3546 3979
rect 3614 4001 3626 4013
rect 3575 3947 3587 3959
rect 3694 4001 3706 4013
rect 3634 3967 3646 3979
rect 3734 4001 3746 4013
rect 3714 3987 3726 3999
rect 3793 3947 3805 3959
rect 3874 3981 3886 3993
rect 3834 3947 3846 3959
rect 3814 3927 3826 3939
rect 3914 3981 3926 3993
rect 3954 3981 3966 3993
rect 3994 3981 4006 3993
rect 4014 3981 4026 3993
rect 4054 3981 4066 3993
rect 4133 3947 4145 3959
rect 4254 4001 4266 4013
rect 4174 3947 4186 3959
rect 4215 3947 4227 3959
rect 4154 3927 4166 3939
rect 4314 4001 4326 4013
rect 4274 3967 4286 3979
rect 4294 3967 4306 3979
rect 4434 3987 4446 3999
rect 4353 3947 4365 3959
rect 4493 3947 4505 3959
rect 4534 3947 4546 3959
rect 4593 3947 4605 3959
rect 4514 3927 4526 3939
rect 4654 4001 4666 4013
rect 4694 4001 4706 4013
rect 4674 3987 4686 3999
rect 4634 3947 4646 3959
rect 4614 3927 4626 3939
rect 35 3741 47 3753
rect 94 3721 106 3733
rect 74 3687 86 3699
rect 221 3764 233 3776
rect 273 3778 285 3790
rect 245 3764 257 3776
rect 193 3732 205 3744
rect 154 3701 166 3713
rect 207 3693 219 3705
rect 261 3660 273 3672
rect 307 3778 319 3790
rect 293 3758 305 3770
rect 325 3744 337 3756
rect 354 3702 366 3714
rect 435 3741 447 3753
rect 334 3688 346 3700
rect 309 3656 321 3668
rect 331 3656 343 3668
rect 374 3701 386 3713
rect 494 3721 506 3733
rect 514 3721 526 3733
rect 474 3687 486 3699
rect 554 3707 566 3719
rect 655 3739 667 3751
rect 674 3721 686 3733
rect 555 3670 567 3682
rect 655 3672 667 3684
rect 694 3701 706 3713
rect 734 3707 746 3719
rect 774 3707 786 3719
rect 881 3778 893 3790
rect 863 3744 875 3756
rect 814 3701 826 3713
rect 834 3702 846 3714
rect 854 3688 866 3700
rect 915 3778 927 3790
rect 895 3758 907 3770
rect 857 3656 869 3668
rect 879 3656 891 3668
rect 943 3764 955 3776
rect 967 3764 979 3776
rect 927 3660 939 3672
rect 995 3732 1007 3744
rect 1065 3738 1077 3750
rect 981 3693 993 3705
rect 1161 3764 1173 3776
rect 1213 3778 1225 3790
rect 1185 3764 1197 3776
rect 1094 3721 1106 3733
rect 1133 3732 1145 3744
rect 1065 3670 1077 3682
rect 1147 3693 1159 3705
rect 1201 3660 1213 3672
rect 1247 3778 1259 3790
rect 1233 3758 1245 3770
rect 1265 3744 1277 3756
rect 1294 3702 1306 3714
rect 1354 3721 1366 3733
rect 1274 3688 1286 3700
rect 1249 3656 1261 3668
rect 1271 3656 1283 3668
rect 1314 3701 1326 3713
rect 1413 3741 1425 3753
rect 1374 3687 1386 3699
rect 1454 3707 1466 3719
rect 1494 3707 1506 3719
rect 1534 3707 1546 3719
rect 1741 3764 1753 3776
rect 1793 3778 1805 3790
rect 1765 3764 1777 3776
rect 1643 3738 1655 3750
rect 1614 3721 1626 3733
rect 1574 3707 1586 3719
rect 1713 3732 1725 3744
rect 1643 3670 1655 3682
rect 1727 3693 1739 3705
rect 1781 3660 1793 3672
rect 1827 3778 1839 3790
rect 1813 3758 1825 3770
rect 1845 3744 1857 3756
rect 1874 3702 1886 3714
rect 1854 3688 1866 3700
rect 1829 3656 1841 3668
rect 1851 3656 1863 3668
rect 1894 3701 1906 3713
rect 1974 3701 1986 3713
rect 2054 3701 2066 3713
rect 2034 3687 2046 3699
rect 2174 3761 2186 3773
rect 2154 3741 2166 3753
rect 2134 3701 2146 3713
rect 2074 3687 2086 3699
rect 2195 3741 2207 3753
rect 2275 3741 2287 3753
rect 2414 3761 2426 3773
rect 2393 3741 2405 3753
rect 2334 3721 2346 3733
rect 2314 3687 2326 3699
rect 2434 3741 2446 3753
rect 2614 3761 2626 3773
rect 2593 3741 2605 3753
rect 2514 3701 2526 3713
rect 2494 3687 2506 3699
rect 2534 3687 2546 3699
rect 2634 3741 2646 3753
rect 2674 3701 2686 3713
rect 2654 3687 2666 3699
rect 2694 3687 2706 3699
rect 2814 3701 2826 3713
rect 2794 3687 2806 3699
rect 3034 3761 3046 3773
rect 3013 3741 3025 3753
rect 2894 3701 2906 3713
rect 2954 3701 2966 3713
rect 2834 3687 2846 3699
rect 3054 3741 3066 3753
rect 3234 3761 3246 3773
rect 3213 3741 3225 3753
rect 3134 3701 3146 3713
rect 3114 3687 3126 3699
rect 3154 3687 3166 3699
rect 3254 3741 3266 3753
rect 3355 3741 3367 3753
rect 3314 3701 3326 3713
rect 3414 3721 3426 3733
rect 3394 3687 3406 3699
rect 3454 3707 3466 3719
rect 3514 3721 3526 3733
rect 3494 3707 3506 3719
rect 3554 3707 3566 3719
rect 3774 3761 3786 3773
rect 3753 3741 3765 3753
rect 3674 3701 3686 3713
rect 3654 3687 3666 3699
rect 3555 3670 3567 3682
rect 3694 3687 3706 3699
rect 3794 3741 3806 3753
rect 3854 3701 3866 3713
rect 3894 3701 3906 3713
rect 3874 3687 3886 3699
rect 3995 3741 4007 3753
rect 3914 3687 3926 3699
rect 4054 3721 4066 3733
rect 4074 3721 4086 3733
rect 4034 3687 4046 3699
rect 4133 3741 4145 3753
rect 4094 3687 4106 3699
rect 4194 3701 4206 3713
rect 4174 3687 4186 3699
rect 4214 3687 4226 3699
rect 4394 3761 4406 3773
rect 4374 3741 4386 3753
rect 4334 3701 4346 3713
rect 4314 3687 4326 3699
rect 4354 3687 4366 3699
rect 4415 3741 4427 3753
rect 4594 3761 4606 3773
rect 4573 3741 4585 3753
rect 4514 3701 4526 3713
rect 4654 3761 4666 3773
rect 4614 3741 4626 3753
rect 4634 3741 4646 3753
rect 4675 3741 4687 3753
rect 34 3507 46 3519
rect 77 3552 89 3564
rect 99 3552 111 3564
rect 74 3520 86 3532
rect 54 3506 66 3518
rect 83 3464 95 3476
rect 115 3450 127 3462
rect 101 3430 113 3442
rect 147 3548 159 3560
rect 201 3515 213 3527
rect 274 3501 286 3513
rect 215 3476 227 3488
rect 163 3444 175 3456
rect 135 3430 147 3442
rect 187 3444 199 3456
rect 314 3501 326 3513
rect 394 3521 406 3533
rect 355 3467 367 3479
rect 454 3501 466 3513
rect 414 3487 426 3499
rect 494 3501 506 3513
rect 553 3467 565 3479
rect 654 3507 666 3519
rect 594 3467 606 3479
rect 574 3447 586 3459
rect 734 3521 746 3533
rect 695 3467 707 3479
rect 754 3487 766 3499
rect 834 3521 846 3533
rect 795 3467 807 3479
rect 874 3507 886 3519
rect 854 3487 866 3499
rect 954 3487 966 3499
rect 994 3487 1006 3499
rect 1047 3515 1059 3527
rect 1033 3476 1045 3488
rect 1101 3548 1113 3560
rect 1061 3444 1073 3456
rect 1085 3444 1097 3456
rect 1149 3552 1161 3564
rect 1171 3552 1183 3564
rect 1133 3450 1145 3462
rect 1113 3430 1125 3442
rect 1174 3520 1186 3532
rect 1194 3506 1206 3518
rect 1214 3507 1226 3519
rect 1254 3507 1266 3519
rect 1165 3464 1177 3476
rect 1147 3430 1159 3442
rect 1414 3521 1426 3533
rect 1314 3487 1326 3499
rect 1354 3487 1366 3499
rect 1394 3487 1406 3499
rect 1605 3538 1617 3550
rect 1494 3501 1506 3513
rect 1453 3467 1465 3479
rect 1534 3501 1546 3513
rect 1694 3507 1706 3519
rect 1634 3487 1646 3499
rect 1605 3470 1617 3482
rect 1747 3515 1759 3527
rect 1733 3476 1745 3488
rect 1801 3548 1813 3560
rect 1761 3444 1773 3456
rect 1785 3444 1797 3456
rect 1849 3552 1861 3564
rect 1871 3552 1883 3564
rect 1833 3450 1845 3462
rect 1813 3430 1825 3442
rect 1874 3520 1886 3532
rect 1894 3506 1906 3518
rect 1914 3507 1926 3519
rect 1865 3464 1877 3476
rect 1847 3430 1859 3442
rect 1974 3521 1986 3533
rect 2010 3521 2022 3533
rect 1954 3487 1966 3499
rect 2074 3501 2086 3513
rect 2033 3487 2045 3499
rect 2194 3521 2206 3533
rect 2114 3501 2126 3513
rect 2234 3521 2246 3533
rect 2214 3507 2226 3519
rect 2293 3467 2305 3479
rect 2394 3507 2406 3519
rect 2334 3467 2346 3479
rect 2314 3447 2326 3459
rect 2453 3467 2465 3479
rect 2494 3467 2506 3479
rect 2553 3467 2565 3479
rect 2474 3447 2486 3459
rect 2674 3521 2686 3533
rect 2594 3467 2606 3479
rect 2635 3467 2647 3479
rect 2574 3447 2586 3459
rect 2734 3521 2746 3533
rect 2694 3487 2706 3499
rect 2714 3487 2726 3499
rect 2814 3501 2826 3513
rect 2773 3467 2785 3479
rect 2854 3501 2866 3513
rect 2914 3521 2926 3533
rect 2894 3487 2906 3499
rect 2994 3487 3006 3499
rect 2953 3467 2965 3479
rect 3034 3487 3046 3499
rect 3134 3521 3146 3533
rect 3095 3467 3107 3479
rect 3195 3521 3207 3533
rect 3233 3521 3245 3533
rect 3154 3487 3166 3499
rect 3175 3487 3187 3499
rect 3294 3501 3306 3513
rect 3254 3487 3266 3499
rect 3334 3501 3346 3513
rect 3374 3501 3386 3513
rect 3414 3501 3426 3513
rect 3454 3501 3466 3513
rect 3494 3501 3506 3513
rect 3614 3501 3626 3513
rect 3534 3487 3546 3499
rect 3574 3487 3586 3499
rect 3654 3501 3666 3513
rect 3694 3501 3706 3513
rect 3734 3501 3746 3513
rect 3794 3501 3806 3513
rect 3834 3501 3846 3513
rect 3934 3501 3946 3513
rect 3874 3487 3886 3499
rect 3914 3487 3926 3499
rect 3974 3501 3986 3513
rect 4014 3501 4026 3513
rect 4054 3501 4066 3513
rect 4114 3521 4126 3533
rect 4094 3487 4106 3499
rect 4153 3467 4165 3479
rect 4233 3467 4245 3479
rect 4274 3467 4286 3479
rect 4294 3467 4306 3479
rect 4254 3447 4266 3459
rect 4394 3521 4406 3533
rect 4434 3521 4446 3533
rect 4414 3507 4426 3519
rect 4335 3467 4347 3479
rect 4314 3447 4326 3459
rect 4494 3507 4506 3519
rect 4593 3467 4605 3479
rect 4634 3467 4646 3479
rect 4654 3467 4666 3479
rect 4614 3447 4626 3459
rect 4695 3467 4707 3479
rect 4674 3447 4686 3459
rect 101 3298 113 3310
rect 83 3264 95 3276
rect 34 3221 46 3233
rect 54 3222 66 3234
rect 74 3208 86 3220
rect 135 3298 147 3310
rect 115 3278 127 3290
rect 77 3176 89 3188
rect 99 3176 111 3188
rect 163 3284 175 3296
rect 187 3284 199 3296
rect 147 3180 159 3192
rect 215 3252 227 3264
rect 201 3213 213 3225
rect 274 3241 286 3253
rect 353 3241 365 3253
rect 295 3207 307 3219
rect 333 3207 345 3219
rect 374 3227 386 3239
rect 454 3241 466 3253
rect 414 3227 426 3239
rect 513 3261 525 3273
rect 474 3207 486 3219
rect 554 3241 566 3253
rect 613 3261 625 3273
rect 574 3207 586 3219
rect 674 3227 686 3239
rect 714 3227 726 3239
rect 734 3221 746 3233
rect 838 3204 850 3216
rect 878 3204 890 3216
rect 918 3204 930 3216
rect 954 3207 966 3219
rect 1014 3207 1026 3219
rect 1050 3204 1062 3216
rect 1090 3204 1102 3216
rect 1130 3204 1142 3216
rect 1301 3284 1313 3296
rect 1353 3298 1365 3310
rect 1325 3284 1337 3296
rect 1273 3252 1285 3264
rect 1234 3221 1246 3233
rect 1287 3213 1299 3225
rect 1341 3180 1353 3192
rect 1387 3298 1399 3310
rect 1373 3278 1385 3290
rect 1405 3264 1417 3276
rect 1434 3222 1446 3234
rect 1494 3241 1506 3253
rect 1414 3208 1426 3220
rect 1389 3176 1401 3188
rect 1411 3176 1423 3188
rect 1454 3221 1466 3233
rect 1553 3261 1565 3273
rect 1615 3261 1627 3273
rect 1514 3207 1526 3219
rect 1715 3261 1727 3273
rect 1674 3241 1686 3253
rect 1654 3207 1666 3219
rect 1774 3241 1786 3253
rect 1754 3207 1766 3219
rect 1875 3261 1887 3273
rect 1834 3221 1846 3233
rect 2101 3284 2113 3296
rect 2153 3298 2165 3310
rect 2125 3284 2137 3296
rect 1975 3261 1987 3273
rect 1934 3241 1946 3253
rect 1914 3207 1926 3219
rect 2034 3241 2046 3253
rect 2073 3252 2085 3264
rect 2014 3207 2026 3219
rect 2087 3213 2099 3225
rect 2141 3180 2153 3192
rect 2187 3298 2199 3310
rect 2173 3278 2185 3290
rect 2205 3264 2217 3276
rect 2234 3222 2246 3234
rect 2474 3281 2486 3293
rect 2453 3261 2465 3273
rect 2214 3208 2226 3220
rect 2189 3176 2201 3188
rect 2211 3176 2223 3188
rect 2254 3221 2266 3233
rect 2334 3221 2346 3233
rect 2394 3221 2406 3233
rect 2494 3261 2506 3273
rect 2534 3221 2546 3233
rect 2514 3207 2526 3219
rect 2554 3207 2566 3219
rect 2695 3261 2707 3273
rect 2654 3221 2666 3233
rect 2754 3241 2766 3253
rect 2774 3241 2786 3253
rect 2814 3241 2826 3253
rect 2854 3241 2866 3253
rect 2734 3207 2746 3219
rect 2913 3261 2925 3273
rect 2874 3207 2886 3219
rect 2954 3227 2966 3239
rect 2994 3227 3006 3239
rect 3034 3227 3046 3239
rect 3074 3227 3086 3239
rect 3274 3281 3286 3293
rect 3253 3261 3265 3273
rect 3174 3221 3186 3233
rect 3154 3207 3166 3219
rect 3194 3207 3206 3219
rect 3294 3261 3306 3273
rect 3335 3261 3347 3273
rect 3394 3241 3406 3253
rect 3374 3207 3386 3219
rect 3494 3241 3506 3253
rect 3454 3227 3466 3239
rect 3453 3190 3465 3202
rect 3514 3227 3526 3239
rect 3554 3227 3566 3239
rect 3674 3241 3686 3253
rect 3714 3241 3726 3253
rect 3634 3227 3646 3239
rect 3633 3190 3645 3202
rect 3793 3241 3805 3253
rect 3735 3207 3747 3219
rect 3773 3207 3785 3219
rect 3834 3227 3846 3239
rect 3894 3241 3906 3253
rect 3874 3227 3886 3239
rect 3953 3261 3965 3273
rect 3914 3207 3926 3219
rect 3994 3227 4006 3239
rect 4034 3227 4046 3239
rect 4154 3241 4166 3253
rect 4114 3227 4126 3239
rect 4113 3190 4125 3202
rect 4174 3227 4186 3239
rect 4254 3241 4266 3253
rect 4214 3227 4226 3239
rect 4294 3227 4306 3239
rect 4374 3221 4386 3233
rect 4354 3207 4366 3219
rect 4295 3190 4307 3202
rect 4454 3241 4466 3253
rect 4394 3207 4406 3219
rect 4513 3261 4525 3273
rect 4474 3207 4486 3219
rect 4554 3241 4566 3253
rect 4714 3281 4726 3293
rect 4613 3261 4625 3273
rect 4693 3261 4705 3273
rect 4574 3207 4586 3219
rect 4734 3261 4746 3273
rect 34 3027 46 3039
rect 77 3072 89 3084
rect 99 3072 111 3084
rect 74 3040 86 3052
rect 54 3026 66 3038
rect 83 2984 95 2996
rect 115 2970 127 2982
rect 101 2950 113 2962
rect 147 3068 159 3080
rect 201 3035 213 3047
rect 215 2996 227 3008
rect 314 3041 326 3053
rect 275 2987 287 2999
rect 163 2964 175 2976
rect 135 2950 147 2962
rect 187 2964 199 2976
rect 374 3021 386 3033
rect 334 3007 346 3019
rect 414 3021 426 3033
rect 467 3035 479 3047
rect 453 2996 465 3008
rect 521 3068 533 3080
rect 481 2964 493 2976
rect 505 2964 517 2976
rect 569 3072 581 3084
rect 591 3072 603 3084
rect 553 2970 565 2982
rect 533 2950 545 2962
rect 594 3040 606 3052
rect 614 3026 626 3038
rect 634 3027 646 3039
rect 694 3027 706 3039
rect 737 3072 749 3084
rect 759 3072 771 3084
rect 734 3040 746 3052
rect 585 2984 597 2996
rect 567 2950 579 2962
rect 714 3026 726 3038
rect 743 2984 755 2996
rect 775 2970 787 2982
rect 761 2950 773 2962
rect 807 3068 819 3080
rect 861 3035 873 3047
rect 914 3027 926 3039
rect 875 2996 887 3008
rect 823 2964 835 2976
rect 795 2950 807 2962
rect 847 2964 859 2976
rect 1074 3021 1086 3033
rect 994 3007 1006 3019
rect 1034 3007 1046 3019
rect 1114 3021 1126 3033
rect 1154 3041 1166 3053
rect 1134 3007 1146 3019
rect 1234 3041 1246 3053
rect 1274 3041 1286 3053
rect 1254 3027 1266 3039
rect 1193 2987 1205 2999
rect 1354 3027 1366 3039
rect 1397 3072 1409 3084
rect 1419 3072 1431 3084
rect 1394 3040 1406 3052
rect 1374 3026 1386 3038
rect 1403 2984 1415 2996
rect 1435 2970 1447 2982
rect 1421 2950 1433 2962
rect 1467 3068 1479 3080
rect 1521 3035 1533 3047
rect 1674 3021 1686 3033
rect 1535 2996 1547 3008
rect 1594 3007 1606 3019
rect 1634 3007 1646 3019
rect 1483 2964 1495 2976
rect 1455 2950 1467 2962
rect 1507 2964 1519 2976
rect 1714 3021 1726 3033
rect 1754 3041 1766 3053
rect 1734 3007 1746 3019
rect 1894 3041 1906 3053
rect 1793 2987 1805 2999
rect 1855 2987 1867 2999
rect 1914 3007 1926 3019
rect 1967 3035 1979 3047
rect 1953 2996 1965 3008
rect 2021 3068 2033 3080
rect 1981 2964 1993 2976
rect 2005 2964 2017 2976
rect 2069 3072 2081 3084
rect 2091 3072 2103 3084
rect 2053 2970 2065 2982
rect 2033 2950 2045 2962
rect 2094 3040 2106 3052
rect 2114 3026 2126 3038
rect 2134 3027 2146 3039
rect 2085 2984 2097 2996
rect 2067 2950 2079 2962
rect 2294 3027 2306 3039
rect 2194 3007 2206 3019
rect 2234 3007 2246 3019
rect 2353 2987 2365 2999
rect 2454 3041 2466 3053
rect 2394 2987 2406 2999
rect 2374 2967 2386 2979
rect 2494 3041 2506 3053
rect 2474 3027 2486 3039
rect 2553 2987 2565 2999
rect 2674 3041 2686 3053
rect 2594 2987 2606 2999
rect 2635 2987 2647 2999
rect 2574 2967 2586 2979
rect 2794 3021 2806 3033
rect 2694 3007 2706 3019
rect 2734 3007 2746 3019
rect 2774 3007 2786 3019
rect 2834 3021 2846 3033
rect 2874 3021 2886 3033
rect 2914 3021 2926 3033
rect 2975 3041 2987 3053
rect 3013 3041 3025 3053
rect 2955 3007 2967 3019
rect 3074 3021 3086 3033
rect 3034 3007 3046 3019
rect 3114 3021 3126 3033
rect 3174 3041 3186 3053
rect 3154 3007 3166 3019
rect 3254 3041 3266 3053
rect 3213 2987 3225 2999
rect 3355 3058 3367 3070
rect 3445 3058 3457 3070
rect 3354 3021 3366 3033
rect 3314 3007 3326 3019
rect 3525 3058 3537 3070
rect 3574 3021 3586 3033
rect 3474 3007 3486 3019
rect 3554 3007 3566 3019
rect 3445 2990 3457 3002
rect 3525 2990 3537 3002
rect 3614 3021 3626 3033
rect 3674 3041 3686 3053
rect 3654 3007 3666 3019
rect 3785 3058 3797 3070
rect 3854 3041 3866 3053
rect 3814 3007 3826 3019
rect 3834 3007 3846 3019
rect 3713 2987 3725 2999
rect 3785 2990 3797 3002
rect 3893 2987 3905 2999
rect 3934 2987 3946 2999
rect 4063 3058 4075 3070
rect 4034 3007 4046 3019
rect 3975 2987 3987 2999
rect 3954 2967 3966 2979
rect 4154 3041 4166 3053
rect 4063 2990 4075 3002
rect 4194 3041 4206 3053
rect 4174 3027 4186 3039
rect 4214 2987 4226 2999
rect 4354 3041 4366 3053
rect 4255 2987 4267 2999
rect 4234 2967 4246 2979
rect 4394 3041 4406 3053
rect 4374 3027 4386 3039
rect 4453 2987 4465 2999
rect 4554 3027 4566 3039
rect 4494 2987 4506 2999
rect 4474 2967 4486 2979
rect 4634 3041 4646 3053
rect 4595 2987 4607 2999
rect 4694 3041 4706 3053
rect 4654 3007 4666 3019
rect 4674 3007 4686 3019
rect 4733 2987 4745 2999
rect 101 2818 113 2830
rect 83 2784 95 2796
rect 34 2741 46 2753
rect 54 2742 66 2754
rect 74 2728 86 2740
rect 135 2818 147 2830
rect 115 2798 127 2810
rect 77 2696 89 2708
rect 99 2696 111 2708
rect 163 2804 175 2816
rect 187 2804 199 2816
rect 147 2700 159 2712
rect 215 2772 227 2784
rect 201 2733 213 2745
rect 274 2761 286 2773
rect 353 2761 365 2773
rect 295 2727 307 2739
rect 333 2727 345 2739
rect 374 2747 386 2759
rect 475 2781 487 2793
rect 414 2747 426 2759
rect 585 2778 597 2790
rect 534 2761 546 2773
rect 614 2761 626 2773
rect 514 2727 526 2739
rect 585 2710 597 2722
rect 634 2747 646 2759
rect 735 2781 747 2793
rect 674 2747 686 2759
rect 794 2761 806 2773
rect 834 2761 846 2773
rect 874 2761 886 2773
rect 774 2727 786 2739
rect 914 2747 926 2759
rect 954 2747 966 2759
rect 974 2741 986 2753
rect 1054 2747 1066 2759
rect 1114 2761 1126 2773
rect 1225 2778 1237 2790
rect 1154 2761 1166 2773
rect 1254 2761 1266 2773
rect 1094 2747 1106 2759
rect 1225 2710 1237 2722
rect 1361 2818 1373 2830
rect 1343 2784 1355 2796
rect 1294 2741 1306 2753
rect 1314 2742 1326 2754
rect 1334 2728 1346 2740
rect 1395 2818 1407 2830
rect 1375 2798 1387 2810
rect 1337 2696 1349 2708
rect 1359 2696 1371 2708
rect 1423 2804 1435 2816
rect 1447 2804 1459 2816
rect 1407 2700 1419 2712
rect 1475 2772 1487 2784
rect 1461 2733 1473 2745
rect 1514 2747 1526 2759
rect 1615 2781 1627 2793
rect 1554 2747 1566 2759
rect 1715 2781 1727 2793
rect 1674 2761 1686 2773
rect 1654 2727 1666 2739
rect 1774 2761 1786 2773
rect 1814 2761 1826 2773
rect 1854 2761 1866 2773
rect 1754 2727 1766 2739
rect 2005 2778 2017 2790
rect 1934 2741 1946 2753
rect 1914 2727 1926 2739
rect 2114 2801 2126 2813
rect 2093 2781 2105 2793
rect 2034 2761 2046 2773
rect 1954 2727 1966 2739
rect 2005 2710 2017 2722
rect 2134 2781 2146 2793
rect 2183 2778 2195 2790
rect 2154 2761 2166 2773
rect 2321 2818 2333 2830
rect 2303 2784 2315 2796
rect 2254 2741 2266 2753
rect 2274 2742 2286 2754
rect 2183 2710 2195 2722
rect 2294 2728 2306 2740
rect 2355 2818 2367 2830
rect 2335 2798 2347 2810
rect 2297 2696 2309 2708
rect 2319 2696 2331 2708
rect 2383 2804 2395 2816
rect 2407 2804 2419 2816
rect 2367 2700 2379 2712
rect 2435 2772 2447 2784
rect 2495 2781 2507 2793
rect 2421 2733 2433 2745
rect 2595 2781 2607 2793
rect 2554 2761 2566 2773
rect 2534 2727 2546 2739
rect 2654 2761 2666 2773
rect 2674 2761 2686 2773
rect 2634 2727 2646 2739
rect 2733 2781 2745 2793
rect 2694 2727 2706 2739
rect 2774 2747 2786 2759
rect 2814 2747 2826 2759
rect 2854 2747 2866 2759
rect 2934 2761 2946 2773
rect 2894 2747 2906 2759
rect 2993 2781 3005 2793
rect 2954 2727 2966 2739
rect 3034 2761 3046 2773
rect 3093 2781 3105 2793
rect 3054 2727 3066 2739
rect 3134 2747 3146 2759
rect 3235 2781 3247 2793
rect 3174 2747 3186 2759
rect 3294 2761 3306 2773
rect 3274 2727 3286 2739
rect 3334 2747 3346 2759
rect 3414 2801 3426 2813
rect 3394 2781 3406 2793
rect 3374 2747 3386 2759
rect 3435 2781 3447 2793
rect 3515 2781 3527 2793
rect 3574 2761 3586 2773
rect 3594 2761 3606 2773
rect 3554 2727 3566 2739
rect 3653 2781 3665 2793
rect 3614 2727 3626 2739
rect 3714 2747 3726 2759
rect 3795 2781 3807 2793
rect 3754 2747 3766 2759
rect 3894 2801 3906 2813
rect 3874 2781 3886 2793
rect 3854 2761 3866 2773
rect 3834 2727 3846 2739
rect 3915 2781 3927 2793
rect 4054 2761 4066 2773
rect 3974 2741 3986 2753
rect 4174 2801 4186 2813
rect 4154 2781 4166 2793
rect 4133 2761 4145 2773
rect 4075 2727 4087 2739
rect 4113 2727 4125 2739
rect 4195 2781 4207 2793
rect 4254 2761 4266 2773
rect 4313 2781 4325 2793
rect 4274 2727 4286 2739
rect 4354 2761 4366 2773
rect 4394 2747 4406 2759
rect 4455 2761 4467 2773
rect 4395 2710 4407 2722
rect 4534 2761 4546 2773
rect 4475 2727 4487 2739
rect 4513 2727 4525 2739
rect 4574 2741 4586 2753
rect 4654 2741 4666 2753
rect 4634 2727 4646 2739
rect 4674 2727 4686 2739
rect 34 2547 46 2559
rect 77 2592 89 2604
rect 99 2592 111 2604
rect 74 2560 86 2572
rect 54 2546 66 2558
rect 83 2504 95 2516
rect 115 2490 127 2502
rect 101 2470 113 2482
rect 147 2588 159 2600
rect 201 2555 213 2567
rect 215 2516 227 2528
rect 314 2561 326 2573
rect 275 2507 287 2519
rect 163 2484 175 2496
rect 135 2470 147 2482
rect 187 2484 199 2496
rect 383 2578 395 2590
rect 434 2541 446 2553
rect 334 2527 346 2539
rect 354 2527 366 2539
rect 383 2510 395 2522
rect 474 2541 486 2553
rect 574 2561 586 2573
rect 535 2507 547 2519
rect 643 2578 655 2590
rect 594 2527 606 2539
rect 614 2527 626 2539
rect 643 2510 655 2522
rect 754 2561 766 2573
rect 715 2507 727 2519
rect 894 2547 906 2559
rect 937 2592 949 2604
rect 959 2592 971 2604
rect 934 2560 946 2572
rect 774 2527 786 2539
rect 794 2527 806 2539
rect 834 2527 846 2539
rect 914 2546 926 2558
rect 943 2504 955 2516
rect 975 2490 987 2502
rect 961 2470 973 2482
rect 1007 2588 1019 2600
rect 1061 2555 1073 2567
rect 1114 2547 1126 2559
rect 1075 2516 1087 2528
rect 1023 2484 1035 2496
rect 995 2470 1007 2482
rect 1047 2484 1059 2496
rect 1194 2561 1206 2573
rect 1174 2527 1186 2539
rect 1274 2547 1286 2559
rect 1233 2507 1245 2519
rect 1334 2541 1346 2553
rect 1374 2541 1386 2553
rect 1447 2555 1459 2567
rect 1433 2516 1445 2528
rect 1501 2588 1513 2600
rect 1461 2484 1473 2496
rect 1485 2484 1497 2496
rect 1549 2592 1561 2604
rect 1571 2592 1583 2604
rect 1533 2490 1545 2502
rect 1513 2470 1525 2482
rect 1574 2560 1586 2572
rect 1594 2546 1606 2558
rect 1614 2547 1626 2559
rect 1565 2504 1577 2516
rect 1547 2470 1559 2482
rect 1674 2561 1686 2573
rect 1654 2527 1666 2539
rect 1787 2555 1799 2567
rect 1713 2507 1725 2519
rect 1773 2516 1785 2528
rect 1841 2588 1853 2600
rect 1801 2484 1813 2496
rect 1825 2484 1837 2496
rect 1889 2592 1901 2604
rect 1911 2592 1923 2604
rect 1873 2490 1885 2502
rect 1853 2470 1865 2482
rect 1914 2560 1926 2572
rect 2014 2561 2026 2573
rect 2050 2564 2062 2576
rect 2090 2564 2102 2576
rect 2130 2564 2142 2576
rect 1934 2546 1946 2558
rect 1954 2547 1966 2559
rect 1905 2504 1917 2516
rect 1887 2470 1899 2482
rect 2214 2547 2226 2559
rect 2257 2592 2269 2604
rect 2279 2592 2291 2604
rect 2254 2560 2266 2572
rect 2234 2546 2246 2558
rect 2263 2504 2275 2516
rect 2295 2490 2307 2502
rect 2281 2470 2293 2482
rect 2327 2588 2339 2600
rect 2381 2555 2393 2567
rect 2454 2541 2466 2553
rect 2395 2516 2407 2528
rect 2343 2484 2355 2496
rect 2315 2470 2327 2482
rect 2367 2484 2379 2496
rect 2494 2541 2506 2553
rect 2514 2547 2526 2559
rect 2634 2561 2646 2573
rect 2595 2507 2607 2519
rect 2674 2547 2686 2559
rect 2654 2527 2666 2539
rect 2754 2541 2766 2553
rect 2794 2541 2806 2553
rect 2874 2561 2886 2573
rect 2835 2507 2847 2519
rect 2955 2578 2967 2590
rect 2954 2541 2966 2553
rect 2894 2527 2906 2539
rect 2914 2527 2926 2539
rect 3034 2561 3046 2573
rect 3014 2527 3026 2539
rect 3134 2541 3146 2553
rect 3073 2507 3085 2519
rect 3174 2541 3186 2553
rect 3235 2578 3247 2590
rect 3234 2541 3246 2553
rect 3194 2527 3206 2539
rect 3333 2507 3345 2519
rect 3394 2547 3406 2559
rect 3374 2507 3386 2519
rect 3354 2487 3366 2499
rect 3454 2541 3466 2553
rect 3494 2541 3506 2553
rect 3575 2578 3587 2590
rect 3574 2541 3586 2553
rect 3534 2527 3546 2539
rect 3663 2578 3675 2590
rect 3714 2547 3726 2559
rect 3634 2527 3646 2539
rect 3663 2510 3675 2522
rect 3813 2578 3825 2590
rect 3814 2541 3826 2553
rect 3915 2561 3927 2573
rect 3953 2561 3965 2573
rect 3854 2527 3866 2539
rect 3894 2527 3906 2539
rect 4014 2541 4026 2553
rect 3973 2527 3985 2539
rect 4054 2541 4066 2553
rect 4094 2541 4106 2553
rect 4134 2541 4146 2553
rect 4174 2561 4186 2573
rect 4154 2527 4166 2539
rect 4254 2541 4266 2553
rect 4213 2507 4225 2519
rect 4294 2541 4306 2553
rect 4373 2507 4385 2519
rect 4414 2507 4426 2519
rect 4473 2507 4485 2519
rect 4394 2487 4406 2499
rect 4534 2561 4546 2573
rect 4574 2561 4586 2573
rect 4554 2547 4566 2559
rect 4514 2507 4526 2519
rect 4494 2487 4506 2499
rect 4673 2507 4685 2519
rect 4714 2507 4726 2519
rect 4694 2487 4706 2499
rect 101 2338 113 2350
rect 83 2304 95 2316
rect 34 2261 46 2273
rect 54 2262 66 2274
rect 74 2248 86 2260
rect 135 2338 147 2350
rect 115 2318 127 2330
rect 77 2216 89 2228
rect 99 2216 111 2228
rect 163 2324 175 2336
rect 187 2324 199 2336
rect 147 2220 159 2232
rect 215 2292 227 2304
rect 201 2253 213 2265
rect 254 2281 266 2293
rect 313 2301 325 2313
rect 274 2247 286 2259
rect 355 2281 367 2293
rect 503 2298 515 2310
rect 434 2281 446 2293
rect 474 2281 486 2293
rect 375 2247 387 2259
rect 413 2247 425 2259
rect 554 2267 566 2279
rect 594 2267 606 2279
rect 694 2281 706 2293
rect 734 2281 746 2293
rect 503 2230 515 2242
rect 674 2261 686 2273
rect 834 2261 846 2273
rect 814 2247 826 2259
rect 874 2281 886 2293
rect 914 2281 926 2293
rect 954 2281 966 2293
rect 994 2281 1006 2293
rect 854 2247 866 2259
rect 1141 2324 1153 2336
rect 1193 2338 1205 2350
rect 1165 2324 1177 2336
rect 1034 2261 1046 2273
rect 1113 2292 1125 2304
rect 1127 2253 1139 2265
rect 1181 2220 1193 2232
rect 1227 2338 1239 2350
rect 1213 2318 1225 2330
rect 1245 2304 1257 2316
rect 1274 2262 1286 2274
rect 1334 2281 1346 2293
rect 1254 2248 1266 2260
rect 1229 2216 1241 2228
rect 1251 2216 1263 2228
rect 1294 2261 1306 2273
rect 1481 2324 1493 2336
rect 1533 2338 1545 2350
rect 1505 2324 1517 2336
rect 1393 2301 1405 2313
rect 1354 2247 1366 2259
rect 1453 2292 1465 2304
rect 1467 2253 1479 2265
rect 1521 2220 1533 2232
rect 1567 2338 1579 2350
rect 1553 2318 1565 2330
rect 1585 2304 1597 2316
rect 1614 2262 1626 2274
rect 1694 2281 1706 2293
rect 1734 2281 1746 2293
rect 1594 2248 1606 2260
rect 1569 2216 1581 2228
rect 1591 2216 1603 2228
rect 1634 2261 1646 2273
rect 1814 2261 1826 2273
rect 1794 2247 1806 2259
rect 1934 2281 1946 2293
rect 1974 2281 1986 2293
rect 1834 2247 1846 2259
rect 1854 2247 1866 2259
rect 2014 2247 2026 2259
rect 2194 2281 2206 2293
rect 2050 2244 2062 2256
rect 2090 2244 2102 2256
rect 2130 2244 2142 2256
rect 2253 2301 2265 2313
rect 2214 2247 2226 2259
rect 2381 2338 2393 2350
rect 2363 2304 2375 2316
rect 2314 2261 2326 2273
rect 2334 2262 2346 2274
rect 2354 2248 2366 2260
rect 2415 2338 2427 2350
rect 2395 2318 2407 2330
rect 2357 2216 2369 2228
rect 2379 2216 2391 2228
rect 2443 2324 2455 2336
rect 2467 2324 2479 2336
rect 2427 2220 2439 2232
rect 2495 2292 2507 2304
rect 2481 2253 2493 2265
rect 2554 2267 2566 2279
rect 2594 2267 2606 2279
rect 2614 2267 2626 2279
rect 2654 2267 2666 2279
rect 2694 2267 2706 2279
rect 2795 2301 2807 2313
rect 2734 2267 2746 2279
rect 2895 2301 2907 2313
rect 2854 2281 2866 2293
rect 2834 2247 2846 2259
rect 2954 2281 2966 2293
rect 2934 2247 2946 2259
rect 3061 2338 3073 2350
rect 3043 2304 3055 2316
rect 2994 2261 3006 2273
rect 3014 2262 3026 2274
rect 3034 2248 3046 2260
rect 3095 2338 3107 2350
rect 3075 2318 3087 2330
rect 3037 2216 3049 2228
rect 3059 2216 3071 2228
rect 3123 2324 3135 2336
rect 3147 2324 3159 2336
rect 3107 2220 3119 2232
rect 3175 2292 3187 2304
rect 3161 2253 3173 2265
rect 3214 2281 3226 2293
rect 3273 2301 3285 2313
rect 3234 2247 3246 2259
rect 3314 2267 3326 2279
rect 3354 2267 3366 2279
rect 3394 2267 3406 2279
rect 3434 2267 3446 2279
rect 3494 2267 3506 2279
rect 3534 2267 3546 2279
rect 3734 2281 3746 2293
rect 3714 2261 3726 2273
rect 3594 2247 3606 2259
rect 3654 2247 3666 2259
rect 3793 2301 3805 2313
rect 3754 2247 3766 2259
rect 3865 2298 3877 2310
rect 3894 2281 3906 2293
rect 3865 2230 3877 2242
rect 3974 2281 3986 2293
rect 3914 2247 3926 2259
rect 4014 2267 4026 2279
rect 4095 2301 4107 2313
rect 4015 2230 4027 2242
rect 4234 2321 4246 2333
rect 4213 2301 4225 2313
rect 4154 2281 4166 2293
rect 4134 2247 4146 2259
rect 4254 2301 4266 2313
rect 4294 2261 4306 2273
rect 4274 2247 4286 2259
rect 4395 2301 4407 2313
rect 4314 2247 4326 2259
rect 4454 2281 4466 2293
rect 4474 2281 4486 2293
rect 4434 2247 4446 2259
rect 4533 2301 4545 2313
rect 4595 2301 4607 2313
rect 4494 2247 4506 2259
rect 4654 2281 4666 2293
rect 4634 2247 4646 2259
rect 4694 2261 4706 2273
rect 4674 2247 4686 2259
rect 4714 2247 4726 2259
rect 34 2081 46 2093
rect 70 2084 82 2096
rect 110 2084 122 2096
rect 150 2084 162 2096
rect 234 2061 246 2073
rect 274 2061 286 2073
rect 354 2081 366 2093
rect 315 2027 327 2039
rect 415 2081 427 2093
rect 453 2081 465 2093
rect 374 2047 386 2059
rect 395 2047 407 2059
rect 534 2067 546 2079
rect 577 2112 589 2124
rect 599 2112 611 2124
rect 574 2080 586 2092
rect 474 2047 486 2059
rect 554 2066 566 2078
rect 583 2024 595 2036
rect 615 2010 627 2022
rect 601 1990 613 2002
rect 647 2108 659 2120
rect 701 2075 713 2087
rect 875 2096 887 2108
rect 774 2061 786 2073
rect 715 2036 727 2048
rect 663 2004 675 2016
rect 635 1990 647 2002
rect 687 2004 699 2016
rect 814 2061 826 2073
rect 914 2067 926 2079
rect 894 2047 906 2059
rect 875 2029 887 2041
rect 934 2061 946 2073
rect 974 2061 986 2073
rect 1114 2081 1126 2093
rect 1014 2047 1026 2059
rect 1054 2047 1066 2059
rect 1094 2047 1106 2059
rect 1194 2061 1206 2073
rect 1153 2027 1165 2039
rect 1234 2061 1246 2073
rect 1274 2047 1286 2059
rect 1314 2047 1326 2059
rect 1387 2075 1399 2087
rect 1373 2036 1385 2048
rect 1441 2108 1453 2120
rect 1401 2004 1413 2016
rect 1425 2004 1437 2016
rect 1489 2112 1501 2124
rect 1511 2112 1523 2124
rect 1473 2010 1485 2022
rect 1453 1990 1465 2002
rect 1514 2080 1526 2092
rect 1634 2081 1646 2093
rect 1534 2066 1546 2078
rect 1554 2067 1566 2079
rect 1505 2024 1517 2036
rect 1487 1990 1499 2002
rect 1725 2098 1737 2110
rect 1674 2081 1686 2093
rect 1654 2067 1666 2079
rect 1754 2047 1766 2059
rect 1807 2075 1819 2087
rect 1725 2030 1737 2042
rect 1793 2036 1805 2048
rect 1861 2108 1873 2120
rect 1821 2004 1833 2016
rect 1845 2004 1857 2016
rect 1909 2112 1921 2124
rect 1931 2112 1943 2124
rect 1893 2010 1905 2022
rect 1873 1990 1885 2002
rect 1934 2080 1946 2092
rect 1954 2066 1966 2078
rect 1974 2067 1986 2079
rect 2054 2067 2066 2079
rect 1925 2024 1937 2036
rect 1907 1990 1919 2002
rect 2094 2061 2106 2073
rect 2134 2061 2146 2073
rect 2183 2098 2195 2110
rect 2234 2061 2246 2073
rect 2154 2047 2166 2059
rect 2183 2030 2195 2042
rect 2274 2061 2286 2073
rect 2374 2081 2386 2093
rect 2335 2027 2347 2039
rect 2434 2061 2446 2073
rect 2394 2047 2406 2059
rect 2474 2061 2486 2073
rect 2514 2061 2526 2073
rect 2554 2061 2566 2073
rect 2634 2081 2646 2093
rect 2595 2027 2607 2039
rect 2654 2047 2666 2059
rect 2734 2081 2746 2093
rect 2695 2027 2707 2039
rect 2794 2067 2806 2079
rect 2837 2112 2849 2124
rect 2859 2112 2871 2124
rect 2834 2080 2846 2092
rect 2754 2047 2766 2059
rect 2814 2066 2826 2078
rect 2843 2024 2855 2036
rect 2875 2010 2887 2022
rect 2861 1990 2873 2002
rect 2907 2108 2919 2120
rect 2961 2075 2973 2087
rect 3055 2098 3067 2110
rect 3054 2061 3066 2073
rect 2975 2036 2987 2048
rect 3014 2047 3026 2059
rect 2923 2004 2935 2016
rect 2895 1990 2907 2002
rect 2947 2004 2959 2016
rect 3174 2081 3186 2093
rect 3135 2027 3147 2039
rect 3194 2047 3206 2059
rect 3274 2081 3286 2093
rect 3235 2027 3247 2039
rect 3314 2061 3326 2073
rect 3294 2047 3306 2059
rect 3354 2061 3366 2073
rect 3454 2081 3466 2093
rect 3415 2027 3427 2039
rect 3474 2047 3486 2059
rect 3494 2027 3506 2039
rect 3594 2067 3606 2079
rect 3535 2027 3547 2039
rect 3514 2007 3526 2019
rect 3654 2027 3666 2039
rect 3754 2061 3766 2073
rect 3695 2027 3707 2039
rect 3674 2007 3686 2019
rect 3794 2061 3806 2073
rect 3863 2098 3875 2110
rect 3934 2081 3946 2093
rect 3834 2047 3846 2059
rect 3914 2047 3926 2059
rect 3863 2030 3875 2042
rect 4034 2061 4046 2073
rect 3973 2027 3985 2039
rect 4074 2061 4086 2073
rect 4114 2061 4126 2073
rect 4154 2061 4166 2073
rect 4194 2061 4206 2073
rect 4234 2061 4246 2073
rect 4295 2098 4307 2110
rect 4294 2061 4306 2073
rect 4254 2047 4266 2059
rect 4354 2081 4366 2093
rect 4394 2081 4406 2093
rect 4374 2067 4386 2079
rect 4494 2081 4506 2093
rect 4534 2081 4546 2093
rect 4514 2067 4526 2079
rect 4554 2027 4566 2039
rect 4595 2027 4607 2039
rect 4654 2027 4666 2039
rect 4574 2007 4586 2019
rect 4695 2027 4707 2039
rect 4674 2007 4686 2019
rect 101 1858 113 1870
rect 83 1824 95 1836
rect 34 1781 46 1793
rect 54 1782 66 1794
rect 74 1768 86 1780
rect 135 1858 147 1870
rect 115 1838 127 1850
rect 77 1736 89 1748
rect 99 1736 111 1748
rect 163 1844 175 1856
rect 187 1844 199 1856
rect 147 1740 159 1752
rect 215 1812 227 1824
rect 201 1773 213 1785
rect 254 1801 266 1813
rect 313 1821 325 1833
rect 375 1821 387 1833
rect 274 1767 286 1779
rect 475 1821 487 1833
rect 434 1801 446 1813
rect 414 1767 426 1779
rect 575 1821 587 1833
rect 534 1801 546 1813
rect 514 1767 526 1779
rect 634 1801 646 1813
rect 614 1767 626 1779
rect 794 1801 806 1813
rect 874 1841 886 1853
rect 854 1821 866 1833
rect 834 1801 846 1813
rect 654 1781 666 1793
rect 714 1781 726 1793
rect 895 1821 907 1833
rect 1041 1858 1053 1870
rect 1023 1824 1035 1836
rect 974 1781 986 1793
rect 994 1782 1006 1794
rect 1014 1768 1026 1780
rect 1075 1858 1087 1870
rect 1055 1838 1067 1850
rect 1017 1736 1029 1748
rect 1039 1736 1051 1748
rect 1103 1844 1115 1856
rect 1127 1844 1139 1856
rect 1087 1740 1099 1752
rect 1155 1812 1167 1824
rect 1141 1773 1153 1785
rect 1194 1787 1206 1799
rect 1295 1821 1307 1833
rect 1234 1787 1246 1799
rect 1354 1801 1366 1813
rect 1334 1767 1346 1779
rect 1661 1858 1673 1870
rect 1643 1824 1655 1836
rect 1594 1781 1606 1793
rect 1614 1782 1626 1794
rect 1418 1764 1430 1776
rect 1458 1764 1470 1776
rect 1498 1764 1510 1776
rect 1534 1767 1546 1779
rect 1634 1768 1646 1780
rect 1695 1858 1707 1870
rect 1675 1838 1687 1850
rect 1637 1736 1649 1748
rect 1659 1736 1671 1748
rect 1723 1844 1735 1856
rect 1747 1844 1759 1856
rect 1707 1740 1719 1752
rect 2321 1844 2333 1856
rect 2373 1858 2385 1870
rect 2345 1844 2357 1856
rect 1775 1812 1787 1824
rect 1761 1773 1773 1785
rect 1874 1781 1886 1793
rect 1854 1767 1866 1779
rect 1914 1801 1926 1813
rect 1954 1801 1966 1813
rect 1894 1767 1906 1779
rect 2054 1781 2066 1793
rect 2034 1767 2046 1779
rect 2114 1801 2126 1813
rect 2154 1801 2166 1813
rect 2074 1767 2086 1779
rect 2194 1781 2206 1793
rect 2174 1767 2186 1779
rect 2214 1767 2226 1779
rect 2293 1812 2305 1824
rect 2307 1773 2319 1785
rect 2361 1740 2373 1752
rect 2407 1858 2419 1870
rect 2393 1838 2405 1850
rect 2425 1824 2437 1836
rect 2454 1782 2466 1794
rect 2601 1858 2613 1870
rect 2583 1824 2595 1836
rect 2434 1768 2446 1780
rect 2409 1736 2421 1748
rect 2431 1736 2443 1748
rect 2474 1781 2486 1793
rect 2534 1781 2546 1793
rect 2554 1782 2566 1794
rect 2574 1768 2586 1780
rect 2635 1858 2647 1870
rect 2615 1838 2627 1850
rect 2577 1736 2589 1748
rect 2599 1736 2611 1748
rect 2663 1844 2675 1856
rect 2687 1844 2699 1856
rect 2647 1740 2659 1752
rect 2715 1812 2727 1824
rect 2701 1773 2713 1785
rect 2841 1858 2853 1870
rect 2823 1824 2835 1836
rect 2774 1781 2786 1793
rect 2794 1782 2806 1794
rect 2814 1768 2826 1780
rect 2875 1858 2887 1870
rect 2855 1838 2867 1850
rect 2817 1736 2829 1748
rect 2839 1736 2851 1748
rect 2903 1844 2915 1856
rect 2927 1844 2939 1856
rect 2887 1740 2899 1752
rect 2955 1812 2967 1824
rect 2941 1773 2953 1785
rect 3074 1787 3086 1799
rect 3034 1767 3046 1779
rect 3114 1787 3126 1799
rect 3214 1781 3226 1793
rect 3174 1767 3186 1779
rect 3194 1767 3206 1779
rect 3294 1801 3306 1813
rect 3334 1801 3346 1813
rect 3234 1767 3246 1779
rect 3454 1801 3466 1813
rect 3414 1787 3426 1799
rect 3413 1750 3425 1762
rect 3554 1801 3566 1813
rect 3474 1767 3486 1779
rect 3633 1801 3645 1813
rect 3575 1767 3587 1779
rect 3613 1767 3625 1779
rect 3734 1801 3746 1813
rect 3823 1818 3835 1830
rect 3774 1801 3786 1813
rect 3794 1801 3806 1813
rect 3874 1801 3886 1813
rect 3694 1767 3706 1779
rect 3823 1750 3835 1762
rect 3914 1787 3926 1799
rect 3994 1801 4006 1813
rect 3915 1750 3927 1762
rect 4073 1801 4085 1813
rect 4095 1801 4107 1813
rect 4015 1767 4027 1779
rect 4053 1767 4065 1779
rect 4174 1801 4186 1813
rect 4115 1767 4127 1779
rect 4153 1767 4165 1779
rect 4214 1787 4226 1799
rect 4294 1801 4306 1813
rect 4254 1787 4266 1799
rect 4334 1787 4346 1799
rect 4395 1801 4407 1813
rect 4335 1750 4347 1762
rect 4474 1801 4486 1813
rect 4415 1767 4427 1779
rect 4453 1767 4465 1779
rect 4574 1801 4586 1813
rect 4554 1781 4566 1793
rect 4633 1821 4645 1833
rect 4594 1767 4606 1779
rect 4674 1781 4686 1793
rect 34 1601 46 1613
rect 70 1604 82 1616
rect 110 1604 122 1616
rect 150 1604 162 1616
rect 325 1618 337 1630
rect 394 1587 406 1599
rect 437 1632 449 1644
rect 459 1632 471 1644
rect 434 1600 446 1612
rect 234 1567 246 1579
rect 274 1567 286 1579
rect 354 1567 366 1579
rect 325 1550 337 1562
rect 414 1586 426 1598
rect 443 1544 455 1556
rect 475 1530 487 1542
rect 461 1510 473 1522
rect 507 1628 519 1640
rect 561 1595 573 1607
rect 634 1587 646 1599
rect 677 1632 689 1644
rect 699 1632 711 1644
rect 674 1600 686 1612
rect 575 1556 587 1568
rect 654 1586 666 1598
rect 523 1524 535 1536
rect 495 1510 507 1522
rect 547 1524 559 1536
rect 683 1544 695 1556
rect 715 1530 727 1542
rect 701 1510 713 1522
rect 747 1628 759 1640
rect 801 1595 813 1607
rect 815 1556 827 1568
rect 887 1595 899 1607
rect 873 1556 885 1568
rect 763 1524 775 1536
rect 735 1510 747 1522
rect 787 1524 799 1536
rect 941 1628 953 1640
rect 901 1524 913 1536
rect 925 1524 937 1536
rect 989 1632 1001 1644
rect 1011 1632 1023 1644
rect 973 1530 985 1542
rect 953 1510 965 1522
rect 1014 1600 1026 1612
rect 1034 1586 1046 1598
rect 1054 1587 1066 1599
rect 1005 1544 1017 1556
rect 987 1510 999 1522
rect 1114 1581 1126 1593
rect 1154 1581 1166 1593
rect 1234 1601 1246 1613
rect 1195 1547 1207 1559
rect 1254 1567 1266 1579
rect 1307 1595 1319 1607
rect 1293 1556 1305 1568
rect 1361 1628 1373 1640
rect 1321 1524 1333 1536
rect 1345 1524 1357 1536
rect 1409 1632 1421 1644
rect 1431 1632 1443 1644
rect 1393 1530 1405 1542
rect 1373 1510 1385 1522
rect 1434 1600 1446 1612
rect 1454 1586 1466 1598
rect 1474 1587 1486 1599
rect 1534 1587 1546 1599
rect 1577 1632 1589 1644
rect 1599 1632 1611 1644
rect 1574 1600 1586 1612
rect 1425 1544 1437 1556
rect 1407 1510 1419 1522
rect 1554 1586 1566 1598
rect 1583 1544 1595 1556
rect 1615 1530 1627 1542
rect 1601 1510 1613 1522
rect 1647 1628 1659 1640
rect 1701 1595 1713 1607
rect 1715 1556 1727 1568
rect 1794 1601 1806 1613
rect 1834 1601 1846 1613
rect 1814 1587 1826 1599
rect 1954 1587 1966 1599
rect 1997 1632 2009 1644
rect 2019 1632 2031 1644
rect 1994 1600 2006 1612
rect 1854 1567 1866 1579
rect 1894 1567 1906 1579
rect 1974 1586 1986 1598
rect 1663 1524 1675 1536
rect 1635 1510 1647 1522
rect 1687 1524 1699 1536
rect 2003 1544 2015 1556
rect 2035 1530 2047 1542
rect 2021 1510 2033 1522
rect 2067 1628 2079 1640
rect 2121 1595 2133 1607
rect 2274 1581 2286 1593
rect 2135 1556 2147 1568
rect 2194 1567 2206 1579
rect 2234 1567 2246 1579
rect 2083 1524 2095 1536
rect 2055 1510 2067 1522
rect 2107 1524 2119 1536
rect 2314 1581 2326 1593
rect 2354 1601 2366 1613
rect 2334 1567 2346 1579
rect 2467 1595 2479 1607
rect 2393 1547 2405 1559
rect 2453 1556 2465 1568
rect 2521 1628 2533 1640
rect 2481 1524 2493 1536
rect 2505 1524 2517 1536
rect 2569 1632 2581 1644
rect 2591 1632 2603 1644
rect 2553 1530 2565 1542
rect 2533 1510 2545 1522
rect 2594 1600 2606 1612
rect 2614 1586 2626 1598
rect 2634 1587 2646 1599
rect 2694 1587 2706 1599
rect 2737 1632 2749 1644
rect 2759 1632 2771 1644
rect 2734 1600 2746 1612
rect 2585 1544 2597 1556
rect 2567 1510 2579 1522
rect 2714 1586 2726 1598
rect 2743 1544 2755 1556
rect 2775 1530 2787 1542
rect 2761 1510 2773 1522
rect 2807 1628 2819 1640
rect 2861 1595 2873 1607
rect 2914 1601 2926 1613
rect 2875 1556 2887 1568
rect 2974 1581 2986 1593
rect 2823 1524 2835 1536
rect 2795 1510 2807 1522
rect 2847 1524 2859 1536
rect 3014 1581 3026 1593
rect 3074 1581 3086 1593
rect 3114 1581 3126 1593
rect 3154 1601 3166 1613
rect 3134 1567 3146 1579
rect 3234 1581 3246 1593
rect 3193 1547 3205 1559
rect 3274 1581 3286 1593
rect 3334 1581 3346 1593
rect 3374 1581 3386 1593
rect 3454 1601 3466 1613
rect 3415 1547 3427 1559
rect 3474 1567 3486 1579
rect 3494 1547 3506 1559
rect 3638 1601 3650 1613
rect 3674 1601 3686 1613
rect 3615 1567 3627 1579
rect 3535 1547 3547 1559
rect 3514 1527 3526 1539
rect 3714 1587 3726 1599
rect 3694 1567 3706 1579
rect 3774 1547 3786 1559
rect 3874 1601 3886 1613
rect 3914 1601 3926 1613
rect 3894 1587 3906 1599
rect 3815 1547 3827 1559
rect 3794 1527 3806 1539
rect 3994 1601 4006 1613
rect 3974 1567 3986 1579
rect 4094 1581 4106 1593
rect 4033 1547 4045 1559
rect 4154 1601 4166 1613
rect 4134 1581 4146 1593
rect 4194 1601 4206 1613
rect 4174 1587 4186 1599
rect 4274 1601 4286 1613
rect 4254 1567 4266 1579
rect 4354 1587 4366 1599
rect 4313 1547 4325 1559
rect 4494 1581 4506 1593
rect 4414 1567 4426 1579
rect 4454 1567 4466 1579
rect 4534 1581 4546 1593
rect 4574 1581 4586 1593
rect 4614 1581 4626 1593
rect 4654 1581 4666 1593
rect 4694 1581 4706 1593
rect 61 1364 73 1376
rect 113 1378 125 1390
rect 85 1364 97 1376
rect 33 1332 45 1344
rect 47 1293 59 1305
rect 101 1260 113 1272
rect 147 1378 159 1390
rect 133 1358 145 1370
rect 165 1344 177 1356
rect 194 1302 206 1314
rect 341 1378 353 1390
rect 323 1344 335 1356
rect 174 1288 186 1300
rect 149 1256 161 1268
rect 171 1256 183 1268
rect 214 1301 226 1313
rect 274 1301 286 1313
rect 294 1302 306 1314
rect 314 1288 326 1300
rect 375 1378 387 1390
rect 355 1358 367 1370
rect 317 1256 329 1268
rect 339 1256 351 1268
rect 403 1364 415 1376
rect 427 1364 439 1376
rect 387 1260 399 1272
rect 455 1332 467 1344
rect 441 1293 453 1305
rect 494 1307 506 1319
rect 595 1341 607 1353
rect 534 1307 546 1319
rect 695 1341 707 1353
rect 654 1321 666 1333
rect 634 1287 646 1299
rect 805 1338 817 1350
rect 754 1321 766 1333
rect 834 1321 846 1333
rect 734 1287 746 1299
rect 805 1270 817 1282
rect 854 1307 866 1319
rect 955 1341 967 1353
rect 894 1307 906 1319
rect 1014 1321 1026 1333
rect 994 1287 1006 1299
rect 1114 1321 1126 1333
rect 1074 1301 1086 1313
rect 1234 1307 1246 1319
rect 1315 1341 1327 1353
rect 1274 1307 1286 1319
rect 1374 1321 1386 1333
rect 1354 1287 1366 1299
rect 1414 1307 1426 1319
rect 1495 1341 1507 1353
rect 1454 1307 1466 1319
rect 1603 1338 1615 1350
rect 1554 1321 1566 1333
rect 1574 1321 1586 1333
rect 1534 1287 1546 1299
rect 1654 1307 1666 1319
rect 1881 1364 1893 1376
rect 1933 1378 1945 1390
rect 1905 1364 1917 1376
rect 1755 1341 1767 1353
rect 1694 1307 1706 1319
rect 1603 1270 1615 1282
rect 1814 1321 1826 1333
rect 1853 1332 1865 1344
rect 1794 1287 1806 1299
rect 1867 1293 1879 1305
rect 1921 1260 1933 1272
rect 1967 1378 1979 1390
rect 1953 1358 1965 1370
rect 1985 1344 1997 1356
rect 2014 1302 2026 1314
rect 2134 1321 2146 1333
rect 1994 1288 2006 1300
rect 1969 1256 1981 1268
rect 1991 1256 2003 1268
rect 2034 1301 2046 1313
rect 2074 1301 2086 1313
rect 2193 1341 2205 1353
rect 2154 1287 2166 1299
rect 2254 1307 2266 1319
rect 2334 1321 2346 1333
rect 2374 1321 2386 1333
rect 2294 1307 2306 1319
rect 2581 1364 2593 1376
rect 2633 1378 2645 1390
rect 2605 1364 2617 1376
rect 2454 1321 2466 1333
rect 2494 1321 2506 1333
rect 2553 1332 2565 1344
rect 2434 1301 2446 1313
rect 2567 1293 2579 1305
rect 2621 1260 2633 1272
rect 2667 1378 2679 1390
rect 2653 1358 2665 1370
rect 2685 1344 2697 1356
rect 2714 1302 2726 1314
rect 2774 1321 2786 1333
rect 2814 1321 2826 1333
rect 2694 1288 2706 1300
rect 2669 1256 2681 1268
rect 2691 1256 2703 1268
rect 2734 1301 2746 1313
rect 2914 1321 2926 1333
rect 2894 1287 2906 1299
rect 2973 1341 2985 1353
rect 2934 1287 2946 1299
rect 3014 1321 3026 1333
rect 3073 1341 3085 1353
rect 3034 1287 3046 1299
rect 3114 1321 3126 1333
rect 3173 1341 3185 1353
rect 3134 1287 3146 1299
rect 3214 1321 3226 1333
rect 3254 1307 3266 1319
rect 3334 1321 3346 1333
rect 3414 1361 3426 1373
rect 3394 1341 3406 1353
rect 3374 1321 3386 1333
rect 3255 1270 3267 1282
rect 3435 1341 3447 1353
rect 3515 1341 3527 1353
rect 3574 1321 3586 1333
rect 3594 1321 3606 1333
rect 3554 1287 3566 1299
rect 3653 1341 3665 1353
rect 3614 1287 3626 1299
rect 3714 1307 3726 1319
rect 3754 1307 3766 1319
rect 3794 1307 3806 1319
rect 3854 1321 3866 1333
rect 3834 1307 3846 1319
rect 3894 1307 3906 1319
rect 3975 1341 3987 1353
rect 3895 1270 3907 1282
rect 4034 1321 4046 1333
rect 4014 1287 4026 1299
rect 4054 1301 4066 1313
rect 4134 1307 4146 1319
rect 4174 1307 4186 1319
rect 4214 1307 4226 1319
rect 4294 1321 4306 1333
rect 4375 1341 4387 1353
rect 4334 1321 4346 1333
rect 4254 1307 4266 1319
rect 4434 1321 4446 1333
rect 4454 1321 4466 1333
rect 4414 1287 4426 1299
rect 4513 1341 4525 1353
rect 4474 1287 4486 1299
rect 4614 1301 4626 1313
rect 4594 1287 4606 1299
rect 4654 1307 4666 1319
rect 4634 1287 4646 1299
rect 4694 1307 4706 1319
rect 14 1107 26 1119
rect 94 1101 106 1113
rect 134 1101 146 1113
rect 214 1121 226 1133
rect 175 1067 187 1079
rect 275 1121 287 1133
rect 313 1121 325 1133
rect 234 1087 246 1099
rect 255 1087 267 1099
rect 414 1121 426 1133
rect 334 1087 346 1099
rect 515 1136 527 1148
rect 454 1121 466 1133
rect 434 1107 446 1119
rect 554 1107 566 1119
rect 534 1087 546 1099
rect 515 1069 527 1081
rect 693 1138 705 1150
rect 574 1087 586 1099
rect 614 1087 626 1099
rect 694 1101 706 1113
rect 785 1138 797 1150
rect 954 1107 966 1119
rect 1014 1107 1026 1119
rect 734 1087 746 1099
rect 814 1087 826 1099
rect 854 1087 866 1099
rect 785 1070 797 1082
rect 894 1087 906 1099
rect 1114 1107 1126 1119
rect 1034 1087 1046 1099
rect 1074 1087 1086 1099
rect 1254 1121 1266 1133
rect 1194 1087 1206 1099
rect 1234 1087 1246 1099
rect 1294 1121 1306 1133
rect 1274 1107 1286 1119
rect 1374 1107 1386 1119
rect 1417 1152 1429 1164
rect 1439 1152 1451 1164
rect 1414 1120 1426 1132
rect 1394 1106 1406 1118
rect 1423 1064 1435 1076
rect 1455 1050 1467 1062
rect 1441 1030 1453 1042
rect 1487 1148 1499 1160
rect 1541 1115 1553 1127
rect 1555 1076 1567 1088
rect 1634 1107 1646 1119
rect 1503 1044 1515 1056
rect 1475 1030 1487 1042
rect 1527 1044 1539 1056
rect 1654 1101 1666 1113
rect 1694 1101 1706 1113
rect 1834 1107 1846 1119
rect 1877 1152 1889 1164
rect 1899 1152 1911 1164
rect 1874 1120 1886 1132
rect 1734 1087 1746 1099
rect 1774 1087 1786 1099
rect 1854 1106 1866 1118
rect 1883 1064 1895 1076
rect 1915 1050 1927 1062
rect 1901 1030 1913 1042
rect 1947 1148 1959 1160
rect 2001 1115 2013 1127
rect 2015 1076 2027 1088
rect 2094 1107 2106 1119
rect 1963 1044 1975 1056
rect 1935 1030 1947 1042
rect 1987 1044 1999 1056
rect 2314 1107 2326 1119
rect 2114 1087 2126 1099
rect 2154 1087 2166 1099
rect 2194 1087 2206 1099
rect 2234 1087 2246 1099
rect 2367 1115 2379 1127
rect 2353 1076 2365 1088
rect 2421 1148 2433 1160
rect 2381 1044 2393 1056
rect 2405 1044 2417 1056
rect 2469 1152 2481 1164
rect 2491 1152 2503 1164
rect 2453 1050 2465 1062
rect 2433 1030 2445 1042
rect 2494 1120 2506 1132
rect 2514 1106 2526 1118
rect 2534 1107 2546 1119
rect 2574 1107 2586 1119
rect 2485 1064 2497 1076
rect 2467 1030 2479 1042
rect 2654 1121 2666 1133
rect 2634 1087 2646 1099
rect 2754 1121 2766 1133
rect 2790 1121 2802 1133
rect 2734 1087 2746 1099
rect 2693 1067 2705 1079
rect 2954 1101 2966 1113
rect 2813 1087 2825 1099
rect 2854 1087 2866 1099
rect 2894 1087 2906 1099
rect 2994 1101 3006 1113
rect 3055 1138 3067 1150
rect 3054 1101 3066 1113
rect 3014 1087 3026 1099
rect 3134 1121 3146 1133
rect 3114 1087 3126 1099
rect 3214 1107 3226 1119
rect 3173 1067 3185 1079
rect 3253 1136 3265 1148
rect 3334 1101 3346 1113
rect 3234 1087 3246 1099
rect 3253 1069 3265 1081
rect 3374 1101 3386 1113
rect 3414 1101 3426 1113
rect 3454 1101 3466 1113
rect 3474 1101 3486 1113
rect 3514 1101 3526 1113
rect 3554 1101 3566 1113
rect 3594 1101 3606 1113
rect 3654 1121 3666 1133
rect 3634 1087 3646 1099
rect 3693 1067 3705 1079
rect 3773 1067 3785 1079
rect 3834 1121 3846 1133
rect 3874 1121 3886 1133
rect 3854 1107 3866 1119
rect 3814 1067 3826 1079
rect 3794 1047 3806 1059
rect 3974 1107 3986 1119
rect 4033 1067 4045 1079
rect 4094 1121 4106 1133
rect 4134 1121 4146 1133
rect 4114 1107 4126 1119
rect 4074 1067 4086 1079
rect 4054 1047 4066 1059
rect 4194 1107 4206 1119
rect 4294 1121 4306 1133
rect 4334 1121 4346 1133
rect 4314 1107 4326 1119
rect 4414 1121 4426 1133
rect 4375 1067 4387 1079
rect 4474 1121 4486 1133
rect 4434 1087 4446 1099
rect 4454 1087 4466 1099
rect 4654 1101 4666 1113
rect 4554 1087 4566 1099
rect 4513 1067 4525 1079
rect 4594 1087 4606 1099
rect 4694 1101 4706 1113
rect 4754 1107 4766 1119
rect 101 898 113 910
rect 83 864 95 876
rect 34 821 46 833
rect 54 822 66 834
rect 74 808 86 820
rect 135 898 147 910
rect 115 878 127 890
rect 77 776 89 788
rect 99 776 111 788
rect 163 884 175 896
rect 187 884 199 896
rect 147 780 159 792
rect 215 852 227 864
rect 201 813 213 825
rect 254 827 266 839
rect 355 861 367 873
rect 294 827 306 839
rect 414 841 426 853
rect 394 807 406 819
rect 521 898 533 910
rect 503 864 515 876
rect 454 821 466 833
rect 474 822 486 834
rect 494 808 506 820
rect 555 898 567 910
rect 535 878 547 890
rect 497 776 509 788
rect 519 776 531 788
rect 583 884 595 896
rect 607 884 619 896
rect 567 780 579 792
rect 635 852 647 864
rect 621 813 633 825
rect 674 827 686 839
rect 775 861 787 873
rect 714 827 726 839
rect 875 861 887 873
rect 834 841 846 853
rect 814 807 826 819
rect 934 841 946 853
rect 914 807 926 819
rect 1034 841 1046 853
rect 1074 841 1086 853
rect 1094 841 1106 853
rect 1134 841 1146 853
rect 994 821 1006 833
rect 1194 827 1206 839
rect 1234 827 1246 839
rect 1274 827 1286 839
rect 1314 827 1326 839
rect 1354 827 1366 839
rect 1394 827 1406 839
rect 1474 821 1486 833
rect 1454 807 1466 819
rect 1494 807 1506 819
rect 1594 841 1606 853
rect 1554 827 1566 839
rect 1553 790 1565 802
rect 1634 821 1646 833
rect 1614 807 1626 819
rect 1654 807 1666 819
rect 1734 807 1746 819
rect 1934 827 1946 839
rect 1770 804 1782 816
rect 1810 804 1822 816
rect 1850 804 1862 816
rect 2014 841 2026 853
rect 2054 841 2066 853
rect 2074 841 2086 853
rect 1974 827 1986 839
rect 2133 861 2145 873
rect 2094 807 2106 819
rect 2174 841 2186 853
rect 2233 861 2245 873
rect 2194 807 2206 819
rect 2274 841 2286 853
rect 2333 861 2345 873
rect 2294 807 2306 819
rect 2374 827 2386 839
rect 2414 827 2426 839
rect 2561 884 2573 896
rect 2613 898 2625 910
rect 2585 884 2597 896
rect 2533 852 2545 864
rect 2494 821 2506 833
rect 2547 813 2559 825
rect 2601 780 2613 792
rect 2647 898 2659 910
rect 2633 878 2645 890
rect 2665 864 2677 876
rect 2694 822 2706 834
rect 2775 861 2787 873
rect 2674 808 2686 820
rect 2649 776 2661 788
rect 2671 776 2683 788
rect 2714 821 2726 833
rect 2834 841 2846 853
rect 2814 807 2826 819
rect 2994 881 3006 893
rect 2974 861 2986 873
rect 2894 821 2906 833
rect 2914 821 2926 833
rect 3015 861 3027 873
rect 3074 821 3086 833
rect 3154 827 3166 839
rect 3194 827 3206 839
rect 3253 859 3265 871
rect 3234 841 3246 853
rect 3214 821 3226 833
rect 3314 827 3326 839
rect 3354 827 3366 839
rect 3394 827 3406 839
rect 3253 792 3265 804
rect 3494 841 3506 853
rect 3534 841 3546 853
rect 3434 827 3446 839
rect 3554 827 3566 839
rect 3694 881 3706 893
rect 3673 861 3685 873
rect 3594 827 3606 839
rect 3794 881 3806 893
rect 3714 861 3726 873
rect 3773 861 3785 873
rect 3814 861 3826 873
rect 3834 827 3846 839
rect 3974 881 3986 893
rect 3953 861 3965 873
rect 3874 827 3886 839
rect 3994 861 4006 873
rect 4095 861 4107 873
rect 4054 821 4066 833
rect 4195 861 4207 873
rect 4154 841 4166 853
rect 4134 807 4146 819
rect 4254 841 4266 853
rect 4234 807 4246 819
rect 4394 881 4406 893
rect 4374 861 4386 873
rect 4334 821 4346 833
rect 4314 807 4326 819
rect 4354 807 4366 819
rect 4415 861 4427 873
rect 4534 881 4546 893
rect 4513 861 4525 873
rect 4554 861 4566 873
rect 4694 881 4706 893
rect 4674 861 4686 873
rect 4634 821 4646 833
rect 4614 807 4626 819
rect 4654 807 4666 819
rect 4715 861 4727 873
rect 34 627 46 639
rect 77 672 89 684
rect 99 672 111 684
rect 74 640 86 652
rect 54 626 66 638
rect 83 584 95 596
rect 115 570 127 582
rect 101 550 113 562
rect 147 668 159 680
rect 201 635 213 647
rect 254 627 266 639
rect 215 596 227 608
rect 163 564 175 576
rect 135 550 147 562
rect 187 564 199 576
rect 334 641 346 653
rect 314 607 326 619
rect 414 621 426 633
rect 373 587 385 599
rect 454 621 466 633
rect 523 658 535 670
rect 494 607 506 619
rect 614 627 626 639
rect 523 590 535 602
rect 667 635 679 647
rect 653 596 665 608
rect 721 668 733 680
rect 681 564 693 576
rect 705 564 717 576
rect 769 672 781 684
rect 791 672 803 684
rect 753 570 765 582
rect 733 550 745 562
rect 794 640 806 652
rect 814 626 826 638
rect 834 627 846 639
rect 785 584 797 596
rect 767 550 779 562
rect 894 641 906 653
rect 874 607 886 619
rect 1054 627 1066 639
rect 994 607 1006 619
rect 933 587 945 599
rect 1034 607 1046 619
rect 1093 656 1105 668
rect 1074 607 1086 619
rect 1093 589 1105 601
rect 1214 641 1226 653
rect 1175 587 1187 599
rect 1293 658 1305 670
rect 1234 607 1246 619
rect 1294 621 1306 633
rect 1463 658 1475 670
rect 1534 627 1546 639
rect 1577 672 1589 684
rect 1599 672 1611 684
rect 1574 640 1586 652
rect 1334 607 1346 619
rect 1354 607 1366 619
rect 1394 607 1406 619
rect 1434 607 1446 619
rect 1463 590 1475 602
rect 1554 626 1566 638
rect 1583 584 1595 596
rect 1615 570 1627 582
rect 1601 550 1613 562
rect 1647 668 1659 680
rect 1701 635 1713 647
rect 1783 658 1795 670
rect 2034 627 2046 639
rect 1715 596 1727 608
rect 1754 607 1766 619
rect 1854 607 1866 619
rect 1663 564 1675 576
rect 1635 550 1647 562
rect 1687 564 1699 576
rect 1783 590 1795 602
rect 1894 607 1906 619
rect 1934 607 1946 619
rect 1974 607 1986 619
rect 2054 607 2066 619
rect 2094 607 2106 619
rect 2167 635 2179 647
rect 2153 596 2165 608
rect 2221 668 2233 680
rect 2181 564 2193 576
rect 2205 564 2217 576
rect 2269 672 2281 684
rect 2291 672 2303 684
rect 2253 570 2265 582
rect 2233 550 2245 562
rect 2294 640 2306 652
rect 2314 626 2326 638
rect 2334 627 2346 639
rect 2285 584 2297 596
rect 2267 550 2279 562
rect 2395 641 2407 653
rect 2433 641 2445 653
rect 2375 607 2387 619
rect 2535 656 2547 668
rect 2634 641 2646 653
rect 2574 627 2586 639
rect 2454 607 2466 619
rect 2554 607 2566 619
rect 2535 589 2547 601
rect 2674 641 2686 653
rect 2734 641 2746 653
rect 2654 627 2666 639
rect 2774 641 2786 653
rect 2754 627 2766 639
rect 2794 627 2806 639
rect 2914 641 2926 653
rect 2875 587 2887 599
rect 2974 641 2986 653
rect 2934 607 2946 619
rect 2954 607 2966 619
rect 3054 621 3066 633
rect 3013 587 3025 599
rect 3094 621 3106 633
rect 3174 627 3186 639
rect 3194 627 3206 639
rect 3293 587 3305 599
rect 3454 641 3466 653
rect 3374 607 3386 619
rect 3334 587 3346 599
rect 3314 567 3326 579
rect 3414 607 3426 619
rect 3434 607 3446 619
rect 3534 641 3546 653
rect 3574 641 3586 653
rect 3554 627 3566 639
rect 3493 587 3505 599
rect 3674 641 3686 653
rect 3714 641 3726 653
rect 3694 627 3706 639
rect 3775 641 3787 653
rect 3813 641 3825 653
rect 3754 607 3766 619
rect 3833 607 3845 619
rect 3893 587 3905 599
rect 3934 587 3946 599
rect 3993 587 4005 599
rect 3914 567 3926 579
rect 4054 627 4066 639
rect 4034 587 4046 599
rect 4014 567 4026 579
rect 4114 587 4126 599
rect 4155 587 4167 599
rect 4214 587 4226 599
rect 4134 567 4146 579
rect 4255 587 4267 599
rect 4234 567 4246 579
rect 4353 587 4365 599
rect 4394 587 4406 599
rect 4453 587 4465 599
rect 4374 567 4386 579
rect 4514 627 4526 639
rect 4494 587 4506 599
rect 4474 567 4486 579
rect 4634 641 4646 653
rect 4595 587 4607 599
rect 4694 641 4706 653
rect 4654 607 4666 619
rect 4674 607 4686 619
rect 4733 587 4745 599
rect 101 418 113 430
rect 83 384 95 396
rect 34 341 46 353
rect 54 342 66 354
rect 74 328 86 340
rect 135 418 147 430
rect 115 398 127 410
rect 77 296 89 308
rect 99 296 111 308
rect 163 404 175 416
rect 187 404 199 416
rect 147 300 159 312
rect 215 372 227 384
rect 201 333 213 345
rect 254 347 266 359
rect 355 381 367 393
rect 294 347 306 359
rect 414 361 426 373
rect 394 327 406 339
rect 434 341 446 353
rect 494 347 506 359
rect 595 381 607 393
rect 534 347 546 359
rect 654 361 666 373
rect 674 361 686 373
rect 634 327 646 339
rect 733 381 745 393
rect 694 327 706 339
rect 774 361 786 373
rect 833 381 845 393
rect 895 381 907 393
rect 794 327 806 339
rect 954 361 966 373
rect 934 327 946 339
rect 974 341 986 353
rect 1034 347 1046 359
rect 1074 347 1086 359
rect 1174 341 1186 353
rect 1154 327 1166 339
rect 1295 381 1307 393
rect 1254 341 1266 353
rect 1194 327 1206 339
rect 1354 361 1366 373
rect 1394 361 1406 373
rect 1434 361 1446 373
rect 1454 361 1466 373
rect 1334 327 1346 339
rect 1513 381 1525 393
rect 1474 327 1486 339
rect 1554 347 1566 359
rect 1681 404 1693 416
rect 1733 418 1745 430
rect 1705 404 1717 416
rect 1653 372 1665 384
rect 1594 347 1606 359
rect 1667 333 1679 345
rect 1721 300 1733 312
rect 1767 418 1779 430
rect 1753 398 1765 410
rect 1785 384 1797 396
rect 1814 342 1826 354
rect 1794 328 1806 340
rect 1769 296 1781 308
rect 1791 296 1803 308
rect 1834 341 1846 353
rect 1894 347 1906 359
rect 1975 381 1987 393
rect 1934 347 1946 359
rect 2034 361 2046 373
rect 2014 327 2026 339
rect 2141 418 2153 430
rect 2123 384 2135 396
rect 2074 341 2086 353
rect 2094 342 2106 354
rect 2114 328 2126 340
rect 2175 418 2187 430
rect 2155 398 2167 410
rect 2117 296 2129 308
rect 2139 296 2151 308
rect 2203 404 2215 416
rect 2227 404 2239 416
rect 2187 300 2199 312
rect 2255 372 2267 384
rect 2241 333 2253 345
rect 2354 361 2366 373
rect 2394 361 2406 373
rect 2334 341 2346 353
rect 2434 341 2446 353
rect 2514 347 2526 359
rect 2621 404 2633 416
rect 2673 418 2685 430
rect 2645 404 2657 416
rect 2593 372 2605 384
rect 2554 347 2566 359
rect 2607 333 2619 345
rect 2661 300 2673 312
rect 2707 418 2719 430
rect 2693 398 2705 410
rect 2725 384 2737 396
rect 2754 342 2766 354
rect 2734 328 2746 340
rect 2709 296 2721 308
rect 2731 296 2743 308
rect 2774 341 2786 353
rect 2814 347 2826 359
rect 2895 361 2907 373
rect 2854 347 2866 359
rect 2974 361 2986 373
rect 3014 361 3026 373
rect 3054 361 3066 373
rect 2915 327 2927 339
rect 2953 327 2965 339
rect 3214 401 3226 413
rect 3193 381 3205 393
rect 3094 341 3106 353
rect 3314 401 3326 413
rect 3234 381 3246 393
rect 3293 381 3305 393
rect 3334 381 3346 393
rect 3354 361 3366 373
rect 3413 381 3425 393
rect 3374 327 3386 339
rect 3494 341 3506 353
rect 3514 347 3526 359
rect 3554 347 3566 359
rect 3594 347 3606 359
rect 3674 361 3686 373
rect 3634 347 3646 359
rect 3733 381 3745 393
rect 3694 327 3706 339
rect 3794 361 3806 373
rect 3834 361 3846 373
rect 3874 361 3886 373
rect 3914 361 3926 373
rect 3934 361 3946 373
rect 3974 347 3986 359
rect 4034 361 4046 373
rect 4074 361 4086 373
rect 3975 310 3987 322
rect 4274 401 4286 413
rect 4253 381 4265 393
rect 4174 341 4186 353
rect 4154 327 4166 339
rect 4194 327 4206 339
rect 4294 381 4306 393
rect 4334 341 4346 353
rect 4314 327 4326 339
rect 4495 381 4507 393
rect 4414 341 4426 353
rect 4354 327 4366 339
rect 4554 361 4566 373
rect 4534 327 4546 339
rect 4574 341 4586 353
rect 4634 341 4646 353
rect 4694 341 4706 353
rect 34 147 46 159
rect 77 192 89 204
rect 99 192 111 204
rect 74 160 86 172
rect 54 146 66 158
rect 83 104 95 116
rect 115 90 127 102
rect 101 70 113 82
rect 147 188 159 200
rect 201 155 213 167
rect 275 161 287 173
rect 313 161 325 173
rect 215 116 227 128
rect 255 127 267 139
rect 595 176 607 188
rect 334 127 346 139
rect 374 127 386 139
rect 414 127 426 139
rect 454 107 466 119
rect 163 84 175 96
rect 135 70 147 82
rect 187 84 199 96
rect 694 161 706 173
rect 634 147 646 159
rect 614 127 626 139
rect 495 107 507 119
rect 474 87 486 99
rect 595 109 607 121
rect 734 161 746 173
rect 714 147 726 159
rect 787 155 799 167
rect 773 116 785 128
rect 841 188 853 200
rect 801 84 813 96
rect 825 84 837 96
rect 889 192 901 204
rect 911 192 923 204
rect 873 90 885 102
rect 853 70 865 82
rect 914 160 926 172
rect 934 146 946 158
rect 954 147 966 159
rect 905 104 917 116
rect 887 70 899 82
rect 1054 161 1066 173
rect 1015 107 1027 119
rect 1134 147 1146 159
rect 1074 127 1086 139
rect 1274 147 1286 159
rect 1174 127 1186 139
rect 1214 127 1226 139
rect 1354 161 1366 173
rect 1315 107 1327 119
rect 1434 147 1446 159
rect 1494 147 1506 159
rect 1374 127 1386 139
rect 1634 161 1646 173
rect 1514 127 1526 139
rect 1554 127 1566 139
rect 1674 161 1686 173
rect 1654 147 1666 159
rect 1714 147 1726 159
rect 1757 192 1769 204
rect 1779 192 1791 204
rect 1754 160 1766 172
rect 1734 146 1746 158
rect 1763 104 1775 116
rect 1795 90 1807 102
rect 1781 70 1793 82
rect 1827 188 1839 200
rect 1881 155 1893 167
rect 1895 116 1907 128
rect 1994 161 2006 173
rect 1955 107 1967 119
rect 1843 84 1855 96
rect 1815 70 1827 82
rect 1867 84 1879 96
rect 2034 147 2046 159
rect 2014 127 2026 139
rect 2454 147 2466 159
rect 2094 127 2106 139
rect 2134 127 2146 139
rect 2174 127 2186 139
rect 2214 127 2226 139
rect 2274 127 2286 139
rect 2314 127 2326 139
rect 2334 127 2346 139
rect 2374 127 2386 139
rect 2507 155 2519 167
rect 2493 116 2505 128
rect 2561 188 2573 200
rect 2521 84 2533 96
rect 2545 84 2557 96
rect 2609 192 2621 204
rect 2631 192 2643 204
rect 2593 90 2605 102
rect 2573 70 2585 82
rect 2634 160 2646 172
rect 2654 146 2666 158
rect 2674 147 2686 159
rect 2625 104 2637 116
rect 2607 70 2619 82
rect 2747 155 2759 167
rect 2733 116 2745 128
rect 2801 188 2813 200
rect 2761 84 2773 96
rect 2785 84 2797 96
rect 2849 192 2861 204
rect 2871 192 2883 204
rect 2833 90 2845 102
rect 2813 70 2825 82
rect 2874 160 2886 172
rect 2894 146 2906 158
rect 2914 147 2926 159
rect 2865 104 2877 116
rect 2847 70 2859 82
rect 2974 161 2986 173
rect 3010 161 3022 173
rect 2954 127 2966 139
rect 3115 176 3127 188
rect 3154 147 3166 159
rect 3033 127 3045 139
rect 3134 127 3146 139
rect 3115 109 3127 121
rect 3194 161 3206 173
rect 3174 127 3186 139
rect 3314 147 3326 159
rect 3233 107 3245 119
rect 3334 141 3346 153
rect 3374 141 3386 153
rect 3453 107 3465 119
rect 3614 161 3626 173
rect 3554 147 3566 159
rect 3494 107 3506 119
rect 3474 87 3486 99
rect 3654 161 3666 173
rect 3634 147 3646 159
rect 3754 147 3766 159
rect 3694 127 3706 139
rect 3734 127 3746 139
rect 3834 161 3846 173
rect 3814 127 3826 139
rect 3914 127 3926 139
rect 3873 107 3885 119
rect 3954 127 3966 139
rect 4033 107 4045 119
rect 4094 141 4106 153
rect 4074 107 4086 119
rect 4054 87 4066 99
rect 4134 141 4146 153
rect 4213 107 4225 119
rect 4294 141 4306 153
rect 4254 107 4266 119
rect 4234 87 4246 99
rect 4334 141 4346 153
rect 4393 107 4405 119
rect 4454 141 4466 153
rect 4434 107 4446 119
rect 4414 87 4426 99
rect 4494 141 4506 153
rect 4534 107 4546 119
rect 4674 161 4686 173
rect 4575 107 4587 119
rect 4554 87 4566 99
rect 4714 161 4726 173
rect 4694 147 4706 159
<< metal1 >>
rect -62 4338 -2 4578
rect 4 4576 4842 4578
rect 4776 4564 4842 4576
rect 4 4562 4842 4564
rect 49 4556 61 4562
rect 149 4556 161 4562
rect 231 4556 243 4562
rect 299 4556 311 4562
rect 371 4556 383 4562
rect 411 4556 423 4562
rect 31 4473 39 4516
rect 71 4510 79 4536
rect 57 4504 79 4510
rect 119 4508 131 4516
rect 57 4498 60 4504
rect 119 4502 143 4508
rect 31 4459 33 4473
rect 31 4424 39 4459
rect 53 4442 60 4498
rect 135 4453 143 4502
rect 195 4502 203 4516
rect 223 4516 251 4522
rect 211 4513 263 4516
rect 281 4510 289 4536
rect 451 4556 463 4562
rect 491 4556 503 4562
rect 539 4556 551 4562
rect 631 4556 643 4562
rect 281 4504 303 4510
rect 195 4495 220 4502
rect 300 4498 303 4504
rect 213 4473 221 4495
rect 57 4436 60 4442
rect 57 4430 83 4436
rect 75 4384 83 4430
rect 135 4384 143 4439
rect 219 4424 227 4459
rect 300 4442 307 4498
rect 321 4473 329 4516
rect 393 4493 400 4536
rect 473 4493 480 4536
rect 521 4510 529 4536
rect 657 4556 669 4562
rect 697 4556 709 4562
rect 737 4556 749 4562
rect 819 4556 831 4562
rect 877 4556 889 4562
rect 925 4556 937 4562
rect 987 4556 999 4562
rect 1057 4556 1069 4562
rect 1159 4556 1171 4562
rect 1217 4556 1229 4562
rect 1265 4556 1277 4562
rect 1327 4556 1339 4562
rect 1397 4556 1409 4562
rect 1501 4556 1513 4562
rect 1563 4556 1575 4562
rect 1611 4556 1623 4562
rect 1669 4556 1681 4562
rect 1719 4556 1731 4562
rect 1819 4556 1831 4562
rect 1877 4556 1889 4562
rect 1925 4556 1937 4562
rect 1987 4556 1999 4562
rect 2057 4556 2069 4562
rect 2230 4556 2242 4562
rect 2311 4556 2323 4562
rect 2391 4556 2403 4562
rect 521 4504 543 4510
rect 540 4498 543 4504
rect 327 4459 329 4473
rect 300 4436 303 4442
rect 277 4430 303 4436
rect 49 4338 61 4344
rect 111 4338 123 4344
rect 151 4338 163 4344
rect 277 4384 285 4430
rect 321 4424 329 4459
rect 393 4431 400 4479
rect 473 4431 480 4479
rect 540 4442 547 4498
rect 561 4473 569 4516
rect 616 4481 624 4536
rect 680 4493 687 4536
rect 567 4459 569 4473
rect 756 4481 764 4536
rect 967 4536 980 4542
rect 851 4530 858 4536
rect 847 4522 858 4530
rect 908 4524 915 4536
rect 973 4530 980 4536
rect 797 4501 805 4516
rect 908 4517 929 4524
rect 887 4506 893 4508
rect 954 4506 961 4512
rect 797 4487 813 4501
rect 887 4500 961 4506
rect 540 4436 543 4442
rect 383 4424 400 4431
rect 463 4424 480 4431
rect 517 4430 543 4436
rect 517 4384 525 4430
rect 561 4424 569 4459
rect 616 4384 624 4467
rect 680 4431 687 4479
rect 680 4424 697 4431
rect 196 4338 208 4344
rect 246 4338 258 4344
rect 299 4338 311 4344
rect 411 4338 423 4344
rect 491 4338 503 4344
rect 539 4338 551 4344
rect 631 4338 643 4344
rect 756 4384 764 4467
rect 797 4424 805 4487
rect 813 4473 827 4487
rect 819 4428 833 4436
rect 887 4428 893 4500
rect 954 4492 961 4500
rect 966 4484 1000 4492
rect 994 4479 1000 4484
rect 947 4466 974 4473
rect 853 4422 893 4428
rect 901 4428 945 4434
rect 853 4404 859 4422
rect 901 4414 907 4428
rect 1013 4432 1019 4516
rect 1049 4516 1077 4522
rect 1037 4513 1089 4516
rect 1307 4536 1320 4542
rect 1191 4530 1198 4536
rect 1187 4522 1198 4530
rect 1248 4524 1255 4536
rect 1313 4530 1320 4536
rect 1097 4502 1105 4516
rect 1080 4495 1105 4502
rect 1137 4501 1145 4516
rect 1248 4517 1269 4524
rect 1227 4506 1233 4508
rect 1294 4506 1301 4512
rect 1079 4473 1087 4495
rect 1137 4487 1153 4501
rect 1227 4500 1301 4506
rect 957 4424 1019 4432
rect 1073 4424 1081 4459
rect 1137 4424 1145 4487
rect 1153 4473 1167 4487
rect 1159 4428 1173 4436
rect 877 4408 907 4414
rect 925 4410 963 4418
rect 955 4404 963 4410
rect 847 4364 859 4398
rect 905 4390 927 4402
rect 955 4390 973 4404
rect 901 4384 913 4390
rect 955 4384 963 4390
rect 1227 4428 1233 4500
rect 1294 4492 1301 4500
rect 1306 4484 1340 4492
rect 1334 4479 1340 4484
rect 1287 4466 1314 4473
rect 1193 4422 1233 4428
rect 1241 4428 1285 4434
rect 1193 4404 1199 4422
rect 1241 4414 1247 4428
rect 1353 4432 1359 4516
rect 1389 4516 1417 4522
rect 1377 4513 1429 4516
rect 1520 4536 1533 4542
rect 1520 4530 1527 4536
rect 1585 4524 1592 4536
rect 1437 4502 1445 4516
rect 1420 4495 1445 4502
rect 1419 4473 1427 4495
rect 1297 4424 1359 4432
rect 1413 4424 1421 4459
rect 1481 4432 1487 4516
rect 1571 4517 1592 4524
rect 1642 4530 1649 4536
rect 1642 4522 1653 4530
rect 1539 4506 1546 4512
rect 1607 4506 1613 4508
rect 1539 4500 1613 4506
rect 1695 4501 1703 4516
rect 1749 4508 1761 4516
rect 1539 4492 1546 4500
rect 1500 4484 1534 4492
rect 1500 4479 1506 4484
rect 1526 4466 1553 4473
rect 1481 4424 1543 4432
rect 1555 4428 1599 4434
rect 1217 4408 1247 4414
rect 1265 4410 1303 4418
rect 1295 4404 1303 4410
rect 1187 4364 1199 4398
rect 1245 4390 1267 4402
rect 1295 4390 1313 4404
rect 1241 4384 1253 4390
rect 1295 4384 1303 4390
rect 1537 4410 1575 4418
rect 1593 4414 1599 4428
rect 1607 4428 1613 4500
rect 1687 4487 1703 4501
rect 1673 4473 1687 4487
rect 1607 4422 1647 4428
rect 1667 4428 1681 4436
rect 1695 4424 1703 4487
rect 1737 4502 1761 4508
rect 1967 4536 1980 4542
rect 1851 4530 1858 4536
rect 1847 4522 1858 4530
rect 1908 4524 1915 4536
rect 1973 4530 1980 4536
rect 1737 4453 1745 4502
rect 1797 4501 1805 4516
rect 1908 4517 1929 4524
rect 1887 4506 1893 4508
rect 1954 4506 1961 4512
rect 1797 4487 1813 4501
rect 1887 4500 1961 4506
rect 1537 4404 1545 4410
rect 1593 4408 1623 4414
rect 1641 4404 1647 4422
rect 1527 4390 1545 4404
rect 1573 4390 1595 4402
rect 1537 4384 1545 4390
rect 1587 4384 1599 4390
rect 1641 4364 1653 4398
rect 1737 4384 1745 4439
rect 1797 4424 1805 4487
rect 1813 4473 1827 4487
rect 1819 4428 1833 4436
rect 1887 4428 1893 4500
rect 1954 4492 1961 4500
rect 1966 4484 2000 4492
rect 1994 4479 2000 4484
rect 1947 4466 1974 4473
rect 1853 4422 1893 4428
rect 1901 4428 1945 4434
rect 1853 4404 1859 4422
rect 1901 4414 1907 4428
rect 2013 4432 2019 4516
rect 2049 4516 2077 4520
rect 2089 4550 2117 4556
rect 2037 4514 2089 4516
rect 2099 4506 2105 4516
rect 2076 4499 2105 4506
rect 2076 4473 2084 4499
rect 2176 4498 2194 4500
rect 2176 4489 2206 4498
rect 2275 4502 2283 4516
rect 2303 4516 2331 4522
rect 2417 4556 2429 4562
rect 2457 4556 2469 4562
rect 2531 4556 2543 4562
rect 2577 4556 2589 4562
rect 2679 4556 2691 4562
rect 2759 4556 2771 4562
rect 2849 4556 2861 4562
rect 2970 4556 2982 4562
rect 3041 4556 3053 4562
rect 3129 4556 3141 4562
rect 3250 4556 3262 4562
rect 2291 4513 2343 4516
rect 2275 4495 2300 4502
rect 2176 4461 2184 4489
rect 2293 4473 2301 4495
rect 2376 4481 2384 4536
rect 2440 4493 2447 4536
rect 1957 4424 2019 4432
rect 2077 4424 2085 4459
rect 2516 4481 2524 4536
rect 2569 4516 2597 4522
rect 2557 4513 2609 4516
rect 2617 4502 2625 4516
rect 2661 4510 2669 4536
rect 2661 4504 2683 4510
rect 2600 4495 2625 4502
rect 2680 4498 2683 4504
rect 1877 4408 1907 4414
rect 1925 4410 1963 4418
rect 1955 4404 1963 4410
rect 1847 4364 1859 4398
rect 1905 4390 1927 4402
rect 1955 4390 1973 4404
rect 1901 4384 1913 4390
rect 1955 4384 1963 4390
rect 2175 4392 2182 4447
rect 2299 4424 2307 4459
rect 2175 4386 2222 4392
rect 2175 4384 2183 4386
rect 2211 4384 2222 4386
rect 657 4338 669 4344
rect 737 4338 749 4344
rect 817 4338 829 4344
rect 875 4338 887 4344
rect 921 4338 933 4344
rect 987 4338 999 4344
rect 1042 4338 1054 4344
rect 1092 4338 1104 4344
rect 1157 4338 1169 4344
rect 1215 4338 1227 4344
rect 1261 4338 1273 4344
rect 1327 4338 1339 4344
rect 1382 4338 1394 4344
rect 1432 4338 1444 4344
rect 1501 4338 1513 4344
rect 1567 4338 1579 4344
rect 1613 4338 1625 4344
rect 1671 4338 1683 4344
rect 1717 4338 1729 4344
rect 1757 4338 1769 4344
rect 1817 4338 1829 4344
rect 1875 4338 1887 4344
rect 1921 4338 1933 4344
rect 1987 4338 1999 4344
rect 2037 4338 2049 4344
rect 2107 4338 2119 4344
rect 2191 4338 2203 4344
rect 2231 4338 2243 4344
rect 2376 4384 2384 4467
rect 2440 4431 2447 4479
rect 2440 4424 2457 4431
rect 2276 4338 2288 4344
rect 2326 4338 2338 4344
rect 2391 4338 2403 4344
rect 2516 4384 2524 4467
rect 2599 4473 2607 4495
rect 2593 4424 2601 4459
rect 2680 4442 2687 4498
rect 2701 4473 2709 4516
rect 2741 4510 2749 4536
rect 2741 4504 2763 4510
rect 2760 4498 2763 4504
rect 2707 4459 2709 4473
rect 2680 4436 2683 4442
rect 2657 4430 2683 4436
rect 2417 4338 2429 4344
rect 2531 4338 2543 4344
rect 2657 4384 2665 4430
rect 2701 4424 2709 4459
rect 2760 4442 2767 4498
rect 2781 4473 2789 4516
rect 2787 4459 2789 4473
rect 2760 4436 2763 4442
rect 2737 4430 2763 4436
rect 2737 4384 2745 4430
rect 2781 4424 2789 4459
rect 2831 4473 2839 4516
rect 2871 4510 2879 4536
rect 2857 4504 2879 4510
rect 2857 4498 2860 4504
rect 2831 4459 2833 4473
rect 2831 4424 2839 4459
rect 2853 4442 2860 4498
rect 2916 4498 2934 4500
rect 2916 4489 2946 4498
rect 3011 4516 3021 4526
rect 2916 4461 2924 4489
rect 3011 4473 3019 4516
rect 3071 4506 3083 4516
rect 3045 4498 3083 4506
rect 3011 4459 3013 4473
rect 2857 4436 2860 4442
rect 2857 4430 2883 4436
rect 2875 4384 2883 4430
rect 2915 4392 2922 4447
rect 3011 4424 3019 4459
rect 2915 4386 2962 4392
rect 2915 4384 2923 4386
rect 2951 4384 2962 4386
rect 3054 4384 3062 4498
rect 3111 4473 3119 4516
rect 3151 4510 3159 4536
rect 3137 4504 3159 4510
rect 3137 4498 3140 4504
rect 3111 4459 3113 4473
rect 3111 4424 3119 4459
rect 3133 4442 3140 4498
rect 3196 4498 3214 4500
rect 3196 4489 3226 4498
rect 3279 4556 3291 4562
rect 3360 4556 3372 4562
rect 3410 4556 3422 4562
rect 3457 4556 3469 4562
rect 3519 4556 3531 4562
rect 3598 4556 3610 4562
rect 3700 4556 3712 4562
rect 3750 4556 3762 4562
rect 3817 4556 3829 4562
rect 3951 4556 3963 4562
rect 4070 4556 4082 4562
rect 4170 4556 4182 4562
rect 3400 4516 3426 4527
rect 3309 4508 3321 4516
rect 3297 4502 3321 4508
rect 3196 4461 3204 4489
rect 3137 4436 3140 4442
rect 3137 4430 3163 4436
rect 3155 4384 3163 4430
rect 3195 4392 3202 4447
rect 3297 4453 3305 4502
rect 3418 4473 3426 4516
rect 3437 4517 3453 4523
rect 3195 4386 3242 4392
rect 3195 4384 3203 4386
rect 3231 4384 3242 4386
rect 3297 4384 3305 4439
rect 3418 4424 3426 4459
rect 3437 4443 3443 4517
rect 3476 4481 3484 4536
rect 3549 4508 3561 4516
rect 3537 4502 3561 4508
rect 3437 4437 3453 4443
rect 3357 4418 3397 4424
rect 3357 4416 3369 4418
rect 2562 4338 2574 4344
rect 2612 4338 2624 4344
rect 2679 4338 2691 4344
rect 2759 4338 2771 4344
rect 2849 4338 2861 4344
rect 2931 4338 2943 4344
rect 2971 4338 2983 4344
rect 3027 4338 3039 4344
rect 3071 4338 3083 4344
rect 3129 4338 3141 4344
rect 3211 4338 3223 4344
rect 3251 4338 3263 4344
rect 3476 4384 3484 4467
rect 3537 4453 3545 4502
rect 3740 4516 3766 4527
rect 3646 4498 3664 4500
rect 3634 4489 3664 4498
rect 3656 4461 3664 4489
rect 3758 4473 3766 4516
rect 3809 4516 3837 4522
rect 3797 4513 3849 4516
rect 3857 4502 3865 4516
rect 3840 4495 3865 4502
rect 3915 4502 3923 4516
rect 3943 4516 3971 4522
rect 3931 4513 3983 4516
rect 3915 4495 3940 4502
rect 4016 4498 4034 4500
rect 3839 4473 3847 4495
rect 3933 4473 3941 4495
rect 4016 4489 4046 4498
rect 4116 4498 4134 4500
rect 4116 4489 4146 4498
rect 4200 4556 4212 4562
rect 4250 4556 4262 4562
rect 4299 4556 4311 4562
rect 4398 4556 4410 4562
rect 4448 4556 4460 4562
rect 4511 4556 4523 4562
rect 4240 4516 4266 4527
rect 4016 4461 4024 4489
rect 4116 4461 4124 4489
rect 4258 4473 4266 4516
rect 4329 4508 4341 4516
rect 4317 4502 4341 4508
rect 4394 4516 4420 4527
rect 4538 4556 4550 4562
rect 4638 4556 4650 4562
rect 3537 4384 3545 4439
rect 3658 4392 3665 4447
rect 3758 4424 3766 4459
rect 3833 4424 3841 4459
rect 3939 4424 3947 4459
rect 3618 4386 3665 4392
rect 3618 4384 3629 4386
rect 3277 4338 3289 4344
rect 3317 4338 3329 4344
rect 3377 4338 3389 4344
rect 3457 4338 3469 4344
rect 3517 4338 3529 4344
rect 3557 4338 3569 4344
rect 3657 4384 3665 4386
rect 3697 4418 3737 4424
rect 3697 4416 3709 4418
rect 3597 4338 3609 4344
rect 3637 4338 3649 4344
rect 3717 4338 3729 4344
rect 3802 4338 3814 4344
rect 3852 4338 3864 4344
rect 4015 4392 4022 4447
rect 4115 4392 4122 4447
rect 4258 4424 4266 4459
rect 4317 4453 4325 4502
rect 4394 4473 4402 4516
rect 4496 4481 4504 4536
rect 4586 4498 4604 4500
rect 4574 4489 4604 4498
rect 4686 4498 4704 4500
rect 4674 4489 4704 4498
rect 4197 4418 4237 4424
rect 4197 4416 4209 4418
rect 4015 4386 4062 4392
rect 4015 4384 4023 4386
rect 4051 4384 4062 4386
rect 4115 4386 4162 4392
rect 4115 4384 4123 4386
rect 4151 4384 4162 4386
rect 4317 4384 4325 4439
rect 4394 4424 4402 4459
rect 4423 4418 4463 4424
rect 4451 4416 4463 4418
rect 4496 4384 4504 4467
rect 4596 4461 4604 4489
rect 4696 4461 4704 4489
rect 4598 4392 4605 4447
rect 4698 4392 4705 4447
rect 4558 4386 4605 4392
rect 4558 4384 4569 4386
rect 3916 4338 3928 4344
rect 3966 4338 3978 4344
rect 4031 4338 4043 4344
rect 4071 4338 4083 4344
rect 4131 4338 4143 4344
rect 4171 4338 4183 4344
rect 4217 4338 4229 4344
rect 4297 4338 4309 4344
rect 4337 4338 4349 4344
rect 4431 4338 4443 4344
rect 4511 4338 4523 4344
rect 4597 4384 4605 4386
rect 4658 4386 4705 4392
rect 4658 4384 4669 4386
rect 4697 4384 4705 4386
rect 4537 4338 4549 4344
rect 4577 4338 4589 4344
rect 4637 4338 4649 4344
rect 4677 4338 4689 4344
rect -62 4336 4776 4338
rect -62 4324 4 4336
rect -62 4322 4776 4324
rect -62 3858 -2 4322
rect 36 4316 48 4322
rect 86 4316 98 4322
rect 147 4316 159 4322
rect 191 4316 203 4322
rect 217 4316 229 4322
rect 351 4316 363 4322
rect 397 4316 409 4322
rect 441 4316 453 4322
rect 551 4316 563 4322
rect 597 4316 609 4322
rect 637 4316 649 4322
rect 717 4316 729 4322
rect 797 4316 809 4322
rect 841 4316 853 4322
rect 916 4316 928 4322
rect 966 4316 978 4322
rect 1031 4316 1043 4322
rect 59 4201 67 4236
rect 131 4201 139 4236
rect 53 4165 61 4187
rect 131 4187 133 4201
rect 35 4158 60 4165
rect 35 4144 43 4158
rect 51 4144 103 4147
rect 63 4138 91 4144
rect 131 4144 139 4187
rect 174 4162 182 4276
rect 371 4242 383 4244
rect 343 4236 383 4242
rect 240 4229 257 4236
rect 240 4181 247 4229
rect 314 4201 322 4236
rect 165 4154 203 4162
rect 191 4144 203 4154
rect 131 4134 141 4144
rect 240 4124 247 4167
rect 314 4144 322 4187
rect 418 4162 426 4276
rect 618 4274 629 4276
rect 657 4274 665 4276
rect 618 4268 665 4274
rect 571 4242 583 4244
rect 543 4236 583 4242
rect 461 4201 469 4236
rect 514 4201 522 4236
rect 658 4213 665 4268
rect 697 4242 709 4244
rect 697 4236 737 4242
rect 467 4187 469 4201
rect 758 4201 766 4236
rect 397 4154 435 4162
rect 397 4144 409 4154
rect 461 4144 469 4187
rect 314 4133 340 4144
rect 71 4098 83 4104
rect 161 4098 173 4104
rect 217 4098 229 4104
rect 257 4098 269 4104
rect 459 4134 469 4144
rect 514 4144 522 4187
rect 656 4171 664 4199
rect 514 4133 540 4144
rect 318 4098 330 4104
rect 368 4098 380 4104
rect 427 4098 439 4104
rect 518 4098 530 4104
rect 568 4098 580 4104
rect 634 4162 664 4171
rect 646 4160 664 4162
rect 758 4144 766 4187
rect 818 4162 826 4276
rect 1057 4316 1069 4322
rect 1137 4316 1149 4322
rect 1217 4316 1229 4322
rect 1297 4316 1309 4322
rect 1377 4316 1389 4322
rect 1435 4316 1447 4322
rect 1481 4316 1493 4322
rect 1547 4316 1559 4322
rect 1602 4316 1614 4322
rect 1652 4316 1664 4322
rect 861 4201 869 4236
rect 939 4201 947 4236
rect 867 4187 869 4201
rect 740 4133 766 4144
rect 797 4154 835 4162
rect 797 4144 809 4154
rect 861 4144 869 4187
rect 933 4165 941 4187
rect 1016 4193 1024 4276
rect 1080 4229 1097 4236
rect 1160 4229 1177 4236
rect 1080 4181 1087 4229
rect 1160 4181 1167 4229
rect 915 4158 940 4165
rect 915 4144 923 4158
rect 859 4134 869 4144
rect 931 4144 983 4147
rect 943 4138 971 4144
rect 1016 4124 1024 4179
rect 1080 4124 1087 4167
rect 1160 4124 1167 4167
rect 1197 4163 1203 4233
rect 1240 4229 1257 4236
rect 1240 4181 1247 4229
rect 1316 4193 1324 4276
rect 1407 4262 1419 4296
rect 1461 4270 1473 4276
rect 1515 4270 1523 4276
rect 1465 4258 1487 4270
rect 1515 4256 1533 4270
rect 1413 4238 1419 4256
rect 1437 4246 1467 4252
rect 1515 4250 1523 4256
rect 1187 4157 1203 4163
rect 1240 4124 1247 4167
rect 1316 4124 1324 4179
rect 1357 4173 1365 4236
rect 1379 4224 1393 4232
rect 1413 4232 1453 4238
rect 1373 4173 1387 4187
rect 1357 4159 1373 4173
rect 1447 4160 1453 4232
rect 1461 4232 1467 4246
rect 1485 4242 1523 4250
rect 1697 4316 1709 4322
rect 1811 4316 1823 4322
rect 1857 4316 1869 4322
rect 1915 4316 1927 4322
rect 1961 4316 1973 4322
rect 2027 4316 2039 4322
rect 2091 4316 2103 4322
rect 2131 4316 2143 4322
rect 2187 4316 2199 4322
rect 2331 4316 2343 4322
rect 2377 4316 2389 4322
rect 2417 4316 2429 4322
rect 1461 4226 1505 4232
rect 1517 4228 1579 4236
rect 1507 4187 1534 4194
rect 1554 4176 1560 4181
rect 1526 4168 1560 4176
rect 1514 4160 1521 4168
rect 1357 4144 1365 4159
rect 1447 4154 1521 4160
rect 1447 4152 1453 4154
rect 598 4098 610 4104
rect 700 4098 712 4104
rect 750 4098 762 4104
rect 827 4098 839 4104
rect 951 4098 963 4104
rect 1031 4098 1043 4104
rect 1057 4098 1069 4104
rect 1097 4098 1109 4104
rect 1137 4098 1149 4104
rect 1177 4098 1189 4104
rect 1217 4098 1229 4104
rect 1257 4098 1269 4104
rect 1514 4148 1521 4154
rect 1407 4130 1418 4138
rect 1411 4124 1418 4130
rect 1468 4136 1489 4143
rect 1573 4144 1579 4228
rect 1633 4201 1641 4236
rect 1720 4229 1737 4236
rect 1639 4165 1647 4187
rect 1720 4181 1727 4229
rect 1796 4193 1804 4276
rect 1887 4262 1899 4296
rect 1941 4270 1953 4276
rect 1995 4270 2003 4276
rect 1945 4258 1967 4270
rect 1995 4256 2013 4270
rect 1893 4238 1899 4256
rect 1917 4246 1947 4252
rect 1995 4250 2003 4256
rect 1640 4158 1665 4165
rect 1468 4124 1475 4136
rect 1533 4124 1540 4130
rect 1527 4118 1540 4124
rect 1597 4144 1649 4147
rect 1609 4138 1637 4144
rect 1657 4144 1665 4158
rect 1720 4124 1727 4167
rect 1796 4124 1804 4179
rect 1837 4173 1845 4236
rect 1859 4224 1873 4232
rect 1893 4232 1933 4238
rect 1853 4173 1867 4187
rect 1837 4159 1853 4173
rect 1927 4160 1933 4232
rect 1941 4232 1947 4246
rect 1965 4242 2003 4250
rect 1941 4226 1985 4232
rect 1997 4228 2059 4236
rect 1987 4187 2014 4194
rect 2034 4176 2040 4181
rect 2006 4168 2040 4176
rect 1994 4160 2001 4168
rect 1837 4144 1845 4159
rect 1927 4154 2001 4160
rect 1927 4152 1933 4154
rect 1994 4148 2001 4154
rect 1887 4130 1898 4138
rect 1891 4124 1898 4130
rect 1948 4136 1969 4143
rect 2053 4144 2059 4228
rect 2115 4221 2123 4276
rect 2219 4237 2223 4246
rect 2157 4228 2165 4236
rect 2157 4220 2193 4228
rect 2115 4158 2123 4207
rect 2198 4164 2204 4219
rect 2214 4193 2223 4237
rect 2283 4310 2311 4316
rect 2323 4238 2351 4244
rect 2476 4316 2488 4322
rect 2526 4316 2538 4322
rect 2611 4316 2623 4322
rect 2657 4316 2669 4322
rect 2791 4316 2803 4322
rect 2859 4316 2871 4322
rect 2951 4316 2963 4322
rect 2991 4316 3003 4322
rect 3051 4316 3063 4322
rect 3091 4316 3103 4322
rect 2292 4230 2304 4236
rect 2292 4224 2319 4230
rect 2313 4201 2319 4224
rect 2397 4221 2405 4276
rect 2637 4242 2649 4244
rect 2637 4236 2677 4242
rect 2811 4242 2823 4244
rect 2783 4236 2823 4242
rect 1948 4124 1955 4136
rect 2013 4124 2020 4130
rect 2007 4118 2020 4124
rect 2099 4152 2123 4158
rect 2183 4152 2193 4158
rect 2099 4144 2111 4152
rect 2183 4124 2189 4152
rect 2220 4144 2227 4179
rect 2320 4144 2327 4187
rect 2397 4158 2405 4207
rect 2499 4201 2507 4236
rect 2583 4229 2600 4236
rect 2493 4165 2501 4187
rect 2593 4181 2600 4229
rect 2698 4201 2706 4236
rect 2754 4201 2762 4236
rect 2837 4230 2845 4276
rect 2935 4274 2943 4276
rect 2971 4274 2982 4276
rect 2935 4268 2982 4274
rect 3035 4274 3043 4276
rect 3117 4316 3129 4322
rect 3157 4316 3169 4322
rect 3231 4316 3243 4322
rect 3291 4316 3303 4322
rect 3331 4316 3343 4322
rect 3391 4316 3403 4322
rect 3431 4316 3443 4322
rect 3491 4316 3503 4322
rect 3531 4316 3543 4322
rect 3591 4316 3603 4322
rect 3631 4316 3643 4322
rect 3071 4274 3082 4276
rect 3035 4268 3082 4274
rect 2837 4224 2863 4230
rect 2860 4218 2863 4224
rect 2475 4158 2500 4165
rect 2397 4152 2421 4158
rect 2409 4144 2421 4152
rect 2475 4144 2483 4158
rect 1297 4098 1309 4104
rect 1379 4098 1391 4104
rect 1437 4098 1449 4104
rect 1485 4098 1497 4104
rect 1547 4098 1559 4104
rect 1617 4098 1629 4104
rect 1697 4098 1709 4104
rect 1737 4098 1749 4104
rect 1811 4098 1823 4104
rect 1859 4098 1871 4104
rect 1917 4098 1929 4104
rect 1965 4098 1977 4104
rect 2027 4098 2039 4104
rect 2129 4098 2141 4104
rect 2157 4098 2165 4104
rect 2197 4098 2209 4104
rect 2292 4098 2304 4104
rect 2348 4098 2360 4104
rect 2491 4144 2543 4147
rect 2503 4138 2531 4144
rect 2593 4124 2600 4167
rect 2698 4144 2706 4187
rect 2379 4098 2391 4104
rect 2511 4098 2523 4104
rect 2571 4098 2583 4104
rect 2611 4098 2623 4104
rect 2680 4133 2706 4144
rect 2754 4144 2762 4187
rect 2860 4162 2867 4218
rect 2881 4201 2889 4236
rect 2935 4213 2942 4268
rect 3007 4257 3023 4263
rect 2887 4187 2889 4201
rect 2860 4156 2863 4162
rect 2841 4150 2863 4156
rect 2754 4133 2780 4144
rect 2640 4098 2652 4104
rect 2690 4098 2702 4104
rect 2841 4124 2849 4150
rect 2881 4144 2889 4187
rect 2936 4171 2944 4199
rect 3017 4183 3023 4257
rect 3035 4213 3042 4268
rect 3137 4221 3145 4276
rect 3007 4177 3023 4183
rect 3036 4171 3044 4199
rect 2936 4162 2966 4171
rect 2936 4160 2954 4162
rect 3036 4162 3066 4171
rect 3036 4160 3054 4162
rect 3137 4158 3145 4207
rect 3216 4193 3224 4276
rect 3275 4274 3283 4276
rect 3311 4274 3322 4276
rect 3275 4268 3322 4274
rect 3375 4274 3383 4276
rect 3411 4274 3422 4276
rect 3375 4268 3422 4274
rect 3475 4274 3483 4276
rect 3511 4274 3522 4276
rect 3475 4268 3522 4274
rect 3575 4274 3583 4276
rect 3657 4316 3669 4322
rect 3697 4316 3709 4322
rect 3777 4316 3789 4322
rect 3862 4316 3874 4322
rect 3912 4316 3924 4322
rect 3611 4274 3622 4276
rect 3575 4268 3622 4274
rect 3678 4274 3689 4276
rect 3717 4274 3725 4276
rect 3678 4268 3725 4274
rect 3275 4213 3282 4268
rect 3137 4152 3161 4158
rect 3149 4144 3161 4152
rect 2758 4098 2770 4104
rect 2808 4098 2820 4104
rect 2859 4098 2871 4104
rect 2990 4098 3002 4104
rect 3090 4098 3102 4104
rect 3216 4124 3224 4179
rect 3276 4171 3284 4199
rect 3357 4183 3363 4233
rect 3375 4213 3382 4268
rect 3475 4213 3482 4268
rect 3575 4213 3582 4268
rect 3718 4213 3725 4268
rect 3757 4242 3769 4244
rect 3757 4236 3797 4242
rect 3957 4316 3969 4322
rect 4037 4316 4049 4322
rect 4151 4316 4163 4322
rect 4191 4316 4203 4322
rect 3818 4201 3826 4236
rect 3893 4201 3901 4236
rect 3327 4177 3363 4183
rect 3376 4171 3384 4199
rect 3476 4171 3484 4199
rect 3576 4171 3584 4199
rect 3716 4171 3724 4199
rect 3276 4162 3306 4171
rect 3276 4160 3294 4162
rect 3376 4162 3406 4171
rect 3376 4160 3394 4162
rect 3476 4162 3506 4171
rect 3476 4160 3494 4162
rect 3576 4162 3606 4171
rect 3576 4160 3594 4162
rect 3119 4098 3131 4104
rect 3231 4098 3243 4104
rect 3330 4098 3342 4104
rect 3430 4098 3442 4104
rect 3530 4098 3542 4104
rect 3630 4098 3642 4104
rect 3694 4162 3724 4171
rect 3706 4160 3724 4162
rect 3818 4144 3826 4187
rect 3976 4193 3984 4276
rect 4017 4242 4029 4244
rect 4017 4236 4057 4242
rect 4135 4274 4143 4276
rect 4217 4316 4229 4322
rect 4257 4316 4269 4322
rect 4337 4316 4349 4322
rect 4422 4316 4434 4322
rect 4472 4316 4484 4322
rect 4537 4316 4549 4322
rect 4691 4316 4703 4322
rect 4171 4274 4182 4276
rect 4135 4268 4182 4274
rect 4238 4274 4249 4276
rect 4277 4274 4285 4276
rect 4238 4268 4285 4274
rect 4078 4201 4086 4236
rect 4135 4213 4142 4268
rect 3899 4165 3907 4187
rect 3900 4158 3925 4165
rect 3800 4133 3826 4144
rect 3857 4144 3909 4147
rect 3869 4138 3897 4144
rect 3917 4144 3925 4158
rect 3976 4124 3984 4179
rect 4278 4213 4285 4268
rect 4317 4242 4329 4244
rect 4317 4236 4357 4242
rect 4529 4238 4557 4244
rect 4569 4310 4597 4316
rect 4378 4201 4386 4236
rect 4453 4201 4461 4236
rect 4576 4230 4588 4236
rect 4561 4224 4588 4230
rect 4663 4229 4680 4236
rect 4561 4201 4567 4224
rect 4078 4144 4086 4187
rect 4136 4171 4144 4199
rect 4276 4171 4284 4199
rect 4136 4162 4166 4171
rect 4136 4160 4154 4162
rect 4060 4133 4086 4144
rect 3658 4098 3670 4104
rect 3760 4098 3772 4104
rect 3810 4098 3822 4104
rect 3877 4098 3889 4104
rect 3957 4098 3969 4104
rect 4020 4098 4032 4104
rect 4070 4098 4082 4104
rect 4190 4098 4202 4104
rect 4254 4162 4284 4171
rect 4266 4160 4284 4162
rect 4378 4144 4386 4187
rect 4459 4165 4467 4187
rect 4460 4158 4485 4165
rect 4360 4133 4386 4144
rect 4417 4144 4469 4147
rect 4429 4138 4457 4144
rect 4477 4144 4485 4158
rect 4553 4144 4560 4187
rect 4673 4181 4680 4229
rect 4673 4124 4680 4167
rect 4218 4098 4230 4104
rect 4320 4098 4332 4104
rect 4370 4098 4382 4104
rect 4437 4098 4449 4104
rect 4520 4098 4532 4104
rect 4576 4098 4588 4104
rect 4651 4098 4663 4104
rect 4691 4098 4703 4104
rect 4782 4098 4842 4562
rect 4 4096 4842 4098
rect 4776 4084 4842 4096
rect 4 4082 4842 4084
rect 69 4076 81 4082
rect 149 4076 161 4082
rect 191 4076 203 4082
rect 231 4076 243 4082
rect 277 4076 289 4082
rect 391 4076 403 4082
rect 451 4076 463 4082
rect 39 4028 51 4036
rect 119 4028 131 4036
rect 39 4022 63 4028
rect 119 4022 143 4028
rect 55 3973 63 4022
rect 135 3973 143 4022
rect 213 4013 220 4056
rect 269 4036 297 4042
rect 257 4033 309 4036
rect 491 4076 503 4082
rect 531 4076 543 4082
rect 587 4076 599 4082
rect 677 4076 689 4082
rect 757 4076 769 4082
rect 837 4076 849 4082
rect 919 4076 931 4082
rect 1031 4076 1043 4082
rect 317 4022 325 4036
rect 300 4015 325 4022
rect 55 3904 63 3959
rect 135 3904 143 3959
rect 213 3951 220 3999
rect 299 3993 307 4015
rect 376 4001 384 4056
rect 436 4001 444 4056
rect 513 4013 520 4056
rect 619 4036 629 4046
rect 557 4026 569 4036
rect 557 4018 595 4026
rect 203 3944 220 3951
rect 293 3944 301 3979
rect 31 3858 43 3864
rect 71 3858 83 3864
rect 111 3858 123 3864
rect 151 3858 163 3864
rect 231 3858 243 3864
rect 376 3904 384 3987
rect 436 3904 444 3987
rect 513 3951 520 3999
rect 503 3944 520 3951
rect 578 3904 586 4018
rect 621 3993 629 4036
rect 669 4036 697 4042
rect 657 4033 709 4036
rect 717 4022 725 4036
rect 700 4015 725 4022
rect 627 3979 629 3993
rect 699 3993 707 4015
rect 776 4001 784 4056
rect 829 4036 857 4042
rect 817 4033 869 4036
rect 1071 4076 1083 4082
rect 1111 4076 1123 4082
rect 1137 4076 1149 4082
rect 1197 4076 1209 4082
rect 1237 4076 1249 4082
rect 1277 4076 1289 4082
rect 1351 4076 1363 4082
rect 1391 4076 1403 4082
rect 1451 4076 1463 4082
rect 1497 4076 1509 4082
rect 1597 4076 1609 4082
rect 1699 4076 1711 4082
rect 1798 4076 1810 4082
rect 1848 4076 1860 4082
rect 877 4022 885 4036
rect 949 4028 961 4036
rect 860 4015 885 4022
rect 937 4022 961 4028
rect 621 3944 629 3979
rect 693 3944 701 3979
rect 262 3858 274 3864
rect 312 3858 324 3864
rect 391 3858 403 3864
rect 451 3858 463 3864
rect 531 3858 543 3864
rect 776 3904 784 3987
rect 859 3993 867 4015
rect 887 3997 903 4003
rect 853 3944 861 3979
rect 897 3947 903 3997
rect 937 3973 945 4022
rect 1016 4001 1024 4056
rect 1093 4013 1100 4056
rect 1156 4001 1164 4056
rect 1220 4013 1227 4056
rect 557 3858 569 3864
rect 601 3858 613 3864
rect 662 3858 674 3864
rect 712 3858 724 3864
rect 937 3904 945 3959
rect 1016 3904 1024 3987
rect 1093 3951 1100 3999
rect 1296 4001 1304 4056
rect 1373 4013 1380 4056
rect 1083 3944 1100 3951
rect 757 3858 769 3864
rect 822 3858 834 3864
rect 872 3858 884 3864
rect 1156 3904 1164 3987
rect 1220 3951 1227 3999
rect 1436 4001 1444 4056
rect 1489 4036 1517 4042
rect 1477 4033 1529 4036
rect 1589 4036 1617 4040
rect 1629 4070 1657 4076
rect 1537 4022 1545 4036
rect 1577 4034 1629 4036
rect 1639 4026 1645 4036
rect 1729 4028 1741 4036
rect 1520 4015 1545 4022
rect 1616 4019 1645 4026
rect 1717 4022 1741 4028
rect 1794 4036 1820 4047
rect 1878 4076 1890 4082
rect 2031 4076 2043 4082
rect 2111 4076 2123 4082
rect 2210 4076 2222 4082
rect 2310 4076 2322 4082
rect 1220 3944 1237 3951
rect 917 3858 929 3864
rect 957 3858 969 3864
rect 1031 3858 1043 3864
rect 1111 3858 1123 3864
rect 1296 3904 1304 3987
rect 1373 3951 1380 3999
rect 1363 3944 1380 3951
rect 1436 3904 1444 3987
rect 1519 3993 1527 4015
rect 1616 3993 1624 4019
rect 1513 3944 1521 3979
rect 1617 3944 1625 3979
rect 1717 3973 1725 4022
rect 1794 3993 1802 4036
rect 1995 4022 2003 4036
rect 2023 4036 2051 4042
rect 2011 4033 2063 4036
rect 1926 4018 1944 4020
rect 1914 4009 1944 4018
rect 1995 4015 2020 4022
rect 1936 3981 1944 4009
rect 2013 3993 2021 4015
rect 2096 4001 2104 4056
rect 2156 4018 2174 4020
rect 1137 3858 1149 3864
rect 1197 3858 1209 3864
rect 1277 3858 1289 3864
rect 1391 3858 1403 3864
rect 1451 3858 1463 3864
rect 1482 3858 1494 3864
rect 1532 3858 1544 3864
rect 1717 3904 1725 3959
rect 1794 3944 1802 3979
rect 2156 4009 2186 4018
rect 2256 4018 2274 4020
rect 2256 4009 2286 4018
rect 2358 4076 2370 4082
rect 2408 4076 2420 4082
rect 2471 4076 2483 4082
rect 2551 4076 2563 4082
rect 2670 4076 2682 4082
rect 2354 4036 2380 4047
rect 1577 3858 1589 3864
rect 1647 3858 1659 3864
rect 1823 3938 1863 3944
rect 1851 3936 1863 3938
rect 1938 3912 1945 3967
rect 2019 3944 2027 3979
rect 1898 3906 1945 3912
rect 1898 3904 1909 3906
rect 1937 3904 1945 3906
rect 2096 3904 2104 3987
rect 2156 3981 2164 4009
rect 2256 3981 2264 4009
rect 2354 3993 2362 4036
rect 2155 3912 2162 3967
rect 2456 4001 2464 4056
rect 2515 4022 2523 4036
rect 2543 4036 2571 4042
rect 2531 4033 2583 4036
rect 2515 4015 2540 4022
rect 2533 3993 2541 4015
rect 2587 4017 2603 4023
rect 2255 3912 2262 3967
rect 2354 3944 2362 3979
rect 2155 3906 2202 3912
rect 2155 3904 2163 3906
rect 2191 3904 2202 3906
rect 2255 3906 2302 3912
rect 2255 3904 2263 3906
rect 2291 3904 2302 3906
rect 2383 3938 2423 3944
rect 2411 3936 2423 3938
rect 2456 3904 2464 3987
rect 2539 3944 2547 3979
rect 2597 3947 2603 4017
rect 2616 4018 2634 4020
rect 2616 4009 2646 4018
rect 2718 4076 2730 4082
rect 2768 4076 2780 4082
rect 2851 4076 2863 4082
rect 2917 4076 2929 4082
rect 3070 4076 3082 4082
rect 3131 4076 3143 4082
rect 3177 4076 3189 4082
rect 3260 4076 3272 4082
rect 3310 4076 3322 4082
rect 3377 4076 3389 4082
rect 3511 4076 3523 4082
rect 3611 4076 3623 4082
rect 3678 4076 3690 4082
rect 3728 4076 3740 4082
rect 3830 4076 3842 4082
rect 3909 4076 3921 4082
rect 3989 4076 4001 4082
rect 2714 4036 2740 4047
rect 2616 3981 2624 4009
rect 1697 3858 1709 3864
rect 1737 3858 1749 3864
rect 1831 3858 1843 3864
rect 1877 3858 1889 3864
rect 1917 3858 1929 3864
rect 1996 3858 2008 3864
rect 2046 3858 2058 3864
rect 2111 3858 2123 3864
rect 2171 3858 2183 3864
rect 2211 3858 2223 3864
rect 2271 3858 2283 3864
rect 2311 3858 2323 3864
rect 2391 3858 2403 3864
rect 2471 3858 2483 3864
rect 2615 3912 2622 3967
rect 2697 3967 2703 4033
rect 2714 3993 2722 4036
rect 2815 4022 2823 4036
rect 2843 4036 2871 4042
rect 2831 4033 2883 4036
rect 2909 4036 2937 4042
rect 2897 4033 2949 4036
rect 2957 4022 2965 4036
rect 2815 4015 2840 4022
rect 2940 4015 2965 4022
rect 3016 4018 3034 4020
rect 2833 3993 2841 4015
rect 2939 3993 2947 4015
rect 3016 4009 3046 4018
rect 3016 3981 3024 4009
rect 3087 3997 3103 4003
rect 3116 4001 3124 4056
rect 3169 4036 3197 4042
rect 3157 4033 3209 4036
rect 3300 4036 3326 4047
rect 3217 4022 3225 4036
rect 3200 4015 3225 4022
rect 2714 3944 2722 3979
rect 2839 3944 2847 3979
rect 2933 3944 2941 3979
rect 2615 3906 2662 3912
rect 2615 3904 2623 3906
rect 2651 3904 2662 3906
rect 2743 3938 2783 3944
rect 2771 3936 2783 3938
rect 2516 3858 2528 3864
rect 2566 3858 2578 3864
rect 2631 3858 2643 3864
rect 2671 3858 2683 3864
rect 2751 3858 2763 3864
rect 2816 3858 2828 3864
rect 2866 3858 2878 3864
rect 3015 3912 3022 3967
rect 3097 3923 3103 3997
rect 3087 3917 3103 3923
rect 3015 3906 3062 3912
rect 3015 3904 3023 3906
rect 3051 3904 3062 3906
rect 3116 3904 3124 3987
rect 3199 3993 3207 4015
rect 3227 3997 3243 4003
rect 3193 3944 3201 3979
rect 3237 3963 3243 3997
rect 3318 3993 3326 4036
rect 3369 4036 3397 4042
rect 3357 4033 3409 4036
rect 3417 4022 3425 4036
rect 3400 4015 3425 4022
rect 3475 4022 3483 4036
rect 3503 4036 3531 4042
rect 3491 4033 3543 4036
rect 3575 4022 3583 4036
rect 3603 4036 3631 4042
rect 3591 4033 3643 4036
rect 3674 4036 3700 4047
rect 3475 4015 3500 4022
rect 3575 4015 3600 4022
rect 3399 3993 3407 4015
rect 3493 3993 3501 4015
rect 3593 3993 3601 4015
rect 3674 3993 3682 4036
rect 3776 4018 3794 4020
rect 3776 4009 3806 4018
rect 4019 4076 4031 4082
rect 4170 4076 4182 4082
rect 4251 4076 4263 4082
rect 4317 4076 4329 4082
rect 4431 4076 4443 4082
rect 4530 4076 4542 4082
rect 4630 4076 4642 4082
rect 3879 4028 3891 4036
rect 3959 4028 3971 4036
rect 4049 4028 4061 4036
rect 3879 4022 3903 4028
rect 3959 4022 3983 4028
rect 3776 3981 3784 4009
rect 3237 3957 3273 3963
rect 3318 3944 3326 3979
rect 3393 3944 3401 3979
rect 3499 3944 3507 3979
rect 3599 3944 3607 3979
rect 3674 3944 3682 3979
rect 2902 3858 2914 3864
rect 2952 3858 2964 3864
rect 3031 3858 3043 3864
rect 3071 3858 3083 3864
rect 3131 3858 3143 3864
rect 3257 3938 3297 3944
rect 3257 3936 3269 3938
rect 3162 3858 3174 3864
rect 3212 3858 3224 3864
rect 3277 3858 3289 3864
rect 3362 3858 3374 3864
rect 3412 3858 3424 3864
rect 3476 3858 3488 3864
rect 3526 3858 3538 3864
rect 3703 3938 3743 3944
rect 3731 3936 3743 3938
rect 3775 3912 3782 3967
rect 3895 3973 3903 4022
rect 3975 3973 3983 4022
rect 4037 4022 4061 4028
rect 4037 3973 4045 4022
rect 4116 4018 4134 4020
rect 4116 4009 4146 4018
rect 4215 4022 4223 4036
rect 4243 4036 4271 4042
rect 4231 4033 4283 4036
rect 4309 4036 4337 4042
rect 4297 4033 4349 4036
rect 4357 4022 4365 4036
rect 4215 4015 4240 4022
rect 4340 4015 4365 4022
rect 4116 3981 4124 4009
rect 4233 3993 4241 4015
rect 4339 3993 4347 4015
rect 4416 4001 4424 4056
rect 4476 4018 4494 4020
rect 4476 4009 4506 4018
rect 4576 4018 4594 4020
rect 4576 4009 4606 4018
rect 4660 4076 4672 4082
rect 4710 4076 4722 4082
rect 4700 4036 4726 4047
rect 3775 3906 3822 3912
rect 3775 3904 3783 3906
rect 3811 3904 3822 3906
rect 3895 3904 3903 3959
rect 3975 3904 3983 3959
rect 4037 3904 4045 3959
rect 4115 3912 4122 3967
rect 4239 3944 4247 3979
rect 4333 3944 4341 3979
rect 4115 3906 4162 3912
rect 4115 3904 4123 3906
rect 3576 3858 3588 3864
rect 3626 3858 3638 3864
rect 3711 3858 3723 3864
rect 3791 3858 3803 3864
rect 3831 3858 3843 3864
rect 3871 3858 3883 3864
rect 3911 3858 3923 3864
rect 3951 3858 3963 3864
rect 3991 3858 4003 3864
rect 4151 3904 4162 3906
rect 4017 3858 4029 3864
rect 4057 3858 4069 3864
rect 4131 3858 4143 3864
rect 4171 3858 4183 3864
rect 4216 3858 4228 3864
rect 4266 3858 4278 3864
rect 4416 3904 4424 3987
rect 4476 3981 4484 4009
rect 4576 3981 4584 4009
rect 4718 3993 4726 4036
rect 4475 3912 4482 3967
rect 4575 3912 4582 3967
rect 4718 3944 4726 3979
rect 4657 3938 4697 3944
rect 4657 3936 4669 3938
rect 4475 3906 4522 3912
rect 4475 3904 4483 3906
rect 4511 3904 4522 3906
rect 4575 3906 4622 3912
rect 4575 3904 4583 3906
rect 4611 3904 4622 3906
rect 4302 3858 4314 3864
rect 4352 3858 4364 3864
rect 4431 3858 4443 3864
rect 4491 3858 4503 3864
rect 4531 3858 4543 3864
rect 4591 3858 4603 3864
rect 4631 3858 4643 3864
rect 4677 3858 4689 3864
rect -62 3856 4776 3858
rect -62 3844 4 3856
rect -62 3842 4776 3844
rect -62 3378 -2 3842
rect 36 3836 48 3842
rect 86 3836 98 3842
rect 151 3836 163 3842
rect 197 3836 209 3842
rect 255 3836 267 3842
rect 301 3836 313 3842
rect 367 3836 379 3842
rect 436 3836 448 3842
rect 486 3836 498 3842
rect 59 3721 67 3756
rect 53 3685 61 3707
rect 136 3713 144 3796
rect 227 3782 239 3816
rect 281 3790 293 3796
rect 335 3790 343 3796
rect 285 3778 307 3790
rect 335 3776 353 3790
rect 233 3758 239 3776
rect 257 3766 287 3772
rect 335 3770 343 3776
rect 35 3678 60 3685
rect 35 3664 43 3678
rect 51 3664 103 3667
rect 63 3658 91 3664
rect 136 3644 144 3699
rect 177 3693 185 3756
rect 199 3744 213 3752
rect 233 3752 273 3758
rect 193 3693 207 3707
rect 177 3679 193 3693
rect 267 3680 273 3752
rect 281 3752 287 3766
rect 305 3762 343 3770
rect 517 3836 529 3842
rect 561 3836 573 3842
rect 661 3836 673 3842
rect 731 3836 743 3842
rect 771 3836 783 3842
rect 821 3836 833 3842
rect 887 3836 899 3842
rect 933 3836 945 3842
rect 991 3836 1003 3842
rect 1069 3836 1081 3842
rect 1137 3836 1149 3842
rect 1195 3836 1207 3842
rect 1241 3836 1253 3842
rect 1307 3836 1319 3842
rect 1362 3836 1374 3842
rect 1412 3836 1424 3842
rect 281 3746 325 3752
rect 337 3748 399 3756
rect 327 3707 354 3714
rect 374 3696 380 3701
rect 346 3688 380 3696
rect 334 3680 341 3688
rect 177 3664 185 3679
rect 267 3674 341 3680
rect 267 3672 273 3674
rect 334 3668 341 3674
rect 227 3650 238 3658
rect 231 3644 238 3650
rect 288 3656 309 3663
rect 393 3664 399 3748
rect 459 3721 467 3756
rect 453 3685 461 3707
rect 435 3678 460 3685
rect 538 3682 546 3796
rect 637 3757 641 3766
rect 581 3721 589 3756
rect 587 3707 589 3721
rect 637 3713 646 3757
rect 695 3748 703 3756
rect 667 3740 703 3748
rect 755 3741 763 3796
rect 857 3790 865 3796
rect 907 3790 919 3796
rect 847 3776 865 3790
rect 893 3778 915 3790
rect 961 3782 973 3816
rect 857 3770 865 3776
rect 857 3762 895 3770
rect 913 3766 943 3772
rect 801 3748 863 3756
rect 435 3664 443 3678
rect 517 3674 555 3682
rect 288 3644 295 3656
rect 353 3644 360 3650
rect 347 3638 360 3644
rect 451 3664 503 3667
rect 463 3658 491 3664
rect 517 3664 529 3674
rect 581 3664 589 3707
rect 633 3664 640 3699
rect 656 3684 662 3739
rect 755 3678 763 3727
rect 667 3672 677 3678
rect 579 3654 589 3664
rect 671 3644 677 3672
rect 739 3672 763 3678
rect 739 3664 751 3672
rect 801 3664 807 3748
rect 913 3752 919 3766
rect 961 3758 967 3776
rect 875 3746 919 3752
rect 927 3752 967 3758
rect 846 3707 873 3714
rect 820 3696 826 3701
rect 820 3688 854 3696
rect 859 3680 866 3688
rect 927 3680 933 3752
rect 987 3744 1001 3752
rect 993 3693 1007 3707
rect 1015 3693 1023 3756
rect 859 3674 933 3680
rect 1007 3679 1023 3693
rect 859 3668 866 3674
rect 927 3672 933 3674
rect 891 3656 912 3663
rect 1015 3664 1023 3679
rect 1051 3721 1059 3756
rect 1095 3750 1103 3796
rect 1077 3744 1103 3750
rect 1167 3782 1179 3816
rect 1221 3790 1233 3796
rect 1275 3790 1283 3796
rect 1225 3778 1247 3790
rect 1275 3776 1293 3790
rect 1173 3758 1179 3776
rect 1197 3766 1227 3772
rect 1275 3770 1283 3776
rect 1077 3738 1080 3744
rect 1051 3707 1053 3721
rect 1051 3664 1059 3707
rect 1073 3682 1080 3738
rect 1077 3676 1080 3682
rect 1117 3693 1125 3756
rect 1139 3744 1153 3752
rect 1173 3752 1213 3758
rect 1133 3693 1147 3707
rect 1117 3679 1133 3693
rect 1207 3680 1213 3752
rect 1221 3752 1227 3766
rect 1245 3762 1283 3770
rect 1457 3836 1469 3842
rect 1497 3836 1509 3842
rect 1537 3836 1549 3842
rect 1577 3836 1589 3842
rect 1639 3836 1651 3842
rect 1717 3836 1729 3842
rect 1775 3836 1787 3842
rect 1821 3836 1833 3842
rect 1887 3836 1899 3842
rect 1971 3836 1983 3842
rect 2051 3836 2063 3842
rect 2131 3836 2143 3842
rect 1221 3746 1265 3752
rect 1277 3748 1339 3756
rect 1267 3707 1294 3714
rect 1314 3696 1320 3701
rect 1286 3688 1320 3696
rect 1274 3680 1281 3688
rect 1077 3670 1099 3676
rect 840 3644 847 3650
rect 905 3644 912 3656
rect 962 3650 973 3658
rect 962 3644 969 3650
rect 840 3638 853 3644
rect 1091 3644 1099 3670
rect 1117 3664 1125 3679
rect 1207 3674 1281 3680
rect 1207 3672 1213 3674
rect 1274 3668 1281 3674
rect 1167 3650 1178 3658
rect 1171 3644 1178 3650
rect 1228 3656 1249 3663
rect 1333 3664 1339 3748
rect 1393 3721 1401 3756
rect 1477 3741 1485 3796
rect 1557 3741 1565 3796
rect 1617 3750 1625 3796
rect 1747 3782 1759 3816
rect 1801 3790 1813 3796
rect 1855 3790 1863 3796
rect 1805 3778 1827 3790
rect 1855 3776 1873 3790
rect 1753 3758 1759 3776
rect 1777 3766 1807 3772
rect 1855 3770 1863 3776
rect 1617 3744 1643 3750
rect 1399 3685 1407 3707
rect 1400 3678 1425 3685
rect 1228 3644 1235 3656
rect 1293 3644 1300 3650
rect 1287 3638 1300 3644
rect 1357 3664 1409 3667
rect 1369 3658 1397 3664
rect 1417 3664 1425 3678
rect 1477 3678 1485 3727
rect 1640 3738 1643 3744
rect 1557 3678 1565 3727
rect 1640 3682 1647 3738
rect 1661 3721 1669 3756
rect 1667 3707 1669 3721
rect 1477 3672 1501 3678
rect 1557 3672 1581 3678
rect 1640 3676 1643 3682
rect 1489 3664 1501 3672
rect 1569 3664 1581 3672
rect 1621 3670 1643 3676
rect 1621 3644 1629 3670
rect 1661 3664 1669 3707
rect 1697 3693 1705 3756
rect 1719 3744 1733 3752
rect 1753 3752 1793 3758
rect 1713 3693 1727 3707
rect 1697 3679 1713 3693
rect 1787 3680 1793 3752
rect 1801 3752 1807 3766
rect 1825 3762 1863 3770
rect 1801 3746 1845 3752
rect 1857 3748 1919 3756
rect 1847 3707 1874 3714
rect 1894 3696 1900 3701
rect 1866 3688 1900 3696
rect 1854 3680 1861 3688
rect 1697 3664 1705 3679
rect 1787 3674 1861 3680
rect 1787 3672 1793 3674
rect 1854 3668 1861 3674
rect 1747 3650 1758 3658
rect 1751 3644 1758 3650
rect 1808 3656 1829 3663
rect 1913 3664 1919 3748
rect 1956 3713 1964 3796
rect 2157 3836 2169 3842
rect 2197 3836 2209 3842
rect 2276 3836 2288 3842
rect 2326 3836 2338 3842
rect 2391 3836 2403 3842
rect 2431 3836 2443 3842
rect 2511 3836 2523 3842
rect 2591 3836 2603 3842
rect 2631 3836 2643 3842
rect 2677 3836 2689 3842
rect 2811 3836 2823 3842
rect 2891 3836 2903 3842
rect 2951 3836 2963 3842
rect 3011 3836 3023 3842
rect 3051 3836 3063 3842
rect 3131 3836 3143 3842
rect 3211 3836 3223 3842
rect 3251 3836 3263 3842
rect 3311 3836 3323 3842
rect 2071 3762 2083 3764
rect 2043 3756 2083 3762
rect 2014 3721 2022 3756
rect 2116 3713 2124 3796
rect 2178 3794 2189 3796
rect 2217 3794 2225 3796
rect 2178 3788 2225 3794
rect 2218 3733 2225 3788
rect 2375 3794 2383 3796
rect 2411 3794 2422 3796
rect 2375 3788 2422 3794
rect 2299 3721 2307 3756
rect 2375 3733 2382 3788
rect 2531 3762 2543 3764
rect 2503 3756 2543 3762
rect 2575 3794 2583 3796
rect 2611 3794 2622 3796
rect 2575 3788 2622 3794
rect 1808 3644 1815 3656
rect 1873 3644 1880 3650
rect 1867 3638 1880 3644
rect 1956 3644 1964 3699
rect 2014 3664 2022 3707
rect 2014 3653 2040 3664
rect 71 3618 83 3624
rect 151 3618 163 3624
rect 199 3618 211 3624
rect 257 3618 269 3624
rect 305 3618 317 3624
rect 367 3618 379 3624
rect 471 3618 483 3624
rect 547 3618 559 3624
rect 651 3618 663 3624
rect 695 3618 703 3624
rect 769 3618 781 3624
rect 821 3618 833 3624
rect 883 3618 895 3624
rect 931 3618 943 3624
rect 989 3618 1001 3624
rect 1069 3618 1081 3624
rect 1139 3618 1151 3624
rect 1197 3618 1209 3624
rect 1245 3618 1257 3624
rect 1307 3618 1319 3624
rect 1377 3618 1389 3624
rect 1459 3618 1471 3624
rect 1539 3618 1551 3624
rect 1639 3618 1651 3624
rect 1719 3618 1731 3624
rect 1777 3618 1789 3624
rect 1825 3618 1837 3624
rect 1887 3618 1899 3624
rect 1971 3618 1983 3624
rect 2116 3644 2124 3699
rect 2216 3691 2224 3719
rect 2018 3618 2030 3624
rect 2068 3618 2080 3624
rect 2131 3618 2143 3624
rect 2194 3682 2224 3691
rect 2293 3685 2301 3707
rect 2474 3721 2482 3756
rect 2575 3733 2582 3788
rect 2657 3762 2669 3764
rect 2657 3756 2697 3762
rect 2831 3762 2843 3764
rect 2803 3756 2843 3762
rect 2376 3691 2384 3719
rect 2206 3680 2224 3682
rect 2275 3678 2300 3685
rect 2376 3682 2406 3691
rect 2376 3680 2394 3682
rect 2275 3664 2283 3678
rect 2291 3664 2343 3667
rect 2303 3658 2331 3664
rect 2474 3664 2482 3707
rect 2557 3687 2563 3733
rect 2718 3721 2726 3756
rect 2774 3721 2782 3756
rect 2576 3691 2584 3719
rect 2576 3682 2606 3691
rect 2576 3680 2594 3682
rect 2474 3653 2500 3664
rect 2158 3618 2170 3624
rect 2311 3618 2323 3624
rect 2430 3618 2442 3624
rect 2718 3664 2726 3707
rect 2478 3618 2490 3624
rect 2528 3618 2540 3624
rect 2630 3618 2642 3624
rect 2700 3653 2726 3664
rect 2774 3664 2782 3707
rect 2857 3667 2863 3733
rect 2876 3713 2884 3796
rect 2936 3713 2944 3796
rect 2995 3794 3003 3796
rect 3031 3794 3042 3796
rect 2995 3788 3042 3794
rect 2995 3733 3002 3788
rect 3151 3762 3163 3764
rect 3123 3756 3163 3762
rect 3195 3794 3203 3796
rect 3356 3836 3368 3842
rect 3406 3836 3418 3842
rect 3231 3794 3242 3796
rect 3195 3788 3242 3794
rect 3094 3721 3102 3756
rect 3195 3733 3202 3788
rect 2774 3653 2800 3664
rect 2660 3618 2672 3624
rect 2710 3618 2722 3624
rect 2876 3644 2884 3699
rect 2936 3644 2944 3699
rect 2996 3691 3004 3719
rect 2996 3682 3026 3691
rect 2996 3680 3014 3682
rect 3094 3664 3102 3707
rect 3196 3691 3204 3719
rect 3296 3713 3304 3796
rect 3451 3836 3463 3842
rect 3491 3836 3503 3842
rect 3517 3836 3529 3842
rect 3561 3836 3573 3842
rect 3671 3836 3683 3842
rect 3751 3836 3763 3842
rect 3791 3836 3803 3842
rect 3851 3836 3863 3842
rect 3897 3836 3909 3842
rect 3996 3836 4008 3842
rect 4046 3836 4058 3842
rect 3379 3721 3387 3756
rect 3475 3741 3483 3796
rect 3196 3682 3226 3691
rect 3196 3680 3214 3682
rect 3094 3653 3120 3664
rect 2778 3618 2790 3624
rect 2828 3618 2840 3624
rect 2891 3618 2903 3624
rect 2951 3618 2963 3624
rect 3050 3618 3062 3624
rect 3296 3644 3304 3699
rect 3373 3685 3381 3707
rect 3355 3678 3380 3685
rect 3475 3678 3483 3727
rect 3538 3682 3546 3796
rect 3691 3762 3703 3764
rect 3663 3756 3703 3762
rect 3735 3794 3743 3796
rect 3771 3794 3782 3796
rect 3735 3788 3782 3794
rect 3581 3721 3589 3756
rect 3634 3721 3642 3756
rect 3735 3733 3742 3788
rect 3807 3777 3823 3783
rect 3587 3707 3589 3721
rect 3355 3664 3363 3678
rect 3459 3672 3483 3678
rect 3517 3674 3555 3682
rect 3371 3664 3423 3667
rect 3383 3658 3411 3664
rect 3459 3664 3471 3672
rect 3517 3664 3529 3674
rect 3581 3664 3589 3707
rect 3579 3654 3589 3664
rect 3634 3664 3642 3707
rect 3736 3691 3744 3719
rect 3736 3682 3766 3691
rect 3736 3680 3754 3682
rect 3634 3653 3660 3664
rect 3817 3667 3823 3777
rect 3836 3713 3844 3796
rect 3877 3762 3889 3764
rect 3877 3756 3917 3762
rect 4082 3836 4094 3842
rect 4132 3836 4144 3842
rect 4197 3836 4209 3842
rect 4331 3836 4343 3842
rect 4377 3836 4389 3842
rect 4417 3836 4429 3842
rect 4511 3836 4523 3842
rect 4571 3836 4583 3842
rect 4611 3836 4623 3842
rect 4177 3762 4189 3764
rect 4177 3756 4217 3762
rect 4398 3794 4409 3796
rect 4437 3794 4445 3796
rect 4398 3788 4445 3794
rect 4351 3762 4363 3764
rect 4323 3756 4363 3762
rect 3938 3721 3946 3756
rect 4019 3721 4027 3756
rect 4113 3721 4121 3756
rect 4238 3721 4246 3756
rect 4294 3721 4302 3756
rect 4438 3733 4445 3788
rect 3836 3644 3844 3699
rect 3938 3664 3946 3707
rect 4013 3685 4021 3707
rect 4119 3685 4127 3707
rect 3995 3678 4020 3685
rect 4120 3678 4145 3685
rect 3995 3664 4003 3678
rect 3098 3618 3110 3624
rect 3148 3618 3160 3624
rect 3250 3618 3262 3624
rect 3311 3618 3323 3624
rect 3391 3618 3403 3624
rect 3489 3618 3501 3624
rect 3547 3618 3559 3624
rect 3638 3618 3650 3624
rect 3688 3618 3700 3624
rect 3790 3618 3802 3624
rect 3851 3618 3863 3624
rect 3920 3653 3946 3664
rect 4011 3664 4063 3667
rect 4023 3658 4051 3664
rect 4077 3664 4129 3667
rect 4089 3658 4117 3664
rect 4137 3664 4145 3678
rect 4238 3664 4246 3707
rect 4220 3653 4246 3664
rect 4294 3664 4302 3707
rect 4436 3691 4444 3719
rect 4496 3713 4504 3796
rect 4555 3794 4563 3796
rect 4637 3836 4649 3842
rect 4677 3836 4689 3842
rect 4591 3794 4602 3796
rect 4555 3788 4602 3794
rect 4658 3794 4669 3796
rect 4697 3794 4705 3796
rect 4658 3788 4705 3794
rect 4555 3733 4562 3788
rect 4698 3733 4705 3788
rect 4294 3653 4320 3664
rect 3880 3618 3892 3624
rect 3930 3618 3942 3624
rect 4031 3618 4043 3624
rect 4097 3618 4109 3624
rect 4180 3618 4192 3624
rect 4230 3618 4242 3624
rect 4298 3618 4310 3624
rect 4348 3618 4360 3624
rect 4414 3682 4444 3691
rect 4426 3680 4444 3682
rect 4496 3644 4504 3699
rect 4556 3691 4564 3719
rect 4696 3691 4704 3719
rect 4556 3682 4586 3691
rect 4556 3680 4574 3682
rect 4378 3618 4390 3624
rect 4511 3618 4523 3624
rect 4610 3618 4622 3624
rect 4674 3682 4704 3691
rect 4686 3680 4704 3682
rect 4638 3618 4650 3624
rect 4782 3618 4842 4082
rect 4 3616 4842 3618
rect 4776 3604 4842 3616
rect 4 3602 4842 3604
rect 41 3596 53 3602
rect 103 3596 115 3602
rect 151 3596 163 3602
rect 209 3596 221 3602
rect 309 3596 321 3602
rect 391 3596 403 3602
rect 489 3596 501 3602
rect 590 3596 602 3602
rect 651 3596 663 3602
rect 731 3596 743 3602
rect 831 3596 843 3602
rect 877 3596 889 3602
rect 951 3596 963 3602
rect 991 3596 1003 3602
rect 1039 3596 1051 3602
rect 1097 3596 1109 3602
rect 1145 3596 1157 3602
rect 1207 3596 1219 3602
rect 1257 3596 1269 3602
rect 1317 3596 1329 3602
rect 1357 3596 1369 3602
rect 1417 3596 1429 3602
rect 1499 3596 1511 3602
rect 1609 3596 1621 3602
rect 1691 3596 1703 3602
rect 1739 3596 1751 3602
rect 1797 3596 1809 3602
rect 1845 3596 1857 3602
rect 1907 3596 1919 3602
rect 1977 3596 1989 3602
rect 2079 3596 2091 3602
rect 2178 3596 2190 3602
rect 2228 3596 2240 3602
rect 2330 3596 2342 3602
rect 2391 3596 2403 3602
rect 2490 3596 2502 3602
rect 2590 3596 2602 3602
rect 2671 3596 2683 3602
rect 2737 3596 2749 3602
rect 2819 3596 2831 3602
rect 2917 3596 2929 3602
rect 2997 3596 3009 3602
rect 3037 3596 3049 3602
rect 3131 3596 3143 3602
rect 3180 3596 3192 3602
rect 3236 3596 3248 3602
rect 60 3576 73 3582
rect 60 3570 67 3576
rect 125 3564 132 3576
rect 21 3472 27 3556
rect 111 3557 132 3564
rect 182 3570 189 3576
rect 182 3562 193 3570
rect 79 3546 86 3552
rect 147 3546 153 3548
rect 79 3540 153 3546
rect 235 3541 243 3556
rect 279 3548 291 3556
rect 279 3542 303 3548
rect 79 3532 86 3540
rect 40 3524 74 3532
rect 40 3519 46 3524
rect 66 3506 93 3513
rect 21 3464 83 3472
rect 95 3468 139 3474
rect 77 3450 115 3458
rect 133 3454 139 3468
rect 147 3468 153 3540
rect 227 3527 243 3541
rect 213 3513 227 3527
rect 147 3462 187 3468
rect 207 3468 221 3476
rect 235 3464 243 3527
rect 295 3493 303 3542
rect 355 3542 363 3556
rect 383 3556 411 3562
rect 371 3553 423 3556
rect 459 3548 471 3556
rect 459 3542 483 3548
rect 355 3535 380 3542
rect 373 3513 381 3535
rect 77 3444 85 3450
rect 133 3448 163 3454
rect 181 3444 187 3462
rect 67 3430 85 3444
rect 113 3430 135 3442
rect 77 3424 85 3430
rect 127 3424 139 3430
rect 181 3404 193 3438
rect 295 3424 303 3479
rect 379 3464 387 3499
rect 475 3493 483 3542
rect 536 3538 554 3540
rect 536 3529 566 3538
rect 536 3501 544 3529
rect 607 3517 623 3523
rect 636 3521 644 3576
rect 695 3542 703 3556
rect 723 3556 751 3562
rect 711 3553 763 3556
rect 795 3542 803 3556
rect 823 3556 851 3562
rect 811 3553 863 3556
rect 695 3535 720 3542
rect 795 3535 820 3542
rect 41 3378 53 3384
rect 107 3378 119 3384
rect 153 3378 165 3384
rect 211 3378 223 3384
rect 271 3378 283 3384
rect 311 3378 323 3384
rect 475 3424 483 3479
rect 535 3432 542 3487
rect 617 3443 623 3517
rect 713 3513 721 3535
rect 607 3437 623 3443
rect 535 3426 582 3432
rect 535 3424 543 3426
rect 356 3378 368 3384
rect 406 3378 418 3384
rect 571 3424 582 3426
rect 636 3424 644 3507
rect 813 3513 821 3535
rect 896 3521 904 3576
rect 973 3533 980 3576
rect 1187 3576 1200 3582
rect 1071 3570 1078 3576
rect 1067 3562 1078 3570
rect 1128 3564 1135 3576
rect 1193 3570 1200 3576
rect 1017 3541 1025 3556
rect 1128 3557 1149 3564
rect 1107 3546 1113 3548
rect 1174 3546 1181 3552
rect 1017 3527 1033 3541
rect 1107 3540 1181 3546
rect 719 3464 727 3499
rect 819 3464 827 3499
rect 451 3378 463 3384
rect 491 3378 503 3384
rect 551 3378 563 3384
rect 591 3378 603 3384
rect 651 3378 663 3384
rect 696 3378 708 3384
rect 746 3378 758 3384
rect 896 3424 904 3507
rect 973 3471 980 3519
rect 963 3464 980 3471
rect 1017 3464 1025 3527
rect 1033 3513 1047 3527
rect 1039 3468 1053 3476
rect 796 3378 808 3384
rect 846 3378 858 3384
rect 1107 3468 1113 3540
rect 1174 3532 1181 3540
rect 1186 3524 1220 3532
rect 1214 3519 1220 3524
rect 1167 3506 1194 3513
rect 1073 3462 1113 3468
rect 1121 3468 1165 3474
rect 1073 3444 1079 3462
rect 1121 3454 1127 3468
rect 1233 3472 1239 3556
rect 1276 3521 1284 3576
rect 1340 3533 1347 3576
rect 1409 3556 1437 3562
rect 1397 3553 1449 3556
rect 1457 3542 1465 3556
rect 1529 3548 1541 3556
rect 1440 3535 1465 3542
rect 1517 3542 1541 3548
rect 1177 3464 1239 3472
rect 1097 3448 1127 3454
rect 1145 3450 1183 3458
rect 1175 3444 1183 3450
rect 1067 3404 1079 3438
rect 1125 3430 1147 3442
rect 1175 3430 1193 3444
rect 1121 3424 1133 3430
rect 1175 3424 1183 3430
rect 1276 3424 1284 3507
rect 1340 3471 1347 3519
rect 1439 3513 1447 3535
rect 1340 3464 1357 3471
rect 1433 3464 1441 3499
rect 1517 3493 1525 3542
rect 1591 3513 1599 3556
rect 1631 3550 1639 3576
rect 1617 3544 1639 3550
rect 1617 3538 1620 3544
rect 1591 3499 1593 3513
rect 1517 3424 1525 3479
rect 1591 3464 1599 3499
rect 1613 3482 1620 3538
rect 1676 3521 1684 3576
rect 1887 3576 1900 3582
rect 1771 3570 1778 3576
rect 1767 3562 1778 3570
rect 1828 3564 1835 3576
rect 1893 3570 1900 3576
rect 1717 3541 1725 3556
rect 1828 3557 1849 3564
rect 1807 3546 1813 3548
rect 1874 3546 1881 3552
rect 1717 3527 1733 3541
rect 1807 3540 1881 3546
rect 1617 3476 1620 3482
rect 1617 3470 1643 3476
rect 877 3378 889 3384
rect 991 3378 1003 3384
rect 1037 3378 1049 3384
rect 1095 3378 1107 3384
rect 1141 3378 1153 3384
rect 1207 3378 1219 3384
rect 1257 3378 1269 3384
rect 1317 3378 1329 3384
rect 1402 3378 1414 3384
rect 1452 3378 1464 3384
rect 1635 3424 1643 3470
rect 1676 3424 1684 3507
rect 1717 3464 1725 3527
rect 1733 3513 1747 3527
rect 1739 3468 1753 3476
rect 1807 3468 1813 3540
rect 1874 3532 1881 3540
rect 1886 3524 1920 3532
rect 1914 3519 1920 3524
rect 1867 3506 1894 3513
rect 1773 3462 1813 3468
rect 1821 3468 1865 3474
rect 1773 3444 1779 3462
rect 1821 3454 1827 3468
rect 1933 3472 1939 3556
rect 1969 3556 1997 3560
rect 2009 3590 2037 3596
rect 1957 3554 2009 3556
rect 2019 3546 2025 3556
rect 2109 3548 2121 3556
rect 1996 3539 2025 3546
rect 2097 3542 2121 3548
rect 2174 3556 2200 3567
rect 1996 3513 2004 3539
rect 1877 3464 1939 3472
rect 1997 3464 2005 3499
rect 2097 3493 2105 3542
rect 2174 3513 2182 3556
rect 2276 3538 2294 3540
rect 2276 3529 2306 3538
rect 2276 3501 2284 3529
rect 2376 3521 2384 3576
rect 2436 3538 2454 3540
rect 2436 3529 2466 3538
rect 2536 3538 2554 3540
rect 2536 3529 2566 3538
rect 2635 3542 2643 3556
rect 2663 3556 2691 3562
rect 2651 3553 2703 3556
rect 2729 3556 2757 3562
rect 2717 3553 2769 3556
rect 2777 3542 2785 3556
rect 2849 3548 2861 3556
rect 2909 3556 2937 3562
rect 2897 3553 2949 3556
rect 2635 3535 2660 3542
rect 2760 3535 2785 3542
rect 2837 3542 2861 3548
rect 2957 3542 2965 3556
rect 1797 3448 1827 3454
rect 1845 3450 1883 3458
rect 1875 3444 1883 3450
rect 1767 3404 1779 3438
rect 1825 3430 1847 3442
rect 1875 3430 1893 3444
rect 1821 3424 1833 3430
rect 1875 3424 1883 3430
rect 2097 3424 2105 3479
rect 2174 3464 2182 3499
rect 1497 3378 1509 3384
rect 1537 3378 1549 3384
rect 1609 3378 1621 3384
rect 1691 3378 1703 3384
rect 1737 3378 1749 3384
rect 1795 3378 1807 3384
rect 1841 3378 1853 3384
rect 1907 3378 1919 3384
rect 1957 3378 1969 3384
rect 2027 3378 2039 3384
rect 2203 3458 2243 3464
rect 2231 3456 2243 3458
rect 2275 3432 2282 3487
rect 2275 3426 2322 3432
rect 2275 3424 2283 3426
rect 2311 3424 2322 3426
rect 2376 3424 2384 3507
rect 2436 3501 2444 3529
rect 2536 3501 2544 3529
rect 2653 3513 2661 3535
rect 2435 3432 2442 3487
rect 2759 3513 2767 3535
rect 2535 3432 2542 3487
rect 2659 3464 2667 3499
rect 2753 3464 2761 3499
rect 2837 3493 2845 3542
rect 2940 3535 2965 3542
rect 2977 3537 2993 3543
rect 2939 3513 2947 3535
rect 2435 3426 2482 3432
rect 2435 3424 2443 3426
rect 2471 3424 2482 3426
rect 2535 3426 2582 3432
rect 2535 3424 2543 3426
rect 2571 3424 2582 3426
rect 2077 3378 2089 3384
rect 2117 3378 2129 3384
rect 2211 3378 2223 3384
rect 2291 3378 2303 3384
rect 2331 3378 2343 3384
rect 2391 3378 2403 3384
rect 2451 3378 2463 3384
rect 2491 3378 2503 3384
rect 2551 3378 2563 3384
rect 2591 3378 2603 3384
rect 2636 3378 2648 3384
rect 2686 3378 2698 3384
rect 2837 3424 2845 3479
rect 2933 3464 2941 3499
rect 2977 3467 2983 3537
rect 3020 3533 3027 3576
rect 3095 3542 3103 3556
rect 3123 3556 3151 3562
rect 3299 3596 3311 3602
rect 3379 3596 3391 3602
rect 3459 3596 3471 3602
rect 3537 3596 3549 3602
rect 3577 3596 3589 3602
rect 3619 3596 3631 3602
rect 3699 3596 3711 3602
rect 3829 3596 3841 3602
rect 3111 3553 3163 3556
rect 3095 3535 3120 3542
rect 3020 3471 3027 3519
rect 3113 3513 3121 3535
rect 3213 3513 3220 3556
rect 3329 3548 3341 3556
rect 3409 3548 3421 3556
rect 3489 3548 3501 3556
rect 3317 3542 3341 3548
rect 3397 3542 3421 3548
rect 3477 3542 3501 3548
rect 2722 3378 2734 3384
rect 2772 3378 2784 3384
rect 2817 3378 2829 3384
rect 2857 3378 2869 3384
rect 3020 3464 3037 3471
rect 3119 3464 3127 3499
rect 3221 3476 3227 3499
rect 3317 3493 3325 3542
rect 3397 3493 3405 3542
rect 3477 3493 3485 3542
rect 3517 3537 3533 3543
rect 3221 3470 3248 3476
rect 3236 3464 3248 3470
rect 2902 3378 2914 3384
rect 2952 3378 2964 3384
rect 3189 3456 3217 3462
rect 3229 3384 3257 3390
rect 3317 3424 3325 3479
rect 3397 3424 3405 3479
rect 3417 3443 3423 3453
rect 3417 3437 3453 3443
rect 3477 3424 3485 3479
rect 3517 3463 3523 3537
rect 3560 3533 3567 3576
rect 3649 3548 3661 3556
rect 3729 3548 3741 3556
rect 3560 3471 3567 3519
rect 3637 3542 3661 3548
rect 3717 3542 3741 3548
rect 3871 3596 3883 3602
rect 3911 3596 3923 3602
rect 3939 3596 3951 3602
rect 4019 3596 4031 3602
rect 4117 3596 4129 3602
rect 4270 3596 4282 3602
rect 3799 3548 3811 3556
rect 3799 3542 3823 3548
rect 3637 3493 3645 3542
rect 3717 3493 3725 3542
rect 3815 3493 3823 3542
rect 3893 3533 3900 3576
rect 3969 3548 3981 3556
rect 4049 3548 4061 3556
rect 4109 3556 4137 3562
rect 4097 3553 4149 3556
rect 3957 3542 3981 3548
rect 4037 3542 4061 3548
rect 4157 3542 4165 3556
rect 3560 3464 3577 3471
rect 3507 3457 3523 3463
rect 2997 3378 3009 3384
rect 3096 3378 3108 3384
rect 3146 3378 3158 3384
rect 3197 3378 3209 3384
rect 3297 3378 3309 3384
rect 3337 3378 3349 3384
rect 3377 3378 3389 3384
rect 3417 3378 3429 3384
rect 3457 3378 3469 3384
rect 3497 3378 3509 3384
rect 3637 3424 3645 3479
rect 3717 3424 3725 3479
rect 3815 3424 3823 3479
rect 3893 3471 3900 3519
rect 3957 3493 3965 3542
rect 4037 3493 4045 3542
rect 4140 3535 4165 3542
rect 4216 3538 4234 3540
rect 4139 3513 4147 3535
rect 4216 3529 4246 3538
rect 4298 3596 4310 3602
rect 4400 3596 4412 3602
rect 4450 3596 4462 3602
rect 4497 3596 4509 3602
rect 4630 3596 4642 3602
rect 4440 3556 4466 3567
rect 4346 3538 4364 3540
rect 4334 3529 4364 3538
rect 4216 3501 4224 3529
rect 4356 3501 4364 3529
rect 4458 3513 4466 3556
rect 4477 3557 4493 3563
rect 3883 3464 3900 3471
rect 3537 3378 3549 3384
rect 3617 3378 3629 3384
rect 3657 3378 3669 3384
rect 3697 3378 3709 3384
rect 3737 3378 3749 3384
rect 3957 3424 3965 3479
rect 4037 3424 4045 3479
rect 4133 3464 4141 3499
rect 3791 3378 3803 3384
rect 3831 3378 3843 3384
rect 3911 3378 3923 3384
rect 3937 3378 3949 3384
rect 3977 3378 3989 3384
rect 4017 3378 4029 3384
rect 4057 3378 4069 3384
rect 4215 3432 4222 3487
rect 4477 3507 4483 3557
rect 4516 3521 4524 3576
rect 4576 3538 4594 3540
rect 4576 3529 4606 3538
rect 4658 3596 4670 3602
rect 4706 3538 4724 3540
rect 4694 3529 4724 3538
rect 4358 3432 4365 3487
rect 4458 3464 4466 3499
rect 4215 3426 4262 3432
rect 4215 3424 4223 3426
rect 4251 3424 4262 3426
rect 4318 3426 4365 3432
rect 4318 3424 4329 3426
rect 4102 3378 4114 3384
rect 4152 3378 4164 3384
rect 4231 3378 4243 3384
rect 4271 3378 4283 3384
rect 4357 3424 4365 3426
rect 4397 3458 4437 3464
rect 4397 3456 4409 3458
rect 4516 3424 4524 3507
rect 4576 3501 4584 3529
rect 4716 3501 4724 3529
rect 4575 3432 4582 3487
rect 4718 3432 4725 3487
rect 4575 3426 4622 3432
rect 4575 3424 4583 3426
rect 4611 3424 4622 3426
rect 4678 3426 4725 3432
rect 4678 3424 4689 3426
rect 4297 3378 4309 3384
rect 4337 3378 4349 3384
rect 4417 3378 4429 3384
rect 4497 3378 4509 3384
rect 4591 3378 4603 3384
rect 4631 3378 4643 3384
rect 4717 3424 4725 3426
rect 4657 3378 4669 3384
rect 4697 3378 4709 3384
rect -62 3376 4776 3378
rect -62 3364 4 3376
rect -62 3362 4776 3364
rect -62 2898 -2 3362
rect 41 3356 53 3362
rect 107 3356 119 3362
rect 153 3356 165 3362
rect 211 3356 223 3362
rect 331 3356 343 3362
rect 377 3356 389 3362
rect 417 3356 429 3362
rect 77 3310 85 3316
rect 127 3310 139 3316
rect 67 3296 85 3310
rect 113 3298 135 3310
rect 181 3302 193 3336
rect 77 3290 85 3296
rect 77 3282 115 3290
rect 133 3286 163 3292
rect 21 3268 83 3276
rect 21 3184 27 3268
rect 133 3272 139 3286
rect 181 3278 187 3296
rect 95 3266 139 3272
rect 147 3272 187 3278
rect 66 3227 93 3234
rect 40 3216 46 3221
rect 40 3208 74 3216
rect 79 3200 86 3208
rect 147 3200 153 3272
rect 283 3350 311 3356
rect 323 3278 351 3284
rect 462 3356 474 3362
rect 512 3356 524 3362
rect 207 3264 221 3272
rect 213 3213 227 3227
rect 235 3213 243 3276
rect 292 3270 304 3276
rect 292 3264 319 3270
rect 313 3241 319 3264
rect 397 3261 405 3316
rect 562 3356 574 3362
rect 612 3356 624 3362
rect 671 3356 683 3362
rect 711 3356 723 3362
rect 737 3356 749 3362
rect 811 3356 823 3362
rect 851 3356 863 3362
rect 891 3356 903 3362
rect 931 3356 943 3362
rect 971 3356 983 3362
rect 79 3194 153 3200
rect 227 3199 243 3213
rect 79 3188 86 3194
rect 147 3192 153 3194
rect 111 3176 132 3183
rect 235 3184 243 3199
rect 320 3184 327 3227
rect 397 3198 405 3247
rect 493 3241 501 3276
rect 593 3241 601 3276
rect 695 3261 703 3316
rect 499 3205 507 3227
rect 599 3205 607 3227
rect 500 3198 525 3205
rect 600 3198 625 3205
rect 695 3198 703 3247
rect 756 3233 764 3316
rect 997 3356 1009 3362
rect 1037 3356 1049 3362
rect 1077 3356 1089 3362
rect 1117 3356 1129 3362
rect 1157 3356 1169 3362
rect 1231 3356 1243 3362
rect 1277 3356 1289 3362
rect 1335 3356 1347 3362
rect 1381 3356 1393 3362
rect 1447 3356 1459 3362
rect 1502 3356 1514 3362
rect 1552 3356 1564 3362
rect 831 3270 843 3276
rect 871 3270 883 3276
rect 911 3270 923 3276
rect 951 3270 963 3276
rect 825 3262 843 3270
rect 858 3262 883 3270
rect 898 3262 923 3270
rect 937 3262 963 3270
rect 1017 3270 1029 3276
rect 1057 3270 1069 3276
rect 1097 3270 1109 3276
rect 1137 3270 1149 3276
rect 1017 3262 1043 3270
rect 1057 3262 1082 3270
rect 1097 3262 1122 3270
rect 1137 3262 1155 3270
rect 825 3233 832 3262
rect 827 3219 832 3233
rect 397 3192 421 3198
rect 409 3184 421 3192
rect 60 3164 67 3170
rect 125 3164 132 3176
rect 182 3170 193 3178
rect 182 3164 189 3170
rect 60 3158 73 3164
rect 41 3138 53 3144
rect 103 3138 115 3144
rect 151 3138 163 3144
rect 209 3138 221 3144
rect 292 3138 304 3144
rect 348 3138 360 3144
rect 457 3184 509 3187
rect 469 3178 497 3184
rect 517 3184 525 3198
rect 557 3184 609 3187
rect 569 3178 597 3184
rect 617 3184 625 3198
rect 679 3192 703 3198
rect 679 3184 691 3192
rect 756 3164 764 3219
rect 825 3198 832 3219
rect 858 3216 866 3262
rect 898 3216 906 3262
rect 937 3216 945 3262
rect 850 3204 866 3216
rect 890 3204 906 3216
rect 930 3204 945 3216
rect 1035 3216 1043 3262
rect 1074 3216 1082 3262
rect 1114 3216 1122 3262
rect 1148 3233 1155 3262
rect 1216 3233 1224 3316
rect 1307 3302 1319 3336
rect 1361 3310 1373 3316
rect 1415 3310 1423 3316
rect 1365 3298 1387 3310
rect 1415 3296 1433 3310
rect 1313 3278 1319 3296
rect 1337 3286 1367 3292
rect 1415 3290 1423 3296
rect 1148 3219 1153 3233
rect 858 3198 866 3204
rect 898 3198 906 3204
rect 937 3198 945 3204
rect 1035 3204 1050 3216
rect 1074 3204 1090 3216
rect 1114 3204 1130 3216
rect 1035 3198 1043 3204
rect 1074 3198 1082 3204
rect 1114 3198 1122 3204
rect 1148 3198 1155 3219
rect 825 3191 844 3198
rect 826 3190 844 3191
rect 858 3190 884 3198
rect 898 3190 923 3198
rect 937 3190 964 3198
rect 832 3184 844 3190
rect 872 3184 884 3190
rect 911 3184 923 3190
rect 952 3184 964 3190
rect 1016 3190 1043 3198
rect 1057 3190 1082 3198
rect 1096 3190 1122 3198
rect 1136 3191 1155 3198
rect 1136 3190 1154 3191
rect 1016 3184 1028 3190
rect 1057 3184 1069 3190
rect 1096 3184 1108 3190
rect 1136 3184 1148 3190
rect 379 3138 391 3144
rect 477 3138 489 3144
rect 577 3138 589 3144
rect 709 3138 721 3144
rect 737 3138 749 3144
rect 811 3138 823 3144
rect 851 3138 863 3144
rect 891 3138 903 3144
rect 931 3138 943 3144
rect 971 3138 983 3144
rect 1216 3164 1224 3219
rect 1257 3213 1265 3276
rect 1279 3264 1293 3272
rect 1313 3272 1353 3278
rect 1273 3213 1287 3227
rect 1257 3199 1273 3213
rect 1347 3200 1353 3272
rect 1361 3272 1367 3286
rect 1385 3282 1423 3290
rect 1616 3356 1628 3362
rect 1666 3356 1678 3362
rect 1716 3356 1728 3362
rect 1766 3356 1778 3362
rect 1831 3356 1843 3362
rect 1876 3356 1888 3362
rect 1926 3356 1938 3362
rect 1361 3266 1405 3272
rect 1417 3268 1479 3276
rect 1407 3227 1434 3234
rect 1454 3216 1460 3221
rect 1426 3208 1460 3216
rect 1414 3200 1421 3208
rect 1257 3184 1265 3199
rect 1347 3194 1421 3200
rect 1347 3192 1353 3194
rect 1414 3188 1421 3194
rect 1307 3170 1318 3178
rect 1311 3164 1318 3170
rect 1368 3176 1389 3183
rect 1473 3184 1479 3268
rect 1533 3241 1541 3276
rect 1639 3241 1647 3276
rect 1739 3241 1747 3276
rect 1539 3205 1547 3227
rect 1633 3205 1641 3227
rect 1733 3205 1741 3227
rect 1816 3233 1824 3316
rect 1976 3356 1988 3362
rect 2026 3356 2038 3362
rect 2077 3356 2089 3362
rect 2135 3356 2147 3362
rect 2181 3356 2193 3362
rect 2247 3356 2259 3362
rect 2331 3356 2343 3362
rect 2391 3356 2403 3362
rect 2451 3356 2463 3362
rect 2491 3356 2503 3362
rect 2537 3356 2549 3362
rect 2651 3356 2663 3362
rect 2107 3302 2119 3336
rect 2161 3310 2173 3316
rect 2215 3310 2223 3316
rect 2165 3298 2187 3310
rect 2215 3296 2233 3310
rect 2113 3278 2119 3296
rect 2137 3286 2167 3292
rect 2215 3290 2223 3296
rect 1899 3241 1907 3276
rect 1999 3241 2007 3276
rect 1540 3198 1565 3205
rect 1368 3164 1375 3176
rect 1433 3164 1440 3170
rect 1427 3158 1440 3164
rect 1497 3184 1549 3187
rect 1509 3178 1537 3184
rect 1557 3184 1565 3198
rect 1615 3198 1640 3205
rect 1715 3198 1740 3205
rect 1615 3184 1623 3198
rect 1631 3184 1683 3187
rect 1715 3184 1723 3198
rect 1643 3178 1671 3184
rect 1731 3184 1783 3187
rect 1743 3178 1771 3184
rect 1816 3164 1824 3219
rect 1893 3205 1901 3227
rect 1993 3205 2001 3227
rect 2057 3213 2065 3276
rect 2079 3264 2093 3272
rect 2113 3272 2153 3278
rect 2073 3213 2087 3227
rect 1875 3198 1900 3205
rect 1975 3198 2000 3205
rect 2057 3199 2073 3213
rect 2147 3200 2153 3272
rect 2161 3272 2167 3286
rect 2185 3282 2223 3290
rect 2161 3266 2205 3272
rect 2217 3268 2279 3276
rect 2207 3227 2234 3234
rect 2254 3216 2260 3221
rect 2226 3208 2260 3216
rect 2214 3200 2221 3208
rect 1875 3184 1883 3198
rect 1891 3184 1943 3187
rect 1975 3184 1983 3198
rect 1903 3178 1931 3184
rect 1991 3184 2043 3187
rect 2003 3178 2031 3184
rect 2057 3184 2065 3199
rect 2147 3194 2221 3200
rect 2147 3192 2153 3194
rect 2214 3188 2221 3194
rect 2107 3170 2118 3178
rect 2111 3164 2118 3170
rect 2168 3176 2189 3183
rect 2273 3184 2279 3268
rect 2316 3233 2324 3316
rect 2376 3233 2384 3316
rect 2435 3314 2443 3316
rect 2471 3314 2482 3316
rect 2435 3308 2482 3314
rect 2435 3253 2442 3308
rect 2517 3282 2529 3284
rect 2517 3276 2557 3282
rect 2696 3356 2708 3362
rect 2746 3356 2758 3362
rect 2578 3241 2586 3276
rect 2168 3164 2175 3176
rect 2233 3164 2240 3170
rect 2227 3158 2240 3164
rect 2316 3164 2324 3219
rect 2376 3164 2384 3219
rect 2436 3211 2444 3239
rect 2436 3202 2466 3211
rect 2636 3233 2644 3316
rect 2777 3356 2789 3362
rect 2862 3356 2874 3362
rect 2912 3356 2924 3362
rect 2957 3356 2969 3362
rect 2997 3356 3009 3362
rect 3037 3356 3049 3362
rect 3077 3356 3089 3362
rect 3171 3356 3183 3362
rect 3251 3356 3263 3362
rect 3291 3356 3303 3362
rect 2937 3277 2953 3283
rect 2719 3241 2727 3276
rect 2800 3269 2817 3276
rect 2436 3200 2454 3202
rect 2578 3184 2586 3227
rect 997 3138 1009 3144
rect 1037 3138 1049 3144
rect 1077 3138 1089 3144
rect 1117 3138 1129 3144
rect 1157 3138 1169 3144
rect 1231 3138 1243 3144
rect 1279 3138 1291 3144
rect 1337 3138 1349 3144
rect 1385 3138 1397 3144
rect 1447 3138 1459 3144
rect 1517 3138 1529 3144
rect 1651 3138 1663 3144
rect 1751 3138 1763 3144
rect 1831 3138 1843 3144
rect 1911 3138 1923 3144
rect 2011 3138 2023 3144
rect 2079 3138 2091 3144
rect 2137 3138 2149 3144
rect 2185 3138 2197 3144
rect 2247 3138 2259 3144
rect 2331 3138 2343 3144
rect 2391 3138 2403 3144
rect 2490 3138 2502 3144
rect 2560 3173 2586 3184
rect 2636 3164 2644 3219
rect 2713 3205 2721 3227
rect 2800 3221 2807 3269
rect 2893 3241 2901 3276
rect 2695 3198 2720 3205
rect 2695 3184 2703 3198
rect 2711 3184 2763 3187
rect 2723 3178 2751 3184
rect 2800 3164 2807 3207
rect 2899 3205 2907 3227
rect 2937 3223 2943 3277
rect 2977 3261 2985 3316
rect 3007 3277 3023 3283
rect 2927 3217 2943 3223
rect 2900 3198 2925 3205
rect 2857 3184 2909 3187
rect 2869 3178 2897 3184
rect 2917 3184 2925 3198
rect 2977 3198 2985 3247
rect 3017 3203 3023 3277
rect 3057 3261 3065 3316
rect 3191 3282 3203 3284
rect 3163 3276 3203 3282
rect 3235 3314 3243 3316
rect 3336 3356 3348 3362
rect 3386 3356 3398 3362
rect 3447 3356 3459 3362
rect 3491 3356 3503 3362
rect 3271 3314 3282 3316
rect 3235 3308 3282 3314
rect 2977 3192 3001 3198
rect 3017 3197 3033 3203
rect 3057 3198 3065 3247
rect 3134 3241 3142 3276
rect 3167 3257 3223 3263
rect 3057 3192 3081 3198
rect 2989 3184 3001 3192
rect 3069 3184 3081 3192
rect 3134 3184 3142 3227
rect 3134 3173 3160 3184
rect 3217 3183 3223 3257
rect 3235 3253 3242 3308
rect 3517 3356 3529 3362
rect 3557 3356 3569 3362
rect 3627 3356 3639 3362
rect 3671 3356 3683 3362
rect 3771 3356 3783 3362
rect 3831 3356 3843 3362
rect 3871 3356 3883 3362
rect 3359 3241 3367 3276
rect 3431 3241 3439 3276
rect 3236 3211 3244 3239
rect 3236 3202 3266 3211
rect 3353 3205 3361 3227
rect 3431 3227 3433 3241
rect 3236 3200 3254 3202
rect 3217 3177 3233 3183
rect 3335 3198 3360 3205
rect 3335 3184 3343 3198
rect 3351 3184 3403 3187
rect 3363 3178 3391 3184
rect 3431 3184 3439 3227
rect 3474 3202 3482 3316
rect 3537 3261 3545 3316
rect 3465 3194 3503 3202
rect 3491 3184 3503 3194
rect 3537 3198 3545 3247
rect 3611 3241 3619 3276
rect 3611 3227 3613 3241
rect 3537 3192 3561 3198
rect 3549 3184 3561 3192
rect 3431 3174 3441 3184
rect 3611 3184 3619 3227
rect 3654 3202 3662 3316
rect 3723 3350 3751 3356
rect 3763 3278 3791 3284
rect 3902 3356 3914 3362
rect 3952 3356 3964 3362
rect 3732 3270 3744 3276
rect 3732 3264 3759 3270
rect 3753 3241 3759 3264
rect 3855 3261 3863 3316
rect 3997 3356 4009 3362
rect 4037 3356 4049 3362
rect 4107 3356 4119 3362
rect 4151 3356 4163 3362
rect 3645 3194 3683 3202
rect 3671 3184 3683 3194
rect 3760 3184 3767 3227
rect 3855 3198 3863 3247
rect 3933 3241 3941 3276
rect 3939 3205 3947 3227
rect 3977 3223 3983 3273
rect 4017 3261 4025 3316
rect 4177 3356 4189 3362
rect 4217 3356 4229 3362
rect 4257 3356 4269 3362
rect 4301 3356 4313 3362
rect 4377 3356 4389 3362
rect 4462 3356 4474 3362
rect 4512 3356 4524 3362
rect 3967 3217 3983 3223
rect 3940 3198 3965 3205
rect 3839 3192 3863 3198
rect 3839 3184 3851 3192
rect 3897 3184 3949 3187
rect 3611 3174 3621 3184
rect 3909 3178 3937 3184
rect 3957 3184 3965 3198
rect 4017 3198 4025 3247
rect 4017 3192 4041 3198
rect 4029 3184 4041 3192
rect 4057 3187 4063 3273
rect 4091 3241 4099 3276
rect 4091 3227 4093 3241
rect 4091 3184 4099 3227
rect 4134 3202 4142 3316
rect 4197 3261 4205 3316
rect 4125 3194 4163 3202
rect 4151 3184 4163 3194
rect 4197 3198 4205 3247
rect 4278 3202 4286 3316
rect 4357 3282 4369 3284
rect 4357 3276 4397 3282
rect 4562 3356 4574 3362
rect 4612 3356 4624 3362
rect 4691 3356 4703 3362
rect 4731 3356 4743 3362
rect 4675 3314 4683 3316
rect 4711 3314 4722 3316
rect 4675 3308 4722 3314
rect 4321 3241 4329 3276
rect 4418 3241 4426 3276
rect 4493 3241 4501 3276
rect 4593 3241 4601 3276
rect 4675 3253 4682 3308
rect 4327 3227 4329 3241
rect 4197 3192 4221 3198
rect 4209 3184 4221 3192
rect 4091 3174 4101 3184
rect 4257 3194 4295 3202
rect 4257 3184 4269 3194
rect 4321 3184 4329 3227
rect 4418 3184 4426 3227
rect 4499 3205 4507 3227
rect 4599 3205 4607 3227
rect 4676 3211 4684 3239
rect 4500 3198 4525 3205
rect 4600 3198 4625 3205
rect 4676 3202 4706 3211
rect 4676 3200 4694 3202
rect 4319 3174 4329 3184
rect 4400 3173 4426 3184
rect 4457 3184 4509 3187
rect 4469 3178 4497 3184
rect 4517 3184 4525 3198
rect 4557 3184 4609 3187
rect 4569 3178 4597 3184
rect 4617 3184 4625 3198
rect 2520 3138 2532 3144
rect 2570 3138 2582 3144
rect 2651 3138 2663 3144
rect 2731 3138 2743 3144
rect 2777 3138 2789 3144
rect 2817 3138 2829 3144
rect 2877 3138 2889 3144
rect 2959 3138 2971 3144
rect 3039 3138 3051 3144
rect 3138 3138 3150 3144
rect 3188 3138 3200 3144
rect 3290 3138 3302 3144
rect 3371 3138 3383 3144
rect 3461 3138 3473 3144
rect 3519 3138 3531 3144
rect 3641 3138 3653 3144
rect 3732 3138 3744 3144
rect 3788 3138 3800 3144
rect 3869 3138 3881 3144
rect 3917 3138 3929 3144
rect 3999 3138 4011 3144
rect 4121 3138 4133 3144
rect 4179 3138 4191 3144
rect 4287 3138 4299 3144
rect 4360 3138 4372 3144
rect 4410 3138 4422 3144
rect 4477 3138 4489 3144
rect 4577 3138 4589 3144
rect 4730 3138 4742 3144
rect 4782 3138 4842 3602
rect 4 3136 4842 3138
rect 4776 3124 4842 3136
rect 4 3122 4842 3124
rect 41 3116 53 3122
rect 103 3116 115 3122
rect 151 3116 163 3122
rect 209 3116 221 3122
rect 311 3116 323 3122
rect 409 3116 421 3122
rect 459 3116 471 3122
rect 517 3116 529 3122
rect 565 3116 577 3122
rect 627 3116 639 3122
rect 701 3116 713 3122
rect 763 3116 775 3122
rect 811 3116 823 3122
rect 869 3116 881 3122
rect 917 3116 929 3122
rect 991 3116 1003 3122
rect 1031 3116 1043 3122
rect 1109 3116 1121 3122
rect 1157 3116 1169 3122
rect 1240 3116 1252 3122
rect 1290 3116 1302 3122
rect 1361 3116 1373 3122
rect 1423 3116 1435 3122
rect 1471 3116 1483 3122
rect 1529 3116 1541 3122
rect 1591 3116 1603 3122
rect 1631 3116 1643 3122
rect 1709 3116 1721 3122
rect 1757 3116 1769 3122
rect 1891 3116 1903 3122
rect 1959 3116 1971 3122
rect 2017 3116 2029 3122
rect 2065 3116 2077 3122
rect 2127 3116 2139 3122
rect 2191 3116 2203 3122
rect 2231 3116 2243 3122
rect 2291 3116 2303 3122
rect 2390 3116 2402 3122
rect 60 3096 73 3102
rect 60 3090 67 3096
rect 125 3084 132 3096
rect 21 2992 27 3076
rect 111 3077 132 3084
rect 182 3090 189 3096
rect 182 3082 193 3090
rect 79 3066 86 3072
rect 147 3066 153 3068
rect 79 3060 153 3066
rect 235 3061 243 3076
rect 79 3052 86 3060
rect 40 3044 74 3052
rect 40 3039 46 3044
rect 66 3026 93 3033
rect 21 2984 83 2992
rect 95 2988 139 2994
rect 77 2970 115 2978
rect 133 2974 139 2988
rect 147 2988 153 3060
rect 227 3047 243 3061
rect 275 3062 283 3076
rect 303 3076 331 3082
rect 291 3073 343 3076
rect 607 3096 620 3102
rect 491 3090 498 3096
rect 487 3082 498 3090
rect 548 3084 555 3096
rect 613 3090 620 3096
rect 379 3068 391 3076
rect 379 3062 403 3068
rect 275 3055 300 3062
rect 213 3033 227 3047
rect 147 2982 187 2988
rect 207 2988 221 2996
rect 235 2984 243 3047
rect 293 3033 301 3055
rect 299 2984 307 3019
rect 395 3013 403 3062
rect 437 3061 445 3076
rect 548 3077 569 3084
rect 527 3066 533 3068
rect 594 3066 601 3072
rect 437 3047 453 3061
rect 527 3060 601 3066
rect 77 2964 85 2970
rect 133 2968 163 2974
rect 181 2964 187 2982
rect 67 2950 85 2964
rect 113 2950 135 2962
rect 77 2944 85 2950
rect 127 2944 139 2950
rect 181 2924 193 2958
rect 395 2944 403 2999
rect 437 2984 445 3047
rect 453 3033 467 3047
rect 459 2988 473 2996
rect 41 2898 53 2904
rect 107 2898 119 2904
rect 153 2898 165 2904
rect 211 2898 223 2904
rect 276 2898 288 2904
rect 326 2898 338 2904
rect 527 2988 533 3060
rect 594 3052 601 3060
rect 606 3044 640 3052
rect 634 3039 640 3044
rect 587 3026 614 3033
rect 493 2982 533 2988
rect 541 2988 585 2994
rect 493 2964 499 2982
rect 541 2974 547 2988
rect 653 2992 659 3076
rect 597 2984 659 2992
rect 517 2968 547 2974
rect 565 2970 603 2978
rect 595 2964 603 2970
rect 487 2924 499 2958
rect 545 2950 567 2962
rect 595 2950 613 2964
rect 541 2944 553 2950
rect 595 2944 603 2950
rect 720 3096 733 3102
rect 720 3090 727 3096
rect 785 3084 792 3096
rect 681 2992 687 3076
rect 771 3077 792 3084
rect 842 3090 849 3096
rect 842 3082 853 3090
rect 739 3066 746 3072
rect 807 3066 813 3068
rect 739 3060 813 3066
rect 895 3061 903 3076
rect 739 3052 746 3060
rect 700 3044 734 3052
rect 700 3039 706 3044
rect 726 3026 753 3033
rect 681 2984 743 2992
rect 755 2988 799 2994
rect 737 2970 775 2978
rect 793 2974 799 2988
rect 807 2988 813 3060
rect 887 3047 903 3061
rect 873 3033 887 3047
rect 807 2982 847 2988
rect 867 2988 881 2996
rect 895 2984 903 3047
rect 936 3041 944 3096
rect 977 3057 993 3063
rect 977 3043 983 3057
rect 1013 3053 1020 3096
rect 1149 3076 1177 3082
rect 1079 3068 1091 3076
rect 1137 3073 1189 3076
rect 1280 3076 1306 3087
rect 1079 3062 1103 3068
rect 1197 3062 1205 3076
rect 957 3037 983 3043
rect 737 2964 745 2970
rect 793 2968 823 2974
rect 841 2964 847 2982
rect 727 2950 745 2964
rect 773 2950 795 2962
rect 737 2944 745 2950
rect 787 2944 799 2950
rect 841 2924 853 2958
rect 936 2944 944 3027
rect 957 2987 963 3037
rect 1013 2991 1020 3039
rect 1095 3013 1103 3062
rect 1180 3055 1205 3062
rect 1179 3033 1187 3055
rect 1298 3033 1306 3076
rect 1380 3096 1393 3102
rect 1380 3090 1387 3096
rect 1445 3084 1452 3096
rect 1003 2984 1020 2991
rect 1095 2944 1103 2999
rect 1173 2984 1181 3019
rect 1298 2984 1306 3019
rect 1341 2992 1347 3076
rect 1431 3077 1452 3084
rect 1502 3090 1509 3096
rect 1502 3082 1513 3090
rect 1399 3066 1406 3072
rect 1467 3066 1473 3068
rect 1399 3060 1473 3066
rect 1555 3061 1563 3076
rect 1399 3052 1406 3060
rect 1360 3044 1394 3052
rect 1360 3039 1366 3044
rect 1386 3026 1413 3033
rect 1341 2984 1403 2992
rect 1415 2988 1459 2994
rect 371 2898 383 2904
rect 411 2898 423 2904
rect 457 2898 469 2904
rect 515 2898 527 2904
rect 561 2898 573 2904
rect 627 2898 639 2904
rect 701 2898 713 2904
rect 767 2898 779 2904
rect 813 2898 825 2904
rect 871 2898 883 2904
rect 917 2898 929 2904
rect 1031 2898 1043 2904
rect 1071 2898 1083 2904
rect 1111 2898 1123 2904
rect 1237 2978 1277 2984
rect 1237 2976 1249 2978
rect 1397 2970 1435 2978
rect 1453 2974 1459 2988
rect 1467 2988 1473 3060
rect 1547 3047 1563 3061
rect 1533 3033 1547 3047
rect 1467 2982 1507 2988
rect 1527 2988 1541 2996
rect 1555 2984 1563 3047
rect 1613 3053 1620 3096
rect 1749 3076 1777 3082
rect 1679 3068 1691 3076
rect 1737 3073 1789 3076
rect 1679 3062 1703 3068
rect 1797 3062 1805 3076
rect 1613 2991 1620 3039
rect 1695 3013 1703 3062
rect 1780 3055 1805 3062
rect 1855 3062 1863 3076
rect 1883 3076 1911 3082
rect 1871 3073 1923 3076
rect 2107 3096 2120 3102
rect 1991 3090 1998 3096
rect 1987 3082 1998 3090
rect 2048 3084 2055 3096
rect 2113 3090 2120 3096
rect 1855 3055 1880 3062
rect 1937 3061 1945 3076
rect 2048 3077 2069 3084
rect 2027 3066 2033 3068
rect 2094 3066 2101 3072
rect 1779 3033 1787 3055
rect 1807 3037 1833 3043
rect 1873 3033 1881 3055
rect 1937 3047 1953 3061
rect 2027 3060 2101 3066
rect 1397 2964 1405 2970
rect 1453 2968 1483 2974
rect 1501 2964 1507 2982
rect 1387 2950 1405 2964
rect 1433 2950 1455 2962
rect 1397 2944 1405 2950
rect 1447 2944 1459 2950
rect 1501 2924 1513 2958
rect 1603 2984 1620 2991
rect 1695 2944 1703 2999
rect 1773 2984 1781 3019
rect 1879 2984 1887 3019
rect 1937 2984 1945 3047
rect 1953 3033 1967 3047
rect 1959 2988 1973 2996
rect 1142 2898 1154 2904
rect 1192 2898 1204 2904
rect 1257 2898 1269 2904
rect 1361 2898 1373 2904
rect 1427 2898 1439 2904
rect 1473 2898 1485 2904
rect 1531 2898 1543 2904
rect 1631 2898 1643 2904
rect 1671 2898 1683 2904
rect 1711 2898 1723 2904
rect 1742 2898 1754 2904
rect 1792 2898 1804 2904
rect 2027 2988 2033 3060
rect 2094 3052 2101 3060
rect 2106 3044 2140 3052
rect 2134 3039 2140 3044
rect 2087 3026 2114 3033
rect 1993 2982 2033 2988
rect 2041 2988 2085 2994
rect 1993 2964 1999 2982
rect 2041 2974 2047 2988
rect 2153 2992 2159 3076
rect 2213 3053 2220 3096
rect 2276 3041 2284 3096
rect 2336 3058 2354 3060
rect 2097 2984 2159 2992
rect 2213 2991 2220 3039
rect 2336 3049 2366 3058
rect 2438 3116 2450 3122
rect 2488 3116 2500 3122
rect 2590 3116 2602 3122
rect 2671 3116 2683 3122
rect 2731 3116 2743 3122
rect 2771 3116 2783 3122
rect 2434 3076 2460 3087
rect 2017 2968 2047 2974
rect 2065 2970 2103 2978
rect 2095 2964 2103 2970
rect 1987 2924 1999 2958
rect 2045 2950 2067 2962
rect 2095 2950 2113 2964
rect 2041 2944 2053 2950
rect 2095 2944 2103 2950
rect 2203 2984 2220 2991
rect 2276 2944 2284 3027
rect 2336 3021 2344 3049
rect 2434 3033 2442 3076
rect 2536 3058 2554 3060
rect 2536 3049 2566 3058
rect 2635 3062 2643 3076
rect 2663 3076 2691 3082
rect 2799 3116 2811 3122
rect 2879 3116 2891 3122
rect 2960 3116 2972 3122
rect 3016 3116 3028 3122
rect 2651 3073 2703 3076
rect 2635 3055 2660 3062
rect 2536 3021 2544 3049
rect 2653 3033 2661 3055
rect 2753 3053 2760 3096
rect 3079 3116 3091 3122
rect 3177 3116 3189 3122
rect 3257 3116 3269 3122
rect 3347 3116 3359 3122
rect 3449 3116 3461 3122
rect 3529 3116 3541 3122
rect 3579 3116 3591 3122
rect 3677 3116 3689 3122
rect 3789 3116 3801 3122
rect 3857 3116 3869 3122
rect 3938 3116 3950 3122
rect 4059 3116 4071 3122
rect 4138 3116 4150 3122
rect 4188 3116 4200 3122
rect 2829 3068 2841 3076
rect 2909 3068 2921 3076
rect 2817 3062 2841 3068
rect 2897 3062 2921 3068
rect 2335 2952 2342 3007
rect 2434 2984 2442 3019
rect 2335 2946 2382 2952
rect 2335 2944 2343 2946
rect 2371 2944 2382 2946
rect 2463 2978 2503 2984
rect 2491 2976 2503 2978
rect 2535 2952 2542 3007
rect 2659 2984 2667 3019
rect 2753 2991 2760 3039
rect 2817 3013 2825 3062
rect 2897 3013 2905 3062
rect 2993 3033 3000 3076
rect 3109 3068 3121 3076
rect 3169 3076 3197 3082
rect 3157 3073 3209 3076
rect 3379 3076 3389 3086
rect 3097 3062 3121 3068
rect 3217 3062 3225 3076
rect 2743 2984 2760 2991
rect 2535 2946 2582 2952
rect 2535 2944 2543 2946
rect 2571 2944 2582 2946
rect 1856 2898 1868 2904
rect 1906 2898 1918 2904
rect 1957 2898 1969 2904
rect 2015 2898 2027 2904
rect 2061 2898 2073 2904
rect 2127 2898 2139 2904
rect 2231 2898 2243 2904
rect 2291 2898 2303 2904
rect 2351 2898 2363 2904
rect 2391 2898 2403 2904
rect 2471 2898 2483 2904
rect 2551 2898 2563 2904
rect 2591 2898 2603 2904
rect 2817 2944 2825 2999
rect 2897 2944 2905 2999
rect 3001 2996 3007 3019
rect 3097 3013 3105 3062
rect 3200 3055 3225 3062
rect 3199 3033 3207 3055
rect 3276 3033 3284 3076
rect 3317 3066 3329 3076
rect 3317 3058 3355 3066
rect 3001 2990 3028 2996
rect 3016 2984 3028 2990
rect 2636 2898 2648 2904
rect 2686 2898 2698 2904
rect 2771 2898 2783 2904
rect 2797 2898 2809 2904
rect 2837 2898 2849 2904
rect 2969 2976 2997 2982
rect 3009 2904 3037 2910
rect 3097 2944 3105 2999
rect 3193 2984 3201 3019
rect 3276 2984 3284 3019
rect 2877 2898 2889 2904
rect 2917 2898 2929 2904
rect 2977 2898 2989 2904
rect 3077 2898 3089 2904
rect 3117 2898 3129 2904
rect 3162 2898 3174 2904
rect 3212 2898 3224 2904
rect 3338 2944 3346 3058
rect 3381 3033 3389 3076
rect 3387 3019 3389 3033
rect 3381 2984 3389 3019
rect 3431 3033 3439 3076
rect 3471 3070 3479 3096
rect 3457 3064 3479 3070
rect 3457 3058 3460 3064
rect 3431 3019 3433 3033
rect 3431 2984 3439 3019
rect 3453 3002 3460 3058
rect 3511 3033 3519 3076
rect 3551 3070 3559 3096
rect 3537 3064 3559 3070
rect 3609 3068 3621 3076
rect 3669 3076 3697 3082
rect 3657 3073 3709 3076
rect 3537 3058 3540 3064
rect 3511 3019 3513 3033
rect 3457 2996 3460 3002
rect 3457 2990 3483 2996
rect 3475 2944 3483 2990
rect 3511 2984 3519 3019
rect 3533 3002 3540 3058
rect 3597 3062 3621 3068
rect 3717 3062 3725 3076
rect 3597 3013 3605 3062
rect 3700 3055 3725 3062
rect 3537 2996 3540 3002
rect 3699 3033 3707 3055
rect 3771 3033 3779 3076
rect 3811 3070 3819 3096
rect 3849 3076 3877 3082
rect 3837 3073 3889 3076
rect 3797 3064 3819 3070
rect 3797 3058 3800 3064
rect 3897 3062 3905 3076
rect 3771 3019 3773 3033
rect 3537 2990 3563 2996
rect 3555 2944 3563 2990
rect 3597 2944 3605 2999
rect 3693 2984 3701 3019
rect 3771 2984 3779 3019
rect 3793 3002 3800 3058
rect 3880 3055 3905 3062
rect 4041 3070 4049 3096
rect 4134 3076 4160 3087
rect 4218 3116 4230 3122
rect 4338 3116 4350 3122
rect 4388 3116 4400 3122
rect 4490 3116 4502 3122
rect 4551 3116 4563 3122
rect 4631 3116 4643 3122
rect 4697 3116 4709 3122
rect 4041 3064 4063 3070
rect 3986 3058 4004 3060
rect 3879 3033 3887 3055
rect 3974 3049 4004 3058
rect 3907 3037 3923 3043
rect 3797 2996 3800 3002
rect 3797 2990 3823 2996
rect 3257 2898 3269 2904
rect 3317 2898 3329 2904
rect 3361 2898 3373 2904
rect 3449 2898 3461 2904
rect 3529 2898 3541 2904
rect 3577 2898 3589 2904
rect 3617 2898 3629 2904
rect 3815 2944 3823 2990
rect 3873 2984 3881 3019
rect 3917 2967 3923 3037
rect 3996 3021 4004 3049
rect 4060 3058 4063 3064
rect 3998 2952 4005 3007
rect 4060 3002 4067 3058
rect 4081 3033 4089 3076
rect 4134 3033 4142 3076
rect 4334 3076 4360 3087
rect 4266 3058 4284 3060
rect 4087 3019 4089 3033
rect 4254 3049 4284 3058
rect 4227 3037 4243 3043
rect 4237 3027 4243 3037
rect 4060 2996 4063 3002
rect 3958 2946 4005 2952
rect 3958 2944 3969 2946
rect 3662 2898 3674 2904
rect 3712 2898 3724 2904
rect 3789 2898 3801 2904
rect 3842 2898 3854 2904
rect 3892 2898 3904 2904
rect 3997 2944 4005 2946
rect 4037 2990 4063 2996
rect 4037 2944 4045 2990
rect 4081 2984 4089 3019
rect 4134 2984 4142 3019
rect 4276 3021 4284 3049
rect 4334 3033 4342 3076
rect 4436 3058 4454 3060
rect 4436 3049 4466 3058
rect 4436 3021 4444 3049
rect 4536 3041 4544 3096
rect 4595 3062 4603 3076
rect 4623 3076 4651 3082
rect 4611 3073 4663 3076
rect 4689 3076 4717 3082
rect 4677 3073 4729 3076
rect 4737 3062 4745 3076
rect 4595 3055 4620 3062
rect 4720 3055 4745 3062
rect 4613 3033 4621 3055
rect 4163 2978 4203 2984
rect 4191 2976 4203 2978
rect 4278 2952 4285 3007
rect 4334 2984 4342 3019
rect 4238 2946 4285 2952
rect 4238 2944 4249 2946
rect 4277 2944 4285 2946
rect 4363 2978 4403 2984
rect 4391 2976 4403 2978
rect 4435 2952 4442 3007
rect 4435 2946 4482 2952
rect 4435 2944 4443 2946
rect 4471 2944 4482 2946
rect 4536 2944 4544 3027
rect 4719 3033 4727 3055
rect 4619 2984 4627 3019
rect 4713 2984 4721 3019
rect 3937 2898 3949 2904
rect 3977 2898 3989 2904
rect 4059 2898 4071 2904
rect 4171 2898 4183 2904
rect 4217 2898 4229 2904
rect 4257 2898 4269 2904
rect 4371 2898 4383 2904
rect 4451 2898 4463 2904
rect 4491 2898 4503 2904
rect 4551 2898 4563 2904
rect 4596 2898 4608 2904
rect 4646 2898 4658 2904
rect 4682 2898 4694 2904
rect 4732 2898 4744 2904
rect -62 2896 4776 2898
rect -62 2884 4 2896
rect -62 2882 4776 2884
rect -62 2418 -2 2882
rect 41 2876 53 2882
rect 107 2876 119 2882
rect 153 2876 165 2882
rect 211 2876 223 2882
rect 331 2876 343 2882
rect 377 2876 389 2882
rect 417 2876 429 2882
rect 77 2830 85 2836
rect 127 2830 139 2836
rect 67 2816 85 2830
rect 113 2818 135 2830
rect 181 2822 193 2856
rect 77 2810 85 2816
rect 77 2802 115 2810
rect 133 2806 163 2812
rect 21 2788 83 2796
rect 21 2704 27 2788
rect 133 2792 139 2806
rect 181 2798 187 2816
rect 95 2786 139 2792
rect 147 2792 187 2798
rect 66 2747 93 2754
rect 40 2736 46 2741
rect 40 2728 74 2736
rect 79 2720 86 2728
rect 147 2720 153 2792
rect 283 2870 311 2876
rect 323 2798 351 2804
rect 476 2876 488 2882
rect 526 2876 538 2882
rect 589 2876 601 2882
rect 637 2876 649 2882
rect 677 2876 689 2882
rect 207 2784 221 2792
rect 213 2733 227 2747
rect 235 2733 243 2796
rect 292 2790 304 2796
rect 292 2784 319 2790
rect 313 2761 319 2784
rect 397 2781 405 2836
rect 736 2876 748 2882
rect 786 2876 798 2882
rect 871 2876 883 2882
rect 79 2714 153 2720
rect 227 2719 243 2733
rect 79 2708 86 2714
rect 147 2712 153 2714
rect 111 2696 132 2703
rect 235 2704 243 2719
rect 320 2704 327 2747
rect 397 2718 405 2767
rect 499 2761 507 2796
rect 571 2761 579 2796
rect 615 2790 623 2836
rect 597 2784 623 2790
rect 597 2778 600 2784
rect 657 2781 665 2836
rect 911 2876 923 2882
rect 951 2876 963 2882
rect 977 2876 989 2882
rect 1051 2876 1063 2882
rect 1091 2876 1103 2882
rect 1117 2876 1129 2882
rect 1229 2876 1241 2882
rect 1301 2876 1313 2882
rect 1367 2876 1379 2882
rect 1413 2876 1425 2882
rect 1471 2876 1483 2882
rect 1517 2876 1529 2882
rect 1557 2876 1569 2882
rect 493 2725 501 2747
rect 571 2747 573 2761
rect 475 2718 500 2725
rect 397 2712 421 2718
rect 409 2704 421 2712
rect 475 2704 483 2718
rect 60 2684 67 2690
rect 125 2684 132 2696
rect 182 2690 193 2698
rect 182 2684 189 2690
rect 60 2678 73 2684
rect 41 2658 53 2664
rect 103 2658 115 2664
rect 151 2658 163 2664
rect 209 2658 221 2664
rect 292 2658 304 2664
rect 348 2658 360 2664
rect 491 2704 543 2707
rect 571 2704 579 2747
rect 593 2722 600 2778
rect 597 2716 600 2722
rect 657 2718 665 2767
rect 759 2761 767 2796
rect 843 2789 860 2796
rect 753 2725 761 2747
rect 853 2741 860 2789
rect 935 2781 943 2836
rect 735 2718 760 2725
rect 597 2710 619 2716
rect 657 2712 681 2718
rect 503 2698 531 2704
rect 611 2684 619 2710
rect 669 2704 681 2712
rect 735 2704 743 2718
rect 751 2704 803 2707
rect 763 2698 791 2704
rect 853 2684 860 2727
rect 935 2718 943 2767
rect 996 2753 1004 2836
rect 1075 2781 1083 2836
rect 1140 2789 1157 2796
rect 919 2712 943 2718
rect 919 2704 931 2712
rect 996 2684 1004 2739
rect 1075 2718 1083 2767
rect 1140 2741 1147 2789
rect 1211 2761 1219 2796
rect 1255 2790 1263 2836
rect 1237 2784 1263 2790
rect 1337 2830 1345 2836
rect 1387 2830 1399 2836
rect 1327 2816 1345 2830
rect 1373 2818 1395 2830
rect 1441 2822 1453 2856
rect 1337 2810 1345 2816
rect 1337 2802 1375 2810
rect 1393 2806 1423 2812
rect 1281 2788 1343 2796
rect 1237 2778 1240 2784
rect 1211 2747 1213 2761
rect 1059 2712 1083 2718
rect 1059 2704 1071 2712
rect 379 2658 391 2664
rect 511 2658 523 2664
rect 589 2658 601 2664
rect 639 2658 651 2664
rect 771 2658 783 2664
rect 831 2658 843 2664
rect 871 2658 883 2664
rect 949 2658 961 2664
rect 1140 2684 1147 2727
rect 1211 2704 1219 2747
rect 1233 2722 1240 2778
rect 1237 2716 1240 2722
rect 1237 2710 1259 2716
rect 977 2658 989 2664
rect 1089 2658 1101 2664
rect 1251 2684 1259 2710
rect 1281 2704 1287 2788
rect 1393 2792 1399 2806
rect 1441 2798 1447 2816
rect 1355 2786 1399 2792
rect 1407 2792 1447 2798
rect 1326 2747 1353 2754
rect 1300 2736 1306 2741
rect 1300 2728 1334 2736
rect 1339 2720 1346 2728
rect 1407 2720 1413 2792
rect 1616 2876 1628 2882
rect 1666 2876 1678 2882
rect 1467 2784 1481 2792
rect 1473 2733 1487 2747
rect 1495 2733 1503 2796
rect 1537 2781 1545 2836
rect 1716 2876 1728 2882
rect 1766 2876 1778 2882
rect 1851 2876 1863 2882
rect 1931 2876 1943 2882
rect 2009 2876 2021 2882
rect 2091 2876 2103 2882
rect 2131 2876 2143 2882
rect 2179 2876 2191 2882
rect 2261 2876 2273 2882
rect 2327 2876 2339 2882
rect 2373 2876 2385 2882
rect 2431 2876 2443 2882
rect 2496 2876 2508 2882
rect 2546 2876 2558 2882
rect 1951 2802 1963 2804
rect 1923 2796 1963 2802
rect 1339 2714 1413 2720
rect 1487 2719 1503 2733
rect 1339 2708 1346 2714
rect 1407 2712 1413 2714
rect 1371 2696 1392 2703
rect 1495 2704 1503 2719
rect 1537 2718 1545 2767
rect 1639 2761 1647 2796
rect 1739 2761 1747 2796
rect 1823 2789 1840 2796
rect 1633 2725 1641 2747
rect 1733 2725 1741 2747
rect 1833 2741 1840 2789
rect 1894 2761 1902 2796
rect 1991 2761 1999 2796
rect 2035 2790 2043 2836
rect 2017 2784 2043 2790
rect 2075 2834 2083 2836
rect 2111 2834 2122 2836
rect 2075 2828 2122 2834
rect 2017 2778 2020 2784
rect 1615 2718 1640 2725
rect 1715 2718 1740 2725
rect 1537 2712 1561 2718
rect 1549 2704 1561 2712
rect 1615 2704 1623 2718
rect 1320 2684 1327 2690
rect 1385 2684 1392 2696
rect 1442 2690 1453 2698
rect 1442 2684 1449 2690
rect 1320 2678 1333 2684
rect 1631 2704 1683 2707
rect 1715 2704 1723 2718
rect 1643 2698 1671 2704
rect 1731 2704 1783 2707
rect 1743 2698 1771 2704
rect 1833 2684 1840 2727
rect 1894 2704 1902 2747
rect 1991 2747 1993 2761
rect 1991 2704 1999 2747
rect 2013 2722 2020 2778
rect 2075 2773 2082 2828
rect 2157 2790 2165 2836
rect 2297 2830 2305 2836
rect 2347 2830 2359 2836
rect 2287 2816 2305 2830
rect 2333 2818 2355 2830
rect 2401 2822 2413 2856
rect 2297 2810 2305 2816
rect 2297 2802 2335 2810
rect 2353 2806 2383 2812
rect 2157 2784 2183 2790
rect 2180 2778 2183 2784
rect 2017 2716 2020 2722
rect 2076 2731 2084 2759
rect 2076 2722 2106 2731
rect 2076 2720 2094 2722
rect 2017 2710 2039 2716
rect 1894 2693 1920 2704
rect 1117 2658 1129 2664
rect 1157 2658 1169 2664
rect 1229 2658 1241 2664
rect 1301 2658 1313 2664
rect 1363 2658 1375 2664
rect 1411 2658 1423 2664
rect 1469 2658 1481 2664
rect 1519 2658 1531 2664
rect 1651 2658 1663 2664
rect 1751 2658 1763 2664
rect 1811 2658 1823 2664
rect 1851 2658 1863 2664
rect 2031 2684 2039 2710
rect 2180 2722 2187 2778
rect 2201 2761 2209 2796
rect 2207 2747 2209 2761
rect 2180 2716 2183 2722
rect 2161 2710 2183 2716
rect 2161 2684 2169 2710
rect 2201 2704 2209 2747
rect 2241 2788 2303 2796
rect 2241 2704 2247 2788
rect 2353 2792 2359 2806
rect 2401 2798 2407 2816
rect 2315 2786 2359 2792
rect 2367 2792 2407 2798
rect 2286 2747 2313 2754
rect 2260 2736 2266 2741
rect 2260 2728 2294 2736
rect 2299 2720 2306 2728
rect 2367 2720 2373 2792
rect 2596 2876 2608 2882
rect 2646 2876 2658 2882
rect 2682 2876 2694 2882
rect 2732 2876 2744 2882
rect 2777 2876 2789 2882
rect 2817 2876 2829 2882
rect 2857 2876 2869 2882
rect 2897 2876 2909 2882
rect 2942 2876 2954 2882
rect 2992 2876 3004 2882
rect 2427 2784 2441 2792
rect 2433 2733 2447 2747
rect 2455 2733 2463 2796
rect 2519 2761 2527 2796
rect 2619 2761 2627 2796
rect 2713 2761 2721 2796
rect 2797 2781 2805 2836
rect 2877 2781 2885 2836
rect 2907 2797 2923 2803
rect 2299 2714 2373 2720
rect 2447 2719 2463 2733
rect 2513 2725 2521 2747
rect 2613 2725 2621 2747
rect 2719 2725 2727 2747
rect 2757 2743 2763 2753
rect 2747 2737 2763 2743
rect 2299 2708 2306 2714
rect 2367 2712 2373 2714
rect 2331 2696 2352 2703
rect 2455 2704 2463 2719
rect 2495 2718 2520 2725
rect 2595 2718 2620 2725
rect 2720 2718 2745 2725
rect 2495 2704 2503 2718
rect 2280 2684 2287 2690
rect 2345 2684 2352 2696
rect 2402 2690 2413 2698
rect 2402 2684 2409 2690
rect 2280 2678 2293 2684
rect 2511 2704 2563 2707
rect 2595 2704 2603 2718
rect 2523 2698 2551 2704
rect 2611 2704 2663 2707
rect 2623 2698 2651 2704
rect 2677 2704 2729 2707
rect 2689 2698 2717 2704
rect 2737 2704 2745 2718
rect 2797 2718 2805 2767
rect 2877 2718 2885 2767
rect 2917 2723 2923 2797
rect 3042 2876 3054 2882
rect 3092 2876 3104 2882
rect 3137 2876 3149 2882
rect 3177 2876 3189 2882
rect 3236 2876 3248 2882
rect 3286 2876 3298 2882
rect 2973 2761 2981 2796
rect 3073 2761 3081 2796
rect 3157 2781 3165 2836
rect 3331 2876 3343 2882
rect 3371 2876 3383 2882
rect 3397 2876 3409 2882
rect 3437 2876 3449 2882
rect 3516 2876 3528 2882
rect 3566 2876 3578 2882
rect 2797 2712 2821 2718
rect 2877 2712 2901 2718
rect 2917 2717 2933 2723
rect 2979 2725 2987 2747
rect 3079 2725 3087 2747
rect 2980 2718 3005 2725
rect 3080 2718 3105 2725
rect 2809 2704 2821 2712
rect 2889 2704 2901 2712
rect 2937 2704 2989 2707
rect 2949 2698 2977 2704
rect 2997 2704 3005 2718
rect 3037 2704 3089 2707
rect 3049 2698 3077 2704
rect 3097 2704 3105 2718
rect 3157 2718 3165 2767
rect 3259 2761 3267 2796
rect 3355 2781 3363 2836
rect 3418 2834 3429 2836
rect 3457 2834 3465 2836
rect 3418 2828 3465 2834
rect 3253 2725 3261 2747
rect 3235 2718 3260 2725
rect 3355 2718 3363 2767
rect 3458 2773 3465 2828
rect 3456 2731 3464 2759
rect 3497 2743 3503 2813
rect 3602 2876 3614 2882
rect 3652 2876 3664 2882
rect 3711 2876 3723 2882
rect 3751 2876 3763 2882
rect 3796 2876 3808 2882
rect 3846 2876 3858 2882
rect 3697 2797 3713 2803
rect 3539 2761 3547 2796
rect 3633 2761 3641 2796
rect 3497 2737 3513 2743
rect 3157 2712 3181 2718
rect 3169 2704 3181 2712
rect 3235 2704 3243 2718
rect 3339 2712 3363 2718
rect 3251 2704 3303 2707
rect 3263 2698 3291 2704
rect 3339 2704 3351 2712
rect 1898 2658 1910 2664
rect 1948 2658 1960 2664
rect 2009 2658 2021 2664
rect 2130 2658 2142 2664
rect 2179 2658 2191 2664
rect 2261 2658 2273 2664
rect 2323 2658 2335 2664
rect 2371 2658 2383 2664
rect 2429 2658 2441 2664
rect 2531 2658 2543 2664
rect 2631 2658 2643 2664
rect 2697 2658 2709 2664
rect 2779 2658 2791 2664
rect 2859 2658 2871 2664
rect 2957 2658 2969 2664
rect 3057 2658 3069 2664
rect 3139 2658 3151 2664
rect 3271 2658 3283 2664
rect 3369 2658 3381 2664
rect 3434 2722 3464 2731
rect 3533 2725 3541 2747
rect 3639 2725 3647 2747
rect 3446 2720 3464 2722
rect 3515 2718 3540 2725
rect 3640 2718 3665 2725
rect 3515 2704 3523 2718
rect 3531 2704 3583 2707
rect 3543 2698 3571 2704
rect 3597 2704 3649 2707
rect 3609 2698 3637 2704
rect 3657 2704 3665 2718
rect 3697 2723 3703 2797
rect 3735 2781 3743 2836
rect 3767 2797 3783 2803
rect 3687 2717 3703 2723
rect 3735 2718 3743 2767
rect 3719 2712 3743 2718
rect 3777 2723 3783 2797
rect 3877 2876 3889 2882
rect 3917 2876 3929 2882
rect 3977 2876 3989 2882
rect 4111 2876 4123 2882
rect 4157 2876 4169 2882
rect 4197 2876 4209 2882
rect 4262 2876 4274 2882
rect 4312 2876 4324 2882
rect 3898 2834 3909 2836
rect 3937 2834 3945 2836
rect 3898 2828 3945 2834
rect 3819 2761 3827 2796
rect 3938 2773 3945 2828
rect 3813 2725 3821 2747
rect 3936 2731 3944 2759
rect 3996 2753 4004 2836
rect 4063 2870 4091 2876
rect 4103 2798 4131 2804
rect 4178 2834 4189 2836
rect 4217 2834 4225 2836
rect 4178 2828 4225 2834
rect 4072 2790 4084 2796
rect 4072 2784 4099 2790
rect 3767 2717 3783 2723
rect 3795 2718 3820 2725
rect 3719 2704 3731 2712
rect 3795 2704 3803 2718
rect 3811 2704 3863 2707
rect 3823 2698 3851 2704
rect 3914 2722 3944 2731
rect 3926 2720 3944 2722
rect 3996 2684 4004 2739
rect 4037 2723 4043 2773
rect 4093 2761 4099 2784
rect 4218 2773 4225 2828
rect 4357 2876 4369 2882
rect 4401 2876 4413 2882
rect 4477 2876 4489 2882
rect 4577 2876 4589 2882
rect 4657 2876 4669 2882
rect 4037 2717 4053 2723
rect 4100 2704 4107 2747
rect 4216 2731 4224 2759
rect 4293 2761 4301 2796
rect 3398 2658 3410 2664
rect 3551 2658 3563 2664
rect 3617 2658 3629 2664
rect 3749 2658 3761 2664
rect 3831 2658 3843 2664
rect 3878 2658 3890 2664
rect 3977 2658 3989 2664
rect 4072 2658 4084 2664
rect 4128 2658 4140 2664
rect 4194 2722 4224 2731
rect 4206 2720 4224 2722
rect 4237 2723 4243 2753
rect 4237 2717 4253 2723
rect 4299 2725 4307 2747
rect 4300 2718 4325 2725
rect 4378 2722 4386 2836
rect 4469 2798 4497 2804
rect 4509 2870 4537 2876
rect 4421 2761 4429 2796
rect 4516 2790 4528 2796
rect 4501 2784 4528 2790
rect 4501 2761 4507 2784
rect 4427 2747 4429 2761
rect 4257 2704 4309 2707
rect 4269 2698 4297 2704
rect 4317 2704 4325 2718
rect 4357 2714 4395 2722
rect 4357 2704 4369 2714
rect 4421 2704 4429 2747
rect 4493 2704 4500 2747
rect 4596 2753 4604 2836
rect 4637 2802 4649 2804
rect 4637 2796 4677 2802
rect 4698 2761 4706 2796
rect 4419 2694 4429 2704
rect 4596 2684 4604 2739
rect 4698 2704 4706 2747
rect 4158 2658 4170 2664
rect 4277 2658 4289 2664
rect 4387 2658 4399 2664
rect 4460 2658 4472 2664
rect 4516 2658 4528 2664
rect 4680 2693 4706 2704
rect 4757 2703 4763 2773
rect 4727 2697 4763 2703
rect 4577 2658 4589 2664
rect 4640 2658 4652 2664
rect 4690 2658 4702 2664
rect 4782 2658 4842 3122
rect 4 2656 4842 2658
rect 4776 2644 4842 2656
rect 4 2642 4842 2644
rect 41 2636 53 2642
rect 103 2636 115 2642
rect 151 2636 163 2642
rect 209 2636 221 2642
rect 311 2636 323 2642
rect 379 2636 391 2642
rect 439 2636 451 2642
rect 571 2636 583 2642
rect 639 2636 651 2642
rect 751 2636 763 2642
rect 797 2636 809 2642
rect 837 2636 849 2642
rect 901 2636 913 2642
rect 963 2636 975 2642
rect 1011 2636 1023 2642
rect 1069 2636 1081 2642
rect 1117 2636 1129 2642
rect 1197 2636 1209 2642
rect 1277 2636 1289 2642
rect 1339 2636 1351 2642
rect 1439 2636 1451 2642
rect 1497 2636 1509 2642
rect 1545 2636 1557 2642
rect 1607 2636 1619 2642
rect 1677 2636 1689 2642
rect 1779 2636 1791 2642
rect 1837 2636 1849 2642
rect 1885 2636 1897 2642
rect 1947 2636 1959 2642
rect 1997 2636 2009 2642
rect 2037 2636 2049 2642
rect 2077 2636 2089 2642
rect 2117 2636 2129 2642
rect 2157 2636 2169 2642
rect 2221 2636 2233 2642
rect 2283 2636 2295 2642
rect 2331 2636 2343 2642
rect 2389 2636 2401 2642
rect 2489 2636 2501 2642
rect 60 2616 73 2622
rect 60 2610 67 2616
rect 125 2604 132 2616
rect 21 2512 27 2596
rect 111 2597 132 2604
rect 182 2610 189 2616
rect 182 2602 193 2610
rect 79 2586 86 2592
rect 147 2586 153 2588
rect 79 2580 153 2586
rect 235 2581 243 2596
rect 79 2572 86 2580
rect 40 2564 74 2572
rect 40 2559 46 2564
rect 66 2546 93 2553
rect 21 2504 83 2512
rect 95 2508 139 2514
rect 77 2490 115 2498
rect 133 2494 139 2508
rect 147 2508 153 2580
rect 227 2567 243 2581
rect 275 2582 283 2596
rect 303 2596 331 2602
rect 291 2593 343 2596
rect 361 2590 369 2616
rect 361 2584 383 2590
rect 275 2575 300 2582
rect 380 2578 383 2584
rect 213 2553 227 2567
rect 147 2502 187 2508
rect 207 2508 221 2516
rect 235 2504 243 2567
rect 293 2553 301 2575
rect 299 2504 307 2539
rect 380 2522 387 2578
rect 401 2553 409 2596
rect 469 2588 481 2596
rect 457 2582 481 2588
rect 535 2582 543 2596
rect 563 2596 591 2602
rect 551 2593 603 2596
rect 621 2590 629 2616
rect 621 2584 643 2590
rect 407 2539 409 2553
rect 380 2516 383 2522
rect 357 2510 383 2516
rect 77 2484 85 2490
rect 133 2488 163 2494
rect 181 2484 187 2502
rect 67 2470 85 2484
rect 113 2470 135 2482
rect 77 2464 85 2470
rect 127 2464 139 2470
rect 181 2444 193 2478
rect 357 2464 365 2510
rect 401 2504 409 2539
rect 457 2533 465 2582
rect 535 2575 560 2582
rect 640 2578 643 2584
rect 553 2553 561 2575
rect 457 2464 465 2519
rect 559 2504 567 2539
rect 640 2522 647 2578
rect 661 2553 669 2596
rect 715 2582 723 2596
rect 743 2596 771 2602
rect 731 2593 783 2596
rect 715 2575 740 2582
rect 667 2539 669 2553
rect 733 2553 741 2575
rect 820 2573 827 2616
rect 640 2516 643 2522
rect 617 2510 643 2516
rect 41 2418 53 2424
rect 107 2418 119 2424
rect 153 2418 165 2424
rect 211 2418 223 2424
rect 276 2418 288 2424
rect 326 2418 338 2424
rect 379 2418 391 2424
rect 437 2418 449 2424
rect 477 2418 489 2424
rect 617 2464 625 2510
rect 661 2504 669 2539
rect 739 2504 747 2539
rect 820 2511 827 2559
rect 920 2616 933 2622
rect 920 2610 927 2616
rect 985 2604 992 2616
rect 881 2512 887 2596
rect 971 2597 992 2604
rect 1042 2610 1049 2616
rect 1042 2602 1053 2610
rect 939 2586 946 2592
rect 1007 2586 1013 2588
rect 939 2580 1013 2586
rect 1095 2581 1103 2596
rect 939 2572 946 2580
rect 900 2564 934 2572
rect 900 2559 906 2564
rect 926 2546 953 2553
rect 820 2504 837 2511
rect 536 2418 548 2424
rect 586 2418 598 2424
rect 639 2418 651 2424
rect 716 2418 728 2424
rect 766 2418 778 2424
rect 881 2504 943 2512
rect 955 2508 999 2514
rect 937 2490 975 2498
rect 993 2494 999 2508
rect 1007 2508 1013 2580
rect 1087 2567 1103 2581
rect 1073 2553 1087 2567
rect 1007 2502 1047 2508
rect 1067 2508 1081 2516
rect 1095 2504 1103 2567
rect 1136 2561 1144 2616
rect 1189 2596 1217 2602
rect 1177 2593 1229 2596
rect 1237 2582 1245 2596
rect 1220 2575 1245 2582
rect 937 2484 945 2490
rect 993 2488 1023 2494
rect 1041 2484 1047 2502
rect 927 2470 945 2484
rect 973 2470 995 2482
rect 937 2464 945 2470
rect 987 2464 999 2470
rect 1041 2444 1053 2478
rect 1136 2464 1144 2547
rect 1219 2553 1227 2575
rect 1296 2561 1304 2616
rect 1369 2588 1381 2596
rect 1357 2582 1381 2588
rect 1587 2616 1600 2622
rect 1471 2610 1478 2616
rect 1467 2602 1478 2610
rect 1528 2604 1535 2616
rect 1593 2610 1600 2616
rect 1213 2504 1221 2539
rect 1296 2464 1304 2547
rect 1357 2533 1365 2582
rect 1417 2581 1425 2596
rect 1528 2597 1549 2604
rect 1507 2586 1513 2588
rect 1574 2586 1581 2592
rect 1417 2567 1433 2581
rect 1507 2580 1581 2586
rect 1357 2464 1365 2519
rect 1417 2504 1425 2567
rect 1433 2553 1447 2567
rect 1439 2508 1453 2516
rect 797 2418 809 2424
rect 901 2418 913 2424
rect 967 2418 979 2424
rect 1013 2418 1025 2424
rect 1071 2418 1083 2424
rect 1117 2418 1129 2424
rect 1182 2418 1194 2424
rect 1232 2418 1244 2424
rect 1507 2508 1513 2580
rect 1574 2572 1581 2580
rect 1586 2564 1620 2572
rect 1614 2559 1620 2564
rect 1567 2546 1594 2553
rect 1473 2502 1513 2508
rect 1521 2508 1565 2514
rect 1473 2484 1479 2502
rect 1521 2494 1527 2508
rect 1633 2512 1639 2596
rect 1669 2596 1697 2602
rect 1657 2593 1709 2596
rect 1927 2616 1940 2622
rect 1811 2610 1818 2616
rect 1807 2602 1818 2610
rect 1868 2604 1875 2616
rect 1933 2610 1940 2616
rect 1717 2582 1725 2596
rect 1700 2575 1725 2582
rect 1757 2581 1765 2596
rect 1868 2597 1889 2604
rect 2240 2616 2253 2622
rect 2240 2610 2247 2616
rect 2305 2604 2312 2616
rect 1847 2586 1853 2588
rect 1914 2586 1921 2592
rect 1699 2553 1707 2575
rect 1757 2567 1773 2581
rect 1847 2580 1921 2586
rect 1577 2504 1639 2512
rect 1693 2504 1701 2539
rect 1757 2504 1765 2567
rect 1773 2553 1787 2567
rect 1779 2508 1793 2516
rect 1497 2488 1527 2494
rect 1545 2490 1583 2498
rect 1575 2484 1583 2490
rect 1467 2444 1479 2478
rect 1525 2470 1547 2482
rect 1575 2470 1593 2484
rect 1521 2464 1533 2470
rect 1575 2464 1583 2470
rect 1847 2508 1853 2580
rect 1914 2572 1921 2580
rect 1926 2564 1960 2572
rect 1954 2559 1960 2564
rect 1907 2546 1934 2553
rect 1813 2502 1853 2508
rect 1861 2508 1905 2514
rect 1813 2484 1819 2502
rect 1861 2494 1867 2508
rect 1973 2512 1979 2596
rect 2016 2590 2028 2596
rect 2057 2590 2069 2596
rect 2096 2590 2108 2596
rect 2136 2590 2148 2596
rect 2016 2582 2043 2590
rect 2057 2582 2082 2590
rect 2096 2582 2122 2590
rect 2136 2589 2154 2590
rect 2136 2582 2155 2589
rect 2035 2576 2043 2582
rect 2074 2576 2082 2582
rect 2114 2576 2122 2582
rect 2035 2564 2050 2576
rect 2074 2564 2090 2576
rect 2114 2564 2130 2576
rect 2035 2518 2043 2564
rect 2074 2518 2082 2564
rect 2114 2518 2122 2564
rect 2148 2561 2155 2582
rect 2148 2547 2153 2561
rect 2148 2518 2155 2547
rect 1917 2504 1979 2512
rect 2017 2510 2043 2518
rect 2057 2510 2082 2518
rect 2097 2510 2122 2518
rect 2137 2510 2155 2518
rect 2201 2512 2207 2596
rect 2291 2597 2312 2604
rect 2362 2610 2369 2616
rect 2362 2602 2373 2610
rect 2259 2586 2266 2592
rect 2327 2586 2333 2588
rect 2259 2580 2333 2586
rect 2415 2581 2423 2596
rect 2517 2636 2529 2642
rect 2631 2636 2643 2642
rect 2677 2636 2689 2642
rect 2789 2636 2801 2642
rect 2871 2636 2883 2642
rect 2947 2636 2959 2642
rect 3037 2636 3049 2642
rect 3169 2636 3181 2642
rect 3227 2636 3239 2642
rect 3370 2636 3382 2642
rect 2459 2588 2471 2596
rect 2459 2582 2483 2588
rect 2259 2572 2266 2580
rect 2220 2564 2254 2572
rect 2220 2559 2226 2564
rect 2246 2546 2273 2553
rect 2017 2504 2029 2510
rect 2057 2504 2069 2510
rect 2097 2504 2109 2510
rect 2137 2504 2149 2510
rect 2201 2504 2263 2512
rect 2275 2508 2319 2514
rect 1837 2488 1867 2494
rect 1885 2490 1923 2498
rect 1915 2484 1923 2490
rect 1807 2444 1819 2478
rect 1865 2470 1887 2482
rect 1915 2470 1933 2484
rect 1861 2464 1873 2470
rect 1915 2464 1923 2470
rect 2257 2490 2295 2498
rect 2313 2494 2319 2508
rect 2327 2508 2333 2580
rect 2407 2567 2423 2581
rect 2393 2553 2407 2567
rect 2327 2502 2367 2508
rect 2387 2508 2401 2516
rect 2415 2504 2423 2567
rect 2475 2533 2483 2582
rect 2536 2561 2544 2616
rect 2595 2582 2603 2596
rect 2623 2596 2651 2602
rect 2611 2593 2663 2596
rect 2595 2575 2620 2582
rect 2613 2553 2621 2575
rect 2257 2484 2265 2490
rect 2313 2488 2343 2494
rect 2361 2484 2367 2502
rect 2247 2470 2265 2484
rect 2293 2470 2315 2482
rect 2257 2464 2265 2470
rect 2307 2464 2319 2470
rect 2361 2444 2373 2478
rect 2475 2464 2483 2519
rect 2536 2464 2544 2547
rect 2696 2561 2704 2616
rect 2759 2588 2771 2596
rect 2759 2582 2783 2588
rect 2619 2504 2627 2539
rect 1277 2418 1289 2424
rect 1337 2418 1349 2424
rect 1377 2418 1389 2424
rect 1437 2418 1449 2424
rect 1495 2418 1507 2424
rect 1541 2418 1553 2424
rect 1607 2418 1619 2424
rect 1662 2418 1674 2424
rect 1712 2418 1724 2424
rect 1777 2418 1789 2424
rect 1835 2418 1847 2424
rect 1881 2418 1893 2424
rect 1947 2418 1959 2424
rect 1997 2418 2009 2424
rect 2037 2418 2049 2424
rect 2077 2418 2089 2424
rect 2117 2418 2129 2424
rect 2157 2418 2169 2424
rect 2221 2418 2233 2424
rect 2287 2418 2299 2424
rect 2333 2418 2345 2424
rect 2391 2418 2403 2424
rect 2451 2418 2463 2424
rect 2491 2418 2503 2424
rect 2696 2464 2704 2547
rect 2775 2533 2783 2582
rect 2835 2582 2843 2596
rect 2863 2596 2891 2602
rect 2851 2593 2903 2596
rect 2979 2596 2989 2606
rect 2917 2586 2929 2596
rect 2835 2575 2860 2582
rect 2917 2578 2955 2586
rect 2853 2553 2861 2575
rect 2775 2464 2783 2519
rect 2859 2504 2867 2539
rect 2517 2418 2529 2424
rect 2596 2418 2608 2424
rect 2646 2418 2658 2424
rect 2677 2418 2689 2424
rect 2751 2418 2763 2424
rect 2791 2418 2803 2424
rect 2938 2464 2946 2578
rect 2981 2553 2989 2596
rect 3029 2596 3057 2602
rect 3017 2593 3069 2596
rect 3259 2596 3269 2606
rect 3077 2582 3085 2596
rect 3139 2588 3151 2596
rect 3139 2582 3163 2588
rect 3060 2575 3085 2582
rect 2987 2539 2989 2553
rect 3059 2553 3067 2575
rect 2981 2504 2989 2539
rect 3053 2504 3061 2539
rect 3155 2533 3163 2582
rect 3197 2586 3209 2596
rect 3197 2578 3235 2586
rect 2836 2418 2848 2424
rect 2886 2418 2898 2424
rect 3155 2464 3163 2519
rect 3218 2464 3226 2578
rect 3261 2553 3269 2596
rect 3267 2539 3269 2553
rect 3316 2578 3334 2580
rect 3316 2569 3346 2578
rect 3397 2636 3409 2642
rect 3459 2636 3471 2642
rect 3567 2636 3579 2642
rect 3659 2636 3671 2642
rect 3717 2636 3729 2642
rect 3821 2636 3833 2642
rect 3912 2636 3924 2642
rect 3968 2636 3980 2642
rect 4049 2636 4061 2642
rect 4129 2636 4141 2642
rect 4177 2636 4189 2642
rect 4259 2636 4271 2642
rect 4410 2636 4422 2642
rect 4510 2636 4522 2642
rect 3316 2541 3324 2569
rect 3416 2561 3424 2616
rect 3489 2588 3501 2596
rect 3477 2582 3501 2588
rect 3599 2596 3609 2606
rect 3537 2586 3549 2596
rect 3261 2504 3269 2539
rect 2917 2418 2929 2424
rect 2961 2418 2973 2424
rect 3022 2418 3034 2424
rect 3072 2418 3084 2424
rect 3131 2418 3143 2424
rect 3171 2418 3183 2424
rect 3315 2472 3322 2527
rect 3315 2466 3362 2472
rect 3315 2464 3323 2466
rect 3351 2464 3362 2466
rect 3416 2464 3424 2547
rect 3477 2533 3485 2582
rect 3537 2578 3575 2586
rect 3477 2464 3485 2519
rect 3558 2464 3566 2578
rect 3601 2553 3609 2596
rect 3641 2590 3649 2616
rect 3641 2584 3663 2590
rect 3660 2578 3663 2584
rect 3607 2539 3609 2553
rect 3601 2504 3609 2539
rect 3660 2522 3667 2578
rect 3681 2553 3689 2596
rect 3736 2561 3744 2616
rect 3791 2596 3801 2606
rect 4169 2596 4197 2602
rect 3687 2539 3689 2553
rect 3791 2553 3799 2596
rect 3851 2586 3863 2596
rect 3825 2578 3863 2586
rect 3660 2516 3663 2522
rect 3637 2510 3663 2516
rect 3197 2418 3209 2424
rect 3241 2418 3253 2424
rect 3331 2418 3343 2424
rect 3371 2418 3383 2424
rect 3397 2418 3409 2424
rect 3457 2418 3469 2424
rect 3497 2418 3509 2424
rect 3637 2464 3645 2510
rect 3681 2504 3689 2539
rect 3736 2464 3744 2547
rect 3791 2539 3793 2553
rect 3791 2504 3799 2539
rect 3834 2464 3842 2578
rect 3940 2553 3947 2596
rect 4019 2588 4031 2596
rect 4099 2588 4111 2596
rect 4157 2593 4209 2596
rect 3987 2577 4003 2583
rect 4019 2582 4043 2588
rect 4099 2582 4123 2588
rect 4217 2582 4225 2596
rect 4289 2588 4301 2596
rect 3997 2547 4003 2577
rect 3933 2516 3939 2539
rect 4035 2533 4043 2582
rect 4115 2533 4123 2582
rect 4200 2575 4225 2582
rect 4277 2582 4301 2588
rect 4199 2553 4207 2575
rect 3912 2510 3939 2516
rect 3912 2504 3924 2510
rect 3903 2424 3931 2430
rect 3943 2496 3971 2502
rect 4035 2464 4043 2519
rect 4115 2464 4123 2519
rect 4193 2504 4201 2539
rect 4277 2533 4285 2582
rect 4356 2578 4374 2580
rect 4356 2569 4386 2578
rect 4456 2578 4474 2580
rect 4456 2569 4486 2578
rect 4540 2636 4552 2642
rect 4590 2636 4602 2642
rect 4710 2636 4722 2642
rect 4580 2596 4606 2607
rect 4356 2541 4364 2569
rect 4456 2541 4464 2569
rect 4598 2553 4606 2596
rect 4656 2578 4674 2580
rect 4656 2569 4686 2578
rect 3537 2418 3549 2424
rect 3581 2418 3593 2424
rect 3659 2418 3671 2424
rect 3717 2418 3729 2424
rect 3807 2418 3819 2424
rect 3851 2418 3863 2424
rect 3951 2418 3963 2424
rect 4011 2418 4023 2424
rect 4051 2418 4063 2424
rect 4091 2418 4103 2424
rect 4131 2418 4143 2424
rect 4277 2464 4285 2519
rect 4355 2472 4362 2527
rect 4656 2541 4664 2569
rect 4455 2472 4462 2527
rect 4598 2504 4606 2539
rect 4537 2498 4577 2504
rect 4537 2496 4549 2498
rect 4355 2466 4402 2472
rect 4355 2464 4363 2466
rect 4162 2418 4174 2424
rect 4212 2418 4224 2424
rect 4391 2464 4402 2466
rect 4455 2466 4502 2472
rect 4455 2464 4463 2466
rect 4491 2464 4502 2466
rect 4655 2472 4662 2527
rect 4655 2466 4702 2472
rect 4655 2464 4663 2466
rect 4691 2464 4702 2466
rect 4257 2418 4269 2424
rect 4297 2418 4309 2424
rect 4371 2418 4383 2424
rect 4411 2418 4423 2424
rect 4471 2418 4483 2424
rect 4511 2418 4523 2424
rect 4557 2418 4569 2424
rect 4671 2418 4683 2424
rect 4711 2418 4723 2424
rect -62 2416 4776 2418
rect -62 2404 4 2416
rect -62 2402 4776 2404
rect -62 1938 -2 2402
rect 41 2396 53 2402
rect 107 2396 119 2402
rect 153 2396 165 2402
rect 211 2396 223 2402
rect 262 2396 274 2402
rect 312 2396 324 2402
rect 377 2396 389 2402
rect 499 2396 511 2402
rect 557 2396 569 2402
rect 597 2396 609 2402
rect 671 2396 683 2402
rect 77 2350 85 2356
rect 127 2350 139 2356
rect 67 2336 85 2350
rect 113 2338 135 2350
rect 181 2342 193 2376
rect 77 2330 85 2336
rect 77 2322 115 2330
rect 133 2326 163 2332
rect 21 2308 83 2316
rect 21 2224 27 2308
rect 133 2312 139 2326
rect 181 2318 187 2336
rect 95 2306 139 2312
rect 147 2312 187 2318
rect 66 2267 93 2274
rect 40 2256 46 2261
rect 40 2248 74 2256
rect 79 2240 86 2248
rect 147 2240 153 2312
rect 369 2318 397 2324
rect 409 2390 437 2396
rect 207 2304 221 2312
rect 213 2253 227 2267
rect 235 2253 243 2316
rect 293 2281 301 2316
rect 416 2310 428 2316
rect 401 2304 428 2310
rect 477 2310 485 2356
rect 697 2396 709 2402
rect 831 2396 843 2402
rect 877 2396 889 2402
rect 957 2396 969 2402
rect 1037 2396 1049 2402
rect 1117 2396 1129 2402
rect 1175 2396 1187 2402
rect 1221 2396 1233 2402
rect 1287 2396 1299 2402
rect 1342 2396 1354 2402
rect 1392 2396 1404 2402
rect 1457 2396 1469 2402
rect 1515 2396 1527 2402
rect 1561 2396 1573 2402
rect 1627 2396 1639 2402
rect 1731 2396 1743 2402
rect 1811 2396 1823 2402
rect 1857 2396 1869 2402
rect 1971 2396 1983 2402
rect 477 2304 503 2310
rect 401 2281 407 2304
rect 500 2298 503 2304
rect 79 2234 153 2240
rect 227 2239 243 2253
rect 299 2245 307 2267
rect 79 2228 86 2234
rect 147 2232 153 2234
rect 111 2216 132 2223
rect 235 2224 243 2239
rect 300 2238 325 2245
rect 60 2204 67 2210
rect 125 2204 132 2216
rect 182 2210 193 2218
rect 182 2204 189 2210
rect 60 2198 73 2204
rect 257 2224 309 2227
rect 269 2218 297 2224
rect 317 2224 325 2238
rect 393 2224 400 2267
rect 500 2242 507 2298
rect 521 2281 529 2316
rect 577 2301 585 2356
rect 527 2267 529 2281
rect 500 2236 503 2242
rect 481 2230 503 2236
rect 481 2204 489 2230
rect 521 2224 529 2267
rect 577 2238 585 2287
rect 656 2273 664 2356
rect 851 2322 863 2324
rect 823 2316 863 2322
rect 720 2309 737 2316
rect 720 2261 727 2309
rect 794 2281 802 2316
rect 900 2309 917 2316
rect 980 2309 997 2316
rect 577 2232 601 2238
rect 589 2224 601 2232
rect 656 2204 664 2259
rect 720 2204 727 2247
rect 794 2224 802 2267
rect 900 2261 907 2309
rect 980 2261 987 2309
rect 1056 2273 1064 2356
rect 1147 2342 1159 2376
rect 1201 2350 1213 2356
rect 1255 2350 1263 2356
rect 1205 2338 1227 2350
rect 1255 2336 1273 2350
rect 1153 2318 1159 2336
rect 1177 2326 1207 2332
rect 1255 2330 1263 2336
rect 794 2213 820 2224
rect 41 2178 53 2184
rect 103 2178 115 2184
rect 151 2178 163 2184
rect 209 2178 221 2184
rect 277 2178 289 2184
rect 360 2178 372 2184
rect 416 2178 428 2184
rect 499 2178 511 2184
rect 559 2178 571 2184
rect 671 2178 683 2184
rect 697 2178 709 2184
rect 737 2178 749 2184
rect 900 2204 907 2247
rect 980 2204 987 2247
rect 1056 2204 1064 2259
rect 1097 2253 1105 2316
rect 1119 2304 1133 2312
rect 1153 2312 1193 2318
rect 1113 2253 1127 2267
rect 1097 2239 1113 2253
rect 1187 2240 1193 2312
rect 1201 2312 1207 2326
rect 1225 2322 1263 2330
rect 1487 2342 1499 2376
rect 1541 2350 1553 2356
rect 1595 2350 1603 2356
rect 1545 2338 1567 2350
rect 1595 2336 1613 2350
rect 1493 2318 1499 2336
rect 1517 2326 1547 2332
rect 1595 2330 1603 2336
rect 1201 2306 1245 2312
rect 1257 2308 1319 2316
rect 1247 2267 1274 2274
rect 1294 2256 1300 2261
rect 1266 2248 1300 2256
rect 1254 2240 1261 2248
rect 1097 2224 1105 2239
rect 1187 2234 1261 2240
rect 1187 2232 1193 2234
rect 798 2178 810 2184
rect 848 2178 860 2184
rect 877 2178 889 2184
rect 917 2178 929 2184
rect 957 2178 969 2184
rect 997 2178 1009 2184
rect 1254 2228 1261 2234
rect 1147 2210 1158 2218
rect 1151 2204 1158 2210
rect 1208 2216 1229 2223
rect 1313 2224 1319 2308
rect 1373 2281 1381 2316
rect 1379 2245 1387 2267
rect 1437 2253 1445 2316
rect 1459 2304 1473 2312
rect 1493 2312 1533 2318
rect 1453 2253 1467 2267
rect 1380 2238 1405 2245
rect 1208 2204 1215 2216
rect 1273 2204 1280 2210
rect 1267 2198 1280 2204
rect 1337 2224 1389 2227
rect 1349 2218 1377 2224
rect 1397 2224 1405 2238
rect 1437 2239 1453 2253
rect 1527 2240 1533 2312
rect 1541 2312 1547 2326
rect 1565 2322 1603 2330
rect 1541 2306 1585 2312
rect 1597 2308 1659 2316
rect 1831 2322 1843 2324
rect 1803 2316 1843 2322
rect 1997 2396 2009 2402
rect 2037 2396 2049 2402
rect 2077 2396 2089 2402
rect 2117 2396 2129 2402
rect 2157 2396 2169 2402
rect 2202 2396 2214 2402
rect 2252 2396 2264 2402
rect 2321 2396 2333 2402
rect 2387 2396 2399 2402
rect 2433 2396 2445 2402
rect 2491 2396 2503 2402
rect 2551 2396 2563 2402
rect 2591 2396 2603 2402
rect 2357 2350 2365 2356
rect 2407 2350 2419 2356
rect 2347 2336 2365 2350
rect 2393 2338 2415 2350
rect 2461 2342 2473 2376
rect 2357 2330 2365 2336
rect 2357 2322 2395 2330
rect 2413 2326 2443 2332
rect 1703 2309 1720 2316
rect 1587 2267 1614 2274
rect 1634 2256 1640 2261
rect 1606 2248 1640 2256
rect 1594 2240 1601 2248
rect 1437 2224 1445 2239
rect 1527 2234 1601 2240
rect 1527 2232 1533 2234
rect 1594 2228 1601 2234
rect 1487 2210 1498 2218
rect 1491 2204 1498 2210
rect 1548 2216 1569 2223
rect 1653 2224 1659 2308
rect 1548 2204 1555 2216
rect 1613 2204 1620 2210
rect 1607 2198 1620 2204
rect 1713 2261 1720 2309
rect 1774 2281 1782 2316
rect 1876 2281 1884 2316
rect 1943 2309 1960 2316
rect 1713 2204 1720 2247
rect 1774 2224 1782 2267
rect 1876 2224 1884 2267
rect 1953 2261 1960 2309
rect 2017 2310 2029 2316
rect 2057 2310 2069 2316
rect 2097 2310 2109 2316
rect 2137 2310 2149 2316
rect 2017 2302 2043 2310
rect 2057 2302 2082 2310
rect 2097 2302 2122 2310
rect 2137 2302 2155 2310
rect 2035 2256 2043 2302
rect 2074 2256 2082 2302
rect 2114 2256 2122 2302
rect 2148 2273 2155 2302
rect 2233 2281 2241 2316
rect 2301 2308 2363 2316
rect 2148 2259 2153 2273
rect 1774 2213 1800 2224
rect 1037 2178 1049 2184
rect 1119 2178 1131 2184
rect 1177 2178 1189 2184
rect 1225 2178 1237 2184
rect 1287 2178 1299 2184
rect 1357 2178 1369 2184
rect 1459 2178 1471 2184
rect 1517 2178 1529 2184
rect 1565 2178 1577 2184
rect 1627 2178 1639 2184
rect 1691 2178 1703 2184
rect 1731 2178 1743 2184
rect 1778 2178 1790 2184
rect 1828 2178 1840 2184
rect 1953 2204 1960 2247
rect 2035 2244 2050 2256
rect 2074 2244 2090 2256
rect 2114 2244 2130 2256
rect 2035 2238 2043 2244
rect 2074 2238 2082 2244
rect 2114 2238 2122 2244
rect 2148 2238 2155 2259
rect 2239 2245 2247 2267
rect 2240 2238 2265 2245
rect 2016 2230 2043 2238
rect 2057 2230 2082 2238
rect 2096 2230 2122 2238
rect 2136 2231 2155 2238
rect 2136 2230 2154 2231
rect 2016 2224 2028 2230
rect 2057 2224 2069 2230
rect 2096 2224 2108 2230
rect 2136 2224 2148 2230
rect 2197 2224 2249 2227
rect 1857 2178 1869 2184
rect 1931 2178 1943 2184
rect 1971 2178 1983 2184
rect 2209 2218 2237 2224
rect 2257 2224 2265 2238
rect 2301 2224 2307 2308
rect 2413 2312 2419 2326
rect 2461 2318 2467 2336
rect 2375 2306 2419 2312
rect 2427 2312 2467 2318
rect 2346 2267 2373 2274
rect 2320 2256 2326 2261
rect 2320 2248 2354 2256
rect 2359 2240 2366 2248
rect 2427 2240 2433 2312
rect 2617 2396 2629 2402
rect 2657 2396 2669 2402
rect 2697 2396 2709 2402
rect 2737 2396 2749 2402
rect 2796 2396 2808 2402
rect 2846 2396 2858 2402
rect 2487 2304 2501 2312
rect 2493 2253 2507 2267
rect 2515 2253 2523 2316
rect 2575 2301 2583 2356
rect 2637 2301 2645 2356
rect 2717 2301 2725 2356
rect 2896 2396 2908 2402
rect 2946 2396 2958 2402
rect 3001 2396 3013 2402
rect 3067 2396 3079 2402
rect 3113 2396 3125 2402
rect 3171 2396 3183 2402
rect 3222 2396 3234 2402
rect 3272 2396 3284 2402
rect 3037 2350 3045 2356
rect 3087 2350 3099 2356
rect 3027 2336 3045 2350
rect 3073 2338 3095 2350
rect 3141 2342 3153 2376
rect 3037 2330 3045 2336
rect 3037 2322 3075 2330
rect 3093 2326 3123 2332
rect 2359 2234 2433 2240
rect 2507 2239 2523 2253
rect 2359 2228 2366 2234
rect 2427 2232 2433 2234
rect 2391 2216 2412 2223
rect 2515 2224 2523 2239
rect 2575 2238 2583 2287
rect 2340 2204 2347 2210
rect 2405 2204 2412 2216
rect 2462 2210 2473 2218
rect 2462 2204 2469 2210
rect 2340 2198 2353 2204
rect 2559 2232 2583 2238
rect 2637 2238 2645 2287
rect 2717 2238 2725 2287
rect 2819 2281 2827 2316
rect 2919 2281 2927 2316
rect 2981 2308 3043 2316
rect 2813 2245 2821 2267
rect 2913 2245 2921 2267
rect 2795 2238 2820 2245
rect 2895 2238 2920 2245
rect 2637 2232 2661 2238
rect 2717 2232 2741 2238
rect 2559 2224 2571 2232
rect 2649 2224 2661 2232
rect 2729 2224 2741 2232
rect 2795 2224 2803 2238
rect 1997 2178 2009 2184
rect 2037 2178 2049 2184
rect 2077 2178 2089 2184
rect 2117 2178 2129 2184
rect 2157 2178 2169 2184
rect 2217 2178 2229 2184
rect 2321 2178 2333 2184
rect 2383 2178 2395 2184
rect 2431 2178 2443 2184
rect 2489 2178 2501 2184
rect 2589 2178 2601 2184
rect 2811 2224 2863 2227
rect 2895 2224 2903 2238
rect 2823 2218 2851 2224
rect 2911 2224 2963 2227
rect 2923 2218 2951 2224
rect 2981 2224 2987 2308
rect 3093 2312 3099 2326
rect 3141 2318 3147 2336
rect 3055 2306 3099 2312
rect 3107 2312 3147 2318
rect 3026 2267 3053 2274
rect 3000 2256 3006 2261
rect 3000 2248 3034 2256
rect 3039 2240 3046 2248
rect 3107 2240 3113 2312
rect 3317 2396 3329 2402
rect 3357 2396 3369 2402
rect 3397 2396 3409 2402
rect 3437 2396 3449 2402
rect 3491 2396 3503 2402
rect 3531 2396 3543 2402
rect 3591 2396 3603 2402
rect 3651 2396 3663 2402
rect 3711 2396 3723 2402
rect 3287 2337 3303 2343
rect 3167 2304 3181 2312
rect 3173 2253 3187 2267
rect 3195 2253 3203 2316
rect 3253 2281 3261 2316
rect 3039 2234 3113 2240
rect 3187 2239 3203 2253
rect 3259 2245 3267 2267
rect 3297 2263 3303 2337
rect 3337 2301 3345 2356
rect 3417 2301 3425 2356
rect 3515 2301 3523 2356
rect 3742 2396 3754 2402
rect 3792 2396 3804 2402
rect 3869 2396 3881 2402
rect 3917 2396 3929 2402
rect 3977 2396 3989 2402
rect 4021 2396 4033 2402
rect 4096 2396 4108 2402
rect 4146 2396 4158 2402
rect 4211 2396 4223 2402
rect 4251 2396 4263 2402
rect 4297 2396 4309 2402
rect 4396 2396 4408 2402
rect 4446 2396 4458 2402
rect 3287 2257 3303 2263
rect 3039 2228 3046 2234
rect 3107 2232 3113 2234
rect 3071 2216 3092 2223
rect 3195 2224 3203 2239
rect 3260 2238 3285 2245
rect 3020 2204 3027 2210
rect 3085 2204 3092 2216
rect 3142 2210 3153 2218
rect 3142 2204 3149 2210
rect 3020 2198 3033 2204
rect 3217 2224 3269 2227
rect 3229 2218 3257 2224
rect 3277 2224 3285 2238
rect 3337 2238 3345 2287
rect 3417 2238 3425 2287
rect 3515 2238 3523 2287
rect 3576 2281 3584 2316
rect 3636 2281 3644 2316
rect 3337 2232 3361 2238
rect 3417 2232 3441 2238
rect 3349 2224 3361 2232
rect 3429 2224 3441 2232
rect 3499 2232 3523 2238
rect 3499 2224 3511 2232
rect 3576 2224 3584 2267
rect 3696 2273 3704 2356
rect 3773 2281 3781 2316
rect 3851 2281 3859 2316
rect 3895 2310 3903 2356
rect 3877 2304 3903 2310
rect 3877 2298 3880 2304
rect 3636 2224 3644 2267
rect 3696 2204 3704 2259
rect 3779 2245 3787 2267
rect 3851 2267 3853 2281
rect 3780 2238 3805 2245
rect 3737 2224 3789 2227
rect 3749 2218 3777 2224
rect 3797 2224 3805 2238
rect 3851 2224 3859 2267
rect 3873 2242 3880 2298
rect 3936 2281 3944 2316
rect 3877 2236 3880 2242
rect 3877 2230 3899 2236
rect 3891 2204 3899 2230
rect 3936 2224 3944 2267
rect 3998 2242 4006 2356
rect 4195 2354 4203 2356
rect 4231 2354 4242 2356
rect 4195 2348 4242 2354
rect 4041 2281 4049 2316
rect 4119 2281 4127 2316
rect 4195 2293 4202 2348
rect 4277 2322 4289 2324
rect 4277 2316 4317 2322
rect 4482 2396 4494 2402
rect 4532 2396 4544 2402
rect 4596 2396 4608 2402
rect 4646 2396 4658 2402
rect 4697 2396 4709 2402
rect 4677 2322 4689 2324
rect 4677 2316 4717 2322
rect 4047 2267 4049 2281
rect 3977 2234 4015 2242
rect 3977 2224 3989 2234
rect 4041 2224 4049 2267
rect 4113 2245 4121 2267
rect 4338 2281 4346 2316
rect 4419 2281 4427 2316
rect 4513 2281 4521 2316
rect 4619 2281 4627 2316
rect 4738 2281 4746 2316
rect 4095 2238 4120 2245
rect 4095 2224 4103 2238
rect 4177 2243 4183 2253
rect 4167 2237 4183 2243
rect 4196 2251 4204 2279
rect 4196 2242 4226 2251
rect 4196 2240 4214 2242
rect 4039 2214 4049 2224
rect 4111 2224 4163 2227
rect 4123 2218 4151 2224
rect 4338 2224 4346 2267
rect 4413 2245 4421 2267
rect 4519 2245 4527 2267
rect 4613 2245 4621 2267
rect 4395 2238 4420 2245
rect 4520 2238 4545 2245
rect 4395 2224 4403 2238
rect 2619 2178 2631 2184
rect 2699 2178 2711 2184
rect 2831 2178 2843 2184
rect 2931 2178 2943 2184
rect 3001 2178 3013 2184
rect 3063 2178 3075 2184
rect 3111 2178 3123 2184
rect 3169 2178 3181 2184
rect 3237 2178 3249 2184
rect 3319 2178 3331 2184
rect 3399 2178 3411 2184
rect 3529 2178 3541 2184
rect 3591 2178 3603 2184
rect 3651 2178 3663 2184
rect 3711 2178 3723 2184
rect 3757 2178 3769 2184
rect 3869 2178 3881 2184
rect 3917 2178 3929 2184
rect 4007 2178 4019 2184
rect 4131 2178 4143 2184
rect 4250 2178 4262 2184
rect 4320 2213 4346 2224
rect 4411 2224 4463 2227
rect 4423 2218 4451 2224
rect 4477 2224 4529 2227
rect 4489 2218 4517 2224
rect 4537 2224 4545 2238
rect 4595 2238 4620 2245
rect 4595 2224 4603 2238
rect 4611 2224 4663 2227
rect 4738 2224 4746 2267
rect 4623 2218 4651 2224
rect 4720 2213 4746 2224
rect 4280 2178 4292 2184
rect 4330 2178 4342 2184
rect 4431 2178 4443 2184
rect 4497 2178 4509 2184
rect 4631 2178 4643 2184
rect 4680 2178 4692 2184
rect 4730 2178 4742 2184
rect 4782 2178 4842 2642
rect 4 2176 4842 2178
rect 4776 2164 4842 2176
rect 4 2162 4842 2164
rect 17 2156 29 2162
rect 57 2156 69 2162
rect 97 2156 109 2162
rect 137 2156 149 2162
rect 177 2156 189 2162
rect 269 2156 281 2162
rect 351 2156 363 2162
rect 400 2156 412 2162
rect 456 2156 468 2162
rect 541 2156 553 2162
rect 603 2156 615 2162
rect 651 2156 663 2162
rect 709 2156 721 2162
rect 809 2156 821 2162
rect 871 2156 883 2162
rect 915 2156 923 2162
rect 36 2110 48 2116
rect 77 2110 89 2116
rect 116 2110 128 2116
rect 156 2110 168 2116
rect 36 2102 63 2110
rect 77 2102 102 2110
rect 116 2102 142 2110
rect 156 2109 174 2110
rect 156 2102 175 2109
rect 239 2108 251 2116
rect 239 2102 263 2108
rect 55 2096 63 2102
rect 94 2096 102 2102
rect 134 2096 142 2102
rect 55 2084 70 2096
rect 94 2084 110 2096
rect 134 2084 150 2096
rect 55 2038 63 2084
rect 94 2038 102 2084
rect 134 2038 142 2084
rect 168 2081 175 2102
rect 168 2067 173 2081
rect 168 2038 175 2067
rect 255 2053 263 2102
rect 315 2102 323 2116
rect 343 2116 371 2122
rect 560 2136 573 2142
rect 560 2130 567 2136
rect 625 2124 632 2136
rect 331 2113 383 2116
rect 315 2095 340 2102
rect 297 2077 313 2083
rect 37 2030 63 2038
rect 77 2030 102 2038
rect 117 2030 142 2038
rect 157 2030 175 2038
rect 37 2024 49 2030
rect 77 2024 89 2030
rect 117 2024 129 2030
rect 157 2024 169 2030
rect 255 1984 263 2039
rect 297 2003 303 2077
rect 333 2073 341 2095
rect 433 2073 440 2116
rect 339 2024 347 2059
rect 441 2036 447 2059
rect 441 2030 468 2036
rect 456 2024 468 2030
rect 521 2032 527 2116
rect 611 2117 632 2124
rect 682 2130 689 2136
rect 682 2122 693 2130
rect 579 2106 586 2112
rect 647 2106 653 2108
rect 579 2100 653 2106
rect 735 2101 743 2116
rect 939 2156 951 2162
rect 1017 2156 1029 2162
rect 1057 2156 1069 2162
rect 1117 2156 1129 2162
rect 1199 2156 1211 2162
rect 1277 2156 1289 2162
rect 1317 2156 1329 2162
rect 1379 2156 1391 2162
rect 1437 2156 1449 2162
rect 1485 2156 1497 2162
rect 1547 2156 1559 2162
rect 1618 2156 1630 2162
rect 1668 2156 1680 2162
rect 1729 2156 1741 2162
rect 1799 2156 1811 2162
rect 1857 2156 1869 2162
rect 1905 2156 1917 2162
rect 1967 2156 1979 2162
rect 2051 2156 2063 2162
rect 2129 2156 2141 2162
rect 2179 2156 2191 2162
rect 2239 2156 2251 2162
rect 2371 2156 2383 2162
rect 2469 2156 2481 2162
rect 2549 2156 2561 2162
rect 2631 2156 2643 2162
rect 2731 2156 2743 2162
rect 2801 2156 2813 2162
rect 2863 2156 2875 2162
rect 2911 2156 2923 2162
rect 2969 2156 2981 2162
rect 3047 2156 3059 2162
rect 3171 2156 3183 2162
rect 3271 2156 3283 2162
rect 3319 2156 3331 2162
rect 3451 2156 3463 2162
rect 3498 2156 3510 2162
rect 3597 2156 3609 2162
rect 3658 2156 3670 2162
rect 3759 2156 3771 2162
rect 3859 2156 3871 2162
rect 3937 2156 3949 2162
rect 4069 2156 4081 2162
rect 4149 2156 4161 2162
rect 4229 2156 4241 2162
rect 4287 2156 4299 2162
rect 4360 2156 4372 2162
rect 4410 2156 4422 2162
rect 779 2108 791 2116
rect 779 2102 803 2108
rect 579 2092 586 2100
rect 540 2084 574 2092
rect 540 2079 546 2084
rect 566 2066 593 2073
rect 521 2024 583 2032
rect 595 2028 639 2034
rect 297 1997 313 2003
rect 17 1938 29 1944
rect 57 1938 69 1944
rect 97 1938 109 1944
rect 137 1938 149 1944
rect 177 1938 189 1944
rect 231 1938 243 1944
rect 271 1938 283 1944
rect 409 2016 437 2022
rect 449 1944 477 1950
rect 577 2010 615 2018
rect 633 2014 639 2028
rect 647 2028 653 2100
rect 727 2087 743 2101
rect 713 2073 727 2087
rect 647 2022 687 2028
rect 707 2028 721 2036
rect 735 2024 743 2087
rect 795 2053 803 2102
rect 853 2081 860 2116
rect 891 2108 897 2136
rect 969 2108 981 2116
rect 887 2102 897 2108
rect 957 2102 981 2108
rect 577 2004 585 2010
rect 633 2008 663 2014
rect 681 2004 687 2022
rect 567 1990 585 2004
rect 613 1990 635 2002
rect 577 1984 585 1990
rect 627 1984 639 1990
rect 681 1964 693 1998
rect 795 1984 803 2039
rect 857 2023 866 2067
rect 876 2041 882 2096
rect 957 2053 965 2102
rect 1040 2093 1047 2136
rect 1109 2116 1137 2122
rect 1097 2113 1149 2116
rect 1157 2102 1165 2116
rect 1229 2108 1241 2116
rect 1140 2095 1165 2102
rect 1217 2102 1241 2108
rect 887 2032 923 2040
rect 915 2024 923 2032
rect 857 2014 861 2023
rect 957 1984 965 2039
rect 1040 2031 1047 2079
rect 1139 2073 1147 2095
rect 1040 2024 1057 2031
rect 1133 2024 1141 2059
rect 1217 2053 1225 2102
rect 1300 2093 1307 2136
rect 316 1938 328 1944
rect 366 1938 378 1944
rect 417 1938 429 1944
rect 541 1938 553 1944
rect 607 1938 619 1944
rect 653 1938 665 1944
rect 711 1938 723 1944
rect 771 1938 783 1944
rect 811 1938 823 1944
rect 881 1938 893 1944
rect 937 1938 949 1944
rect 977 1938 989 1944
rect 1217 1984 1225 2039
rect 1300 2031 1307 2079
rect 1527 2136 1540 2142
rect 1411 2130 1418 2136
rect 1407 2122 1418 2130
rect 1468 2124 1475 2136
rect 1533 2130 1540 2136
rect 1357 2101 1365 2116
rect 1468 2117 1489 2124
rect 1447 2106 1453 2108
rect 1514 2106 1521 2112
rect 1357 2087 1373 2101
rect 1447 2100 1521 2106
rect 1300 2024 1317 2031
rect 1017 1938 1029 1944
rect 1102 1938 1114 1944
rect 1152 1938 1164 1944
rect 1197 1938 1209 1944
rect 1237 1938 1249 1944
rect 1357 2024 1365 2087
rect 1373 2073 1387 2087
rect 1379 2028 1393 2036
rect 1447 2028 1453 2100
rect 1514 2092 1521 2100
rect 1526 2084 1560 2092
rect 1554 2079 1560 2084
rect 1507 2066 1534 2073
rect 1413 2022 1453 2028
rect 1461 2028 1505 2034
rect 1413 2004 1419 2022
rect 1461 2014 1467 2028
rect 1573 2032 1579 2116
rect 1614 2116 1640 2127
rect 1614 2073 1622 2116
rect 1711 2073 1719 2116
rect 1751 2110 1759 2136
rect 1737 2104 1759 2110
rect 1947 2136 1960 2142
rect 1831 2130 1838 2136
rect 1827 2122 1838 2130
rect 1888 2124 1895 2136
rect 1953 2130 1960 2136
rect 1737 2098 1740 2104
rect 1711 2059 1713 2073
rect 1517 2024 1579 2032
rect 1614 2024 1622 2059
rect 1711 2024 1719 2059
rect 1733 2042 1740 2098
rect 1777 2101 1785 2116
rect 1888 2117 1909 2124
rect 1867 2106 1873 2108
rect 1934 2106 1941 2112
rect 1777 2087 1793 2101
rect 1867 2100 1941 2106
rect 1737 2036 1740 2042
rect 1737 2030 1763 2036
rect 1437 2008 1467 2014
rect 1485 2010 1523 2018
rect 1515 2004 1523 2010
rect 1407 1964 1419 1998
rect 1465 1990 1487 2002
rect 1515 1990 1533 2004
rect 1461 1984 1473 1990
rect 1515 1984 1523 1990
rect 1643 2018 1683 2024
rect 1671 2016 1683 2018
rect 1755 1984 1763 2030
rect 1777 2024 1785 2087
rect 1793 2073 1807 2087
rect 1799 2028 1813 2036
rect 1867 2028 1873 2100
rect 1934 2092 1941 2100
rect 1946 2084 1980 2092
rect 1974 2079 1980 2084
rect 1927 2066 1954 2073
rect 1833 2022 1873 2028
rect 1881 2028 1925 2034
rect 1833 2004 1839 2022
rect 1881 2014 1887 2028
rect 1993 2032 1999 2116
rect 2036 2081 2044 2136
rect 2099 2108 2111 2116
rect 2161 2110 2169 2136
rect 2099 2102 2123 2108
rect 2161 2104 2183 2110
rect 1937 2024 1999 2032
rect 1857 2008 1887 2014
rect 1905 2010 1943 2018
rect 1935 2004 1943 2010
rect 1827 1964 1839 1998
rect 1885 1990 1907 2002
rect 1935 1990 1953 2004
rect 1881 1984 1893 1990
rect 1935 1984 1943 1990
rect 2036 1984 2044 2067
rect 2115 2053 2123 2102
rect 2180 2098 2183 2104
rect 2180 2042 2187 2098
rect 2201 2073 2209 2116
rect 2269 2108 2281 2116
rect 2257 2102 2281 2108
rect 2335 2102 2343 2116
rect 2363 2116 2391 2122
rect 2351 2113 2403 2116
rect 2439 2108 2451 2116
rect 2519 2108 2531 2116
rect 2439 2102 2463 2108
rect 2207 2059 2209 2073
rect 2115 1984 2123 2039
rect 2180 2036 2183 2042
rect 2157 2030 2183 2036
rect 2157 1984 2165 2030
rect 2201 2024 2209 2059
rect 2257 2053 2265 2102
rect 2335 2095 2360 2102
rect 2353 2073 2361 2095
rect 1277 1938 1289 1944
rect 1377 1938 1389 1944
rect 1435 1938 1447 1944
rect 1481 1938 1493 1944
rect 1547 1938 1559 1944
rect 1651 1938 1663 1944
rect 1729 1938 1741 1944
rect 1797 1938 1809 1944
rect 1855 1938 1867 1944
rect 1901 1938 1913 1944
rect 1967 1938 1979 1944
rect 2051 1938 2063 1944
rect 2257 1984 2265 2039
rect 2359 2024 2367 2059
rect 2455 2053 2463 2102
rect 2487 2097 2503 2103
rect 2519 2102 2543 2108
rect 2091 1938 2103 1944
rect 2131 1938 2143 1944
rect 2179 1938 2191 1944
rect 2237 1938 2249 1944
rect 2277 1938 2289 1944
rect 2455 1984 2463 2039
rect 2497 2023 2503 2097
rect 2535 2053 2543 2102
rect 2595 2102 2603 2116
rect 2623 2116 2651 2122
rect 2611 2113 2663 2116
rect 2695 2102 2703 2116
rect 2723 2116 2751 2122
rect 2711 2113 2763 2116
rect 2820 2136 2833 2142
rect 2820 2130 2827 2136
rect 2885 2124 2892 2136
rect 2595 2095 2620 2102
rect 2695 2095 2720 2102
rect 2613 2073 2621 2095
rect 2713 2073 2721 2095
rect 2497 2017 2513 2023
rect 2535 1984 2543 2039
rect 2619 2024 2627 2059
rect 2719 2024 2727 2059
rect 2781 2032 2787 2116
rect 2871 2117 2892 2124
rect 2942 2130 2949 2136
rect 2942 2122 2953 2130
rect 2839 2106 2846 2112
rect 2907 2106 2913 2108
rect 2839 2100 2913 2106
rect 2995 2101 3003 2116
rect 2839 2092 2846 2100
rect 2800 2084 2834 2092
rect 2800 2079 2806 2084
rect 2826 2066 2853 2073
rect 2781 2024 2843 2032
rect 2855 2028 2899 2034
rect 2336 1938 2348 1944
rect 2386 1938 2398 1944
rect 2431 1938 2443 1944
rect 2471 1938 2483 1944
rect 2511 1938 2523 1944
rect 2551 1938 2563 1944
rect 2596 1938 2608 1944
rect 2646 1938 2658 1944
rect 2837 2010 2875 2018
rect 2893 2014 2899 2028
rect 2907 2028 2913 2100
rect 2987 2087 3003 2101
rect 3079 2116 3089 2126
rect 3017 2106 3029 2116
rect 3017 2098 3055 2106
rect 2973 2073 2987 2087
rect 2907 2022 2947 2028
rect 2967 2028 2981 2036
rect 2995 2024 3003 2087
rect 2837 2004 2845 2010
rect 2893 2008 2923 2014
rect 2941 2004 2947 2022
rect 2827 1990 2845 2004
rect 2873 1990 2895 2002
rect 2837 1984 2845 1990
rect 2887 1984 2899 1990
rect 2941 1964 2953 1998
rect 3038 1984 3046 2098
rect 3081 2073 3089 2116
rect 3135 2102 3143 2116
rect 3163 2116 3191 2122
rect 3151 2113 3203 2116
rect 3235 2102 3243 2116
rect 3263 2116 3291 2122
rect 3251 2113 3303 2116
rect 3349 2108 3361 2116
rect 3337 2102 3361 2108
rect 3415 2102 3423 2116
rect 3443 2116 3471 2122
rect 3431 2113 3483 2116
rect 3135 2095 3160 2102
rect 3235 2095 3260 2102
rect 3087 2059 3089 2073
rect 3081 2024 3089 2059
rect 3117 2077 3133 2083
rect 3117 2027 3123 2077
rect 3153 2073 3161 2095
rect 3253 2073 3261 2095
rect 3159 2024 3167 2059
rect 3259 2024 3267 2059
rect 3337 2053 3345 2102
rect 3415 2095 3440 2102
rect 3546 2098 3564 2100
rect 3433 2073 3441 2095
rect 3534 2089 3564 2098
rect 2696 1938 2708 1944
rect 2746 1938 2758 1944
rect 2801 1938 2813 1944
rect 2867 1938 2879 1944
rect 2913 1938 2925 1944
rect 2971 1938 2983 1944
rect 3017 1938 3029 1944
rect 3061 1938 3073 1944
rect 3136 1938 3148 1944
rect 3186 1938 3198 1944
rect 3337 1984 3345 2039
rect 3377 2023 3383 2073
rect 3556 2061 3564 2089
rect 3616 2081 3624 2136
rect 3789 2108 3801 2116
rect 3777 2102 3801 2108
rect 3841 2110 3849 2136
rect 3929 2116 3957 2122
rect 3841 2104 3863 2110
rect 3706 2098 3724 2100
rect 3694 2089 3724 2098
rect 3637 2077 3653 2083
rect 3439 2024 3447 2059
rect 3367 2017 3383 2023
rect 3236 1938 3248 1944
rect 3286 1938 3298 1944
rect 3317 1938 3329 1944
rect 3357 1938 3369 1944
rect 3558 1992 3565 2047
rect 3518 1986 3565 1992
rect 3518 1984 3529 1986
rect 3416 1938 3428 1944
rect 3466 1938 3478 1944
rect 3557 1984 3565 1986
rect 3616 1984 3624 2067
rect 3637 2007 3643 2077
rect 3716 2061 3724 2089
rect 3777 2053 3785 2102
rect 3860 2098 3863 2104
rect 3718 1992 3725 2047
rect 3860 2042 3867 2098
rect 3881 2073 3889 2116
rect 3917 2113 3969 2116
rect 4319 2116 4329 2126
rect 4478 2156 4490 2162
rect 4528 2156 4540 2162
rect 4400 2116 4426 2127
rect 3977 2102 3985 2116
rect 4039 2108 4051 2116
rect 4119 2108 4131 2116
rect 4199 2108 4211 2116
rect 4039 2102 4063 2108
rect 4119 2102 4143 2108
rect 3960 2095 3985 2102
rect 3887 2059 3889 2073
rect 3959 2073 3967 2095
rect 3678 1986 3725 1992
rect 3678 1984 3689 1986
rect 3717 1984 3725 1986
rect 3777 1984 3785 2039
rect 3860 2036 3863 2042
rect 3837 2030 3863 2036
rect 3837 1984 3845 2030
rect 3881 2024 3889 2059
rect 3953 2024 3961 2059
rect 4055 2053 4063 2102
rect 4135 2053 4143 2102
rect 4167 2097 4183 2103
rect 4199 2102 4223 2108
rect 3987 1997 3993 2003
rect 4007 1997 4033 2003
rect 4055 1984 4063 2039
rect 4135 1984 4143 2039
rect 4177 2023 4183 2097
rect 4215 2053 4223 2102
rect 4257 2106 4269 2116
rect 4257 2098 4295 2106
rect 4167 2017 4183 2023
rect 4215 1984 4223 2039
rect 4278 1984 4286 2098
rect 4321 2073 4329 2116
rect 4327 2059 4329 2073
rect 4418 2073 4426 2116
rect 4474 2116 4500 2127
rect 4558 2156 4570 2162
rect 4658 2156 4670 2162
rect 4474 2073 4482 2116
rect 4606 2098 4624 2100
rect 4594 2089 4624 2098
rect 4706 2098 4724 2100
rect 4694 2089 4724 2098
rect 4616 2061 4624 2089
rect 4716 2061 4724 2089
rect 4321 2024 4329 2059
rect 4418 2024 4426 2059
rect 4474 2024 4482 2059
rect 3497 1938 3509 1944
rect 3537 1938 3549 1944
rect 3597 1938 3609 1944
rect 3657 1938 3669 1944
rect 3697 1938 3709 1944
rect 3757 1938 3769 1944
rect 3797 1938 3809 1944
rect 3859 1938 3871 1944
rect 3922 1938 3934 1944
rect 3972 1938 3984 1944
rect 4031 1938 4043 1944
rect 4071 1938 4083 1944
rect 4111 1938 4123 1944
rect 4151 1938 4163 1944
rect 4191 1938 4203 1944
rect 4231 1938 4243 1944
rect 4357 2018 4397 2024
rect 4357 2016 4369 2018
rect 4503 2018 4543 2024
rect 4531 2016 4543 2018
rect 4618 1992 4625 2047
rect 4718 1992 4725 2047
rect 4578 1986 4625 1992
rect 4578 1984 4589 1986
rect 4617 1984 4625 1986
rect 4678 1986 4725 1992
rect 4678 1984 4689 1986
rect 4717 1984 4725 1986
rect 4257 1938 4269 1944
rect 4301 1938 4313 1944
rect 4377 1938 4389 1944
rect 4511 1938 4523 1944
rect 4557 1938 4569 1944
rect 4597 1938 4609 1944
rect 4657 1938 4669 1944
rect 4697 1938 4709 1944
rect -62 1936 4776 1938
rect -62 1924 4 1936
rect -62 1922 4776 1924
rect -62 1458 -2 1922
rect 41 1916 53 1922
rect 107 1916 119 1922
rect 153 1916 165 1922
rect 211 1916 223 1922
rect 262 1916 274 1922
rect 312 1916 324 1922
rect 77 1870 85 1876
rect 127 1870 139 1876
rect 67 1856 85 1870
rect 113 1858 135 1870
rect 181 1862 193 1896
rect 77 1850 85 1856
rect 77 1842 115 1850
rect 133 1846 163 1852
rect 21 1828 83 1836
rect 21 1744 27 1828
rect 133 1832 139 1846
rect 181 1838 187 1856
rect 95 1826 139 1832
rect 147 1832 187 1838
rect 66 1787 93 1794
rect 40 1776 46 1781
rect 40 1768 74 1776
rect 79 1760 86 1768
rect 147 1760 153 1832
rect 376 1916 388 1922
rect 426 1916 438 1922
rect 337 1857 373 1863
rect 207 1824 221 1832
rect 213 1773 227 1787
rect 235 1773 243 1836
rect 293 1801 301 1836
rect 79 1754 153 1760
rect 227 1759 243 1773
rect 299 1765 307 1787
rect 337 1783 343 1857
rect 476 1916 488 1922
rect 526 1916 538 1922
rect 576 1916 588 1922
rect 626 1916 638 1922
rect 657 1916 669 1922
rect 717 1916 729 1922
rect 831 1916 843 1922
rect 399 1801 407 1836
rect 499 1801 507 1836
rect 599 1801 607 1836
rect 327 1777 343 1783
rect 393 1765 401 1787
rect 493 1765 501 1787
rect 593 1765 601 1787
rect 676 1793 684 1876
rect 736 1793 744 1876
rect 857 1916 869 1922
rect 897 1916 909 1922
rect 981 1916 993 1922
rect 1047 1916 1059 1922
rect 1093 1916 1105 1922
rect 1151 1916 1163 1922
rect 1197 1916 1209 1922
rect 1237 1916 1249 1922
rect 878 1874 889 1876
rect 917 1874 925 1876
rect 878 1868 925 1874
rect 803 1829 820 1836
rect 79 1748 86 1754
rect 147 1752 153 1754
rect 111 1736 132 1743
rect 235 1744 243 1759
rect 300 1758 325 1765
rect 60 1724 67 1730
rect 125 1724 132 1736
rect 182 1730 193 1738
rect 182 1724 189 1730
rect 60 1718 73 1724
rect 257 1744 309 1747
rect 269 1738 297 1744
rect 317 1744 325 1758
rect 375 1758 400 1765
rect 475 1758 500 1765
rect 575 1758 600 1765
rect 375 1744 383 1758
rect 391 1744 443 1747
rect 475 1744 483 1758
rect 403 1738 431 1744
rect 491 1744 543 1747
rect 575 1744 583 1758
rect 503 1738 531 1744
rect 591 1744 643 1747
rect 603 1738 631 1744
rect 676 1724 684 1779
rect 813 1781 820 1829
rect 918 1813 925 1868
rect 1017 1870 1025 1876
rect 1067 1870 1079 1876
rect 1007 1856 1025 1870
rect 1053 1858 1075 1870
rect 1121 1862 1133 1896
rect 1017 1850 1025 1856
rect 1017 1842 1055 1850
rect 1073 1846 1103 1852
rect 961 1828 1023 1836
rect 736 1724 744 1779
rect 916 1771 924 1799
rect 813 1724 820 1767
rect 41 1698 53 1704
rect 103 1698 115 1704
rect 151 1698 163 1704
rect 209 1698 221 1704
rect 277 1698 289 1704
rect 411 1698 423 1704
rect 511 1698 523 1704
rect 611 1698 623 1704
rect 657 1698 669 1704
rect 717 1698 729 1704
rect 791 1698 803 1704
rect 831 1698 843 1704
rect 894 1762 924 1771
rect 906 1760 924 1762
rect 961 1744 967 1828
rect 1073 1832 1079 1846
rect 1121 1838 1127 1856
rect 1035 1826 1079 1832
rect 1087 1832 1127 1838
rect 1006 1787 1033 1794
rect 980 1776 986 1781
rect 980 1768 1014 1776
rect 1019 1760 1026 1768
rect 1087 1760 1093 1832
rect 1296 1916 1308 1922
rect 1346 1916 1358 1922
rect 1147 1824 1161 1832
rect 1153 1773 1167 1787
rect 1175 1773 1183 1836
rect 1217 1821 1225 1876
rect 1391 1916 1403 1922
rect 1431 1916 1443 1922
rect 1471 1916 1483 1922
rect 1511 1916 1523 1922
rect 1551 1916 1563 1922
rect 1601 1916 1613 1922
rect 1667 1916 1679 1922
rect 1713 1916 1725 1922
rect 1771 1916 1783 1922
rect 1871 1916 1883 1922
rect 1917 1916 1929 1922
rect 2051 1916 2063 1922
rect 2151 1916 2163 1922
rect 2197 1916 2209 1922
rect 2297 1916 2309 1922
rect 2355 1916 2367 1922
rect 2401 1916 2413 1922
rect 2467 1916 2479 1922
rect 2541 1916 2553 1922
rect 2607 1916 2619 1922
rect 2653 1916 2665 1922
rect 2711 1916 2723 1922
rect 2781 1916 2793 1922
rect 2847 1916 2859 1922
rect 2893 1916 2905 1922
rect 2951 1916 2963 1922
rect 3031 1916 3043 1922
rect 1637 1870 1645 1876
rect 1687 1870 1699 1876
rect 1627 1856 1645 1870
rect 1673 1858 1695 1870
rect 1741 1862 1753 1896
rect 1637 1850 1645 1856
rect 1637 1842 1675 1850
rect 1693 1846 1723 1852
rect 1019 1754 1093 1760
rect 1167 1759 1183 1773
rect 1019 1748 1026 1754
rect 1087 1752 1093 1754
rect 1051 1736 1072 1743
rect 1175 1744 1183 1759
rect 1217 1758 1225 1807
rect 1319 1801 1327 1836
rect 1411 1830 1423 1836
rect 1451 1830 1463 1836
rect 1491 1830 1503 1836
rect 1531 1830 1543 1836
rect 1405 1822 1423 1830
rect 1438 1822 1463 1830
rect 1478 1822 1503 1830
rect 1517 1822 1543 1830
rect 1581 1828 1643 1836
rect 1313 1765 1321 1787
rect 1405 1793 1412 1822
rect 1407 1779 1412 1793
rect 1295 1758 1320 1765
rect 1405 1758 1412 1779
rect 1438 1776 1446 1822
rect 1478 1776 1486 1822
rect 1517 1776 1525 1822
rect 1430 1764 1446 1776
rect 1470 1764 1486 1776
rect 1510 1764 1525 1776
rect 1438 1758 1446 1764
rect 1478 1758 1486 1764
rect 1517 1758 1525 1764
rect 1217 1752 1241 1758
rect 1229 1744 1241 1752
rect 1295 1744 1303 1758
rect 1405 1751 1424 1758
rect 1406 1750 1424 1751
rect 1438 1750 1464 1758
rect 1478 1750 1503 1758
rect 1517 1750 1544 1758
rect 1000 1724 1007 1730
rect 1065 1724 1072 1736
rect 1122 1730 1133 1738
rect 1122 1724 1129 1730
rect 1000 1718 1013 1724
rect 1311 1744 1363 1747
rect 1412 1744 1424 1750
rect 1452 1744 1464 1750
rect 1491 1744 1503 1750
rect 1532 1744 1544 1750
rect 1581 1744 1587 1828
rect 1693 1832 1699 1846
rect 1741 1838 1747 1856
rect 1655 1826 1699 1832
rect 1707 1832 1747 1838
rect 1626 1787 1653 1794
rect 1600 1776 1606 1781
rect 1600 1768 1634 1776
rect 1639 1760 1646 1768
rect 1707 1760 1713 1832
rect 1891 1842 1903 1844
rect 1863 1836 1903 1842
rect 2071 1842 2083 1844
rect 2043 1836 2083 1842
rect 2177 1842 2189 1844
rect 2177 1836 2217 1842
rect 2327 1862 2339 1896
rect 2381 1870 2393 1876
rect 2435 1870 2443 1876
rect 2385 1858 2407 1870
rect 2435 1856 2453 1870
rect 2333 1838 2339 1856
rect 2357 1846 2387 1852
rect 2435 1850 2443 1856
rect 1767 1824 1781 1832
rect 1773 1773 1787 1787
rect 1795 1773 1803 1836
rect 1834 1801 1842 1836
rect 1940 1829 1957 1836
rect 1639 1754 1713 1760
rect 1787 1759 1803 1773
rect 1639 1748 1646 1754
rect 1707 1752 1713 1754
rect 1323 1738 1351 1744
rect 1671 1736 1692 1743
rect 1795 1744 1803 1759
rect 1620 1724 1627 1730
rect 1685 1724 1692 1736
rect 1742 1730 1753 1738
rect 1742 1724 1749 1730
rect 1620 1718 1633 1724
rect 1834 1744 1842 1787
rect 1940 1781 1947 1829
rect 2014 1801 2022 1836
rect 2123 1829 2140 1836
rect 1834 1733 1860 1744
rect 1940 1724 1947 1767
rect 2014 1744 2022 1787
rect 2133 1781 2140 1829
rect 2238 1801 2246 1836
rect 2014 1733 2040 1744
rect 858 1698 870 1704
rect 981 1698 993 1704
rect 1043 1698 1055 1704
rect 1091 1698 1103 1704
rect 1149 1698 1161 1704
rect 1199 1698 1211 1704
rect 1331 1698 1343 1704
rect 1391 1698 1403 1704
rect 1431 1698 1443 1704
rect 1471 1698 1483 1704
rect 1511 1698 1523 1704
rect 1551 1698 1563 1704
rect 1601 1698 1613 1704
rect 1663 1698 1675 1704
rect 1711 1698 1723 1704
rect 1769 1698 1781 1704
rect 1838 1698 1850 1704
rect 1888 1698 1900 1704
rect 1917 1698 1929 1704
rect 1957 1698 1969 1704
rect 2133 1724 2140 1767
rect 2238 1744 2246 1787
rect 2018 1698 2030 1704
rect 2068 1698 2080 1704
rect 2111 1698 2123 1704
rect 2151 1698 2163 1704
rect 2220 1733 2246 1744
rect 2277 1773 2285 1836
rect 2299 1824 2313 1832
rect 2333 1832 2373 1838
rect 2293 1773 2307 1787
rect 2277 1759 2293 1773
rect 2367 1760 2373 1832
rect 2381 1832 2387 1846
rect 2405 1842 2443 1850
rect 2381 1826 2425 1832
rect 2437 1828 2499 1836
rect 2427 1787 2454 1794
rect 2474 1776 2480 1781
rect 2446 1768 2480 1776
rect 2434 1760 2441 1768
rect 2277 1744 2285 1759
rect 2367 1754 2441 1760
rect 2367 1752 2373 1754
rect 2434 1748 2441 1754
rect 2327 1730 2338 1738
rect 2331 1724 2338 1730
rect 2388 1736 2409 1743
rect 2493 1744 2499 1828
rect 2388 1724 2395 1736
rect 2453 1724 2460 1730
rect 2447 1718 2460 1724
rect 2577 1870 2585 1876
rect 2627 1870 2639 1876
rect 2567 1856 2585 1870
rect 2613 1858 2635 1870
rect 2681 1862 2693 1896
rect 2577 1850 2585 1856
rect 2577 1842 2615 1850
rect 2633 1846 2663 1852
rect 2521 1828 2583 1836
rect 2521 1744 2527 1828
rect 2633 1832 2639 1846
rect 2681 1838 2687 1856
rect 2595 1826 2639 1832
rect 2647 1832 2687 1838
rect 2566 1787 2593 1794
rect 2540 1776 2546 1781
rect 2540 1768 2574 1776
rect 2579 1760 2586 1768
rect 2647 1760 2653 1832
rect 2707 1824 2721 1832
rect 2713 1773 2727 1787
rect 2735 1773 2743 1836
rect 2579 1754 2653 1760
rect 2727 1759 2743 1773
rect 2579 1748 2586 1754
rect 2647 1752 2653 1754
rect 2611 1736 2632 1743
rect 2735 1744 2743 1759
rect 2560 1724 2567 1730
rect 2625 1724 2632 1736
rect 2682 1730 2693 1738
rect 2682 1724 2689 1730
rect 2560 1718 2573 1724
rect 2817 1870 2825 1876
rect 2867 1870 2879 1876
rect 2807 1856 2825 1870
rect 2853 1858 2875 1870
rect 2921 1862 2933 1896
rect 2817 1850 2825 1856
rect 2817 1842 2855 1850
rect 2873 1846 2903 1852
rect 2761 1828 2823 1836
rect 2761 1744 2767 1828
rect 2873 1832 2879 1846
rect 2921 1838 2927 1856
rect 2835 1826 2879 1832
rect 2887 1832 2927 1838
rect 2806 1787 2833 1794
rect 2780 1776 2786 1781
rect 2780 1768 2814 1776
rect 2819 1760 2826 1768
rect 2887 1760 2893 1832
rect 3071 1916 3083 1922
rect 3111 1916 3123 1922
rect 3171 1916 3183 1922
rect 3217 1916 3229 1922
rect 3297 1916 3309 1922
rect 3407 1916 3419 1922
rect 3451 1916 3463 1922
rect 2947 1824 2961 1832
rect 2953 1773 2967 1787
rect 2975 1773 2983 1836
rect 3016 1801 3024 1836
rect 3095 1821 3103 1876
rect 3197 1842 3209 1844
rect 3197 1836 3237 1842
rect 3477 1916 3489 1922
rect 3611 1916 3623 1922
rect 3691 1916 3703 1922
rect 3771 1916 3783 1922
rect 3819 1916 3831 1922
rect 3877 1916 3889 1922
rect 3921 1916 3933 1922
rect 4051 1916 4063 1922
rect 4117 1916 4129 1922
rect 4217 1916 4229 1922
rect 4257 1916 4269 1922
rect 2819 1754 2893 1760
rect 2967 1759 2983 1773
rect 2819 1748 2826 1754
rect 2887 1752 2893 1754
rect 2851 1736 2872 1743
rect 2975 1744 2983 1759
rect 3016 1744 3024 1787
rect 3095 1758 3103 1807
rect 3156 1801 3164 1836
rect 3187 1817 3213 1823
rect 3258 1801 3266 1836
rect 3320 1829 3337 1836
rect 3079 1752 3103 1758
rect 3079 1744 3091 1752
rect 3156 1744 3164 1787
rect 3258 1744 3266 1787
rect 3320 1781 3327 1829
rect 3391 1801 3399 1836
rect 3391 1787 3393 1801
rect 2800 1724 2807 1730
rect 2865 1724 2872 1736
rect 2922 1730 2933 1738
rect 2922 1724 2929 1730
rect 2800 1718 2813 1724
rect 2180 1698 2192 1704
rect 2230 1698 2242 1704
rect 2299 1698 2311 1704
rect 2357 1698 2369 1704
rect 2405 1698 2417 1704
rect 2467 1698 2479 1704
rect 2541 1698 2553 1704
rect 2603 1698 2615 1704
rect 2651 1698 2663 1704
rect 2709 1698 2721 1704
rect 2781 1698 2793 1704
rect 2843 1698 2855 1704
rect 2891 1698 2903 1704
rect 2949 1698 2961 1704
rect 3031 1698 3043 1704
rect 3109 1698 3121 1704
rect 3171 1698 3183 1704
rect 3240 1733 3266 1744
rect 3320 1724 3327 1767
rect 3391 1744 3399 1787
rect 3434 1762 3442 1876
rect 3563 1910 3591 1916
rect 3603 1838 3631 1844
rect 3496 1801 3504 1836
rect 3572 1830 3584 1836
rect 3572 1824 3599 1830
rect 3593 1801 3599 1824
rect 3676 1801 3684 1836
rect 3743 1829 3760 1836
rect 3425 1754 3463 1762
rect 3451 1744 3463 1754
rect 3496 1744 3504 1787
rect 3600 1744 3607 1787
rect 3676 1744 3684 1787
rect 3753 1781 3760 1829
rect 3797 1830 3805 1876
rect 3797 1824 3823 1830
rect 3820 1818 3823 1824
rect 3391 1734 3401 1744
rect 3200 1698 3212 1704
rect 3250 1698 3262 1704
rect 3753 1724 3760 1767
rect 3820 1762 3827 1818
rect 3841 1801 3849 1836
rect 3847 1787 3849 1801
rect 3820 1756 3823 1762
rect 3801 1750 3823 1756
rect 3801 1724 3809 1750
rect 3841 1744 3849 1787
rect 3898 1762 3906 1876
rect 4003 1910 4031 1916
rect 4043 1838 4071 1844
rect 4109 1838 4137 1844
rect 4149 1910 4177 1916
rect 4297 1916 4309 1922
rect 4341 1916 4353 1922
rect 4417 1916 4429 1922
rect 4551 1916 4563 1922
rect 3941 1801 3949 1836
rect 4012 1830 4024 1836
rect 4156 1830 4168 1836
rect 4012 1824 4039 1830
rect 4033 1801 4039 1824
rect 4141 1824 4168 1830
rect 4141 1801 4147 1824
rect 4237 1821 4245 1876
rect 3947 1787 3949 1801
rect 3877 1754 3915 1762
rect 3877 1744 3889 1754
rect 3941 1744 3949 1787
rect 4040 1744 4047 1787
rect 4133 1744 4140 1787
rect 4237 1758 4245 1807
rect 4318 1762 4326 1876
rect 4409 1838 4437 1844
rect 4449 1910 4477 1916
rect 4582 1916 4594 1922
rect 4632 1916 4644 1922
rect 4361 1801 4369 1836
rect 4456 1830 4468 1836
rect 4441 1824 4468 1830
rect 4441 1801 4447 1824
rect 4367 1787 4369 1801
rect 4237 1752 4261 1758
rect 4249 1744 4261 1752
rect 3297 1698 3309 1704
rect 3337 1698 3349 1704
rect 3421 1698 3433 1704
rect 3477 1698 3489 1704
rect 3572 1698 3584 1704
rect 3628 1698 3640 1704
rect 3691 1698 3703 1704
rect 3939 1734 3949 1744
rect 3731 1698 3743 1704
rect 3771 1698 3783 1704
rect 3819 1698 3831 1704
rect 3907 1698 3919 1704
rect 4012 1698 4024 1704
rect 4068 1698 4080 1704
rect 4100 1698 4112 1704
rect 4156 1698 4168 1704
rect 4297 1754 4335 1762
rect 4297 1744 4309 1754
rect 4361 1744 4369 1787
rect 4433 1744 4440 1787
rect 4536 1793 4544 1876
rect 4677 1916 4689 1922
rect 4613 1801 4621 1836
rect 4359 1734 4369 1744
rect 4536 1724 4544 1779
rect 4696 1793 4704 1876
rect 4619 1765 4627 1787
rect 4657 1783 4663 1793
rect 4647 1777 4663 1783
rect 4620 1758 4645 1765
rect 4577 1744 4629 1747
rect 4589 1738 4617 1744
rect 4637 1744 4645 1758
rect 4696 1724 4704 1779
rect 4219 1698 4231 1704
rect 4327 1698 4339 1704
rect 4400 1698 4412 1704
rect 4456 1698 4468 1704
rect 4551 1698 4563 1704
rect 4597 1698 4609 1704
rect 4677 1698 4689 1704
rect 4782 1698 4842 2162
rect 4 1696 4842 1698
rect 4776 1684 4842 1696
rect 4 1682 4842 1684
rect 17 1676 29 1682
rect 57 1676 69 1682
rect 97 1676 109 1682
rect 137 1676 149 1682
rect 177 1676 189 1682
rect 231 1676 243 1682
rect 271 1676 283 1682
rect 329 1676 341 1682
rect 401 1676 413 1682
rect 463 1676 475 1682
rect 511 1676 523 1682
rect 569 1676 581 1682
rect 641 1676 653 1682
rect 703 1676 715 1682
rect 751 1676 763 1682
rect 809 1676 821 1682
rect 879 1676 891 1682
rect 937 1676 949 1682
rect 985 1676 997 1682
rect 1047 1676 1059 1682
rect 1149 1676 1161 1682
rect 1231 1676 1243 1682
rect 1299 1676 1311 1682
rect 1357 1676 1369 1682
rect 1405 1676 1417 1682
rect 1467 1676 1479 1682
rect 1541 1676 1553 1682
rect 1603 1676 1615 1682
rect 1651 1676 1663 1682
rect 1709 1676 1721 1682
rect 1778 1676 1790 1682
rect 1828 1676 1840 1682
rect 36 1630 48 1636
rect 77 1630 89 1636
rect 116 1630 128 1636
rect 156 1630 168 1636
rect 36 1622 63 1630
rect 77 1622 102 1630
rect 116 1622 142 1630
rect 156 1629 174 1630
rect 156 1622 175 1629
rect 55 1616 63 1622
rect 94 1616 102 1622
rect 134 1616 142 1622
rect 55 1604 70 1616
rect 94 1604 110 1616
rect 134 1604 150 1616
rect 55 1558 63 1604
rect 94 1558 102 1604
rect 134 1558 142 1604
rect 168 1601 175 1622
rect 253 1613 260 1656
rect 168 1587 173 1601
rect 168 1558 175 1587
rect 37 1550 63 1558
rect 77 1550 102 1558
rect 117 1550 142 1558
rect 157 1550 175 1558
rect 253 1551 260 1599
rect 311 1593 319 1636
rect 351 1630 359 1656
rect 337 1624 359 1630
rect 420 1656 433 1662
rect 420 1650 427 1656
rect 485 1644 492 1656
rect 337 1618 340 1624
rect 311 1579 313 1593
rect 37 1544 49 1550
rect 77 1544 89 1550
rect 117 1544 129 1550
rect 157 1544 169 1550
rect 243 1544 260 1551
rect 311 1544 319 1579
rect 333 1562 340 1618
rect 337 1556 340 1562
rect 337 1550 363 1556
rect 355 1504 363 1550
rect 381 1552 387 1636
rect 471 1637 492 1644
rect 542 1650 549 1656
rect 542 1642 553 1650
rect 439 1626 446 1632
rect 507 1626 513 1628
rect 439 1620 513 1626
rect 595 1621 603 1636
rect 439 1612 446 1620
rect 400 1604 434 1612
rect 400 1599 406 1604
rect 426 1586 453 1593
rect 381 1544 443 1552
rect 455 1548 499 1554
rect 437 1530 475 1538
rect 493 1534 499 1548
rect 507 1548 513 1620
rect 587 1607 603 1621
rect 573 1593 587 1607
rect 507 1542 547 1548
rect 567 1548 581 1556
rect 595 1544 603 1607
rect 437 1524 445 1530
rect 493 1528 523 1534
rect 541 1524 547 1542
rect 427 1510 445 1524
rect 473 1510 495 1522
rect 437 1504 445 1510
rect 487 1504 499 1510
rect 541 1484 553 1518
rect 660 1656 673 1662
rect 660 1650 667 1656
rect 725 1644 732 1656
rect 621 1552 627 1636
rect 711 1637 732 1644
rect 782 1650 789 1656
rect 782 1642 793 1650
rect 679 1626 686 1632
rect 747 1626 753 1628
rect 679 1620 753 1626
rect 835 1621 843 1636
rect 679 1612 686 1620
rect 640 1604 674 1612
rect 640 1599 646 1604
rect 666 1586 693 1593
rect 621 1544 683 1552
rect 695 1548 739 1554
rect 677 1530 715 1538
rect 733 1534 739 1548
rect 747 1548 753 1620
rect 827 1607 843 1621
rect 813 1593 827 1607
rect 747 1542 787 1548
rect 807 1548 821 1556
rect 835 1544 843 1607
rect 677 1524 685 1530
rect 733 1528 763 1534
rect 781 1524 787 1542
rect 667 1510 685 1524
rect 713 1510 735 1522
rect 677 1504 685 1510
rect 727 1504 739 1510
rect 781 1484 793 1518
rect 1027 1656 1040 1662
rect 911 1650 918 1656
rect 907 1642 918 1650
rect 968 1644 975 1656
rect 1033 1650 1040 1656
rect 857 1621 865 1636
rect 968 1637 989 1644
rect 947 1626 953 1628
rect 1014 1626 1021 1632
rect 857 1607 873 1621
rect 947 1620 1021 1626
rect 857 1544 865 1607
rect 873 1593 887 1607
rect 879 1548 893 1556
rect 947 1548 953 1620
rect 1014 1612 1021 1620
rect 1026 1604 1060 1612
rect 1054 1599 1060 1604
rect 1007 1586 1034 1593
rect 913 1542 953 1548
rect 961 1548 1005 1554
rect 913 1524 919 1542
rect 961 1534 967 1548
rect 1073 1552 1079 1636
rect 1119 1628 1131 1636
rect 1119 1622 1143 1628
rect 1135 1573 1143 1622
rect 1195 1622 1203 1636
rect 1223 1636 1251 1642
rect 1211 1633 1263 1636
rect 1447 1656 1460 1662
rect 1331 1650 1338 1656
rect 1327 1642 1338 1650
rect 1388 1644 1395 1656
rect 1453 1650 1460 1656
rect 1195 1615 1220 1622
rect 1277 1621 1285 1636
rect 1388 1637 1409 1644
rect 1367 1626 1373 1628
rect 1434 1626 1441 1632
rect 1213 1593 1221 1615
rect 1277 1607 1293 1621
rect 1367 1620 1441 1626
rect 1017 1544 1079 1552
rect 937 1528 967 1534
rect 985 1530 1023 1538
rect 1015 1524 1023 1530
rect 907 1484 919 1518
rect 965 1510 987 1522
rect 1015 1510 1033 1524
rect 961 1504 973 1510
rect 1015 1504 1023 1510
rect 1135 1504 1143 1559
rect 1219 1544 1227 1579
rect 1277 1544 1285 1607
rect 1293 1593 1307 1607
rect 1299 1548 1313 1556
rect 17 1458 29 1464
rect 57 1458 69 1464
rect 97 1458 109 1464
rect 137 1458 149 1464
rect 177 1458 189 1464
rect 271 1458 283 1464
rect 329 1458 341 1464
rect 401 1458 413 1464
rect 467 1458 479 1464
rect 513 1458 525 1464
rect 571 1458 583 1464
rect 641 1458 653 1464
rect 707 1458 719 1464
rect 753 1458 765 1464
rect 811 1458 823 1464
rect 877 1458 889 1464
rect 935 1458 947 1464
rect 981 1458 993 1464
rect 1047 1458 1059 1464
rect 1111 1458 1123 1464
rect 1151 1458 1163 1464
rect 1367 1548 1373 1620
rect 1434 1612 1441 1620
rect 1446 1604 1480 1612
rect 1474 1599 1480 1604
rect 1427 1586 1454 1593
rect 1333 1542 1373 1548
rect 1381 1548 1425 1554
rect 1333 1524 1339 1542
rect 1381 1534 1387 1548
rect 1493 1552 1499 1636
rect 1437 1544 1499 1552
rect 1357 1528 1387 1534
rect 1405 1530 1443 1538
rect 1435 1524 1443 1530
rect 1327 1484 1339 1518
rect 1385 1510 1407 1522
rect 1435 1510 1453 1524
rect 1381 1504 1393 1510
rect 1435 1504 1443 1510
rect 1560 1656 1573 1662
rect 1560 1650 1567 1656
rect 1625 1644 1632 1656
rect 1521 1552 1527 1636
rect 1611 1637 1632 1644
rect 1682 1650 1689 1656
rect 1682 1642 1693 1650
rect 1579 1626 1586 1632
rect 1647 1626 1653 1628
rect 1579 1620 1653 1626
rect 1735 1621 1743 1636
rect 1579 1612 1586 1620
rect 1540 1604 1574 1612
rect 1540 1599 1546 1604
rect 1566 1586 1593 1593
rect 1521 1544 1583 1552
rect 1595 1548 1639 1554
rect 1577 1530 1615 1538
rect 1633 1534 1639 1548
rect 1647 1548 1653 1620
rect 1727 1607 1743 1621
rect 1713 1593 1727 1607
rect 1647 1542 1687 1548
rect 1707 1548 1721 1556
rect 1735 1544 1743 1607
rect 1774 1636 1800 1647
rect 1857 1676 1869 1682
rect 1897 1676 1909 1682
rect 1961 1676 1973 1682
rect 2023 1676 2035 1682
rect 2071 1676 2083 1682
rect 2129 1676 2141 1682
rect 2191 1676 2203 1682
rect 2231 1676 2243 1682
rect 2309 1676 2321 1682
rect 2357 1676 2369 1682
rect 2459 1676 2471 1682
rect 2517 1676 2529 1682
rect 2565 1676 2577 1682
rect 2627 1676 2639 1682
rect 2701 1676 2713 1682
rect 2763 1676 2775 1682
rect 2811 1676 2823 1682
rect 2869 1676 2881 1682
rect 2917 1676 2929 1682
rect 2979 1676 2991 1682
rect 3109 1676 3121 1682
rect 3157 1676 3169 1682
rect 3239 1676 3251 1682
rect 3369 1676 3381 1682
rect 3451 1676 3463 1682
rect 3498 1676 3510 1682
rect 3671 1676 3683 1682
rect 3717 1676 3729 1682
rect 3778 1676 3790 1682
rect 3880 1676 3892 1682
rect 3930 1676 3942 1682
rect 3997 1676 4009 1682
rect 4129 1676 4141 1682
rect 1774 1593 1782 1636
rect 1880 1613 1887 1656
rect 1774 1544 1782 1579
rect 1880 1551 1887 1599
rect 1980 1656 1993 1662
rect 1980 1650 1987 1656
rect 2045 1644 2052 1656
rect 1941 1552 1947 1636
rect 2031 1637 2052 1644
rect 2102 1650 2109 1656
rect 2102 1642 2113 1650
rect 1999 1626 2006 1632
rect 2067 1626 2073 1628
rect 1999 1620 2073 1626
rect 2155 1621 2163 1636
rect 1999 1612 2006 1620
rect 1960 1604 1994 1612
rect 1960 1599 1966 1604
rect 1986 1586 2013 1593
rect 1880 1544 1897 1551
rect 1577 1524 1585 1530
rect 1633 1528 1663 1534
rect 1681 1524 1687 1542
rect 1567 1510 1585 1524
rect 1613 1510 1635 1522
rect 1577 1504 1585 1510
rect 1627 1504 1639 1510
rect 1681 1484 1693 1518
rect 1803 1538 1843 1544
rect 1831 1536 1843 1538
rect 1941 1544 2003 1552
rect 2015 1548 2059 1554
rect 1997 1530 2035 1538
rect 2053 1534 2059 1548
rect 2067 1548 2073 1620
rect 2147 1607 2163 1621
rect 2133 1593 2147 1607
rect 2067 1542 2107 1548
rect 2127 1548 2141 1556
rect 2155 1544 2163 1607
rect 2213 1613 2220 1656
rect 2349 1636 2377 1642
rect 2279 1628 2291 1636
rect 2337 1633 2389 1636
rect 2607 1656 2620 1662
rect 2491 1650 2498 1656
rect 2487 1642 2498 1650
rect 2548 1644 2555 1656
rect 2613 1650 2620 1656
rect 2279 1622 2303 1628
rect 2397 1622 2405 1636
rect 2213 1551 2220 1599
rect 2295 1573 2303 1622
rect 2380 1615 2405 1622
rect 2437 1621 2445 1636
rect 2548 1637 2569 1644
rect 2527 1626 2533 1628
rect 2594 1626 2601 1632
rect 2379 1593 2387 1615
rect 2437 1607 2453 1621
rect 2527 1620 2601 1626
rect 1997 1524 2005 1530
rect 2053 1528 2083 1534
rect 2101 1524 2107 1542
rect 1987 1510 2005 1524
rect 2033 1510 2055 1522
rect 1997 1504 2005 1510
rect 2047 1504 2059 1510
rect 2101 1484 2113 1518
rect 2203 1544 2220 1551
rect 2295 1504 2303 1559
rect 2373 1544 2381 1579
rect 2437 1544 2445 1607
rect 2453 1593 2467 1607
rect 2459 1548 2473 1556
rect 1196 1458 1208 1464
rect 1246 1458 1258 1464
rect 1297 1458 1309 1464
rect 1355 1458 1367 1464
rect 1401 1458 1413 1464
rect 1467 1458 1479 1464
rect 1541 1458 1553 1464
rect 1607 1458 1619 1464
rect 1653 1458 1665 1464
rect 1711 1458 1723 1464
rect 1811 1458 1823 1464
rect 1857 1458 1869 1464
rect 1961 1458 1973 1464
rect 2027 1458 2039 1464
rect 2073 1458 2085 1464
rect 2131 1458 2143 1464
rect 2231 1458 2243 1464
rect 2271 1458 2283 1464
rect 2311 1458 2323 1464
rect 2527 1548 2533 1620
rect 2594 1612 2601 1620
rect 2606 1604 2640 1612
rect 2634 1599 2640 1604
rect 2587 1586 2614 1593
rect 2493 1542 2533 1548
rect 2541 1548 2585 1554
rect 2493 1524 2499 1542
rect 2541 1534 2547 1548
rect 2653 1552 2659 1636
rect 2597 1544 2659 1552
rect 2517 1528 2547 1534
rect 2565 1530 2603 1538
rect 2595 1524 2603 1530
rect 2487 1484 2499 1518
rect 2545 1510 2567 1522
rect 2595 1510 2613 1524
rect 2541 1504 2553 1510
rect 2595 1504 2603 1510
rect 2720 1656 2733 1662
rect 2720 1650 2727 1656
rect 2785 1644 2792 1656
rect 2681 1552 2687 1636
rect 2771 1637 2792 1644
rect 2842 1650 2849 1656
rect 2842 1642 2853 1650
rect 2739 1626 2746 1632
rect 2807 1626 2813 1628
rect 2739 1620 2813 1626
rect 2895 1621 2903 1636
rect 2739 1612 2746 1620
rect 2700 1604 2734 1612
rect 2700 1599 2706 1604
rect 2726 1586 2753 1593
rect 2681 1544 2743 1552
rect 2755 1548 2799 1554
rect 2737 1530 2775 1538
rect 2793 1534 2799 1548
rect 2807 1548 2813 1620
rect 2887 1607 2903 1621
rect 2873 1593 2887 1607
rect 2807 1542 2847 1548
rect 2867 1548 2881 1556
rect 2895 1544 2903 1607
rect 2936 1593 2944 1636
rect 3009 1628 3021 1636
rect 2997 1622 3021 1628
rect 3149 1636 3177 1642
rect 3079 1628 3091 1636
rect 3137 1633 3189 1636
rect 3079 1622 3103 1628
rect 3197 1622 3205 1636
rect 3269 1628 3281 1636
rect 2936 1544 2944 1579
rect 2997 1573 3005 1622
rect 3095 1573 3103 1622
rect 3180 1615 3205 1622
rect 3257 1622 3281 1628
rect 3339 1628 3351 1636
rect 3179 1593 3187 1615
rect 2737 1524 2745 1530
rect 2793 1528 2823 1534
rect 2841 1524 2847 1542
rect 2727 1510 2745 1524
rect 2773 1510 2795 1522
rect 2737 1504 2745 1510
rect 2787 1504 2799 1510
rect 2841 1484 2853 1518
rect 2997 1504 3005 1559
rect 3095 1504 3103 1559
rect 3173 1544 3181 1579
rect 3257 1573 3265 1622
rect 3339 1622 3363 1628
rect 2342 1458 2354 1464
rect 2392 1458 2404 1464
rect 2457 1458 2469 1464
rect 2515 1458 2527 1464
rect 2561 1458 2573 1464
rect 2627 1458 2639 1464
rect 2701 1458 2713 1464
rect 2767 1458 2779 1464
rect 2813 1458 2825 1464
rect 2871 1458 2883 1464
rect 2917 1458 2929 1464
rect 2977 1458 2989 1464
rect 3017 1458 3029 1464
rect 3071 1458 3083 1464
rect 3111 1458 3123 1464
rect 3257 1504 3265 1559
rect 3317 1543 3323 1613
rect 3355 1573 3363 1622
rect 3387 1617 3403 1623
rect 3317 1537 3333 1543
rect 3355 1504 3363 1559
rect 3397 1527 3403 1617
rect 3415 1622 3423 1636
rect 3443 1636 3471 1642
rect 3431 1633 3483 1636
rect 3415 1615 3440 1622
rect 3623 1670 3651 1676
rect 3663 1636 3691 1640
rect 3635 1626 3641 1636
rect 3651 1634 3703 1636
rect 3546 1618 3564 1620
rect 3635 1619 3664 1626
rect 3433 1593 3441 1615
rect 3534 1609 3564 1618
rect 3556 1581 3564 1609
rect 3439 1544 3447 1579
rect 3656 1593 3664 1619
rect 3736 1601 3744 1656
rect 3920 1636 3946 1647
rect 3826 1618 3844 1620
rect 3814 1609 3844 1618
rect 3142 1458 3154 1464
rect 3192 1458 3204 1464
rect 3237 1458 3249 1464
rect 3277 1458 3289 1464
rect 3331 1458 3343 1464
rect 3371 1458 3383 1464
rect 3558 1512 3565 1567
rect 3655 1544 3663 1579
rect 3518 1506 3565 1512
rect 3518 1504 3529 1506
rect 3416 1458 3428 1464
rect 3466 1458 3478 1464
rect 3557 1504 3565 1506
rect 3736 1504 3744 1587
rect 3836 1581 3844 1609
rect 3938 1593 3946 1636
rect 3989 1636 4017 1642
rect 3977 1633 4029 1636
rect 4160 1676 4172 1682
rect 4210 1676 4222 1682
rect 4277 1676 4289 1682
rect 4357 1676 4369 1682
rect 4417 1676 4429 1682
rect 4457 1676 4469 1682
rect 4200 1636 4226 1647
rect 4037 1622 4045 1636
rect 4099 1628 4111 1636
rect 4099 1622 4123 1628
rect 4020 1615 4045 1622
rect 4019 1593 4027 1615
rect 3838 1512 3845 1567
rect 3938 1544 3946 1579
rect 4013 1544 4021 1579
rect 4115 1573 4123 1622
rect 4218 1593 4226 1636
rect 4269 1636 4297 1642
rect 4257 1633 4309 1636
rect 4499 1676 4511 1682
rect 4579 1676 4591 1682
rect 4659 1676 4671 1682
rect 4317 1622 4325 1636
rect 4300 1615 4325 1622
rect 4299 1593 4307 1615
rect 4376 1601 4384 1656
rect 4440 1613 4447 1656
rect 4529 1628 4541 1636
rect 4609 1628 4621 1636
rect 4689 1628 4701 1636
rect 3798 1506 3845 1512
rect 3798 1504 3809 1506
rect 3497 1458 3509 1464
rect 3537 1458 3549 1464
rect 3621 1458 3633 1464
rect 3691 1458 3703 1464
rect 3837 1504 3845 1506
rect 3877 1538 3917 1544
rect 3877 1536 3889 1538
rect 4115 1504 4123 1559
rect 4218 1544 4226 1579
rect 4293 1544 4301 1579
rect 4157 1538 4197 1544
rect 4157 1536 4169 1538
rect 3717 1458 3729 1464
rect 3777 1458 3789 1464
rect 3817 1458 3829 1464
rect 3897 1458 3909 1464
rect 3982 1458 3994 1464
rect 4032 1458 4044 1464
rect 4376 1504 4384 1587
rect 4440 1551 4447 1599
rect 4517 1622 4541 1628
rect 4597 1622 4621 1628
rect 4517 1573 4525 1622
rect 4597 1573 4605 1622
rect 4677 1622 4701 1628
rect 4440 1544 4457 1551
rect 4091 1458 4103 1464
rect 4131 1458 4143 1464
rect 4177 1458 4189 1464
rect 4262 1458 4274 1464
rect 4312 1458 4324 1464
rect 4517 1504 4525 1559
rect 4597 1504 4605 1559
rect 4637 1543 4643 1613
rect 4677 1573 4685 1622
rect 4627 1537 4643 1543
rect 4677 1504 4685 1559
rect 4357 1458 4369 1464
rect 4417 1458 4429 1464
rect 4497 1458 4509 1464
rect 4537 1458 4549 1464
rect 4577 1458 4589 1464
rect 4617 1458 4629 1464
rect 4657 1458 4669 1464
rect 4697 1458 4709 1464
rect -62 1456 4776 1458
rect -62 1444 4 1456
rect -62 1442 4776 1444
rect -62 978 -2 1442
rect 37 1436 49 1442
rect 95 1436 107 1442
rect 141 1436 153 1442
rect 207 1436 219 1442
rect 281 1436 293 1442
rect 347 1436 359 1442
rect 393 1436 405 1442
rect 451 1436 463 1442
rect 497 1436 509 1442
rect 537 1436 549 1442
rect 67 1382 79 1416
rect 121 1390 133 1396
rect 175 1390 183 1396
rect 125 1378 147 1390
rect 175 1376 193 1390
rect 73 1358 79 1376
rect 97 1366 127 1372
rect 175 1370 183 1376
rect 17 1293 25 1356
rect 39 1344 53 1352
rect 73 1352 113 1358
rect 33 1293 47 1307
rect 17 1279 33 1293
rect 107 1280 113 1352
rect 121 1352 127 1366
rect 145 1362 183 1370
rect 121 1346 165 1352
rect 177 1348 239 1356
rect 167 1307 194 1314
rect 214 1296 220 1301
rect 186 1288 220 1296
rect 174 1280 181 1288
rect 17 1264 25 1279
rect 107 1274 181 1280
rect 107 1272 113 1274
rect 174 1268 181 1274
rect 67 1250 78 1258
rect 71 1244 78 1250
rect 128 1256 149 1263
rect 233 1264 239 1348
rect 128 1244 135 1256
rect 193 1244 200 1250
rect 187 1238 200 1244
rect 317 1390 325 1396
rect 367 1390 379 1396
rect 307 1376 325 1390
rect 353 1378 375 1390
rect 421 1382 433 1416
rect 317 1370 325 1376
rect 317 1362 355 1370
rect 373 1366 403 1372
rect 261 1348 323 1356
rect 261 1264 267 1348
rect 373 1352 379 1366
rect 421 1358 427 1376
rect 335 1346 379 1352
rect 387 1352 427 1358
rect 306 1307 333 1314
rect 280 1296 286 1301
rect 280 1288 314 1296
rect 319 1280 326 1288
rect 387 1280 393 1352
rect 596 1436 608 1442
rect 646 1436 658 1442
rect 447 1344 461 1352
rect 453 1293 467 1307
rect 475 1293 483 1356
rect 517 1341 525 1396
rect 696 1436 708 1442
rect 746 1436 758 1442
rect 809 1436 821 1442
rect 857 1436 869 1442
rect 897 1436 909 1442
rect 956 1436 968 1442
rect 1006 1436 1018 1442
rect 1071 1436 1083 1442
rect 319 1274 393 1280
rect 467 1279 483 1293
rect 319 1268 326 1274
rect 387 1272 393 1274
rect 351 1256 372 1263
rect 475 1264 483 1279
rect 517 1278 525 1327
rect 619 1321 627 1356
rect 719 1321 727 1356
rect 791 1321 799 1356
rect 835 1350 843 1396
rect 817 1344 843 1350
rect 817 1338 820 1344
rect 877 1341 885 1396
rect 1097 1436 1109 1442
rect 1137 1436 1149 1442
rect 1177 1436 1189 1442
rect 613 1285 621 1307
rect 713 1285 721 1307
rect 791 1307 793 1321
rect 595 1278 620 1285
rect 695 1278 720 1285
rect 517 1272 541 1278
rect 529 1264 541 1272
rect 595 1264 603 1278
rect 300 1244 307 1250
rect 365 1244 372 1256
rect 422 1250 433 1258
rect 422 1244 429 1250
rect 300 1238 313 1244
rect 611 1264 663 1267
rect 695 1264 703 1278
rect 623 1258 651 1264
rect 711 1264 763 1267
rect 791 1264 799 1307
rect 813 1282 820 1338
rect 817 1276 820 1282
rect 877 1278 885 1327
rect 979 1321 987 1356
rect 973 1285 981 1307
rect 1056 1313 1064 1396
rect 1231 1436 1243 1442
rect 1271 1436 1283 1442
rect 1316 1436 1328 1442
rect 1366 1436 1378 1442
rect 1117 1350 1129 1356
rect 1157 1350 1165 1356
rect 1117 1344 1165 1350
rect 1157 1321 1165 1344
rect 1255 1341 1263 1396
rect 1411 1436 1423 1442
rect 1451 1436 1463 1442
rect 1496 1436 1508 1442
rect 1546 1436 1558 1442
rect 1599 1436 1611 1442
rect 1657 1436 1669 1442
rect 1697 1436 1709 1442
rect 955 1278 980 1285
rect 817 1270 839 1276
rect 877 1272 901 1278
rect 723 1258 751 1264
rect 831 1244 839 1270
rect 889 1264 901 1272
rect 955 1264 963 1278
rect 971 1264 1023 1267
rect 983 1258 1011 1264
rect 1056 1244 1064 1299
rect 1157 1278 1165 1307
rect 1255 1278 1263 1327
rect 1339 1321 1347 1356
rect 1435 1341 1443 1396
rect 1333 1285 1341 1307
rect 1117 1270 1165 1278
rect 1117 1264 1125 1270
rect 1157 1264 1165 1270
rect 1239 1272 1263 1278
rect 1315 1278 1340 1285
rect 1435 1278 1443 1327
rect 1519 1321 1527 1356
rect 1577 1350 1585 1396
rect 1756 1436 1768 1442
rect 1806 1436 1818 1442
rect 1857 1436 1869 1442
rect 1915 1436 1927 1442
rect 1961 1436 1973 1442
rect 2027 1436 2039 1442
rect 2077 1436 2089 1442
rect 2142 1436 2154 1442
rect 2192 1436 2204 1442
rect 1577 1344 1603 1350
rect 1600 1338 1603 1344
rect 1513 1285 1521 1307
rect 1239 1264 1251 1272
rect 1315 1264 1323 1278
rect 1419 1272 1443 1278
rect 1495 1278 1520 1285
rect 1600 1282 1607 1338
rect 1621 1321 1629 1356
rect 1677 1341 1685 1396
rect 1887 1382 1899 1416
rect 1941 1390 1953 1396
rect 1995 1390 2003 1396
rect 1945 1378 1967 1390
rect 1995 1376 2013 1390
rect 1893 1358 1899 1376
rect 1917 1366 1947 1372
rect 1995 1370 2003 1376
rect 1627 1307 1629 1321
rect 39 1218 51 1224
rect 97 1218 109 1224
rect 145 1218 157 1224
rect 207 1218 219 1224
rect 281 1218 293 1224
rect 343 1218 355 1224
rect 391 1218 403 1224
rect 449 1218 461 1224
rect 499 1218 511 1224
rect 631 1218 643 1224
rect 731 1218 743 1224
rect 809 1218 821 1224
rect 859 1218 871 1224
rect 991 1218 1003 1224
rect 1071 1218 1083 1224
rect 1331 1264 1383 1267
rect 1343 1258 1371 1264
rect 1419 1264 1431 1272
rect 1495 1264 1503 1278
rect 1600 1276 1603 1282
rect 1581 1270 1603 1276
rect 1511 1264 1563 1267
rect 1523 1258 1551 1264
rect 1581 1244 1589 1270
rect 1621 1264 1629 1307
rect 1677 1278 1685 1327
rect 1779 1321 1787 1356
rect 1773 1285 1781 1307
rect 1837 1293 1845 1356
rect 1859 1344 1873 1352
rect 1893 1352 1933 1358
rect 1853 1293 1867 1307
rect 1755 1278 1780 1285
rect 1837 1279 1853 1293
rect 1927 1280 1933 1352
rect 1941 1352 1947 1366
rect 1965 1362 2003 1370
rect 1941 1346 1985 1352
rect 1997 1348 2059 1356
rect 1987 1307 2014 1314
rect 2034 1296 2040 1301
rect 2006 1288 2040 1296
rect 1994 1280 2001 1288
rect 1677 1272 1701 1278
rect 1689 1264 1701 1272
rect 1755 1264 1763 1278
rect 1771 1264 1823 1267
rect 1783 1258 1811 1264
rect 1837 1264 1845 1279
rect 1927 1274 2001 1280
rect 1927 1272 1933 1274
rect 1994 1268 2001 1274
rect 1887 1250 1898 1258
rect 1891 1244 1898 1250
rect 1948 1256 1969 1263
rect 2053 1264 2059 1348
rect 2096 1313 2104 1396
rect 2251 1436 2263 1442
rect 2291 1436 2303 1442
rect 2371 1436 2383 1442
rect 2431 1436 2443 1442
rect 2173 1321 2181 1356
rect 2275 1341 2283 1396
rect 2457 1436 2469 1442
rect 2557 1436 2569 1442
rect 2615 1436 2627 1442
rect 2661 1436 2673 1442
rect 2727 1436 2739 1442
rect 2777 1436 2789 1442
rect 2891 1436 2903 1442
rect 2343 1349 2360 1356
rect 1948 1244 1955 1256
rect 2013 1244 2020 1250
rect 2007 1238 2020 1244
rect 2096 1244 2104 1299
rect 2179 1285 2187 1307
rect 2180 1278 2205 1285
rect 2275 1278 2283 1327
rect 2137 1264 2189 1267
rect 2149 1258 2177 1264
rect 2197 1264 2205 1278
rect 2259 1272 2283 1278
rect 2353 1301 2360 1349
rect 2416 1313 2424 1396
rect 2480 1349 2497 1356
rect 2587 1382 2599 1416
rect 2641 1390 2653 1396
rect 2695 1390 2703 1396
rect 2645 1378 2667 1390
rect 2695 1376 2713 1390
rect 2593 1358 2599 1376
rect 2617 1366 2647 1372
rect 2695 1370 2703 1376
rect 2480 1301 2487 1349
rect 2259 1264 2271 1272
rect 2353 1244 2360 1287
rect 2416 1244 2424 1299
rect 2480 1244 2487 1287
rect 2537 1293 2545 1356
rect 2559 1344 2573 1352
rect 2593 1352 2633 1358
rect 2553 1293 2567 1307
rect 2537 1279 2553 1293
rect 2627 1280 2633 1352
rect 2641 1352 2647 1366
rect 2665 1362 2703 1370
rect 2922 1436 2934 1442
rect 2972 1436 2984 1442
rect 3022 1436 3034 1442
rect 3072 1436 3084 1442
rect 3122 1436 3134 1442
rect 3172 1436 3184 1442
rect 3217 1436 3229 1442
rect 3261 1436 3273 1442
rect 3371 1436 3383 1442
rect 2641 1346 2685 1352
rect 2697 1348 2759 1356
rect 2687 1307 2714 1314
rect 2734 1296 2740 1301
rect 2706 1288 2740 1296
rect 2694 1280 2701 1288
rect 2537 1264 2545 1279
rect 2627 1274 2701 1280
rect 2627 1272 2633 1274
rect 1097 1218 1109 1224
rect 1137 1218 1149 1224
rect 1177 1218 1189 1224
rect 1269 1218 1281 1224
rect 1351 1218 1363 1224
rect 1449 1218 1461 1224
rect 1531 1218 1543 1224
rect 1599 1218 1611 1224
rect 1659 1218 1671 1224
rect 1791 1218 1803 1224
rect 1859 1218 1871 1224
rect 1917 1218 1929 1224
rect 1965 1218 1977 1224
rect 2027 1218 2039 1224
rect 2077 1218 2089 1224
rect 2157 1218 2169 1224
rect 2289 1218 2301 1224
rect 2331 1218 2343 1224
rect 2371 1218 2383 1224
rect 2431 1218 2443 1224
rect 2694 1268 2701 1274
rect 2587 1250 2598 1258
rect 2591 1244 2598 1250
rect 2648 1256 2669 1263
rect 2753 1264 2759 1348
rect 2800 1349 2817 1356
rect 2800 1301 2807 1349
rect 2876 1321 2884 1356
rect 2953 1321 2961 1356
rect 3053 1321 3061 1356
rect 3153 1321 3161 1356
rect 2648 1244 2655 1256
rect 2713 1244 2720 1250
rect 2707 1238 2720 1244
rect 2800 1244 2807 1287
rect 2876 1264 2884 1307
rect 2959 1285 2967 1307
rect 3059 1285 3067 1307
rect 3159 1285 3167 1307
rect 2960 1278 2985 1285
rect 3060 1278 3085 1285
rect 3160 1278 3185 1285
rect 3238 1282 3246 1396
rect 3397 1436 3409 1442
rect 3437 1436 3449 1442
rect 3516 1436 3528 1442
rect 3566 1436 3578 1442
rect 3418 1394 3429 1396
rect 3457 1394 3465 1396
rect 3418 1388 3465 1394
rect 3281 1321 3289 1356
rect 3343 1349 3360 1356
rect 3287 1307 3289 1321
rect 2917 1264 2969 1267
rect 2929 1258 2957 1264
rect 2977 1264 2985 1278
rect 3017 1264 3069 1267
rect 3029 1258 3057 1264
rect 3077 1264 3085 1278
rect 3117 1264 3169 1267
rect 3129 1258 3157 1264
rect 3177 1264 3185 1278
rect 3217 1274 3255 1282
rect 3217 1264 3229 1274
rect 3281 1264 3289 1307
rect 3279 1254 3289 1264
rect 3353 1301 3360 1349
rect 3458 1333 3465 1388
rect 3602 1436 3614 1442
rect 3652 1436 3664 1442
rect 3711 1436 3723 1442
rect 3751 1436 3763 1442
rect 3791 1436 3803 1442
rect 3831 1436 3843 1442
rect 3857 1436 3869 1442
rect 3901 1436 3913 1442
rect 3976 1436 3988 1442
rect 4026 1436 4038 1442
rect 3539 1321 3547 1356
rect 3633 1321 3641 1356
rect 3735 1341 3743 1396
rect 3815 1341 3823 1396
rect 3456 1291 3464 1319
rect 3353 1244 3360 1287
rect 2457 1218 2469 1224
rect 2497 1218 2509 1224
rect 2559 1218 2571 1224
rect 2617 1218 2629 1224
rect 2665 1218 2677 1224
rect 2727 1218 2739 1224
rect 2777 1218 2789 1224
rect 2817 1218 2829 1224
rect 2891 1218 2903 1224
rect 2937 1218 2949 1224
rect 3037 1218 3049 1224
rect 3137 1218 3149 1224
rect 3247 1218 3259 1224
rect 3331 1218 3343 1224
rect 3371 1218 3383 1224
rect 3434 1282 3464 1291
rect 3533 1285 3541 1307
rect 3639 1285 3647 1307
rect 3446 1280 3464 1282
rect 3515 1278 3540 1285
rect 3640 1278 3665 1285
rect 3735 1278 3743 1327
rect 3815 1278 3823 1327
rect 3878 1282 3886 1396
rect 4057 1436 4069 1442
rect 4131 1436 4143 1442
rect 4171 1436 4183 1442
rect 4211 1436 4223 1442
rect 4251 1436 4263 1442
rect 4331 1436 4343 1442
rect 3921 1321 3929 1356
rect 3999 1321 4007 1356
rect 3927 1307 3929 1321
rect 3515 1264 3523 1278
rect 3531 1264 3583 1267
rect 3543 1258 3571 1264
rect 3597 1264 3649 1267
rect 3609 1258 3637 1264
rect 3657 1264 3665 1278
rect 3719 1272 3743 1278
rect 3799 1272 3823 1278
rect 3857 1274 3895 1282
rect 3719 1264 3731 1272
rect 3799 1264 3811 1272
rect 3857 1264 3869 1274
rect 3921 1264 3929 1307
rect 3993 1285 4001 1307
rect 4076 1313 4084 1396
rect 4155 1341 4163 1396
rect 4235 1341 4243 1396
rect 4376 1436 4388 1442
rect 4426 1436 4438 1442
rect 4303 1349 4320 1356
rect 3975 1278 4000 1285
rect 3975 1264 3983 1278
rect 3919 1254 3929 1264
rect 3991 1264 4043 1267
rect 4003 1258 4031 1264
rect 4076 1244 4084 1299
rect 4155 1278 4163 1327
rect 4235 1278 4243 1327
rect 4139 1272 4163 1278
rect 4219 1272 4243 1278
rect 4313 1301 4320 1349
rect 4139 1264 4151 1272
rect 4219 1264 4231 1272
rect 4313 1244 4320 1287
rect 4357 1283 4363 1373
rect 4462 1436 4474 1442
rect 4512 1436 4524 1442
rect 4611 1436 4623 1442
rect 4657 1436 4669 1442
rect 4697 1436 4709 1442
rect 4631 1362 4643 1364
rect 4603 1356 4643 1362
rect 4399 1321 4407 1356
rect 4493 1321 4501 1356
rect 4574 1321 4582 1356
rect 4677 1341 4685 1396
rect 4393 1285 4401 1307
rect 4499 1285 4507 1307
rect 4347 1277 4363 1283
rect 4375 1278 4400 1285
rect 4500 1278 4525 1285
rect 4375 1264 4383 1278
rect 3398 1218 3410 1224
rect 3551 1218 3563 1224
rect 3617 1218 3629 1224
rect 3749 1218 3761 1224
rect 3829 1218 3841 1224
rect 3887 1218 3899 1224
rect 4011 1218 4023 1224
rect 4057 1218 4069 1224
rect 4169 1218 4181 1224
rect 4249 1218 4261 1224
rect 4391 1264 4443 1267
rect 4403 1258 4431 1264
rect 4457 1264 4509 1267
rect 4469 1258 4497 1264
rect 4517 1264 4525 1278
rect 4574 1264 4582 1307
rect 4677 1278 4685 1327
rect 4677 1272 4701 1278
rect 4689 1264 4701 1272
rect 4574 1253 4600 1264
rect 4291 1218 4303 1224
rect 4331 1218 4343 1224
rect 4411 1218 4423 1224
rect 4477 1218 4489 1224
rect 4578 1218 4590 1224
rect 4628 1218 4640 1224
rect 4659 1218 4671 1224
rect 4782 1218 4842 1682
rect 4 1216 4842 1218
rect 4776 1204 4842 1216
rect 4 1202 4842 1204
rect 17 1196 29 1202
rect 129 1196 141 1202
rect 211 1196 223 1202
rect 260 1196 272 1202
rect 316 1196 328 1202
rect 36 1121 44 1176
rect 99 1148 111 1156
rect 99 1142 123 1148
rect 36 1024 44 1107
rect 115 1093 123 1142
rect 175 1142 183 1156
rect 203 1156 231 1162
rect 398 1196 410 1202
rect 448 1196 460 1202
rect 511 1196 523 1202
rect 555 1196 563 1202
rect 394 1156 420 1167
rect 577 1196 589 1202
rect 617 1196 629 1202
rect 701 1196 713 1202
rect 789 1196 801 1202
rect 851 1196 863 1202
rect 891 1196 903 1202
rect 951 1196 963 1202
rect 1011 1196 1023 1202
rect 191 1153 243 1156
rect 175 1135 200 1142
rect 157 1117 173 1123
rect 115 1024 123 1079
rect 157 1043 163 1117
rect 193 1113 201 1135
rect 293 1113 300 1156
rect 394 1113 402 1156
rect 493 1121 500 1156
rect 531 1148 537 1176
rect 527 1142 537 1148
rect 199 1064 207 1099
rect 301 1076 307 1099
rect 301 1070 328 1076
rect 316 1064 328 1070
rect 394 1064 402 1099
rect 157 1037 173 1043
rect 17 978 29 984
rect 91 978 103 984
rect 131 978 143 984
rect 269 1056 297 1062
rect 309 984 337 990
rect 423 1058 463 1064
rect 451 1056 463 1058
rect 497 1063 506 1107
rect 516 1081 522 1136
rect 600 1133 607 1176
rect 527 1072 563 1080
rect 555 1064 563 1072
rect 600 1071 607 1119
rect 671 1156 681 1166
rect 1037 1196 1049 1202
rect 1077 1196 1089 1202
rect 1117 1196 1129 1202
rect 1191 1196 1203 1202
rect 1231 1196 1243 1202
rect 1260 1196 1272 1202
rect 1310 1196 1322 1202
rect 1381 1196 1393 1202
rect 1443 1196 1455 1202
rect 1491 1196 1503 1202
rect 1549 1196 1561 1202
rect 1631 1196 1643 1202
rect 671 1113 679 1156
rect 731 1146 743 1156
rect 705 1138 743 1146
rect 671 1099 673 1113
rect 600 1064 617 1071
rect 671 1064 679 1099
rect 497 1054 501 1063
rect 714 1024 722 1138
rect 771 1113 779 1156
rect 811 1150 819 1176
rect 797 1144 819 1150
rect 797 1138 800 1144
rect 771 1099 773 1113
rect 771 1064 779 1099
rect 793 1082 800 1138
rect 873 1133 880 1176
rect 936 1121 944 1176
rect 797 1076 800 1082
rect 797 1070 823 1076
rect 873 1071 880 1119
rect 996 1121 1004 1176
rect 1060 1133 1067 1176
rect 1136 1121 1144 1176
rect 1213 1133 1220 1176
rect 1300 1156 1326 1167
rect 815 1024 823 1070
rect 863 1064 880 1071
rect 936 1024 944 1107
rect 996 1024 1004 1107
rect 1060 1071 1067 1119
rect 1060 1064 1077 1071
rect 176 978 188 984
rect 226 978 238 984
rect 277 978 289 984
rect 431 978 443 984
rect 521 978 533 984
rect 577 978 589 984
rect 687 978 699 984
rect 731 978 743 984
rect 789 978 801 984
rect 891 978 903 984
rect 951 978 963 984
rect 1011 978 1023 984
rect 1136 1024 1144 1107
rect 1213 1071 1220 1119
rect 1318 1113 1326 1156
rect 1400 1176 1413 1182
rect 1400 1170 1407 1176
rect 1465 1164 1472 1176
rect 1203 1064 1220 1071
rect 1318 1064 1326 1099
rect 1361 1072 1367 1156
rect 1451 1157 1472 1164
rect 1522 1170 1529 1176
rect 1522 1162 1533 1170
rect 1419 1146 1426 1152
rect 1659 1196 1671 1202
rect 1737 1196 1749 1202
rect 1777 1196 1789 1202
rect 1841 1196 1853 1202
rect 1903 1196 1915 1202
rect 1951 1196 1963 1202
rect 2009 1196 2021 1202
rect 2091 1196 2103 1202
rect 1487 1146 1493 1148
rect 1419 1140 1493 1146
rect 1575 1141 1583 1156
rect 1419 1132 1426 1140
rect 1380 1124 1414 1132
rect 1380 1119 1386 1124
rect 1406 1106 1433 1113
rect 1361 1064 1423 1072
rect 1435 1068 1479 1074
rect 1257 1058 1297 1064
rect 1257 1056 1269 1058
rect 1417 1050 1455 1058
rect 1473 1054 1479 1068
rect 1487 1068 1493 1140
rect 1567 1127 1583 1141
rect 1553 1113 1567 1127
rect 1487 1062 1527 1068
rect 1547 1068 1561 1076
rect 1575 1064 1583 1127
rect 1616 1121 1624 1176
rect 1689 1148 1701 1156
rect 1677 1142 1701 1148
rect 1417 1044 1425 1050
rect 1473 1048 1503 1054
rect 1521 1044 1527 1062
rect 1407 1030 1425 1044
rect 1453 1030 1475 1042
rect 1417 1024 1425 1030
rect 1467 1024 1479 1030
rect 1521 1004 1533 1038
rect 1616 1024 1624 1107
rect 1677 1093 1685 1142
rect 1760 1133 1767 1176
rect 1677 1024 1685 1079
rect 1760 1071 1767 1119
rect 1860 1176 1873 1182
rect 1860 1170 1867 1176
rect 1925 1164 1932 1176
rect 1821 1072 1827 1156
rect 1911 1157 1932 1164
rect 1982 1170 1989 1176
rect 1982 1162 1993 1170
rect 1879 1146 1886 1152
rect 2117 1196 2129 1202
rect 2157 1196 2169 1202
rect 2197 1196 2209 1202
rect 2237 1196 2249 1202
rect 2311 1196 2323 1202
rect 2359 1196 2371 1202
rect 2417 1196 2429 1202
rect 2465 1196 2477 1202
rect 2527 1196 2539 1202
rect 2577 1196 2589 1202
rect 2657 1196 2669 1202
rect 2757 1196 2769 1202
rect 2857 1196 2869 1202
rect 2897 1196 2909 1202
rect 2989 1196 3001 1202
rect 3047 1196 3059 1202
rect 3137 1196 3149 1202
rect 3217 1196 3225 1202
rect 3257 1196 3269 1202
rect 3369 1196 3381 1202
rect 3449 1196 3461 1202
rect 1947 1146 1953 1148
rect 1879 1140 1953 1146
rect 2035 1141 2043 1156
rect 1879 1132 1886 1140
rect 1840 1124 1874 1132
rect 1840 1119 1846 1124
rect 1866 1106 1893 1113
rect 1760 1064 1777 1071
rect 1037 978 1049 984
rect 1117 978 1129 984
rect 1231 978 1243 984
rect 1277 978 1289 984
rect 1381 978 1393 984
rect 1447 978 1459 984
rect 1493 978 1505 984
rect 1551 978 1563 984
rect 1631 978 1643 984
rect 1657 978 1669 984
rect 1697 978 1709 984
rect 1821 1064 1883 1072
rect 1895 1068 1939 1074
rect 1877 1050 1915 1058
rect 1933 1054 1939 1068
rect 1947 1068 1953 1140
rect 2027 1127 2043 1141
rect 2013 1113 2027 1127
rect 1947 1062 1987 1068
rect 2007 1068 2021 1076
rect 2035 1064 2043 1127
rect 2076 1121 2084 1176
rect 2140 1133 2147 1176
rect 2220 1133 2227 1176
rect 2296 1121 2304 1176
rect 2507 1176 2520 1182
rect 2391 1170 2398 1176
rect 2387 1162 2398 1170
rect 2448 1164 2455 1176
rect 2513 1170 2520 1176
rect 2337 1141 2345 1156
rect 2448 1157 2469 1164
rect 2427 1146 2433 1148
rect 2494 1146 2501 1152
rect 1877 1044 1885 1050
rect 1933 1048 1963 1054
rect 1981 1044 1987 1062
rect 1867 1030 1885 1044
rect 1913 1030 1935 1042
rect 1877 1024 1885 1030
rect 1927 1024 1939 1030
rect 1981 1004 1993 1038
rect 2076 1024 2084 1107
rect 2140 1071 2147 1119
rect 2220 1071 2227 1119
rect 2337 1127 2353 1141
rect 2427 1140 2501 1146
rect 2140 1064 2157 1071
rect 2220 1064 2237 1071
rect 1737 978 1749 984
rect 1841 978 1853 984
rect 1907 978 1919 984
rect 1953 978 1965 984
rect 2011 978 2023 984
rect 2091 978 2103 984
rect 2296 1024 2304 1107
rect 2337 1064 2345 1127
rect 2353 1113 2367 1127
rect 2359 1068 2373 1076
rect 2427 1068 2433 1140
rect 2494 1132 2501 1140
rect 2506 1124 2540 1132
rect 2534 1119 2540 1124
rect 2487 1106 2514 1113
rect 2393 1062 2433 1068
rect 2441 1068 2485 1074
rect 2393 1044 2399 1062
rect 2441 1054 2447 1068
rect 2553 1072 2559 1156
rect 2596 1121 2604 1176
rect 2649 1156 2677 1162
rect 2637 1153 2689 1156
rect 2749 1156 2777 1160
rect 2789 1190 2817 1196
rect 2697 1142 2705 1156
rect 2737 1154 2789 1156
rect 2799 1146 2805 1156
rect 2680 1135 2705 1142
rect 2776 1139 2805 1146
rect 2497 1064 2559 1072
rect 2417 1048 2447 1054
rect 2465 1050 2503 1058
rect 2495 1044 2503 1050
rect 2387 1004 2399 1038
rect 2445 1030 2467 1042
rect 2495 1030 2513 1044
rect 2441 1024 2453 1030
rect 2495 1024 2503 1030
rect 2596 1024 2604 1107
rect 2679 1113 2687 1135
rect 2707 1117 2723 1123
rect 2673 1064 2681 1099
rect 2717 1067 2723 1117
rect 2776 1113 2784 1139
rect 2880 1133 2887 1176
rect 3079 1156 3089 1166
rect 2959 1148 2971 1156
rect 2959 1142 2983 1148
rect 2777 1064 2785 1099
rect 2880 1071 2887 1119
rect 2975 1093 2983 1142
rect 3017 1146 3029 1156
rect 3017 1138 3055 1146
rect 2880 1064 2897 1071
rect 2117 978 2129 984
rect 2197 978 2209 984
rect 2311 978 2323 984
rect 2357 978 2369 984
rect 2415 978 2427 984
rect 2461 978 2473 984
rect 2527 978 2539 984
rect 2577 978 2589 984
rect 2642 978 2654 984
rect 2692 978 2704 984
rect 2737 978 2749 984
rect 2807 978 2819 984
rect 2975 1024 2983 1079
rect 3038 1024 3046 1138
rect 3081 1113 3089 1156
rect 3129 1156 3157 1162
rect 3117 1153 3169 1156
rect 3177 1142 3185 1156
rect 3243 1148 3249 1176
rect 3479 1196 3491 1202
rect 3559 1196 3571 1202
rect 3657 1196 3669 1202
rect 3810 1196 3822 1202
rect 3243 1142 3253 1148
rect 3160 1135 3185 1142
rect 3087 1099 3089 1113
rect 3159 1113 3167 1135
rect 3187 1117 3203 1123
rect 3081 1064 3089 1099
rect 3153 1064 3161 1099
rect 2857 978 2869 984
rect 2951 978 2963 984
rect 2991 978 3003 984
rect 3197 1043 3203 1117
rect 3258 1081 3264 1136
rect 3280 1121 3287 1156
rect 3339 1148 3351 1156
rect 3419 1148 3431 1156
rect 3509 1148 3521 1156
rect 3589 1148 3601 1156
rect 3649 1156 3677 1162
rect 3637 1153 3689 1156
rect 3339 1142 3363 1148
rect 3419 1142 3443 1148
rect 3187 1037 3203 1043
rect 3217 1072 3253 1080
rect 3217 1064 3225 1072
rect 3274 1063 3283 1107
rect 3355 1093 3363 1142
rect 3435 1093 3443 1142
rect 3497 1142 3521 1148
rect 3497 1093 3505 1142
rect 3577 1142 3601 1148
rect 3697 1142 3705 1156
rect 3279 1054 3283 1063
rect 3355 1024 3363 1079
rect 3435 1024 3443 1079
rect 3497 1024 3505 1079
rect 3537 1063 3543 1133
rect 3577 1093 3585 1142
rect 3680 1135 3705 1142
rect 3756 1138 3774 1140
rect 3679 1113 3687 1135
rect 3756 1129 3786 1138
rect 3840 1196 3852 1202
rect 3890 1196 3902 1202
rect 3971 1196 3983 1202
rect 4070 1196 4082 1202
rect 3880 1156 3906 1167
rect 3756 1101 3764 1129
rect 3898 1113 3906 1156
rect 3956 1121 3964 1176
rect 4016 1138 4034 1140
rect 3527 1057 3543 1063
rect 3577 1024 3585 1079
rect 3673 1064 3681 1099
rect 4016 1129 4046 1138
rect 4100 1196 4112 1202
rect 4150 1196 4162 1202
rect 4197 1196 4209 1202
rect 4278 1196 4290 1202
rect 4328 1196 4340 1202
rect 4411 1196 4423 1202
rect 4477 1196 4489 1202
rect 4557 1196 4569 1202
rect 4597 1196 4609 1202
rect 4689 1196 4701 1202
rect 4751 1196 4763 1202
rect 4140 1156 4166 1167
rect 3017 978 3029 984
rect 3061 978 3073 984
rect 3122 978 3134 984
rect 3172 978 3184 984
rect 3247 978 3259 984
rect 3331 978 3343 984
rect 3371 978 3383 984
rect 3411 978 3423 984
rect 3451 978 3463 984
rect 3477 978 3489 984
rect 3517 978 3529 984
rect 3557 978 3569 984
rect 3597 978 3609 984
rect 3755 1032 3762 1087
rect 3898 1064 3906 1099
rect 3837 1058 3877 1064
rect 3837 1056 3849 1058
rect 3755 1026 3802 1032
rect 3755 1024 3763 1026
rect 3791 1024 3802 1026
rect 3956 1024 3964 1107
rect 4016 1101 4024 1129
rect 4158 1113 4166 1156
rect 4216 1121 4224 1176
rect 4274 1156 4300 1167
rect 4274 1113 4282 1156
rect 4375 1142 4383 1156
rect 4403 1156 4431 1162
rect 4391 1153 4443 1156
rect 4469 1156 4497 1162
rect 4457 1153 4509 1156
rect 4517 1142 4525 1156
rect 4375 1135 4400 1142
rect 4500 1135 4525 1142
rect 4015 1032 4022 1087
rect 4158 1064 4166 1099
rect 4097 1058 4137 1064
rect 4097 1056 4109 1058
rect 4015 1026 4062 1032
rect 4015 1024 4023 1026
rect 4051 1024 4062 1026
rect 4216 1024 4224 1107
rect 4393 1113 4401 1135
rect 4499 1113 4507 1135
rect 4580 1133 4587 1176
rect 4659 1148 4671 1156
rect 4659 1142 4683 1148
rect 4274 1064 4282 1099
rect 4399 1064 4407 1099
rect 4493 1064 4501 1099
rect 4580 1071 4587 1119
rect 4675 1093 4683 1142
rect 4707 1137 4723 1143
rect 4717 1087 4723 1137
rect 4736 1121 4744 1176
rect 4580 1064 4597 1071
rect 4303 1058 4343 1064
rect 4331 1056 4343 1058
rect 3642 978 3654 984
rect 3692 978 3704 984
rect 3771 978 3783 984
rect 3811 978 3823 984
rect 3857 978 3869 984
rect 3971 978 3983 984
rect 4031 978 4043 984
rect 4071 978 4083 984
rect 4117 978 4129 984
rect 4197 978 4209 984
rect 4311 978 4323 984
rect 4376 978 4388 984
rect 4426 978 4438 984
rect 4462 978 4474 984
rect 4512 978 4524 984
rect 4675 1024 4683 1079
rect 4736 1024 4744 1107
rect 4557 978 4569 984
rect 4651 978 4663 984
rect 4691 978 4703 984
rect 4751 978 4763 984
rect -62 976 4776 978
rect -62 964 4 976
rect -62 962 4776 964
rect -62 498 -2 962
rect 41 956 53 962
rect 107 956 119 962
rect 153 956 165 962
rect 211 956 223 962
rect 257 956 269 962
rect 297 956 309 962
rect 77 910 85 916
rect 127 910 139 916
rect 67 896 85 910
rect 113 898 135 910
rect 181 902 193 936
rect 77 890 85 896
rect 77 882 115 890
rect 133 886 163 892
rect 21 868 83 876
rect 21 784 27 868
rect 133 872 139 886
rect 181 878 187 896
rect 95 866 139 872
rect 147 872 187 878
rect 66 827 93 834
rect 40 816 46 821
rect 40 808 74 816
rect 79 800 86 808
rect 147 800 153 872
rect 356 956 368 962
rect 406 956 418 962
rect 461 956 473 962
rect 527 956 539 962
rect 573 956 585 962
rect 631 956 643 962
rect 677 956 689 962
rect 717 956 729 962
rect 207 864 221 872
rect 213 813 227 827
rect 235 813 243 876
rect 277 861 285 916
rect 497 910 505 916
rect 547 910 559 916
rect 487 896 505 910
rect 533 898 555 910
rect 601 902 613 936
rect 497 890 505 896
rect 497 882 535 890
rect 553 886 583 892
rect 79 794 153 800
rect 227 799 243 813
rect 79 788 86 794
rect 147 792 153 794
rect 111 776 132 783
rect 235 784 243 799
rect 277 798 285 847
rect 379 841 387 876
rect 441 868 503 876
rect 373 805 381 827
rect 355 798 380 805
rect 277 792 301 798
rect 289 784 301 792
rect 355 784 363 798
rect 60 764 67 770
rect 125 764 132 776
rect 182 770 193 778
rect 182 764 189 770
rect 60 758 73 764
rect 371 784 423 787
rect 383 778 411 784
rect 441 784 447 868
rect 553 872 559 886
rect 601 878 607 896
rect 515 866 559 872
rect 567 872 607 878
rect 486 827 513 834
rect 460 816 466 821
rect 460 808 494 816
rect 499 800 506 808
rect 567 800 573 872
rect 776 956 788 962
rect 826 956 838 962
rect 627 864 641 872
rect 633 813 647 827
rect 655 813 663 876
rect 697 861 705 916
rect 876 956 888 962
rect 926 956 938 962
rect 991 956 1003 962
rect 1071 956 1083 962
rect 499 794 573 800
rect 647 799 663 813
rect 499 788 506 794
rect 567 792 573 794
rect 531 776 552 783
rect 655 784 663 799
rect 697 798 705 847
rect 799 841 807 876
rect 899 841 907 876
rect 793 805 801 827
rect 893 805 901 827
rect 976 833 984 916
rect 1097 956 1109 962
rect 1191 956 1203 962
rect 1231 956 1243 962
rect 1271 956 1283 962
rect 1311 956 1323 962
rect 1351 956 1363 962
rect 1391 956 1403 962
rect 1471 956 1483 962
rect 1547 956 1559 962
rect 1591 956 1603 962
rect 1637 956 1649 962
rect 1717 956 1729 962
rect 1757 956 1769 962
rect 1797 956 1809 962
rect 1837 956 1849 962
rect 1877 956 1889 962
rect 1043 869 1060 876
rect 1053 821 1060 869
rect 1120 869 1137 876
rect 1120 821 1127 869
rect 1215 861 1223 916
rect 1295 861 1303 916
rect 1375 861 1383 916
rect 1491 882 1503 884
rect 1463 876 1503 882
rect 775 798 800 805
rect 875 798 900 805
rect 697 792 721 798
rect 709 784 721 792
rect 775 784 783 798
rect 480 764 487 770
rect 545 764 552 776
rect 602 770 613 778
rect 602 764 609 770
rect 480 758 493 764
rect 791 784 843 787
rect 875 784 883 798
rect 803 778 831 784
rect 891 784 943 787
rect 903 778 931 784
rect 976 764 984 819
rect 1053 764 1060 807
rect 1120 764 1127 807
rect 1215 798 1223 847
rect 1295 798 1303 847
rect 1375 798 1383 847
rect 1434 841 1442 876
rect 1531 841 1539 876
rect 1199 792 1223 798
rect 1279 792 1303 798
rect 1359 792 1383 798
rect 1199 784 1211 792
rect 1279 784 1291 792
rect 1359 784 1371 792
rect 1434 784 1442 827
rect 1531 827 1533 841
rect 1531 784 1539 827
rect 1574 802 1582 916
rect 1617 882 1629 884
rect 1617 876 1657 882
rect 1931 956 1943 962
rect 1971 956 1983 962
rect 2051 956 2063 962
rect 1678 841 1686 876
rect 1737 870 1749 876
rect 1777 870 1789 876
rect 1817 870 1829 876
rect 1857 870 1869 876
rect 1737 862 1763 870
rect 1777 862 1802 870
rect 1817 862 1842 870
rect 1857 862 1875 870
rect 1565 794 1603 802
rect 1591 784 1603 794
rect 1678 784 1686 827
rect 1755 816 1763 862
rect 1794 816 1802 862
rect 1834 816 1842 862
rect 1868 833 1875 862
rect 1955 861 1963 916
rect 2082 956 2094 962
rect 2132 956 2144 962
rect 2182 956 2194 962
rect 2232 956 2244 962
rect 2282 956 2294 962
rect 2332 956 2344 962
rect 2377 956 2389 962
rect 2417 956 2429 962
rect 2491 956 2503 962
rect 2537 956 2549 962
rect 2595 956 2607 962
rect 2641 956 2653 962
rect 2707 956 2719 962
rect 2776 956 2788 962
rect 2826 956 2838 962
rect 2891 956 2903 962
rect 2023 869 2040 876
rect 1868 819 1873 833
rect 1755 804 1770 816
rect 1794 804 1810 816
rect 1834 804 1850 816
rect 1755 798 1763 804
rect 1794 798 1802 804
rect 1834 798 1842 804
rect 1868 798 1875 819
rect 1955 798 1963 847
rect 1736 790 1763 798
rect 1777 790 1802 798
rect 1816 790 1842 798
rect 1856 791 1875 798
rect 1939 792 1963 798
rect 2033 821 2040 869
rect 2113 841 2121 876
rect 2213 841 2221 876
rect 2313 841 2321 876
rect 2397 861 2405 916
rect 1856 790 1874 791
rect 1736 784 1748 790
rect 1777 784 1789 790
rect 1816 784 1828 790
rect 1856 784 1868 790
rect 1939 784 1951 792
rect 41 738 53 744
rect 103 738 115 744
rect 151 738 163 744
rect 209 738 221 744
rect 259 738 271 744
rect 391 738 403 744
rect 461 738 473 744
rect 523 738 535 744
rect 571 738 583 744
rect 629 738 641 744
rect 679 738 691 744
rect 811 738 823 744
rect 911 738 923 744
rect 991 738 1003 744
rect 1031 738 1043 744
rect 1071 738 1083 744
rect 1434 773 1460 784
rect 1097 738 1109 744
rect 1137 738 1149 744
rect 1229 738 1241 744
rect 1309 738 1321 744
rect 1389 738 1401 744
rect 1531 774 1541 784
rect 1660 773 1686 784
rect 1438 738 1450 744
rect 1488 738 1500 744
rect 1561 738 1573 744
rect 1620 738 1632 744
rect 1670 738 1682 744
rect 2033 764 2040 807
rect 2119 805 2127 827
rect 2219 805 2227 827
rect 2319 805 2327 827
rect 2120 798 2145 805
rect 2220 798 2245 805
rect 2320 798 2345 805
rect 2077 784 2129 787
rect 1717 738 1729 744
rect 1757 738 1769 744
rect 1797 738 1809 744
rect 1837 738 1849 744
rect 1877 738 1889 744
rect 1969 738 1981 744
rect 2089 778 2117 784
rect 2137 784 2145 798
rect 2177 784 2229 787
rect 2189 778 2217 784
rect 2237 784 2245 798
rect 2277 784 2329 787
rect 2289 778 2317 784
rect 2337 784 2345 798
rect 2397 798 2405 847
rect 2476 833 2484 916
rect 2567 902 2579 936
rect 2621 910 2633 916
rect 2675 910 2683 916
rect 2625 898 2647 910
rect 2675 896 2693 910
rect 2573 878 2579 896
rect 2597 886 2627 892
rect 2675 890 2683 896
rect 2397 792 2421 798
rect 2409 784 2421 792
rect 2476 764 2484 819
rect 2517 813 2525 876
rect 2539 864 2553 872
rect 2573 872 2613 878
rect 2533 813 2547 827
rect 2517 799 2533 813
rect 2607 800 2613 872
rect 2621 872 2627 886
rect 2645 882 2683 890
rect 2917 956 2929 962
rect 2977 956 2989 962
rect 3017 956 3029 962
rect 3077 956 3089 962
rect 3151 956 3163 962
rect 3191 956 3203 962
rect 3247 956 3259 962
rect 3317 956 3329 962
rect 3357 956 3369 962
rect 2621 866 2665 872
rect 2677 868 2739 876
rect 2667 827 2694 834
rect 2714 816 2720 821
rect 2686 808 2720 816
rect 2674 800 2681 808
rect 2517 784 2525 799
rect 2607 794 2681 800
rect 2607 792 2613 794
rect 2674 788 2681 794
rect 2567 770 2578 778
rect 2571 764 2578 770
rect 2628 776 2649 783
rect 2733 784 2739 868
rect 2799 841 2807 876
rect 2793 805 2801 827
rect 2876 833 2884 916
rect 2936 833 2944 916
rect 2998 914 3009 916
rect 3037 914 3045 916
rect 2998 908 3045 914
rect 3038 853 3045 908
rect 2775 798 2800 805
rect 2775 784 2783 798
rect 2628 764 2635 776
rect 2693 764 2700 770
rect 2687 758 2700 764
rect 2791 784 2843 787
rect 2803 778 2831 784
rect 2876 764 2884 819
rect 2936 764 2944 819
rect 3036 811 3044 839
rect 3096 833 3104 916
rect 3175 861 3183 916
rect 3397 956 3409 962
rect 3437 956 3449 962
rect 3531 956 3543 962
rect 3279 877 3283 886
rect 3217 868 3225 876
rect 3217 860 3253 868
rect 2011 738 2023 744
rect 2051 738 2063 744
rect 2097 738 2109 744
rect 2197 738 2209 744
rect 2297 738 2309 744
rect 2379 738 2391 744
rect 2491 738 2503 744
rect 2539 738 2551 744
rect 2597 738 2609 744
rect 2645 738 2657 744
rect 2707 738 2719 744
rect 2811 738 2823 744
rect 2891 738 2903 744
rect 3014 802 3044 811
rect 3026 800 3044 802
rect 3096 764 3104 819
rect 3175 798 3183 847
rect 3258 804 3264 859
rect 3274 833 3283 877
rect 3159 792 3183 798
rect 3243 792 3253 798
rect 3159 784 3171 792
rect 3243 764 3249 792
rect 3280 784 3287 819
rect 3297 803 3303 893
rect 3337 861 3345 916
rect 3417 861 3425 916
rect 3557 956 3569 962
rect 3597 956 3609 962
rect 3671 956 3683 962
rect 3711 956 3723 962
rect 3771 956 3783 962
rect 3811 956 3823 962
rect 3503 869 3520 876
rect 3297 797 3313 803
rect 3337 798 3345 847
rect 3417 798 3425 847
rect 3513 821 3520 869
rect 3577 861 3585 916
rect 3655 914 3663 916
rect 3691 914 3702 916
rect 3655 908 3702 914
rect 3755 914 3763 916
rect 3837 956 3849 962
rect 3877 956 3889 962
rect 3951 956 3963 962
rect 3991 956 4003 962
rect 4051 956 4063 962
rect 3791 914 3802 916
rect 3755 908 3802 914
rect 3655 853 3662 908
rect 3337 792 3361 798
rect 3417 792 3441 798
rect 3349 784 3361 792
rect 3429 784 3441 792
rect 2917 738 2929 744
rect 2978 738 2990 744
rect 3077 738 3089 744
rect 3189 738 3201 744
rect 3513 764 3520 807
rect 3577 798 3585 847
rect 3755 853 3762 908
rect 3857 861 3865 916
rect 3935 914 3943 916
rect 4096 956 4108 962
rect 4146 956 4158 962
rect 3971 914 3982 916
rect 3935 908 3982 914
rect 3656 811 3664 839
rect 3756 811 3764 839
rect 3656 802 3686 811
rect 3656 800 3674 802
rect 3577 792 3601 798
rect 3589 784 3601 792
rect 3217 738 3225 744
rect 3257 738 3269 744
rect 3319 738 3331 744
rect 3399 738 3411 744
rect 3491 738 3503 744
rect 3531 738 3543 744
rect 3756 802 3786 811
rect 3756 800 3774 802
rect 3857 798 3865 847
rect 3857 792 3881 798
rect 3869 784 3881 792
rect 3559 738 3571 744
rect 3710 738 3722 744
rect 3810 738 3822 744
rect 3917 783 3923 873
rect 3935 853 3942 908
rect 4007 897 4023 903
rect 4017 847 4023 897
rect 3936 811 3944 839
rect 4036 833 4044 916
rect 4196 956 4208 962
rect 4246 956 4258 962
rect 4331 956 4343 962
rect 4377 956 4389 962
rect 4417 956 4429 962
rect 4511 956 4523 962
rect 4551 956 4563 962
rect 4631 956 4643 962
rect 4677 956 4689 962
rect 4717 956 4729 962
rect 4119 841 4127 876
rect 3936 802 3966 811
rect 3936 800 3954 802
rect 3917 777 3933 783
rect 4036 764 4044 819
rect 4113 805 4121 827
rect 4177 827 4183 893
rect 4398 914 4409 916
rect 4437 914 4445 916
rect 4398 908 4445 914
rect 4351 882 4363 884
rect 4323 876 4363 882
rect 4219 841 4227 876
rect 4213 805 4221 827
rect 4277 807 4283 853
rect 4294 841 4302 876
rect 4438 853 4445 908
rect 4495 914 4503 916
rect 4531 914 4542 916
rect 4495 908 4542 914
rect 4095 798 4120 805
rect 4195 798 4220 805
rect 4095 784 4103 798
rect 4111 784 4163 787
rect 4195 784 4203 798
rect 4123 778 4151 784
rect 4211 784 4263 787
rect 4223 778 4251 784
rect 4294 784 4302 827
rect 4436 811 4444 839
rect 4294 773 4320 784
rect 3839 738 3851 744
rect 3990 738 4002 744
rect 4051 738 4063 744
rect 4131 738 4143 744
rect 4231 738 4243 744
rect 4298 738 4310 744
rect 4348 738 4360 744
rect 4414 802 4444 811
rect 4477 807 4483 893
rect 4495 853 4502 908
rect 4698 914 4709 916
rect 4737 914 4745 916
rect 4698 908 4745 914
rect 4651 882 4663 884
rect 4623 876 4663 882
rect 4594 841 4602 876
rect 4738 853 4745 908
rect 4496 811 4504 839
rect 4426 800 4444 802
rect 4496 802 4526 811
rect 4496 800 4514 802
rect 4594 784 4602 827
rect 4736 811 4744 839
rect 4594 773 4620 784
rect 4378 738 4390 744
rect 4550 738 4562 744
rect 4598 738 4610 744
rect 4648 738 4660 744
rect 4714 802 4744 811
rect 4726 800 4744 802
rect 4678 738 4690 744
rect 4782 738 4842 1202
rect 4 736 4842 738
rect 4776 724 4842 736
rect 4 722 4842 724
rect 41 716 53 722
rect 103 716 115 722
rect 151 716 163 722
rect 209 716 221 722
rect 257 716 269 722
rect 337 716 349 722
rect 419 716 431 722
rect 519 716 531 722
rect 611 716 623 722
rect 659 716 671 722
rect 717 716 729 722
rect 765 716 777 722
rect 827 716 839 722
rect 897 716 909 722
rect 991 716 1003 722
rect 1031 716 1043 722
rect 60 696 73 702
rect 60 690 67 696
rect 125 684 132 696
rect 21 592 27 676
rect 111 677 132 684
rect 182 690 189 696
rect 182 682 193 690
rect 79 666 86 672
rect 147 666 153 668
rect 79 660 153 666
rect 235 661 243 676
rect 79 652 86 660
rect 40 644 74 652
rect 40 639 46 644
rect 66 626 93 633
rect 21 584 83 592
rect 95 588 139 594
rect 77 570 115 578
rect 133 574 139 588
rect 147 588 153 660
rect 227 647 243 661
rect 213 633 227 647
rect 147 582 187 588
rect 207 588 221 596
rect 235 584 243 647
rect 276 641 284 696
rect 329 676 357 682
rect 317 673 369 676
rect 377 662 385 676
rect 449 668 461 676
rect 360 655 385 662
rect 437 662 461 668
rect 501 670 509 696
rect 501 664 523 670
rect 77 564 85 570
rect 133 568 163 574
rect 181 564 187 582
rect 67 550 85 564
rect 113 550 135 562
rect 77 544 85 550
rect 127 544 139 550
rect 181 524 193 558
rect 276 544 284 627
rect 359 633 367 655
rect 353 584 361 619
rect 437 613 445 662
rect 520 658 523 664
rect 520 602 527 658
rect 541 633 549 676
rect 596 641 604 696
rect 807 696 820 702
rect 691 690 698 696
rect 687 682 698 690
rect 748 684 755 696
rect 813 690 820 696
rect 637 661 645 676
rect 748 677 769 684
rect 727 666 733 668
rect 794 666 801 672
rect 547 619 549 633
rect 637 647 653 661
rect 727 660 801 666
rect 437 544 445 599
rect 520 596 523 602
rect 497 590 523 596
rect 497 544 505 590
rect 541 584 549 619
rect 41 498 53 504
rect 107 498 119 504
rect 153 498 165 504
rect 211 498 223 504
rect 257 498 269 504
rect 322 498 334 504
rect 372 498 384 504
rect 596 544 604 627
rect 637 584 645 647
rect 653 633 667 647
rect 659 588 673 596
rect 727 588 733 660
rect 794 652 801 660
rect 806 644 840 652
rect 834 639 840 644
rect 787 626 814 633
rect 693 582 733 588
rect 741 588 785 594
rect 693 564 699 582
rect 741 574 747 588
rect 853 592 859 676
rect 889 676 917 682
rect 877 673 929 676
rect 1057 716 1065 722
rect 1097 716 1109 722
rect 1211 716 1223 722
rect 1301 716 1313 722
rect 1357 716 1369 722
rect 1397 716 1409 722
rect 1459 716 1471 722
rect 1541 716 1553 722
rect 1603 716 1615 722
rect 1651 716 1663 722
rect 1709 716 1721 722
rect 1779 716 1791 722
rect 1851 716 1863 722
rect 1891 716 1903 722
rect 937 662 945 676
rect 920 655 945 662
rect 919 633 927 655
rect 1013 653 1020 696
rect 1083 668 1089 696
rect 1083 662 1093 668
rect 797 584 859 592
rect 913 584 921 619
rect 1013 591 1020 639
rect 1098 601 1104 656
rect 1120 641 1127 676
rect 1175 662 1183 676
rect 1203 676 1231 682
rect 1191 673 1243 676
rect 1271 676 1281 686
rect 1175 655 1200 662
rect 1193 633 1201 655
rect 1003 584 1020 591
rect 1057 592 1093 600
rect 1057 584 1065 592
rect 717 568 747 574
rect 765 570 803 578
rect 795 564 803 570
rect 687 524 699 558
rect 745 550 767 562
rect 795 550 813 564
rect 741 544 753 550
rect 795 544 803 550
rect 1114 583 1123 627
rect 1271 633 1279 676
rect 1331 666 1343 676
rect 1305 658 1343 666
rect 1271 619 1273 633
rect 1199 584 1207 619
rect 1271 584 1279 619
rect 1119 574 1123 583
rect 1314 544 1322 658
rect 1380 653 1387 696
rect 1441 670 1449 696
rect 1560 696 1573 702
rect 1560 690 1567 696
rect 1625 684 1632 696
rect 1441 664 1463 670
rect 1380 591 1387 639
rect 1460 658 1463 664
rect 1460 602 1467 658
rect 1481 633 1489 676
rect 1487 619 1489 633
rect 1460 596 1463 602
rect 1380 584 1397 591
rect 417 498 429 504
rect 457 498 469 504
rect 519 498 531 504
rect 611 498 623 504
rect 657 498 669 504
rect 715 498 727 504
rect 761 498 773 504
rect 827 498 839 504
rect 882 498 894 504
rect 932 498 944 504
rect 1031 498 1043 504
rect 1087 498 1099 504
rect 1176 498 1188 504
rect 1226 498 1238 504
rect 1287 498 1299 504
rect 1331 498 1343 504
rect 1437 590 1463 596
rect 1437 544 1445 590
rect 1481 584 1489 619
rect 1521 592 1527 676
rect 1611 677 1632 684
rect 1682 690 1689 696
rect 1682 682 1693 690
rect 1579 666 1586 672
rect 1647 666 1653 668
rect 1579 660 1653 666
rect 1735 661 1743 676
rect 1761 670 1769 696
rect 1931 716 1943 722
rect 1971 716 1983 722
rect 2031 716 2043 722
rect 2057 716 2069 722
rect 2097 716 2109 722
rect 2159 716 2171 722
rect 2217 716 2229 722
rect 2265 716 2277 722
rect 2327 716 2339 722
rect 2380 716 2392 722
rect 2436 716 2448 722
rect 2531 716 2543 722
rect 2575 716 2583 722
rect 1761 664 1783 670
rect 1579 652 1586 660
rect 1540 644 1574 652
rect 1540 639 1546 644
rect 1566 626 1593 633
rect 1521 584 1583 592
rect 1595 588 1639 594
rect 1577 570 1615 578
rect 1633 574 1639 588
rect 1647 588 1653 660
rect 1727 647 1743 661
rect 1713 633 1727 647
rect 1647 582 1687 588
rect 1707 588 1721 596
rect 1735 584 1743 647
rect 1780 658 1783 664
rect 1780 602 1787 658
rect 1801 633 1809 676
rect 1873 653 1880 696
rect 1953 653 1960 696
rect 2016 641 2024 696
rect 2080 653 2087 696
rect 1807 619 1809 633
rect 1780 596 1783 602
rect 1577 564 1585 570
rect 1633 568 1663 574
rect 1681 564 1687 582
rect 1567 550 1585 564
rect 1613 550 1635 562
rect 1577 544 1585 550
rect 1627 544 1639 550
rect 1681 524 1693 558
rect 1757 590 1783 596
rect 1757 544 1765 590
rect 1801 584 1809 619
rect 1873 591 1880 639
rect 1953 591 1960 639
rect 1863 584 1880 591
rect 1943 584 1960 591
rect 2016 544 2024 627
rect 2080 591 2087 639
rect 2307 696 2320 702
rect 2191 690 2198 696
rect 2187 682 2198 690
rect 2248 684 2255 696
rect 2313 690 2320 696
rect 2137 661 2145 676
rect 2248 677 2269 684
rect 2618 716 2630 722
rect 2668 716 2680 722
rect 2227 666 2233 668
rect 2294 666 2301 672
rect 2137 647 2153 661
rect 2227 660 2301 666
rect 2080 584 2097 591
rect 1357 498 1369 504
rect 1459 498 1471 504
rect 1541 498 1553 504
rect 1607 498 1619 504
rect 1653 498 1665 504
rect 1711 498 1723 504
rect 1779 498 1791 504
rect 1891 498 1903 504
rect 1971 498 1983 504
rect 2031 498 2043 504
rect 2137 584 2145 647
rect 2153 633 2167 647
rect 2159 588 2173 596
rect 2227 588 2233 660
rect 2294 652 2301 660
rect 2306 644 2340 652
rect 2334 639 2340 644
rect 2287 626 2314 633
rect 2193 582 2233 588
rect 2241 588 2285 594
rect 2193 564 2199 582
rect 2241 574 2247 588
rect 2353 592 2359 676
rect 2413 633 2420 676
rect 2513 641 2520 676
rect 2551 668 2557 696
rect 2547 662 2557 668
rect 2614 676 2640 687
rect 2718 716 2730 722
rect 2768 716 2780 722
rect 2714 676 2740 687
rect 2797 716 2809 722
rect 2911 716 2923 722
rect 2977 716 2989 722
rect 3059 716 3071 722
rect 3171 716 3183 722
rect 2297 584 2359 592
rect 2421 596 2427 619
rect 2421 590 2448 596
rect 2436 584 2448 590
rect 2217 568 2247 574
rect 2265 570 2303 578
rect 2295 564 2303 570
rect 2187 524 2199 558
rect 2245 550 2267 562
rect 2295 550 2313 564
rect 2241 544 2253 550
rect 2295 544 2303 550
rect 2389 576 2417 582
rect 2429 504 2457 510
rect 2517 583 2526 627
rect 2536 601 2542 656
rect 2614 633 2622 676
rect 2714 633 2722 676
rect 2816 641 2824 696
rect 2875 662 2883 676
rect 2903 676 2931 682
rect 2891 673 2943 676
rect 2969 676 2997 682
rect 2957 673 3009 676
rect 3197 716 3209 722
rect 3330 716 3342 722
rect 3017 662 3025 676
rect 3089 668 3101 676
rect 2875 655 2900 662
rect 3000 655 3025 662
rect 3077 662 3101 668
rect 2893 633 2901 655
rect 2547 592 2583 600
rect 2575 584 2583 592
rect 2614 584 2622 619
rect 2714 584 2722 619
rect 2517 574 2521 583
rect 2643 578 2683 584
rect 2671 576 2683 578
rect 2743 578 2783 584
rect 2771 576 2783 578
rect 2816 544 2824 627
rect 2999 633 3007 655
rect 2899 584 2907 619
rect 2993 584 3001 619
rect 3077 613 3085 662
rect 3156 641 3164 696
rect 3216 641 3224 696
rect 3276 658 3294 660
rect 3276 649 3306 658
rect 3371 716 3383 722
rect 3411 716 3423 722
rect 3457 716 3469 722
rect 3540 716 3552 722
rect 3590 716 3602 722
rect 3393 653 3400 696
rect 3449 676 3477 682
rect 3437 673 3489 676
rect 3658 716 3670 722
rect 3708 716 3720 722
rect 3580 676 3606 687
rect 3497 662 3505 676
rect 3480 655 3505 662
rect 2057 498 2069 504
rect 2157 498 2169 504
rect 2215 498 2227 504
rect 2261 498 2273 504
rect 2327 498 2339 504
rect 2397 498 2409 504
rect 2541 498 2553 504
rect 2651 498 2663 504
rect 2751 498 2763 504
rect 2797 498 2809 504
rect 2876 498 2888 504
rect 2926 498 2938 504
rect 3077 544 3085 599
rect 3156 544 3164 627
rect 3216 544 3224 627
rect 3276 621 3284 649
rect 3275 552 3282 607
rect 3393 591 3400 639
rect 3479 633 3487 655
rect 3507 637 3523 643
rect 3383 584 3400 591
rect 3473 584 3481 619
rect 3517 603 3523 637
rect 3598 633 3606 676
rect 3654 676 3680 687
rect 3772 716 3784 722
rect 3828 716 3840 722
rect 3930 716 3942 722
rect 4030 716 4042 722
rect 3654 633 3662 676
rect 3800 633 3807 676
rect 3876 658 3894 660
rect 3876 649 3906 658
rect 3976 658 3994 660
rect 3976 649 4006 658
rect 4057 716 4069 722
rect 4118 716 4130 722
rect 4218 716 4230 722
rect 4390 716 4402 722
rect 4490 716 4502 722
rect 3876 621 3884 649
rect 3976 621 3984 649
rect 4076 641 4084 696
rect 4166 658 4184 660
rect 4154 649 4184 658
rect 4266 658 4284 660
rect 4254 649 4284 658
rect 3517 597 3553 603
rect 3598 584 3606 619
rect 3654 584 3662 619
rect 3793 596 3799 619
rect 3772 590 3799 596
rect 3772 584 3784 590
rect 3275 546 3322 552
rect 3275 544 3283 546
rect 2962 498 2974 504
rect 3012 498 3024 504
rect 3057 498 3069 504
rect 3097 498 3109 504
rect 3171 498 3183 504
rect 3311 544 3322 546
rect 3197 498 3209 504
rect 3291 498 3303 504
rect 3331 498 3343 504
rect 3411 498 3423 504
rect 3537 578 3577 584
rect 3537 576 3549 578
rect 3683 578 3723 584
rect 3711 576 3723 578
rect 3763 504 3791 510
rect 3803 576 3831 582
rect 3875 552 3882 607
rect 3975 552 3982 607
rect 3875 546 3922 552
rect 3875 544 3883 546
rect 3911 544 3922 546
rect 3975 546 4022 552
rect 3975 544 3983 546
rect 4011 544 4022 546
rect 4076 544 4084 627
rect 4176 621 4184 649
rect 4276 621 4284 649
rect 4336 658 4354 660
rect 4336 649 4366 658
rect 4436 658 4454 660
rect 4436 649 4466 658
rect 4517 716 4529 722
rect 4631 716 4643 722
rect 4697 716 4709 722
rect 4336 621 4344 649
rect 4436 621 4444 649
rect 4536 641 4544 696
rect 4595 662 4603 676
rect 4623 676 4651 682
rect 4611 673 4663 676
rect 4689 676 4717 682
rect 4677 673 4729 676
rect 4737 662 4745 676
rect 4595 655 4620 662
rect 4720 655 4745 662
rect 4613 633 4621 655
rect 4178 552 4185 607
rect 4278 552 4285 607
rect 4297 597 4313 603
rect 4297 587 4303 597
rect 4138 546 4185 552
rect 4138 544 4149 546
rect 3442 498 3454 504
rect 3492 498 3504 504
rect 3557 498 3569 504
rect 3691 498 3703 504
rect 3811 498 3823 504
rect 3891 498 3903 504
rect 3931 498 3943 504
rect 3991 498 4003 504
rect 4031 498 4043 504
rect 4177 544 4185 546
rect 4238 546 4285 552
rect 4238 544 4249 546
rect 4277 544 4285 546
rect 4335 552 4342 607
rect 4435 552 4442 607
rect 4335 546 4382 552
rect 4335 544 4343 546
rect 4371 544 4382 546
rect 4435 546 4482 552
rect 4435 544 4443 546
rect 4471 544 4482 546
rect 4536 544 4544 627
rect 4719 633 4727 655
rect 4619 584 4627 619
rect 4713 584 4721 619
rect 4057 498 4069 504
rect 4117 498 4129 504
rect 4157 498 4169 504
rect 4217 498 4229 504
rect 4257 498 4269 504
rect 4351 498 4363 504
rect 4391 498 4403 504
rect 4451 498 4463 504
rect 4491 498 4503 504
rect 4517 498 4529 504
rect 4596 498 4608 504
rect 4646 498 4658 504
rect 4682 498 4694 504
rect 4732 498 4744 504
rect -62 496 4776 498
rect -62 484 4 496
rect -62 482 4776 484
rect -62 18 -2 482
rect 41 476 53 482
rect 107 476 119 482
rect 153 476 165 482
rect 211 476 223 482
rect 257 476 269 482
rect 297 476 309 482
rect 77 430 85 436
rect 127 430 139 436
rect 67 416 85 430
rect 113 418 135 430
rect 181 422 193 456
rect 77 410 85 416
rect 77 402 115 410
rect 133 406 163 412
rect 21 388 83 396
rect 21 304 27 388
rect 133 392 139 406
rect 181 398 187 416
rect 95 386 139 392
rect 147 392 187 398
rect 66 347 93 354
rect 40 336 46 341
rect 40 328 74 336
rect 79 320 86 328
rect 147 320 153 392
rect 356 476 368 482
rect 406 476 418 482
rect 207 384 221 392
rect 213 333 227 347
rect 235 333 243 396
rect 277 381 285 436
rect 437 476 449 482
rect 497 476 509 482
rect 537 476 549 482
rect 596 476 608 482
rect 646 476 658 482
rect 79 314 153 320
rect 227 319 243 333
rect 79 308 86 314
rect 147 312 153 314
rect 111 296 132 303
rect 235 304 243 319
rect 277 318 285 367
rect 379 361 387 396
rect 373 325 381 347
rect 456 353 464 436
rect 517 381 525 436
rect 682 476 694 482
rect 732 476 744 482
rect 782 476 794 482
rect 832 476 844 482
rect 355 318 380 325
rect 277 312 301 318
rect 289 304 301 312
rect 355 304 363 318
rect 60 284 67 290
rect 125 284 132 296
rect 182 290 193 298
rect 182 284 189 290
rect 60 278 73 284
rect 371 304 423 307
rect 383 298 411 304
rect 456 284 464 339
rect 517 318 525 367
rect 619 361 627 396
rect 713 361 721 396
rect 896 476 908 482
rect 946 476 958 482
rect 977 476 989 482
rect 1037 476 1049 482
rect 1077 476 1089 482
rect 1171 476 1183 482
rect 1251 476 1263 482
rect 613 325 621 347
rect 719 325 727 347
rect 757 343 763 393
rect 813 361 821 396
rect 919 361 927 396
rect 747 337 763 343
rect 819 325 827 347
rect 913 325 921 347
rect 996 353 1004 436
rect 1057 381 1065 436
rect 1296 476 1308 482
rect 1346 476 1358 482
rect 1431 476 1443 482
rect 1191 402 1203 404
rect 1163 396 1203 402
rect 595 318 620 325
rect 720 318 745 325
rect 820 318 845 325
rect 517 312 541 318
rect 529 304 541 312
rect 595 304 603 318
rect 611 304 663 307
rect 623 298 651 304
rect 677 304 729 307
rect 689 298 717 304
rect 737 304 745 318
rect 777 304 829 307
rect 789 298 817 304
rect 837 304 845 318
rect 895 318 920 325
rect 895 304 903 318
rect 911 304 963 307
rect 923 298 951 304
rect 996 284 1004 339
rect 1057 318 1065 367
rect 1134 361 1142 396
rect 1236 353 1244 436
rect 1462 476 1474 482
rect 1512 476 1524 482
rect 1557 476 1569 482
rect 1597 476 1609 482
rect 1657 476 1669 482
rect 1715 476 1727 482
rect 1761 476 1773 482
rect 1827 476 1839 482
rect 1891 476 1903 482
rect 1931 476 1943 482
rect 1319 361 1327 396
rect 1403 389 1420 396
rect 1057 312 1081 318
rect 1069 304 1081 312
rect 1134 304 1142 347
rect 1134 293 1160 304
rect 1236 284 1244 339
rect 1313 325 1321 347
rect 1413 341 1420 389
rect 1493 361 1501 396
rect 1577 381 1585 436
rect 1687 422 1699 456
rect 1741 430 1753 436
rect 1795 430 1803 436
rect 1745 418 1767 430
rect 1795 416 1813 430
rect 1693 398 1699 416
rect 1717 406 1747 412
rect 1795 410 1803 416
rect 1295 318 1320 325
rect 1295 304 1303 318
rect 1311 304 1363 307
rect 1323 298 1351 304
rect 1413 284 1420 327
rect 1499 325 1507 347
rect 1500 318 1525 325
rect 1457 304 1509 307
rect 1469 298 1497 304
rect 1517 304 1525 318
rect 1577 318 1585 367
rect 1637 333 1645 396
rect 1659 384 1673 392
rect 1693 392 1733 398
rect 1653 333 1667 347
rect 1637 319 1653 333
rect 1727 320 1733 392
rect 1741 392 1747 406
rect 1765 402 1803 410
rect 1976 476 1988 482
rect 2026 476 2038 482
rect 2081 476 2093 482
rect 2147 476 2159 482
rect 2193 476 2205 482
rect 2251 476 2263 482
rect 2331 476 2343 482
rect 1741 386 1785 392
rect 1797 388 1859 396
rect 1787 347 1814 354
rect 1834 336 1840 341
rect 1806 328 1840 336
rect 1794 320 1801 328
rect 1577 312 1601 318
rect 1589 304 1601 312
rect 1637 304 1645 319
rect 1727 314 1801 320
rect 1727 312 1733 314
rect 1794 308 1801 314
rect 1687 290 1698 298
rect 1691 284 1698 290
rect 1748 296 1769 303
rect 1853 304 1859 388
rect 1915 381 1923 436
rect 2117 430 2125 436
rect 2167 430 2179 436
rect 2107 416 2125 430
rect 2153 418 2175 430
rect 2221 422 2233 456
rect 2117 410 2125 416
rect 2117 402 2155 410
rect 2173 406 2203 412
rect 1915 318 1923 367
rect 1999 361 2007 396
rect 2061 388 2123 396
rect 1993 325 2001 347
rect 1748 284 1755 296
rect 1813 284 1820 290
rect 1807 278 1820 284
rect 1899 312 1923 318
rect 1975 318 2000 325
rect 1899 304 1911 312
rect 1975 304 1983 318
rect 1991 304 2043 307
rect 2003 298 2031 304
rect 2061 304 2067 388
rect 2173 392 2179 406
rect 2221 398 2227 416
rect 2135 386 2179 392
rect 2187 392 2227 398
rect 2106 347 2133 354
rect 2080 336 2086 341
rect 2080 328 2114 336
rect 2119 320 2126 328
rect 2187 320 2193 392
rect 2357 476 2369 482
rect 2437 476 2449 482
rect 2511 476 2523 482
rect 2551 476 2563 482
rect 2597 476 2609 482
rect 2655 476 2667 482
rect 2701 476 2713 482
rect 2767 476 2779 482
rect 2817 476 2829 482
rect 2857 476 2869 482
rect 2917 476 2929 482
rect 3017 476 3029 482
rect 3097 476 3109 482
rect 3191 476 3203 482
rect 3231 476 3243 482
rect 3291 476 3303 482
rect 3331 476 3343 482
rect 2247 384 2261 392
rect 2253 333 2267 347
rect 2275 333 2283 396
rect 2316 353 2324 436
rect 2380 389 2397 396
rect 2380 341 2387 389
rect 2456 353 2464 436
rect 2535 381 2543 436
rect 2627 422 2639 456
rect 2681 430 2693 436
rect 2735 430 2743 436
rect 2685 418 2707 430
rect 2735 416 2753 430
rect 2633 398 2639 416
rect 2657 406 2687 412
rect 2735 410 2743 416
rect 2119 314 2193 320
rect 2267 319 2283 333
rect 2119 308 2126 314
rect 2187 312 2193 314
rect 2151 296 2172 303
rect 2275 304 2283 319
rect 2100 284 2107 290
rect 2165 284 2172 296
rect 2222 290 2233 298
rect 2222 284 2229 290
rect 2100 278 2113 284
rect 2316 284 2324 339
rect 2380 284 2387 327
rect 2456 284 2464 339
rect 2535 318 2543 367
rect 2519 312 2543 318
rect 2577 333 2585 396
rect 2599 384 2613 392
rect 2633 392 2673 398
rect 2593 333 2607 347
rect 2577 319 2593 333
rect 2667 320 2673 392
rect 2681 392 2687 406
rect 2705 402 2743 410
rect 2681 386 2725 392
rect 2737 388 2799 396
rect 2727 347 2754 354
rect 2774 336 2780 341
rect 2746 328 2780 336
rect 2734 320 2741 328
rect 2519 304 2531 312
rect 2577 304 2585 319
rect 2667 314 2741 320
rect 2667 312 2673 314
rect 41 258 53 264
rect 103 258 115 264
rect 151 258 163 264
rect 209 258 221 264
rect 259 258 271 264
rect 391 258 403 264
rect 437 258 449 264
rect 499 258 511 264
rect 631 258 643 264
rect 697 258 709 264
rect 797 258 809 264
rect 931 258 943 264
rect 977 258 989 264
rect 1039 258 1051 264
rect 1138 258 1150 264
rect 1188 258 1200 264
rect 1251 258 1263 264
rect 1331 258 1343 264
rect 1391 258 1403 264
rect 1431 258 1443 264
rect 1477 258 1489 264
rect 1559 258 1571 264
rect 1659 258 1671 264
rect 1717 258 1729 264
rect 1765 258 1777 264
rect 1827 258 1839 264
rect 1929 258 1941 264
rect 2011 258 2023 264
rect 2081 258 2093 264
rect 2143 258 2155 264
rect 2191 258 2203 264
rect 2249 258 2261 264
rect 2331 258 2343 264
rect 2357 258 2369 264
rect 2397 258 2409 264
rect 2734 308 2741 314
rect 2627 290 2638 298
rect 2631 284 2638 290
rect 2688 296 2709 303
rect 2793 304 2799 388
rect 2837 381 2845 436
rect 2909 398 2937 404
rect 2949 470 2977 476
rect 2956 390 2968 396
rect 2941 384 2968 390
rect 3040 389 3057 396
rect 2837 318 2845 367
rect 2941 361 2947 384
rect 2837 312 2861 318
rect 2849 304 2861 312
rect 2933 304 2940 347
rect 3040 341 3047 389
rect 3116 353 3124 436
rect 3175 434 3183 436
rect 3211 434 3222 436
rect 3175 428 3222 434
rect 3275 434 3283 436
rect 3362 476 3374 482
rect 3412 476 3424 482
rect 3491 476 3503 482
rect 3311 434 3322 436
rect 3275 428 3322 434
rect 3175 373 3182 428
rect 3275 373 3282 428
rect 3517 476 3529 482
rect 3557 476 3569 482
rect 3597 476 3609 482
rect 3637 476 3649 482
rect 3682 476 3694 482
rect 3732 476 3744 482
rect 3831 476 3843 482
rect 3911 476 3923 482
rect 3393 361 3401 396
rect 2688 284 2695 296
rect 2753 284 2760 290
rect 2747 278 2760 284
rect 3040 284 3047 327
rect 3116 284 3124 339
rect 3176 331 3184 359
rect 3276 331 3284 359
rect 3476 353 3484 436
rect 3537 381 3545 436
rect 3617 381 3625 436
rect 3647 397 3663 403
rect 3176 322 3206 331
rect 3176 320 3194 322
rect 2437 258 2449 264
rect 2549 258 2561 264
rect 2599 258 2611 264
rect 2657 258 2669 264
rect 2705 258 2717 264
rect 2767 258 2779 264
rect 2819 258 2831 264
rect 2900 258 2912 264
rect 2956 258 2968 264
rect 3017 258 3029 264
rect 3057 258 3069 264
rect 3276 322 3306 331
rect 3399 325 3407 347
rect 3276 320 3294 322
rect 3400 318 3425 325
rect 3357 304 3409 307
rect 3369 298 3397 304
rect 3417 304 3425 318
rect 3476 284 3484 339
rect 3537 318 3545 367
rect 3617 318 3625 367
rect 3657 327 3663 397
rect 3937 476 3949 482
rect 3981 476 3993 482
rect 4037 476 4049 482
rect 4171 476 4183 482
rect 4251 476 4263 482
rect 4291 476 4303 482
rect 4337 476 4349 482
rect 4417 476 4429 482
rect 4496 476 4508 482
rect 4546 476 4558 482
rect 3713 361 3721 396
rect 3803 389 3820 396
rect 3883 389 3900 396
rect 3537 312 3561 318
rect 3617 312 3641 318
rect 3719 325 3727 347
rect 3813 341 3820 389
rect 3893 341 3900 389
rect 3720 318 3745 325
rect 3549 304 3561 312
rect 3629 304 3641 312
rect 3097 258 3109 264
rect 3230 258 3242 264
rect 3330 258 3342 264
rect 3377 258 3389 264
rect 3491 258 3503 264
rect 3677 304 3729 307
rect 3689 298 3717 304
rect 3737 304 3745 318
rect 3813 284 3820 327
rect 3893 284 3900 327
rect 3958 322 3966 436
rect 4191 402 4203 404
rect 4163 396 4203 402
rect 4235 434 4243 436
rect 4271 434 4282 436
rect 4235 428 4282 434
rect 4001 361 4009 396
rect 4060 389 4077 396
rect 4007 347 4009 361
rect 3937 314 3975 322
rect 3937 304 3949 314
rect 4001 304 4009 347
rect 4060 341 4067 389
rect 4134 361 4142 396
rect 4235 373 4242 428
rect 4317 402 4329 404
rect 4317 396 4357 402
rect 4378 361 4386 396
rect 3519 258 3531 264
rect 3599 258 3611 264
rect 3697 258 3709 264
rect 3791 258 3803 264
rect 3831 258 3843 264
rect 3999 294 4009 304
rect 4060 284 4067 327
rect 4134 304 4142 347
rect 4236 331 4244 359
rect 4236 322 4266 331
rect 4436 353 4444 436
rect 4577 476 4589 482
rect 4637 476 4649 482
rect 4697 476 4709 482
rect 4519 361 4527 396
rect 4236 320 4254 322
rect 4134 293 4160 304
rect 3871 258 3883 264
rect 3911 258 3923 264
rect 3967 258 3979 264
rect 4037 258 4049 264
rect 4077 258 4089 264
rect 4378 304 4386 347
rect 4138 258 4150 264
rect 4188 258 4200 264
rect 4290 258 4302 264
rect 4360 293 4386 304
rect 4436 284 4444 339
rect 4513 325 4521 347
rect 4596 353 4604 436
rect 4656 353 4664 436
rect 4716 353 4724 436
rect 4495 318 4520 325
rect 4495 304 4503 318
rect 4320 258 4332 264
rect 4370 258 4382 264
rect 4511 304 4563 307
rect 4523 298 4551 304
rect 4596 284 4604 339
rect 4656 284 4664 339
rect 4716 284 4724 339
rect 4417 258 4429 264
rect 4531 258 4543 264
rect 4577 258 4589 264
rect 4637 258 4649 264
rect 4697 258 4709 264
rect 4782 258 4842 722
rect 4 256 4842 258
rect 4776 244 4842 256
rect 4 242 4842 244
rect 41 236 53 242
rect 103 236 115 242
rect 151 236 163 242
rect 209 236 221 242
rect 260 236 272 242
rect 316 236 328 242
rect 60 216 73 222
rect 60 210 67 216
rect 125 204 132 216
rect 21 112 27 196
rect 111 197 132 204
rect 182 210 189 216
rect 182 202 193 210
rect 79 186 86 192
rect 377 236 389 242
rect 417 236 429 242
rect 458 236 470 242
rect 591 236 603 242
rect 635 236 643 242
rect 147 186 153 188
rect 79 180 153 186
rect 235 181 243 196
rect 79 172 86 180
rect 40 164 74 172
rect 40 159 46 164
rect 66 146 93 153
rect 21 104 83 112
rect 95 108 139 114
rect 77 90 115 98
rect 133 94 139 108
rect 147 108 153 180
rect 227 167 243 181
rect 213 153 227 167
rect 147 102 187 108
rect 207 108 221 116
rect 235 104 243 167
rect 293 153 300 196
rect 400 173 407 216
rect 678 236 690 242
rect 728 236 740 242
rect 779 236 791 242
rect 837 236 849 242
rect 885 236 897 242
rect 947 236 959 242
rect 1051 236 1063 242
rect 1131 236 1143 242
rect 506 178 524 180
rect 494 169 524 178
rect 301 116 307 139
rect 301 110 328 116
rect 316 104 328 110
rect 400 111 407 159
rect 516 141 524 169
rect 573 161 580 196
rect 611 188 617 216
rect 607 182 617 188
rect 674 196 700 207
rect 927 216 940 222
rect 811 210 818 216
rect 807 202 818 210
rect 868 204 875 216
rect 933 210 940 216
rect 400 104 417 111
rect 77 84 85 90
rect 133 88 163 94
rect 181 84 187 102
rect 67 70 85 84
rect 113 70 135 82
rect 77 64 85 70
rect 127 64 139 70
rect 181 44 193 78
rect 269 96 297 102
rect 309 24 337 30
rect 518 72 525 127
rect 577 103 586 147
rect 596 121 602 176
rect 674 153 682 196
rect 757 181 765 196
rect 868 197 889 204
rect 847 186 853 188
rect 914 186 921 192
rect 757 167 773 181
rect 847 180 921 186
rect 607 112 643 120
rect 635 104 643 112
rect 674 104 682 139
rect 757 104 765 167
rect 773 153 787 167
rect 779 108 793 116
rect 577 94 581 103
rect 478 66 525 72
rect 478 64 489 66
rect 517 64 525 66
rect 703 98 743 104
rect 731 96 743 98
rect 847 108 853 180
rect 914 172 921 180
rect 926 164 960 172
rect 954 159 960 164
rect 907 146 934 153
rect 813 102 853 108
rect 861 108 905 114
rect 813 84 819 102
rect 861 94 867 108
rect 973 112 979 196
rect 1015 182 1023 196
rect 1043 196 1071 202
rect 1171 236 1183 242
rect 1211 236 1223 242
rect 1271 236 1283 242
rect 1351 236 1363 242
rect 1431 236 1443 242
rect 1491 236 1503 242
rect 1031 193 1083 196
rect 1015 175 1040 182
rect 1033 153 1041 175
rect 1116 161 1124 216
rect 1193 173 1200 216
rect 1256 161 1264 216
rect 1315 182 1323 196
rect 1343 196 1371 202
rect 1517 236 1529 242
rect 1557 236 1569 242
rect 1618 236 1630 242
rect 1668 236 1680 242
rect 1721 236 1733 242
rect 1783 236 1795 242
rect 1831 236 1843 242
rect 1889 236 1901 242
rect 1991 236 2003 242
rect 2037 236 2049 242
rect 2097 236 2109 242
rect 2137 236 2149 242
rect 1331 193 1383 196
rect 1315 175 1340 182
rect 917 104 979 112
rect 1039 104 1047 139
rect 837 88 867 94
rect 885 90 923 98
rect 915 84 923 90
rect 807 44 819 78
rect 865 70 887 82
rect 915 70 933 84
rect 861 64 873 70
rect 915 64 923 70
rect 1116 64 1124 147
rect 1193 111 1200 159
rect 1333 153 1341 175
rect 1416 161 1424 216
rect 1183 104 1200 111
rect 1256 64 1264 147
rect 1476 161 1484 216
rect 1540 173 1547 216
rect 1339 104 1347 139
rect 41 18 53 24
rect 107 18 119 24
rect 153 18 165 24
rect 211 18 223 24
rect 277 18 289 24
rect 377 18 389 24
rect 457 18 469 24
rect 497 18 509 24
rect 601 18 613 24
rect 711 18 723 24
rect 777 18 789 24
rect 835 18 847 24
rect 881 18 893 24
rect 947 18 959 24
rect 1016 18 1028 24
rect 1066 18 1078 24
rect 1131 18 1143 24
rect 1211 18 1223 24
rect 1271 18 1283 24
rect 1416 64 1424 147
rect 1476 64 1484 147
rect 1540 111 1547 159
rect 1614 196 1640 207
rect 1740 216 1753 222
rect 1740 210 1747 216
rect 1805 204 1812 216
rect 1614 153 1622 196
rect 1540 104 1557 111
rect 1614 104 1622 139
rect 1701 112 1707 196
rect 1791 197 1812 204
rect 1862 210 1869 216
rect 1862 202 1873 210
rect 1759 186 1766 192
rect 1827 186 1833 188
rect 1759 180 1833 186
rect 1915 181 1923 196
rect 1759 172 1766 180
rect 1720 164 1754 172
rect 1720 159 1726 164
rect 1746 146 1773 153
rect 1701 104 1763 112
rect 1775 108 1819 114
rect 1316 18 1328 24
rect 1366 18 1378 24
rect 1431 18 1443 24
rect 1491 18 1503 24
rect 1643 98 1683 104
rect 1671 96 1683 98
rect 1757 90 1795 98
rect 1813 94 1819 108
rect 1827 108 1833 180
rect 1907 167 1923 181
rect 1955 182 1963 196
rect 1983 196 2011 202
rect 2177 236 2189 242
rect 2217 236 2229 242
rect 2271 236 2283 242
rect 2311 236 2323 242
rect 2337 236 2349 242
rect 2377 236 2389 242
rect 2451 236 2463 242
rect 2499 236 2511 242
rect 2557 236 2569 242
rect 2605 236 2617 242
rect 2667 236 2679 242
rect 2739 236 2751 242
rect 2797 236 2809 242
rect 2845 236 2857 242
rect 2907 236 2919 242
rect 2977 236 2989 242
rect 3111 236 3123 242
rect 3155 236 3163 242
rect 3197 236 3209 242
rect 3311 236 3323 242
rect 1971 193 2023 196
rect 1955 175 1980 182
rect 1893 153 1907 167
rect 1827 102 1867 108
rect 1887 108 1901 116
rect 1915 104 1923 167
rect 1973 153 1981 175
rect 2056 161 2064 216
rect 2120 173 2127 216
rect 2200 173 2207 216
rect 1979 104 1987 139
rect 1757 84 1765 90
rect 1813 88 1843 94
rect 1861 84 1867 102
rect 1747 70 1765 84
rect 1793 70 1815 82
rect 1757 64 1765 70
rect 1807 64 1819 70
rect 1861 44 1873 78
rect 2056 64 2064 147
rect 2120 111 2127 159
rect 2200 111 2207 159
rect 2293 173 2300 216
rect 2360 173 2367 216
rect 2436 161 2444 216
rect 2647 216 2660 222
rect 2531 210 2538 216
rect 2527 202 2538 210
rect 2588 204 2595 216
rect 2653 210 2660 216
rect 2477 181 2485 196
rect 2588 197 2609 204
rect 2567 186 2573 188
rect 2634 186 2641 192
rect 2293 111 2300 159
rect 2120 104 2137 111
rect 2200 104 2217 111
rect 1517 18 1529 24
rect 1651 18 1663 24
rect 1721 18 1733 24
rect 1787 18 1799 24
rect 1833 18 1845 24
rect 1891 18 1903 24
rect 1956 18 1968 24
rect 2006 18 2018 24
rect 2283 104 2300 111
rect 2360 111 2367 159
rect 2477 167 2493 181
rect 2567 180 2641 186
rect 2360 104 2377 111
rect 2037 18 2049 24
rect 2097 18 2109 24
rect 2177 18 2189 24
rect 2311 18 2323 24
rect 2436 64 2444 147
rect 2477 104 2485 167
rect 2493 153 2507 167
rect 2499 108 2513 116
rect 2567 108 2573 180
rect 2634 172 2641 180
rect 2646 164 2680 172
rect 2674 159 2680 164
rect 2627 146 2654 153
rect 2533 102 2573 108
rect 2581 108 2625 114
rect 2533 84 2539 102
rect 2581 94 2587 108
rect 2693 112 2699 196
rect 2637 104 2699 112
rect 2557 88 2587 94
rect 2605 90 2643 98
rect 2635 84 2643 90
rect 2527 44 2539 78
rect 2585 70 2607 82
rect 2635 70 2653 84
rect 2581 64 2593 70
rect 2635 64 2643 70
rect 2887 216 2900 222
rect 2771 210 2778 216
rect 2767 202 2778 210
rect 2828 204 2835 216
rect 2893 210 2900 216
rect 2717 181 2725 196
rect 2828 197 2849 204
rect 2807 186 2813 188
rect 2874 186 2881 192
rect 2717 167 2733 181
rect 2807 180 2881 186
rect 2717 104 2725 167
rect 2733 153 2747 167
rect 2739 108 2753 116
rect 2807 108 2813 180
rect 2874 172 2881 180
rect 2886 164 2920 172
rect 2914 159 2920 164
rect 2867 146 2894 153
rect 2773 102 2813 108
rect 2821 108 2865 114
rect 2773 84 2779 102
rect 2821 94 2827 108
rect 2933 112 2939 196
rect 2969 196 2997 200
rect 3009 230 3037 236
rect 2957 194 3009 196
rect 3019 186 3025 196
rect 2996 179 3025 186
rect 2996 153 3004 179
rect 3093 161 3100 196
rect 3131 188 3137 216
rect 3189 196 3217 202
rect 3177 193 3229 196
rect 3339 236 3351 242
rect 3490 236 3502 242
rect 3551 236 3563 242
rect 3127 182 3137 188
rect 3237 182 3245 196
rect 2877 104 2939 112
rect 2997 104 3005 139
rect 2797 88 2827 94
rect 2845 90 2883 98
rect 2875 84 2883 90
rect 2767 44 2779 78
rect 2825 70 2847 82
rect 2875 70 2893 84
rect 2821 64 2833 70
rect 2875 64 2883 70
rect 3097 103 3106 147
rect 3116 121 3122 176
rect 3220 175 3245 182
rect 3219 153 3227 175
rect 3296 161 3304 216
rect 3369 188 3381 196
rect 3357 182 3381 188
rect 3127 112 3163 120
rect 3155 104 3163 112
rect 3213 104 3221 139
rect 3097 94 3101 103
rect 3296 64 3304 147
rect 3357 133 3365 182
rect 3436 178 3454 180
rect 3436 169 3466 178
rect 3598 236 3610 242
rect 3648 236 3660 242
rect 3436 141 3444 169
rect 3536 161 3544 216
rect 3594 196 3620 207
rect 3691 236 3703 242
rect 3731 236 3743 242
rect 3757 236 3769 242
rect 3837 236 3849 242
rect 3917 236 3929 242
rect 3957 236 3969 242
rect 4070 236 4082 242
rect 3594 153 3602 196
rect 3713 173 3720 216
rect 3357 64 3365 119
rect 3435 72 3442 127
rect 3435 66 3482 72
rect 3435 64 3443 66
rect 2337 18 2349 24
rect 2451 18 2463 24
rect 2497 18 2509 24
rect 2555 18 2567 24
rect 2601 18 2613 24
rect 2667 18 2679 24
rect 2737 18 2749 24
rect 2795 18 2807 24
rect 2841 18 2853 24
rect 2907 18 2919 24
rect 2957 18 2969 24
rect 3027 18 3039 24
rect 3121 18 3133 24
rect 3182 18 3194 24
rect 3232 18 3244 24
rect 3311 18 3323 24
rect 3471 64 3482 66
rect 3536 64 3544 147
rect 3776 161 3784 216
rect 3829 196 3857 202
rect 3817 193 3869 196
rect 3877 182 3885 196
rect 3860 175 3885 182
rect 3594 104 3602 139
rect 3713 111 3720 159
rect 3703 104 3720 111
rect 3623 98 3663 104
rect 3651 96 3663 98
rect 3776 64 3784 147
rect 3859 153 3867 175
rect 3940 173 3947 216
rect 3853 104 3861 139
rect 3940 111 3947 159
rect 4016 178 4034 180
rect 4016 169 4046 178
rect 4099 236 4111 242
rect 4250 236 4262 242
rect 4329 236 4341 242
rect 4430 236 4442 242
rect 4129 188 4141 196
rect 4117 182 4141 188
rect 4016 141 4024 169
rect 3940 104 3957 111
rect 3337 18 3349 24
rect 3377 18 3389 24
rect 3451 18 3463 24
rect 3491 18 3503 24
rect 3551 18 3563 24
rect 3631 18 3643 24
rect 3731 18 3743 24
rect 3757 18 3769 24
rect 3822 18 3834 24
rect 3872 18 3884 24
rect 4015 72 4022 127
rect 4117 133 4125 182
rect 4196 178 4214 180
rect 4196 169 4226 178
rect 4299 188 4311 196
rect 4299 182 4323 188
rect 4196 141 4204 169
rect 4015 66 4062 72
rect 4015 64 4023 66
rect 4051 64 4062 66
rect 4117 64 4125 119
rect 4195 72 4202 127
rect 4315 133 4323 182
rect 4376 178 4394 180
rect 4376 169 4406 178
rect 4459 236 4471 242
rect 4538 236 4550 242
rect 4658 236 4670 242
rect 4708 236 4720 242
rect 4489 188 4501 196
rect 4477 182 4501 188
rect 4376 141 4384 169
rect 4195 66 4242 72
rect 4195 64 4203 66
rect 3917 18 3929 24
rect 4031 18 4043 24
rect 4071 18 4083 24
rect 4231 64 4242 66
rect 4315 64 4323 119
rect 4375 72 4382 127
rect 4477 133 4485 182
rect 4654 196 4680 207
rect 4586 178 4604 180
rect 4574 169 4604 178
rect 4596 141 4604 169
rect 4654 153 4662 196
rect 4375 66 4422 72
rect 4375 64 4383 66
rect 4097 18 4109 24
rect 4137 18 4149 24
rect 4211 18 4223 24
rect 4251 18 4263 24
rect 4411 64 4422 66
rect 4477 64 4485 119
rect 4598 72 4605 127
rect 4654 104 4662 139
rect 4558 66 4605 72
rect 4558 64 4569 66
rect 4291 18 4303 24
rect 4331 18 4343 24
rect 4391 18 4403 24
rect 4431 18 4443 24
rect 4457 18 4469 24
rect 4497 18 4509 24
rect 4597 64 4605 66
rect 4683 98 4723 104
rect 4711 96 4723 98
rect 4537 18 4549 24
rect 4577 18 4589 24
rect 4691 18 4703 24
rect -62 16 4776 18
rect -62 4 4 16
rect -62 2 4776 4
rect 4782 2 4842 242
<< m2contact >>
rect 33 4459 47 4473
rect 73 4459 87 4473
rect 113 4447 127 4461
rect 133 4439 147 4453
rect 153 4447 167 4461
rect 213 4459 227 4473
rect 233 4467 247 4481
rect 253 4459 267 4473
rect 273 4459 287 4473
rect 193 4439 207 4453
rect 393 4479 407 4493
rect 473 4479 487 4493
rect 313 4459 327 4473
rect 373 4459 387 4473
rect 413 4459 427 4473
rect 453 4459 467 4473
rect 493 4459 507 4473
rect 513 4459 527 4473
rect 553 4459 567 4473
rect 613 4467 627 4481
rect 633 4479 647 4493
rect 673 4479 687 4493
rect 733 4479 747 4493
rect 833 4516 847 4530
rect 973 4516 987 4530
rect 813 4487 827 4501
rect 653 4459 667 4473
rect 693 4459 707 4473
rect 753 4467 767 4481
rect 833 4422 847 4436
rect 893 4459 907 4473
rect 933 4459 947 4473
rect 1173 4516 1187 4530
rect 1313 4516 1327 4530
rect 1033 4459 1047 4473
rect 1053 4467 1067 4481
rect 1073 4459 1087 4473
rect 1153 4487 1167 4501
rect 1093 4439 1107 4453
rect 833 4384 847 4398
rect 973 4390 987 4404
rect 1173 4422 1187 4436
rect 1233 4459 1247 4473
rect 1273 4459 1287 4473
rect 1513 4516 1527 4530
rect 1373 4459 1387 4473
rect 1393 4467 1407 4481
rect 1413 4459 1427 4473
rect 1433 4439 1447 4453
rect 1653 4516 1667 4530
rect 1553 4459 1567 4473
rect 1593 4459 1607 4473
rect 1173 4384 1187 4398
rect 1313 4390 1327 4404
rect 1673 4487 1687 4501
rect 1653 4422 1667 4436
rect 1833 4516 1847 4530
rect 1713 4447 1727 4461
rect 1973 4516 1987 4530
rect 1813 4487 1827 4501
rect 1733 4439 1747 4453
rect 1753 4447 1767 4461
rect 1513 4390 1527 4404
rect 1653 4384 1667 4398
rect 1833 4422 1847 4436
rect 1893 4459 1907 4473
rect 1933 4459 1947 4473
rect 2033 4459 2047 4473
rect 2053 4467 2067 4481
rect 2073 4459 2087 4473
rect 2093 4467 2107 4481
rect 2113 4459 2127 4473
rect 2173 4447 2187 4461
rect 2293 4459 2307 4473
rect 2313 4467 2327 4481
rect 2333 4459 2347 4473
rect 2373 4467 2387 4481
rect 2393 4479 2407 4493
rect 2433 4479 2447 4493
rect 1833 4384 1847 4398
rect 1973 4390 1987 4404
rect 2193 4439 2207 4453
rect 2233 4439 2247 4453
rect 2273 4439 2287 4453
rect 2213 4419 2227 4433
rect 2413 4459 2427 4473
rect 2453 4459 2467 4473
rect 2513 4467 2527 4481
rect 2533 4479 2547 4493
rect 2553 4459 2567 4473
rect 2573 4467 2587 4481
rect 2593 4459 2607 4473
rect 2653 4459 2667 4473
rect 2613 4439 2627 4453
rect 2693 4459 2707 4473
rect 2733 4459 2747 4473
rect 2773 4459 2787 4473
rect 2833 4459 2847 4473
rect 2873 4459 2887 4473
rect 2913 4447 2927 4461
rect 3013 4459 3027 4473
rect 2933 4439 2947 4453
rect 2973 4439 2987 4453
rect 2953 4419 2967 4433
rect 3033 4447 3047 4461
rect 3073 4459 3087 4473
rect 3113 4459 3127 4473
rect 3153 4459 3167 4473
rect 3193 4447 3207 4461
rect 3213 4439 3227 4453
rect 3253 4439 3267 4453
rect 3273 4447 3287 4461
rect 3353 4467 3367 4481
rect 3373 4479 3387 4493
rect 3393 4467 3407 4481
rect 3293 4439 3307 4453
rect 3313 4447 3327 4461
rect 3413 4459 3427 4473
rect 3233 4419 3247 4433
rect 3453 4513 3467 4527
rect 3453 4479 3467 4493
rect 3473 4467 3487 4481
rect 3453 4433 3467 4447
rect 3513 4447 3527 4461
rect 3693 4467 3707 4481
rect 3713 4479 3727 4493
rect 3733 4467 3747 4481
rect 3533 4439 3547 4453
rect 3553 4447 3567 4461
rect 3593 4439 3607 4453
rect 3633 4439 3647 4453
rect 3653 4447 3667 4461
rect 3753 4459 3767 4473
rect 3793 4459 3807 4473
rect 3813 4467 3827 4481
rect 3833 4459 3847 4473
rect 3933 4459 3947 4473
rect 3953 4467 3967 4481
rect 3973 4459 3987 4473
rect 4193 4467 4207 4481
rect 4213 4479 4227 4493
rect 4233 4467 4247 4481
rect 3613 4419 3627 4433
rect 3853 4439 3867 4453
rect 3913 4439 3927 4453
rect 4013 4447 4027 4461
rect 4033 4439 4047 4453
rect 4073 4439 4087 4453
rect 4113 4447 4127 4461
rect 4253 4459 4267 4473
rect 4053 4419 4067 4433
rect 4133 4439 4147 4453
rect 4173 4439 4187 4453
rect 4153 4419 4167 4433
rect 4293 4447 4307 4461
rect 4313 4439 4327 4453
rect 4333 4447 4347 4461
rect 4393 4459 4407 4473
rect 4413 4467 4427 4481
rect 4433 4479 4447 4493
rect 4453 4467 4467 4481
rect 4493 4467 4507 4481
rect 4513 4479 4527 4493
rect 4533 4439 4547 4453
rect 4573 4439 4587 4453
rect 4593 4447 4607 4461
rect 4553 4419 4567 4433
rect 4633 4439 4647 4453
rect 4673 4439 4687 4453
rect 4693 4447 4707 4461
rect 4653 4419 4667 4433
rect 33 4207 47 4221
rect 53 4187 67 4201
rect 73 4179 87 4193
rect 93 4187 107 4201
rect 133 4187 147 4201
rect 153 4199 167 4213
rect 193 4187 207 4201
rect 213 4187 227 4201
rect 253 4187 267 4201
rect 313 4187 327 4201
rect 233 4167 247 4181
rect 333 4179 347 4193
rect 353 4167 367 4181
rect 373 4179 387 4193
rect 393 4187 407 4201
rect 433 4199 447 4213
rect 613 4227 627 4241
rect 593 4207 607 4221
rect 633 4207 647 4221
rect 453 4187 467 4201
rect 513 4187 527 4201
rect 653 4199 667 4213
rect 533 4179 547 4193
rect 553 4167 567 4181
rect 573 4179 587 4193
rect 693 4179 707 4193
rect 713 4167 727 4181
rect 733 4179 747 4193
rect 753 4187 767 4201
rect 793 4187 807 4201
rect 833 4199 847 4213
rect 913 4207 927 4221
rect 853 4187 867 4201
rect 933 4187 947 4201
rect 953 4179 967 4193
rect 973 4187 987 4201
rect 1193 4233 1207 4247
rect 1013 4179 1027 4193
rect 1053 4187 1067 4201
rect 1093 4187 1107 4201
rect 1133 4187 1147 4201
rect 1173 4187 1187 4201
rect 1033 4167 1047 4181
rect 1073 4167 1087 4181
rect 1153 4167 1167 4181
rect 1173 4153 1187 4167
rect 1213 4187 1227 4201
rect 1253 4187 1267 4201
rect 1393 4262 1407 4276
rect 1533 4256 1547 4270
rect 1233 4167 1247 4181
rect 1293 4167 1307 4181
rect 1313 4179 1327 4193
rect 1393 4224 1407 4238
rect 1373 4159 1387 4173
rect 1453 4187 1467 4201
rect 1493 4187 1507 4201
rect 1393 4130 1407 4144
rect 1653 4207 1667 4221
rect 1593 4187 1607 4201
rect 1613 4179 1627 4193
rect 1633 4187 1647 4201
rect 1693 4187 1707 4201
rect 1733 4187 1747 4201
rect 1873 4262 1887 4276
rect 2013 4256 2027 4270
rect 1713 4167 1727 4181
rect 1793 4179 1807 4193
rect 1533 4130 1547 4144
rect 1813 4167 1827 4181
rect 1873 4224 1887 4238
rect 1853 4159 1867 4173
rect 1933 4187 1947 4201
rect 1973 4187 1987 4201
rect 1873 4130 1887 4144
rect 2093 4199 2107 4213
rect 2113 4207 2127 4221
rect 2133 4199 2147 4213
rect 2173 4187 2187 4201
rect 2153 4167 2167 4181
rect 2213 4179 2227 4193
rect 2273 4187 2287 4201
rect 2293 4179 2307 4193
rect 2313 4187 2327 4201
rect 2013 4130 2027 4144
rect 2333 4179 2347 4193
rect 2353 4187 2367 4201
rect 2373 4199 2387 4213
rect 2393 4207 2407 4221
rect 2413 4199 2427 4213
rect 2473 4207 2487 4221
rect 2493 4187 2507 4201
rect 2513 4179 2527 4193
rect 2533 4187 2547 4201
rect 2573 4187 2587 4201
rect 2613 4187 2627 4201
rect 2593 4167 2607 4181
rect 2633 4179 2647 4193
rect 2653 4167 2667 4181
rect 2673 4179 2687 4193
rect 2693 4187 2707 4201
rect 2753 4187 2767 4201
rect 2773 4179 2787 4193
rect 2793 4167 2807 4181
rect 2813 4179 2827 4193
rect 2833 4187 2847 4201
rect 2993 4253 3007 4267
rect 2973 4227 2987 4241
rect 2873 4187 2887 4201
rect 2933 4199 2947 4213
rect 2953 4207 2967 4221
rect 2993 4207 3007 4221
rect 2993 4173 3007 4187
rect 3073 4227 3087 4241
rect 3033 4199 3047 4213
rect 3053 4207 3067 4221
rect 3093 4207 3107 4221
rect 3113 4199 3127 4213
rect 3133 4207 3147 4221
rect 3153 4199 3167 4213
rect 3313 4227 3327 4241
rect 3353 4233 3367 4247
rect 3273 4199 3287 4213
rect 3293 4207 3307 4221
rect 3333 4207 3347 4221
rect 3213 4179 3227 4193
rect 3233 4167 3247 4181
rect 3313 4173 3327 4187
rect 3413 4227 3427 4241
rect 3373 4199 3387 4213
rect 3393 4207 3407 4221
rect 3433 4207 3447 4221
rect 3513 4227 3527 4241
rect 3473 4199 3487 4213
rect 3493 4207 3507 4221
rect 3533 4207 3547 4221
rect 3613 4227 3627 4241
rect 3673 4227 3687 4241
rect 3573 4199 3587 4213
rect 3593 4207 3607 4221
rect 3633 4207 3647 4221
rect 3653 4207 3667 4221
rect 3693 4207 3707 4221
rect 3713 4199 3727 4213
rect 3913 4207 3927 4221
rect 3753 4179 3767 4193
rect 3773 4167 3787 4181
rect 3793 4179 3807 4193
rect 3813 4187 3827 4201
rect 3853 4187 3867 4201
rect 3873 4179 3887 4193
rect 3893 4187 3907 4201
rect 4173 4227 4187 4241
rect 4233 4227 4247 4241
rect 3953 4167 3967 4181
rect 3973 4179 3987 4193
rect 4013 4179 4027 4193
rect 4033 4167 4047 4181
rect 4053 4179 4067 4193
rect 4073 4187 4087 4201
rect 4133 4199 4147 4213
rect 4153 4207 4167 4221
rect 4193 4207 4207 4221
rect 4213 4207 4227 4221
rect 4253 4207 4267 4221
rect 4273 4199 4287 4213
rect 4473 4207 4487 4221
rect 4313 4179 4327 4193
rect 4333 4167 4347 4181
rect 4353 4179 4367 4193
rect 4373 4187 4387 4201
rect 4413 4187 4427 4201
rect 4433 4179 4447 4193
rect 4453 4187 4467 4201
rect 4513 4187 4527 4201
rect 4533 4179 4547 4193
rect 4553 4187 4567 4201
rect 4573 4179 4587 4193
rect 4593 4187 4607 4201
rect 4653 4187 4667 4201
rect 4693 4187 4707 4201
rect 4673 4167 4687 4181
rect 33 3967 47 3981
rect 53 3959 67 3973
rect 73 3967 87 3981
rect 113 3967 127 3981
rect 213 3999 227 4013
rect 133 3959 147 3973
rect 153 3967 167 3981
rect 193 3979 207 3993
rect 233 3979 247 3993
rect 253 3979 267 3993
rect 273 3987 287 4001
rect 293 3979 307 3993
rect 373 3987 387 4001
rect 393 3999 407 4013
rect 433 3987 447 4001
rect 453 3999 467 4013
rect 513 3999 527 4013
rect 313 3959 327 3973
rect 493 3979 507 3993
rect 533 3979 547 3993
rect 553 3979 567 3993
rect 593 3967 607 3981
rect 613 3979 627 3993
rect 653 3979 667 3993
rect 673 3987 687 4001
rect 753 3999 767 4013
rect 693 3979 707 3993
rect 773 3987 787 4001
rect 713 3959 727 3973
rect 813 3979 827 3993
rect 833 3987 847 4001
rect 873 3993 887 4007
rect 853 3979 867 3993
rect 873 3959 887 3973
rect 913 3967 927 3981
rect 1013 3987 1027 4001
rect 1033 3999 1047 4013
rect 1093 3999 1107 4013
rect 1133 3999 1147 4013
rect 933 3959 947 3973
rect 953 3967 967 3981
rect 893 3933 907 3947
rect 1073 3979 1087 3993
rect 1113 3979 1127 3993
rect 1153 3987 1167 4001
rect 1213 3999 1227 4013
rect 1273 3999 1287 4013
rect 1193 3979 1207 3993
rect 1233 3979 1247 3993
rect 1293 3987 1307 4001
rect 1373 3999 1387 4013
rect 1353 3979 1367 3993
rect 1393 3979 1407 3993
rect 1433 3987 1447 4001
rect 1453 3999 1467 4013
rect 1473 3979 1487 3993
rect 1493 3987 1507 4001
rect 1513 3979 1527 3993
rect 1573 3979 1587 3993
rect 1593 3987 1607 4001
rect 1613 3979 1627 3993
rect 1633 3987 1647 4001
rect 1653 3979 1667 3993
rect 1533 3959 1547 3973
rect 1693 3967 1707 3981
rect 1713 3959 1727 3973
rect 1733 3967 1747 3981
rect 1793 3979 1807 3993
rect 1813 3987 1827 4001
rect 1833 3999 1847 4013
rect 1853 3987 1867 4001
rect 1873 3959 1887 3973
rect 1913 3959 1927 3973
rect 1933 3967 1947 3981
rect 2013 3979 2027 3993
rect 2033 3987 2047 4001
rect 2053 3979 2067 3993
rect 2093 3987 2107 4001
rect 2113 3999 2127 4013
rect 1893 3939 1907 3953
rect 1993 3959 2007 3973
rect 2153 3967 2167 3981
rect 2173 3959 2187 3973
rect 2213 3959 2227 3973
rect 2253 3967 2267 3981
rect 2353 3979 2367 3993
rect 2373 3987 2387 4001
rect 2393 3999 2407 4013
rect 2413 3987 2427 4001
rect 2453 3987 2467 4001
rect 2473 3999 2487 4013
rect 2573 4013 2587 4027
rect 2193 3939 2207 3953
rect 2273 3959 2287 3973
rect 2313 3959 2327 3973
rect 2293 3939 2307 3953
rect 2533 3979 2547 3993
rect 2553 3987 2567 4001
rect 2573 3979 2587 3993
rect 2513 3959 2527 3973
rect 2693 4033 2707 4047
rect 2613 3967 2627 3981
rect 2593 3933 2607 3947
rect 2633 3959 2647 3973
rect 2673 3959 2687 3973
rect 2713 3979 2727 3993
rect 2733 3987 2747 4001
rect 2753 3999 2767 4013
rect 2773 3987 2787 4001
rect 2833 3979 2847 3993
rect 2853 3987 2867 4001
rect 2873 3979 2887 3993
rect 2893 3979 2907 3993
rect 2913 3987 2927 4001
rect 2933 3979 2947 3993
rect 3073 3993 3087 4007
rect 2653 3939 2667 3953
rect 2693 3953 2707 3967
rect 2813 3959 2827 3973
rect 2953 3959 2967 3973
rect 3013 3967 3027 3981
rect 3033 3959 3047 3973
rect 3073 3959 3087 3973
rect 3053 3939 3067 3953
rect 3073 3913 3087 3927
rect 3113 3987 3127 4001
rect 3133 3999 3147 4013
rect 3153 3979 3167 3993
rect 3173 3987 3187 4001
rect 3213 3993 3227 4007
rect 3193 3979 3207 3993
rect 3213 3959 3227 3973
rect 3253 3987 3267 4001
rect 3273 3999 3287 4013
rect 3293 3987 3307 4001
rect 3313 3979 3327 3993
rect 3353 3979 3367 3993
rect 3373 3987 3387 4001
rect 3393 3979 3407 3993
rect 3493 3979 3507 3993
rect 3513 3987 3527 4001
rect 3533 3979 3547 3993
rect 3593 3979 3607 3993
rect 3613 3987 3627 4001
rect 3633 3979 3647 3993
rect 3673 3979 3687 3993
rect 3693 3987 3707 4001
rect 3713 3999 3727 4013
rect 3733 3987 3747 4001
rect 3273 3953 3287 3967
rect 3413 3959 3427 3973
rect 3473 3959 3487 3973
rect 3573 3959 3587 3973
rect 3773 3967 3787 3981
rect 3793 3959 3807 3973
rect 3833 3959 3847 3973
rect 3873 3967 3887 3981
rect 3893 3959 3907 3973
rect 3913 3967 3927 3981
rect 3953 3967 3967 3981
rect 3973 3959 3987 3973
rect 3993 3967 4007 3981
rect 4013 3967 4027 3981
rect 4033 3959 4047 3973
rect 4053 3967 4067 3981
rect 4113 3967 4127 3981
rect 4233 3979 4247 3993
rect 4253 3987 4267 4001
rect 4273 3979 4287 3993
rect 4293 3979 4307 3993
rect 4313 3987 4327 4001
rect 4333 3979 4347 3993
rect 4413 3987 4427 4001
rect 4433 3999 4447 4013
rect 3813 3939 3827 3953
rect 4133 3959 4147 3973
rect 4173 3959 4187 3973
rect 4213 3959 4227 3973
rect 4153 3939 4167 3953
rect 4353 3959 4367 3973
rect 4653 3987 4667 4001
rect 4673 3999 4687 4013
rect 4693 3987 4707 4001
rect 4473 3967 4487 3981
rect 4493 3959 4507 3973
rect 4533 3959 4547 3973
rect 4573 3967 4587 3981
rect 4713 3979 4727 3993
rect 4513 3939 4527 3953
rect 4593 3959 4607 3973
rect 4633 3959 4647 3973
rect 4613 3939 4627 3953
rect 33 3727 47 3741
rect 53 3707 67 3721
rect 73 3699 87 3713
rect 93 3707 107 3721
rect 213 3782 227 3796
rect 353 3776 367 3790
rect 133 3699 147 3713
rect 153 3687 167 3701
rect 213 3744 227 3758
rect 193 3679 207 3693
rect 273 3707 287 3721
rect 313 3707 327 3721
rect 213 3650 227 3664
rect 433 3727 447 3741
rect 453 3707 467 3721
rect 473 3699 487 3713
rect 493 3707 507 3721
rect 513 3707 527 3721
rect 553 3719 567 3733
rect 573 3707 587 3721
rect 833 3776 847 3790
rect 973 3782 987 3796
rect 353 3650 367 3664
rect 633 3699 647 3713
rect 673 3707 687 3721
rect 733 3719 747 3733
rect 753 3727 767 3741
rect 693 3687 707 3701
rect 773 3719 787 3733
rect 873 3707 887 3721
rect 913 3707 927 3721
rect 973 3744 987 3758
rect 993 3679 1007 3693
rect 833 3650 847 3664
rect 1153 3782 1167 3796
rect 1293 3776 1307 3790
rect 1053 3707 1067 3721
rect 1093 3707 1107 3721
rect 1153 3744 1167 3758
rect 1133 3679 1147 3693
rect 1213 3707 1227 3721
rect 1253 3707 1267 3721
rect 973 3650 987 3664
rect 1153 3650 1167 3664
rect 1733 3782 1747 3796
rect 1873 3776 1887 3790
rect 1413 3727 1427 3741
rect 1353 3707 1367 3721
rect 1373 3699 1387 3713
rect 1393 3707 1407 3721
rect 1453 3719 1467 3733
rect 1473 3727 1487 3741
rect 1293 3650 1307 3664
rect 1493 3719 1507 3733
rect 1533 3719 1547 3733
rect 1553 3727 1567 3741
rect 1573 3719 1587 3733
rect 1613 3707 1627 3721
rect 1653 3707 1667 3721
rect 1733 3744 1747 3758
rect 1713 3679 1727 3693
rect 1793 3707 1807 3721
rect 1833 3707 1847 3721
rect 1733 3650 1747 3664
rect 1953 3699 1967 3713
rect 2013 3707 2027 3721
rect 2173 3747 2187 3761
rect 2153 3727 2167 3741
rect 2193 3727 2207 3741
rect 2213 3719 2227 3733
rect 2273 3727 2287 3741
rect 2413 3747 2427 3761
rect 1873 3650 1887 3664
rect 1973 3687 1987 3701
rect 2033 3699 2047 3713
rect 2053 3687 2067 3701
rect 2073 3699 2087 3713
rect 2113 3699 2127 3713
rect 2133 3687 2147 3701
rect 2293 3707 2307 3721
rect 2313 3699 2327 3713
rect 2333 3707 2347 3721
rect 2373 3719 2387 3733
rect 2393 3727 2407 3741
rect 2433 3727 2447 3741
rect 2553 3733 2567 3747
rect 2613 3747 2627 3761
rect 2473 3707 2487 3721
rect 2493 3699 2507 3713
rect 2513 3687 2527 3701
rect 2533 3699 2547 3713
rect 2573 3719 2587 3733
rect 2593 3727 2607 3741
rect 2633 3727 2647 3741
rect 2853 3733 2867 3747
rect 2653 3699 2667 3713
rect 2553 3673 2567 3687
rect 2673 3687 2687 3701
rect 2693 3699 2707 3713
rect 2713 3707 2727 3721
rect 2773 3707 2787 3721
rect 2793 3699 2807 3713
rect 2813 3687 2827 3701
rect 2833 3699 2847 3713
rect 3033 3747 3047 3761
rect 2993 3719 3007 3733
rect 3013 3727 3027 3741
rect 3053 3727 3067 3741
rect 3233 3747 3247 3761
rect 2873 3699 2887 3713
rect 2853 3653 2867 3667
rect 2893 3687 2907 3701
rect 2933 3699 2947 3713
rect 2953 3687 2967 3701
rect 3093 3707 3107 3721
rect 3193 3719 3207 3733
rect 3213 3727 3227 3741
rect 3253 3727 3267 3741
rect 3113 3699 3127 3713
rect 3133 3687 3147 3701
rect 3153 3699 3167 3713
rect 3353 3727 3367 3741
rect 3293 3699 3307 3713
rect 3373 3707 3387 3721
rect 3313 3687 3327 3701
rect 3393 3699 3407 3713
rect 3413 3707 3427 3721
rect 3453 3719 3467 3733
rect 3473 3727 3487 3741
rect 3493 3719 3507 3733
rect 3513 3707 3527 3721
rect 3553 3719 3567 3733
rect 3793 3773 3807 3787
rect 3773 3747 3787 3761
rect 3573 3707 3587 3721
rect 3633 3707 3647 3721
rect 3733 3719 3747 3733
rect 3753 3727 3767 3741
rect 3793 3727 3807 3741
rect 3653 3699 3667 3713
rect 3673 3687 3687 3701
rect 3693 3699 3707 3713
rect 3993 3727 4007 3741
rect 4133 3727 4147 3741
rect 4393 3747 4407 3761
rect 4373 3727 4387 3741
rect 4413 3727 4427 3741
rect 3833 3699 3847 3713
rect 3813 3653 3827 3667
rect 3853 3687 3867 3701
rect 3873 3699 3887 3713
rect 3893 3687 3907 3701
rect 3913 3699 3927 3713
rect 3933 3707 3947 3721
rect 4013 3707 4027 3721
rect 4033 3699 4047 3713
rect 4053 3707 4067 3721
rect 4073 3707 4087 3721
rect 4093 3699 4107 3713
rect 4113 3707 4127 3721
rect 4173 3699 4187 3713
rect 4193 3687 4207 3701
rect 4213 3699 4227 3713
rect 4233 3707 4247 3721
rect 4293 3707 4307 3721
rect 4433 3719 4447 3733
rect 4313 3699 4327 3713
rect 4333 3687 4347 3701
rect 4353 3699 4367 3713
rect 4593 3747 4607 3761
rect 4653 3747 4667 3761
rect 4553 3719 4567 3733
rect 4573 3727 4587 3741
rect 4613 3727 4627 3741
rect 4633 3727 4647 3741
rect 4673 3727 4687 3741
rect 4693 3719 4707 3733
rect 4493 3699 4507 3713
rect 4513 3687 4527 3701
rect 53 3556 67 3570
rect 193 3556 207 3570
rect 93 3499 107 3513
rect 133 3499 147 3513
rect 213 3527 227 3541
rect 193 3462 207 3476
rect 273 3487 287 3501
rect 293 3479 307 3493
rect 313 3487 327 3501
rect 373 3499 387 3513
rect 393 3507 407 3521
rect 413 3499 427 3513
rect 353 3479 367 3493
rect 53 3430 67 3444
rect 193 3424 207 3438
rect 453 3487 467 3501
rect 593 3513 607 3527
rect 473 3479 487 3493
rect 493 3487 507 3501
rect 533 3487 547 3501
rect 553 3479 567 3493
rect 593 3479 607 3493
rect 573 3459 587 3473
rect 593 3433 607 3447
rect 633 3507 647 3521
rect 653 3519 667 3533
rect 713 3499 727 3513
rect 733 3507 747 3521
rect 753 3499 767 3513
rect 813 3499 827 3513
rect 833 3507 847 3521
rect 873 3519 887 3533
rect 1053 3556 1067 3570
rect 1193 3556 1207 3570
rect 853 3499 867 3513
rect 893 3507 907 3521
rect 973 3519 987 3533
rect 1033 3527 1047 3541
rect 693 3479 707 3493
rect 793 3479 807 3493
rect 953 3499 967 3513
rect 993 3499 1007 3513
rect 1053 3462 1067 3476
rect 1113 3499 1127 3513
rect 1153 3499 1167 3513
rect 1253 3519 1267 3533
rect 1273 3507 1287 3521
rect 1333 3519 1347 3533
rect 1053 3424 1067 3438
rect 1193 3430 1207 3444
rect 1313 3499 1327 3513
rect 1353 3499 1367 3513
rect 1393 3499 1407 3513
rect 1413 3507 1427 3521
rect 1433 3499 1447 3513
rect 1453 3479 1467 3493
rect 1493 3487 1507 3501
rect 1513 3479 1527 3493
rect 1533 3487 1547 3501
rect 1593 3499 1607 3513
rect 1753 3556 1767 3570
rect 1893 3556 1907 3570
rect 1633 3499 1647 3513
rect 1673 3507 1687 3521
rect 1693 3519 1707 3533
rect 1733 3527 1747 3541
rect 1753 3462 1767 3476
rect 1813 3499 1827 3513
rect 1853 3499 1867 3513
rect 1953 3499 1967 3513
rect 1973 3507 1987 3521
rect 1993 3499 2007 3513
rect 2013 3507 2027 3521
rect 2033 3499 2047 3513
rect 2073 3487 2087 3501
rect 2093 3479 2107 3493
rect 2113 3487 2127 3501
rect 2173 3499 2187 3513
rect 2193 3507 2207 3521
rect 2213 3519 2227 3533
rect 2233 3507 2247 3521
rect 2373 3507 2387 3521
rect 2393 3519 2407 3533
rect 1753 3424 1767 3438
rect 1893 3430 1907 3444
rect 2273 3487 2287 3501
rect 2293 3479 2307 3493
rect 2333 3479 2347 3493
rect 2313 3459 2327 3473
rect 2433 3487 2447 3501
rect 2453 3479 2467 3493
rect 2493 3479 2507 3493
rect 2533 3487 2547 3501
rect 2653 3499 2667 3513
rect 2673 3507 2687 3521
rect 2693 3499 2707 3513
rect 2713 3499 2727 3513
rect 2733 3507 2747 3521
rect 2753 3499 2767 3513
rect 2473 3459 2487 3473
rect 2553 3479 2567 3493
rect 2593 3479 2607 3493
rect 2633 3479 2647 3493
rect 2573 3459 2587 3473
rect 2773 3479 2787 3493
rect 2813 3487 2827 3501
rect 2833 3479 2847 3493
rect 2853 3487 2867 3501
rect 2893 3499 2907 3513
rect 2913 3507 2927 3521
rect 2933 3499 2947 3513
rect 2953 3479 2967 3493
rect 2993 3533 3007 3547
rect 3013 3519 3027 3533
rect 2993 3499 3007 3513
rect 3033 3499 3047 3513
rect 3113 3499 3127 3513
rect 3133 3507 3147 3521
rect 3153 3499 3167 3513
rect 3173 3499 3187 3513
rect 3193 3507 3207 3521
rect 3213 3499 3227 3513
rect 3233 3507 3247 3521
rect 3253 3499 3267 3513
rect 3093 3479 3107 3493
rect 2973 3453 2987 3467
rect 3293 3487 3307 3501
rect 3313 3479 3327 3493
rect 3333 3487 3347 3501
rect 3373 3487 3387 3501
rect 3393 3479 3407 3493
rect 3413 3487 3427 3501
rect 3453 3487 3467 3501
rect 3473 3479 3487 3493
rect 3493 3487 3507 3501
rect 3413 3453 3427 3467
rect 3453 3433 3467 3447
rect 3493 3453 3507 3467
rect 3533 3533 3547 3547
rect 3553 3519 3567 3533
rect 3533 3499 3547 3513
rect 3573 3499 3587 3513
rect 3613 3487 3627 3501
rect 3633 3479 3647 3493
rect 3653 3487 3667 3501
rect 3693 3487 3707 3501
rect 3713 3479 3727 3493
rect 3733 3487 3747 3501
rect 3793 3487 3807 3501
rect 3893 3519 3907 3533
rect 3813 3479 3827 3493
rect 3833 3487 3847 3501
rect 3873 3499 3887 3513
rect 3913 3499 3927 3513
rect 3933 3487 3947 3501
rect 3953 3479 3967 3493
rect 3973 3487 3987 3501
rect 4013 3487 4027 3501
rect 4033 3479 4047 3493
rect 4053 3487 4067 3501
rect 4093 3499 4107 3513
rect 4113 3507 4127 3521
rect 4133 3499 4147 3513
rect 4393 3507 4407 3521
rect 4413 3519 4427 3533
rect 4433 3507 4447 3521
rect 4153 3479 4167 3493
rect 4213 3487 4227 3501
rect 4233 3479 4247 3493
rect 4273 3479 4287 3493
rect 4293 3479 4307 3493
rect 4333 3479 4347 3493
rect 4353 3487 4367 3501
rect 4453 3499 4467 3513
rect 4493 3553 4507 3567
rect 4493 3519 4507 3533
rect 4513 3507 4527 3521
rect 4253 3459 4267 3473
rect 4313 3459 4327 3473
rect 4473 3493 4487 3507
rect 4573 3487 4587 3501
rect 4593 3479 4607 3493
rect 4633 3479 4647 3493
rect 4653 3479 4667 3493
rect 4693 3479 4707 3493
rect 4713 3487 4727 3501
rect 4613 3459 4627 3473
rect 4673 3459 4687 3473
rect 53 3296 67 3310
rect 193 3302 207 3316
rect 93 3227 107 3241
rect 133 3227 147 3241
rect 193 3264 207 3278
rect 273 3227 287 3241
rect 293 3219 307 3233
rect 313 3227 327 3241
rect 213 3199 227 3213
rect 53 3170 67 3184
rect 333 3219 347 3233
rect 353 3227 367 3241
rect 373 3239 387 3253
rect 393 3247 407 3261
rect 413 3239 427 3253
rect 513 3247 527 3261
rect 613 3247 627 3261
rect 453 3227 467 3241
rect 473 3219 487 3233
rect 493 3227 507 3241
rect 553 3227 567 3241
rect 573 3219 587 3233
rect 593 3227 607 3241
rect 673 3239 687 3253
rect 693 3247 707 3261
rect 713 3239 727 3253
rect 733 3207 747 3221
rect 753 3219 767 3233
rect 813 3219 827 3233
rect 193 3170 207 3184
rect 953 3219 967 3233
rect 1013 3219 1027 3233
rect 1293 3302 1307 3316
rect 1433 3296 1447 3310
rect 1153 3219 1167 3233
rect 1213 3219 1227 3233
rect 1233 3207 1247 3221
rect 1293 3264 1307 3278
rect 1273 3199 1287 3213
rect 1353 3227 1367 3241
rect 1393 3227 1407 3241
rect 1293 3170 1307 3184
rect 1553 3247 1567 3261
rect 1613 3247 1627 3261
rect 1713 3247 1727 3261
rect 1493 3227 1507 3241
rect 1513 3219 1527 3233
rect 1533 3227 1547 3241
rect 1633 3227 1647 3241
rect 1653 3219 1667 3233
rect 1673 3227 1687 3241
rect 1733 3227 1747 3241
rect 1753 3219 1767 3233
rect 1773 3227 1787 3241
rect 2093 3302 2107 3316
rect 2233 3296 2247 3310
rect 1873 3247 1887 3261
rect 1973 3247 1987 3261
rect 1813 3219 1827 3233
rect 1893 3227 1907 3241
rect 1433 3170 1447 3184
rect 1833 3207 1847 3221
rect 1913 3219 1927 3233
rect 1933 3227 1947 3241
rect 1993 3227 2007 3241
rect 2013 3219 2027 3233
rect 2033 3227 2047 3241
rect 2093 3264 2107 3278
rect 2073 3199 2087 3213
rect 2153 3227 2167 3241
rect 2193 3227 2207 3241
rect 2093 3170 2107 3184
rect 2473 3267 2487 3281
rect 2433 3239 2447 3253
rect 2453 3247 2467 3261
rect 2493 3247 2507 3261
rect 2313 3219 2327 3233
rect 2233 3170 2247 3184
rect 2333 3207 2347 3221
rect 2373 3219 2387 3233
rect 2393 3207 2407 3221
rect 2513 3219 2527 3233
rect 2533 3207 2547 3221
rect 2553 3219 2567 3233
rect 2573 3227 2587 3241
rect 2693 3247 2707 3261
rect 2633 3219 2647 3233
rect 2713 3227 2727 3241
rect 2653 3207 2667 3221
rect 2733 3219 2747 3233
rect 2753 3227 2767 3241
rect 2773 3227 2787 3241
rect 2913 3247 2927 3261
rect 2813 3227 2827 3241
rect 2853 3227 2867 3241
rect 2793 3207 2807 3221
rect 2873 3219 2887 3233
rect 2893 3227 2907 3241
rect 2913 3213 2927 3227
rect 2953 3273 2967 3287
rect 2993 3273 3007 3287
rect 2953 3239 2967 3253
rect 2973 3247 2987 3261
rect 2993 3239 3007 3253
rect 3033 3239 3047 3253
rect 3053 3247 3067 3261
rect 3033 3193 3047 3207
rect 3073 3239 3087 3253
rect 3153 3253 3167 3267
rect 3133 3227 3147 3241
rect 3153 3219 3167 3233
rect 3173 3207 3187 3221
rect 3193 3219 3207 3233
rect 3273 3267 3287 3281
rect 3233 3239 3247 3253
rect 3253 3247 3267 3261
rect 3293 3247 3307 3261
rect 3333 3247 3347 3261
rect 3353 3227 3367 3241
rect 3373 3219 3387 3233
rect 3393 3227 3407 3241
rect 3433 3227 3447 3241
rect 3453 3239 3467 3253
rect 3233 3173 3247 3187
rect 3493 3227 3507 3241
rect 3513 3239 3527 3253
rect 3533 3247 3547 3261
rect 3553 3239 3567 3253
rect 3613 3227 3627 3241
rect 3633 3239 3647 3253
rect 3673 3227 3687 3241
rect 3713 3227 3727 3241
rect 3733 3219 3747 3233
rect 3753 3227 3767 3241
rect 3773 3219 3787 3233
rect 3793 3227 3807 3241
rect 3833 3239 3847 3253
rect 3853 3247 3867 3261
rect 3873 3239 3887 3253
rect 3973 3273 3987 3287
rect 3953 3247 3967 3261
rect 3893 3227 3907 3241
rect 3913 3219 3927 3233
rect 3933 3227 3947 3241
rect 3953 3213 3967 3227
rect 4053 3273 4067 3287
rect 3993 3239 4007 3253
rect 4013 3247 4027 3261
rect 4033 3239 4047 3253
rect 4093 3227 4107 3241
rect 4113 3239 4127 3253
rect 4053 3173 4067 3187
rect 4153 3227 4167 3241
rect 4173 3239 4187 3253
rect 4193 3247 4207 3261
rect 4213 3239 4227 3253
rect 4253 3227 4267 3241
rect 4293 3239 4307 3253
rect 4513 3247 4527 3261
rect 4613 3247 4627 3261
rect 4713 3267 4727 3281
rect 4313 3227 4327 3241
rect 4353 3219 4367 3233
rect 4373 3207 4387 3221
rect 4393 3219 4407 3233
rect 4413 3227 4427 3241
rect 4453 3227 4467 3241
rect 4473 3219 4487 3233
rect 4493 3227 4507 3241
rect 4553 3227 4567 3241
rect 4573 3219 4587 3233
rect 4593 3227 4607 3241
rect 4673 3239 4687 3253
rect 4693 3247 4707 3261
rect 4733 3247 4747 3261
rect 53 3076 67 3090
rect 193 3076 207 3090
rect 93 3019 107 3033
rect 133 3019 147 3033
rect 213 3047 227 3061
rect 473 3076 487 3090
rect 193 2982 207 2996
rect 293 3019 307 3033
rect 313 3027 327 3041
rect 333 3019 347 3033
rect 273 2999 287 3013
rect 373 3007 387 3021
rect 613 3076 627 3090
rect 453 3047 467 3061
rect 393 2999 407 3013
rect 413 3007 427 3021
rect 53 2950 67 2964
rect 193 2944 207 2958
rect 473 2982 487 2996
rect 533 3019 547 3033
rect 573 3019 587 3033
rect 473 2944 487 2958
rect 613 2950 627 2964
rect 713 3076 727 3090
rect 853 3076 867 3090
rect 753 3019 767 3033
rect 793 3019 807 3033
rect 873 3047 887 3061
rect 853 2982 867 2996
rect 913 3039 927 3053
rect 993 3053 1007 3067
rect 933 3027 947 3041
rect 1013 3039 1027 3053
rect 713 2950 727 2964
rect 853 2944 867 2958
rect 993 3019 1007 3033
rect 1033 3019 1047 3033
rect 1073 3007 1087 3021
rect 1093 2999 1107 3013
rect 1113 3007 1127 3021
rect 1133 3019 1147 3033
rect 1153 3027 1167 3041
rect 1173 3019 1187 3033
rect 1233 3027 1247 3041
rect 1253 3039 1267 3053
rect 1273 3027 1287 3041
rect 1373 3076 1387 3090
rect 1293 3019 1307 3033
rect 953 2973 967 2987
rect 1193 2999 1207 3013
rect 1513 3076 1527 3090
rect 1413 3019 1427 3033
rect 1453 3019 1467 3033
rect 1533 3047 1547 3061
rect 1513 2982 1527 2996
rect 1613 3039 1627 3053
rect 1593 3019 1607 3033
rect 1633 3019 1647 3033
rect 1673 3007 1687 3021
rect 1973 3076 1987 3090
rect 2113 3076 2127 3090
rect 1693 2999 1707 3013
rect 1713 3007 1727 3021
rect 1733 3019 1747 3033
rect 1753 3027 1767 3041
rect 1793 3033 1807 3047
rect 1833 3033 1847 3047
rect 1953 3047 1967 3061
rect 1773 3019 1787 3033
rect 1873 3019 1887 3033
rect 1893 3027 1907 3041
rect 1913 3019 1927 3033
rect 1373 2950 1387 2964
rect 1513 2944 1527 2958
rect 1793 2999 1807 3013
rect 1853 2999 1867 3013
rect 1973 2982 1987 2996
rect 2033 3019 2047 3033
rect 2073 3019 2087 3033
rect 2213 3039 2227 3053
rect 2193 3019 2207 3033
rect 2233 3019 2247 3033
rect 2273 3027 2287 3041
rect 2293 3039 2307 3053
rect 1973 2944 1987 2958
rect 2113 2950 2127 2964
rect 2333 3007 2347 3021
rect 2433 3019 2447 3033
rect 2453 3027 2467 3041
rect 2473 3039 2487 3053
rect 2493 3027 2507 3041
rect 2353 2999 2367 3013
rect 2393 2999 2407 3013
rect 2373 2979 2387 2993
rect 2533 3007 2547 3021
rect 2653 3019 2667 3033
rect 2673 3027 2687 3041
rect 2753 3039 2767 3053
rect 2693 3019 2707 3033
rect 2733 3019 2747 3033
rect 2553 2999 2567 3013
rect 2593 2999 2607 3013
rect 2633 2999 2647 3013
rect 2573 2979 2587 2993
rect 2773 3019 2787 3033
rect 2793 3007 2807 3021
rect 2813 2999 2827 3013
rect 2833 3007 2847 3021
rect 2873 3007 2887 3021
rect 2893 2999 2907 3013
rect 2913 3007 2927 3021
rect 2953 3019 2967 3033
rect 2973 3027 2987 3041
rect 2993 3019 3007 3033
rect 3013 3027 3027 3041
rect 3033 3019 3047 3033
rect 3073 3007 3087 3021
rect 3093 2999 3107 3013
rect 3113 3007 3127 3021
rect 3153 3019 3167 3033
rect 3173 3027 3187 3041
rect 3193 3019 3207 3033
rect 3253 3027 3267 3041
rect 3273 3019 3287 3033
rect 3313 3019 3327 3033
rect 3213 2999 3227 3013
rect 3353 3007 3367 3021
rect 3373 3019 3387 3033
rect 3433 3019 3447 3033
rect 3473 3019 3487 3033
rect 3513 3019 3527 3033
rect 3553 3019 3567 3033
rect 3573 3007 3587 3021
rect 3593 2999 3607 3013
rect 3613 3007 3627 3021
rect 3653 3019 3667 3033
rect 3673 3027 3687 3041
rect 3693 3019 3707 3033
rect 3773 3019 3787 3033
rect 3713 2999 3727 3013
rect 3813 3019 3827 3033
rect 3833 3019 3847 3033
rect 3853 3027 3867 3041
rect 3893 3033 3907 3047
rect 3873 3019 3887 3033
rect 3893 2999 3907 3013
rect 3933 2999 3947 3013
rect 3973 2999 3987 3013
rect 3993 3007 4007 3021
rect 4033 3019 4047 3033
rect 3953 2979 3967 2993
rect 3913 2953 3927 2967
rect 4073 3019 4087 3033
rect 4133 3019 4147 3033
rect 4153 3027 4167 3041
rect 4173 3039 4187 3053
rect 4193 3027 4207 3041
rect 4213 3033 4227 3047
rect 4233 3013 4247 3027
rect 4213 2999 4227 3013
rect 4253 2999 4267 3013
rect 4273 3007 4287 3021
rect 4333 3019 4347 3033
rect 4353 3027 4367 3041
rect 4373 3039 4387 3053
rect 4393 3027 4407 3041
rect 4533 3027 4547 3041
rect 4553 3039 4567 3053
rect 4233 2979 4247 2993
rect 4433 3007 4447 3021
rect 4453 2999 4467 3013
rect 4493 2999 4507 3013
rect 4473 2979 4487 2993
rect 4613 3019 4627 3033
rect 4633 3027 4647 3041
rect 4653 3019 4667 3033
rect 4673 3019 4687 3033
rect 4693 3027 4707 3041
rect 4713 3019 4727 3033
rect 4593 2999 4607 3013
rect 4733 2999 4747 3013
rect 53 2816 67 2830
rect 193 2822 207 2836
rect 93 2747 107 2761
rect 133 2747 147 2761
rect 193 2784 207 2798
rect 273 2747 287 2761
rect 293 2739 307 2753
rect 313 2747 327 2761
rect 213 2719 227 2733
rect 53 2690 67 2704
rect 333 2739 347 2753
rect 353 2747 367 2761
rect 373 2759 387 2773
rect 393 2767 407 2781
rect 413 2759 427 2773
rect 473 2767 487 2781
rect 493 2747 507 2761
rect 513 2739 527 2753
rect 533 2747 547 2761
rect 573 2747 587 2761
rect 193 2690 207 2704
rect 613 2747 627 2761
rect 633 2759 647 2773
rect 653 2767 667 2781
rect 673 2759 687 2773
rect 733 2767 747 2781
rect 753 2747 767 2761
rect 773 2739 787 2753
rect 793 2747 807 2761
rect 833 2747 847 2761
rect 873 2747 887 2761
rect 913 2759 927 2773
rect 933 2767 947 2781
rect 853 2727 867 2741
rect 953 2759 967 2773
rect 1053 2759 1067 2773
rect 1073 2767 1087 2781
rect 973 2727 987 2741
rect 993 2739 1007 2753
rect 1093 2759 1107 2773
rect 1113 2747 1127 2761
rect 1313 2816 1327 2830
rect 1453 2822 1467 2836
rect 1153 2747 1167 2761
rect 1213 2747 1227 2761
rect 1133 2727 1147 2741
rect 1253 2747 1267 2761
rect 1353 2747 1367 2761
rect 1393 2747 1407 2761
rect 1453 2784 1467 2798
rect 1513 2759 1527 2773
rect 1533 2767 1547 2781
rect 1473 2719 1487 2733
rect 1313 2690 1327 2704
rect 1553 2759 1567 2773
rect 1613 2767 1627 2781
rect 1713 2767 1727 2781
rect 1633 2747 1647 2761
rect 1653 2739 1667 2753
rect 1673 2747 1687 2761
rect 1733 2747 1747 2761
rect 1753 2739 1767 2753
rect 1773 2747 1787 2761
rect 1813 2747 1827 2761
rect 1853 2747 1867 2761
rect 1893 2747 1907 2761
rect 1833 2727 1847 2741
rect 1453 2690 1467 2704
rect 1913 2739 1927 2753
rect 1933 2727 1947 2741
rect 1953 2739 1967 2753
rect 1993 2747 2007 2761
rect 2113 2787 2127 2801
rect 2273 2816 2287 2830
rect 2413 2822 2427 2836
rect 2033 2747 2047 2761
rect 2073 2759 2087 2773
rect 2093 2767 2107 2781
rect 2133 2767 2147 2781
rect 2153 2747 2167 2761
rect 2193 2747 2207 2761
rect 2313 2747 2327 2761
rect 2353 2747 2367 2761
rect 2413 2784 2427 2798
rect 2493 2767 2507 2781
rect 2593 2767 2607 2781
rect 2893 2793 2907 2807
rect 2733 2767 2747 2781
rect 2433 2719 2447 2733
rect 2513 2747 2527 2761
rect 2533 2739 2547 2753
rect 2553 2747 2567 2761
rect 2613 2747 2627 2761
rect 2633 2739 2647 2753
rect 2653 2747 2667 2761
rect 2673 2747 2687 2761
rect 2693 2739 2707 2753
rect 2713 2747 2727 2761
rect 2753 2753 2767 2767
rect 2773 2759 2787 2773
rect 2793 2767 2807 2781
rect 2733 2733 2747 2747
rect 2273 2690 2287 2704
rect 2413 2690 2427 2704
rect 2813 2759 2827 2773
rect 2853 2759 2867 2773
rect 2873 2767 2887 2781
rect 2893 2759 2907 2773
rect 2993 2767 3007 2781
rect 3093 2767 3107 2781
rect 2933 2747 2947 2761
rect 2953 2739 2967 2753
rect 2973 2747 2987 2761
rect 3033 2747 3047 2761
rect 2933 2713 2947 2727
rect 3053 2739 3067 2753
rect 3073 2747 3087 2761
rect 3133 2759 3147 2773
rect 3153 2767 3167 2781
rect 3173 2759 3187 2773
rect 3233 2767 3247 2781
rect 3413 2787 3427 2801
rect 3253 2747 3267 2761
rect 3273 2739 3287 2753
rect 3293 2747 3307 2761
rect 3333 2759 3347 2773
rect 3353 2767 3367 2781
rect 3373 2759 3387 2773
rect 3393 2767 3407 2781
rect 3433 2767 3447 2781
rect 3493 2813 3507 2827
rect 3453 2759 3467 2773
rect 3513 2767 3527 2781
rect 3653 2767 3667 2781
rect 3533 2747 3547 2761
rect 3513 2733 3527 2747
rect 3553 2739 3567 2753
rect 3573 2747 3587 2761
rect 3593 2747 3607 2761
rect 3613 2739 3627 2753
rect 3633 2747 3647 2761
rect 3673 2713 3687 2727
rect 3713 2793 3727 2807
rect 3753 2793 3767 2807
rect 3713 2759 3727 2773
rect 3733 2767 3747 2781
rect 3753 2759 3767 2773
rect 3753 2713 3767 2727
rect 3793 2767 3807 2781
rect 3893 2787 3907 2801
rect 3873 2767 3887 2781
rect 3913 2767 3927 2781
rect 3813 2747 3827 2761
rect 3833 2739 3847 2753
rect 3853 2747 3867 2761
rect 3933 2759 3947 2773
rect 4033 2773 4047 2787
rect 3973 2727 3987 2741
rect 3993 2739 4007 2753
rect 4173 2787 4187 2801
rect 4153 2767 4167 2781
rect 4193 2767 4207 2781
rect 4053 2747 4067 2761
rect 4073 2739 4087 2753
rect 4093 2747 4107 2761
rect 4053 2713 4067 2727
rect 4113 2739 4127 2753
rect 4133 2747 4147 2761
rect 4213 2759 4227 2773
rect 4233 2753 4247 2767
rect 4313 2767 4327 2781
rect 4253 2747 4267 2761
rect 4273 2739 4287 2753
rect 4293 2747 4307 2761
rect 4353 2747 4367 2761
rect 4253 2713 4267 2727
rect 4393 2759 4407 2773
rect 4413 2747 4427 2761
rect 4453 2747 4467 2761
rect 4473 2739 4487 2753
rect 4493 2747 4507 2761
rect 4513 2739 4527 2753
rect 4533 2747 4547 2761
rect 4753 2773 4767 2787
rect 4573 2727 4587 2741
rect 4593 2739 4607 2753
rect 4633 2739 4647 2753
rect 4653 2727 4667 2741
rect 4673 2739 4687 2753
rect 4693 2747 4707 2761
rect 4713 2693 4727 2707
rect 53 2596 67 2610
rect 193 2596 207 2610
rect 93 2539 107 2553
rect 133 2539 147 2553
rect 213 2567 227 2581
rect 193 2502 207 2516
rect 293 2539 307 2553
rect 313 2547 327 2561
rect 333 2539 347 2553
rect 353 2539 367 2553
rect 273 2519 287 2533
rect 393 2539 407 2553
rect 53 2470 67 2484
rect 193 2464 207 2478
rect 433 2527 447 2541
rect 453 2519 467 2533
rect 473 2527 487 2541
rect 553 2539 567 2553
rect 573 2547 587 2561
rect 593 2539 607 2553
rect 613 2539 627 2553
rect 533 2519 547 2533
rect 653 2539 667 2553
rect 733 2539 747 2553
rect 753 2547 767 2561
rect 813 2559 827 2573
rect 773 2539 787 2553
rect 793 2539 807 2553
rect 713 2519 727 2533
rect 913 2596 927 2610
rect 833 2539 847 2553
rect 1053 2596 1067 2610
rect 953 2539 967 2553
rect 993 2539 1007 2553
rect 1073 2567 1087 2581
rect 1053 2502 1067 2516
rect 1113 2559 1127 2573
rect 1133 2547 1147 2561
rect 913 2470 927 2484
rect 1053 2464 1067 2478
rect 1173 2539 1187 2553
rect 1193 2547 1207 2561
rect 1273 2559 1287 2573
rect 1453 2596 1467 2610
rect 1213 2539 1227 2553
rect 1293 2547 1307 2561
rect 1233 2519 1247 2533
rect 1333 2527 1347 2541
rect 1593 2596 1607 2610
rect 1433 2567 1447 2581
rect 1353 2519 1367 2533
rect 1373 2527 1387 2541
rect 1453 2502 1467 2516
rect 1513 2539 1527 2553
rect 1553 2539 1567 2553
rect 1793 2596 1807 2610
rect 1933 2596 1947 2610
rect 2233 2596 2247 2610
rect 1653 2539 1667 2553
rect 1673 2547 1687 2561
rect 1693 2539 1707 2553
rect 1773 2567 1787 2581
rect 1713 2519 1727 2533
rect 1453 2464 1467 2478
rect 1593 2470 1607 2484
rect 1793 2502 1807 2516
rect 1853 2539 1867 2553
rect 1893 2539 1907 2553
rect 2013 2547 2027 2561
rect 2153 2547 2167 2561
rect 2373 2596 2387 2610
rect 2273 2539 2287 2553
rect 2313 2539 2327 2553
rect 1793 2464 1807 2478
rect 1933 2470 1947 2484
rect 2393 2567 2407 2581
rect 2373 2502 2387 2516
rect 2453 2527 2467 2541
rect 2513 2559 2527 2573
rect 2533 2547 2547 2561
rect 2473 2519 2487 2533
rect 2493 2527 2507 2541
rect 2233 2470 2247 2484
rect 2373 2464 2387 2478
rect 2613 2539 2627 2553
rect 2633 2547 2647 2561
rect 2673 2559 2687 2573
rect 2653 2539 2667 2553
rect 2693 2547 2707 2561
rect 2593 2519 2607 2533
rect 2753 2527 2767 2541
rect 2773 2519 2787 2533
rect 2793 2527 2807 2541
rect 2853 2539 2867 2553
rect 2873 2547 2887 2561
rect 2893 2539 2907 2553
rect 2913 2539 2927 2553
rect 2833 2519 2847 2533
rect 2953 2527 2967 2541
rect 2973 2539 2987 2553
rect 3013 2539 3027 2553
rect 3033 2547 3047 2561
rect 3053 2539 3067 2553
rect 3073 2519 3087 2533
rect 3133 2527 3147 2541
rect 3153 2519 3167 2533
rect 3173 2527 3187 2541
rect 3193 2539 3207 2553
rect 3233 2527 3247 2541
rect 3253 2539 3267 2553
rect 3393 2559 3407 2573
rect 3413 2547 3427 2561
rect 3313 2527 3327 2541
rect 3333 2519 3347 2533
rect 3373 2519 3387 2533
rect 3353 2499 3367 2513
rect 3453 2527 3467 2541
rect 3473 2519 3487 2533
rect 3493 2527 3507 2541
rect 3533 2539 3547 2553
rect 3573 2527 3587 2541
rect 3593 2539 3607 2553
rect 3633 2539 3647 2553
rect 3713 2559 3727 2573
rect 3673 2539 3687 2553
rect 3733 2547 3747 2561
rect 3793 2539 3807 2553
rect 3813 2527 3827 2541
rect 3853 2539 3867 2553
rect 3893 2539 3907 2553
rect 3913 2547 3927 2561
rect 3973 2573 3987 2587
rect 3933 2539 3947 2553
rect 3953 2547 3967 2561
rect 3973 2539 3987 2553
rect 3993 2533 4007 2547
rect 4013 2527 4027 2541
rect 4033 2519 4047 2533
rect 4053 2527 4067 2541
rect 4093 2527 4107 2541
rect 4113 2519 4127 2533
rect 4133 2527 4147 2541
rect 4153 2539 4167 2553
rect 4173 2547 4187 2561
rect 4193 2539 4207 2553
rect 4213 2519 4227 2533
rect 4253 2527 4267 2541
rect 4533 2547 4547 2561
rect 4553 2559 4567 2573
rect 4573 2547 4587 2561
rect 4273 2519 4287 2533
rect 4293 2527 4307 2541
rect 4353 2527 4367 2541
rect 4373 2519 4387 2533
rect 4413 2519 4427 2533
rect 4453 2527 4467 2541
rect 4593 2539 4607 2553
rect 4393 2499 4407 2513
rect 4473 2519 4487 2533
rect 4513 2519 4527 2533
rect 4493 2499 4507 2513
rect 4653 2527 4667 2541
rect 4673 2519 4687 2533
rect 4713 2519 4727 2533
rect 4693 2499 4707 2513
rect 53 2336 67 2350
rect 193 2342 207 2356
rect 93 2267 107 2281
rect 133 2267 147 2281
rect 193 2304 207 2318
rect 313 2287 327 2301
rect 253 2267 267 2281
rect 273 2259 287 2273
rect 293 2267 307 2281
rect 353 2267 367 2281
rect 213 2239 227 2253
rect 373 2259 387 2273
rect 393 2267 407 2281
rect 53 2210 67 2224
rect 193 2210 207 2224
rect 413 2259 427 2273
rect 433 2267 447 2281
rect 473 2267 487 2281
rect 513 2267 527 2281
rect 553 2279 567 2293
rect 573 2287 587 2301
rect 593 2279 607 2293
rect 653 2259 667 2273
rect 693 2267 707 2281
rect 733 2267 747 2281
rect 793 2267 807 2281
rect 673 2247 687 2261
rect 713 2247 727 2261
rect 813 2259 827 2273
rect 833 2247 847 2261
rect 853 2259 867 2273
rect 873 2267 887 2281
rect 913 2267 927 2281
rect 953 2267 967 2281
rect 993 2267 1007 2281
rect 1133 2342 1147 2356
rect 1273 2336 1287 2350
rect 893 2247 907 2261
rect 973 2247 987 2261
rect 1033 2247 1047 2261
rect 1053 2259 1067 2273
rect 1133 2304 1147 2318
rect 1113 2239 1127 2253
rect 1473 2342 1487 2356
rect 1613 2336 1627 2350
rect 1193 2267 1207 2281
rect 1233 2267 1247 2281
rect 1133 2210 1147 2224
rect 1393 2287 1407 2301
rect 1333 2267 1347 2281
rect 1353 2259 1367 2273
rect 1373 2267 1387 2281
rect 1473 2304 1487 2318
rect 1273 2210 1287 2224
rect 1453 2239 1467 2253
rect 2333 2336 2347 2350
rect 2473 2342 2487 2356
rect 1533 2267 1547 2281
rect 1573 2267 1587 2281
rect 1473 2210 1487 2224
rect 1693 2267 1707 2281
rect 1613 2210 1627 2224
rect 1733 2267 1747 2281
rect 1773 2267 1787 2281
rect 1713 2247 1727 2261
rect 1793 2259 1807 2273
rect 1813 2247 1827 2261
rect 1833 2259 1847 2273
rect 1853 2259 1867 2273
rect 1873 2267 1887 2281
rect 1933 2267 1947 2281
rect 1973 2267 1987 2281
rect 1953 2247 1967 2261
rect 2013 2259 2027 2273
rect 2253 2287 2267 2301
rect 2153 2259 2167 2273
rect 2193 2267 2207 2281
rect 2213 2259 2227 2273
rect 2233 2267 2247 2281
rect 2373 2267 2387 2281
rect 2413 2267 2427 2281
rect 2473 2304 2487 2318
rect 3013 2336 3027 2350
rect 3153 2342 3167 2356
rect 2553 2279 2567 2293
rect 2573 2287 2587 2301
rect 2493 2239 2507 2253
rect 2333 2210 2347 2224
rect 2593 2279 2607 2293
rect 2613 2279 2627 2293
rect 2633 2287 2647 2301
rect 2473 2210 2487 2224
rect 2653 2279 2667 2293
rect 2693 2279 2707 2293
rect 2713 2287 2727 2301
rect 2733 2279 2747 2293
rect 2793 2287 2807 2301
rect 2893 2287 2907 2301
rect 2813 2267 2827 2281
rect 2833 2259 2847 2273
rect 2853 2267 2867 2281
rect 2913 2267 2927 2281
rect 2933 2259 2947 2273
rect 2953 2267 2967 2281
rect 3053 2267 3067 2281
rect 3093 2267 3107 2281
rect 3153 2304 3167 2318
rect 3273 2333 3287 2347
rect 3273 2287 3287 2301
rect 3213 2267 3227 2281
rect 3233 2259 3247 2273
rect 3253 2267 3267 2281
rect 3173 2239 3187 2253
rect 3273 2253 3287 2267
rect 3313 2279 3327 2293
rect 3333 2287 3347 2301
rect 3013 2210 3027 2224
rect 3153 2210 3167 2224
rect 3353 2279 3367 2293
rect 3393 2279 3407 2293
rect 3413 2287 3427 2301
rect 3433 2279 3447 2293
rect 3493 2279 3507 2293
rect 3513 2287 3527 2301
rect 3533 2279 3547 2293
rect 3573 2267 3587 2281
rect 3593 2259 3607 2273
rect 3633 2267 3647 2281
rect 3793 2287 3807 2301
rect 3653 2259 3667 2273
rect 3693 2259 3707 2273
rect 3733 2267 3747 2281
rect 3713 2247 3727 2261
rect 3753 2259 3767 2273
rect 3773 2267 3787 2281
rect 3853 2267 3867 2281
rect 3893 2267 3907 2281
rect 3913 2259 3927 2273
rect 3933 2267 3947 2281
rect 3973 2267 3987 2281
rect 4013 2279 4027 2293
rect 4093 2287 4107 2301
rect 4233 2307 4247 2321
rect 4033 2267 4047 2281
rect 4113 2267 4127 2281
rect 4133 2259 4147 2273
rect 4153 2267 4167 2281
rect 4193 2279 4207 2293
rect 4213 2287 4227 2301
rect 4253 2287 4267 2301
rect 4393 2287 4407 2301
rect 4533 2287 4547 2301
rect 4593 2287 4607 2301
rect 4173 2253 4187 2267
rect 4153 2233 4167 2247
rect 4273 2259 4287 2273
rect 4293 2247 4307 2261
rect 4313 2259 4327 2273
rect 4333 2267 4347 2281
rect 4413 2267 4427 2281
rect 4433 2259 4447 2273
rect 4453 2267 4467 2281
rect 4473 2267 4487 2281
rect 4493 2259 4507 2273
rect 4513 2267 4527 2281
rect 4613 2267 4627 2281
rect 4633 2259 4647 2273
rect 4653 2267 4667 2281
rect 4673 2259 4687 2273
rect 4693 2247 4707 2261
rect 4713 2259 4727 2273
rect 4733 2267 4747 2281
rect 33 2067 47 2081
rect 173 2067 187 2081
rect 233 2047 247 2061
rect 553 2116 567 2130
rect 253 2039 267 2053
rect 273 2047 287 2061
rect 313 2073 327 2087
rect 333 2059 347 2073
rect 353 2067 367 2081
rect 373 2059 387 2073
rect 393 2059 407 2073
rect 413 2067 427 2081
rect 433 2059 447 2073
rect 453 2067 467 2081
rect 473 2059 487 2073
rect 313 2039 327 2053
rect 693 2116 707 2130
rect 593 2059 607 2073
rect 633 2059 647 2073
rect 313 1993 327 2007
rect 713 2087 727 2101
rect 693 2022 707 2036
rect 773 2047 787 2061
rect 853 2067 867 2081
rect 793 2039 807 2053
rect 813 2047 827 2061
rect 553 1990 567 2004
rect 693 1984 707 1998
rect 913 2079 927 2093
rect 893 2059 907 2073
rect 933 2047 947 2061
rect 1033 2079 1047 2093
rect 953 2039 967 2053
rect 973 2047 987 2061
rect 1013 2059 1027 2073
rect 1053 2059 1067 2073
rect 1093 2059 1107 2073
rect 1113 2067 1127 2081
rect 1133 2059 1147 2073
rect 1153 2039 1167 2053
rect 1193 2047 1207 2061
rect 1293 2079 1307 2093
rect 1213 2039 1227 2053
rect 1233 2047 1247 2061
rect 1273 2059 1287 2073
rect 1393 2116 1407 2130
rect 1533 2116 1547 2130
rect 1373 2087 1387 2101
rect 1313 2059 1327 2073
rect 1393 2022 1407 2036
rect 1453 2059 1467 2073
rect 1493 2059 1507 2073
rect 1613 2059 1627 2073
rect 1633 2067 1647 2081
rect 1653 2079 1667 2093
rect 1673 2067 1687 2081
rect 1813 2116 1827 2130
rect 1713 2059 1727 2073
rect 1953 2116 1967 2130
rect 1793 2087 1807 2101
rect 1753 2059 1767 2073
rect 1393 1984 1407 1998
rect 1533 1990 1547 2004
rect 1813 2022 1827 2036
rect 1873 2059 1887 2073
rect 1913 2059 1927 2073
rect 2033 2067 2047 2081
rect 2053 2079 2067 2093
rect 1813 1984 1827 1998
rect 1953 1990 1967 2004
rect 2093 2047 2107 2061
rect 2113 2039 2127 2053
rect 2133 2047 2147 2061
rect 2153 2059 2167 2073
rect 2193 2059 2207 2073
rect 2233 2047 2247 2061
rect 2253 2039 2267 2053
rect 2273 2047 2287 2061
rect 2353 2059 2367 2073
rect 2373 2067 2387 2081
rect 2393 2059 2407 2073
rect 2333 2039 2347 2053
rect 2433 2047 2447 2061
rect 2473 2093 2487 2107
rect 2453 2039 2467 2053
rect 2473 2047 2487 2061
rect 2513 2047 2527 2061
rect 2813 2116 2827 2130
rect 2533 2039 2547 2053
rect 2553 2047 2567 2061
rect 2613 2059 2627 2073
rect 2633 2067 2647 2081
rect 2653 2059 2667 2073
rect 2713 2059 2727 2073
rect 2733 2067 2747 2081
rect 2753 2059 2767 2073
rect 2593 2039 2607 2053
rect 2513 2013 2527 2027
rect 2693 2039 2707 2053
rect 2953 2116 2967 2130
rect 2853 2059 2867 2073
rect 2893 2059 2907 2073
rect 2973 2087 2987 2101
rect 2953 2022 2967 2036
rect 3013 2059 3027 2073
rect 2813 1990 2827 2004
rect 2953 1984 2967 1998
rect 3053 2047 3067 2061
rect 3073 2059 3087 2073
rect 3133 2073 3147 2087
rect 3153 2059 3167 2073
rect 3173 2067 3187 2081
rect 3193 2059 3207 2073
rect 3253 2059 3267 2073
rect 3273 2067 3287 2081
rect 3293 2059 3307 2073
rect 3133 2039 3147 2053
rect 3113 2013 3127 2027
rect 3233 2039 3247 2053
rect 3313 2047 3327 2061
rect 3373 2073 3387 2087
rect 3333 2039 3347 2053
rect 3353 2047 3367 2061
rect 3353 2013 3367 2027
rect 3433 2059 3447 2073
rect 3453 2067 3467 2081
rect 3473 2059 3487 2073
rect 3593 2079 3607 2093
rect 3613 2067 3627 2081
rect 3413 2039 3427 2053
rect 3493 2039 3507 2053
rect 3533 2039 3547 2053
rect 3553 2047 3567 2061
rect 3513 2019 3527 2033
rect 3653 2073 3667 2087
rect 3653 2039 3667 2053
rect 3693 2039 3707 2053
rect 3713 2047 3727 2061
rect 3753 2047 3767 2061
rect 3673 2019 3687 2033
rect 3633 1993 3647 2007
rect 3773 2039 3787 2053
rect 3793 2047 3807 2061
rect 3833 2059 3847 2073
rect 3873 2059 3887 2073
rect 3913 2059 3927 2073
rect 3933 2067 3947 2081
rect 3953 2059 3967 2073
rect 3973 2039 3987 2053
rect 4033 2047 4047 2061
rect 4053 2039 4067 2053
rect 4073 2047 4087 2061
rect 4113 2047 4127 2061
rect 4153 2093 4167 2107
rect 4133 2039 4147 2053
rect 4153 2047 4167 2061
rect 3973 1993 3987 2007
rect 3993 1993 4007 2007
rect 4033 1993 4047 2007
rect 4153 2013 4167 2027
rect 4193 2047 4207 2061
rect 4213 2039 4227 2053
rect 4233 2047 4247 2061
rect 4253 2059 4267 2073
rect 4293 2047 4307 2061
rect 4313 2059 4327 2073
rect 4353 2067 4367 2081
rect 4373 2079 4387 2093
rect 4393 2067 4407 2081
rect 4413 2059 4427 2073
rect 4473 2059 4487 2073
rect 4493 2067 4507 2081
rect 4513 2079 4527 2093
rect 4533 2067 4547 2081
rect 4553 2039 4567 2053
rect 4593 2039 4607 2053
rect 4613 2047 4627 2061
rect 4573 2019 4587 2033
rect 4653 2039 4667 2053
rect 4693 2039 4707 2053
rect 4713 2047 4727 2061
rect 4673 2019 4687 2033
rect 53 1856 67 1870
rect 193 1862 207 1876
rect 93 1787 107 1801
rect 133 1787 147 1801
rect 193 1824 207 1838
rect 313 1807 327 1821
rect 253 1787 267 1801
rect 273 1779 287 1793
rect 293 1787 307 1801
rect 213 1759 227 1773
rect 313 1773 327 1787
rect 373 1853 387 1867
rect 373 1807 387 1821
rect 473 1807 487 1821
rect 573 1807 587 1821
rect 393 1787 407 1801
rect 413 1779 427 1793
rect 433 1787 447 1801
rect 493 1787 507 1801
rect 513 1779 527 1793
rect 533 1787 547 1801
rect 593 1787 607 1801
rect 613 1779 627 1793
rect 633 1787 647 1801
rect 653 1767 667 1781
rect 673 1779 687 1793
rect 53 1730 67 1744
rect 193 1730 207 1744
rect 713 1767 727 1781
rect 733 1779 747 1793
rect 793 1787 807 1801
rect 873 1827 887 1841
rect 853 1807 867 1821
rect 893 1807 907 1821
rect 993 1856 1007 1870
rect 1133 1862 1147 1876
rect 833 1787 847 1801
rect 913 1799 927 1813
rect 813 1767 827 1781
rect 1033 1787 1047 1801
rect 1073 1787 1087 1801
rect 1133 1824 1147 1838
rect 1613 1856 1627 1870
rect 1753 1862 1767 1876
rect 1193 1799 1207 1813
rect 1213 1807 1227 1821
rect 1153 1759 1167 1773
rect 993 1730 1007 1744
rect 1233 1799 1247 1813
rect 1293 1807 1307 1821
rect 1313 1787 1327 1801
rect 1333 1779 1347 1793
rect 1353 1787 1367 1801
rect 1393 1779 1407 1793
rect 1533 1779 1547 1793
rect 1133 1730 1147 1744
rect 1653 1787 1667 1801
rect 1693 1787 1707 1801
rect 1753 1824 1767 1838
rect 2313 1862 2327 1876
rect 2453 1856 2467 1870
rect 1833 1787 1847 1801
rect 1773 1759 1787 1773
rect 1613 1730 1627 1744
rect 1753 1730 1767 1744
rect 1853 1779 1867 1793
rect 1873 1767 1887 1781
rect 1893 1779 1907 1793
rect 1913 1787 1927 1801
rect 1953 1787 1967 1801
rect 2013 1787 2027 1801
rect 1933 1767 1947 1781
rect 2033 1779 2047 1793
rect 2053 1767 2067 1781
rect 2073 1779 2087 1793
rect 2113 1787 2127 1801
rect 2153 1787 2167 1801
rect 2133 1767 2147 1781
rect 2173 1779 2187 1793
rect 2193 1767 2207 1781
rect 2213 1779 2227 1793
rect 2233 1787 2247 1801
rect 2313 1824 2327 1838
rect 2293 1759 2307 1773
rect 2373 1787 2387 1801
rect 2413 1787 2427 1801
rect 2313 1730 2327 1744
rect 2453 1730 2467 1744
rect 2553 1856 2567 1870
rect 2693 1862 2707 1876
rect 2593 1787 2607 1801
rect 2633 1787 2647 1801
rect 2693 1824 2707 1838
rect 2713 1759 2727 1773
rect 2553 1730 2567 1744
rect 2693 1730 2707 1744
rect 2793 1856 2807 1870
rect 2933 1862 2947 1876
rect 2833 1787 2847 1801
rect 2873 1787 2887 1801
rect 2933 1824 2947 1838
rect 3013 1787 3027 1801
rect 3073 1799 3087 1813
rect 3093 1807 3107 1821
rect 2953 1759 2967 1773
rect 2793 1730 2807 1744
rect 3033 1779 3047 1793
rect 3113 1799 3127 1813
rect 3173 1813 3187 1827
rect 3213 1813 3227 1827
rect 3153 1787 3167 1801
rect 3173 1779 3187 1793
rect 3193 1779 3207 1793
rect 3213 1767 3227 1781
rect 3233 1779 3247 1793
rect 3253 1787 3267 1801
rect 3293 1787 3307 1801
rect 3333 1787 3347 1801
rect 3393 1787 3407 1801
rect 3413 1799 3427 1813
rect 3313 1767 3327 1781
rect 2933 1730 2947 1744
rect 3453 1787 3467 1801
rect 3473 1779 3487 1793
rect 3493 1787 3507 1801
rect 3553 1787 3567 1801
rect 3573 1779 3587 1793
rect 3593 1787 3607 1801
rect 3613 1779 3627 1793
rect 3633 1787 3647 1801
rect 3673 1787 3687 1801
rect 3693 1779 3707 1793
rect 3733 1787 3747 1801
rect 3773 1787 3787 1801
rect 3793 1787 3807 1801
rect 3753 1767 3767 1781
rect 3833 1787 3847 1801
rect 3873 1787 3887 1801
rect 3913 1799 3927 1813
rect 3933 1787 3947 1801
rect 3993 1787 4007 1801
rect 4013 1779 4027 1793
rect 4033 1787 4047 1801
rect 4053 1779 4067 1793
rect 4073 1787 4087 1801
rect 4093 1787 4107 1801
rect 4113 1779 4127 1793
rect 4133 1787 4147 1801
rect 4153 1779 4167 1793
rect 4173 1787 4187 1801
rect 4213 1799 4227 1813
rect 4233 1807 4247 1821
rect 4253 1799 4267 1813
rect 4293 1787 4307 1801
rect 4333 1799 4347 1813
rect 4353 1787 4367 1801
rect 4393 1787 4407 1801
rect 4413 1779 4427 1793
rect 4433 1787 4447 1801
rect 4453 1779 4467 1793
rect 4473 1787 4487 1801
rect 4633 1807 4647 1821
rect 4533 1779 4547 1793
rect 4573 1787 4587 1801
rect 4553 1767 4567 1781
rect 4593 1779 4607 1793
rect 4613 1787 4627 1801
rect 4653 1793 4667 1807
rect 4633 1773 4647 1787
rect 4673 1767 4687 1781
rect 4693 1779 4707 1793
rect 33 1587 47 1601
rect 173 1587 187 1601
rect 253 1599 267 1613
rect 233 1579 247 1593
rect 413 1636 427 1650
rect 273 1579 287 1593
rect 313 1579 327 1593
rect 353 1579 367 1593
rect 553 1636 567 1650
rect 453 1579 467 1593
rect 493 1579 507 1593
rect 573 1607 587 1621
rect 553 1542 567 1556
rect 413 1510 427 1524
rect 553 1504 567 1518
rect 653 1636 667 1650
rect 793 1636 807 1650
rect 693 1579 707 1593
rect 733 1579 747 1593
rect 813 1607 827 1621
rect 793 1542 807 1556
rect 653 1510 667 1524
rect 793 1504 807 1518
rect 893 1636 907 1650
rect 1033 1636 1047 1650
rect 873 1607 887 1621
rect 893 1542 907 1556
rect 953 1579 967 1593
rect 993 1579 1007 1593
rect 1113 1567 1127 1581
rect 1313 1636 1327 1650
rect 1453 1636 1467 1650
rect 1293 1607 1307 1621
rect 1133 1559 1147 1573
rect 1153 1567 1167 1581
rect 1213 1579 1227 1593
rect 1233 1587 1247 1601
rect 1253 1579 1267 1593
rect 1193 1559 1207 1573
rect 893 1504 907 1518
rect 1033 1510 1047 1524
rect 1313 1542 1327 1556
rect 1373 1579 1387 1593
rect 1413 1579 1427 1593
rect 1313 1504 1327 1518
rect 1453 1510 1467 1524
rect 1553 1636 1567 1650
rect 1693 1636 1707 1650
rect 1593 1579 1607 1593
rect 1633 1579 1647 1593
rect 1713 1607 1727 1621
rect 1693 1542 1707 1556
rect 1773 1579 1787 1593
rect 1793 1587 1807 1601
rect 1813 1599 1827 1613
rect 1833 1587 1847 1601
rect 1873 1599 1887 1613
rect 1853 1579 1867 1593
rect 1973 1636 1987 1650
rect 1893 1579 1907 1593
rect 2113 1636 2127 1650
rect 2013 1579 2027 1593
rect 2053 1579 2067 1593
rect 1553 1510 1567 1524
rect 1693 1504 1707 1518
rect 2133 1607 2147 1621
rect 2113 1542 2127 1556
rect 2473 1636 2487 1650
rect 2213 1599 2227 1613
rect 2193 1579 2207 1593
rect 2233 1579 2247 1593
rect 2273 1567 2287 1581
rect 2613 1636 2627 1650
rect 2293 1559 2307 1573
rect 2313 1567 2327 1581
rect 2333 1579 2347 1593
rect 2353 1587 2367 1601
rect 2373 1579 2387 1593
rect 2453 1607 2467 1621
rect 1973 1510 1987 1524
rect 2113 1504 2127 1518
rect 2393 1559 2407 1573
rect 2473 1542 2487 1556
rect 2533 1579 2547 1593
rect 2573 1579 2587 1593
rect 2473 1504 2487 1518
rect 2613 1510 2627 1524
rect 2713 1636 2727 1650
rect 2853 1636 2867 1650
rect 2753 1579 2767 1593
rect 2793 1579 2807 1593
rect 2873 1607 2887 1621
rect 2853 1542 2867 1556
rect 2913 1587 2927 1601
rect 2933 1579 2947 1593
rect 2973 1567 2987 1581
rect 2993 1559 3007 1573
rect 3013 1567 3027 1581
rect 3073 1567 3087 1581
rect 3093 1559 3107 1573
rect 3113 1567 3127 1581
rect 3133 1579 3147 1593
rect 3153 1587 3167 1601
rect 3173 1579 3187 1593
rect 2713 1510 2727 1524
rect 2853 1504 2867 1518
rect 3193 1559 3207 1573
rect 3233 1567 3247 1581
rect 3313 1613 3327 1627
rect 3253 1559 3267 1573
rect 3273 1567 3287 1581
rect 3333 1567 3347 1581
rect 3373 1613 3387 1627
rect 3353 1559 3367 1573
rect 3373 1567 3387 1581
rect 3333 1533 3347 1547
rect 3433 1579 3447 1593
rect 3453 1587 3467 1601
rect 3473 1579 3487 1593
rect 3413 1559 3427 1573
rect 3493 1559 3507 1573
rect 3533 1559 3547 1573
rect 3553 1567 3567 1581
rect 3613 1579 3627 1593
rect 3633 1587 3647 1601
rect 3653 1579 3667 1593
rect 3673 1587 3687 1601
rect 3713 1599 3727 1613
rect 3693 1579 3707 1593
rect 3733 1587 3747 1601
rect 3393 1513 3407 1527
rect 3513 1539 3527 1553
rect 3873 1587 3887 1601
rect 3893 1599 3907 1613
rect 3913 1587 3927 1601
rect 3773 1559 3787 1573
rect 3813 1559 3827 1573
rect 3833 1567 3847 1581
rect 3933 1579 3947 1593
rect 3973 1579 3987 1593
rect 3993 1587 4007 1601
rect 4013 1579 4027 1593
rect 3793 1539 3807 1553
rect 4033 1559 4047 1573
rect 4093 1567 4107 1581
rect 4153 1587 4167 1601
rect 4173 1599 4187 1613
rect 4193 1587 4207 1601
rect 4113 1559 4127 1573
rect 4133 1567 4147 1581
rect 4213 1579 4227 1593
rect 4253 1579 4267 1593
rect 4273 1587 4287 1601
rect 4353 1599 4367 1613
rect 4293 1579 4307 1593
rect 4373 1587 4387 1601
rect 4433 1599 4447 1613
rect 4313 1559 4327 1573
rect 4413 1579 4427 1593
rect 4453 1579 4467 1593
rect 4493 1567 4507 1581
rect 4513 1559 4527 1573
rect 4533 1567 4547 1581
rect 4573 1567 4587 1581
rect 4633 1613 4647 1627
rect 4593 1559 4607 1573
rect 4613 1567 4627 1581
rect 4613 1533 4627 1547
rect 4653 1567 4667 1581
rect 4673 1559 4687 1573
rect 4693 1567 4707 1581
rect 53 1382 67 1396
rect 193 1376 207 1390
rect 53 1344 67 1358
rect 33 1279 47 1293
rect 113 1307 127 1321
rect 153 1307 167 1321
rect 53 1250 67 1264
rect 193 1250 207 1264
rect 293 1376 307 1390
rect 433 1382 447 1396
rect 333 1307 347 1321
rect 373 1307 387 1321
rect 433 1344 447 1358
rect 493 1319 507 1333
rect 513 1327 527 1341
rect 453 1279 467 1293
rect 293 1250 307 1264
rect 533 1319 547 1333
rect 593 1327 607 1341
rect 693 1327 707 1341
rect 613 1307 627 1321
rect 633 1299 647 1313
rect 653 1307 667 1321
rect 713 1307 727 1321
rect 733 1299 747 1313
rect 753 1307 767 1321
rect 793 1307 807 1321
rect 433 1250 447 1264
rect 833 1307 847 1321
rect 853 1319 867 1333
rect 873 1327 887 1341
rect 893 1319 907 1333
rect 953 1327 967 1341
rect 973 1307 987 1321
rect 993 1299 1007 1313
rect 1013 1307 1027 1321
rect 1053 1299 1067 1313
rect 1113 1307 1127 1321
rect 1153 1307 1167 1321
rect 1233 1319 1247 1333
rect 1253 1327 1267 1341
rect 1073 1287 1087 1301
rect 1273 1319 1287 1333
rect 1313 1327 1327 1341
rect 1333 1307 1347 1321
rect 1353 1299 1367 1313
rect 1373 1307 1387 1321
rect 1413 1319 1427 1333
rect 1433 1327 1447 1341
rect 1453 1319 1467 1333
rect 1493 1327 1507 1341
rect 1513 1307 1527 1321
rect 1533 1299 1547 1313
rect 1553 1307 1567 1321
rect 1573 1307 1587 1321
rect 1873 1382 1887 1396
rect 2013 1376 2027 1390
rect 1613 1307 1627 1321
rect 1653 1319 1667 1333
rect 1673 1327 1687 1341
rect 1693 1319 1707 1333
rect 1753 1327 1767 1341
rect 1773 1307 1787 1321
rect 1793 1299 1807 1313
rect 1813 1307 1827 1321
rect 1873 1344 1887 1358
rect 1853 1279 1867 1293
rect 1933 1307 1947 1321
rect 1973 1307 1987 1321
rect 1873 1250 1887 1264
rect 2193 1327 2207 1341
rect 2073 1287 2087 1301
rect 2093 1299 2107 1313
rect 2133 1307 2147 1321
rect 2153 1299 2167 1313
rect 2173 1307 2187 1321
rect 2253 1319 2267 1333
rect 2273 1327 2287 1341
rect 2013 1250 2027 1264
rect 2293 1319 2307 1333
rect 2333 1307 2347 1321
rect 2373 1307 2387 1321
rect 2573 1382 2587 1396
rect 2713 1376 2727 1390
rect 2353 1287 2367 1301
rect 2413 1299 2427 1313
rect 2453 1307 2467 1321
rect 2493 1307 2507 1321
rect 2433 1287 2447 1301
rect 2473 1287 2487 1301
rect 2573 1344 2587 1358
rect 2553 1279 2567 1293
rect 2633 1307 2647 1321
rect 2673 1307 2687 1321
rect 2573 1250 2587 1264
rect 2773 1307 2787 1321
rect 2973 1327 2987 1341
rect 3073 1327 3087 1341
rect 3173 1327 3187 1341
rect 2813 1307 2827 1321
rect 2873 1307 2887 1321
rect 2793 1287 2807 1301
rect 2713 1250 2727 1264
rect 2893 1299 2907 1313
rect 2913 1307 2927 1321
rect 2933 1299 2947 1313
rect 2953 1307 2967 1321
rect 3013 1307 3027 1321
rect 3033 1299 3047 1313
rect 3053 1307 3067 1321
rect 3113 1307 3127 1321
rect 3133 1299 3147 1313
rect 3153 1307 3167 1321
rect 3213 1307 3227 1321
rect 3253 1319 3267 1333
rect 3273 1307 3287 1321
rect 3333 1307 3347 1321
rect 3413 1347 3427 1361
rect 3393 1327 3407 1341
rect 3433 1327 3447 1341
rect 3373 1307 3387 1321
rect 3453 1319 3467 1333
rect 3513 1327 3527 1341
rect 3653 1327 3667 1341
rect 3353 1287 3367 1301
rect 3533 1307 3547 1321
rect 3553 1299 3567 1313
rect 3573 1307 3587 1321
rect 3593 1307 3607 1321
rect 3613 1299 3627 1313
rect 3633 1307 3647 1321
rect 3713 1319 3727 1333
rect 3733 1327 3747 1341
rect 3753 1319 3767 1333
rect 3793 1319 3807 1333
rect 3813 1327 3827 1341
rect 3833 1319 3847 1333
rect 3853 1307 3867 1321
rect 3893 1319 3907 1333
rect 3973 1327 3987 1341
rect 3913 1307 3927 1321
rect 3993 1307 4007 1321
rect 4013 1299 4027 1313
rect 4033 1307 4047 1321
rect 4353 1373 4367 1387
rect 4133 1319 4147 1333
rect 4153 1327 4167 1341
rect 4053 1287 4067 1301
rect 4073 1299 4087 1313
rect 4173 1319 4187 1333
rect 4213 1319 4227 1333
rect 4233 1327 4247 1341
rect 4253 1319 4267 1333
rect 4293 1307 4307 1321
rect 4333 1307 4347 1321
rect 4313 1287 4327 1301
rect 4333 1273 4347 1287
rect 4373 1327 4387 1341
rect 4513 1327 4527 1341
rect 4393 1307 4407 1321
rect 4413 1299 4427 1313
rect 4433 1307 4447 1321
rect 4453 1307 4467 1321
rect 4473 1299 4487 1313
rect 4493 1307 4507 1321
rect 4573 1307 4587 1321
rect 4653 1319 4667 1333
rect 4673 1327 4687 1341
rect 4593 1299 4607 1313
rect 4613 1287 4627 1301
rect 4633 1299 4647 1313
rect 4693 1319 4707 1333
rect 13 1119 27 1133
rect 33 1107 47 1121
rect 93 1087 107 1101
rect 113 1079 127 1093
rect 133 1087 147 1101
rect 173 1113 187 1127
rect 193 1099 207 1113
rect 213 1107 227 1121
rect 233 1099 247 1113
rect 253 1099 267 1113
rect 273 1107 287 1121
rect 293 1099 307 1113
rect 313 1107 327 1121
rect 333 1099 347 1113
rect 393 1099 407 1113
rect 413 1107 427 1121
rect 433 1119 447 1133
rect 453 1107 467 1121
rect 493 1107 507 1121
rect 173 1079 187 1093
rect 173 1033 187 1047
rect 553 1119 567 1133
rect 593 1119 607 1133
rect 533 1099 547 1113
rect 573 1099 587 1113
rect 613 1099 627 1113
rect 673 1099 687 1113
rect 693 1087 707 1101
rect 733 1099 747 1113
rect 773 1099 787 1113
rect 873 1119 887 1133
rect 813 1099 827 1113
rect 853 1099 867 1113
rect 893 1099 907 1113
rect 933 1107 947 1121
rect 953 1119 967 1133
rect 993 1107 1007 1121
rect 1013 1119 1027 1133
rect 1053 1119 1067 1133
rect 1113 1119 1127 1133
rect 1033 1099 1047 1113
rect 1073 1099 1087 1113
rect 1133 1107 1147 1121
rect 1213 1119 1227 1133
rect 1193 1099 1207 1113
rect 1233 1099 1247 1113
rect 1253 1107 1267 1121
rect 1273 1119 1287 1133
rect 1293 1107 1307 1121
rect 1393 1156 1407 1170
rect 1313 1099 1327 1113
rect 1533 1156 1547 1170
rect 1433 1099 1447 1113
rect 1473 1099 1487 1113
rect 1553 1127 1567 1141
rect 1533 1062 1547 1076
rect 1613 1107 1627 1121
rect 1633 1119 1647 1133
rect 1393 1030 1407 1044
rect 1533 1024 1547 1038
rect 1653 1087 1667 1101
rect 1753 1119 1767 1133
rect 1673 1079 1687 1093
rect 1693 1087 1707 1101
rect 1733 1099 1747 1113
rect 1853 1156 1867 1170
rect 1773 1099 1787 1113
rect 1993 1156 2007 1170
rect 1893 1099 1907 1113
rect 1933 1099 1947 1113
rect 2013 1127 2027 1141
rect 1993 1062 2007 1076
rect 2073 1107 2087 1121
rect 2093 1119 2107 1133
rect 2133 1119 2147 1133
rect 2213 1119 2227 1133
rect 2373 1156 2387 1170
rect 2513 1156 2527 1170
rect 1853 1030 1867 1044
rect 1993 1024 2007 1038
rect 2113 1099 2127 1113
rect 2153 1099 2167 1113
rect 2193 1099 2207 1113
rect 2233 1099 2247 1113
rect 2293 1107 2307 1121
rect 2313 1119 2327 1133
rect 2353 1127 2367 1141
rect 2373 1062 2387 1076
rect 2433 1099 2447 1113
rect 2473 1099 2487 1113
rect 2573 1119 2587 1133
rect 2593 1107 2607 1121
rect 2373 1024 2387 1038
rect 2513 1030 2527 1044
rect 2633 1099 2647 1113
rect 2653 1107 2667 1121
rect 2693 1113 2707 1127
rect 2673 1099 2687 1113
rect 2693 1079 2707 1093
rect 2733 1099 2747 1113
rect 2753 1107 2767 1121
rect 2773 1099 2787 1113
rect 2793 1107 2807 1121
rect 2873 1119 2887 1133
rect 2813 1099 2827 1113
rect 2853 1099 2867 1113
rect 2713 1053 2727 1067
rect 2893 1099 2907 1113
rect 2953 1087 2967 1101
rect 2973 1079 2987 1093
rect 2993 1087 3007 1101
rect 3013 1099 3027 1113
rect 3053 1087 3067 1101
rect 3073 1099 3087 1113
rect 3113 1099 3127 1113
rect 3133 1107 3147 1121
rect 3173 1113 3187 1127
rect 3213 1119 3227 1133
rect 3153 1099 3167 1113
rect 3173 1079 3187 1093
rect 3173 1033 3187 1047
rect 3233 1099 3247 1113
rect 3273 1107 3287 1121
rect 3333 1087 3347 1101
rect 3353 1079 3367 1093
rect 3373 1087 3387 1101
rect 3413 1087 3427 1101
rect 3433 1079 3447 1093
rect 3453 1087 3467 1101
rect 3473 1087 3487 1101
rect 3533 1133 3547 1147
rect 3493 1079 3507 1093
rect 3513 1087 3527 1101
rect 3513 1053 3527 1067
rect 3553 1087 3567 1101
rect 3573 1079 3587 1093
rect 3593 1087 3607 1101
rect 3633 1099 3647 1113
rect 3653 1107 3667 1121
rect 3673 1099 3687 1113
rect 3833 1107 3847 1121
rect 3853 1119 3867 1133
rect 3873 1107 3887 1121
rect 3693 1079 3707 1093
rect 3753 1087 3767 1101
rect 3893 1099 3907 1113
rect 3953 1107 3967 1121
rect 3973 1119 3987 1133
rect 3773 1079 3787 1093
rect 3813 1079 3827 1093
rect 3793 1059 3807 1073
rect 4093 1107 4107 1121
rect 4113 1119 4127 1133
rect 4133 1107 4147 1121
rect 4193 1119 4207 1133
rect 4013 1087 4027 1101
rect 4153 1099 4167 1113
rect 4213 1107 4227 1121
rect 4033 1079 4047 1093
rect 4073 1079 4087 1093
rect 4053 1059 4067 1073
rect 4273 1099 4287 1113
rect 4293 1107 4307 1121
rect 4313 1119 4327 1133
rect 4333 1107 4347 1121
rect 4393 1099 4407 1113
rect 4413 1107 4427 1121
rect 4433 1099 4447 1113
rect 4453 1099 4467 1113
rect 4473 1107 4487 1121
rect 4573 1119 4587 1133
rect 4493 1099 4507 1113
rect 4553 1099 4567 1113
rect 4373 1079 4387 1093
rect 4513 1079 4527 1093
rect 4593 1099 4607 1113
rect 4653 1087 4667 1101
rect 4693 1133 4707 1147
rect 4673 1079 4687 1093
rect 4693 1087 4707 1101
rect 4733 1107 4747 1121
rect 4753 1119 4767 1133
rect 4713 1073 4727 1087
rect 53 896 67 910
rect 193 902 207 916
rect 93 827 107 841
rect 133 827 147 841
rect 193 864 207 878
rect 473 896 487 910
rect 613 902 627 916
rect 253 839 267 853
rect 273 847 287 861
rect 213 799 227 813
rect 53 770 67 784
rect 293 839 307 853
rect 353 847 367 861
rect 373 827 387 841
rect 393 819 407 833
rect 413 827 427 841
rect 193 770 207 784
rect 513 827 527 841
rect 553 827 567 841
rect 613 864 627 878
rect 673 839 687 853
rect 693 847 707 861
rect 633 799 647 813
rect 473 770 487 784
rect 713 839 727 853
rect 773 847 787 861
rect 873 847 887 861
rect 793 827 807 841
rect 813 819 827 833
rect 833 827 847 841
rect 893 827 907 841
rect 913 819 927 833
rect 933 827 947 841
rect 973 819 987 833
rect 1033 827 1047 841
rect 1073 827 1087 841
rect 1093 827 1107 841
rect 1133 827 1147 841
rect 1193 839 1207 853
rect 1213 847 1227 861
rect 613 770 627 784
rect 993 807 1007 821
rect 1053 807 1067 821
rect 1113 807 1127 821
rect 1233 839 1247 853
rect 1273 839 1287 853
rect 1293 847 1307 861
rect 1313 839 1327 853
rect 1353 839 1367 853
rect 1373 847 1387 861
rect 1393 839 1407 853
rect 1433 827 1447 841
rect 1453 819 1467 833
rect 1473 807 1487 821
rect 1493 819 1507 833
rect 1533 827 1547 841
rect 1553 839 1567 853
rect 1593 827 1607 841
rect 1613 819 1627 833
rect 1633 807 1647 821
rect 1653 819 1667 833
rect 1673 827 1687 841
rect 1733 819 1747 833
rect 1933 839 1947 853
rect 1953 847 1967 861
rect 1873 819 1887 833
rect 1973 839 1987 853
rect 2013 827 2027 841
rect 2133 847 2147 861
rect 2233 847 2247 861
rect 2333 847 2347 861
rect 2053 827 2067 841
rect 2073 827 2087 841
rect 2033 807 2047 821
rect 2093 819 2107 833
rect 2113 827 2127 841
rect 2173 827 2187 841
rect 2193 819 2207 833
rect 2213 827 2227 841
rect 2273 827 2287 841
rect 2293 819 2307 833
rect 2313 827 2327 841
rect 2373 839 2387 853
rect 2393 847 2407 861
rect 2413 839 2427 853
rect 2553 902 2567 916
rect 2693 896 2707 910
rect 2473 819 2487 833
rect 2493 807 2507 821
rect 2553 864 2567 878
rect 2533 799 2547 813
rect 2613 827 2627 841
rect 2653 827 2667 841
rect 2553 770 2567 784
rect 2773 847 2787 861
rect 2793 827 2807 841
rect 2813 819 2827 833
rect 2833 827 2847 841
rect 2993 867 3007 881
rect 2973 847 2987 861
rect 3013 847 3027 861
rect 3033 839 3047 853
rect 2873 819 2887 833
rect 2693 770 2707 784
rect 2893 807 2907 821
rect 2913 807 2927 821
rect 2933 819 2947 833
rect 3293 893 3307 907
rect 3153 839 3167 853
rect 3173 847 3187 861
rect 3073 807 3087 821
rect 3093 819 3107 833
rect 3193 839 3207 853
rect 3233 827 3247 841
rect 3213 807 3227 821
rect 3273 819 3287 833
rect 3313 839 3327 853
rect 3333 847 3347 861
rect 3313 793 3327 807
rect 3353 839 3367 853
rect 3393 839 3407 853
rect 3413 847 3427 861
rect 3433 839 3447 853
rect 3493 827 3507 841
rect 3533 827 3547 841
rect 3553 839 3567 853
rect 3573 847 3587 861
rect 3693 867 3707 881
rect 3513 807 3527 821
rect 3593 839 3607 853
rect 3653 839 3667 853
rect 3673 847 3687 861
rect 3713 847 3727 861
rect 3793 867 3807 881
rect 3913 873 3927 887
rect 3753 839 3767 853
rect 3773 847 3787 861
rect 3813 847 3827 861
rect 3833 839 3847 853
rect 3853 847 3867 861
rect 3873 839 3887 853
rect 3993 893 4007 907
rect 3973 867 3987 881
rect 3933 839 3947 853
rect 3953 847 3967 861
rect 3993 847 4007 861
rect 4013 833 4027 847
rect 4173 893 4187 907
rect 4093 847 4107 861
rect 4033 819 4047 833
rect 4113 827 4127 841
rect 3933 773 3947 787
rect 4053 807 4067 821
rect 4133 819 4147 833
rect 4153 827 4167 841
rect 4193 847 4207 861
rect 4273 853 4287 867
rect 4213 827 4227 841
rect 4173 813 4187 827
rect 4233 819 4247 833
rect 4253 827 4267 841
rect 4393 867 4407 881
rect 4373 847 4387 861
rect 4413 847 4427 861
rect 4473 893 4487 907
rect 4293 827 4307 841
rect 4433 839 4447 853
rect 4273 793 4287 807
rect 4313 819 4327 833
rect 4333 807 4347 821
rect 4353 819 4367 833
rect 4533 867 4547 881
rect 4493 839 4507 853
rect 4513 847 4527 861
rect 4553 847 4567 861
rect 4693 867 4707 881
rect 4673 847 4687 861
rect 4713 847 4727 861
rect 4593 827 4607 841
rect 4733 839 4747 853
rect 4473 793 4487 807
rect 4613 819 4627 833
rect 4633 807 4647 821
rect 4653 819 4667 833
rect 53 676 67 690
rect 193 676 207 690
rect 93 619 107 633
rect 133 619 147 633
rect 213 647 227 661
rect 193 582 207 596
rect 253 639 267 653
rect 273 627 287 641
rect 53 550 67 564
rect 193 544 207 558
rect 313 619 327 633
rect 333 627 347 641
rect 353 619 367 633
rect 373 599 387 613
rect 413 607 427 621
rect 433 599 447 613
rect 453 607 467 621
rect 493 619 507 633
rect 673 676 687 690
rect 813 676 827 690
rect 533 619 547 633
rect 593 627 607 641
rect 613 639 627 653
rect 653 647 667 661
rect 673 582 687 596
rect 733 619 747 633
rect 773 619 787 633
rect 873 619 887 633
rect 893 627 907 641
rect 1013 639 1027 653
rect 1053 639 1067 653
rect 913 619 927 633
rect 993 619 1007 633
rect 933 599 947 613
rect 1033 619 1047 633
rect 1073 619 1087 633
rect 1113 627 1127 641
rect 673 544 687 558
rect 813 550 827 564
rect 1193 619 1207 633
rect 1213 627 1227 641
rect 1233 619 1247 633
rect 1273 619 1287 633
rect 1173 599 1187 613
rect 1293 607 1307 621
rect 1553 676 1567 690
rect 1373 639 1387 653
rect 1333 619 1347 633
rect 1353 619 1367 633
rect 1393 619 1407 633
rect 1433 619 1447 633
rect 1473 619 1487 633
rect 1693 676 1707 690
rect 1593 619 1607 633
rect 1633 619 1647 633
rect 1713 647 1727 661
rect 1693 582 1707 596
rect 1753 619 1767 633
rect 1873 639 1887 653
rect 1953 639 1967 653
rect 1793 619 1807 633
rect 1853 619 1867 633
rect 1553 550 1567 564
rect 1693 544 1707 558
rect 1893 619 1907 633
rect 1933 619 1947 633
rect 1973 619 1987 633
rect 2013 627 2027 641
rect 2033 639 2047 653
rect 2073 639 2087 653
rect 2053 619 2067 633
rect 2173 676 2187 690
rect 2313 676 2327 690
rect 2153 647 2167 661
rect 2093 619 2107 633
rect 2173 582 2187 596
rect 2233 619 2247 633
rect 2273 619 2287 633
rect 2373 619 2387 633
rect 2393 627 2407 641
rect 2413 619 2427 633
rect 2433 627 2447 641
rect 2453 619 2467 633
rect 2513 627 2527 641
rect 2173 544 2187 558
rect 2313 550 2327 564
rect 2573 639 2587 653
rect 2553 619 2567 633
rect 2613 619 2627 633
rect 2633 627 2647 641
rect 2653 639 2667 653
rect 2673 627 2687 641
rect 2713 619 2727 633
rect 2733 627 2747 641
rect 2753 639 2767 653
rect 2773 627 2787 641
rect 2793 639 2807 653
rect 2813 627 2827 641
rect 2893 619 2907 633
rect 2913 627 2927 641
rect 2933 619 2947 633
rect 2953 619 2967 633
rect 2973 627 2987 641
rect 2993 619 3007 633
rect 2873 599 2887 613
rect 3013 599 3027 613
rect 3053 607 3067 621
rect 3153 627 3167 641
rect 3173 639 3187 653
rect 3193 639 3207 653
rect 3213 627 3227 641
rect 3073 599 3087 613
rect 3093 607 3107 621
rect 3393 639 3407 653
rect 3273 607 3287 621
rect 3373 619 3387 633
rect 3293 599 3307 613
rect 3333 599 3347 613
rect 3313 579 3327 593
rect 3413 619 3427 633
rect 3433 619 3447 633
rect 3453 627 3467 641
rect 3493 633 3507 647
rect 3473 619 3487 633
rect 3493 599 3507 613
rect 3533 627 3547 641
rect 3553 639 3567 653
rect 3573 627 3587 641
rect 3593 619 3607 633
rect 3653 619 3667 633
rect 3673 627 3687 641
rect 3693 639 3707 653
rect 3713 627 3727 641
rect 3753 619 3767 633
rect 3773 627 3787 641
rect 3793 619 3807 633
rect 3813 627 3827 641
rect 3833 619 3847 633
rect 4053 639 4067 653
rect 4073 627 4087 641
rect 3553 593 3567 607
rect 3873 607 3887 621
rect 3893 599 3907 613
rect 3933 599 3947 613
rect 3973 607 3987 621
rect 3913 579 3927 593
rect 3993 599 4007 613
rect 4033 599 4047 613
rect 4013 579 4027 593
rect 4513 639 4527 653
rect 4533 627 4547 641
rect 4113 599 4127 613
rect 4153 599 4167 613
rect 4173 607 4187 621
rect 4133 579 4147 593
rect 4213 599 4227 613
rect 4253 599 4267 613
rect 4273 607 4287 621
rect 4333 607 4347 621
rect 4233 579 4247 593
rect 4313 593 4327 607
rect 4293 573 4307 587
rect 4353 599 4367 613
rect 4393 599 4407 613
rect 4433 607 4447 621
rect 4373 579 4387 593
rect 4453 599 4467 613
rect 4493 599 4507 613
rect 4473 579 4487 593
rect 4613 619 4627 633
rect 4633 627 4647 641
rect 4653 619 4667 633
rect 4673 619 4687 633
rect 4693 627 4707 641
rect 4713 619 4727 633
rect 4593 599 4607 613
rect 4733 599 4747 613
rect 53 416 67 430
rect 193 422 207 436
rect 93 347 107 361
rect 133 347 147 361
rect 193 384 207 398
rect 253 359 267 373
rect 273 367 287 381
rect 213 319 227 333
rect 53 290 67 304
rect 293 359 307 373
rect 353 367 367 381
rect 373 347 387 361
rect 393 339 407 353
rect 413 347 427 361
rect 493 359 507 373
rect 513 367 527 381
rect 433 327 447 341
rect 453 339 467 353
rect 193 290 207 304
rect 533 359 547 373
rect 593 367 607 381
rect 753 393 767 407
rect 733 367 747 381
rect 613 347 627 361
rect 633 339 647 353
rect 653 347 667 361
rect 673 347 687 361
rect 693 339 707 353
rect 713 347 727 361
rect 733 333 747 347
rect 833 367 847 381
rect 893 367 907 381
rect 773 347 787 361
rect 793 339 807 353
rect 813 347 827 361
rect 913 347 927 361
rect 933 339 947 353
rect 953 347 967 361
rect 1033 359 1047 373
rect 1053 367 1067 381
rect 973 327 987 341
rect 993 339 1007 353
rect 1073 359 1087 373
rect 1133 347 1147 361
rect 1293 367 1307 381
rect 1153 339 1167 353
rect 1173 327 1187 341
rect 1193 339 1207 353
rect 1233 339 1247 353
rect 1313 347 1327 361
rect 1253 327 1267 341
rect 1333 339 1347 353
rect 1353 347 1367 361
rect 1393 347 1407 361
rect 1673 422 1687 436
rect 1813 416 1827 430
rect 1513 367 1527 381
rect 1433 347 1447 361
rect 1453 347 1467 361
rect 1413 327 1427 341
rect 1473 339 1487 353
rect 1493 347 1507 361
rect 1553 359 1567 373
rect 1573 367 1587 381
rect 1593 359 1607 373
rect 1673 384 1687 398
rect 1653 319 1667 333
rect 1733 347 1747 361
rect 1773 347 1787 361
rect 1673 290 1687 304
rect 2093 416 2107 430
rect 2233 422 2247 436
rect 1893 359 1907 373
rect 1913 367 1927 381
rect 1933 359 1947 373
rect 1973 367 1987 381
rect 1993 347 2007 361
rect 2013 339 2027 353
rect 2033 347 2047 361
rect 1813 290 1827 304
rect 2133 347 2147 361
rect 2173 347 2187 361
rect 2233 384 2247 398
rect 2313 339 2327 353
rect 2353 347 2367 361
rect 2393 347 2407 361
rect 2613 422 2627 436
rect 2753 416 2767 430
rect 2513 359 2527 373
rect 2533 367 2547 381
rect 2253 319 2267 333
rect 2093 290 2107 304
rect 2233 290 2247 304
rect 2333 327 2347 341
rect 2373 327 2387 341
rect 2433 327 2447 341
rect 2453 339 2467 353
rect 2553 359 2567 373
rect 2613 384 2627 398
rect 2593 319 2607 333
rect 2673 347 2687 361
rect 2713 347 2727 361
rect 2613 290 2627 304
rect 2813 359 2827 373
rect 2833 367 2847 381
rect 2853 359 2867 373
rect 2893 347 2907 361
rect 2913 339 2927 353
rect 2933 347 2947 361
rect 2953 339 2967 353
rect 2973 347 2987 361
rect 3013 347 3027 361
rect 3053 347 3067 361
rect 3213 387 3227 401
rect 3173 359 3187 373
rect 3193 367 3207 381
rect 3233 367 3247 381
rect 3313 387 3327 401
rect 3273 359 3287 373
rect 3293 367 3307 381
rect 3333 367 3347 381
rect 3413 367 3427 381
rect 3033 327 3047 341
rect 3093 327 3107 341
rect 3113 339 3127 353
rect 2753 290 2767 304
rect 3353 347 3367 361
rect 3373 339 3387 353
rect 3393 347 3407 361
rect 3633 393 3647 407
rect 3513 359 3527 373
rect 3533 367 3547 381
rect 3473 339 3487 353
rect 3493 327 3507 341
rect 3553 359 3567 373
rect 3593 359 3607 373
rect 3613 367 3627 381
rect 3633 359 3647 373
rect 3733 367 3747 381
rect 3673 347 3687 361
rect 3693 339 3707 353
rect 3713 347 3727 361
rect 3793 347 3807 361
rect 3653 313 3667 327
rect 3833 347 3847 361
rect 3873 347 3887 361
rect 3913 347 3927 361
rect 3933 347 3947 361
rect 3813 327 3827 341
rect 3893 327 3907 341
rect 3973 359 3987 373
rect 3993 347 4007 361
rect 4033 347 4047 361
rect 4273 387 4287 401
rect 4073 347 4087 361
rect 4133 347 4147 361
rect 4233 359 4247 373
rect 4253 367 4267 381
rect 4293 367 4307 381
rect 4053 327 4067 341
rect 4153 339 4167 353
rect 4173 327 4187 341
rect 4193 339 4207 353
rect 4313 339 4327 353
rect 4333 327 4347 341
rect 4353 339 4367 353
rect 4373 347 4387 361
rect 4493 367 4507 381
rect 4413 327 4427 341
rect 4433 339 4447 353
rect 4513 347 4527 361
rect 4533 339 4547 353
rect 4553 347 4567 361
rect 4573 327 4587 341
rect 4593 339 4607 353
rect 4633 327 4647 341
rect 4653 339 4667 353
rect 4693 327 4707 341
rect 4713 339 4727 353
rect 53 196 67 210
rect 193 196 207 210
rect 93 139 107 153
rect 133 139 147 153
rect 213 167 227 181
rect 193 102 207 116
rect 253 139 267 153
rect 273 147 287 161
rect 293 139 307 153
rect 313 147 327 161
rect 393 159 407 173
rect 333 139 347 153
rect 373 139 387 153
rect 413 139 427 153
rect 793 196 807 210
rect 573 147 587 161
rect 453 119 467 133
rect 493 119 507 133
rect 513 127 527 141
rect 53 70 67 84
rect 193 64 207 78
rect 473 99 487 113
rect 633 159 647 173
rect 613 139 627 153
rect 933 196 947 210
rect 673 139 687 153
rect 693 147 707 161
rect 713 159 727 173
rect 773 167 787 181
rect 733 147 747 161
rect 793 102 807 116
rect 853 139 867 153
rect 893 139 907 153
rect 1033 139 1047 153
rect 1053 147 1067 161
rect 1073 139 1087 153
rect 1113 147 1127 161
rect 1133 159 1147 173
rect 1193 159 1207 173
rect 1013 119 1027 133
rect 793 64 807 78
rect 933 70 947 84
rect 1173 139 1187 153
rect 1213 139 1227 153
rect 1253 147 1267 161
rect 1273 159 1287 173
rect 1333 139 1347 153
rect 1353 147 1367 161
rect 1373 139 1387 153
rect 1413 147 1427 161
rect 1433 159 1447 173
rect 1473 147 1487 161
rect 1493 159 1507 173
rect 1533 159 1547 173
rect 1313 119 1327 133
rect 1513 139 1527 153
rect 1733 196 1747 210
rect 1553 139 1567 153
rect 1613 139 1627 153
rect 1633 147 1647 161
rect 1653 159 1667 173
rect 1673 147 1687 161
rect 1873 196 1887 210
rect 1773 139 1787 153
rect 1813 139 1827 153
rect 1893 167 1907 181
rect 1873 102 1887 116
rect 1973 139 1987 153
rect 1993 147 2007 161
rect 2033 159 2047 173
rect 2013 139 2027 153
rect 2053 147 2067 161
rect 2113 159 2127 173
rect 2193 159 2207 173
rect 1953 119 1967 133
rect 1733 70 1747 84
rect 1873 64 1887 78
rect 2093 139 2107 153
rect 2133 139 2147 153
rect 2173 139 2187 153
rect 2293 159 2307 173
rect 2353 159 2367 173
rect 2513 196 2527 210
rect 2653 196 2667 210
rect 2213 139 2227 153
rect 2273 139 2287 153
rect 2313 139 2327 153
rect 2333 139 2347 153
rect 2373 139 2387 153
rect 2433 147 2447 161
rect 2453 159 2467 173
rect 2493 167 2507 181
rect 2513 102 2527 116
rect 2573 139 2587 153
rect 2613 139 2627 153
rect 2513 64 2527 78
rect 2653 70 2667 84
rect 2753 196 2767 210
rect 2893 196 2907 210
rect 2733 167 2747 181
rect 2753 102 2767 116
rect 2813 139 2827 153
rect 2853 139 2867 153
rect 2953 139 2967 153
rect 2973 147 2987 161
rect 2993 139 3007 153
rect 3013 147 3027 161
rect 3033 139 3047 153
rect 3093 147 3107 161
rect 2753 64 2767 78
rect 2893 70 2907 84
rect 3153 159 3167 173
rect 3133 139 3147 153
rect 3173 139 3187 153
rect 3193 147 3207 161
rect 3213 139 3227 153
rect 3293 147 3307 161
rect 3313 159 3327 173
rect 3233 119 3247 133
rect 3333 127 3347 141
rect 3533 147 3547 161
rect 3553 159 3567 173
rect 3353 119 3367 133
rect 3373 127 3387 141
rect 3433 127 3447 141
rect 3453 119 3467 133
rect 3493 119 3507 133
rect 3473 99 3487 113
rect 3593 139 3607 153
rect 3613 147 3627 161
rect 3633 159 3647 173
rect 3653 147 3667 161
rect 3713 159 3727 173
rect 3753 159 3767 173
rect 3693 139 3707 153
rect 3733 139 3747 153
rect 3773 147 3787 161
rect 3813 139 3827 153
rect 3833 147 3847 161
rect 3933 159 3947 173
rect 3853 139 3867 153
rect 3913 139 3927 153
rect 3873 119 3887 133
rect 3953 139 3967 153
rect 4013 127 4027 141
rect 4033 119 4047 133
rect 4073 119 4087 133
rect 4093 127 4107 141
rect 4113 119 4127 133
rect 4133 127 4147 141
rect 4193 127 4207 141
rect 4053 99 4067 113
rect 4213 119 4227 133
rect 4253 119 4267 133
rect 4293 127 4307 141
rect 4313 119 4327 133
rect 4333 127 4347 141
rect 4373 127 4387 141
rect 4233 99 4247 113
rect 4393 119 4407 133
rect 4433 119 4447 133
rect 4453 127 4467 141
rect 4473 119 4487 133
rect 4493 127 4507 141
rect 4533 119 4547 133
rect 4573 119 4587 133
rect 4593 127 4607 141
rect 4653 139 4667 153
rect 4673 147 4687 161
rect 4693 159 4707 173
rect 4713 147 4727 161
rect 4413 99 4427 113
rect 4553 99 4567 113
<< metal2 >>
rect 36 4487 43 4623
rect 316 4487 323 4573
rect 496 4567 503 4623
rect 536 4587 543 4623
rect 556 4616 583 4623
rect 2756 4616 2783 4623
rect 33 4473 47 4487
rect 73 4483 87 4487
rect 73 4476 103 4483
rect 73 4473 87 4476
rect 96 4223 103 4476
rect 113 4433 127 4447
rect 153 4433 167 4447
rect 233 4453 247 4467
rect 273 4483 287 4487
rect 273 4476 303 4483
rect 273 4473 287 4476
rect 236 4447 243 4453
rect 116 4407 123 4433
rect 156 4427 163 4433
rect 156 4227 163 4393
rect 96 4216 123 4223
rect 33 4193 47 4207
rect 36 4127 43 4193
rect 53 4173 67 4187
rect 93 4173 107 4187
rect 16 3963 23 4013
rect 56 4007 63 4173
rect 96 4147 103 4173
rect 33 3963 47 3967
rect 16 3956 47 3963
rect 33 3953 47 3956
rect 96 3943 103 4113
rect 116 4007 123 4216
rect 176 4187 183 4213
rect 276 4207 283 4413
rect 193 4173 207 4187
rect 196 4167 203 4173
rect 256 4167 263 4173
rect 233 4153 247 4167
rect 236 4147 243 4153
rect 276 4127 283 4193
rect 153 3963 167 3967
rect 176 3963 183 4093
rect 196 4007 203 4113
rect 216 4027 223 4093
rect 213 4013 227 4027
rect 256 4007 263 4053
rect 296 4047 303 4476
rect 313 4473 327 4487
rect 373 4483 387 4487
rect 356 4476 387 4483
rect 416 4487 423 4513
rect 336 4247 343 4453
rect 356 4447 363 4476
rect 373 4473 387 4476
rect 436 4443 443 4553
rect 456 4487 463 4493
rect 453 4473 467 4487
rect 496 4487 503 4493
rect 556 4487 563 4616
rect 493 4473 507 4487
rect 513 4483 527 4487
rect 513 4476 543 4483
rect 513 4473 527 4476
rect 416 4436 443 4443
rect 393 4173 407 4187
rect 353 4153 367 4167
rect 356 4107 363 4153
rect 396 4107 403 4173
rect 296 4007 303 4013
rect 233 4003 247 4007
rect 253 4003 267 4007
rect 233 3996 267 4003
rect 233 3993 247 3996
rect 253 3993 267 3996
rect 293 3993 307 4007
rect 153 3956 183 3963
rect 153 3953 167 3956
rect 76 3936 103 3943
rect 16 3723 23 3933
rect 76 3727 83 3936
rect 216 3827 223 3973
rect 217 3758 225 3782
rect 33 3723 47 3727
rect 16 3716 47 3723
rect 33 3713 47 3716
rect 133 3723 147 3727
rect 93 3703 107 3707
rect 116 3716 147 3723
rect 116 3703 123 3716
rect 93 3696 123 3703
rect 133 3713 147 3716
rect 193 3703 207 3707
rect 93 3693 107 3696
rect 153 3683 167 3687
rect 176 3696 207 3703
rect 176 3683 183 3696
rect 153 3676 183 3683
rect 193 3693 207 3696
rect 153 3673 167 3676
rect 16 2507 23 3673
rect 56 3444 64 3556
rect 133 3523 147 3527
rect 156 3523 163 3613
rect 133 3516 163 3523
rect 133 3513 147 3516
rect 56 3184 64 3296
rect 56 2964 64 3076
rect 116 3047 123 3293
rect 133 3223 147 3227
rect 156 3223 163 3516
rect 133 3216 163 3223
rect 133 3213 147 3216
rect 136 3107 143 3213
rect 136 3047 143 3093
rect 133 3033 147 3047
rect 176 3023 183 3676
rect 217 3664 225 3744
rect 195 3476 203 3556
rect 213 3513 227 3527
rect 216 3487 223 3513
rect 195 3438 203 3462
rect 195 3278 203 3302
rect 195 3184 203 3264
rect 216 3227 223 3253
rect 213 3213 227 3227
rect 156 3016 183 3023
rect 36 2287 43 2873
rect 56 2704 64 2816
rect 93 2733 107 2747
rect 96 2707 103 2733
rect 56 2484 64 2596
rect 96 2567 103 2613
rect 116 2567 123 2973
rect 156 2787 163 3016
rect 195 2996 203 3076
rect 213 3033 227 3047
rect 133 2733 147 2747
rect 136 2567 143 2733
rect 93 2553 107 2567
rect 133 2563 147 2567
rect 133 2556 163 2563
rect 133 2553 147 2556
rect 76 2467 83 2513
rect 96 2447 103 2513
rect 16 2247 23 2273
rect 56 2224 64 2336
rect 116 2243 123 2553
rect 133 2263 147 2267
rect 156 2263 163 2556
rect 133 2256 163 2263
rect 133 2253 147 2256
rect 116 2236 143 2243
rect 16 1583 23 2053
rect 56 1987 63 2093
rect 56 1744 64 1856
rect 93 1783 107 1787
rect 116 1783 123 2073
rect 136 1967 143 2236
rect 156 2167 163 2256
rect 176 2183 183 2993
rect 195 2958 203 2982
rect 216 2863 223 3033
rect 236 2887 243 3933
rect 256 3307 263 3813
rect 273 3693 287 3707
rect 276 3627 283 3693
rect 273 3473 287 3487
rect 276 3467 283 3473
rect 256 3147 263 3273
rect 316 3263 323 3473
rect 336 3287 343 4033
rect 396 4027 403 4033
rect 393 4013 407 4027
rect 416 3983 423 4436
rect 476 4227 483 4453
rect 536 4267 543 4476
rect 553 4473 567 4487
rect 596 4463 603 4513
rect 736 4507 743 4533
rect 633 4503 647 4507
rect 633 4496 663 4503
rect 633 4493 647 4496
rect 656 4487 663 4496
rect 613 4463 627 4467
rect 596 4456 627 4463
rect 696 4487 703 4493
rect 693 4473 707 4487
rect 613 4453 627 4456
rect 756 4447 763 4453
rect 837 4436 845 4516
rect 896 4487 903 4493
rect 893 4473 907 4487
rect 933 4483 947 4487
rect 933 4476 963 4483
rect 933 4473 947 4476
rect 956 4427 963 4476
rect 837 4398 845 4422
rect 976 4404 984 4516
rect 996 4467 1003 4513
rect 1076 4487 1083 4513
rect 1033 4483 1047 4487
rect 1016 4476 1047 4483
rect 1016 4447 1023 4476
rect 1033 4473 1047 4476
rect 1073 4473 1087 4487
rect 1016 4327 1023 4433
rect 1116 4427 1123 4513
rect 1136 4483 1143 4533
rect 1153 4483 1167 4487
rect 1136 4476 1167 4483
rect 1153 4473 1167 4476
rect 1177 4436 1185 4516
rect 1236 4487 1243 4493
rect 1276 4487 1283 4513
rect 1233 4473 1247 4487
rect 1273 4473 1287 4487
rect 1177 4398 1185 4422
rect 1316 4404 1324 4516
rect 453 4173 467 4187
rect 456 4167 463 4173
rect 476 4047 483 4193
rect 496 4023 503 4253
rect 536 4207 543 4233
rect 613 4213 627 4227
rect 653 4223 667 4227
rect 513 4173 527 4187
rect 533 4193 547 4207
rect 593 4193 607 4207
rect 516 4047 523 4173
rect 596 4167 603 4193
rect 616 4167 623 4213
rect 653 4216 683 4223
rect 653 4213 667 4216
rect 396 3976 423 3983
rect 476 4016 503 4023
rect 356 3664 364 3776
rect 396 3687 403 3976
rect 433 3973 447 3987
rect 416 3727 423 3813
rect 436 3787 443 3973
rect 476 3807 483 4016
rect 527 4016 563 4023
rect 556 4007 563 4016
rect 553 3993 567 4007
rect 576 3987 583 4073
rect 596 4007 603 4033
rect 616 4007 623 4153
rect 613 3993 627 4007
rect 593 3953 607 3967
rect 636 3963 643 4193
rect 676 4187 683 4216
rect 696 4207 703 4233
rect 693 4193 707 4207
rect 753 4183 767 4187
rect 776 4183 783 4213
rect 753 4176 783 4183
rect 753 4173 767 4176
rect 816 4167 823 4193
rect 853 4173 867 4187
rect 656 4027 663 4133
rect 756 4027 763 4073
rect 856 4047 863 4173
rect 753 4013 767 4027
rect 656 4007 663 4013
rect 653 3993 667 4007
rect 716 3987 723 4013
rect 627 3956 643 3963
rect 596 3947 603 3953
rect 476 3727 483 3753
rect 433 3723 447 3727
rect 427 3716 447 3723
rect 433 3713 447 3716
rect 453 3693 467 3707
rect 473 3713 487 3727
rect 513 3703 527 3707
rect 536 3703 543 3753
rect 556 3747 563 3773
rect 513 3696 543 3703
rect 513 3693 527 3696
rect 573 3693 587 3707
rect 393 3493 407 3507
rect 456 3523 463 3693
rect 436 3516 463 3523
rect 396 3483 403 3493
rect 396 3476 413 3483
rect 416 3267 423 3453
rect 436 3287 443 3516
rect 493 3483 507 3487
rect 516 3483 523 3533
rect 576 3527 583 3693
rect 596 3527 603 3793
rect 616 3667 623 3953
rect 676 3767 683 3973
rect 736 3747 743 3993
rect 776 3747 783 3933
rect 733 3743 747 3747
rect 716 3736 747 3743
rect 633 3723 647 3727
rect 633 3716 663 3723
rect 633 3713 647 3716
rect 656 3583 663 3716
rect 693 3683 707 3687
rect 716 3683 723 3736
rect 733 3733 747 3736
rect 753 3713 767 3727
rect 693 3676 723 3683
rect 693 3673 707 3676
rect 656 3576 683 3583
rect 656 3547 663 3553
rect 653 3533 667 3547
rect 493 3476 523 3483
rect 493 3473 507 3476
rect 316 3256 343 3263
rect 296 3247 303 3253
rect 336 3247 343 3256
rect 413 3263 427 3267
rect 273 3213 287 3227
rect 293 3233 307 3247
rect 313 3213 327 3227
rect 333 3233 347 3247
rect 413 3256 443 3263
rect 413 3253 427 3256
rect 353 3213 367 3227
rect 436 3223 443 3256
rect 476 3247 483 3253
rect 453 3223 467 3227
rect 436 3216 467 3223
rect 473 3233 487 3247
rect 276 3127 283 3213
rect 216 2856 243 2863
rect 195 2798 203 2822
rect 195 2704 203 2784
rect 216 2747 223 2793
rect 213 2733 227 2747
rect 236 2607 243 2856
rect 256 2743 263 3113
rect 316 3067 323 3213
rect 356 3167 363 3213
rect 336 3067 343 3133
rect 276 3027 283 3053
rect 333 3043 347 3047
rect 273 3013 287 3027
rect 333 3036 363 3043
rect 333 3033 347 3036
rect 316 2787 323 2993
rect 356 2987 363 3036
rect 396 3027 403 3133
rect 373 2993 387 3007
rect 393 3013 407 3027
rect 376 2867 383 2993
rect 436 2867 443 3216
rect 453 3213 467 3216
rect 536 3223 543 3273
rect 576 3247 583 3273
rect 596 3267 603 3433
rect 616 3287 623 3513
rect 676 3527 683 3576
rect 716 3527 723 3653
rect 756 3583 763 3713
rect 796 3607 803 4033
rect 896 4007 903 4313
rect 1196 4227 1203 4233
rect 1016 4207 1023 4213
rect 933 4173 947 4187
rect 1013 4193 1027 4207
rect 973 4173 987 4187
rect 916 4107 923 4173
rect 936 4167 943 4173
rect 976 4167 983 4173
rect 853 4003 867 4007
rect 833 3973 847 3987
rect 853 3996 873 4003
rect 853 3993 867 3996
rect 836 3967 843 3973
rect 896 3963 903 3993
rect 976 3987 983 4033
rect 996 4027 1003 4193
rect 1053 4173 1067 4187
rect 1056 4167 1063 4173
rect 1116 4183 1123 4213
rect 1107 4176 1123 4183
rect 1133 4173 1147 4187
rect 1173 4183 1187 4187
rect 1196 4183 1203 4193
rect 1033 4163 1047 4167
rect 1016 4156 1047 4163
rect 1016 4107 1023 4156
rect 1033 4153 1047 4156
rect 1073 4153 1087 4167
rect 1036 4063 1043 4093
rect 1016 4056 1043 4063
rect 1016 4047 1023 4056
rect 1036 4027 1043 4033
rect 1076 4023 1083 4153
rect 1136 4107 1143 4173
rect 1173 4176 1203 4183
rect 1173 4173 1187 4176
rect 1213 4173 1227 4187
rect 1153 4163 1167 4167
rect 1153 4156 1173 4163
rect 1153 4153 1167 4156
rect 1216 4143 1223 4173
rect 1256 4167 1263 4173
rect 1336 4167 1343 4493
rect 1416 4487 1423 4513
rect 1393 4453 1407 4467
rect 1413 4473 1427 4487
rect 1433 4463 1447 4467
rect 1433 4456 1463 4463
rect 1433 4453 1447 4456
rect 1396 4447 1403 4453
rect 1456 4427 1463 4456
rect 1397 4238 1405 4262
rect 1196 4136 1223 4143
rect 1096 4027 1103 4053
rect 1196 4047 1203 4136
rect 1216 4027 1223 4113
rect 1276 4027 1283 4073
rect 913 3963 927 3967
rect 896 3956 927 3963
rect 976 3967 983 3973
rect 913 3953 927 3956
rect 953 3953 967 3967
rect 916 3947 923 3953
rect 816 3707 823 3733
rect 836 3664 844 3776
rect 873 3703 887 3707
rect 896 3703 903 3933
rect 916 3827 923 3933
rect 956 3727 963 3953
rect 975 3758 983 3782
rect 873 3696 903 3703
rect 873 3693 887 3696
rect 913 3693 927 3707
rect 916 3687 923 3693
rect 756 3576 783 3583
rect 756 3527 763 3553
rect 776 3527 783 3576
rect 816 3527 823 3533
rect 856 3527 863 3553
rect 713 3513 727 3527
rect 693 3503 707 3507
rect 676 3496 707 3503
rect 656 3263 663 3493
rect 676 3487 683 3496
rect 693 3493 707 3496
rect 753 3513 767 3527
rect 813 3513 827 3527
rect 793 3503 807 3507
rect 787 3496 807 3503
rect 793 3493 807 3496
rect 853 3513 867 3527
rect 893 3493 907 3507
rect 676 3467 683 3473
rect 716 3267 723 3473
rect 673 3263 687 3267
rect 656 3256 687 3263
rect 673 3253 687 3256
rect 553 3223 567 3227
rect 536 3216 567 3223
rect 573 3233 587 3247
rect 613 3233 627 3247
rect 553 3213 567 3216
rect 593 3213 607 3227
rect 453 3033 467 3047
rect 456 3007 463 3033
rect 477 2996 485 3076
rect 536 3047 543 3093
rect 596 3083 603 3213
rect 616 3147 623 3233
rect 576 3076 603 3083
rect 576 3047 583 3076
rect 573 3033 587 3047
rect 336 2787 343 2793
rect 296 2767 303 2773
rect 336 2767 343 2773
rect 273 2743 287 2747
rect 256 2736 287 2743
rect 293 2753 307 2767
rect 195 2516 203 2596
rect 213 2553 227 2567
rect 216 2527 223 2553
rect 195 2478 203 2502
rect 195 2318 203 2342
rect 195 2224 203 2304
rect 216 2267 223 2293
rect 213 2253 227 2267
rect 176 2176 203 2183
rect 156 2063 163 2153
rect 173 2063 187 2067
rect 156 2056 187 2063
rect 173 2053 187 2056
rect 93 1776 123 1783
rect 93 1773 107 1776
rect 33 1583 47 1587
rect 16 1576 47 1583
rect 33 1573 47 1576
rect 36 1527 43 1573
rect 57 1358 65 1382
rect 33 1303 47 1307
rect 16 1296 47 1303
rect 16 1147 23 1296
rect 33 1293 47 1296
rect 57 1264 65 1344
rect 113 1293 127 1307
rect 116 1287 123 1293
rect 136 1227 143 1753
rect 156 1567 163 2033
rect 176 1787 183 2053
rect 196 2027 203 2176
rect 236 2123 243 2533
rect 256 2327 263 2736
rect 273 2733 287 2736
rect 313 2733 327 2747
rect 333 2753 347 2767
rect 436 2747 443 2853
rect 353 2733 367 2747
rect 276 2547 283 2573
rect 296 2567 303 2713
rect 316 2587 323 2733
rect 356 2727 363 2733
rect 356 2567 363 2573
rect 376 2567 383 2613
rect 396 2567 403 2733
rect 456 2627 463 2993
rect 477 2958 485 2982
rect 616 2964 624 3076
rect 636 2827 643 3253
rect 713 3253 727 3267
rect 756 3247 763 3433
rect 753 3233 767 3247
rect 776 3207 783 3493
rect 816 3247 823 3473
rect 896 3467 903 3493
rect 916 3487 923 3673
rect 975 3664 983 3744
rect 996 3707 1003 3993
rect 1056 4016 1083 4023
rect 1056 3747 1063 4016
rect 1093 4013 1107 4027
rect 1133 4023 1147 4027
rect 1116 4016 1147 4023
rect 1116 4007 1123 4016
rect 1133 4013 1147 4016
rect 1213 4013 1227 4027
rect 1193 4003 1207 4007
rect 1153 3983 1167 3987
rect 1176 3996 1207 4003
rect 1176 3983 1183 3996
rect 1153 3976 1183 3983
rect 1193 3993 1207 3996
rect 1153 3973 1167 3976
rect 993 3693 1007 3707
rect 1053 3703 1067 3707
rect 1076 3703 1083 3933
rect 1053 3696 1083 3703
rect 1136 3707 1143 3973
rect 1157 3758 1165 3782
rect 1176 3747 1183 3976
rect 1053 3693 1067 3696
rect 1093 3693 1107 3707
rect 1133 3693 1147 3707
rect 1096 3683 1103 3693
rect 1076 3676 1103 3683
rect 936 3507 943 3533
rect 956 3527 963 3573
rect 976 3547 983 3553
rect 973 3533 987 3547
rect 953 3513 967 3527
rect 996 3527 1003 3533
rect 1057 3476 1065 3556
rect 1076 3467 1083 3676
rect 1157 3664 1165 3744
rect 1057 3438 1065 3462
rect 813 3243 827 3247
rect 796 3236 827 3243
rect 493 2733 507 2747
rect 533 2743 547 2747
rect 556 2743 563 2773
rect 533 2736 563 2743
rect 533 2733 547 2736
rect 573 2733 587 2747
rect 496 2707 503 2733
rect 293 2553 307 2567
rect 273 2533 287 2547
rect 353 2553 367 2567
rect 393 2553 407 2567
rect 253 2253 267 2267
rect 313 2273 327 2287
rect 216 2116 243 2123
rect 216 2047 223 2116
rect 256 2107 263 2253
rect 316 2227 323 2273
rect 336 2207 343 2493
rect 376 2287 383 2513
rect 416 2347 423 2613
rect 496 2367 503 2633
rect 536 2627 543 2733
rect 576 2727 583 2733
rect 576 2687 583 2713
rect 596 2647 603 2813
rect 636 2787 643 2793
rect 633 2773 647 2787
rect 613 2733 627 2747
rect 516 2527 523 2613
rect 596 2567 603 2613
rect 616 2607 623 2733
rect 676 2667 683 2733
rect 696 2727 703 3153
rect 716 2964 724 3076
rect 736 2923 743 3193
rect 796 3187 803 3236
rect 813 3233 827 3236
rect 756 3047 763 3073
rect 796 3047 803 3173
rect 753 3033 767 3047
rect 855 2996 863 3076
rect 913 3063 927 3067
rect 873 3043 887 3047
rect 896 3056 927 3063
rect 896 3043 903 3056
rect 873 3036 903 3043
rect 913 3053 927 3056
rect 1013 3063 1027 3067
rect 1007 3056 1027 3063
rect 1013 3053 1027 3056
rect 873 3033 887 3036
rect 933 3023 947 3027
rect 956 3023 963 3033
rect 933 3016 963 3023
rect 933 3013 947 3016
rect 956 3007 963 3016
rect 976 2987 983 3053
rect 1036 3047 1043 3053
rect 1033 3033 1047 3047
rect 1056 3003 1063 3233
rect 1096 3107 1103 3593
rect 1113 3523 1127 3527
rect 1136 3523 1143 3633
rect 1156 3527 1163 3553
rect 1113 3516 1143 3523
rect 1113 3513 1127 3516
rect 1136 3483 1143 3516
rect 1153 3513 1167 3527
rect 1136 3476 1163 3483
rect 1156 3247 1163 3476
rect 1153 3233 1167 3247
rect 1176 3167 1183 3713
rect 1213 3693 1227 3707
rect 1216 3687 1223 3693
rect 1296 3664 1304 3776
rect 1336 3647 1343 4153
rect 1356 4007 1363 4213
rect 1397 4144 1405 4224
rect 1453 4173 1467 4187
rect 1456 4167 1463 4173
rect 1376 4027 1383 4053
rect 1476 4047 1483 4473
rect 1516 4404 1524 4516
rect 1596 4487 1603 4493
rect 1553 4483 1567 4487
rect 1536 4476 1567 4483
rect 1536 4303 1543 4476
rect 1553 4473 1567 4476
rect 1593 4473 1607 4487
rect 1655 4436 1663 4516
rect 1516 4296 1543 4303
rect 1456 4027 1463 4033
rect 1373 4013 1387 4027
rect 1353 3993 1367 4007
rect 1453 4013 1467 4027
rect 1393 4003 1407 4007
rect 1393 3996 1423 4003
rect 1393 3993 1407 3996
rect 1416 3983 1423 3996
rect 1476 4007 1483 4013
rect 1516 4007 1523 4296
rect 1536 4144 1544 4256
rect 1616 4207 1623 4433
rect 1753 4433 1767 4447
rect 1655 4398 1663 4422
rect 1576 4183 1583 4193
rect 1593 4183 1607 4187
rect 1576 4176 1607 4183
rect 1613 4193 1627 4207
rect 1653 4193 1667 4207
rect 1593 4173 1607 4176
rect 1616 4007 1623 4133
rect 1656 4107 1663 4193
rect 1676 4027 1683 4393
rect 1693 4173 1707 4187
rect 1696 4047 1703 4173
rect 1733 4173 1747 4187
rect 1736 4167 1743 4173
rect 1713 4153 1727 4167
rect 1716 4127 1723 4153
rect 1416 3976 1433 3983
rect 1473 3993 1487 4007
rect 1513 3993 1527 4007
rect 1533 3983 1547 3987
rect 1533 3976 1563 3983
rect 1533 3973 1547 3976
rect 1556 3767 1563 3976
rect 1593 3973 1607 3987
rect 1613 3993 1627 4007
rect 1596 3967 1603 3973
rect 1676 3967 1683 4013
rect 1693 3963 1707 3967
rect 1687 3956 1707 3963
rect 1693 3953 1707 3956
rect 1376 3727 1383 3733
rect 1353 3693 1367 3707
rect 1373 3713 1387 3727
rect 1436 3736 1453 3743
rect 1356 3687 1363 3693
rect 1436 3687 1443 3736
rect 1493 3743 1507 3747
rect 1493 3736 1523 3743
rect 1493 3733 1507 3736
rect 1516 3707 1523 3736
rect 1573 3743 1587 3747
rect 1573 3736 1603 3743
rect 1573 3733 1587 3736
rect 1196 3444 1204 3556
rect 1313 3523 1327 3527
rect 1296 3516 1327 3523
rect 1396 3527 1403 3673
rect 1436 3527 1443 3553
rect 1353 3523 1367 3527
rect 1296 3507 1303 3516
rect 1313 3513 1327 3516
rect 1273 3503 1287 3507
rect 1273 3496 1293 3503
rect 1273 3493 1287 3496
rect 1353 3516 1383 3523
rect 1353 3513 1367 3516
rect 1196 3236 1213 3243
rect 1176 3047 1183 3073
rect 1196 3067 1203 3236
rect 1256 3067 1263 3333
rect 1297 3278 1305 3302
rect 1297 3184 1305 3264
rect 1253 3053 1267 3067
rect 1036 2996 1063 3003
rect 855 2958 863 2982
rect 716 2916 743 2923
rect 716 2703 723 2916
rect 956 2827 963 2973
rect 956 2787 963 2813
rect 913 2783 927 2787
rect 896 2776 927 2783
rect 793 2743 807 2747
rect 833 2743 847 2747
rect 793 2736 847 2743
rect 793 2733 807 2736
rect 696 2696 723 2703
rect 616 2567 623 2573
rect 613 2563 627 2567
rect 613 2556 643 2563
rect 613 2553 627 2556
rect 636 2527 643 2556
rect 676 2547 683 2613
rect 416 2287 423 2293
rect 373 2273 387 2287
rect 393 2253 407 2267
rect 413 2273 427 2287
rect 433 2263 447 2267
rect 456 2263 463 2313
rect 433 2256 463 2263
rect 433 2253 447 2256
rect 273 2033 287 2047
rect 195 1838 203 1862
rect 176 1647 183 1773
rect 195 1744 203 1824
rect 216 1787 223 1993
rect 213 1773 227 1787
rect 236 1767 243 2013
rect 276 2007 283 2033
rect 296 1827 303 2113
rect 316 2087 323 2133
rect 356 2103 363 2253
rect 396 2147 403 2253
rect 456 2103 463 2256
rect 473 2253 487 2267
rect 476 2127 483 2253
rect 356 2096 403 2103
rect 456 2096 483 2103
rect 396 2087 403 2096
rect 476 2087 483 2096
rect 353 2053 367 2067
rect 393 2073 407 2087
rect 413 2053 427 2067
rect 473 2073 487 2087
rect 496 2067 503 2333
rect 513 2253 527 2267
rect 516 2207 523 2253
rect 316 1847 323 1993
rect 253 1773 267 1787
rect 313 1793 327 1807
rect 316 1787 323 1793
rect 256 1627 263 1773
rect 336 1627 343 2033
rect 356 2027 363 2053
rect 376 1867 383 2033
rect 416 2007 423 2053
rect 356 1803 363 1833
rect 536 1827 543 2353
rect 596 2307 603 2513
rect 696 2507 703 2696
rect 716 2547 723 2653
rect 736 2567 743 2633
rect 816 2587 823 2736
rect 833 2733 847 2736
rect 876 2707 883 2733
rect 896 2727 903 2776
rect 913 2773 927 2776
rect 933 2753 947 2767
rect 953 2773 967 2787
rect 996 2767 1003 2773
rect 993 2753 1007 2767
rect 936 2667 943 2753
rect 1016 2727 1023 2813
rect 813 2573 827 2587
rect 733 2553 747 2567
rect 773 2563 787 2567
rect 713 2533 727 2547
rect 773 2556 793 2563
rect 773 2553 787 2556
rect 833 2563 847 2567
rect 856 2563 863 2573
rect 833 2556 863 2563
rect 833 2553 847 2556
rect 856 2547 863 2556
rect 573 2273 587 2287
rect 593 2293 607 2307
rect 576 2227 583 2273
rect 616 2247 623 2333
rect 716 2287 723 2353
rect 653 2283 667 2287
rect 636 2276 667 2283
rect 636 2187 643 2276
rect 653 2273 667 2276
rect 693 2253 707 2267
rect 673 2243 687 2247
rect 696 2243 703 2253
rect 673 2236 703 2243
rect 733 2253 747 2267
rect 673 2233 687 2236
rect 713 2233 727 2247
rect 636 2147 643 2153
rect 556 2004 564 2116
rect 596 2087 603 2113
rect 636 2087 643 2133
rect 676 2087 683 2233
rect 716 2167 723 2233
rect 736 2207 743 2253
rect 593 2073 607 2087
rect 633 2073 647 2087
rect 695 2036 703 2116
rect 736 2027 743 2073
rect 695 1998 703 2022
rect 373 1803 387 1807
rect 356 1796 387 1803
rect 373 1793 387 1796
rect 393 1773 407 1787
rect 433 1773 447 1787
rect 396 1767 403 1773
rect 436 1767 443 1773
rect 456 1743 463 1793
rect 556 1803 563 1833
rect 616 1807 623 1813
rect 573 1803 587 1807
rect 556 1796 587 1803
rect 573 1793 587 1796
rect 533 1773 547 1787
rect 613 1793 627 1807
rect 536 1763 543 1773
rect 636 1767 643 1773
rect 436 1736 463 1743
rect 516 1756 543 1763
rect 253 1613 267 1627
rect 233 1603 247 1607
rect 216 1596 247 1603
rect 316 1607 323 1613
rect 356 1607 363 1653
rect 153 1303 167 1307
rect 153 1296 183 1303
rect 153 1293 167 1296
rect 13 1133 27 1147
rect 36 1087 43 1093
rect 56 784 64 896
rect 116 823 123 893
rect 133 823 147 827
rect 116 816 147 823
rect 133 813 147 816
rect 56 564 64 676
rect 136 647 143 813
rect 93 643 107 647
rect 93 636 123 643
rect 93 633 107 636
rect 56 304 64 416
rect 76 343 83 413
rect 116 347 123 636
rect 156 627 163 1253
rect 176 1207 183 1296
rect 196 1264 204 1376
rect 216 1267 223 1596
rect 233 1593 247 1596
rect 313 1593 327 1607
rect 176 1127 183 1173
rect 196 1127 203 1213
rect 236 1187 243 1553
rect 296 1427 303 1593
rect 353 1593 367 1607
rect 256 1227 263 1413
rect 296 1264 304 1376
rect 373 1303 387 1307
rect 396 1303 403 1573
rect 416 1524 424 1636
rect 436 1563 443 1736
rect 493 1603 507 1607
rect 476 1596 507 1603
rect 476 1587 483 1596
rect 493 1593 507 1596
rect 516 1587 523 1756
rect 653 1763 667 1767
rect 696 1763 703 1833
rect 736 1807 743 1953
rect 713 1763 727 1767
rect 653 1756 683 1763
rect 696 1756 727 1763
rect 653 1753 667 1756
rect 436 1556 463 1563
rect 435 1358 443 1382
rect 456 1347 463 1556
rect 536 1367 543 1613
rect 555 1556 563 1636
rect 573 1603 587 1607
rect 596 1603 603 1613
rect 573 1596 603 1603
rect 573 1593 587 1596
rect 555 1518 563 1542
rect 373 1296 403 1303
rect 373 1293 387 1296
rect 376 1287 383 1293
rect 256 1143 263 1213
rect 236 1136 263 1143
rect 236 1127 243 1136
rect 296 1127 303 1193
rect 193 1113 207 1127
rect 213 1093 227 1107
rect 233 1113 247 1127
rect 293 1113 307 1127
rect 313 1093 327 1107
rect 176 787 183 1033
rect 195 878 203 902
rect 216 867 223 1093
rect 316 1067 323 1093
rect 195 784 203 864
rect 216 827 223 853
rect 213 813 227 827
rect 176 423 183 633
rect 195 596 203 676
rect 253 663 267 667
rect 213 633 227 647
rect 236 656 267 663
rect 216 627 223 633
rect 236 607 243 656
rect 253 653 267 656
rect 273 613 287 627
rect 195 558 203 582
rect 156 416 183 423
rect 93 343 107 347
rect 76 336 107 343
rect 93 333 107 336
rect 133 343 147 347
rect 156 343 163 416
rect 195 398 203 422
rect 133 336 163 343
rect 133 333 147 336
rect 56 84 64 196
rect 136 167 143 333
rect 176 167 183 393
rect 256 387 263 613
rect 276 407 283 613
rect 296 387 303 793
rect 316 647 323 1013
rect 356 907 363 1273
rect 435 1264 443 1344
rect 456 1307 463 1333
rect 453 1293 467 1307
rect 376 1087 383 1213
rect 396 1127 403 1153
rect 393 1113 407 1127
rect 476 1107 483 1353
rect 536 1347 543 1353
rect 533 1333 547 1347
rect 556 1267 563 1473
rect 576 1303 583 1573
rect 656 1524 664 1636
rect 676 1607 683 1756
rect 713 1753 727 1756
rect 756 1667 763 2513
rect 776 2263 783 2493
rect 876 2303 883 2633
rect 916 2484 924 2596
rect 953 2563 967 2567
rect 936 2556 967 2563
rect 936 2527 943 2556
rect 953 2553 967 2556
rect 976 2367 983 2673
rect 993 2563 1007 2567
rect 993 2556 1023 2563
rect 993 2553 1007 2556
rect 856 2296 883 2303
rect 816 2287 823 2293
rect 856 2287 863 2296
rect 793 2263 807 2267
rect 776 2256 807 2263
rect 813 2273 827 2287
rect 793 2253 807 2256
rect 873 2253 887 2267
rect 833 2233 847 2247
rect 836 2227 843 2233
rect 796 2067 803 2073
rect 793 2053 807 2067
rect 836 2047 843 2213
rect 856 2107 863 2233
rect 876 2167 883 2253
rect 913 2253 927 2267
rect 916 2247 923 2253
rect 936 2247 943 2293
rect 953 2253 967 2267
rect 1016 2267 1023 2556
rect 1036 2307 1043 2996
rect 1153 3013 1167 3027
rect 1173 3033 1187 3047
rect 1193 3023 1207 3027
rect 1193 3016 1223 3023
rect 1193 3013 1207 3016
rect 1113 2993 1127 3007
rect 1156 3003 1163 3013
rect 1156 2996 1183 3003
rect 1116 2987 1123 2993
rect 1136 2787 1143 2993
rect 1176 2787 1183 2996
rect 1216 2947 1223 3016
rect 1233 3013 1247 3027
rect 1073 2753 1087 2767
rect 1076 2627 1083 2753
rect 1113 2733 1127 2747
rect 1055 2516 1063 2596
rect 1116 2587 1123 2733
rect 1153 2733 1167 2747
rect 1133 2713 1147 2727
rect 1136 2707 1143 2713
rect 1156 2627 1163 2733
rect 1176 2647 1183 2773
rect 1213 2733 1227 2747
rect 1216 2647 1223 2733
rect 1236 2687 1243 3013
rect 1316 3003 1323 3453
rect 1376 3447 1383 3516
rect 1433 3513 1447 3527
rect 1476 3483 1483 3513
rect 1493 3483 1507 3487
rect 1476 3476 1507 3483
rect 1353 3213 1367 3227
rect 1393 3213 1407 3227
rect 1356 3187 1363 3213
rect 1396 3187 1403 3213
rect 1436 3184 1444 3296
rect 1476 3223 1483 3476
rect 1493 3473 1507 3476
rect 1533 3473 1547 3487
rect 1536 3427 1543 3473
rect 1493 3223 1507 3227
rect 1476 3216 1507 3223
rect 1553 3233 1567 3247
rect 1493 3213 1507 3216
rect 1533 3213 1547 3227
rect 1536 3187 1543 3213
rect 1556 3187 1563 3233
rect 1356 3087 1363 3173
rect 1336 3027 1343 3053
rect 1296 2996 1323 3003
rect 1296 2747 1303 2996
rect 1376 2964 1384 3076
rect 1113 2583 1127 2587
rect 1073 2563 1087 2567
rect 1096 2576 1127 2583
rect 1096 2563 1103 2576
rect 1073 2556 1103 2563
rect 1113 2573 1127 2576
rect 1176 2567 1183 2633
rect 1073 2553 1087 2556
rect 1173 2553 1187 2567
rect 1156 2527 1163 2553
rect 1055 2478 1063 2502
rect 893 2233 907 2247
rect 896 2227 903 2233
rect 813 2033 827 2047
rect 816 2007 823 2033
rect 876 2027 883 2093
rect 896 2087 903 2213
rect 956 2187 963 2253
rect 1033 2233 1047 2247
rect 1036 2207 1043 2233
rect 893 2073 907 2087
rect 916 2007 923 2053
rect 973 2033 987 2047
rect 976 2027 983 2033
rect 996 1967 1003 2093
rect 1016 2087 1023 2153
rect 1076 2107 1083 2353
rect 1137 2318 1145 2342
rect 1113 2263 1127 2267
rect 1096 2256 1127 2263
rect 1096 2207 1103 2256
rect 1113 2253 1127 2256
rect 1137 2224 1145 2304
rect 1156 2227 1163 2433
rect 1233 2253 1247 2267
rect 1056 2096 1073 2103
rect 1056 2087 1063 2096
rect 1136 2087 1143 2113
rect 1156 2087 1163 2173
rect 1196 2147 1203 2253
rect 1236 2247 1243 2253
rect 1053 2073 1067 2087
rect 1093 2083 1107 2087
rect 1076 2076 1107 2083
rect 1076 2047 1083 2076
rect 1093 2073 1107 2076
rect 1133 2073 1147 2087
rect 1193 2043 1207 2047
rect 1187 2036 1207 2043
rect 1193 2033 1207 2036
rect 816 1847 823 1953
rect 696 1607 703 1613
rect 736 1607 743 1633
rect 693 1593 707 1607
rect 733 1593 747 1607
rect 776 1487 783 1813
rect 816 1807 823 1833
rect 873 1813 887 1827
rect 853 1793 867 1807
rect 836 1767 843 1773
rect 813 1753 827 1767
rect 816 1727 823 1753
rect 795 1556 803 1636
rect 856 1627 863 1793
rect 876 1787 883 1813
rect 996 1744 1004 1856
rect 813 1593 827 1607
rect 795 1518 803 1542
rect 816 1427 823 1593
rect 897 1556 905 1636
rect 897 1518 905 1542
rect 776 1327 783 1353
rect 896 1347 903 1473
rect 576 1296 603 1303
rect 453 1093 467 1107
rect 456 1087 463 1093
rect 516 1087 523 1193
rect 556 1147 563 1193
rect 553 1133 567 1147
rect 536 1127 543 1133
rect 533 1113 547 1127
rect 576 1127 583 1213
rect 596 1147 603 1296
rect 653 1303 667 1307
rect 713 1303 727 1307
rect 653 1296 727 1303
rect 653 1293 667 1296
rect 713 1293 727 1296
rect 776 1283 783 1313
rect 793 1303 807 1307
rect 816 1303 823 1333
rect 793 1296 823 1303
rect 873 1313 887 1327
rect 893 1333 907 1347
rect 793 1293 807 1296
rect 756 1276 783 1283
rect 593 1133 607 1147
rect 573 1113 587 1127
rect 376 1027 383 1073
rect 636 1067 643 1153
rect 676 1127 683 1273
rect 673 1113 687 1127
rect 336 807 343 853
rect 413 813 427 827
rect 416 807 423 813
rect 356 647 363 773
rect 456 743 463 833
rect 476 784 484 896
rect 536 823 543 893
rect 615 878 623 902
rect 553 823 567 827
rect 536 816 567 823
rect 553 813 567 816
rect 596 807 603 873
rect 456 736 483 743
rect 333 613 347 627
rect 353 633 367 647
rect 336 607 343 613
rect 396 603 403 633
rect 413 603 427 607
rect 396 596 427 603
rect 413 593 427 596
rect 195 304 203 384
rect 253 373 267 387
rect 293 383 307 387
rect 293 376 323 383
rect 293 373 307 376
rect 213 343 227 347
rect 213 336 243 343
rect 213 333 227 336
rect 236 287 243 336
rect 93 163 107 167
rect 93 156 123 163
rect 93 153 107 156
rect 116 147 123 156
rect 133 153 147 167
rect 195 116 203 196
rect 213 163 227 167
rect 236 163 243 213
rect 316 187 323 376
rect 336 227 343 593
rect 476 387 483 736
rect 496 647 503 733
rect 536 647 543 793
rect 615 784 623 864
rect 636 827 643 853
rect 633 813 647 827
rect 656 767 663 1113
rect 716 1067 723 1253
rect 733 1123 747 1127
rect 756 1123 763 1276
rect 836 1203 843 1293
rect 876 1203 883 1313
rect 916 1307 923 1413
rect 936 1287 943 1653
rect 956 1607 963 1633
rect 953 1593 967 1607
rect 993 1603 1007 1607
rect 1016 1603 1023 2033
rect 1033 1773 1047 1787
rect 1036 1767 1043 1773
rect 993 1596 1023 1603
rect 993 1593 1007 1596
rect 1036 1524 1044 1636
rect 1056 1427 1063 2013
rect 1135 1838 1143 1862
rect 1073 1773 1087 1787
rect 1076 1647 1083 1773
rect 1096 1387 1103 1813
rect 1135 1744 1143 1824
rect 1156 1787 1163 1813
rect 1153 1773 1167 1787
rect 1153 1553 1167 1567
rect 1156 1547 1163 1553
rect 1156 1487 1163 1533
rect 996 1327 1003 1353
rect 1096 1347 1103 1353
rect 973 1293 987 1307
rect 993 1313 1007 1327
rect 1013 1293 1027 1307
rect 1096 1303 1103 1333
rect 1113 1303 1127 1307
rect 816 1196 843 1203
rect 856 1196 883 1203
rect 816 1127 823 1196
rect 856 1143 863 1196
rect 876 1147 883 1173
rect 836 1136 863 1143
rect 733 1116 763 1123
rect 733 1113 747 1116
rect 756 1067 763 1116
rect 773 1123 787 1127
rect 773 1116 803 1123
rect 773 1113 787 1116
rect 676 867 683 1053
rect 716 867 723 873
rect 713 853 727 867
rect 613 663 627 667
rect 613 656 643 663
rect 613 653 627 656
rect 493 633 507 647
rect 533 633 547 647
rect 636 643 643 656
rect 653 643 667 647
rect 636 636 667 643
rect 653 633 667 636
rect 596 607 603 613
rect 677 596 685 676
rect 736 647 743 893
rect 796 867 803 1116
rect 813 1113 827 1127
rect 836 863 843 1136
rect 873 1133 887 1147
rect 896 1127 903 1133
rect 916 1087 923 1273
rect 976 1207 983 1293
rect 1016 1247 1023 1293
rect 1096 1296 1127 1303
rect 1113 1293 1127 1296
rect 1073 1273 1087 1287
rect 956 1147 963 1153
rect 953 1133 967 1147
rect 933 1093 947 1107
rect 936 1087 943 1093
rect 976 907 983 1173
rect 1036 1127 1043 1233
rect 1076 1187 1083 1273
rect 1056 1147 1063 1153
rect 1053 1133 1067 1147
rect 1033 1113 1047 1127
rect 1076 1127 1083 1173
rect 1073 1113 1087 1127
rect 1096 867 1103 1153
rect 1116 1147 1123 1153
rect 1113 1133 1127 1147
rect 1136 1143 1143 1373
rect 1176 1367 1183 2033
rect 1256 2027 1263 2733
rect 1316 2704 1324 2816
rect 1353 2743 1367 2747
rect 1376 2743 1383 2813
rect 1353 2736 1383 2743
rect 1353 2733 1367 2736
rect 1393 2733 1407 2747
rect 1276 2587 1283 2613
rect 1273 2573 1287 2587
rect 1316 2523 1323 2633
rect 1396 2627 1403 2733
rect 1436 2647 1443 3093
rect 1456 3047 1463 3073
rect 1453 3033 1467 3047
rect 1455 2798 1463 2822
rect 1455 2704 1463 2784
rect 1476 2747 1483 3093
rect 1496 2727 1503 3133
rect 1576 3107 1583 3693
rect 1596 3667 1603 3736
rect 1613 3693 1627 3707
rect 1653 3703 1667 3707
rect 1676 3703 1683 3953
rect 1737 3758 1745 3782
rect 1713 3703 1727 3707
rect 1653 3696 1683 3703
rect 1696 3696 1727 3703
rect 1653 3693 1667 3696
rect 1616 3523 1623 3693
rect 1696 3587 1703 3696
rect 1713 3693 1727 3696
rect 1737 3664 1745 3744
rect 1696 3547 1703 3573
rect 1693 3533 1707 3547
rect 1633 3523 1647 3527
rect 1616 3516 1647 3523
rect 1616 3467 1623 3516
rect 1633 3513 1647 3516
rect 1716 3523 1723 3653
rect 1756 3627 1763 4433
rect 1776 4167 1783 4473
rect 1837 4436 1845 4516
rect 1896 4487 1903 4493
rect 1893 4473 1907 4487
rect 1837 4398 1845 4422
rect 1796 4227 1803 4333
rect 1877 4238 1885 4262
rect 1796 4207 1803 4213
rect 1793 4193 1807 4207
rect 1853 4183 1867 4187
rect 1836 4176 1867 4183
rect 1836 4087 1843 4176
rect 1853 4173 1867 4176
rect 1877 4144 1885 4224
rect 1916 4183 1923 4493
rect 1976 4404 1984 4516
rect 2393 4503 2407 4507
rect 2393 4496 2423 4503
rect 2393 4493 2407 4496
rect 2116 4487 2123 4493
rect 2033 4483 2047 4487
rect 2016 4476 2047 4483
rect 2016 4347 2023 4476
rect 2033 4473 2047 4476
rect 2053 4453 2067 4467
rect 2113 4473 2127 4487
rect 2333 4483 2347 4487
rect 2056 4407 2063 4453
rect 2173 4433 2187 4447
rect 2233 4463 2247 4467
rect 2273 4463 2287 4467
rect 2233 4456 2287 4463
rect 2233 4453 2247 4456
rect 2176 4427 2183 4433
rect 2056 4387 2063 4393
rect 1933 4183 1947 4187
rect 1916 4176 1947 4183
rect 1933 4173 1947 4176
rect 1876 3987 1883 4053
rect 1896 4007 1903 4013
rect 1853 3983 1867 3987
rect 1873 3983 1887 3987
rect 1853 3976 1887 3983
rect 1853 3973 1867 3976
rect 1873 3973 1887 3976
rect 1816 3947 1823 3973
rect 1896 3967 1903 3993
rect 1893 3953 1907 3967
rect 1956 3963 1963 4193
rect 1973 4173 1987 4187
rect 1976 4147 1983 4173
rect 2016 4144 2024 4256
rect 2113 4193 2127 4207
rect 2216 4207 2223 4393
rect 2256 4387 2263 4456
rect 2273 4453 2287 4456
rect 2313 4453 2327 4467
rect 2333 4476 2363 4483
rect 2333 4473 2347 4476
rect 2356 4463 2363 4476
rect 2416 4487 2423 4496
rect 2456 4487 2463 4493
rect 2373 4463 2387 4467
rect 2356 4456 2387 4463
rect 2316 4407 2323 4453
rect 2356 4447 2363 4456
rect 2373 4453 2387 4456
rect 2453 4473 2467 4487
rect 2696 4487 2703 4553
rect 2776 4487 2783 4616
rect 2513 4453 2527 4467
rect 2573 4453 2587 4467
rect 2653 4483 2667 4487
rect 2636 4476 2667 4483
rect 2396 4427 2403 4453
rect 2116 4167 2123 4193
rect 2136 4067 2143 4173
rect 2173 4173 2187 4187
rect 2213 4193 2227 4207
rect 2236 4187 2243 4213
rect 2176 4167 2183 4173
rect 2256 4147 2263 4373
rect 2336 4207 2343 4253
rect 2396 4247 2403 4413
rect 2516 4407 2523 4453
rect 2576 4407 2583 4453
rect 2416 4267 2423 4353
rect 2416 4227 2423 4253
rect 2333 4193 2347 4207
rect 2393 4193 2407 4207
rect 2413 4213 2427 4227
rect 2396 4167 2403 4193
rect 1947 3956 1963 3963
rect 2136 3963 2143 4053
rect 2176 3987 2183 4033
rect 2336 4027 2343 4073
rect 2216 3987 2223 4013
rect 2276 3987 2283 4013
rect 2153 3963 2167 3967
rect 2136 3956 2167 3963
rect 2173 3973 2187 3987
rect 2213 3983 2227 3987
rect 2213 3976 2243 3983
rect 2213 3973 2227 3976
rect 2153 3953 2167 3956
rect 2236 3963 2243 3976
rect 2253 3963 2267 3967
rect 2236 3956 2267 3963
rect 2273 3973 2287 3987
rect 2253 3953 2267 3956
rect 1793 3693 1807 3707
rect 1833 3693 1847 3707
rect 1796 3647 1803 3693
rect 1733 3523 1747 3527
rect 1716 3516 1747 3523
rect 1733 3513 1747 3516
rect 1673 3493 1687 3507
rect 1676 3447 1683 3493
rect 1515 2996 1523 3076
rect 1596 3047 1603 3413
rect 1656 3247 1663 3273
rect 1653 3233 1667 3247
rect 1673 3213 1687 3227
rect 1636 3047 1643 3053
rect 1633 3033 1647 3047
rect 1515 2958 1523 2982
rect 1516 2787 1523 2913
rect 1656 2907 1663 3073
rect 1676 3067 1683 3213
rect 1696 3207 1703 3493
rect 1736 3267 1743 3513
rect 1757 3476 1765 3556
rect 1757 3438 1765 3462
rect 1713 3233 1727 3247
rect 1716 3227 1723 3233
rect 1733 3213 1747 3227
rect 1773 3213 1787 3227
rect 1736 3207 1743 3213
rect 1696 3027 1703 3173
rect 1776 3147 1783 3213
rect 1736 3047 1743 3053
rect 1796 3047 1803 3613
rect 1816 3527 1823 3633
rect 1836 3547 1843 3693
rect 1876 3664 1884 3776
rect 1956 3727 1963 3933
rect 1953 3713 1967 3727
rect 1996 3703 2003 3933
rect 2213 3743 2227 3747
rect 2013 3703 2027 3707
rect 1996 3696 2027 3703
rect 2073 3723 2087 3727
rect 2073 3716 2103 3723
rect 2073 3713 2087 3716
rect 2013 3693 2027 3696
rect 1973 3673 1987 3687
rect 2053 3673 2067 3687
rect 1976 3587 1983 3673
rect 2056 3607 2063 3673
rect 2096 3647 2103 3716
rect 2153 3713 2167 3727
rect 2156 3647 2163 3713
rect 2176 3687 2183 3733
rect 2193 3713 2207 3727
rect 2213 3736 2243 3743
rect 2213 3733 2227 3736
rect 2196 3607 2203 3713
rect 1813 3513 1827 3527
rect 1853 3523 1867 3527
rect 1836 3516 1867 3523
rect 1836 3507 1843 3516
rect 1853 3513 1867 3516
rect 1896 3444 1904 3556
rect 1996 3527 2003 3533
rect 1953 3523 1967 3527
rect 1936 3516 1967 3523
rect 1936 3447 1943 3516
rect 1953 3513 1967 3516
rect 1993 3513 2007 3527
rect 1976 3487 1983 3493
rect 2056 3467 2063 3573
rect 2113 3473 2127 3487
rect 2116 3467 2123 3473
rect 1916 3267 1923 3273
rect 1916 3247 1923 3253
rect 1873 3233 1887 3247
rect 1833 3193 1847 3207
rect 1836 3127 1843 3193
rect 1733 3033 1747 3047
rect 1673 2993 1687 3007
rect 1693 3013 1707 3027
rect 1753 3013 1767 3027
rect 1796 3027 1803 3033
rect 1793 3013 1807 3027
rect 1713 2993 1727 3007
rect 1676 2927 1683 2993
rect 1716 2983 1723 2993
rect 1696 2976 1723 2983
rect 1556 2787 1563 2793
rect 1533 2753 1547 2767
rect 1553 2773 1567 2787
rect 1576 2767 1583 2813
rect 1656 2767 1663 2893
rect 1613 2753 1627 2767
rect 1356 2567 1363 2613
rect 1316 2516 1333 2523
rect 1373 2513 1387 2527
rect 1457 2516 1465 2596
rect 1276 2224 1284 2336
rect 1336 2303 1343 2513
rect 1376 2427 1383 2513
rect 1457 2478 1465 2502
rect 1336 2296 1363 2303
rect 1356 2287 1363 2296
rect 1353 2273 1367 2287
rect 1393 2283 1407 2287
rect 1416 2283 1423 2353
rect 1393 2276 1423 2283
rect 1393 2273 1407 2276
rect 1373 2253 1387 2267
rect 1376 2247 1383 2253
rect 1276 2087 1283 2093
rect 1273 2073 1287 2087
rect 1376 2047 1383 2073
rect 1397 2036 1405 2116
rect 1416 2067 1423 2093
rect 1397 1998 1405 2022
rect 1213 1793 1227 1807
rect 1216 1787 1223 1793
rect 1256 1607 1263 1833
rect 1293 1793 1307 1807
rect 1253 1593 1267 1607
rect 1276 1587 1283 1793
rect 1296 1787 1303 1793
rect 1313 1773 1327 1787
rect 1393 1803 1407 1807
rect 1353 1773 1367 1787
rect 1376 1796 1407 1803
rect 1316 1767 1323 1773
rect 1356 1767 1363 1773
rect 1293 1593 1307 1607
rect 1236 1567 1243 1573
rect 1153 1293 1167 1307
rect 1156 1287 1163 1293
rect 1196 1167 1203 1393
rect 1236 1387 1243 1553
rect 1296 1547 1303 1593
rect 1317 1556 1325 1636
rect 1376 1627 1383 1796
rect 1393 1793 1407 1796
rect 1416 1623 1423 1813
rect 1396 1616 1423 1623
rect 1376 1607 1383 1613
rect 1373 1593 1387 1607
rect 1317 1518 1325 1542
rect 1236 1347 1243 1373
rect 1233 1333 1247 1347
rect 1273 1343 1287 1347
rect 1273 1336 1303 1343
rect 1273 1333 1287 1336
rect 1136 1136 1163 1143
rect 1133 1093 1147 1107
rect 836 856 863 863
rect 833 813 847 827
rect 836 807 843 813
rect 733 643 747 647
rect 733 636 763 643
rect 733 633 747 636
rect 677 558 685 582
rect 756 447 763 636
rect 816 564 824 676
rect 856 663 863 856
rect 1136 863 1143 1093
rect 1156 903 1163 1136
rect 1193 1123 1207 1127
rect 1176 1116 1207 1123
rect 1236 1127 1243 1153
rect 1276 1147 1283 1173
rect 1296 1147 1303 1336
rect 1356 1327 1363 1373
rect 1333 1293 1347 1307
rect 1353 1313 1367 1327
rect 1373 1303 1387 1307
rect 1396 1303 1403 1616
rect 1436 1407 1443 2373
rect 1456 2287 1463 2413
rect 1476 2387 1483 2633
rect 1477 2318 1485 2342
rect 1456 2267 1463 2273
rect 1453 2253 1467 2267
rect 1477 2224 1485 2304
rect 1496 2267 1503 2613
rect 1516 2567 1523 2613
rect 1513 2553 1527 2567
rect 1536 2367 1543 2753
rect 1616 2747 1623 2753
rect 1653 2753 1667 2767
rect 1673 2733 1687 2747
rect 1676 2727 1683 2733
rect 1596 2484 1604 2596
rect 1573 2253 1587 2267
rect 1576 2207 1583 2253
rect 1453 2083 1467 2087
rect 1476 2083 1483 2093
rect 1453 2076 1483 2083
rect 1453 2073 1467 2076
rect 1456 1524 1464 1636
rect 1476 1627 1483 2076
rect 1536 2004 1544 2116
rect 1596 1807 1603 2293
rect 1616 2224 1624 2336
rect 1636 2127 1643 2713
rect 1696 2687 1703 2976
rect 1736 2967 1743 2993
rect 1756 2907 1763 3013
rect 1776 2783 1783 2993
rect 1756 2776 1783 2783
rect 1756 2767 1763 2776
rect 1713 2753 1727 2767
rect 1716 2747 1723 2753
rect 1753 2753 1767 2767
rect 1773 2733 1787 2747
rect 1776 2723 1783 2733
rect 1756 2716 1783 2723
rect 1656 2567 1663 2573
rect 1653 2553 1667 2567
rect 1673 2533 1687 2547
rect 1716 2547 1723 2573
rect 1713 2533 1727 2547
rect 1676 2527 1683 2533
rect 1733 2253 1747 2267
rect 1736 2223 1743 2253
rect 1716 2216 1743 2223
rect 1716 2147 1723 2216
rect 1756 2187 1763 2716
rect 1776 2707 1783 2716
rect 1796 2667 1803 2893
rect 1816 2787 1823 3053
rect 1856 3047 1863 3233
rect 1876 3187 1883 3233
rect 1913 3233 1927 3247
rect 1933 3213 1947 3227
rect 1876 3167 1883 3173
rect 1936 3067 1943 3213
rect 1956 3087 1963 3253
rect 1973 3233 1987 3247
rect 1976 3227 1983 3233
rect 1993 3213 2007 3227
rect 2033 3223 2047 3227
rect 2056 3223 2063 3333
rect 2097 3278 2105 3302
rect 2033 3216 2063 3223
rect 2033 3213 2047 3216
rect 1996 3207 2003 3213
rect 1913 3043 1927 3047
rect 1836 2987 1843 3033
rect 1893 3013 1907 3027
rect 1913 3036 1943 3043
rect 1913 3033 1927 3036
rect 1896 3007 1903 3013
rect 1916 2967 1923 2993
rect 1813 2733 1827 2747
rect 1816 2687 1823 2733
rect 1876 2743 1883 2773
rect 1936 2767 1943 3036
rect 1953 3033 1967 3047
rect 1956 2987 1963 3033
rect 1977 2996 1985 3076
rect 1977 2958 1985 2982
rect 1996 2807 2003 3053
rect 2036 3047 2043 3153
rect 2033 3043 2047 3047
rect 2016 3036 2047 3043
rect 1956 2767 1963 2773
rect 1867 2736 1883 2743
rect 1893 2733 1907 2747
rect 1953 2763 1967 2767
rect 1953 2756 1983 2763
rect 1953 2753 1967 2756
rect 1797 2516 1805 2596
rect 1816 2567 1823 2673
rect 1856 2567 1863 2613
rect 1896 2567 1903 2733
rect 1976 2743 1983 2756
rect 1993 2743 2007 2747
rect 1976 2736 2007 2743
rect 1993 2733 2007 2736
rect 1933 2713 1947 2727
rect 1893 2553 1907 2567
rect 1797 2478 1805 2502
rect 1773 2253 1787 2267
rect 1776 2207 1783 2253
rect 1896 2247 1903 2313
rect 1813 2233 1827 2247
rect 1816 2167 1823 2233
rect 1656 2107 1663 2113
rect 1653 2093 1667 2107
rect 1716 2087 1723 2133
rect 1713 2083 1727 2087
rect 1673 2063 1687 2067
rect 1696 2076 1727 2083
rect 1696 2063 1703 2076
rect 1673 2056 1703 2063
rect 1713 2073 1727 2076
rect 1673 2053 1687 2056
rect 1736 1947 1743 2113
rect 1756 2087 1763 2113
rect 1776 2087 1783 2153
rect 1836 2147 1843 2233
rect 1753 2073 1767 2087
rect 1817 2036 1825 2116
rect 1856 2087 1863 2233
rect 1916 2167 1923 2713
rect 1936 2707 1943 2713
rect 1936 2484 1944 2596
rect 1996 2267 2003 2653
rect 2016 2627 2023 3036
rect 2033 3033 2047 3036
rect 2013 2533 2027 2547
rect 2016 2307 2023 2533
rect 2016 2287 2023 2293
rect 2013 2273 2027 2287
rect 1973 2253 1987 2267
rect 1876 2087 1883 2093
rect 1873 2073 1887 2087
rect 1817 1998 1825 2022
rect 1416 1347 1423 1373
rect 1413 1333 1427 1347
rect 1373 1296 1403 1303
rect 1373 1293 1387 1296
rect 1336 1147 1343 1293
rect 1273 1133 1287 1147
rect 1176 1087 1183 1116
rect 1193 1113 1207 1116
rect 1233 1113 1247 1127
rect 1313 1123 1327 1127
rect 1313 1116 1343 1123
rect 1313 1113 1327 1116
rect 1296 1087 1303 1093
rect 1156 896 1183 903
rect 1156 863 1163 873
rect 1136 856 1163 863
rect 916 847 923 853
rect 876 667 883 833
rect 893 813 907 827
rect 913 833 927 847
rect 973 843 987 847
rect 933 823 947 827
rect 956 836 987 843
rect 956 823 963 836
rect 933 816 963 823
rect 973 833 987 836
rect 1016 823 1023 853
rect 1033 823 1047 827
rect 933 813 947 816
rect 896 807 903 813
rect 1016 816 1047 823
rect 1033 813 1047 816
rect 993 793 1007 807
rect 1093 813 1107 827
rect 1133 823 1147 827
rect 1156 823 1163 856
rect 1053 793 1067 807
rect 996 787 1003 793
rect 836 656 863 663
rect 756 407 763 413
rect 836 407 843 656
rect 873 643 887 647
rect 856 636 887 643
rect 856 627 863 636
rect 873 633 887 636
rect 936 627 943 693
rect 1016 667 1023 673
rect 1056 667 1063 793
rect 1096 787 1103 813
rect 1133 816 1163 823
rect 1133 813 1147 816
rect 1013 653 1027 667
rect 956 627 963 653
rect 996 647 1003 653
rect 993 633 1007 647
rect 933 613 947 627
rect 1076 647 1083 653
rect 496 387 503 393
rect 493 373 507 387
rect 453 363 467 367
rect 413 333 427 347
rect 453 356 483 363
rect 453 353 467 356
rect 416 323 423 333
rect 396 316 423 323
rect 476 327 483 356
rect 556 343 563 393
rect 536 336 563 343
rect 336 167 343 193
rect 356 167 363 173
rect 376 167 383 273
rect 396 187 403 316
rect 433 313 447 327
rect 436 287 443 313
rect 393 173 407 187
rect 213 156 243 163
rect 213 153 227 156
rect 273 133 287 147
rect 333 153 347 167
rect 373 153 387 167
rect 416 167 423 173
rect 276 127 283 133
rect 356 127 363 153
rect 413 153 427 167
rect 436 147 443 213
rect 456 147 463 273
rect 516 187 523 213
rect 496 147 503 173
rect 453 133 467 147
rect 513 123 527 127
rect 536 123 543 336
rect 576 307 583 373
rect 636 367 643 393
rect 796 387 803 393
rect 633 353 647 367
rect 673 333 687 347
rect 713 343 727 347
rect 713 336 733 343
rect 713 333 727 336
rect 656 327 663 333
rect 676 327 683 333
rect 756 327 763 373
rect 796 367 803 373
rect 793 353 807 367
rect 813 333 827 347
rect 816 307 823 333
rect 836 307 843 333
rect 556 143 563 193
rect 616 167 623 193
rect 636 187 643 213
rect 716 187 723 193
rect 633 173 647 187
rect 713 173 727 187
rect 573 143 587 147
rect 556 136 587 143
rect 613 153 627 167
rect 676 167 683 173
rect 673 153 687 167
rect 573 133 587 136
rect 733 143 747 147
rect 756 143 763 213
rect 773 153 787 167
rect 733 136 763 143
rect 733 133 747 136
rect 513 116 543 123
rect 513 113 527 116
rect 195 78 203 102
rect 776 107 783 153
rect 797 116 805 196
rect 856 167 863 433
rect 876 363 883 393
rect 1036 387 1043 593
rect 1096 403 1103 633
rect 1113 613 1127 627
rect 1116 407 1123 613
rect 1076 396 1103 403
rect 1076 387 1083 396
rect 1136 387 1143 673
rect 1176 647 1183 896
rect 1196 867 1203 893
rect 1193 853 1207 867
rect 1213 833 1227 847
rect 1216 827 1223 833
rect 1256 827 1263 1053
rect 1313 863 1327 867
rect 1336 863 1343 1116
rect 1396 1044 1404 1156
rect 1356 867 1363 893
rect 1396 867 1403 893
rect 1293 833 1307 847
rect 1313 856 1343 863
rect 1313 853 1327 856
rect 1353 853 1367 867
rect 1393 853 1407 867
rect 1196 647 1203 693
rect 1236 647 1243 713
rect 1296 667 1303 833
rect 1416 803 1423 1273
rect 1436 1127 1443 1133
rect 1476 1127 1483 1613
rect 1556 1524 1564 1636
rect 1576 1563 1583 1793
rect 1616 1744 1624 1856
rect 1693 1773 1707 1787
rect 1696 1707 1703 1773
rect 1736 1767 1743 1933
rect 1755 1838 1763 1862
rect 1896 1827 1903 2153
rect 1916 2087 1923 2133
rect 1913 2073 1927 2087
rect 1936 2067 1943 2173
rect 1976 2147 1983 2253
rect 1956 2004 1964 2116
rect 1976 2047 1983 2133
rect 2036 2103 2043 2653
rect 2056 2123 2063 3216
rect 2097 3184 2105 3264
rect 2116 3187 2123 3213
rect 2116 2964 2124 3076
rect 2136 2987 2143 3553
rect 2156 3263 2163 3573
rect 2236 3547 2243 3736
rect 2256 3707 2263 3933
rect 2336 3907 2343 4013
rect 2413 3973 2427 3987
rect 2416 3907 2423 3973
rect 2436 3767 2443 4313
rect 2473 4193 2487 4207
rect 2476 4147 2483 4193
rect 2493 4173 2507 4187
rect 2533 4173 2547 4187
rect 2496 4107 2503 4173
rect 2536 4127 2543 4173
rect 2556 4087 2563 4213
rect 2596 4207 2603 4433
rect 2636 4387 2643 4476
rect 2653 4473 2667 4476
rect 2693 4473 2707 4487
rect 2733 4483 2747 4487
rect 2733 4476 2763 4483
rect 2733 4473 2747 4476
rect 2636 4207 2643 4213
rect 2613 4173 2627 4187
rect 2633 4193 2647 4207
rect 2456 3967 2463 3973
rect 2496 3947 2503 3993
rect 2516 3987 2523 4013
rect 2536 4007 2543 4033
rect 2576 4007 2583 4013
rect 2533 3993 2547 4007
rect 2513 3973 2527 3987
rect 2573 3993 2587 4007
rect 2596 3967 2603 4133
rect 2616 4087 2623 4173
rect 2693 4183 2707 4187
rect 2716 4183 2723 4273
rect 2756 4223 2763 4476
rect 2773 4473 2787 4487
rect 2693 4176 2723 4183
rect 2736 4216 2763 4223
rect 2693 4173 2707 4176
rect 2653 4153 2667 4167
rect 2656 4147 2663 4153
rect 2613 3953 2627 3967
rect 2656 3967 2663 4053
rect 2676 4007 2683 4153
rect 2736 4107 2743 4216
rect 2796 4207 2803 4573
rect 2836 4487 2843 4623
rect 2876 4587 2883 4623
rect 2833 4473 2847 4487
rect 2873 4483 2887 4487
rect 2856 4476 2887 4483
rect 2856 4327 2863 4476
rect 2873 4473 2887 4476
rect 2816 4207 2823 4293
rect 2896 4263 2903 4473
rect 2936 4467 2943 4533
rect 3076 4487 3083 4533
rect 3116 4487 3123 4623
rect 3156 4567 3163 4623
rect 3456 4507 3463 4513
rect 3453 4493 3467 4507
rect 2913 4433 2927 4447
rect 2933 4453 2947 4467
rect 2987 4456 3003 4463
rect 3073 4473 3087 4487
rect 2996 4447 3003 4456
rect 3113 4473 3127 4487
rect 3153 4483 3167 4487
rect 3153 4476 3183 4483
rect 3153 4473 3167 4476
rect 2916 4307 2923 4433
rect 2896 4256 2923 4263
rect 2753 4173 2767 4187
rect 2756 4127 2763 4173
rect 2833 4173 2847 4187
rect 2696 4047 2703 4093
rect 2836 4067 2843 4173
rect 2716 4023 2723 4033
rect 2756 4027 2763 4033
rect 2696 4016 2723 4023
rect 2673 3983 2687 3987
rect 2696 3983 2703 4016
rect 2856 4023 2863 4253
rect 2896 4167 2903 4233
rect 2916 4207 2923 4256
rect 2936 4227 2943 4293
rect 2996 4267 3003 4293
rect 2933 4213 2947 4227
rect 2973 4213 2987 4227
rect 2896 4087 2903 4093
rect 2673 3976 2703 3983
rect 2836 4016 2863 4023
rect 2836 4007 2843 4016
rect 2896 4007 2903 4073
rect 2916 4027 2923 4173
rect 2976 4147 2983 4213
rect 2993 4203 3007 4207
rect 3016 4203 3023 4413
rect 3036 4247 3043 4433
rect 3116 4227 3123 4253
rect 3156 4227 3163 4393
rect 2993 4196 3023 4203
rect 2993 4193 3007 4196
rect 3093 4193 3107 4207
rect 3113 4213 3127 4227
rect 3153 4213 3167 4227
rect 3096 4187 3103 4193
rect 2976 4087 2983 4133
rect 2833 3993 2847 4007
rect 2673 3973 2687 3976
rect 2773 3973 2787 3987
rect 2813 3983 2827 3987
rect 2796 3976 2827 3983
rect 2596 3927 2603 3933
rect 2616 3907 2623 3953
rect 2696 3787 2703 3953
rect 2333 3693 2347 3707
rect 2336 3567 2343 3693
rect 2356 3663 2363 3753
rect 2393 3713 2407 3727
rect 2396 3667 2403 3713
rect 2416 3687 2423 3733
rect 2356 3656 2383 3663
rect 2213 3543 2227 3547
rect 2213 3536 2233 3543
rect 2213 3533 2227 3536
rect 2296 3507 2303 3533
rect 2233 3493 2247 3507
rect 2196 3287 2203 3493
rect 2236 3487 2243 3493
rect 2273 3473 2287 3487
rect 2293 3493 2307 3507
rect 2356 3503 2363 3633
rect 2376 3547 2383 3656
rect 2396 3567 2403 3613
rect 2396 3547 2403 3553
rect 2436 3547 2443 3713
rect 2456 3587 2463 3753
rect 2556 3747 2563 3773
rect 2533 3723 2547 3727
rect 2533 3716 2563 3723
rect 2613 3733 2627 3747
rect 2533 3713 2547 3716
rect 2556 3703 2563 3716
rect 2593 3713 2607 3727
rect 2596 3707 2603 3713
rect 2556 3696 2583 3703
rect 2393 3533 2407 3547
rect 2373 3503 2387 3507
rect 2356 3496 2387 3503
rect 2373 3493 2387 3496
rect 2276 3467 2283 3473
rect 2416 3327 2423 3533
rect 2456 3507 2463 3553
rect 2496 3507 2503 3613
rect 2516 3507 2523 3673
rect 2556 3627 2563 3673
rect 2576 3667 2583 3696
rect 2596 3667 2603 3693
rect 2616 3687 2623 3733
rect 2696 3727 2703 3733
rect 2693 3713 2707 3727
rect 2736 3707 2743 3973
rect 2713 3693 2727 3707
rect 2576 3587 2583 3653
rect 2556 3507 2563 3513
rect 2453 3493 2467 3507
rect 2493 3493 2507 3507
rect 2553 3493 2567 3507
rect 2576 3487 2583 3573
rect 2573 3473 2587 3487
rect 2156 3256 2183 3263
rect 2153 3213 2167 3227
rect 2156 3167 2163 3213
rect 2176 2847 2183 3256
rect 2193 3213 2207 3227
rect 2196 3207 2203 3213
rect 2216 3083 2223 3273
rect 2236 3184 2244 3296
rect 2196 3076 2223 3083
rect 2196 3047 2203 3076
rect 2193 3033 2207 3047
rect 2236 3047 2243 3053
rect 2233 3033 2247 3047
rect 2216 2927 2223 3013
rect 2256 3003 2263 3293
rect 2296 3103 2303 3313
rect 2316 3247 2323 3273
rect 2433 3263 2447 3267
rect 2416 3256 2447 3263
rect 2313 3233 2327 3247
rect 2333 3193 2347 3207
rect 2393 3193 2407 3207
rect 2296 3096 2323 3103
rect 2296 3067 2303 3073
rect 2293 3053 2307 3067
rect 2273 3013 2287 3027
rect 2316 3023 2323 3096
rect 2336 3047 2343 3193
rect 2296 3016 2323 3023
rect 2236 2996 2263 3003
rect 2076 2787 2083 2813
rect 2073 2773 2087 2787
rect 2113 2773 2127 2787
rect 2116 2767 2123 2773
rect 2133 2753 2147 2767
rect 2136 2743 2143 2753
rect 2116 2736 2143 2743
rect 2116 2527 2123 2736
rect 2156 2723 2163 2733
rect 2136 2716 2163 2723
rect 2136 2607 2143 2716
rect 2056 2116 2083 2123
rect 2016 2096 2043 2103
rect 1755 1744 1763 1824
rect 1896 1807 1903 1813
rect 1773 1783 1787 1787
rect 1773 1776 1803 1783
rect 1773 1773 1787 1776
rect 1796 1767 1803 1776
rect 1893 1793 1907 1807
rect 1913 1773 1927 1787
rect 1916 1767 1923 1773
rect 1953 1773 1967 1787
rect 1873 1753 1887 1767
rect 1876 1727 1883 1753
rect 1636 1627 1643 1693
rect 1636 1607 1643 1613
rect 1633 1593 1647 1607
rect 1576 1556 1603 1563
rect 1695 1556 1703 1636
rect 1816 1627 1823 1713
rect 1876 1627 1883 1633
rect 1813 1613 1827 1627
rect 1713 1593 1727 1607
rect 1716 1587 1723 1593
rect 1873 1613 1887 1627
rect 1793 1573 1807 1587
rect 1896 1607 1903 1713
rect 1916 1667 1923 1753
rect 1956 1727 1963 1773
rect 1976 1687 1983 1853
rect 2016 1827 2023 2096
rect 2036 1867 2043 2053
rect 2076 1847 2083 2116
rect 2116 2067 2123 2193
rect 2136 2127 2143 2593
rect 2176 2587 2183 2813
rect 2216 2787 2223 2853
rect 2193 2733 2207 2747
rect 2196 2707 2203 2733
rect 2216 2527 2223 2713
rect 2236 2667 2243 2996
rect 2256 2727 2263 2973
rect 2276 2867 2283 3013
rect 2296 2867 2303 3016
rect 2333 2993 2347 3007
rect 2376 3007 2383 3133
rect 2396 3127 2403 3193
rect 2416 3107 2423 3256
rect 2433 3253 2447 3256
rect 2473 3253 2487 3267
rect 2476 3187 2483 3253
rect 2493 3243 2507 3247
rect 2513 3243 2527 3247
rect 2493 3236 2527 3243
rect 2493 3233 2507 3236
rect 2513 3233 2527 3236
rect 2496 3227 2503 3233
rect 2573 3223 2587 3227
rect 2596 3223 2603 3453
rect 2573 3216 2603 3223
rect 2573 3213 2587 3216
rect 2533 3193 2547 3207
rect 2536 3187 2543 3193
rect 2556 3167 2563 3193
rect 2476 3067 2483 3093
rect 2473 3053 2487 3067
rect 2436 3047 2443 3053
rect 2433 3033 2447 3047
rect 2393 3023 2407 3027
rect 2393 3016 2423 3023
rect 2393 3013 2407 3016
rect 2373 2993 2387 3007
rect 2336 2947 2343 2993
rect 2416 2967 2423 3016
rect 2516 2987 2523 3093
rect 2556 3027 2563 3093
rect 2576 3027 2583 3153
rect 2596 3067 2603 3073
rect 2596 3047 2603 3053
rect 2596 3027 2603 3033
rect 2593 3013 2607 3027
rect 2276 2704 2284 2816
rect 2236 2484 2244 2596
rect 2276 2567 2283 2593
rect 2273 2553 2287 2567
rect 2156 2287 2163 2293
rect 2153 2273 2167 2287
rect 2176 2247 2183 2313
rect 2216 2287 2223 2373
rect 2193 2253 2207 2267
rect 2213 2273 2227 2287
rect 2253 2273 2267 2287
rect 2156 2087 2163 2113
rect 2153 2073 2167 2087
rect 2093 2033 2107 2047
rect 2113 2053 2127 2067
rect 2176 2047 2183 2233
rect 2196 2147 2203 2253
rect 2256 2207 2263 2273
rect 2193 2083 2207 2087
rect 2193 2076 2223 2083
rect 2193 2073 2207 2076
rect 2096 2027 2103 2033
rect 2096 1987 2103 2013
rect 2216 2007 2223 2076
rect 2233 2033 2247 2047
rect 2236 2027 2243 2033
rect 2076 1807 2083 1833
rect 2176 1807 2183 1933
rect 2296 1807 2303 2833
rect 2313 2733 2327 2747
rect 2353 2733 2367 2747
rect 2316 2687 2323 2733
rect 2356 2567 2363 2733
rect 2396 2603 2403 2893
rect 2415 2798 2423 2822
rect 2415 2704 2423 2784
rect 2436 2747 2443 2933
rect 2456 2627 2463 2853
rect 2536 2767 2543 2833
rect 2556 2787 2563 2813
rect 2616 2807 2623 3613
rect 2656 3527 2663 3593
rect 2716 3527 2723 3693
rect 2756 3627 2763 3973
rect 2776 3967 2783 3973
rect 2796 3947 2803 3976
rect 2813 3973 2827 3976
rect 2853 3973 2867 3987
rect 2893 3993 2907 4007
rect 2956 3987 2963 4013
rect 2953 3973 2967 3987
rect 2856 3963 2863 3973
rect 2856 3956 2883 3963
rect 2796 3847 2803 3933
rect 2876 3927 2883 3956
rect 2856 3747 2863 3793
rect 2876 3787 2883 3913
rect 2836 3727 2843 3733
rect 2936 3727 2943 3733
rect 2956 3727 2963 3853
rect 2976 3807 2983 4053
rect 2996 3867 3003 4173
rect 3176 4027 3183 4476
rect 3216 4467 3223 4493
rect 3256 4467 3263 4473
rect 3296 4467 3303 4493
rect 3193 4433 3207 4447
rect 3213 4453 3227 4467
rect 3253 4453 3267 4467
rect 3273 4433 3287 4447
rect 3293 4453 3307 4467
rect 3353 4463 3367 4467
rect 3313 4433 3327 4447
rect 3336 4456 3367 4463
rect 3196 4367 3203 4433
rect 3196 4107 3203 4293
rect 3216 4207 3223 4373
rect 3276 4287 3283 4433
rect 3316 4407 3323 4433
rect 3336 4387 3343 4456
rect 3353 4453 3367 4456
rect 3256 4207 3263 4273
rect 3356 4247 3363 4433
rect 3376 4227 3383 4273
rect 3436 4243 3443 4493
rect 3636 4476 3683 4483
rect 3456 4427 3463 4433
rect 3496 4407 3503 4453
rect 3513 4433 3527 4447
rect 3593 4463 3607 4467
rect 3576 4456 3607 4463
rect 3516 4407 3523 4433
rect 3516 4287 3523 4393
rect 3556 4303 3563 4433
rect 3576 4407 3583 4456
rect 3593 4453 3607 4456
rect 3616 4447 3623 4473
rect 3636 4467 3643 4476
rect 3676 4467 3683 4476
rect 3796 4487 3803 4513
rect 3936 4487 3943 4533
rect 4136 4516 4263 4523
rect 3976 4487 3983 4513
rect 4136 4507 4143 4516
rect 3633 4453 3647 4467
rect 3693 4453 3707 4467
rect 3793 4473 3807 4487
rect 3933 4473 3947 4487
rect 3913 4463 3927 4467
rect 3653 4443 3667 4447
rect 3653 4436 3673 4443
rect 3653 4433 3667 4436
rect 3656 4423 3663 4433
rect 3647 4416 3663 4423
rect 3696 4407 3703 4453
rect 3556 4296 3583 4303
rect 3436 4236 3463 4243
rect 3313 4213 3327 4227
rect 3373 4223 3387 4227
rect 3316 4187 3323 4213
rect 3333 4203 3347 4207
rect 3356 4216 3387 4223
rect 3356 4203 3363 4216
rect 3333 4196 3363 4203
rect 3373 4213 3387 4216
rect 3333 4193 3347 4196
rect 3393 4193 3407 4207
rect 3433 4193 3447 4207
rect 3396 4127 3403 4193
rect 3416 4043 3423 4193
rect 3436 4187 3443 4193
rect 3456 4167 3463 4236
rect 3556 4227 3563 4273
rect 3576 4227 3583 4296
rect 3736 4267 3743 4453
rect 3896 4456 3927 4463
rect 3896 4427 3903 4456
rect 3913 4453 3927 4456
rect 3973 4473 3987 4487
rect 3996 4447 4003 4473
rect 4036 4467 4043 4473
rect 4056 4467 4063 4493
rect 4136 4467 4143 4473
rect 4013 4433 4027 4447
rect 4033 4453 4047 4467
rect 4073 4463 4087 4467
rect 4073 4456 4103 4463
rect 4073 4453 4087 4456
rect 3513 4213 3527 4227
rect 3493 4193 3507 4207
rect 3396 4036 3423 4043
rect 3133 4023 3147 4027
rect 3133 4016 3163 4023
rect 3133 4013 3147 4016
rect 3067 3996 3073 4003
rect 2833 3713 2847 3727
rect 2873 3723 2887 3727
rect 2856 3716 2887 3723
rect 2856 3687 2863 3716
rect 2873 3713 2887 3716
rect 2933 3713 2947 3727
rect 2893 3673 2907 3687
rect 2756 3527 2763 3553
rect 2653 3513 2667 3527
rect 2693 3523 2707 3527
rect 2713 3523 2727 3527
rect 2636 3507 2643 3513
rect 2693 3516 2727 3523
rect 2693 3513 2707 3516
rect 2713 3513 2727 3516
rect 2753 3513 2767 3527
rect 2776 3507 2783 3533
rect 2656 3267 2663 3313
rect 2656 3247 2663 3253
rect 2636 3027 2643 3113
rect 2656 3087 2663 3193
rect 2676 3187 2683 3473
rect 2736 3447 2743 3493
rect 2756 3267 2763 3473
rect 2796 3247 2803 3533
rect 2816 3527 2823 3613
rect 2856 3547 2863 3653
rect 2896 3567 2903 3673
rect 2896 3527 2903 3553
rect 2916 3547 2923 3713
rect 2976 3687 2983 3773
rect 2996 3747 3003 3833
rect 2993 3733 3007 3747
rect 3013 3713 3027 3727
rect 3016 3707 3023 3713
rect 2953 3673 2967 3687
rect 2956 3607 2963 3673
rect 2936 3527 2943 3573
rect 2893 3513 2907 3527
rect 2836 3507 2843 3513
rect 2813 3473 2827 3487
rect 2833 3493 2847 3507
rect 2853 3473 2867 3487
rect 2816 3367 2823 3473
rect 2856 3467 2863 3473
rect 2753 3213 2767 3227
rect 2773 3213 2787 3227
rect 2676 3063 2683 3093
rect 2656 3056 2683 3063
rect 2656 3047 2663 3056
rect 2696 3047 2703 3073
rect 2716 3047 2723 3173
rect 2736 3047 2743 3173
rect 2756 3127 2763 3213
rect 2776 3187 2783 3213
rect 2793 3193 2807 3207
rect 2796 3167 2803 3193
rect 2836 3187 2843 3393
rect 2876 3287 2883 3513
rect 2913 3493 2927 3507
rect 2933 3513 2947 3527
rect 2956 3507 2963 3593
rect 2976 3587 2983 3653
rect 2996 3547 3003 3693
rect 3016 3627 3023 3673
rect 3036 3667 3043 3733
rect 3056 3687 3063 3713
rect 2916 3487 2923 3493
rect 2976 3487 2983 3533
rect 3036 3527 3043 3533
rect 3033 3513 3047 3527
rect 2896 3263 2903 3413
rect 2976 3283 2983 3453
rect 2996 3287 3003 3453
rect 3016 3287 3023 3493
rect 3076 3463 3083 3913
rect 3096 3907 3103 4013
rect 3156 4007 3163 4016
rect 3196 4007 3203 4033
rect 3216 4007 3223 4013
rect 3173 3973 3187 3987
rect 3193 3993 3207 4007
rect 3213 3983 3227 3987
rect 3236 3983 3243 4013
rect 3213 3976 3243 3983
rect 3213 3973 3227 3976
rect 3116 3947 3123 3973
rect 3176 3963 3183 3973
rect 3176 3956 3203 3963
rect 3196 3947 3203 3956
rect 3096 3767 3103 3893
rect 3176 3727 3183 3933
rect 3236 3887 3243 3976
rect 3316 4007 3323 4013
rect 3396 4007 3403 4036
rect 3416 4007 3423 4036
rect 3293 3973 3307 3987
rect 3313 3993 3327 4007
rect 3393 3993 3407 4007
rect 3093 3693 3107 3707
rect 3233 3733 3247 3747
rect 3236 3727 3243 3733
rect 3213 3713 3227 3727
rect 3096 3627 3103 3693
rect 3216 3703 3223 3713
rect 3216 3696 3243 3703
rect 3133 3673 3147 3687
rect 3096 3507 3103 3573
rect 3116 3527 3123 3673
rect 3136 3667 3143 3673
rect 3176 3667 3183 3693
rect 3156 3527 3163 3593
rect 3176 3527 3183 3593
rect 3236 3567 3243 3696
rect 3216 3527 3223 3553
rect 3113 3513 3127 3527
rect 3093 3493 3107 3507
rect 3153 3513 3167 3527
rect 3173 3513 3187 3527
rect 3193 3493 3207 3507
rect 3233 3493 3247 3507
rect 3196 3467 3203 3493
rect 3056 3456 3083 3463
rect 3036 3287 3043 3433
rect 3056 3307 3063 3456
rect 2967 3276 2983 3283
rect 2953 3263 2967 3267
rect 2876 3256 2903 3263
rect 2876 3247 2883 3256
rect 2853 3213 2867 3227
rect 2873 3233 2887 3247
rect 2936 3256 2967 3263
rect 2993 3263 3007 3267
rect 3033 3263 3047 3267
rect 2856 3207 2863 3213
rect 2653 3033 2667 3047
rect 2633 3013 2647 3027
rect 2693 3033 2707 3047
rect 2776 3047 2783 3053
rect 2836 3047 2843 3133
rect 2773 3033 2787 3047
rect 2816 3027 2823 3033
rect 2493 2763 2507 2767
rect 2476 2756 2507 2763
rect 2396 2596 2423 2603
rect 2375 2516 2383 2596
rect 2393 2553 2407 2567
rect 2375 2478 2383 2502
rect 2396 2407 2403 2553
rect 2316 2207 2323 2293
rect 2336 2224 2344 2336
rect 2356 2307 2363 2333
rect 2416 2303 2423 2596
rect 2396 2296 2423 2303
rect 2396 2107 2403 2296
rect 2413 2263 2427 2267
rect 2436 2263 2443 2553
rect 2476 2547 2483 2756
rect 2493 2753 2507 2756
rect 2513 2733 2527 2747
rect 2533 2753 2547 2767
rect 2553 2733 2567 2747
rect 2516 2687 2523 2733
rect 2556 2707 2563 2733
rect 2576 2707 2583 2773
rect 2636 2767 2643 2913
rect 2716 2827 2723 3013
rect 2793 2993 2807 3007
rect 2776 2807 2783 2993
rect 2796 2867 2803 2993
rect 2856 2983 2863 3193
rect 2916 3043 2923 3213
rect 2936 3207 2943 3256
rect 2953 3253 2967 3256
rect 2993 3256 3047 3263
rect 3073 3263 3087 3267
rect 3096 3263 3103 3373
rect 3116 3347 3123 3433
rect 3236 3423 3243 3493
rect 3216 3416 3243 3423
rect 2993 3253 3007 3256
rect 3016 3207 3023 3256
rect 3033 3253 3047 3256
rect 3073 3256 3103 3263
rect 3073 3253 3087 3256
rect 2956 3047 2963 3193
rect 3016 3087 3023 3193
rect 2996 3047 3003 3073
rect 3036 3067 3043 3193
rect 3056 3167 3063 3233
rect 2953 3043 2967 3047
rect 2907 3036 2923 3043
rect 2936 3036 2967 3043
rect 2913 2993 2927 3007
rect 2836 2976 2863 2983
rect 2756 2767 2763 2793
rect 2816 2787 2823 2813
rect 2836 2787 2843 2976
rect 2876 2963 2883 2993
rect 2916 2987 2923 2993
rect 2867 2956 2883 2963
rect 2856 2787 2863 2953
rect 2896 2807 2903 2973
rect 2916 2847 2923 2873
rect 2936 2867 2943 3036
rect 2953 3033 2967 3036
rect 2993 3033 3007 3047
rect 3056 3027 3063 3133
rect 3076 3107 3083 3213
rect 3096 3183 3103 3256
rect 3116 3223 3123 3273
rect 3156 3267 3163 3333
rect 3176 3247 3183 3293
rect 3216 3267 3223 3416
rect 3276 3347 3283 3953
rect 3296 3947 3303 3973
rect 3336 3967 3343 3973
rect 3296 3727 3303 3873
rect 3336 3723 3343 3953
rect 3376 3747 3383 3953
rect 3396 3727 3403 3933
rect 3416 3907 3423 3933
rect 3353 3723 3367 3727
rect 3336 3716 3367 3723
rect 3353 3713 3367 3716
rect 3313 3673 3327 3687
rect 3316 3627 3323 3673
rect 3356 3627 3363 3713
rect 3316 3507 3323 3573
rect 3336 3547 3343 3573
rect 3376 3567 3383 3673
rect 3416 3667 3423 3693
rect 3396 3527 3403 3593
rect 3416 3527 3423 3633
rect 3293 3473 3307 3487
rect 3313 3493 3327 3507
rect 3333 3473 3347 3487
rect 3296 3463 3303 3473
rect 3296 3456 3323 3463
rect 3296 3347 3303 3373
rect 3236 3267 3243 3313
rect 3316 3267 3323 3456
rect 3336 3387 3343 3473
rect 3356 3287 3363 3513
rect 3436 3507 3443 4153
rect 3476 4087 3483 4173
rect 3496 4143 3503 4193
rect 3516 4167 3523 4213
rect 3573 4213 3587 4227
rect 3533 4193 3547 4207
rect 3593 4193 3607 4207
rect 3536 4147 3543 4193
rect 3496 4136 3523 4143
rect 3496 4007 3503 4113
rect 3516 4027 3523 4136
rect 3536 4007 3543 4113
rect 3596 4107 3603 4193
rect 3493 3993 3507 4007
rect 3476 3987 3483 3993
rect 3473 3973 3487 3987
rect 3513 3973 3527 3987
rect 3533 3993 3547 4007
rect 3456 3927 3463 3953
rect 3516 3927 3523 3973
rect 3556 3767 3563 4073
rect 3576 3987 3583 4013
rect 3596 4007 3603 4093
rect 3616 4047 3623 4213
rect 3633 4193 3647 4207
rect 3673 4213 3687 4227
rect 3713 4223 3727 4227
rect 3636 4187 3643 4193
rect 3676 4167 3683 4213
rect 3713 4216 3743 4223
rect 3713 4213 3727 4216
rect 3636 4007 3643 4113
rect 3593 3993 3607 4007
rect 3573 3973 3587 3987
rect 3613 3973 3627 3987
rect 3576 3747 3583 3913
rect 3596 3903 3603 3953
rect 3616 3927 3623 3973
rect 3656 3967 3663 4133
rect 3676 4027 3683 4153
rect 3696 4147 3703 4193
rect 3736 4187 3743 4216
rect 3796 4207 3803 4213
rect 3793 4193 3807 4207
rect 3836 4047 3843 4293
rect 3853 4173 3867 4187
rect 3913 4193 3927 4207
rect 3893 4173 3907 4187
rect 3856 4087 3863 4173
rect 3896 4147 3903 4173
rect 3916 4167 3923 4193
rect 3693 3973 3707 3987
rect 3596 3896 3623 3903
rect 3553 3743 3567 3747
rect 3547 3736 3567 3743
rect 3553 3733 3567 3736
rect 3513 3703 3527 3707
rect 3507 3696 3527 3703
rect 3513 3693 3527 3696
rect 3476 3507 3483 3613
rect 3496 3527 3503 3693
rect 3536 3623 3543 3733
rect 3573 3703 3587 3707
rect 3596 3703 3603 3753
rect 3573 3696 3603 3703
rect 3573 3693 3587 3696
rect 3516 3616 3543 3623
rect 3373 3473 3387 3487
rect 3453 3473 3467 3487
rect 3473 3493 3487 3507
rect 3376 3307 3383 3473
rect 3456 3467 3463 3473
rect 3396 3367 3403 3453
rect 3416 3447 3423 3453
rect 3496 3447 3503 3453
rect 3456 3367 3463 3433
rect 3516 3427 3523 3616
rect 3536 3547 3543 3573
rect 3556 3547 3563 3553
rect 3616 3547 3623 3896
rect 3636 3747 3643 3953
rect 3696 3907 3703 3973
rect 3553 3533 3567 3547
rect 3536 3527 3543 3533
rect 3533 3513 3547 3527
rect 3573 3523 3587 3527
rect 3573 3516 3603 3523
rect 3573 3513 3587 3516
rect 3596 3507 3603 3516
rect 3636 3507 3643 3533
rect 3233 3253 3247 3267
rect 3196 3247 3203 3253
rect 3133 3223 3147 3227
rect 3116 3216 3147 3223
rect 3193 3233 3207 3247
rect 3133 3213 3147 3216
rect 3096 3176 3143 3183
rect 3096 3027 3103 3113
rect 2976 2987 2983 3013
rect 3093 3013 3107 3027
rect 3113 3003 3127 3007
rect 3136 3003 3143 3176
rect 3156 3167 3163 3193
rect 3216 3167 3223 3233
rect 3176 3087 3183 3113
rect 3196 3047 3203 3093
rect 3173 3013 3187 3027
rect 3193 3033 3207 3047
rect 3216 3027 3223 3093
rect 3213 3013 3227 3027
rect 3113 2996 3143 3003
rect 3176 3003 3183 3013
rect 3176 2996 3203 3003
rect 3113 2993 3127 2996
rect 2633 2753 2647 2767
rect 2653 2733 2667 2747
rect 2673 2733 2687 2747
rect 2813 2773 2827 2787
rect 2873 2753 2887 2767
rect 2713 2743 2727 2747
rect 2713 2736 2733 2743
rect 2713 2733 2727 2736
rect 2656 2707 2663 2733
rect 2556 2687 2563 2693
rect 2676 2687 2683 2733
rect 2716 2687 2723 2693
rect 2516 2587 2523 2653
rect 2656 2647 2663 2673
rect 2453 2513 2467 2527
rect 2473 2533 2487 2547
rect 2533 2533 2547 2547
rect 2493 2513 2507 2527
rect 2456 2467 2463 2513
rect 2456 2427 2463 2453
rect 2496 2347 2503 2513
rect 2516 2367 2523 2533
rect 2536 2387 2543 2533
rect 2556 2363 2563 2533
rect 2576 2407 2583 2573
rect 2616 2567 2623 2593
rect 2656 2567 2663 2633
rect 2613 2553 2627 2567
rect 2653 2553 2667 2567
rect 2536 2356 2563 2363
rect 2475 2318 2483 2342
rect 2516 2323 2523 2353
rect 2496 2316 2523 2323
rect 2413 2256 2443 2263
rect 2413 2253 2427 2256
rect 2475 2224 2483 2304
rect 2496 2267 2503 2316
rect 2536 2287 2543 2356
rect 2596 2307 2603 2333
rect 2616 2307 2623 2413
rect 2716 2387 2723 2673
rect 2756 2603 2763 2733
rect 2836 2667 2843 2753
rect 2876 2727 2883 2753
rect 2916 2743 2923 2833
rect 2956 2767 2963 2833
rect 2896 2736 2923 2743
rect 2876 2707 2883 2713
rect 2896 2667 2903 2736
rect 2953 2753 2967 2767
rect 2993 2753 3007 2767
rect 2736 2596 2763 2603
rect 2736 2403 2743 2596
rect 2793 2513 2807 2527
rect 2756 2427 2763 2513
rect 2736 2396 2763 2403
rect 2656 2307 2663 2313
rect 2593 2293 2607 2307
rect 2613 2293 2627 2307
rect 2633 2273 2647 2287
rect 2653 2293 2667 2307
rect 2493 2253 2507 2267
rect 2636 2247 2643 2273
rect 2476 2107 2483 2113
rect 2316 1927 2323 2093
rect 2393 2083 2407 2087
rect 2373 2053 2387 2067
rect 2393 2076 2423 2083
rect 2393 2073 2407 2076
rect 2376 2047 2383 2053
rect 2416 1887 2423 2076
rect 2456 2067 2463 2073
rect 2453 2053 2467 2067
rect 2496 2047 2503 2213
rect 2553 2033 2567 2047
rect 2436 1987 2443 2033
rect 2317 1838 2325 1862
rect 2013 1783 2027 1787
rect 1996 1776 2027 1783
rect 2073 1793 2087 1807
rect 1893 1593 1907 1607
rect 1596 1527 1603 1556
rect 1695 1518 1703 1542
rect 1536 1327 1543 1373
rect 1513 1293 1527 1307
rect 1533 1313 1547 1327
rect 1553 1293 1567 1307
rect 1433 1113 1447 1127
rect 1473 1113 1487 1127
rect 1456 847 1463 893
rect 1496 847 1503 873
rect 1453 833 1467 847
rect 1493 833 1507 847
rect 1416 796 1443 803
rect 1436 747 1443 796
rect 1193 633 1207 647
rect 1233 633 1247 647
rect 1293 603 1307 607
rect 1316 603 1323 673
rect 1336 647 1343 693
rect 1356 647 1363 673
rect 1376 667 1383 713
rect 1373 653 1387 667
rect 1333 633 1347 647
rect 1353 633 1367 647
rect 1396 647 1403 693
rect 1436 647 1443 733
rect 1516 647 1523 1293
rect 1556 1267 1563 1293
rect 1535 1076 1543 1156
rect 1535 1038 1543 1062
rect 1556 927 1563 1113
rect 1576 1047 1583 1293
rect 1596 1067 1603 1513
rect 1656 1367 1663 1373
rect 1716 1363 1723 1573
rect 1796 1567 1803 1573
rect 1696 1356 1723 1363
rect 1656 1347 1663 1353
rect 1696 1347 1703 1356
rect 1653 1333 1667 1347
rect 1693 1333 1707 1347
rect 1676 1107 1683 1133
rect 1673 1093 1687 1107
rect 1553 863 1567 867
rect 1553 856 1583 863
rect 1553 853 1567 856
rect 1533 813 1547 827
rect 1536 807 1543 813
rect 1576 687 1583 856
rect 1616 847 1623 873
rect 1656 847 1663 853
rect 1593 813 1607 827
rect 1613 833 1627 847
rect 1653 833 1667 847
rect 1596 807 1603 813
rect 1673 813 1687 827
rect 1596 787 1603 793
rect 1393 633 1407 647
rect 1433 633 1447 647
rect 1473 643 1487 647
rect 1473 636 1503 643
rect 1473 633 1487 636
rect 1293 596 1323 603
rect 1293 593 1307 596
rect 1496 407 1503 636
rect 1556 564 1564 676
rect 1636 647 1643 653
rect 1633 633 1647 647
rect 1033 383 1047 387
rect 1016 376 1047 383
rect 893 363 907 367
rect 876 356 907 363
rect 893 353 907 356
rect 913 343 927 347
rect 896 336 927 343
rect 896 167 903 336
rect 913 333 927 336
rect 956 327 963 333
rect 1016 347 1023 376
rect 1033 373 1047 376
rect 1053 353 1067 367
rect 1073 373 1087 387
rect 973 313 987 327
rect 853 153 867 167
rect 816 127 823 153
rect 893 153 907 167
rect 797 78 805 102
rect 936 84 944 196
rect 976 107 983 313
rect 1056 307 1063 353
rect 1096 347 1103 373
rect 1016 147 1023 273
rect 1116 247 1123 373
rect 1196 367 1203 393
rect 1336 367 1343 373
rect 1193 353 1207 367
rect 1293 353 1307 367
rect 1173 323 1187 327
rect 1296 327 1303 353
rect 1333 353 1347 367
rect 1353 333 1367 347
rect 1376 343 1383 393
rect 1596 387 1603 393
rect 1656 387 1663 753
rect 1676 707 1683 813
rect 1696 767 1703 1073
rect 1716 683 1723 1333
rect 1773 1293 1787 1307
rect 1736 1127 1743 1213
rect 1776 1207 1783 1293
rect 1816 1287 1823 1293
rect 1836 1267 1843 1573
rect 1916 1567 1923 1633
rect 1936 1587 1943 1673
rect 1877 1358 1885 1382
rect 1877 1264 1885 1344
rect 1933 1303 1947 1307
rect 1956 1303 1963 1613
rect 1976 1524 1984 1636
rect 1996 1603 2003 1776
rect 2013 1773 2027 1776
rect 2053 1753 2067 1767
rect 2056 1727 2063 1753
rect 2096 1747 2103 1793
rect 2113 1773 2127 1787
rect 2116 1727 2123 1773
rect 2153 1773 2167 1787
rect 2173 1793 2187 1807
rect 2156 1767 2163 1773
rect 2293 1783 2307 1787
rect 2276 1776 2307 1783
rect 2276 1767 2283 1776
rect 2293 1773 2307 1776
rect 2193 1753 2207 1767
rect 2013 1603 2027 1607
rect 1996 1596 2027 1603
rect 2013 1593 2027 1596
rect 1933 1296 1963 1303
rect 1933 1293 1947 1296
rect 1896 1227 1903 1293
rect 1756 1147 1763 1153
rect 1753 1133 1767 1147
rect 1773 1123 1787 1127
rect 1773 1116 1803 1123
rect 1773 1113 1787 1116
rect 1796 1087 1803 1116
rect 1736 847 1743 1053
rect 1856 1044 1864 1156
rect 1896 1127 1903 1193
rect 1893 1113 1907 1127
rect 1733 833 1747 847
rect 1716 676 1743 683
rect 1695 596 1703 676
rect 1713 643 1727 647
rect 1736 643 1743 676
rect 1756 647 1763 1033
rect 1873 843 1887 847
rect 1856 836 1887 843
rect 1713 636 1743 643
rect 1713 633 1727 636
rect 1695 558 1703 582
rect 1677 398 1685 422
rect 1393 343 1407 347
rect 1376 336 1407 343
rect 1393 333 1407 336
rect 1173 316 1203 323
rect 1173 313 1187 316
rect 1073 163 1087 167
rect 1013 133 1027 147
rect 1073 156 1103 163
rect 1073 153 1087 156
rect 1096 143 1103 156
rect 1156 147 1163 233
rect 1176 167 1183 193
rect 1196 187 1203 316
rect 1253 313 1267 327
rect 1173 153 1187 167
rect 1216 167 1223 293
rect 1256 287 1263 313
rect 1356 307 1363 333
rect 1433 333 1447 347
rect 1593 373 1607 387
rect 1736 387 1743 636
rect 1753 633 1767 647
rect 1656 347 1663 373
rect 1653 333 1667 347
rect 1113 143 1127 147
rect 1096 136 1127 143
rect 1113 133 1127 136
rect 1236 143 1243 193
rect 1336 167 1343 213
rect 1376 167 1383 213
rect 1436 187 1443 333
rect 1677 304 1685 384
rect 1776 383 1783 653
rect 1836 643 1843 693
rect 1856 667 1863 836
rect 1873 833 1887 836
rect 1916 827 1923 1133
rect 1936 1127 1943 1293
rect 1933 1113 1947 1127
rect 1976 927 1983 1273
rect 2016 1264 2024 1376
rect 1995 1076 2003 1156
rect 1995 1038 2003 1062
rect 1936 867 1943 913
rect 1976 867 1983 913
rect 2036 887 2043 1653
rect 2056 1607 2063 1613
rect 2053 1593 2067 1607
rect 2115 1556 2123 1636
rect 2156 1567 2163 1753
rect 2196 1727 2203 1753
rect 2317 1744 2325 1824
rect 2373 1773 2387 1787
rect 2376 1767 2383 1773
rect 2396 1747 2403 1793
rect 2196 1607 2203 1713
rect 2216 1627 2223 1733
rect 2213 1613 2227 1627
rect 2193 1593 2207 1607
rect 2115 1518 2123 1542
rect 2256 1347 2263 1593
rect 2296 1587 2303 1613
rect 2293 1573 2307 1587
rect 2353 1573 2367 1587
rect 2396 1587 2403 1613
rect 2393 1573 2407 1587
rect 2316 1387 2323 1553
rect 2356 1447 2363 1573
rect 2296 1347 2303 1373
rect 2056 1107 2063 1313
rect 2133 1293 2147 1307
rect 2253 1333 2267 1347
rect 2293 1333 2307 1347
rect 2396 1323 2403 1433
rect 2436 1367 2443 1813
rect 2456 1744 2464 1856
rect 2453 1593 2467 1607
rect 2456 1347 2463 1593
rect 2477 1556 2485 1636
rect 2477 1518 2485 1542
rect 2496 1407 2503 1873
rect 2516 1787 2523 2013
rect 2556 2007 2563 2033
rect 2536 1643 2543 1813
rect 2556 1744 2564 1856
rect 2576 1727 2583 2093
rect 2616 2087 2623 2113
rect 2656 2087 2663 2173
rect 2676 2107 2683 2333
rect 2736 2307 2743 2313
rect 2733 2293 2747 2307
rect 2756 2187 2763 2396
rect 2613 2073 2627 2087
rect 2596 2067 2603 2073
rect 2593 2053 2607 2067
rect 2633 2053 2647 2067
rect 2653 2073 2667 2087
rect 2636 1987 2643 2053
rect 2676 2007 2683 2093
rect 2756 2087 2763 2093
rect 2733 2053 2747 2067
rect 2753 2073 2767 2087
rect 2736 2007 2743 2053
rect 2636 1767 2643 1773
rect 2516 1636 2543 1643
rect 2413 1323 2427 1327
rect 2333 1293 2347 1307
rect 2373 1303 2387 1307
rect 2396 1316 2427 1323
rect 2396 1303 2403 1316
rect 2136 1287 2143 1293
rect 2073 1273 2087 1287
rect 2076 1227 2083 1273
rect 2336 1167 2343 1293
rect 2373 1296 2403 1303
rect 2413 1313 2427 1316
rect 2373 1293 2387 1296
rect 2353 1273 2367 1287
rect 2433 1283 2447 1287
rect 2456 1283 2463 1293
rect 2433 1276 2463 1283
rect 2433 1273 2447 1276
rect 2473 1273 2487 1287
rect 2356 1187 2363 1273
rect 2093 1143 2107 1147
rect 2093 1136 2123 1143
rect 2093 1133 2107 1136
rect 2116 1127 2123 1136
rect 2156 1127 2163 1153
rect 2316 1147 2323 1153
rect 2153 1113 2167 1127
rect 1933 853 1947 867
rect 1953 833 1967 847
rect 1973 853 1987 867
rect 1876 667 1883 673
rect 1873 653 1887 667
rect 1853 643 1867 647
rect 1836 636 1867 643
rect 1896 647 1903 673
rect 1936 647 1943 733
rect 1956 723 1963 833
rect 1996 823 2003 853
rect 2013 823 2027 827
rect 1996 816 2027 823
rect 2013 813 2027 816
rect 2073 813 2087 827
rect 2133 833 2147 847
rect 2076 787 2083 813
rect 1956 716 1983 723
rect 1956 667 1963 693
rect 1976 667 1983 716
rect 1953 653 1967 667
rect 1853 633 1867 636
rect 1893 633 1907 647
rect 1933 633 1947 647
rect 1973 643 1987 647
rect 1996 643 2003 773
rect 2096 747 2103 793
rect 2136 787 2143 833
rect 2156 827 2163 893
rect 2176 867 2183 1133
rect 2313 1143 2327 1147
rect 2313 1136 2343 1143
rect 2313 1133 2327 1136
rect 2233 1123 2247 1127
rect 2233 1116 2263 1123
rect 2233 1113 2247 1116
rect 2256 1107 2263 1116
rect 2336 1123 2343 1136
rect 2353 1123 2367 1127
rect 2336 1116 2367 1123
rect 2353 1113 2367 1116
rect 2296 1087 2303 1093
rect 2377 1076 2385 1156
rect 2436 1127 2443 1253
rect 2476 1247 2483 1273
rect 2496 1227 2503 1293
rect 2516 1287 2523 1636
rect 2536 1607 2543 1613
rect 2533 1593 2547 1607
rect 2596 1547 2603 1673
rect 2616 1524 2624 1636
rect 2636 1627 2643 1753
rect 2577 1358 2585 1382
rect 2577 1264 2585 1344
rect 2433 1113 2447 1127
rect 2377 1038 2385 1062
rect 2173 813 2187 827
rect 2213 813 2227 827
rect 2256 823 2263 913
rect 2376 867 2383 913
rect 2416 867 2423 873
rect 2496 867 2503 1193
rect 2516 1044 2524 1156
rect 2556 943 2563 1173
rect 2576 1147 2583 1213
rect 2596 1187 2603 1513
rect 2633 1303 2647 1307
rect 2656 1303 2663 1613
rect 2676 1467 2683 1953
rect 2695 1838 2703 1862
rect 2695 1744 2703 1824
rect 2713 1783 2727 1787
rect 2713 1776 2743 1783
rect 2713 1773 2727 1776
rect 2736 1707 2743 1776
rect 2633 1296 2663 1303
rect 2696 1307 2703 1573
rect 2716 1524 2724 1636
rect 2756 1607 2763 2013
rect 2753 1593 2767 1607
rect 2776 1487 2783 2453
rect 2796 2347 2803 2513
rect 2816 2307 2823 2593
rect 2856 2567 2863 2613
rect 2896 2567 2903 2633
rect 2916 2583 2923 2713
rect 2936 2607 2943 2713
rect 2996 2707 3003 2753
rect 3016 2603 3023 2953
rect 3096 2807 3103 2973
rect 3116 2783 3123 2853
rect 3136 2807 3143 2833
rect 3156 2807 3163 2953
rect 3196 2927 3203 2996
rect 3196 2847 3203 2913
rect 3133 2783 3147 2787
rect 3033 2733 3047 2747
rect 3116 2776 3147 2783
rect 3096 2747 3103 2753
rect 3073 2733 3087 2747
rect 3036 2687 3043 2733
rect 3076 2723 3083 2733
rect 3116 2723 3123 2776
rect 3133 2773 3147 2776
rect 3056 2716 3083 2723
rect 3096 2716 3123 2723
rect 3056 2707 3063 2716
rect 2996 2596 3023 2603
rect 2916 2576 2943 2583
rect 2853 2553 2867 2567
rect 2873 2533 2887 2547
rect 2893 2553 2907 2567
rect 2876 2527 2883 2533
rect 2936 2523 2943 2576
rect 2953 2523 2967 2527
rect 2936 2516 2967 2523
rect 2953 2513 2967 2516
rect 2956 2447 2963 2513
rect 2836 2287 2843 2313
rect 2936 2287 2943 2313
rect 2813 2263 2827 2267
rect 2796 2256 2827 2263
rect 2833 2273 2847 2287
rect 2893 2273 2907 2287
rect 2796 1963 2803 2256
rect 2813 2253 2827 2256
rect 2896 2263 2903 2273
rect 2876 2256 2903 2263
rect 2816 2004 2824 2116
rect 2856 2103 2863 2253
rect 2876 2247 2883 2256
rect 2933 2273 2947 2287
rect 2953 2253 2967 2267
rect 2896 2207 2903 2233
rect 2836 2096 2863 2103
rect 2796 1956 2823 1963
rect 2796 1744 2804 1856
rect 2816 1783 2823 1956
rect 2836 1827 2843 2096
rect 2896 2087 2903 2193
rect 2893 2083 2907 2087
rect 2876 2076 2907 2083
rect 2833 1783 2847 1787
rect 2816 1776 2847 1783
rect 2833 1773 2847 1776
rect 2796 1607 2803 1633
rect 2793 1593 2807 1607
rect 2816 1507 2823 1713
rect 2856 1683 2863 1833
rect 2876 1823 2883 2076
rect 2893 2073 2907 2076
rect 2876 1816 2903 1823
rect 2896 1783 2903 1816
rect 2887 1776 2903 1783
rect 2836 1676 2863 1683
rect 2836 1527 2843 1676
rect 2876 1647 2883 1773
rect 2855 1556 2863 1636
rect 2896 1583 2903 1693
rect 2916 1623 2923 2173
rect 2936 1967 2943 2213
rect 2956 2207 2963 2253
rect 2976 2207 2983 2513
rect 2996 2507 3003 2596
rect 3016 2567 3023 2573
rect 3056 2567 3063 2613
rect 3076 2567 3083 2693
rect 3013 2553 3027 2567
rect 3053 2553 3067 2567
rect 3096 2563 3103 2716
rect 3136 2567 3143 2713
rect 3096 2556 3123 2563
rect 3076 2547 3083 2553
rect 3073 2533 3087 2547
rect 2955 2036 2963 2116
rect 2955 1998 2963 2022
rect 2996 1907 3003 2293
rect 3016 2224 3024 2336
rect 3016 2087 3023 2113
rect 3036 2043 3043 2493
rect 3076 2267 3083 2333
rect 3096 2307 3103 2533
rect 3116 2487 3123 2556
rect 3156 2547 3163 2733
rect 3176 2707 3183 2733
rect 3196 2587 3203 2793
rect 3153 2533 3167 2547
rect 3173 2513 3187 2527
rect 3176 2487 3183 2513
rect 3093 2253 3107 2267
rect 3096 2247 3103 2253
rect 3116 2227 3123 2433
rect 3176 2407 3183 2473
rect 3216 2467 3223 2913
rect 3236 2807 3243 3173
rect 3276 3147 3283 3253
rect 3396 3263 3403 3313
rect 3293 3243 3307 3247
rect 3376 3256 3403 3263
rect 3376 3247 3383 3256
rect 3293 3236 3323 3243
rect 3293 3233 3307 3236
rect 3256 2947 3263 3013
rect 3276 2767 3283 2893
rect 3296 2827 3303 3193
rect 3316 3127 3323 3236
rect 3336 3127 3343 3233
rect 3373 3233 3387 3247
rect 3393 3213 3407 3227
rect 3396 3183 3403 3213
rect 3416 3207 3423 3273
rect 3436 3267 3443 3353
rect 3456 3267 3463 3293
rect 3453 3253 3467 3267
rect 3433 3213 3447 3227
rect 3396 3176 3423 3183
rect 3316 3047 3323 3113
rect 3376 3047 3383 3153
rect 3416 3067 3423 3176
rect 3436 3127 3443 3213
rect 3476 3187 3483 3413
rect 3556 3407 3563 3493
rect 3613 3473 3627 3487
rect 3633 3493 3647 3507
rect 3653 3473 3667 3487
rect 3496 3267 3503 3313
rect 3516 3267 3523 3273
rect 3556 3267 3563 3293
rect 3513 3253 3527 3267
rect 3553 3253 3567 3267
rect 3576 3247 3583 3453
rect 3436 3047 3443 3073
rect 3313 3033 3327 3047
rect 3373 3043 3387 3047
rect 3373 3036 3403 3043
rect 3373 3033 3387 3036
rect 3353 2993 3367 3007
rect 3316 2887 3323 2993
rect 3356 2967 3363 2993
rect 3376 2867 3383 2993
rect 3396 2827 3403 3036
rect 3433 3033 3447 3047
rect 3456 3003 3463 3173
rect 3476 3047 3483 3073
rect 3473 3033 3487 3047
rect 3496 3007 3503 3213
rect 3536 3103 3543 3133
rect 3516 3096 3543 3103
rect 3516 3047 3523 3096
rect 3556 3047 3563 3053
rect 3576 3047 3583 3213
rect 3596 3147 3603 3413
rect 3616 3387 3623 3473
rect 3656 3427 3663 3473
rect 3616 3267 3623 3373
rect 3656 3347 3663 3393
rect 3636 3267 3643 3293
rect 3633 3253 3647 3267
rect 3656 3223 3663 3333
rect 3676 3267 3683 3653
rect 3716 3627 3723 3973
rect 3736 3927 3743 3973
rect 3756 3767 3763 4033
rect 3796 3987 3803 3993
rect 3793 3973 3807 3987
rect 3833 3983 3847 3987
rect 3833 3976 3863 3983
rect 3833 3973 3847 3976
rect 3816 3967 3823 3973
rect 3813 3953 3827 3967
rect 3796 3787 3803 3913
rect 3856 3907 3863 3976
rect 3913 3953 3927 3967
rect 3936 3963 3943 4233
rect 3996 4223 4003 4273
rect 4016 4247 4023 4433
rect 4096 4387 4103 4456
rect 4133 4453 4147 4467
rect 4156 4447 4163 4493
rect 4256 4487 4263 4516
rect 4396 4487 4403 4513
rect 4233 4453 4247 4467
rect 4253 4473 4267 4487
rect 4393 4473 4407 4487
rect 3996 4216 4023 4223
rect 4016 4207 4023 4216
rect 4013 4193 4027 4207
rect 4073 4173 4087 4187
rect 4076 4167 4083 4173
rect 4033 4153 4047 4167
rect 4036 4107 4043 4153
rect 4036 3987 4043 4033
rect 3953 3963 3967 3967
rect 3936 3956 3967 3963
rect 3993 3963 4007 3967
rect 4013 3963 4027 3967
rect 3953 3953 3967 3956
rect 3993 3956 4027 3963
rect 4033 3973 4047 3987
rect 3993 3953 4007 3956
rect 4013 3953 4027 3956
rect 4053 3953 4067 3967
rect 3916 3907 3923 3953
rect 3773 3733 3787 3747
rect 3776 3727 3783 3733
rect 3793 3713 3807 3727
rect 3756 3587 3763 3713
rect 3776 3707 3783 3713
rect 3796 3707 3803 3713
rect 3796 3687 3803 3693
rect 3816 3687 3823 3893
rect 3716 3507 3723 3553
rect 3693 3473 3707 3487
rect 3713 3493 3727 3507
rect 3636 3216 3663 3223
rect 3616 3107 3623 3213
rect 3513 3033 3527 3047
rect 3553 3043 3567 3047
rect 3536 3036 3567 3043
rect 3456 2996 3483 3003
rect 3436 2847 3443 2873
rect 3253 2733 3267 2747
rect 3273 2753 3287 2767
rect 3293 2733 3307 2747
rect 3256 2723 3263 2733
rect 3256 2716 3283 2723
rect 3256 2567 3263 2693
rect 3276 2687 3283 2716
rect 3296 2667 3303 2733
rect 3296 2607 3303 2653
rect 3253 2553 3267 2567
rect 3236 2447 3243 2513
rect 3155 2318 3163 2342
rect 3136 2227 3143 2293
rect 3155 2224 3163 2304
rect 3176 2267 3183 2293
rect 3196 2287 3203 2373
rect 3256 2307 3263 2433
rect 3276 2347 3283 2573
rect 3316 2567 3323 2813
rect 3396 2803 3403 2813
rect 3376 2796 3403 2803
rect 3376 2787 3383 2796
rect 3456 2787 3463 2833
rect 3373 2773 3387 2787
rect 3413 2773 3427 2787
rect 3393 2753 3407 2767
rect 3396 2687 3403 2753
rect 3296 2327 3303 2553
rect 3336 2547 3343 2633
rect 3333 2533 3347 2547
rect 3356 2527 3363 2613
rect 3416 2587 3423 2773
rect 3453 2773 3467 2787
rect 3476 2747 3483 2996
rect 3496 2947 3503 2993
rect 3516 2867 3523 2933
rect 3507 2816 3513 2823
rect 3393 2583 3407 2587
rect 3376 2576 3407 2583
rect 3376 2547 3383 2576
rect 3393 2573 3407 2576
rect 3373 2543 3387 2547
rect 3373 2536 3403 2543
rect 3373 2533 3387 2536
rect 3353 2513 3367 2527
rect 3396 2503 3403 2536
rect 3436 2527 3443 2733
rect 3496 2687 3503 2793
rect 3536 2787 3543 3036
rect 3553 3033 3567 3036
rect 3636 3007 3643 3216
rect 3673 3213 3687 3227
rect 3676 3207 3683 3213
rect 3696 3207 3703 3473
rect 3736 3407 3743 3473
rect 3756 3347 3763 3513
rect 3776 3403 3783 3653
rect 3796 3527 3803 3673
rect 3816 3647 3823 3653
rect 3856 3627 3863 3673
rect 3916 3663 3923 3673
rect 3956 3667 3963 3933
rect 4016 3887 4023 3953
rect 4056 3907 4063 3953
rect 4076 3947 4083 4093
rect 4096 3827 4103 4353
rect 4116 4067 4123 4413
rect 4196 4287 4203 4453
rect 4236 4447 4243 4453
rect 4236 4427 4243 4433
rect 4136 4227 4143 4273
rect 4216 4247 4223 4393
rect 4276 4247 4283 4453
rect 4293 4433 4307 4447
rect 4513 4503 4527 4507
rect 4513 4496 4543 4503
rect 4513 4493 4527 4496
rect 4413 4453 4427 4467
rect 4536 4467 4543 4496
rect 4493 4453 4507 4467
rect 4533 4463 4547 4467
rect 4516 4456 4547 4463
rect 4416 4447 4423 4453
rect 4333 4433 4347 4447
rect 4296 4407 4303 4433
rect 4336 4407 4343 4433
rect 4133 4213 4147 4227
rect 4173 4213 4187 4227
rect 4153 4193 4167 4207
rect 4136 4047 4143 4173
rect 4156 4167 4163 4193
rect 4176 4167 4183 4213
rect 4213 4203 4227 4207
rect 4253 4203 4267 4207
rect 4207 4196 4227 4203
rect 4213 4193 4227 4196
rect 4236 4196 4267 4203
rect 4156 4127 4163 4153
rect 4136 4007 4143 4033
rect 4176 3987 4183 4013
rect 4136 3807 4143 3933
rect 3993 3713 4007 3727
rect 3896 3656 3923 3663
rect 3816 3507 3823 3613
rect 3856 3567 3863 3613
rect 3896 3547 3903 3656
rect 3893 3533 3907 3547
rect 3873 3523 3887 3527
rect 3856 3516 3887 3523
rect 3793 3473 3807 3487
rect 3813 3493 3827 3507
rect 3833 3483 3847 3487
rect 3856 3483 3863 3516
rect 3873 3513 3887 3516
rect 3956 3507 3963 3633
rect 3976 3583 3983 3713
rect 3996 3707 4003 3713
rect 4013 3693 4027 3707
rect 4053 3703 4067 3707
rect 4073 3703 4087 3707
rect 4053 3696 4087 3703
rect 4133 3713 4147 3727
rect 4053 3693 4067 3696
rect 4073 3693 4087 3696
rect 3996 3607 4003 3693
rect 4016 3667 4023 3693
rect 3976 3576 4003 3583
rect 3833 3476 3863 3483
rect 3833 3473 3847 3476
rect 3796 3427 3803 3473
rect 3776 3396 3803 3403
rect 3736 3247 3743 3273
rect 3776 3247 3783 3293
rect 3796 3267 3803 3396
rect 3856 3287 3863 3476
rect 3953 3493 3967 3507
rect 3973 3473 3987 3487
rect 3896 3267 3903 3333
rect 3833 3263 3847 3267
rect 3816 3256 3847 3263
rect 3816 3247 3823 3256
rect 3833 3253 3847 3256
rect 3713 3213 3727 3227
rect 3733 3233 3747 3247
rect 3916 3247 3923 3313
rect 3936 3267 3943 3473
rect 3976 3387 3983 3473
rect 3996 3407 4003 3576
rect 4036 3567 4043 3573
rect 4036 3507 4043 3553
rect 4056 3527 4063 3673
rect 4013 3473 4027 3487
rect 4033 3493 4047 3507
rect 4053 3473 4067 3487
rect 4016 3427 4023 3473
rect 4056 3387 4063 3473
rect 4076 3447 4083 3693
rect 4096 3527 4103 3613
rect 4136 3547 4143 3713
rect 4156 3687 4163 3833
rect 4176 3727 4183 3793
rect 4196 3727 4203 4173
rect 4236 4147 4243 4196
rect 4253 4193 4267 4196
rect 4216 3987 4223 4133
rect 4236 4007 4243 4053
rect 4256 4027 4263 4173
rect 4276 4167 4283 4173
rect 4276 4027 4283 4153
rect 4296 4107 4303 4253
rect 4396 4183 4403 4413
rect 4416 4267 4423 4433
rect 4456 4347 4463 4453
rect 4496 4427 4503 4453
rect 4516 4447 4523 4456
rect 4533 4453 4547 4456
rect 4556 4447 4563 4493
rect 4633 4463 4647 4467
rect 4593 4433 4607 4447
rect 4616 4456 4647 4463
rect 4413 4183 4427 4187
rect 4396 4176 4427 4183
rect 4413 4173 4427 4176
rect 4453 4173 4467 4187
rect 4333 4163 4347 4167
rect 4316 4156 4347 4163
rect 4316 4047 4323 4156
rect 4333 4153 4347 4156
rect 4336 4007 4343 4093
rect 4233 3993 4247 4007
rect 4213 3973 4227 3987
rect 4333 3993 4347 4007
rect 4356 3987 4363 4113
rect 4433 4023 4447 4027
rect 4456 4023 4463 4173
rect 4496 4107 4503 4333
rect 4536 4227 4543 4413
rect 4596 4387 4603 4433
rect 4596 4227 4603 4373
rect 4536 4207 4543 4213
rect 4553 4173 4567 4187
rect 4593 4173 4607 4187
rect 4433 4016 4463 4023
rect 4433 4013 4447 4016
rect 4353 3973 4367 3987
rect 4316 3963 4323 3973
rect 4316 3956 4343 3963
rect 4216 3727 4223 3933
rect 4256 3707 4263 3953
rect 4316 3727 4323 3733
rect 4336 3727 4343 3956
rect 4396 3867 4403 4013
rect 4456 4007 4463 4016
rect 4473 3953 4487 3967
rect 4516 3967 4523 4133
rect 4536 3987 4543 4153
rect 4556 4127 4563 4173
rect 4596 4167 4603 4173
rect 4616 4107 4623 4456
rect 4633 4453 4647 4456
rect 4693 4433 4707 4447
rect 4696 4227 4703 4433
rect 4716 4367 4723 4453
rect 4636 4147 4643 4193
rect 4653 4173 4667 4187
rect 4656 4127 4663 4173
rect 4693 4173 4707 4187
rect 4673 4153 4687 4167
rect 4436 3747 4443 3853
rect 4233 3693 4247 3707
rect 4236 3687 4243 3693
rect 4193 3673 4207 3687
rect 4136 3527 4143 3533
rect 4093 3513 4107 3527
rect 4113 3493 4127 3507
rect 4133 3513 4147 3527
rect 4156 3507 4163 3553
rect 4153 3493 4167 3507
rect 4116 3483 4123 3493
rect 4096 3476 4123 3483
rect 3987 3276 3993 3283
rect 4036 3267 4043 3293
rect 4056 3287 4063 3333
rect 3993 3263 4007 3267
rect 3793 3213 3807 3227
rect 3716 3207 3723 3213
rect 3796 3207 3803 3213
rect 3816 3167 3823 3233
rect 3893 3213 3907 3227
rect 3913 3233 3927 3247
rect 3976 3256 4007 3263
rect 4033 3263 4047 3267
rect 3976 3227 3983 3256
rect 3993 3253 4007 3256
rect 4033 3256 4053 3263
rect 4033 3253 4047 3256
rect 3656 3047 3663 3113
rect 3696 3047 3703 3093
rect 3653 3033 3667 3047
rect 3693 3033 3707 3047
rect 3716 3027 3723 3133
rect 3713 3023 3727 3027
rect 3713 3016 3743 3023
rect 3713 3013 3727 3016
rect 3613 2993 3627 3007
rect 3616 2967 3623 2993
rect 3556 2827 3563 2893
rect 3556 2767 3563 2813
rect 3513 2753 3527 2767
rect 3516 2747 3523 2753
rect 3533 2733 3547 2747
rect 3553 2753 3567 2767
rect 3573 2743 3587 2747
rect 3593 2743 3607 2747
rect 3573 2736 3607 2743
rect 3573 2733 3587 2736
rect 3593 2733 3607 2736
rect 3633 2733 3647 2747
rect 3676 2743 3683 2993
rect 3716 2807 3723 2953
rect 3736 2847 3743 3016
rect 3756 2987 3763 3113
rect 3776 3047 3783 3153
rect 3836 3107 3843 3213
rect 3876 3087 3883 3213
rect 3896 3187 3903 3213
rect 3816 3047 3823 3053
rect 3896 3047 3903 3173
rect 3773 3033 3787 3047
rect 3813 3033 3827 3047
rect 3796 2947 3803 3033
rect 3853 3013 3867 3027
rect 3936 3027 3943 3033
rect 3956 3027 3963 3213
rect 3976 3207 3983 3213
rect 4056 3203 4063 3253
rect 4076 3223 4083 3413
rect 4096 3347 4103 3476
rect 4116 3323 4123 3453
rect 4136 3347 4143 3473
rect 4176 3467 4183 3673
rect 4196 3647 4203 3673
rect 4116 3316 4143 3323
rect 4093 3223 4107 3227
rect 4076 3216 4107 3223
rect 4093 3213 4107 3216
rect 4056 3196 4083 3203
rect 4016 3047 4023 3193
rect 4036 3047 4043 3053
rect 4033 3033 4047 3047
rect 3893 3023 3907 3027
rect 3893 3016 3923 3023
rect 3893 3013 3907 3016
rect 3856 3003 3863 3013
rect 3836 2996 3863 3003
rect 3816 2967 3823 2993
rect 3756 2807 3763 2893
rect 3713 2783 3727 2787
rect 3696 2776 3727 2783
rect 3696 2767 3703 2776
rect 3713 2773 3727 2776
rect 3733 2753 3747 2767
rect 3656 2736 3683 2743
rect 3536 2667 3543 2733
rect 3476 2547 3483 2633
rect 3576 2607 3583 2733
rect 3616 2663 3623 2713
rect 3636 2687 3643 2733
rect 3616 2656 3643 2663
rect 3453 2513 3467 2527
rect 3473 2533 3487 2547
rect 3493 2513 3507 2527
rect 3376 2496 3403 2503
rect 3173 2253 3187 2267
rect 3253 2263 3267 2267
rect 3253 2256 3273 2263
rect 3253 2253 3267 2256
rect 3136 2143 3143 2213
rect 3116 2136 3143 2143
rect 3073 2083 3087 2087
rect 3073 2076 3103 2083
rect 3073 2073 3087 2076
rect 3053 2043 3067 2047
rect 3036 2036 3067 2043
rect 3053 2033 3067 2036
rect 3016 1887 3023 2033
rect 2935 1838 2943 1862
rect 2935 1744 2943 1824
rect 3016 1823 3023 1873
rect 3056 1867 3063 2033
rect 3096 2027 3103 2076
rect 3116 2047 3123 2136
rect 3196 2123 3203 2233
rect 3176 2116 3203 2123
rect 3176 2107 3183 2116
rect 3276 2103 3283 2233
rect 3296 2127 3303 2313
rect 3316 2307 3323 2333
rect 3356 2307 3363 2353
rect 3313 2293 3327 2307
rect 3353 2293 3367 2307
rect 3376 2287 3383 2496
rect 3456 2407 3463 2513
rect 3396 2307 3403 2353
rect 3496 2307 3503 2513
rect 3516 2487 3523 2573
rect 3596 2567 3603 2593
rect 3616 2587 3623 2613
rect 3636 2567 3643 2656
rect 3593 2553 3607 2567
rect 3616 2527 3623 2553
rect 3573 2513 3587 2527
rect 3536 2427 3543 2513
rect 3576 2507 3583 2513
rect 3536 2307 3543 2413
rect 3393 2293 3407 2307
rect 3456 2207 3463 2293
rect 3513 2273 3527 2287
rect 3533 2293 3547 2307
rect 3596 2287 3603 2493
rect 3336 2147 3343 2193
rect 3276 2096 3303 2103
rect 3196 2087 3203 2093
rect 3296 2087 3303 2096
rect 3376 2087 3383 2193
rect 3136 2067 3143 2073
rect 3133 2053 3147 2067
rect 3173 2053 3187 2067
rect 3193 2073 3207 2087
rect 3233 2063 3247 2067
rect 3216 2056 3247 2063
rect 3176 2047 3183 2053
rect 3216 2027 3223 2056
rect 3233 2053 3247 2056
rect 3273 2053 3287 2067
rect 3293 2073 3307 2087
rect 3276 2043 3283 2053
rect 3256 2036 3283 2043
rect 3116 1987 3123 2013
rect 2996 1816 3023 1823
rect 2996 1783 3003 1816
rect 3036 1807 3043 1813
rect 3013 1783 3027 1787
rect 2996 1776 3027 1783
rect 3033 1793 3047 1807
rect 3013 1773 3027 1776
rect 2916 1616 2943 1623
rect 2936 1607 2943 1616
rect 2913 1583 2927 1587
rect 2896 1576 2927 1583
rect 2913 1573 2927 1576
rect 2916 1567 2923 1573
rect 2855 1518 2863 1542
rect 2896 1487 2903 1533
rect 2633 1293 2647 1296
rect 2673 1293 2687 1307
rect 2636 1267 2643 1293
rect 2573 1133 2587 1147
rect 2616 1123 2623 1153
rect 2676 1127 2683 1293
rect 2716 1264 2724 1376
rect 2756 1187 2763 1353
rect 2813 1303 2827 1307
rect 2836 1303 2843 1353
rect 2813 1296 2843 1303
rect 2813 1293 2827 1296
rect 2793 1273 2807 1287
rect 2856 1283 2863 1473
rect 2896 1327 2903 1473
rect 2936 1327 2943 1353
rect 2956 1347 2963 1633
rect 3013 1553 3027 1567
rect 3016 1547 3023 1553
rect 2996 1427 3003 1533
rect 3016 1527 3023 1533
rect 3016 1343 3023 1453
rect 3036 1387 3043 1573
rect 3056 1527 3063 1833
rect 3076 1827 3083 1953
rect 3156 1827 3163 1973
rect 3176 1827 3183 1953
rect 3073 1813 3087 1827
rect 3127 1816 3143 1823
rect 3076 1687 3083 1773
rect 3096 1767 3103 1793
rect 3096 1587 3103 1633
rect 3136 1627 3143 1816
rect 3176 1807 3183 1813
rect 3196 1807 3203 1893
rect 3216 1807 3223 1813
rect 3236 1807 3243 1833
rect 3256 1827 3263 2036
rect 3313 2033 3327 2047
rect 3296 1967 3303 2033
rect 3316 2027 3323 2033
rect 3173 1793 3187 1807
rect 3193 1793 3207 1807
rect 3233 1793 3247 1807
rect 3156 1727 3163 1773
rect 3253 1773 3267 1787
rect 3213 1753 3227 1767
rect 3216 1747 3223 1753
rect 3236 1687 3243 1753
rect 3256 1667 3263 1773
rect 3073 1553 3087 1567
rect 3093 1573 3107 1587
rect 3153 1573 3167 1587
rect 3196 1587 3203 1633
rect 3193 1573 3207 1587
rect 3076 1467 3083 1553
rect 2873 1293 2887 1307
rect 2893 1313 2907 1327
rect 2913 1293 2927 1307
rect 2933 1313 2947 1327
rect 2996 1336 3023 1343
rect 2953 1293 2967 1307
rect 2876 1287 2883 1293
rect 2836 1276 2863 1283
rect 2796 1147 2803 1273
rect 2816 1127 2823 1153
rect 2633 1123 2647 1127
rect 2593 1103 2607 1107
rect 2616 1116 2647 1123
rect 2616 1103 2623 1116
rect 2593 1096 2623 1103
rect 2633 1113 2647 1116
rect 2593 1093 2607 1096
rect 2673 1113 2687 1127
rect 2733 1123 2747 1127
rect 2716 1116 2747 1123
rect 2696 1107 2703 1113
rect 2693 1093 2707 1107
rect 2556 936 2583 943
rect 2557 878 2565 902
rect 2373 853 2387 867
rect 2273 823 2287 827
rect 2256 816 2287 823
rect 2273 813 2287 816
rect 2313 813 2327 827
rect 1916 607 1923 633
rect 1973 636 2003 643
rect 2033 663 2047 667
rect 2056 663 2063 713
rect 2076 667 2083 673
rect 2033 656 2063 663
rect 2033 653 2047 656
rect 1973 633 1987 636
rect 1996 623 2003 636
rect 2056 647 2063 656
rect 2073 653 2087 667
rect 2013 623 2027 627
rect 1996 616 2027 623
rect 2096 647 2103 673
rect 2093 633 2107 647
rect 2013 613 2027 616
rect 1756 376 1783 383
rect 1733 343 1747 347
rect 1756 343 1763 376
rect 1733 336 1763 343
rect 1733 333 1747 336
rect 1756 327 1763 336
rect 1496 187 1503 193
rect 1333 153 1347 167
rect 1253 143 1267 147
rect 1313 143 1327 147
rect 1236 136 1267 143
rect 1253 133 1267 136
rect 1296 136 1327 143
rect 1156 127 1163 133
rect 1296 107 1303 136
rect 1313 133 1327 136
rect 1353 133 1367 147
rect 1373 153 1387 167
rect 1356 127 1363 133
rect 1396 127 1403 173
rect 1493 173 1507 187
rect 1516 167 1523 213
rect 1473 133 1487 147
rect 1513 153 1527 167
rect 1556 167 1563 193
rect 1616 167 1623 273
rect 1656 187 1663 193
rect 1653 173 1667 187
rect 1553 153 1567 167
rect 1613 153 1627 167
rect 1696 167 1703 233
rect 1476 107 1483 133
rect 1676 127 1683 133
rect 1736 84 1744 196
rect 1756 167 1763 313
rect 1816 304 1824 416
rect 1916 403 1923 593
rect 1916 396 1943 403
rect 1936 387 1943 396
rect 1913 353 1927 367
rect 1956 363 1963 613
rect 1973 363 1987 367
rect 1956 356 1987 363
rect 1973 353 1987 356
rect 1773 163 1787 167
rect 1773 156 1803 163
rect 1773 153 1787 156
rect 1796 127 1803 156
rect 1875 116 1883 196
rect 1916 107 1923 353
rect 2033 343 2047 347
rect 2056 343 2063 373
rect 2033 336 2063 343
rect 2033 333 2047 336
rect 2036 203 2043 333
rect 2096 304 2104 416
rect 2136 387 2143 753
rect 2176 727 2183 813
rect 2216 787 2223 813
rect 2236 687 2243 813
rect 2316 787 2323 813
rect 2177 596 2185 676
rect 2276 647 2283 773
rect 2233 643 2247 647
rect 2216 636 2247 643
rect 2177 558 2185 582
rect 2173 333 2187 347
rect 2176 327 2183 333
rect 2216 327 2223 636
rect 2233 633 2247 636
rect 2273 633 2287 647
rect 2316 564 2324 676
rect 2356 447 2363 853
rect 2413 853 2427 867
rect 2473 843 2487 847
rect 2456 836 2487 843
rect 2376 667 2383 733
rect 2376 647 2383 653
rect 2416 647 2423 773
rect 2456 667 2463 836
rect 2473 833 2487 836
rect 2533 823 2547 827
rect 2493 803 2507 807
rect 2516 816 2547 823
rect 2516 803 2523 816
rect 2493 796 2523 803
rect 2533 813 2547 816
rect 2493 793 2507 796
rect 2496 687 2503 793
rect 2557 784 2565 864
rect 2576 707 2583 936
rect 2656 927 2663 1093
rect 2716 1087 2723 1116
rect 2733 1113 2747 1116
rect 2793 1093 2807 1107
rect 2813 1113 2827 1127
rect 2727 1056 2743 1063
rect 2613 823 2627 827
rect 2596 816 2627 823
rect 2373 633 2387 647
rect 2393 613 2407 627
rect 2413 633 2427 647
rect 2453 643 2467 647
rect 2453 636 2483 643
rect 2453 633 2467 636
rect 2476 627 2483 636
rect 2235 398 2243 422
rect 2396 407 2403 613
rect 2536 467 2543 693
rect 2556 647 2563 673
rect 2553 633 2567 647
rect 2596 623 2603 816
rect 2613 813 2627 816
rect 2653 813 2667 827
rect 2656 787 2663 813
rect 2696 784 2704 896
rect 2716 787 2723 873
rect 2656 687 2663 693
rect 2656 667 2663 673
rect 2736 667 2743 1056
rect 2756 843 2763 1093
rect 2776 887 2783 1073
rect 2796 867 2803 1093
rect 2836 1007 2843 1276
rect 2916 1267 2923 1293
rect 2876 1147 2883 1153
rect 2873 1133 2887 1147
rect 2896 1127 2903 1173
rect 2816 847 2823 853
rect 2876 847 2883 1093
rect 2916 1067 2923 1113
rect 2936 1083 2943 1133
rect 2956 1127 2963 1293
rect 2976 1147 2983 1313
rect 2996 1207 3003 1336
rect 3036 1327 3043 1353
rect 3013 1293 3027 1307
rect 3033 1313 3047 1327
rect 3073 1313 3087 1327
rect 3053 1293 3067 1307
rect 3016 1287 3023 1293
rect 3056 1187 3063 1293
rect 3076 1287 3083 1313
rect 2976 1107 2983 1113
rect 2953 1083 2967 1087
rect 2936 1076 2967 1083
rect 3036 1107 3043 1133
rect 3076 1127 3083 1153
rect 3073 1113 3087 1127
rect 2953 1073 2967 1076
rect 2993 1073 3007 1087
rect 3053 1073 3067 1087
rect 2916 847 2923 933
rect 2936 847 2943 853
rect 2773 843 2787 847
rect 2756 836 2787 843
rect 2773 833 2787 836
rect 2813 833 2827 847
rect 2873 843 2887 847
rect 2833 813 2847 827
rect 2856 836 2887 843
rect 2836 807 2843 813
rect 2796 667 2803 753
rect 2653 653 2667 667
rect 2576 616 2603 623
rect 2516 387 2523 393
rect 2216 307 2223 313
rect 2235 304 2243 384
rect 2513 373 2527 387
rect 2253 343 2267 347
rect 2253 336 2283 343
rect 2253 333 2267 336
rect 2276 327 2283 336
rect 2393 343 2407 347
rect 2416 343 2423 353
rect 2393 336 2423 343
rect 2393 333 2407 336
rect 2416 327 2423 336
rect 2373 313 2387 327
rect 2433 313 2447 327
rect 2276 227 2283 233
rect 2016 196 2043 203
rect 2016 167 2023 196
rect 2116 187 2123 213
rect 2196 187 2203 193
rect 2113 173 2127 187
rect 1973 163 1987 167
rect 1936 156 1987 163
rect 1936 127 1943 156
rect 1973 153 1987 156
rect 1993 133 2007 147
rect 2013 153 2027 167
rect 2096 167 2103 173
rect 2053 133 2067 147
rect 2093 153 2107 167
rect 2193 173 2207 187
rect 2173 163 2187 167
rect 2156 156 2187 163
rect 2216 167 2223 173
rect 2236 167 2243 193
rect 2276 167 2283 213
rect 2296 187 2303 193
rect 2293 173 2307 187
rect 1996 127 2003 133
rect 2056 127 2063 133
rect 2156 127 2163 156
rect 2173 153 2187 156
rect 2213 153 2227 167
rect 2273 153 2287 167
rect 2316 167 2323 193
rect 2336 167 2343 313
rect 2376 227 2383 313
rect 2436 207 2443 313
rect 2576 307 2583 616
rect 2633 613 2647 627
rect 2673 623 2687 627
rect 2696 623 2703 653
rect 2716 647 2723 653
rect 2673 616 2703 623
rect 2713 633 2727 647
rect 2793 653 2807 667
rect 2673 613 2687 616
rect 2733 613 2747 627
rect 2636 427 2643 613
rect 2736 567 2743 613
rect 2756 467 2763 613
rect 2776 547 2783 613
rect 2836 587 2843 673
rect 2856 667 2863 836
rect 2873 833 2887 836
rect 2933 833 2947 847
rect 2956 843 2963 1073
rect 2996 1047 3003 1073
rect 3016 887 3023 1073
rect 3056 1067 3063 1073
rect 3096 1027 3103 1513
rect 3156 1507 3163 1573
rect 3136 1327 3143 1373
rect 3173 1323 3187 1327
rect 3196 1323 3203 1413
rect 3216 1343 3223 1653
rect 3256 1587 3263 1633
rect 3276 1607 3283 1853
rect 3356 1847 3363 2013
rect 3376 1987 3383 2053
rect 3396 2007 3403 2093
rect 3416 2087 3423 2113
rect 3476 2107 3483 2193
rect 3516 2143 3523 2273
rect 3573 2253 3587 2267
rect 3593 2273 3607 2287
rect 3576 2247 3583 2253
rect 3496 2136 3523 2143
rect 3496 2107 3503 2136
rect 3476 2087 3483 2093
rect 3453 2053 3467 2067
rect 3473 2073 3487 2087
rect 3496 2067 3503 2093
rect 3493 2053 3507 2067
rect 3333 1783 3347 1787
rect 3333 1776 3363 1783
rect 3333 1773 3347 1776
rect 3313 1753 3327 1767
rect 3316 1667 3323 1753
rect 3253 1573 3267 1587
rect 3276 1547 3283 1553
rect 3256 1347 3263 1453
rect 3276 1347 3283 1473
rect 3296 1447 3303 1633
rect 3316 1627 3323 1633
rect 3216 1336 3243 1343
rect 3173 1316 3203 1323
rect 3173 1313 3187 1316
rect 3153 1293 3167 1307
rect 3116 1127 3123 1293
rect 3156 1287 3163 1293
rect 3156 1147 3163 1273
rect 3216 1167 3223 1293
rect 3176 1127 3183 1153
rect 3236 1143 3243 1336
rect 3253 1333 3267 1347
rect 3296 1307 3303 1433
rect 3316 1387 3323 1593
rect 3356 1587 3363 1776
rect 3376 1627 3383 1833
rect 3436 1787 3443 2033
rect 3456 2027 3463 2053
rect 3516 2047 3523 2073
rect 3536 2067 3543 2113
rect 3556 2087 3563 2233
rect 3596 2167 3603 2233
rect 3533 2053 3547 2067
rect 3513 2033 3527 2047
rect 3553 2043 3567 2047
rect 3576 2043 3583 2113
rect 3616 2107 3623 2393
rect 3656 2347 3663 2736
rect 3676 2627 3683 2713
rect 3696 2707 3703 2753
rect 3716 2683 3723 2733
rect 3696 2676 3723 2683
rect 3676 2567 3683 2573
rect 3673 2553 3687 2567
rect 3656 2287 3663 2313
rect 3653 2273 3667 2287
rect 3636 2207 3643 2253
rect 3656 2067 3663 2073
rect 3676 2067 3683 2333
rect 3696 2307 3703 2676
rect 3716 2587 3723 2653
rect 3736 2627 3743 2753
rect 3756 2587 3763 2713
rect 3733 2533 3747 2547
rect 3716 2287 3723 2533
rect 3736 2487 3743 2533
rect 3736 2443 3743 2473
rect 3756 2467 3763 2553
rect 3736 2436 3763 2443
rect 3756 2287 3763 2436
rect 3776 2307 3783 2833
rect 3796 2803 3803 2933
rect 3836 2827 3843 2996
rect 3796 2796 3823 2803
rect 3816 2787 3823 2796
rect 3836 2767 3843 2813
rect 3876 2807 3883 2993
rect 3916 2987 3923 3016
rect 3933 3013 3947 3027
rect 3916 2807 3923 2953
rect 3936 2787 3943 2933
rect 3956 2827 3963 2873
rect 3796 2607 3803 2753
rect 3813 2733 3827 2747
rect 3833 2753 3847 2767
rect 3873 2753 3887 2767
rect 3913 2753 3927 2767
rect 3933 2773 3947 2787
rect 3816 2687 3823 2733
rect 3796 2567 3803 2573
rect 3793 2553 3807 2567
rect 3813 2513 3827 2527
rect 3796 2327 3803 2513
rect 3816 2507 3823 2513
rect 3733 2253 3747 2267
rect 3753 2273 3767 2287
rect 3793 2283 3807 2287
rect 3816 2283 3823 2353
rect 3793 2276 3823 2283
rect 3793 2273 3807 2276
rect 3773 2253 3787 2267
rect 3836 2263 3843 2713
rect 3876 2707 3883 2753
rect 3896 2727 3903 2753
rect 3876 2647 3883 2693
rect 3916 2687 3923 2753
rect 3936 2687 3943 2733
rect 3956 2683 3963 2773
rect 3976 2767 3983 2953
rect 3996 2767 4003 2973
rect 3993 2753 4007 2767
rect 3973 2713 3987 2727
rect 3976 2707 3983 2713
rect 3956 2676 3983 2683
rect 3976 2587 3983 2676
rect 3853 2563 3867 2567
rect 3893 2563 3907 2567
rect 3853 2556 3907 2563
rect 3853 2553 3867 2556
rect 3876 2527 3883 2556
rect 3893 2553 3907 2556
rect 3973 2563 3987 2567
rect 3996 2563 4003 2713
rect 4016 2627 4023 3013
rect 4036 2787 4043 2973
rect 4056 2967 4063 3173
rect 4076 3047 4083 3196
rect 4073 3033 4087 3047
rect 4096 2947 4103 3173
rect 4116 2787 4123 3213
rect 4136 3187 4143 3316
rect 4156 3267 4163 3433
rect 4196 3307 4203 3533
rect 4216 3527 4223 3613
rect 4236 3507 4243 3593
rect 4256 3507 4263 3633
rect 4276 3527 4283 3713
rect 4313 3713 4327 3727
rect 4373 3713 4387 3727
rect 4376 3687 4383 3713
rect 4376 3567 4383 3673
rect 4396 3547 4403 3733
rect 4433 3733 4447 3747
rect 4416 3667 4423 3713
rect 4416 3547 4423 3653
rect 4456 3647 4463 3913
rect 4476 3907 4483 3953
rect 4556 3947 4563 4093
rect 4676 4087 4683 4153
rect 4696 4023 4703 4173
rect 4696 4016 4723 4023
rect 4573 3953 4587 3967
rect 4616 3967 4623 4013
rect 4636 3987 4643 3993
rect 4716 4007 4723 4016
rect 4633 3973 4647 3987
rect 4713 3993 4727 4007
rect 4413 3533 4427 3547
rect 4296 3507 4303 3533
rect 4233 3493 4247 3507
rect 4293 3493 4307 3507
rect 4316 3487 4323 3513
rect 4313 3473 4327 3487
rect 4176 3267 4183 3273
rect 4216 3267 4223 3453
rect 4173 3253 4187 3267
rect 4193 3233 4207 3247
rect 4176 3147 4183 3213
rect 4196 3167 4203 3233
rect 4136 3047 4143 3113
rect 4133 3033 4147 3047
rect 4216 3047 4223 3053
rect 4236 3047 4243 3373
rect 4253 3213 4267 3227
rect 4256 3187 4263 3213
rect 4276 3127 4283 3393
rect 4296 3287 4303 3453
rect 4356 3447 4363 3453
rect 4153 3013 4167 3027
rect 4193 3023 4207 3027
rect 4176 3016 4207 3023
rect 4156 3007 4163 3013
rect 4156 2887 4163 2993
rect 4176 2967 4183 3016
rect 4193 3013 4207 3016
rect 4236 3007 4243 3013
rect 4273 3003 4287 3007
rect 4296 3003 4303 3213
rect 4316 3127 4323 3193
rect 4336 3187 4343 3273
rect 4356 3247 4363 3433
rect 4376 3427 4383 3513
rect 4456 3527 4463 3553
rect 4476 3527 4483 3813
rect 4536 3703 4543 3933
rect 4556 3747 4563 3913
rect 4576 3887 4583 3953
rect 4656 3827 4663 3973
rect 4553 3733 4567 3747
rect 4696 3747 4703 3953
rect 4573 3713 4587 3727
rect 4536 3696 4563 3703
rect 4513 3683 4527 3687
rect 4513 3676 4543 3683
rect 4513 3673 4527 3676
rect 4496 3567 4503 3633
rect 4433 3503 4447 3507
rect 4416 3496 4447 3503
rect 4453 3513 4467 3527
rect 4536 3507 4543 3676
rect 4556 3663 4563 3696
rect 4576 3687 4583 3713
rect 4556 3656 4583 3663
rect 4376 3407 4383 3413
rect 4396 3383 4403 3493
rect 4416 3467 4423 3496
rect 4433 3493 4447 3496
rect 4513 3493 4527 3507
rect 4376 3376 4403 3383
rect 4376 3247 4383 3376
rect 4396 3247 4403 3293
rect 4416 3267 4423 3353
rect 4436 3267 4443 3473
rect 4476 3287 4483 3493
rect 4496 3447 4503 3493
rect 4516 3467 4523 3493
rect 4393 3233 4407 3247
rect 4273 2996 4303 3003
rect 4273 2993 4287 2996
rect 4316 2987 4323 3113
rect 4336 3047 4343 3133
rect 4333 3033 4347 3047
rect 4353 3013 4367 3027
rect 4176 2907 4183 2953
rect 4216 2787 4223 2973
rect 4036 2667 4043 2753
rect 4053 2733 4067 2747
rect 4153 2753 4167 2767
rect 4213 2773 4227 2787
rect 4236 2767 4243 2873
rect 4276 2767 4283 2813
rect 4056 2727 4063 2733
rect 4036 2567 4043 2653
rect 4056 2567 4063 2633
rect 4076 2587 4083 2693
rect 3953 2533 3967 2547
rect 3973 2556 4003 2563
rect 3973 2553 3987 2556
rect 3876 2447 3883 2513
rect 3956 2507 3963 2533
rect 3996 2507 4003 2533
rect 4013 2513 4027 2527
rect 3816 2256 3843 2263
rect 3713 2233 3727 2247
rect 3716 2167 3723 2233
rect 3736 2187 3743 2253
rect 3776 2187 3783 2253
rect 3796 2087 3803 2253
rect 3816 2207 3823 2256
rect 3836 2227 3843 2233
rect 3613 2053 3627 2067
rect 3653 2053 3667 2067
rect 3553 2036 3583 2043
rect 3553 2033 3567 2036
rect 3476 1807 3483 1833
rect 3473 1793 3487 1807
rect 3493 1773 3507 1787
rect 3373 1553 3387 1567
rect 3316 1303 3323 1353
rect 3336 1347 3343 1533
rect 3376 1487 3383 1553
rect 3396 1547 3403 1713
rect 3456 1627 3463 1773
rect 3496 1687 3503 1773
rect 3516 1667 3523 1993
rect 3596 1827 3603 2053
rect 3616 2047 3623 2053
rect 3636 2027 3643 2053
rect 3636 1967 3643 1993
rect 3536 1787 3543 1813
rect 3616 1807 3623 1873
rect 3553 1773 3567 1787
rect 3593 1773 3607 1787
rect 3613 1793 3627 1807
rect 3556 1767 3563 1773
rect 3596 1703 3603 1773
rect 3596 1696 3623 1703
rect 3496 1643 3503 1653
rect 3496 1636 3523 1643
rect 3453 1573 3467 1587
rect 3496 1587 3503 1613
rect 3516 1587 3523 1636
rect 3536 1587 3543 1633
rect 3596 1587 3603 1673
rect 3616 1647 3623 1696
rect 3636 1687 3643 1733
rect 3656 1727 3663 2013
rect 3736 1987 3743 2053
rect 3753 2033 3767 2047
rect 3756 1987 3763 2033
rect 3796 2007 3803 2033
rect 3696 1867 3703 1873
rect 3696 1807 3703 1853
rect 3693 1793 3707 1807
rect 3616 1607 3623 1633
rect 3656 1607 3663 1673
rect 3676 1627 3683 1773
rect 3716 1767 3723 1853
rect 3733 1773 3747 1787
rect 3736 1747 3743 1773
rect 3773 1773 3787 1787
rect 3793 1783 3807 1787
rect 3816 1783 3823 2193
rect 3836 2087 3843 2213
rect 3833 2073 3847 2087
rect 3836 1907 3843 2033
rect 3856 1887 3863 2233
rect 3876 2087 3883 2293
rect 3916 2287 3923 2493
rect 3893 2253 3907 2267
rect 3933 2263 3947 2267
rect 3956 2263 3963 2273
rect 3933 2256 3963 2263
rect 3933 2253 3947 2256
rect 3973 2253 3987 2267
rect 3896 2207 3903 2253
rect 3896 2083 3903 2133
rect 3936 2107 3943 2253
rect 3976 2247 3983 2253
rect 3956 2087 3963 2193
rect 3913 2083 3927 2087
rect 3896 2076 3927 2083
rect 3793 1776 3823 1783
rect 3793 1773 3807 1776
rect 3753 1753 3767 1767
rect 3756 1747 3763 1753
rect 3696 1607 3703 1653
rect 3716 1627 3723 1633
rect 3713 1613 3727 1627
rect 3613 1593 3627 1607
rect 3493 1573 3507 1587
rect 3533 1573 3547 1587
rect 3356 1327 3363 1373
rect 3396 1363 3403 1513
rect 3456 1507 3463 1573
rect 3633 1573 3647 1587
rect 3653 1593 3667 1607
rect 3693 1593 3707 1607
rect 3553 1553 3567 1567
rect 3556 1527 3563 1553
rect 3376 1356 3403 1363
rect 3376 1347 3383 1356
rect 3413 1333 3427 1347
rect 3333 1303 3347 1307
rect 3316 1296 3347 1303
rect 3333 1293 3347 1296
rect 3276 1147 3283 1293
rect 3373 1293 3387 1307
rect 3376 1287 3383 1293
rect 3353 1273 3367 1287
rect 3236 1136 3263 1143
rect 3113 1113 3127 1127
rect 3136 1047 3143 1053
rect 2973 843 2987 847
rect 2956 836 2987 843
rect 2913 793 2927 807
rect 2916 787 2923 793
rect 2876 647 2883 773
rect 2956 767 2963 836
rect 2973 833 2987 836
rect 2936 647 2943 653
rect 2956 647 2963 733
rect 2996 727 3003 833
rect 2996 647 3003 673
rect 2873 623 2887 627
rect 2856 616 2887 623
rect 2856 607 2863 616
rect 2873 613 2887 616
rect 2933 633 2947 647
rect 2973 613 2987 627
rect 2993 633 3007 647
rect 3016 627 3023 793
rect 3036 743 3043 813
rect 3056 767 3063 913
rect 3036 736 3063 743
rect 3013 613 3027 627
rect 2916 603 2923 613
rect 2976 603 2983 613
rect 2916 596 2983 603
rect 2617 398 2625 422
rect 2636 407 2643 413
rect 2596 347 2603 373
rect 2593 333 2607 347
rect 2617 304 2625 384
rect 2673 333 2687 347
rect 2676 307 2683 333
rect 2356 187 2363 193
rect 2353 173 2367 187
rect 2313 153 2327 167
rect 2333 153 2347 167
rect 2376 167 2383 193
rect 2453 183 2467 187
rect 2453 176 2483 183
rect 2453 173 2467 176
rect 2416 143 2423 173
rect 2476 147 2483 176
rect 2433 143 2447 147
rect 2416 136 2447 143
rect 2433 133 2447 136
rect 2517 116 2525 196
rect 2576 167 2583 293
rect 2616 167 2623 193
rect 2573 153 2587 167
rect 2613 153 2627 167
rect 1875 78 1883 102
rect 2517 78 2525 102
rect 2656 84 2664 196
rect 2696 47 2703 453
rect 2756 304 2764 416
rect 2733 153 2747 167
rect 2736 147 2743 153
rect 2757 116 2765 196
rect 2757 78 2765 102
rect 2776 67 2783 433
rect 2856 403 2863 593
rect 2896 407 2903 593
rect 2856 396 2883 403
rect 2813 383 2827 387
rect 2796 376 2827 383
rect 2796 367 2803 376
rect 2813 373 2827 376
rect 2833 353 2847 367
rect 2836 347 2843 353
rect 2876 307 2883 396
rect 2916 367 2923 413
rect 3036 407 3043 713
rect 3056 647 3063 736
rect 3076 627 3083 633
rect 3053 593 3067 607
rect 3073 613 3087 627
rect 3093 603 3107 607
rect 3116 603 3123 853
rect 3136 747 3143 1033
rect 3156 867 3163 913
rect 3176 883 3183 1033
rect 3196 927 3203 1113
rect 3196 883 3203 893
rect 3176 876 3203 883
rect 3196 867 3203 876
rect 3153 853 3167 867
rect 3173 833 3187 847
rect 3193 853 3207 867
rect 3216 847 3223 913
rect 3176 827 3183 833
rect 3176 807 3183 813
rect 3233 813 3247 827
rect 3236 807 3243 813
rect 3213 793 3227 807
rect 3216 767 3223 793
rect 3176 667 3183 673
rect 3173 653 3187 667
rect 3153 613 3167 627
rect 3213 613 3227 627
rect 3093 596 3123 603
rect 3093 593 3107 596
rect 3056 587 3063 593
rect 2893 333 2907 347
rect 2913 353 2927 367
rect 2933 333 2947 347
rect 2973 333 2987 347
rect 2996 343 3003 393
rect 3013 343 3027 347
rect 2996 336 3027 343
rect 3013 333 3027 336
rect 2896 327 2903 333
rect 2816 167 2823 293
rect 2813 153 2827 167
rect 2876 147 2883 293
rect 2936 207 2943 333
rect 2976 287 2983 333
rect 2896 84 2904 196
rect 2956 167 2963 173
rect 3036 167 3043 193
rect 2953 153 2967 167
rect 3033 153 3047 167
rect 3056 127 3063 273
rect 3076 27 3083 393
rect 3116 383 3123 596
rect 3156 567 3163 613
rect 3176 487 3183 613
rect 3116 376 3143 383
rect 3136 327 3143 376
rect 3156 203 3163 393
rect 3176 387 3183 453
rect 3196 407 3203 613
rect 3216 607 3223 613
rect 3236 427 3243 713
rect 3173 373 3187 387
rect 3213 373 3227 387
rect 3193 353 3207 367
rect 3196 347 3203 353
rect 3216 287 3223 373
rect 3256 367 3263 1136
rect 3296 987 3303 1153
rect 3316 1047 3323 1273
rect 3356 1247 3363 1273
rect 3416 1247 3423 1333
rect 3433 1313 3447 1327
rect 3336 1127 3343 1153
rect 3373 1083 3387 1087
rect 3396 1083 3403 1173
rect 3436 1107 3443 1313
rect 3456 1247 3463 1293
rect 3476 1267 3483 1413
rect 3536 1347 3543 1373
rect 3496 1227 3503 1333
rect 3556 1327 3563 1433
rect 3576 1427 3583 1573
rect 3596 1563 3603 1573
rect 3636 1567 3643 1573
rect 3596 1556 3623 1563
rect 3596 1347 3603 1393
rect 3616 1367 3623 1556
rect 3616 1327 3623 1353
rect 3533 1293 3547 1307
rect 3553 1313 3567 1327
rect 3573 1293 3587 1307
rect 3613 1313 3627 1327
rect 3653 1313 3667 1327
rect 3536 1267 3543 1293
rect 3496 1107 3503 1153
rect 3536 1147 3543 1233
rect 3556 1123 3563 1193
rect 3576 1127 3583 1293
rect 3596 1287 3603 1293
rect 3636 1187 3643 1293
rect 3656 1267 3663 1313
rect 3676 1147 3683 1533
rect 3716 1527 3723 1573
rect 3756 1467 3763 1713
rect 3776 1667 3783 1773
rect 3776 1587 3783 1613
rect 3796 1587 3803 1733
rect 3816 1647 3823 1776
rect 3833 1783 3847 1787
rect 3856 1783 3863 1833
rect 3876 1827 3883 2033
rect 3833 1776 3863 1783
rect 3896 1787 3903 2076
rect 3913 2073 3927 2076
rect 3953 2073 3967 2087
rect 3996 2083 4003 2433
rect 4016 2307 4023 2513
rect 4056 2247 4063 2513
rect 4076 2487 4083 2573
rect 4116 2547 4123 2573
rect 4136 2567 4143 2733
rect 4156 2727 4163 2753
rect 4156 2587 4163 2613
rect 4176 2587 4183 2713
rect 4196 2647 4203 2753
rect 4253 2743 4267 2747
rect 4236 2736 4267 2743
rect 4273 2753 4287 2767
rect 4236 2687 4243 2736
rect 4253 2733 4267 2736
rect 4293 2733 4307 2747
rect 4156 2567 4163 2573
rect 4153 2553 4167 2567
rect 4093 2513 4107 2527
rect 4113 2533 4127 2547
rect 4173 2533 4187 2547
rect 4176 2523 4183 2533
rect 4156 2516 4183 2523
rect 4076 2367 4083 2473
rect 4076 2083 4083 2353
rect 4096 2347 4103 2513
rect 4136 2407 4143 2513
rect 4156 2467 4163 2516
rect 4156 2387 4163 2413
rect 4136 2287 4143 2333
rect 4156 2307 4163 2373
rect 4093 2273 4107 2287
rect 4096 2267 4103 2273
rect 4113 2253 4127 2267
rect 4176 2267 4183 2493
rect 4196 2407 4203 2513
rect 4236 2427 4243 2673
rect 4256 2627 4263 2713
rect 4296 2687 4303 2733
rect 4316 2527 4323 2733
rect 4336 2547 4343 2993
rect 4356 2967 4363 3013
rect 4376 2807 4383 3013
rect 4396 3007 4403 3013
rect 4416 2927 4423 3193
rect 4436 3147 4443 3233
rect 4453 3213 4467 3227
rect 4456 3187 4463 3213
rect 4496 3087 4503 3213
rect 4536 3167 4543 3493
rect 4556 3267 4563 3533
rect 4576 3527 4583 3656
rect 4596 3627 4603 3733
rect 4633 3713 4647 3727
rect 4673 3713 4687 3727
rect 4693 3733 4707 3747
rect 4596 3507 4603 3513
rect 4573 3473 4587 3487
rect 4593 3493 4607 3507
rect 4616 3487 4623 3573
rect 4636 3507 4643 3713
rect 4656 3547 4663 3713
rect 4676 3687 4683 3713
rect 4696 3627 4703 3693
rect 4656 3507 4663 3533
rect 4613 3473 4627 3487
rect 4653 3493 4667 3507
rect 4676 3487 4683 3573
rect 4716 3527 4723 3953
rect 4736 3847 4743 4393
rect 4756 3967 4763 4433
rect 4736 3707 4743 3813
rect 4696 3507 4703 3513
rect 4576 3447 4583 3473
rect 4673 3473 4687 3487
rect 4713 3473 4727 3487
rect 4596 3267 4603 3333
rect 4636 3247 4643 3413
rect 4656 3267 4663 3453
rect 4676 3267 4683 3433
rect 4696 3287 4703 3453
rect 4716 3447 4723 3473
rect 4736 3427 4743 3673
rect 4756 3647 4763 3933
rect 4776 3747 4783 4213
rect 4756 3447 4763 3613
rect 4736 3307 4743 3373
rect 4673 3253 4687 3267
rect 4593 3213 4607 3227
rect 4496 3027 4503 3053
rect 4433 2993 4447 3007
rect 4516 3023 4523 3133
rect 4556 3067 4563 3093
rect 4576 3067 4583 3173
rect 4553 3053 4567 3067
rect 4596 3043 4603 3213
rect 4616 3047 4623 3193
rect 4656 3187 4663 3253
rect 4693 3233 4707 3247
rect 4696 3227 4703 3233
rect 4656 3067 4663 3093
rect 4676 3047 4683 3073
rect 4696 3067 4703 3213
rect 4716 3047 4723 3233
rect 4736 3103 4743 3233
rect 4756 3127 4763 3393
rect 4776 3207 4783 3573
rect 4736 3096 4763 3103
rect 4576 3036 4603 3043
rect 4533 3023 4547 3027
rect 4516 3016 4547 3023
rect 4533 3013 4547 3016
rect 4436 2987 4443 2993
rect 4496 2787 4503 2973
rect 4516 2967 4523 2993
rect 4536 2963 4543 2993
rect 4556 2987 4563 3013
rect 4536 2956 4563 2963
rect 4393 2783 4407 2787
rect 4376 2776 4407 2783
rect 4353 2733 4367 2747
rect 4356 2727 4363 2733
rect 4376 2667 4383 2776
rect 4393 2773 4407 2776
rect 4516 2767 4523 2953
rect 4396 2627 4403 2713
rect 4436 2707 4443 2753
rect 4493 2733 4507 2747
rect 4293 2513 4307 2527
rect 4396 2527 4403 2553
rect 4416 2547 4423 2613
rect 4413 2533 4427 2547
rect 4296 2487 4303 2513
rect 4196 2307 4203 2373
rect 4256 2347 4263 2453
rect 4336 2347 4343 2513
rect 4193 2293 4207 2307
rect 4233 2293 4247 2307
rect 4236 2287 4243 2293
rect 4213 2273 4227 2287
rect 4253 2273 4267 2287
rect 4096 2247 4103 2253
rect 4116 2227 4123 2253
rect 4096 2107 4103 2213
rect 4156 2107 4163 2233
rect 3996 2076 4023 2083
rect 4076 2076 4103 2083
rect 3973 2063 3987 2067
rect 3973 2056 4003 2063
rect 3973 2053 3987 2056
rect 3916 1827 3923 2033
rect 3936 1967 3943 2053
rect 3996 2007 4003 2056
rect 3833 1773 3847 1776
rect 3873 1773 3887 1787
rect 3876 1767 3883 1773
rect 3896 1667 3903 1773
rect 3916 1727 3923 1773
rect 3956 1647 3963 1893
rect 3976 1787 3983 1993
rect 4016 1843 4023 2076
rect 4033 2033 4047 2047
rect 4073 2043 4087 2047
rect 4096 2043 4103 2076
rect 4136 2067 4143 2073
rect 4073 2036 4103 2043
rect 4073 2033 4087 2036
rect 4113 2033 4127 2047
rect 4133 2053 4147 2067
rect 4153 2033 4167 2047
rect 4036 2007 4043 2033
rect 4016 1836 4043 1843
rect 4036 1827 4043 1836
rect 4016 1807 4023 1813
rect 4056 1807 4063 1833
rect 4076 1827 4083 2033
rect 4116 2027 4123 2033
rect 4156 2027 4163 2033
rect 4116 1807 4123 2013
rect 4156 1867 4163 2013
rect 4156 1807 4163 1833
rect 4176 1823 4183 2233
rect 4196 2227 4203 2253
rect 4216 2187 4223 2273
rect 4236 2207 4243 2273
rect 4256 2267 4263 2273
rect 4256 2183 4263 2253
rect 4356 2247 4363 2413
rect 4376 2387 4383 2493
rect 4293 2233 4307 2247
rect 4296 2187 4303 2233
rect 4236 2176 4263 2183
rect 4216 2067 4223 2113
rect 4236 2087 4243 2176
rect 4256 2087 4263 2133
rect 4316 2087 4323 2233
rect 4376 2147 4383 2353
rect 4416 2327 4423 2493
rect 4436 2327 4443 2633
rect 4496 2567 4503 2733
rect 4536 2723 4543 2733
rect 4516 2716 4543 2723
rect 4516 2687 4523 2716
rect 4536 2587 4543 2673
rect 4556 2667 4563 2956
rect 4576 2787 4583 3036
rect 4613 3033 4627 3047
rect 4653 3043 4667 3047
rect 4673 3043 4687 3047
rect 4653 3036 4687 3043
rect 4653 3033 4667 3036
rect 4673 3033 4687 3036
rect 4713 3033 4727 3047
rect 4736 3027 4743 3053
rect 4733 3013 4747 3027
rect 4616 2847 4623 2993
rect 4516 2547 4523 2553
rect 4596 2567 4603 2693
rect 4453 2513 4467 2527
rect 4533 2533 4547 2547
rect 4573 2543 4587 2547
rect 4556 2536 4587 2543
rect 4593 2553 4607 2567
rect 4456 2447 4463 2513
rect 4536 2487 4543 2533
rect 4556 2507 4563 2536
rect 4573 2533 4587 2536
rect 4496 2307 4503 2473
rect 4556 2427 4563 2493
rect 4516 2307 4523 2393
rect 4453 2263 4467 2267
rect 4473 2263 4487 2267
rect 4453 2256 4487 2263
rect 4453 2253 4467 2256
rect 4473 2253 4487 2256
rect 4513 2253 4527 2267
rect 4373 2103 4387 2107
rect 4416 2103 4423 2253
rect 4373 2096 4423 2103
rect 4373 2093 4387 2096
rect 4253 2083 4267 2087
rect 4253 2076 4283 2083
rect 4253 2073 4267 2076
rect 4193 2033 4207 2047
rect 4213 2053 4227 2067
rect 4233 2033 4247 2047
rect 4196 2027 4203 2033
rect 4236 2007 4243 2033
rect 4276 2027 4283 2076
rect 4393 2053 4407 2067
rect 4293 2033 4307 2047
rect 4296 2007 4303 2033
rect 4216 1827 4223 1873
rect 4256 1827 4263 1833
rect 4176 1816 4203 1823
rect 3993 1773 4007 1787
rect 4013 1793 4027 1807
rect 4033 1773 4047 1787
rect 4053 1793 4067 1807
rect 4113 1793 4127 1807
rect 4133 1773 4147 1787
rect 4153 1793 4167 1807
rect 4196 1787 4203 1816
rect 4233 1793 4247 1807
rect 4253 1813 4267 1827
rect 4173 1773 4187 1787
rect 3996 1767 4003 1773
rect 3996 1707 4003 1753
rect 4016 1667 4023 1753
rect 4036 1727 4043 1773
rect 3816 1587 3823 1593
rect 3813 1573 3827 1587
rect 3796 1567 3803 1573
rect 3793 1553 3807 1567
rect 3833 1553 3847 1567
rect 3713 1343 3727 1347
rect 3696 1336 3727 1343
rect 3696 1307 3703 1336
rect 3713 1333 3727 1336
rect 3733 1313 3747 1327
rect 3736 1307 3743 1313
rect 3716 1227 3723 1293
rect 3776 1227 3783 1353
rect 3796 1347 3803 1393
rect 3836 1347 3843 1553
rect 3793 1333 3807 1347
rect 3813 1313 3827 1327
rect 3856 1343 3863 1633
rect 3913 1573 3927 1587
rect 3896 1367 3903 1573
rect 3916 1567 3923 1573
rect 3856 1336 3883 1343
rect 3816 1287 3823 1313
rect 3696 1147 3703 1213
rect 3536 1116 3563 1123
rect 3373 1076 3403 1083
rect 3373 1073 3387 1076
rect 3413 1073 3427 1087
rect 3433 1093 3447 1107
rect 3493 1093 3507 1107
rect 3513 1073 3527 1087
rect 3416 1067 3423 1073
rect 3516 1067 3523 1073
rect 3536 1067 3543 1116
rect 3576 1107 3583 1113
rect 3573 1093 3587 1107
rect 3593 1073 3607 1087
rect 3287 896 3293 903
rect 3316 883 3323 1033
rect 3296 876 3323 883
rect 3276 847 3283 873
rect 3273 833 3287 847
rect 3276 647 3283 753
rect 3296 667 3303 876
rect 3356 867 3363 873
rect 3333 833 3347 847
rect 3353 853 3367 867
rect 3336 823 3343 833
rect 3336 816 3363 823
rect 3327 796 3333 803
rect 3356 727 3363 816
rect 3376 767 3383 1013
rect 3433 863 3447 867
rect 3413 833 3427 847
rect 3433 856 3463 863
rect 3433 853 3447 856
rect 3416 827 3423 833
rect 3316 667 3323 693
rect 3293 623 3307 627
rect 3316 623 3323 653
rect 3336 627 3343 673
rect 3293 616 3323 623
rect 3293 613 3307 616
rect 3333 613 3347 627
rect 3356 607 3363 693
rect 3376 647 3383 713
rect 3396 687 3403 813
rect 3416 787 3423 813
rect 3456 787 3463 856
rect 3456 707 3463 773
rect 3373 633 3387 647
rect 3436 647 3443 673
rect 3476 667 3483 993
rect 3496 867 3503 1053
rect 3516 947 3523 1053
rect 3556 987 3563 1073
rect 3596 1067 3603 1073
rect 3616 927 3623 1133
rect 3653 1093 3667 1107
rect 3696 1107 3703 1133
rect 3693 1093 3707 1107
rect 3656 1047 3663 1093
rect 3556 867 3563 873
rect 3553 853 3567 867
rect 3573 833 3587 847
rect 3576 827 3583 833
rect 3513 793 3527 807
rect 3496 647 3503 793
rect 3516 747 3523 793
rect 3433 633 3447 647
rect 3493 623 3507 627
rect 3516 623 3523 693
rect 3556 667 3563 733
rect 3616 707 3623 873
rect 3636 747 3643 1013
rect 3716 947 3723 1113
rect 3776 1107 3783 1173
rect 3876 1147 3883 1336
rect 3913 1293 3927 1307
rect 3916 1187 3923 1293
rect 3853 1143 3867 1147
rect 3847 1136 3867 1143
rect 3853 1133 3867 1136
rect 3816 1107 3823 1133
rect 3893 1123 3907 1127
rect 3753 1073 3767 1087
rect 3813 1093 3827 1107
rect 3893 1116 3923 1123
rect 3893 1113 3907 1116
rect 3756 883 3763 1073
rect 3876 1067 3883 1093
rect 3656 867 3663 873
rect 3653 853 3667 867
rect 3693 853 3707 867
rect 3736 876 3763 883
rect 3673 833 3687 847
rect 3676 767 3683 833
rect 3676 667 3683 753
rect 3696 707 3703 853
rect 3713 833 3727 847
rect 3716 827 3723 833
rect 3696 667 3703 693
rect 3716 667 3723 813
rect 3553 653 3567 667
rect 3693 653 3707 667
rect 3493 616 3523 623
rect 3593 643 3607 647
rect 3653 643 3667 647
rect 3493 613 3507 616
rect 3533 613 3547 627
rect 3593 636 3623 643
rect 3593 633 3607 636
rect 3456 607 3463 613
rect 3276 407 3283 593
rect 3536 547 3543 613
rect 3356 387 3363 433
rect 3233 353 3247 367
rect 3293 353 3307 367
rect 3333 353 3347 367
rect 3236 307 3243 353
rect 3136 196 3183 203
rect 3136 167 3143 196
rect 3093 133 3107 147
rect 3133 153 3147 167
rect 3176 167 3183 196
rect 3216 167 3223 193
rect 3193 133 3207 147
rect 3213 153 3227 167
rect 3236 147 3243 293
rect 3296 187 3303 353
rect 3336 307 3343 353
rect 3353 333 3367 347
rect 3356 307 3363 333
rect 3316 187 3323 193
rect 3313 173 3327 187
rect 3233 133 3247 147
rect 3096 127 3103 133
rect 3196 107 3203 133
rect 3256 107 3263 173
rect 3276 127 3283 153
rect 3356 147 3363 193
rect 3396 147 3403 333
rect 3353 133 3367 147
rect 3373 113 3387 127
rect 3416 123 3423 173
rect 3436 167 3443 393
rect 3456 207 3463 533
rect 3556 467 3563 593
rect 3556 387 3563 393
rect 3533 353 3547 367
rect 3553 373 3567 387
rect 3536 287 3543 353
rect 3576 307 3583 613
rect 3616 407 3623 636
rect 3636 636 3667 643
rect 3636 607 3643 636
rect 3653 633 3667 636
rect 3716 547 3723 613
rect 3736 587 3743 876
rect 3773 833 3787 847
rect 3853 833 3867 847
rect 3776 807 3783 833
rect 3756 647 3763 793
rect 3796 667 3803 833
rect 3856 807 3863 833
rect 3816 667 3823 713
rect 3876 707 3883 813
rect 3896 647 3903 1073
rect 3916 887 3923 1116
rect 3936 1027 3943 1473
rect 3956 1143 3963 1613
rect 3976 1607 3983 1653
rect 4016 1607 4023 1613
rect 3973 1593 3987 1607
rect 4013 1593 4027 1607
rect 4036 1603 4043 1633
rect 4056 1627 4063 1733
rect 4076 1627 4083 1753
rect 4136 1723 4143 1773
rect 4136 1716 4163 1723
rect 4036 1596 4063 1603
rect 4016 1527 4023 1553
rect 3996 1347 4003 1393
rect 4016 1327 4023 1413
rect 4056 1347 4063 1596
rect 4076 1447 4083 1613
rect 4096 1607 4103 1653
rect 4116 1587 4123 1633
rect 4136 1607 4143 1693
rect 4156 1667 4163 1716
rect 4176 1707 4183 1773
rect 4196 1627 4203 1653
rect 4216 1627 4223 1753
rect 4236 1663 4243 1793
rect 4276 1767 4283 1793
rect 4293 1773 4307 1787
rect 4296 1707 4303 1773
rect 4316 1747 4323 1953
rect 4336 1867 4343 2053
rect 4376 1883 4383 2053
rect 4396 1907 4403 2053
rect 4436 2007 4443 2213
rect 4356 1876 4383 1883
rect 4336 1827 4343 1833
rect 4356 1827 4363 1876
rect 4333 1813 4347 1827
rect 4353 1773 4367 1787
rect 4356 1767 4363 1773
rect 4376 1767 4383 1853
rect 4456 1827 4463 2093
rect 4476 2087 4483 2253
rect 4496 2127 4503 2233
rect 4516 2207 4523 2253
rect 4536 2227 4543 2253
rect 4556 2187 4563 2333
rect 4576 2283 4583 2513
rect 4616 2367 4623 2773
rect 4676 2767 4683 2793
rect 4696 2787 4703 3013
rect 4673 2753 4687 2767
rect 4716 2727 4723 2813
rect 4653 2713 4667 2727
rect 4636 2467 4643 2713
rect 4656 2687 4663 2713
rect 4656 2567 4663 2653
rect 4716 2647 4723 2693
rect 4736 2687 4743 2793
rect 4756 2787 4763 3096
rect 4696 2527 4703 2613
rect 4713 2543 4727 2547
rect 4713 2536 4743 2543
rect 4713 2533 4727 2536
rect 4636 2287 4643 2313
rect 4656 2307 4663 2453
rect 4676 2387 4683 2493
rect 4676 2287 4683 2373
rect 4696 2287 4703 2473
rect 4716 2447 4723 2493
rect 4736 2407 4743 2536
rect 4716 2287 4723 2393
rect 4593 2283 4607 2287
rect 4576 2276 4607 2283
rect 4576 2143 4583 2276
rect 4593 2273 4607 2276
rect 4613 2253 4627 2267
rect 4633 2273 4647 2287
rect 4673 2273 4687 2287
rect 4713 2273 4727 2287
rect 4616 2187 4623 2253
rect 4656 2247 4663 2253
rect 4707 2236 4723 2243
rect 4556 2136 4583 2143
rect 4516 2107 4523 2113
rect 4513 2093 4527 2107
rect 4473 2073 4487 2087
rect 4556 2087 4563 2136
rect 4493 2053 4507 2067
rect 4533 2053 4547 2067
rect 4496 2047 4503 2053
rect 4496 1807 4503 2033
rect 4516 1867 4523 2053
rect 4536 2027 4543 2053
rect 4576 2047 4583 2113
rect 4596 2087 4603 2173
rect 4573 2033 4587 2047
rect 4536 1847 4543 2013
rect 4433 1773 4447 1787
rect 4236 1656 4263 1663
rect 4093 1553 4107 1567
rect 4113 1573 4127 1587
rect 4153 1573 4167 1587
rect 4236 1587 4243 1633
rect 4256 1607 4263 1656
rect 4253 1593 4267 1607
rect 4096 1547 4103 1553
rect 4116 1463 4123 1533
rect 4156 1527 4163 1573
rect 4096 1456 4123 1463
rect 4076 1327 4083 1373
rect 4096 1367 4103 1456
rect 3993 1293 4007 1307
rect 4073 1313 4087 1327
rect 3996 1247 4003 1293
rect 4053 1273 4067 1287
rect 4056 1267 4063 1273
rect 3973 1143 3987 1147
rect 3956 1136 3987 1143
rect 3973 1133 3987 1136
rect 3976 903 3983 1093
rect 3996 927 4003 1193
rect 4016 1127 4023 1213
rect 4096 1167 4103 1333
rect 4116 1307 4123 1433
rect 4156 1387 4163 1513
rect 4136 1347 4143 1373
rect 4176 1347 4183 1433
rect 4133 1333 4147 1347
rect 4153 1313 4167 1327
rect 4173 1333 4187 1347
rect 4136 1267 4143 1293
rect 4096 1143 4103 1153
rect 4136 1147 4143 1213
rect 4156 1207 4163 1313
rect 4176 1147 4183 1293
rect 4196 1227 4203 1453
rect 4216 1367 4223 1513
rect 4236 1427 4243 1573
rect 4276 1467 4283 1553
rect 4216 1347 4223 1353
rect 4213 1333 4227 1347
rect 4253 1343 4267 1347
rect 4276 1343 4283 1453
rect 4336 1407 4343 1673
rect 4356 1627 4363 1653
rect 4436 1647 4443 1773
rect 4353 1613 4367 1627
rect 4356 1387 4363 1453
rect 4316 1347 4323 1373
rect 4376 1367 4383 1553
rect 4396 1527 4403 1633
rect 4456 1607 4463 1633
rect 4453 1593 4467 1607
rect 4436 1547 4443 1573
rect 4233 1313 4247 1327
rect 4253 1336 4283 1343
rect 4253 1333 4267 1336
rect 4236 1243 4243 1313
rect 4256 1267 4263 1293
rect 4276 1247 4283 1313
rect 4356 1307 4363 1353
rect 4416 1327 4423 1373
rect 4456 1343 4463 1553
rect 4476 1367 4483 1733
rect 4516 1607 4523 1813
rect 4556 1807 4563 1873
rect 4576 1827 4583 1993
rect 4636 1887 4643 2113
rect 4656 2067 4663 2233
rect 4653 2053 4667 2067
rect 4676 2063 4683 2193
rect 4696 2087 4703 2173
rect 4716 2107 4723 2236
rect 4736 2183 4743 2233
rect 4756 2207 4763 2753
rect 4776 2707 4783 3073
rect 4776 2467 4783 2673
rect 4776 2287 4783 2313
rect 4736 2176 4763 2183
rect 4693 2063 4707 2067
rect 4676 2056 4707 2063
rect 4693 2053 4707 2056
rect 4713 2033 4727 2047
rect 4636 1847 4643 1873
rect 4696 1863 4703 2013
rect 4716 2007 4723 2033
rect 4676 1856 4703 1863
rect 4596 1816 4613 1823
rect 4596 1807 4603 1816
rect 4656 1807 4663 1853
rect 4676 1807 4683 1856
rect 4696 1807 4703 1833
rect 4573 1773 4587 1787
rect 4593 1793 4607 1807
rect 4693 1793 4707 1807
rect 4576 1767 4583 1773
rect 4616 1627 4623 1753
rect 4636 1627 4643 1773
rect 4656 1647 4663 1773
rect 4673 1753 4687 1767
rect 4676 1727 4683 1753
rect 4696 1727 4703 1753
rect 4656 1603 4663 1633
rect 4647 1596 4663 1603
rect 4493 1553 4507 1567
rect 4496 1547 4503 1553
rect 4496 1507 4503 1533
rect 4536 1347 4543 1533
rect 4456 1336 4483 1343
rect 4476 1327 4483 1336
rect 4373 1313 4387 1327
rect 4333 1293 4347 1307
rect 4336 1287 4343 1293
rect 4376 1287 4383 1313
rect 4393 1293 4407 1307
rect 4413 1313 4427 1327
rect 4453 1293 4467 1307
rect 4493 1293 4507 1307
rect 4313 1273 4327 1287
rect 4316 1267 4323 1273
rect 4216 1236 4243 1243
rect 4196 1147 4203 1153
rect 4216 1147 4223 1236
rect 4076 1136 4103 1143
rect 4013 1073 4027 1087
rect 4056 1087 4063 1133
rect 4076 1127 4083 1136
rect 4193 1133 4207 1147
rect 4076 1107 4083 1113
rect 4153 1123 4167 1127
rect 4073 1093 4087 1107
rect 4107 1096 4123 1103
rect 4016 907 4023 1073
rect 3976 896 3993 903
rect 4016 867 4023 893
rect 3933 863 3947 867
rect 3916 856 3947 863
rect 3916 687 3923 856
rect 3933 853 3947 856
rect 4036 847 4043 853
rect 4056 847 4063 893
rect 3993 833 4007 847
rect 4033 833 4047 847
rect 3996 827 4003 833
rect 3936 727 3943 773
rect 3753 633 3767 647
rect 3833 643 3847 647
rect 3813 613 3827 627
rect 3833 636 3863 643
rect 3833 633 3847 636
rect 3816 607 3823 613
rect 3636 407 3643 433
rect 3633 383 3647 387
rect 3613 353 3627 367
rect 3633 376 3663 383
rect 3633 373 3647 376
rect 3556 227 3563 293
rect 3596 247 3603 333
rect 3616 307 3623 353
rect 3656 347 3663 376
rect 3696 367 3703 393
rect 3673 333 3687 347
rect 3693 353 3707 367
rect 3733 353 3747 367
rect 3676 327 3683 333
rect 3656 307 3663 313
rect 3676 307 3683 313
rect 3553 183 3567 187
rect 3576 183 3583 233
rect 3736 207 3743 353
rect 3756 267 3763 593
rect 3856 567 3863 636
rect 3936 627 3943 653
rect 3933 613 3947 627
rect 3636 187 3643 193
rect 3756 187 3763 213
rect 3553 176 3583 183
rect 3553 173 3567 176
rect 3496 147 3503 173
rect 3633 173 3647 187
rect 3593 163 3607 167
rect 3433 123 3447 127
rect 3416 116 3447 123
rect 3493 133 3507 147
rect 3533 133 3547 147
rect 3576 156 3607 163
rect 3433 113 3447 116
rect 3536 127 3543 133
rect 3376 107 3383 113
rect 3576 107 3583 156
rect 3593 153 3607 156
rect 3613 133 3627 147
rect 3653 143 3667 147
rect 3676 143 3683 173
rect 3653 136 3683 143
rect 3753 173 3767 187
rect 3776 183 3783 473
rect 3793 333 3807 347
rect 3796 287 3803 333
rect 3833 333 3847 347
rect 3856 343 3863 413
rect 3873 343 3887 347
rect 3856 336 3887 343
rect 3873 333 3887 336
rect 3813 313 3827 327
rect 3816 247 3823 313
rect 3836 227 3843 333
rect 3876 327 3883 333
rect 3933 333 3947 347
rect 3936 327 3943 333
rect 3893 313 3907 327
rect 3896 227 3903 313
rect 3776 176 3803 183
rect 3653 133 3667 136
rect 3773 133 3787 147
rect 3616 87 3623 133
rect 3776 107 3783 133
rect 3496 -24 3503 13
rect 3576 -24 3583 33
rect 3616 -24 3623 53
rect 3796 27 3803 176
rect 3833 133 3847 147
rect 3876 147 3883 173
rect 3896 163 3903 213
rect 3956 183 3963 633
rect 3996 627 4003 673
rect 4016 667 4023 833
rect 4076 667 4083 913
rect 4096 887 4103 1073
rect 4116 1067 4123 1096
rect 4153 1116 4183 1123
rect 4153 1113 4167 1116
rect 4156 1027 4163 1073
rect 4116 867 4123 953
rect 4156 867 4163 933
rect 4176 907 4183 1116
rect 4213 1093 4227 1107
rect 4196 1007 4203 1093
rect 4216 927 4223 1093
rect 4236 1087 4243 1213
rect 4113 813 4127 827
rect 4176 843 4183 873
rect 4256 867 4263 1233
rect 4276 1127 4283 1193
rect 4316 1167 4323 1253
rect 4356 1167 4363 1173
rect 4273 1113 4287 1127
rect 4333 1103 4347 1107
rect 4356 1103 4363 1153
rect 4376 1107 4383 1233
rect 4396 1187 4403 1293
rect 4456 1287 4463 1293
rect 4456 1127 4463 1233
rect 4496 1147 4503 1293
rect 4536 1287 4543 1313
rect 4516 1127 4523 1173
rect 4556 1143 4563 1593
rect 4573 1553 4587 1567
rect 4613 1563 4627 1567
rect 4636 1563 4643 1593
rect 4613 1556 4643 1563
rect 4613 1553 4627 1556
rect 4653 1553 4667 1567
rect 4693 1553 4707 1567
rect 4576 1467 4583 1553
rect 4596 1347 4603 1533
rect 4616 1327 4623 1533
rect 4636 1447 4643 1533
rect 4656 1507 4663 1553
rect 4676 1407 4683 1533
rect 4696 1527 4703 1553
rect 4636 1327 4643 1393
rect 4676 1363 4683 1393
rect 4676 1356 4703 1363
rect 4696 1347 4703 1356
rect 4573 1293 4587 1307
rect 4633 1313 4647 1327
rect 4673 1313 4687 1327
rect 4693 1333 4707 1347
rect 4576 1247 4583 1293
rect 4576 1147 4583 1213
rect 4536 1136 4563 1143
rect 4433 1123 4447 1127
rect 4453 1123 4467 1127
rect 4333 1096 4363 1103
rect 4333 1093 4347 1096
rect 4413 1093 4427 1107
rect 4433 1116 4467 1123
rect 4433 1113 4447 1116
rect 4453 1113 4467 1116
rect 4473 1093 4487 1107
rect 4316 1067 4323 1093
rect 4276 867 4283 1013
rect 4336 987 4343 1093
rect 4416 1087 4423 1093
rect 4316 847 4323 913
rect 4356 847 4363 1053
rect 4416 1047 4423 1073
rect 4436 927 4443 1073
rect 4456 963 4463 1073
rect 4476 1047 4483 1093
rect 4456 956 4483 963
rect 4436 867 4443 893
rect 4193 843 4207 847
rect 4176 836 4207 843
rect 4193 833 4207 836
rect 4153 823 4167 827
rect 4153 816 4173 823
rect 4153 813 4167 816
rect 4213 813 4227 827
rect 4253 823 4267 827
rect 4276 823 4283 833
rect 4253 816 4283 823
rect 4253 813 4267 816
rect 4293 813 4307 827
rect 4373 833 4387 847
rect 4116 787 4123 813
rect 4016 647 4023 653
rect 3973 593 3987 607
rect 3976 547 3983 593
rect 3976 407 3983 533
rect 4056 527 4063 593
rect 4096 547 4103 733
rect 4176 647 4183 733
rect 4173 593 4187 607
rect 4176 567 4183 593
rect 3996 287 4003 333
rect 4073 333 4087 347
rect 4053 313 4067 327
rect 3956 176 3983 183
rect 3913 163 3927 167
rect 3896 156 3927 163
rect 3913 153 3927 156
rect 3873 133 3887 147
rect 3836 107 3843 133
rect 3896 87 3903 133
rect 3976 47 3983 176
rect 3996 167 4003 213
rect 4036 147 4043 233
rect 4056 227 4063 313
rect 4076 207 4083 333
rect 4096 227 4103 393
rect 4116 343 4123 373
rect 4196 367 4203 813
rect 4216 767 4223 813
rect 4236 747 4243 793
rect 4276 767 4283 793
rect 4296 787 4303 813
rect 4376 827 4383 833
rect 4396 807 4403 853
rect 4433 853 4447 867
rect 4216 627 4223 733
rect 4213 613 4227 627
rect 4236 607 4243 653
rect 4273 603 4287 607
rect 4296 603 4303 693
rect 4316 607 4323 633
rect 4356 627 4363 693
rect 4376 627 4383 753
rect 4396 647 4403 773
rect 4416 747 4423 793
rect 4436 767 4443 813
rect 4456 667 4463 933
rect 4476 907 4483 956
rect 4496 883 4503 913
rect 4536 907 4543 1136
rect 4573 1133 4587 1147
rect 4596 1143 4603 1273
rect 4596 1136 4623 1143
rect 4576 927 4583 1093
rect 4596 907 4603 1073
rect 4616 947 4623 1136
rect 4476 876 4503 883
rect 4476 827 4483 876
rect 4533 853 4547 867
rect 4513 833 4527 847
rect 4516 827 4523 833
rect 4396 627 4403 633
rect 4273 596 4303 603
rect 4273 593 4287 596
rect 4353 613 4367 627
rect 4393 613 4407 627
rect 4416 587 4423 653
rect 4456 627 4463 633
rect 4433 593 4447 607
rect 4453 613 4467 627
rect 4476 623 4483 793
rect 4536 747 4543 853
rect 4553 833 4567 847
rect 4556 787 4563 833
rect 4496 627 4503 633
rect 4493 623 4507 627
rect 4476 616 4507 623
rect 4493 613 4507 616
rect 4533 613 4547 627
rect 4296 407 4303 573
rect 4316 387 4323 573
rect 4436 527 4443 593
rect 4133 343 4147 347
rect 4116 336 4147 343
rect 4193 363 4207 367
rect 4193 356 4223 363
rect 4193 353 4207 356
rect 4133 333 4147 336
rect 4173 313 4187 327
rect 4033 133 4047 147
rect 4056 127 4063 173
rect 4076 167 4083 193
rect 4076 147 4083 153
rect 4116 147 4123 293
rect 4176 287 4183 313
rect 4216 307 4223 356
rect 4276 347 4283 373
rect 4293 363 4307 367
rect 4313 363 4327 367
rect 4336 363 4343 393
rect 4356 367 4363 453
rect 4293 356 4343 363
rect 4293 353 4307 356
rect 4313 353 4327 356
rect 4236 287 4243 333
rect 4316 303 4323 313
rect 4376 303 4383 333
rect 4316 296 4383 303
rect 4396 227 4403 513
rect 4516 407 4523 613
rect 4536 547 4543 613
rect 4556 427 4563 753
rect 4576 387 4583 893
rect 4616 847 4623 893
rect 4636 847 4643 1193
rect 4656 1147 4663 1193
rect 4676 1127 4683 1313
rect 4696 1147 4703 1293
rect 4716 1103 4723 1933
rect 4736 1167 4743 2133
rect 4756 1147 4763 2176
rect 4776 2167 4783 2233
rect 4776 1927 4783 2033
rect 4776 1487 4783 1893
rect 4776 1207 4783 1433
rect 4753 1133 4767 1147
rect 4733 1103 4747 1107
rect 4716 1096 4747 1103
rect 4733 1093 4747 1096
rect 4693 1073 4707 1087
rect 4656 867 4663 1013
rect 4696 987 4703 1073
rect 4716 907 4723 1073
rect 4736 907 4743 1073
rect 4756 1027 4763 1093
rect 4756 943 4763 993
rect 4776 967 4783 1153
rect 4756 936 4783 943
rect 4736 867 4743 873
rect 4756 867 4763 913
rect 4593 813 4607 827
rect 4673 833 4687 847
rect 4596 807 4603 813
rect 4633 793 4647 807
rect 4616 767 4623 793
rect 4636 787 4643 793
rect 4596 667 4603 693
rect 4596 627 4603 653
rect 4616 647 4623 673
rect 4656 667 4663 793
rect 4676 767 4683 833
rect 4696 787 4703 853
rect 4733 853 4747 867
rect 4716 747 4723 833
rect 4676 647 4683 713
rect 4716 647 4723 653
rect 4613 633 4627 647
rect 4653 643 4667 647
rect 4673 643 4687 647
rect 4593 613 4607 627
rect 4653 636 4687 643
rect 4653 633 4667 636
rect 4673 633 4687 636
rect 4713 633 4727 647
rect 4736 627 4743 633
rect 4733 613 4747 627
rect 4696 603 4703 613
rect 4696 596 4723 603
rect 4513 333 4527 347
rect 4413 313 4427 327
rect 4416 307 4423 313
rect 4053 113 4067 127
rect 4113 133 4127 147
rect 4156 127 4163 173
rect 4216 147 4223 193
rect 4213 133 4227 147
rect 4236 127 4243 213
rect 4256 147 4263 213
rect 4316 147 4323 173
rect 4313 133 4327 147
rect 4356 123 4363 153
rect 4396 147 4403 173
rect 4476 147 4483 193
rect 4516 147 4523 333
rect 4556 327 4563 333
rect 4573 313 4587 327
rect 4536 147 4543 293
rect 4576 287 4583 313
rect 4373 123 4387 127
rect 4356 116 4387 123
rect 4393 133 4407 147
rect 4373 113 4387 116
rect 4473 133 4487 147
rect 4533 133 4547 147
rect 4556 127 4563 273
rect 4596 163 4603 293
rect 4576 156 4603 163
rect 4576 147 4583 156
rect 4573 133 4587 147
rect 4553 113 4567 127
rect 4496 107 4503 113
rect 4136 -24 4143 13
rect 4176 -24 4183 33
rect 4616 27 4623 373
rect 4676 323 4683 593
rect 4716 367 4723 596
rect 4756 587 4763 653
rect 4713 353 4727 367
rect 4693 323 4707 327
rect 4676 316 4707 323
rect 4693 313 4707 316
rect 4656 167 4663 253
rect 4653 153 4667 167
rect 4713 143 4727 147
rect 4736 143 4743 413
rect 4756 147 4763 393
rect 4776 187 4783 936
rect 4713 136 4743 143
rect 4713 133 4727 136
rect 4216 -24 4223 13
<< m3contact >>
rect 313 4573 327 4587
rect 533 4573 547 4587
rect 433 4553 447 4567
rect 493 4553 507 4567
rect 413 4513 427 4527
rect 393 4493 407 4507
rect 213 4473 227 4487
rect 133 4453 147 4467
rect 193 4453 207 4467
rect 253 4473 267 4487
rect 233 4433 247 4447
rect 153 4413 167 4427
rect 273 4413 287 4427
rect 113 4393 127 4407
rect 153 4393 167 4407
rect 73 4193 87 4207
rect 33 4113 47 4127
rect 13 4013 27 4027
rect 93 4133 107 4147
rect 93 4113 107 4127
rect 53 3993 67 4007
rect 53 3973 67 3987
rect 73 3953 87 3967
rect 13 3933 27 3947
rect 153 4213 167 4227
rect 173 4213 187 4227
rect 133 4173 147 4187
rect 173 4173 187 4187
rect 213 4173 227 4187
rect 273 4193 287 4207
rect 253 4173 267 4187
rect 193 4153 207 4167
rect 253 4153 267 4167
rect 233 4133 247 4147
rect 193 4113 207 4127
rect 273 4113 287 4127
rect 173 4093 187 4107
rect 113 3993 127 4007
rect 113 3953 127 3967
rect 133 3973 147 3987
rect 213 4093 227 4107
rect 253 4053 267 4067
rect 193 3993 207 4007
rect 333 4453 347 4467
rect 413 4473 427 4487
rect 353 4433 367 4447
rect 453 4493 467 4507
rect 473 4493 487 4507
rect 493 4493 507 4507
rect 2693 4553 2707 4567
rect 733 4533 747 4547
rect 1133 4533 1147 4547
rect 593 4513 607 4527
rect 473 4453 487 4467
rect 333 4233 347 4247
rect 313 4173 327 4187
rect 333 4193 347 4207
rect 373 4193 387 4207
rect 353 4093 367 4107
rect 393 4093 407 4107
rect 293 4033 307 4047
rect 333 4033 347 4047
rect 393 4033 407 4047
rect 293 4013 307 4027
rect 213 3973 227 3987
rect 273 3973 287 3987
rect 313 3973 327 3987
rect 233 3933 247 3947
rect 213 3813 227 3827
rect 53 3693 67 3707
rect 73 3713 87 3727
rect 13 3673 27 3687
rect 153 3613 167 3627
rect 93 3513 107 3527
rect 113 3293 127 3307
rect 93 3213 107 3227
rect 133 3093 147 3107
rect 93 3033 107 3047
rect 113 3033 127 3047
rect 213 3473 227 3487
rect 213 3253 227 3267
rect 113 2973 127 2987
rect 33 2873 47 2887
rect 13 2493 27 2507
rect 93 2693 107 2707
rect 93 2613 107 2627
rect 173 2993 187 3007
rect 153 2773 167 2787
rect 113 2553 127 2567
rect 73 2513 87 2527
rect 93 2513 107 2527
rect 73 2453 87 2467
rect 93 2433 107 2447
rect 13 2273 27 2287
rect 33 2273 47 2287
rect 13 2233 27 2247
rect 93 2253 107 2267
rect 53 2093 67 2107
rect 13 2053 27 2067
rect 33 2053 47 2067
rect 113 2073 127 2087
rect 53 1973 67 1987
rect 253 3813 267 3827
rect 313 3693 327 3707
rect 273 3613 287 3627
rect 293 3493 307 3507
rect 313 3473 327 3487
rect 273 3453 287 3467
rect 253 3293 267 3307
rect 253 3273 267 3287
rect 293 3253 307 3267
rect 373 3973 387 3987
rect 673 4493 687 4507
rect 693 4493 707 4507
rect 733 4493 747 4507
rect 653 4473 667 4487
rect 813 4473 827 4487
rect 753 4453 767 4467
rect 753 4433 767 4447
rect 893 4493 907 4507
rect 953 4413 967 4427
rect 993 4513 1007 4527
rect 1073 4513 1087 4527
rect 1113 4513 1127 4527
rect 993 4453 1007 4467
rect 1053 4453 1067 4467
rect 1093 4453 1107 4467
rect 1013 4433 1027 4447
rect 1273 4513 1287 4527
rect 1233 4493 1247 4507
rect 1113 4413 1127 4427
rect 1413 4513 1427 4527
rect 1333 4493 1347 4507
rect 893 4313 907 4327
rect 1013 4313 1027 4327
rect 493 4253 507 4267
rect 533 4253 547 4267
rect 433 4213 447 4227
rect 473 4213 487 4227
rect 473 4193 487 4207
rect 453 4153 467 4167
rect 473 4033 487 4047
rect 453 4013 467 4027
rect 533 4233 547 4247
rect 693 4233 707 4247
rect 573 4193 587 4207
rect 633 4193 647 4207
rect 553 4153 567 4167
rect 593 4153 607 4167
rect 613 4153 627 4167
rect 573 4073 587 4087
rect 513 4033 527 4047
rect 413 3813 427 3827
rect 513 4013 527 4027
rect 493 3993 507 4007
rect 533 3993 547 4007
rect 593 4033 607 4047
rect 593 3993 607 4007
rect 573 3973 587 3987
rect 613 3953 627 3967
rect 773 4213 787 4227
rect 833 4213 847 4227
rect 673 4173 687 4187
rect 733 4193 747 4207
rect 813 4193 827 4207
rect 793 4173 807 4187
rect 713 4153 727 4167
rect 813 4153 827 4167
rect 653 4133 667 4147
rect 753 4073 767 4087
rect 793 4033 807 4047
rect 853 4033 867 4047
rect 653 4013 667 4027
rect 713 4013 727 4027
rect 673 3973 687 3987
rect 693 3993 707 4007
rect 733 3993 747 4007
rect 713 3973 727 3987
rect 593 3933 607 3947
rect 473 3793 487 3807
rect 593 3793 607 3807
rect 433 3773 447 3787
rect 553 3773 567 3787
rect 473 3753 487 3767
rect 533 3753 547 3767
rect 413 3713 427 3727
rect 493 3693 507 3707
rect 553 3733 567 3747
rect 393 3673 407 3687
rect 373 3513 387 3527
rect 353 3493 367 3507
rect 413 3513 427 3527
rect 513 3533 527 3547
rect 413 3473 427 3487
rect 413 3453 427 3467
rect 333 3273 347 3287
rect 453 3473 467 3487
rect 473 3493 487 3507
rect 673 3753 687 3767
rect 773 3973 787 3987
rect 773 3933 787 3947
rect 613 3653 627 3667
rect 673 3693 687 3707
rect 773 3733 787 3747
rect 713 3653 727 3667
rect 653 3553 667 3567
rect 573 3513 587 3527
rect 613 3513 627 3527
rect 533 3473 547 3487
rect 553 3493 567 3507
rect 593 3493 607 3507
rect 573 3473 587 3487
rect 433 3273 447 3287
rect 533 3273 547 3287
rect 573 3273 587 3287
rect 373 3253 387 3267
rect 393 3233 407 3247
rect 473 3253 487 3267
rect 513 3233 527 3247
rect 253 3133 267 3147
rect 253 3113 267 3127
rect 273 3113 287 3127
rect 233 2873 247 2887
rect 213 2793 227 2807
rect 353 3153 367 3167
rect 333 3133 347 3147
rect 393 3133 407 3147
rect 273 3053 287 3067
rect 313 3053 327 3067
rect 333 3053 347 3067
rect 293 3033 307 3047
rect 313 3013 327 3027
rect 313 2993 327 3007
rect 413 2993 427 3007
rect 353 2973 367 2987
rect 493 3213 507 3227
rect 1013 4213 1027 4227
rect 1113 4213 1127 4227
rect 1193 4213 1207 4227
rect 913 4193 927 4207
rect 913 4173 927 4187
rect 953 4193 967 4207
rect 993 4193 1007 4207
rect 933 4153 947 4167
rect 973 4153 987 4167
rect 913 4093 927 4107
rect 973 4033 987 4047
rect 813 3993 827 4007
rect 893 3993 907 4007
rect 873 3973 887 3987
rect 833 3953 847 3967
rect 1093 4173 1107 4187
rect 1193 4193 1207 4207
rect 1053 4153 1067 4167
rect 1013 4093 1027 4107
rect 1033 4093 1047 4107
rect 1013 4033 1027 4047
rect 1033 4033 1047 4047
rect 993 4013 1007 4027
rect 1033 4013 1047 4027
rect 1253 4173 1267 4187
rect 1313 4193 1327 4207
rect 1373 4473 1387 4487
rect 1473 4473 1487 4487
rect 1393 4433 1407 4447
rect 1453 4413 1467 4427
rect 1353 4213 1367 4227
rect 1233 4153 1247 4167
rect 1253 4153 1267 4167
rect 1293 4153 1307 4167
rect 1333 4153 1347 4167
rect 1133 4093 1147 4107
rect 1093 4053 1107 4067
rect 1213 4113 1227 4127
rect 1193 4033 1207 4047
rect 1273 4073 1287 4087
rect 993 3993 1007 4007
rect 933 3973 947 3987
rect 973 3973 987 3987
rect 973 3953 987 3967
rect 913 3933 927 3947
rect 813 3733 827 3747
rect 813 3693 827 3707
rect 913 3813 927 3827
rect 953 3713 967 3727
rect 913 3673 927 3687
rect 793 3593 807 3607
rect 753 3553 767 3567
rect 853 3553 867 3567
rect 813 3533 827 3547
rect 873 3533 887 3547
rect 673 3513 687 3527
rect 633 3493 647 3507
rect 653 3493 667 3507
rect 613 3273 627 3287
rect 593 3253 607 3267
rect 633 3253 647 3267
rect 733 3493 747 3507
rect 773 3513 787 3527
rect 773 3493 787 3507
rect 833 3493 847 3507
rect 673 3473 687 3487
rect 713 3473 727 3487
rect 673 3453 687 3467
rect 753 3433 767 3447
rect 533 3093 547 3107
rect 453 2993 467 3007
rect 613 3133 627 3147
rect 533 3033 547 3047
rect 373 2853 387 2867
rect 433 2853 447 2867
rect 333 2793 347 2807
rect 293 2773 307 2787
rect 313 2773 327 2787
rect 333 2773 347 2787
rect 373 2773 387 2787
rect 233 2593 247 2607
rect 233 2533 247 2547
rect 213 2513 227 2527
rect 213 2293 227 2307
rect 153 2153 167 2167
rect 153 2033 167 2047
rect 133 1953 147 1967
rect 133 1773 147 1787
rect 133 1753 147 1767
rect 33 1513 47 1527
rect 113 1273 127 1287
rect 393 2753 407 2767
rect 413 2773 427 2787
rect 393 2733 407 2747
rect 433 2733 447 2747
rect 293 2713 307 2727
rect 273 2573 287 2587
rect 353 2713 367 2727
rect 373 2613 387 2627
rect 313 2573 327 2587
rect 353 2573 367 2587
rect 693 3233 707 3247
rect 813 3473 827 3487
rect 1013 3973 1027 3987
rect 1073 3993 1087 4007
rect 1113 3993 1127 4007
rect 1133 3973 1147 3987
rect 1273 4013 1287 4027
rect 1233 3993 1247 4007
rect 1073 3933 1087 3947
rect 1053 3733 1067 3747
rect 1293 3973 1307 3987
rect 953 3573 967 3587
rect 933 3533 947 3547
rect 973 3553 987 3567
rect 993 3533 1007 3547
rect 933 3493 947 3507
rect 993 3513 1007 3527
rect 1033 3513 1047 3527
rect 913 3473 927 3487
rect 893 3453 907 3467
rect 1173 3733 1187 3747
rect 1173 3713 1187 3727
rect 1133 3633 1147 3647
rect 1093 3593 1107 3607
rect 1073 3453 1087 3467
rect 733 3193 747 3207
rect 773 3193 787 3207
rect 693 3153 707 3167
rect 593 2813 607 2827
rect 633 2813 647 2827
rect 553 2773 567 2787
rect 473 2753 487 2767
rect 513 2753 527 2767
rect 493 2693 507 2707
rect 493 2633 507 2647
rect 413 2613 427 2627
rect 453 2613 467 2627
rect 313 2533 327 2547
rect 333 2553 347 2567
rect 373 2553 387 2567
rect 373 2513 387 2527
rect 333 2493 347 2507
rect 253 2313 267 2327
rect 273 2273 287 2287
rect 293 2253 307 2267
rect 313 2213 327 2227
rect 433 2513 447 2527
rect 453 2533 467 2547
rect 473 2513 487 2527
rect 573 2713 587 2727
rect 573 2673 587 2687
rect 633 2793 647 2807
rect 653 2753 667 2767
rect 673 2773 687 2787
rect 673 2733 687 2747
rect 593 2633 607 2647
rect 513 2613 527 2627
rect 533 2613 547 2627
rect 593 2613 607 2627
rect 953 3233 967 3247
rect 1013 3233 1027 3247
rect 1053 3233 1067 3247
rect 793 3173 807 3187
rect 753 3073 767 3087
rect 793 3033 807 3047
rect 973 3053 987 3067
rect 1033 3053 1047 3067
rect 953 3033 967 3047
rect 953 2993 967 3007
rect 993 3033 1007 3047
rect 1153 3553 1167 3567
rect 1253 3693 1267 3707
rect 1213 3673 1227 3687
rect 1373 4173 1387 4187
rect 1453 4153 1467 4167
rect 1373 4053 1387 4067
rect 1593 4493 1607 4507
rect 1613 4433 1627 4447
rect 1673 4473 1687 4487
rect 1773 4473 1787 4487
rect 1813 4473 1827 4487
rect 1493 4173 1507 4187
rect 1453 4033 1467 4047
rect 1473 4033 1487 4047
rect 1473 4013 1487 4027
rect 1713 4433 1727 4447
rect 1733 4453 1747 4467
rect 1673 4393 1687 4407
rect 1573 4193 1587 4207
rect 1633 4173 1647 4187
rect 1613 4133 1627 4147
rect 1653 4093 1667 4107
rect 1733 4153 1747 4167
rect 1713 4113 1727 4127
rect 1693 4033 1707 4047
rect 1673 4013 1687 4027
rect 1433 3973 1447 3987
rect 1493 3973 1507 3987
rect 1573 3993 1587 4007
rect 1633 3973 1647 3987
rect 1653 3993 1667 4007
rect 1593 3953 1607 3967
rect 1673 3953 1687 3967
rect 1713 3973 1727 3987
rect 1733 3953 1747 3967
rect 1553 3753 1567 3767
rect 1373 3733 1387 3747
rect 1413 3713 1427 3727
rect 1393 3693 1407 3707
rect 1453 3733 1467 3747
rect 1473 3713 1487 3727
rect 1533 3733 1547 3747
rect 1553 3713 1567 3727
rect 1513 3693 1527 3707
rect 1573 3693 1587 3707
rect 1353 3673 1367 3687
rect 1393 3673 1407 3687
rect 1433 3673 1447 3687
rect 1333 3633 1347 3647
rect 1253 3533 1267 3547
rect 1333 3533 1347 3547
rect 1433 3553 1447 3567
rect 1293 3493 1307 3507
rect 1313 3453 1327 3467
rect 1253 3333 1267 3347
rect 1173 3153 1187 3167
rect 1093 3093 1107 3107
rect 1173 3073 1187 3087
rect 1213 3233 1227 3247
rect 1233 3193 1247 3207
rect 1273 3213 1287 3227
rect 1193 3053 1207 3067
rect 1133 3033 1147 3047
rect 973 2973 987 2987
rect 693 2713 707 2727
rect 953 2813 967 2827
rect 1013 2813 1027 2827
rect 733 2753 747 2767
rect 753 2733 767 2747
rect 773 2753 787 2767
rect 673 2653 687 2667
rect 673 2613 687 2627
rect 613 2593 627 2607
rect 613 2573 627 2587
rect 553 2553 567 2567
rect 533 2533 547 2547
rect 573 2533 587 2547
rect 593 2553 607 2567
rect 513 2513 527 2527
rect 653 2553 667 2567
rect 673 2533 687 2547
rect 593 2513 607 2527
rect 633 2513 647 2527
rect 493 2353 507 2367
rect 533 2353 547 2367
rect 413 2333 427 2347
rect 493 2333 507 2347
rect 453 2313 467 2327
rect 413 2293 427 2307
rect 353 2253 367 2267
rect 333 2193 347 2207
rect 313 2133 327 2147
rect 293 2113 307 2127
rect 253 2093 267 2107
rect 213 2033 227 2047
rect 233 2033 247 2047
rect 253 2053 267 2067
rect 193 2013 207 2027
rect 233 2013 247 2027
rect 213 1993 227 2007
rect 173 1773 187 1787
rect 273 1993 287 2007
rect 393 2133 407 2147
rect 473 2113 487 2127
rect 333 2073 347 2087
rect 313 2053 327 2067
rect 373 2073 387 2087
rect 433 2073 447 2087
rect 453 2053 467 2067
rect 513 2193 527 2207
rect 493 2053 507 2067
rect 333 2033 347 2047
rect 313 1833 327 1847
rect 293 1813 307 1827
rect 273 1793 287 1807
rect 293 1773 307 1787
rect 233 1753 247 1767
rect 173 1633 187 1647
rect 373 2033 387 2047
rect 353 2013 367 2027
rect 413 1993 427 2007
rect 353 1833 367 1847
rect 713 2653 727 2667
rect 733 2633 747 2647
rect 873 2733 887 2747
rect 853 2713 867 2727
rect 993 2773 1007 2787
rect 893 2713 907 2727
rect 873 2693 887 2707
rect 973 2713 987 2727
rect 1013 2713 1027 2727
rect 973 2673 987 2687
rect 933 2653 947 2667
rect 873 2633 887 2647
rect 853 2573 867 2587
rect 753 2533 767 2547
rect 793 2553 807 2567
rect 853 2533 867 2547
rect 753 2513 767 2527
rect 693 2493 707 2507
rect 713 2353 727 2367
rect 613 2333 627 2347
rect 553 2293 567 2307
rect 613 2233 627 2247
rect 573 2213 587 2227
rect 713 2273 727 2287
rect 633 2173 647 2187
rect 633 2153 647 2167
rect 633 2133 647 2147
rect 593 2113 607 2127
rect 733 2193 747 2207
rect 713 2153 727 2167
rect 673 2073 687 2087
rect 713 2073 727 2087
rect 733 2073 747 2087
rect 733 2013 747 2027
rect 733 1953 747 1967
rect 553 1833 567 1847
rect 693 1833 707 1847
rect 533 1813 547 1827
rect 413 1793 427 1807
rect 453 1793 467 1807
rect 473 1793 487 1807
rect 393 1753 407 1767
rect 433 1753 447 1767
rect 493 1773 507 1787
rect 513 1793 527 1807
rect 613 1813 627 1827
rect 593 1773 607 1787
rect 633 1773 647 1787
rect 673 1793 687 1807
rect 353 1653 367 1667
rect 313 1613 327 1627
rect 333 1613 347 1627
rect 173 1573 187 1587
rect 153 1553 167 1567
rect 153 1253 167 1267
rect 133 1213 147 1227
rect 33 1093 47 1107
rect 33 1073 47 1087
rect 93 1073 107 1087
rect 113 1093 127 1107
rect 133 1073 147 1087
rect 113 893 127 907
rect 93 813 107 827
rect 73 413 87 427
rect 133 633 147 647
rect 273 1593 287 1607
rect 293 1593 307 1607
rect 233 1553 247 1567
rect 213 1253 227 1267
rect 193 1213 207 1227
rect 173 1193 187 1207
rect 173 1173 187 1187
rect 393 1573 407 1587
rect 253 1413 267 1427
rect 293 1413 307 1427
rect 333 1293 347 1307
rect 453 1593 467 1607
rect 473 1573 487 1587
rect 633 1753 647 1767
rect 733 1793 747 1807
rect 533 1613 547 1627
rect 513 1573 527 1587
rect 593 1613 607 1627
rect 573 1573 587 1587
rect 553 1473 567 1487
rect 473 1353 487 1367
rect 533 1353 547 1367
rect 353 1273 367 1287
rect 373 1273 387 1287
rect 253 1213 267 1227
rect 233 1173 247 1187
rect 293 1193 307 1207
rect 173 1093 187 1107
rect 253 1113 267 1127
rect 273 1093 287 1107
rect 333 1113 347 1127
rect 313 1053 327 1067
rect 313 1013 327 1027
rect 173 773 187 787
rect 213 853 227 867
rect 253 853 267 867
rect 273 833 287 847
rect 293 853 307 867
rect 293 793 307 807
rect 173 633 187 647
rect 153 613 167 627
rect 213 613 227 627
rect 253 613 267 627
rect 233 593 247 607
rect 113 333 127 347
rect 173 393 187 407
rect 273 393 287 407
rect 453 1333 467 1347
rect 373 1213 387 1227
rect 393 1153 407 1167
rect 433 1133 447 1147
rect 413 1093 427 1107
rect 493 1333 507 1347
rect 513 1313 527 1327
rect 773 2493 787 2507
rect 813 2293 827 2307
rect 933 2513 947 2527
rect 973 2353 987 2367
rect 933 2293 947 2307
rect 853 2273 867 2287
rect 853 2233 867 2247
rect 833 2213 847 2227
rect 793 2073 807 2087
rect 773 2033 787 2047
rect 1073 2993 1087 3007
rect 1093 3013 1107 3027
rect 1133 2993 1147 3007
rect 1113 2973 1127 2987
rect 1273 3013 1287 3027
rect 1293 3033 1307 3047
rect 1213 2933 1227 2947
rect 1053 2773 1067 2787
rect 1093 2773 1107 2787
rect 1133 2773 1147 2787
rect 1173 2773 1187 2787
rect 1073 2613 1087 2627
rect 1133 2693 1147 2707
rect 1393 3513 1407 3527
rect 1413 3493 1427 3507
rect 1473 3513 1487 3527
rect 1453 3493 1467 3507
rect 1513 3493 1527 3507
rect 1373 3433 1387 3447
rect 1353 3173 1367 3187
rect 1393 3173 1407 3187
rect 1533 3413 1547 3427
rect 1513 3233 1527 3247
rect 1533 3173 1547 3187
rect 1553 3173 1567 3187
rect 1493 3133 1507 3147
rect 1433 3093 1447 3107
rect 1473 3093 1487 3107
rect 1353 3073 1367 3087
rect 1333 3053 1347 3067
rect 1333 3013 1347 3027
rect 1413 3033 1427 3047
rect 1253 2733 1267 2747
rect 1293 2733 1307 2747
rect 1233 2673 1247 2687
rect 1173 2633 1187 2647
rect 1213 2633 1227 2647
rect 1153 2613 1167 2627
rect 1153 2553 1167 2567
rect 1133 2533 1147 2547
rect 1193 2533 1207 2547
rect 1213 2553 1227 2567
rect 1233 2533 1247 2547
rect 1153 2513 1167 2527
rect 1153 2433 1167 2447
rect 1073 2353 1087 2367
rect 1033 2293 1047 2307
rect 1053 2273 1067 2287
rect 913 2233 927 2247
rect 933 2233 947 2247
rect 893 2213 907 2227
rect 873 2153 887 2167
rect 853 2093 867 2107
rect 873 2093 887 2107
rect 853 2053 867 2067
rect 833 2033 847 2047
rect 993 2253 1007 2267
rect 1013 2253 1027 2267
rect 973 2233 987 2247
rect 1033 2193 1047 2207
rect 953 2173 967 2187
rect 1013 2153 1027 2167
rect 913 2093 927 2107
rect 993 2093 1007 2107
rect 913 2053 927 2067
rect 873 2013 887 2027
rect 933 2033 947 2047
rect 953 2053 967 2067
rect 973 2013 987 2027
rect 813 1993 827 2007
rect 913 1993 927 2007
rect 1193 2253 1207 2267
rect 1153 2213 1167 2227
rect 1093 2193 1107 2207
rect 1153 2173 1167 2187
rect 1133 2113 1147 2127
rect 1033 2093 1047 2107
rect 1013 2073 1027 2087
rect 1073 2093 1087 2107
rect 1233 2233 1247 2247
rect 1193 2133 1207 2147
rect 1113 2053 1127 2067
rect 1153 2073 1167 2087
rect 1153 2053 1167 2067
rect 1013 2033 1027 2047
rect 1073 2033 1087 2047
rect 1173 2033 1187 2047
rect 1213 2053 1227 2067
rect 1233 2033 1247 2047
rect 813 1953 827 1967
rect 993 1953 1007 1967
rect 813 1833 827 1847
rect 773 1813 787 1827
rect 753 1653 767 1667
rect 733 1633 747 1647
rect 693 1613 707 1627
rect 673 1593 687 1607
rect 813 1793 827 1807
rect 793 1773 807 1787
rect 833 1773 847 1787
rect 833 1753 847 1767
rect 813 1713 827 1727
rect 893 1793 907 1807
rect 913 1813 927 1827
rect 873 1773 887 1787
rect 933 1653 947 1667
rect 853 1613 867 1627
rect 873 1593 887 1607
rect 773 1473 787 1487
rect 893 1473 907 1487
rect 813 1413 827 1427
rect 773 1353 787 1367
rect 913 1413 927 1427
rect 813 1333 827 1347
rect 853 1333 867 1347
rect 593 1313 607 1327
rect 553 1253 567 1267
rect 573 1213 587 1227
rect 513 1193 527 1207
rect 553 1193 567 1207
rect 473 1093 487 1107
rect 493 1093 507 1107
rect 533 1133 547 1147
rect 613 1293 627 1307
rect 633 1313 647 1327
rect 693 1313 707 1327
rect 733 1313 747 1327
rect 773 1313 787 1327
rect 753 1293 767 1307
rect 673 1273 687 1287
rect 833 1293 847 1307
rect 633 1153 647 1167
rect 613 1113 627 1127
rect 373 1073 387 1087
rect 453 1073 467 1087
rect 513 1073 527 1087
rect 713 1253 727 1267
rect 653 1113 667 1127
rect 633 1053 647 1067
rect 373 1013 387 1027
rect 353 893 367 907
rect 333 853 347 867
rect 353 833 367 847
rect 373 813 387 827
rect 393 833 407 847
rect 453 833 467 847
rect 333 793 347 807
rect 413 793 427 807
rect 353 773 367 787
rect 533 893 547 907
rect 513 813 527 827
rect 593 873 607 887
rect 533 793 547 807
rect 593 793 607 807
rect 313 633 327 647
rect 393 633 407 647
rect 373 613 387 627
rect 333 593 347 607
rect 433 613 447 627
rect 453 593 467 607
rect 273 353 287 367
rect 233 273 247 287
rect 233 213 247 227
rect 173 153 187 167
rect 113 133 127 147
rect 493 733 507 747
rect 633 853 647 867
rect 693 1073 707 1087
rect 913 1293 927 1307
rect 953 1633 967 1647
rect 1053 2013 1067 2027
rect 1033 1753 1047 1767
rect 1093 1813 1107 1827
rect 1073 1633 1087 1647
rect 1053 1413 1067 1427
rect 1153 1813 1167 1827
rect 1113 1553 1127 1567
rect 1133 1573 1147 1587
rect 1153 1533 1167 1547
rect 1153 1473 1167 1487
rect 1093 1373 1107 1387
rect 1133 1373 1147 1387
rect 993 1353 1007 1367
rect 1093 1353 1107 1367
rect 1093 1333 1107 1347
rect 953 1313 967 1327
rect 1053 1313 1067 1327
rect 913 1273 927 1287
rect 933 1273 947 1287
rect 873 1173 887 1187
rect 673 1053 687 1067
rect 713 1053 727 1067
rect 753 1053 767 1067
rect 733 893 747 907
rect 713 873 727 887
rect 673 853 687 867
rect 693 833 707 847
rect 653 753 667 767
rect 593 613 607 627
rect 593 593 607 607
rect 793 853 807 867
rect 893 1133 907 1147
rect 853 1113 867 1127
rect 893 1113 907 1127
rect 1013 1233 1027 1247
rect 1033 1233 1047 1247
rect 973 1193 987 1207
rect 973 1173 987 1187
rect 953 1153 967 1167
rect 913 1073 927 1087
rect 933 1073 947 1087
rect 1013 1133 1027 1147
rect 1073 1173 1087 1187
rect 1053 1153 1067 1167
rect 993 1093 1007 1107
rect 1093 1153 1107 1167
rect 1113 1153 1127 1167
rect 973 893 987 907
rect 1373 2813 1387 2827
rect 1313 2633 1327 2647
rect 1273 2613 1287 2627
rect 1293 2533 1307 2547
rect 1453 3073 1467 3087
rect 1473 2733 1487 2747
rect 1593 3653 1607 3667
rect 1593 3513 1607 3527
rect 1713 3653 1727 3667
rect 1693 3573 1707 3587
rect 1893 4493 1907 4507
rect 1913 4493 1927 4507
rect 1793 4333 1807 4347
rect 1793 4213 1807 4227
rect 1773 4153 1787 4167
rect 1813 4153 1827 4167
rect 1933 4473 1947 4487
rect 2113 4493 2127 4507
rect 2073 4473 2087 4487
rect 2093 4453 2107 4467
rect 2293 4473 2307 4487
rect 2193 4453 2207 4467
rect 2213 4433 2227 4447
rect 2173 4413 2187 4427
rect 2053 4393 2067 4407
rect 2213 4393 2227 4407
rect 2053 4373 2067 4387
rect 2013 4333 2027 4347
rect 1953 4193 1967 4207
rect 1833 4073 1847 4087
rect 1873 4053 1887 4067
rect 1833 4013 1847 4027
rect 1793 3993 1807 4007
rect 1813 3973 1827 3987
rect 1893 4013 1907 4027
rect 1893 3993 1907 4007
rect 1913 3973 1927 3987
rect 1933 3953 1947 3967
rect 1973 4133 1987 4147
rect 2093 4213 2107 4227
rect 2133 4213 2147 4227
rect 2433 4493 2447 4507
rect 2453 4493 2467 4507
rect 2533 4493 2547 4507
rect 2413 4473 2427 4487
rect 2393 4453 2407 4467
rect 2793 4573 2807 4587
rect 2553 4473 2567 4487
rect 2593 4473 2607 4487
rect 2613 4453 2627 4467
rect 2353 4433 2367 4447
rect 2393 4413 2407 4427
rect 2313 4393 2327 4407
rect 2253 4373 2267 4387
rect 2233 4213 2247 4227
rect 2133 4173 2147 4187
rect 2113 4153 2127 4167
rect 2233 4173 2247 4187
rect 2153 4153 2167 4167
rect 2173 4153 2187 4167
rect 2333 4253 2347 4267
rect 2593 4433 2607 4447
rect 2513 4393 2527 4407
rect 2573 4393 2587 4407
rect 2413 4353 2427 4367
rect 2433 4313 2447 4327
rect 2413 4253 2427 4267
rect 2393 4233 2407 4247
rect 2373 4213 2387 4227
rect 2273 4173 2287 4187
rect 2293 4193 2307 4207
rect 2313 4173 2327 4187
rect 2353 4173 2367 4187
rect 2393 4153 2407 4167
rect 2253 4133 2267 4147
rect 2333 4073 2347 4087
rect 2133 4053 2147 4067
rect 2113 4013 2127 4027
rect 2013 3993 2027 4007
rect 1993 3973 2007 3987
rect 2033 3973 2047 3987
rect 2053 3993 2067 4007
rect 2093 3973 2107 3987
rect 2173 4033 2187 4047
rect 2213 4013 2227 4027
rect 2273 4013 2287 4027
rect 2333 4013 2347 4027
rect 2393 4013 2407 4027
rect 2193 3953 2207 3967
rect 2313 3973 2327 3987
rect 2293 3953 2307 3967
rect 1813 3933 1827 3947
rect 1953 3933 1967 3947
rect 1993 3933 2007 3947
rect 2253 3933 2267 3947
rect 1793 3633 1807 3647
rect 1813 3633 1827 3647
rect 1753 3613 1767 3627
rect 1793 3613 1807 3627
rect 1693 3493 1707 3507
rect 1613 3453 1627 3467
rect 1673 3433 1687 3447
rect 1593 3413 1607 3427
rect 1573 3093 1587 3107
rect 1653 3273 1667 3287
rect 1613 3233 1627 3247
rect 1633 3213 1647 3227
rect 1653 3073 1667 3087
rect 1613 3053 1627 3067
rect 1633 3053 1647 3067
rect 1533 3033 1547 3047
rect 1593 3033 1607 3047
rect 1513 2913 1527 2927
rect 1733 3253 1747 3267
rect 1713 3213 1727 3227
rect 1753 3233 1767 3247
rect 1693 3193 1707 3207
rect 1733 3193 1747 3207
rect 1693 3173 1707 3187
rect 1673 3053 1687 3067
rect 1773 3133 1787 3147
rect 1733 3053 1747 3067
rect 2173 3733 2187 3747
rect 2033 3713 2047 3727
rect 2113 3713 2127 3727
rect 2133 3673 2147 3687
rect 2173 3673 2187 3687
rect 2093 3633 2107 3647
rect 2153 3633 2167 3647
rect 2053 3593 2067 3607
rect 2193 3593 2207 3607
rect 1973 3573 1987 3587
rect 2053 3573 2067 3587
rect 2153 3573 2167 3587
rect 1833 3533 1847 3547
rect 1833 3493 1847 3507
rect 1993 3533 2007 3547
rect 1973 3493 1987 3507
rect 2013 3493 2027 3507
rect 2033 3513 2047 3527
rect 1973 3473 1987 3487
rect 2133 3553 2147 3567
rect 2073 3473 2087 3487
rect 2093 3493 2107 3507
rect 2053 3453 2067 3467
rect 2113 3453 2127 3467
rect 1933 3433 1947 3447
rect 2053 3333 2067 3347
rect 1913 3273 1927 3287
rect 1913 3253 1927 3267
rect 1953 3253 1967 3267
rect 1813 3233 1827 3247
rect 1853 3233 1867 3247
rect 1833 3113 1847 3127
rect 1813 3053 1827 3067
rect 1773 3033 1787 3047
rect 1733 2993 1747 3007
rect 1673 2913 1687 2927
rect 1653 2893 1667 2907
rect 1573 2813 1587 2827
rect 1553 2793 1567 2807
rect 1513 2773 1527 2787
rect 1573 2753 1587 2767
rect 1493 2713 1507 2727
rect 1433 2633 1447 2647
rect 1473 2633 1487 2647
rect 1353 2613 1367 2627
rect 1393 2613 1407 2627
rect 1353 2553 1367 2567
rect 1433 2553 1447 2567
rect 1333 2513 1347 2527
rect 1353 2533 1367 2547
rect 1373 2413 1387 2427
rect 1453 2413 1467 2427
rect 1433 2373 1447 2387
rect 1413 2353 1427 2367
rect 1333 2253 1347 2267
rect 1373 2233 1387 2247
rect 1273 2093 1287 2107
rect 1293 2093 1307 2107
rect 1313 2073 1327 2087
rect 1373 2073 1387 2087
rect 1373 2033 1387 2047
rect 1413 2093 1427 2107
rect 1413 2053 1427 2067
rect 1253 2013 1267 2027
rect 1253 1833 1267 1847
rect 1193 1813 1207 1827
rect 1233 1813 1247 1827
rect 1213 1773 1227 1787
rect 1413 1813 1427 1827
rect 1273 1793 1287 1807
rect 1213 1593 1227 1607
rect 1193 1573 1207 1587
rect 1233 1573 1247 1587
rect 1293 1773 1307 1787
rect 1333 1793 1347 1807
rect 1313 1753 1327 1767
rect 1353 1753 1367 1767
rect 1273 1573 1287 1587
rect 1233 1553 1247 1567
rect 1193 1393 1207 1407
rect 1173 1353 1187 1367
rect 1153 1273 1167 1287
rect 1373 1613 1387 1627
rect 1293 1533 1307 1547
rect 1233 1373 1247 1387
rect 1353 1373 1367 1387
rect 1253 1313 1267 1327
rect 1273 1173 1287 1187
rect 1193 1153 1207 1167
rect 1233 1153 1247 1167
rect 773 833 787 847
rect 793 813 807 827
rect 813 833 827 847
rect 833 793 847 807
rect 773 633 787 647
rect 913 853 927 867
rect 1013 853 1027 867
rect 1093 853 1107 867
rect 1213 1133 1227 1147
rect 1313 1313 1327 1327
rect 1413 1593 1427 1607
rect 1493 2613 1507 2627
rect 1513 2613 1527 2627
rect 1473 2373 1487 2387
rect 1453 2273 1467 2287
rect 1613 2733 1627 2747
rect 1633 2733 1647 2747
rect 1633 2713 1647 2727
rect 1673 2713 1687 2727
rect 1553 2553 1567 2567
rect 1533 2353 1547 2367
rect 1593 2293 1607 2307
rect 1493 2253 1507 2267
rect 1533 2253 1547 2267
rect 1573 2193 1587 2207
rect 1473 2093 1487 2107
rect 1493 2073 1507 2087
rect 1733 2953 1747 2967
rect 1773 2993 1787 3007
rect 1753 2893 1767 2907
rect 1793 2893 1807 2907
rect 1713 2733 1727 2747
rect 1733 2733 1747 2747
rect 1693 2673 1707 2687
rect 1653 2573 1667 2587
rect 1713 2573 1727 2587
rect 1693 2553 1707 2567
rect 1673 2513 1687 2527
rect 1693 2253 1707 2267
rect 1713 2233 1727 2247
rect 1773 2693 1787 2707
rect 1893 3213 1907 3227
rect 1873 3173 1887 3187
rect 1873 3153 1887 3167
rect 1973 3213 1987 3227
rect 2013 3233 2027 3247
rect 1993 3193 2007 3207
rect 2033 3153 2047 3167
rect 1953 3073 1967 3087
rect 1933 3053 1947 3067
rect 1853 3033 1867 3047
rect 1873 3033 1887 3047
rect 1853 3013 1867 3027
rect 1893 2993 1907 3007
rect 1913 2993 1927 3007
rect 1833 2973 1847 2987
rect 1913 2953 1927 2967
rect 1813 2773 1827 2787
rect 1873 2773 1887 2787
rect 1853 2733 1867 2747
rect 1993 3053 2007 3067
rect 1953 2973 1967 2987
rect 1993 2793 2007 2807
rect 1953 2773 1967 2787
rect 1913 2753 1927 2767
rect 1933 2753 1947 2767
rect 1833 2713 1847 2727
rect 1813 2673 1827 2687
rect 1793 2653 1807 2667
rect 1773 2553 1787 2567
rect 1853 2613 1867 2627
rect 1913 2713 1927 2727
rect 1813 2553 1827 2567
rect 1853 2553 1867 2567
rect 1893 2313 1907 2327
rect 1793 2273 1807 2287
rect 1833 2273 1847 2287
rect 1853 2273 1867 2287
rect 1873 2253 1887 2267
rect 1833 2233 1847 2247
rect 1853 2233 1867 2247
rect 1893 2233 1907 2247
rect 1773 2193 1787 2207
rect 1753 2173 1767 2187
rect 1773 2153 1787 2167
rect 1813 2153 1827 2167
rect 1713 2133 1727 2147
rect 1633 2113 1647 2127
rect 1653 2113 1667 2127
rect 1613 2073 1627 2087
rect 1733 2113 1747 2127
rect 1753 2113 1767 2127
rect 1633 2053 1647 2067
rect 1833 2133 1847 2147
rect 1773 2073 1787 2087
rect 1793 2073 1807 2087
rect 1933 2693 1947 2707
rect 1993 2653 2007 2667
rect 1933 2253 1947 2267
rect 2033 2733 2047 2747
rect 2033 2653 2047 2667
rect 2013 2613 2027 2627
rect 2013 2293 2027 2307
rect 1993 2253 2007 2267
rect 1953 2233 1967 2247
rect 1933 2173 1947 2187
rect 1893 2153 1907 2167
rect 1913 2153 1927 2167
rect 1873 2093 1887 2107
rect 1853 2073 1867 2087
rect 1733 1933 1747 1947
rect 1533 1793 1547 1807
rect 1573 1793 1587 1807
rect 1593 1793 1607 1807
rect 1473 1613 1487 1627
rect 1433 1393 1447 1407
rect 1413 1373 1427 1387
rect 1433 1313 1447 1327
rect 1453 1333 1467 1347
rect 1413 1273 1427 1287
rect 1293 1133 1307 1147
rect 1333 1133 1347 1147
rect 1253 1093 1267 1107
rect 1293 1093 1307 1107
rect 1173 1073 1187 1087
rect 1293 1073 1307 1087
rect 1253 1053 1267 1067
rect 1153 873 1167 887
rect 873 833 887 847
rect 893 793 907 807
rect 1073 813 1087 827
rect 993 773 1007 787
rect 933 693 947 707
rect 753 433 767 447
rect 753 413 767 427
rect 873 653 887 667
rect 853 613 867 627
rect 893 613 907 627
rect 913 633 927 647
rect 1013 673 1027 687
rect 1113 793 1127 807
rect 1093 773 1107 787
rect 1133 673 1147 687
rect 953 653 967 667
rect 993 653 1007 667
rect 1053 653 1067 667
rect 1073 653 1087 667
rect 953 613 967 627
rect 1033 633 1047 647
rect 1073 633 1087 647
rect 1093 633 1107 647
rect 1033 593 1047 607
rect 853 433 867 447
rect 493 393 507 407
rect 553 393 567 407
rect 633 393 647 407
rect 793 393 807 407
rect 833 393 847 407
rect 473 373 487 387
rect 353 353 367 367
rect 373 333 387 347
rect 393 353 407 367
rect 513 353 527 367
rect 533 373 547 387
rect 573 373 587 387
rect 373 273 387 287
rect 333 213 347 227
rect 333 193 347 207
rect 313 173 327 187
rect 353 173 367 187
rect 473 313 487 327
rect 433 273 447 287
rect 453 273 467 287
rect 433 213 447 227
rect 413 173 427 187
rect 253 153 267 167
rect 293 153 307 167
rect 313 133 327 147
rect 353 153 367 167
rect 513 213 527 227
rect 493 173 507 187
rect 513 173 527 187
rect 433 133 447 147
rect 273 113 287 127
rect 353 113 367 127
rect 493 133 507 147
rect 473 113 487 127
rect 753 373 767 387
rect 793 373 807 387
rect 593 353 607 367
rect 613 333 627 347
rect 653 333 667 347
rect 693 353 707 367
rect 733 353 747 367
rect 773 333 787 347
rect 833 353 847 367
rect 833 333 847 347
rect 653 313 667 327
rect 673 313 687 327
rect 753 313 767 327
rect 573 293 587 307
rect 813 293 827 307
rect 833 293 847 307
rect 633 213 647 227
rect 753 213 767 227
rect 553 193 567 207
rect 613 193 627 207
rect 713 193 727 207
rect 673 173 687 187
rect 693 133 707 147
rect 873 393 887 407
rect 1113 393 1127 407
rect 1193 893 1207 907
rect 1233 853 1247 867
rect 1273 853 1287 867
rect 1353 893 1367 907
rect 1393 893 1407 907
rect 1373 833 1387 847
rect 1213 813 1227 827
rect 1253 813 1267 827
rect 1233 713 1247 727
rect 1193 693 1207 707
rect 1433 1133 1447 1147
rect 1653 1773 1667 1787
rect 1913 2133 1927 2147
rect 1973 2133 1987 2147
rect 1933 2053 1947 2067
rect 2073 3213 2087 3227
rect 2113 3213 2127 3227
rect 2113 3173 2127 3187
rect 2073 3033 2087 3047
rect 2353 3993 2367 4007
rect 2373 3973 2387 3987
rect 2333 3893 2347 3907
rect 2413 3893 2427 3907
rect 2553 4213 2567 4227
rect 2513 4193 2527 4207
rect 2473 4133 2487 4147
rect 2533 4113 2547 4127
rect 2493 4093 2507 4107
rect 2633 4373 2647 4387
rect 2713 4273 2727 4287
rect 2633 4213 2647 4227
rect 2593 4193 2607 4207
rect 2573 4173 2587 4187
rect 2673 4193 2687 4207
rect 2593 4153 2607 4167
rect 2593 4133 2607 4147
rect 2553 4073 2567 4087
rect 2533 4033 2547 4047
rect 2473 4013 2487 4027
rect 2513 4013 2527 4027
rect 2493 3993 2507 4007
rect 2453 3973 2467 3987
rect 2453 3953 2467 3967
rect 2553 3973 2567 3987
rect 2673 4153 2687 4167
rect 2653 4133 2667 4147
rect 2613 4073 2627 4087
rect 2653 4053 2667 4067
rect 2593 3953 2607 3967
rect 2633 3973 2647 3987
rect 2873 4573 2887 4587
rect 2933 4533 2947 4547
rect 3073 4533 3087 4547
rect 2893 4473 2907 4487
rect 2853 4313 2867 4327
rect 2813 4293 2827 4307
rect 2853 4253 2867 4267
rect 3153 4553 3167 4567
rect 3933 4533 3947 4547
rect 3793 4513 3807 4527
rect 3213 4493 3227 4507
rect 3293 4493 3307 4507
rect 3373 4493 3387 4507
rect 3433 4493 3447 4507
rect 3013 4473 3027 4487
rect 2973 4453 2987 4467
rect 2953 4433 2967 4447
rect 2993 4433 3007 4447
rect 3033 4433 3047 4447
rect 3013 4413 3027 4427
rect 2913 4293 2927 4307
rect 2933 4293 2947 4307
rect 2993 4293 3007 4307
rect 2773 4193 2787 4207
rect 2793 4193 2807 4207
rect 2813 4193 2827 4207
rect 2793 4153 2807 4167
rect 2753 4113 2767 4127
rect 2693 4093 2707 4107
rect 2733 4093 2747 4107
rect 2833 4053 2847 4067
rect 2713 4033 2727 4047
rect 2753 4033 2767 4047
rect 2673 3993 2687 4007
rect 2753 4013 2767 4027
rect 2893 4233 2907 4247
rect 2873 4173 2887 4187
rect 2913 4193 2927 4207
rect 2953 4193 2967 4207
rect 2913 4173 2927 4187
rect 2893 4153 2907 4167
rect 2893 4093 2907 4107
rect 2893 4073 2907 4087
rect 2713 3993 2727 4007
rect 3153 4393 3167 4407
rect 3113 4253 3127 4267
rect 3033 4233 3047 4247
rect 3033 4213 3047 4227
rect 3073 4213 3087 4227
rect 3053 4193 3067 4207
rect 3133 4193 3147 4207
rect 3093 4173 3107 4187
rect 2973 4133 2987 4147
rect 2973 4073 2987 4087
rect 2973 4053 2987 4067
rect 2913 4013 2927 4027
rect 2953 4013 2967 4027
rect 2733 3973 2747 3987
rect 2753 3973 2767 3987
rect 2653 3953 2667 3967
rect 2493 3933 2507 3947
rect 2593 3913 2607 3927
rect 2613 3893 2627 3907
rect 2553 3773 2567 3787
rect 2693 3773 2707 3787
rect 2353 3753 2367 3767
rect 2273 3713 2287 3727
rect 2253 3693 2267 3707
rect 2293 3693 2307 3707
rect 2313 3713 2327 3727
rect 2433 3753 2447 3767
rect 2453 3753 2467 3767
rect 2373 3733 2387 3747
rect 2413 3733 2427 3747
rect 2433 3713 2447 3727
rect 2413 3673 2427 3687
rect 2353 3633 2367 3647
rect 2333 3553 2347 3567
rect 2233 3533 2247 3547
rect 2293 3533 2307 3547
rect 2173 3513 2187 3527
rect 2193 3493 2207 3507
rect 2233 3473 2247 3487
rect 2333 3493 2347 3507
rect 2393 3653 2407 3667
rect 2393 3613 2407 3627
rect 2393 3553 2407 3567
rect 2573 3733 2587 3747
rect 2473 3693 2487 3707
rect 2493 3713 2507 3727
rect 2513 3673 2527 3687
rect 2493 3613 2507 3627
rect 2453 3573 2467 3587
rect 2453 3553 2467 3567
rect 2373 3533 2387 3547
rect 2413 3533 2427 3547
rect 2433 3533 2447 3547
rect 2313 3473 2327 3487
rect 2273 3453 2287 3467
rect 2593 3693 2607 3707
rect 2693 3733 2707 3747
rect 2633 3713 2647 3727
rect 2653 3713 2667 3727
rect 2733 3693 2747 3707
rect 2613 3673 2627 3687
rect 2673 3673 2687 3687
rect 2573 3653 2587 3667
rect 2593 3653 2607 3667
rect 2553 3613 2567 3627
rect 2613 3613 2627 3627
rect 2573 3573 2587 3587
rect 2553 3513 2567 3527
rect 2433 3473 2447 3487
rect 2513 3493 2527 3507
rect 2473 3473 2487 3487
rect 2533 3473 2547 3487
rect 2593 3493 2607 3507
rect 2593 3453 2607 3467
rect 2293 3313 2307 3327
rect 2413 3313 2427 3327
rect 2193 3273 2207 3287
rect 2213 3273 2227 3287
rect 2153 3153 2167 3167
rect 2133 2973 2147 2987
rect 2193 3193 2207 3207
rect 2253 3293 2267 3307
rect 2213 3053 2227 3067
rect 2233 3053 2247 3067
rect 2213 3013 2227 3027
rect 2313 3273 2327 3287
rect 2373 3233 2387 3247
rect 2293 3073 2307 3087
rect 2373 3133 2387 3147
rect 2333 3033 2347 3047
rect 2213 2913 2227 2927
rect 2213 2853 2227 2867
rect 2173 2833 2187 2847
rect 2073 2813 2087 2827
rect 2173 2813 2187 2827
rect 2093 2753 2107 2767
rect 2113 2753 2127 2767
rect 2153 2733 2167 2747
rect 2133 2593 2147 2607
rect 2113 2513 2127 2527
rect 2113 2193 2127 2207
rect 1973 2033 1987 2047
rect 1973 1853 1987 1867
rect 1733 1753 1747 1767
rect 1893 1813 1907 1827
rect 1833 1773 1847 1787
rect 1853 1793 1867 1807
rect 1793 1753 1807 1767
rect 1913 1753 1927 1767
rect 1933 1753 1947 1767
rect 1813 1713 1827 1727
rect 1873 1713 1887 1727
rect 1893 1713 1907 1727
rect 1633 1693 1647 1707
rect 1693 1693 1707 1707
rect 1633 1613 1647 1627
rect 1593 1593 1607 1607
rect 1873 1633 1887 1647
rect 1773 1593 1787 1607
rect 1713 1573 1727 1587
rect 1833 1573 1847 1587
rect 1853 1593 1867 1607
rect 1953 1713 1967 1727
rect 2053 2093 2067 2107
rect 2033 2053 2047 2067
rect 2033 1853 2047 1867
rect 2213 2773 2227 2787
rect 2213 2713 2227 2727
rect 2193 2693 2207 2707
rect 2173 2573 2187 2587
rect 2153 2533 2167 2547
rect 2253 2973 2267 2987
rect 2353 3013 2367 3027
rect 2393 3113 2407 3127
rect 2453 3233 2467 3247
rect 2493 3213 2507 3227
rect 2553 3233 2567 3247
rect 2553 3193 2567 3207
rect 2473 3173 2487 3187
rect 2533 3173 2547 3187
rect 2553 3153 2567 3167
rect 2573 3153 2587 3167
rect 2413 3093 2427 3107
rect 2473 3093 2487 3107
rect 2513 3093 2527 3107
rect 2553 3093 2567 3107
rect 2433 3053 2447 3067
rect 2453 3013 2467 3027
rect 2493 3013 2507 3027
rect 2593 3073 2607 3087
rect 2593 3053 2607 3067
rect 2593 3033 2607 3047
rect 2533 2993 2547 3007
rect 2553 3013 2567 3027
rect 2573 3013 2587 3027
rect 2573 2993 2587 3007
rect 2513 2973 2527 2987
rect 2413 2953 2427 2967
rect 2333 2933 2347 2947
rect 2433 2933 2447 2947
rect 2393 2893 2407 2907
rect 2273 2853 2287 2867
rect 2293 2853 2307 2867
rect 2293 2833 2307 2847
rect 2253 2713 2267 2727
rect 2233 2653 2247 2667
rect 2213 2513 2227 2527
rect 2273 2593 2287 2607
rect 2213 2373 2227 2387
rect 2173 2313 2187 2327
rect 2153 2293 2167 2307
rect 2233 2253 2247 2267
rect 2173 2233 2187 2247
rect 2133 2113 2147 2127
rect 2153 2113 2167 2127
rect 2253 2193 2267 2207
rect 2193 2133 2207 2147
rect 2133 2033 2147 2047
rect 2173 2033 2187 2047
rect 2093 2013 2107 2027
rect 2253 2053 2267 2067
rect 2273 2033 2287 2047
rect 2233 2013 2247 2027
rect 2213 1993 2227 2007
rect 2093 1973 2107 1987
rect 2173 1933 2187 1947
rect 2073 1833 2087 1847
rect 2013 1813 2027 1827
rect 2313 2673 2327 2687
rect 2453 2853 2467 2867
rect 2433 2733 2447 2747
rect 2533 2833 2547 2847
rect 2553 2813 2567 2827
rect 2653 3593 2667 3607
rect 2773 3953 2787 3967
rect 2873 3993 2887 4007
rect 2913 3973 2927 3987
rect 2933 3993 2947 4007
rect 2793 3933 2807 3947
rect 2873 3913 2887 3927
rect 2793 3833 2807 3847
rect 2853 3793 2867 3807
rect 2953 3853 2967 3867
rect 2873 3773 2887 3787
rect 2833 3733 2847 3747
rect 2933 3733 2947 3747
rect 3253 4473 3267 4487
rect 3233 4433 3247 4447
rect 3213 4373 3227 4387
rect 3193 4353 3207 4367
rect 3193 4293 3207 4307
rect 3313 4393 3327 4407
rect 3393 4453 3407 4467
rect 3413 4473 3427 4487
rect 3353 4433 3367 4447
rect 3333 4373 3347 4387
rect 3253 4273 3267 4287
rect 3273 4273 3287 4287
rect 3373 4273 3387 4287
rect 3713 4493 3727 4507
rect 3613 4473 3627 4487
rect 3473 4453 3487 4467
rect 3493 4453 3507 4467
rect 3453 4413 3467 4427
rect 3533 4453 3547 4467
rect 3553 4433 3567 4447
rect 3493 4393 3507 4407
rect 3513 4393 3527 4407
rect 3973 4513 3987 4527
rect 4053 4493 4067 4507
rect 4133 4493 4147 4507
rect 4153 4493 4167 4507
rect 4213 4493 4227 4507
rect 3613 4433 3627 4447
rect 3673 4453 3687 4467
rect 3733 4453 3747 4467
rect 3753 4473 3767 4487
rect 3813 4453 3827 4467
rect 3833 4473 3847 4487
rect 3853 4453 3867 4467
rect 3673 4433 3687 4447
rect 3633 4413 3647 4427
rect 3573 4393 3587 4407
rect 3693 4393 3707 4407
rect 3513 4273 3527 4287
rect 3553 4273 3567 4287
rect 3273 4213 3287 4227
rect 3213 4193 3227 4207
rect 3253 4193 3267 4207
rect 3293 4193 3307 4207
rect 3413 4213 3427 4227
rect 3413 4193 3427 4207
rect 3233 4153 3247 4167
rect 3393 4113 3407 4127
rect 3193 4093 3207 4107
rect 3193 4033 3207 4047
rect 3433 4173 3447 4187
rect 3953 4453 3967 4467
rect 3993 4473 4007 4487
rect 4033 4473 4047 4487
rect 4133 4473 4147 4487
rect 3993 4433 4007 4447
rect 4053 4453 4067 4467
rect 4053 4433 4067 4447
rect 3893 4413 3907 4427
rect 3833 4293 3847 4307
rect 3733 4253 3747 4267
rect 3473 4213 3487 4227
rect 3473 4173 3487 4187
rect 3433 4153 3447 4167
rect 3453 4153 3467 4167
rect 3093 4013 3107 4027
rect 3053 3993 3067 4007
rect 3013 3953 3027 3967
rect 3033 3973 3047 3987
rect 3073 3973 3087 3987
rect 3053 3953 3067 3967
rect 2993 3853 3007 3867
rect 2993 3833 3007 3847
rect 2973 3793 2987 3807
rect 2973 3773 2987 3787
rect 2773 3693 2787 3707
rect 2793 3713 2807 3727
rect 2913 3713 2927 3727
rect 2953 3713 2967 3727
rect 2813 3673 2827 3687
rect 2853 3673 2867 3687
rect 2753 3613 2767 3627
rect 2813 3613 2827 3627
rect 2753 3553 2767 3567
rect 2773 3533 2787 3547
rect 2793 3533 2807 3547
rect 2633 3513 2647 3527
rect 2633 3493 2647 3507
rect 2673 3493 2687 3507
rect 2733 3493 2747 3507
rect 2773 3493 2787 3507
rect 2673 3473 2687 3487
rect 2653 3313 2667 3327
rect 2653 3253 2667 3267
rect 2633 3233 2647 3247
rect 2653 3233 2667 3247
rect 2653 3193 2667 3207
rect 2633 3113 2647 3127
rect 2753 3473 2767 3487
rect 2733 3433 2747 3447
rect 2753 3253 2767 3267
rect 2893 3553 2907 3567
rect 2853 3533 2867 3547
rect 3033 3733 3047 3747
rect 2993 3693 3007 3707
rect 3013 3693 3027 3707
rect 2973 3673 2987 3687
rect 2973 3653 2987 3667
rect 2953 3593 2967 3607
rect 2933 3573 2947 3587
rect 2913 3533 2927 3547
rect 2813 3513 2827 3527
rect 2833 3513 2847 3527
rect 2873 3513 2887 3527
rect 2853 3453 2867 3467
rect 2833 3393 2847 3407
rect 2813 3353 2827 3367
rect 2693 3233 2707 3247
rect 2713 3213 2727 3227
rect 2733 3233 2747 3247
rect 2793 3233 2807 3247
rect 2673 3173 2687 3187
rect 2713 3173 2727 3187
rect 2733 3173 2747 3187
rect 2673 3093 2687 3107
rect 2653 3073 2667 3087
rect 2693 3073 2707 3087
rect 2813 3213 2827 3227
rect 2773 3173 2787 3187
rect 2973 3573 2987 3587
rect 3013 3673 3027 3687
rect 3053 3713 3067 3727
rect 3053 3673 3067 3687
rect 3033 3653 3047 3667
rect 3013 3613 3027 3627
rect 2973 3533 2987 3547
rect 3013 3533 3027 3547
rect 3033 3533 3047 3547
rect 2953 3493 2967 3507
rect 2913 3473 2927 3487
rect 2993 3513 3007 3527
rect 3013 3493 3027 3507
rect 2973 3473 2987 3487
rect 2993 3453 3007 3467
rect 2893 3413 2907 3427
rect 2873 3273 2887 3287
rect 3173 4013 3187 4027
rect 3213 4013 3227 4027
rect 3233 4013 3247 4027
rect 3273 4013 3287 4027
rect 3313 4013 3327 4027
rect 3113 3973 3127 3987
rect 3153 3993 3167 4007
rect 3113 3933 3127 3947
rect 3173 3933 3187 3947
rect 3193 3933 3207 3947
rect 3093 3893 3107 3907
rect 3093 3753 3107 3767
rect 3253 3973 3267 3987
rect 3353 3993 3367 4007
rect 3333 3973 3347 3987
rect 3373 3973 3387 3987
rect 3413 3993 3427 4007
rect 3413 3973 3427 3987
rect 3233 3873 3247 3887
rect 3193 3733 3207 3747
rect 3113 3713 3127 3727
rect 3153 3713 3167 3727
rect 3173 3713 3187 3727
rect 3233 3713 3247 3727
rect 3253 3713 3267 3727
rect 3173 3693 3187 3707
rect 3113 3673 3127 3687
rect 3093 3613 3107 3627
rect 3093 3573 3107 3587
rect 3133 3653 3147 3667
rect 3173 3653 3187 3667
rect 3153 3593 3167 3607
rect 3173 3593 3187 3607
rect 3213 3553 3227 3567
rect 3233 3553 3247 3567
rect 3133 3493 3147 3507
rect 3213 3513 3227 3527
rect 3253 3513 3267 3527
rect 3033 3433 3047 3447
rect 3193 3453 3207 3467
rect 3113 3433 3127 3447
rect 3093 3373 3107 3387
rect 3053 3293 3067 3307
rect 3013 3273 3027 3287
rect 3033 3273 3047 3287
rect 2913 3233 2927 3247
rect 2893 3213 2907 3227
rect 2853 3193 2867 3207
rect 2833 3173 2847 3187
rect 2793 3153 2807 3167
rect 2833 3133 2847 3147
rect 2753 3113 2767 3127
rect 2753 3053 2767 3067
rect 2773 3053 2787 3067
rect 2673 3013 2687 3027
rect 2713 3033 2727 3047
rect 2733 3033 2747 3047
rect 2713 3013 2727 3027
rect 2813 3033 2827 3047
rect 2833 3033 2847 3047
rect 2633 2913 2647 2927
rect 2613 2793 2627 2807
rect 2553 2773 2567 2787
rect 2573 2773 2587 2787
rect 2453 2613 2467 2627
rect 2313 2553 2327 2567
rect 2353 2553 2367 2567
rect 2393 2393 2407 2407
rect 2313 2293 2327 2307
rect 2353 2333 2367 2347
rect 2353 2293 2367 2307
rect 2433 2553 2447 2567
rect 2373 2253 2387 2267
rect 2313 2193 2327 2207
rect 2773 2993 2787 3007
rect 2813 3013 2827 3027
rect 2833 2993 2847 3007
rect 2713 2813 2727 2827
rect 2893 3033 2907 3047
rect 2973 3233 2987 3247
rect 3113 3333 3127 3347
rect 3153 3333 3167 3347
rect 3113 3273 3127 3287
rect 3053 3233 3067 3247
rect 2933 3193 2947 3207
rect 2953 3193 2967 3207
rect 3013 3193 3027 3207
rect 2993 3073 3007 3087
rect 3013 3073 3027 3087
rect 3073 3213 3087 3227
rect 3053 3153 3067 3167
rect 3053 3133 3067 3147
rect 3033 3053 3047 3067
rect 2873 2993 2887 3007
rect 2893 3013 2907 3027
rect 2793 2853 2807 2867
rect 2813 2813 2827 2827
rect 2753 2793 2767 2807
rect 2773 2793 2787 2807
rect 2853 2953 2867 2967
rect 2893 2973 2907 2987
rect 2913 2973 2927 2987
rect 2913 2873 2927 2887
rect 2973 3013 2987 3027
rect 3013 3013 3027 3027
rect 3033 3033 3047 3047
rect 3173 3293 3187 3307
rect 3333 3953 3347 3967
rect 3373 3953 3387 3967
rect 3293 3933 3307 3947
rect 3293 3873 3307 3887
rect 3293 3713 3307 3727
rect 3393 3933 3407 3947
rect 3413 3933 3427 3947
rect 3373 3733 3387 3747
rect 3413 3893 3427 3907
rect 3373 3693 3387 3707
rect 3393 3713 3407 3727
rect 3413 3693 3427 3707
rect 3373 3673 3387 3687
rect 3313 3613 3327 3627
rect 3353 3613 3367 3627
rect 3313 3573 3327 3587
rect 3333 3573 3347 3587
rect 3413 3653 3427 3667
rect 3413 3633 3427 3647
rect 3393 3593 3407 3607
rect 3373 3553 3387 3567
rect 3333 3533 3347 3547
rect 3353 3513 3367 3527
rect 3393 3513 3407 3527
rect 3413 3513 3427 3527
rect 3293 3373 3307 3387
rect 3273 3333 3287 3347
rect 3293 3333 3307 3347
rect 3233 3313 3247 3327
rect 3333 3373 3347 3387
rect 3553 4213 3567 4227
rect 3613 4213 3627 4227
rect 3513 4153 3527 4167
rect 3493 4113 3507 4127
rect 3473 4073 3487 4087
rect 3533 4133 3547 4147
rect 3533 4113 3547 4127
rect 3513 4013 3527 4027
rect 3593 4093 3607 4107
rect 3553 4073 3567 4087
rect 3473 3993 3487 4007
rect 3453 3953 3467 3967
rect 3453 3913 3467 3927
rect 3513 3913 3527 3927
rect 3573 4013 3587 4027
rect 3653 4193 3667 4207
rect 3633 4173 3647 4187
rect 3693 4193 3707 4207
rect 3673 4153 3687 4167
rect 3653 4133 3667 4147
rect 3633 4113 3647 4127
rect 3613 4033 3627 4047
rect 3633 3993 3647 4007
rect 3593 3953 3607 3967
rect 3573 3913 3587 3927
rect 3553 3753 3567 3767
rect 3793 4213 3807 4227
rect 3753 4193 3767 4207
rect 3733 4173 3747 4187
rect 3813 4173 3827 4187
rect 3773 4153 3787 4167
rect 3693 4133 3707 4147
rect 3993 4273 4007 4287
rect 3933 4233 3947 4247
rect 3873 4193 3887 4207
rect 3913 4153 3927 4167
rect 3893 4133 3907 4147
rect 3853 4073 3867 4087
rect 3753 4033 3767 4047
rect 3833 4033 3847 4047
rect 3673 4013 3687 4027
rect 3713 4013 3727 4027
rect 3673 3993 3687 4007
rect 3713 3973 3727 3987
rect 3733 3973 3747 3987
rect 3633 3953 3647 3967
rect 3653 3953 3667 3967
rect 3613 3913 3627 3927
rect 3593 3753 3607 3767
rect 3453 3733 3467 3747
rect 3473 3713 3487 3727
rect 3493 3733 3507 3747
rect 3533 3733 3547 3747
rect 3573 3733 3587 3747
rect 3493 3693 3507 3707
rect 3473 3613 3487 3627
rect 3493 3513 3507 3527
rect 3393 3493 3407 3507
rect 3433 3493 3447 3507
rect 3413 3473 3427 3487
rect 3493 3473 3507 3487
rect 3393 3453 3407 3467
rect 3453 3453 3467 3467
rect 3413 3433 3427 3447
rect 3493 3433 3507 3447
rect 3533 3573 3547 3587
rect 3553 3553 3567 3567
rect 3693 3893 3707 3907
rect 3633 3733 3647 3747
rect 3633 3693 3647 3707
rect 3653 3713 3667 3727
rect 3693 3713 3707 3727
rect 3673 3673 3687 3687
rect 3673 3653 3687 3667
rect 3613 3533 3627 3547
rect 3633 3533 3647 3547
rect 3553 3493 3567 3507
rect 3593 3493 3607 3507
rect 3473 3413 3487 3427
rect 3513 3413 3527 3427
rect 3393 3353 3407 3367
rect 3433 3353 3447 3367
rect 3453 3353 3467 3367
rect 3393 3313 3407 3327
rect 3373 3293 3387 3307
rect 3353 3273 3367 3287
rect 3193 3253 3207 3267
rect 3213 3253 3227 3267
rect 3153 3233 3167 3247
rect 3173 3233 3187 3247
rect 3213 3233 3227 3247
rect 3273 3253 3287 3267
rect 3253 3233 3267 3247
rect 3153 3193 3167 3207
rect 3173 3193 3187 3207
rect 3093 3113 3107 3127
rect 3073 3093 3087 3107
rect 3053 3013 3067 3027
rect 3073 2993 3087 3007
rect 3153 3153 3167 3167
rect 3213 3153 3227 3167
rect 3173 3113 3187 3127
rect 3193 3093 3207 3107
rect 3213 3093 3227 3107
rect 3173 3073 3187 3087
rect 3153 3033 3167 3047
rect 2973 2973 2987 2987
rect 3093 2973 3107 2987
rect 3013 2953 3027 2967
rect 2933 2853 2947 2867
rect 2913 2833 2927 2847
rect 2953 2833 2967 2847
rect 2773 2773 2787 2787
rect 2593 2753 2607 2767
rect 2613 2733 2627 2747
rect 2693 2753 2707 2767
rect 2733 2753 2747 2767
rect 2793 2753 2807 2767
rect 2833 2773 2847 2787
rect 2853 2773 2867 2787
rect 2833 2753 2847 2767
rect 2893 2773 2907 2787
rect 2753 2733 2767 2747
rect 2553 2693 2567 2707
rect 2573 2693 2587 2707
rect 2653 2693 2667 2707
rect 2713 2693 2727 2707
rect 2513 2673 2527 2687
rect 2553 2673 2567 2687
rect 2653 2673 2667 2687
rect 2673 2673 2687 2687
rect 2713 2673 2727 2687
rect 2513 2653 2527 2667
rect 2653 2633 2667 2647
rect 2613 2593 2627 2607
rect 2513 2573 2527 2587
rect 2573 2573 2587 2587
rect 2513 2533 2527 2547
rect 2553 2533 2567 2547
rect 2453 2453 2467 2467
rect 2453 2413 2467 2427
rect 2533 2373 2547 2387
rect 2513 2353 2527 2367
rect 2673 2573 2687 2587
rect 2593 2533 2607 2547
rect 2633 2533 2647 2547
rect 2693 2533 2707 2547
rect 2613 2413 2627 2427
rect 2573 2393 2587 2407
rect 2493 2333 2507 2347
rect 2593 2333 2607 2347
rect 2873 2713 2887 2727
rect 2873 2693 2887 2707
rect 2933 2733 2947 2747
rect 2973 2733 2987 2747
rect 2913 2713 2927 2727
rect 2833 2653 2847 2667
rect 2893 2653 2907 2667
rect 2893 2633 2907 2647
rect 2853 2613 2867 2627
rect 2813 2593 2827 2607
rect 2753 2513 2767 2527
rect 2773 2533 2787 2547
rect 2773 2453 2787 2467
rect 2753 2413 2767 2427
rect 2713 2373 2727 2387
rect 2673 2333 2687 2347
rect 2653 2313 2667 2327
rect 2553 2293 2567 2307
rect 2533 2273 2547 2287
rect 2573 2273 2587 2287
rect 2633 2233 2647 2247
rect 2493 2213 2507 2227
rect 2473 2113 2487 2127
rect 2313 2093 2327 2107
rect 2393 2093 2407 2107
rect 2353 2073 2367 2087
rect 2333 2053 2347 2067
rect 2373 2033 2387 2047
rect 2313 1913 2327 1927
rect 2453 2073 2467 2087
rect 2433 2033 2447 2047
rect 2653 2173 2667 2187
rect 2613 2113 2627 2127
rect 2573 2093 2587 2107
rect 2473 2033 2487 2047
rect 2493 2033 2507 2047
rect 2513 2033 2527 2047
rect 2533 2053 2547 2067
rect 2433 1973 2447 1987
rect 2413 1873 2427 1887
rect 2493 1873 2507 1887
rect 2033 1793 2047 1807
rect 2093 1793 2107 1807
rect 1933 1673 1947 1687
rect 1973 1673 1987 1687
rect 1913 1653 1927 1667
rect 1913 1633 1927 1647
rect 1593 1513 1607 1527
rect 1533 1373 1547 1387
rect 1493 1313 1507 1327
rect 1573 1293 1587 1307
rect 1453 893 1467 907
rect 1493 873 1507 887
rect 1433 813 1447 827
rect 1473 793 1487 807
rect 1433 733 1447 747
rect 1373 713 1387 727
rect 1333 693 1347 707
rect 1313 673 1327 687
rect 1293 653 1307 667
rect 1173 633 1187 647
rect 1173 613 1187 627
rect 1213 613 1227 627
rect 1273 633 1287 647
rect 1353 673 1367 687
rect 1393 693 1407 707
rect 1553 1253 1567 1267
rect 1553 1113 1567 1127
rect 1653 1373 1667 1387
rect 1653 1353 1667 1367
rect 1793 1553 1807 1567
rect 1673 1313 1687 1327
rect 1713 1333 1727 1347
rect 1613 1293 1627 1307
rect 1633 1133 1647 1147
rect 1673 1133 1687 1147
rect 1613 1093 1627 1107
rect 1653 1073 1667 1087
rect 1693 1073 1707 1087
rect 1593 1053 1607 1067
rect 1573 1033 1587 1047
rect 1553 913 1567 927
rect 1613 873 1627 887
rect 1533 793 1547 807
rect 1653 853 1667 867
rect 1593 793 1607 807
rect 1633 793 1647 807
rect 1593 773 1607 787
rect 1653 753 1667 767
rect 1513 633 1527 647
rect 1573 673 1587 687
rect 1633 653 1647 667
rect 1593 633 1607 647
rect 1193 393 1207 407
rect 1373 393 1387 407
rect 1493 393 1507 407
rect 1593 393 1607 407
rect 933 353 947 367
rect 953 333 967 347
rect 993 353 1007 367
rect 1093 373 1107 387
rect 1113 373 1127 387
rect 1133 373 1147 387
rect 1013 333 1027 347
rect 953 313 967 327
rect 813 153 827 167
rect 773 93 787 107
rect 813 113 827 127
rect 1093 333 1107 347
rect 1053 293 1067 307
rect 1013 273 1027 287
rect 1333 373 1347 387
rect 1133 333 1147 347
rect 1153 353 1167 367
rect 1233 353 1247 367
rect 1313 333 1327 347
rect 1693 753 1707 767
rect 1673 693 1687 707
rect 1753 1313 1767 1327
rect 1793 1313 1807 1327
rect 1813 1293 1827 1307
rect 1733 1213 1747 1227
rect 1813 1273 1827 1287
rect 1953 1613 1967 1627
rect 1933 1573 1947 1587
rect 1913 1553 1927 1567
rect 1853 1293 1867 1307
rect 1833 1253 1847 1267
rect 1893 1293 1907 1307
rect 2093 1733 2107 1747
rect 2213 1793 2227 1807
rect 2293 1793 2307 1807
rect 2233 1773 2247 1787
rect 2133 1753 2147 1767
rect 2153 1753 2167 1767
rect 2273 1753 2287 1767
rect 2053 1713 2067 1727
rect 2113 1713 2127 1727
rect 2033 1653 2047 1667
rect 1973 1293 1987 1307
rect 1893 1213 1907 1227
rect 1773 1193 1787 1207
rect 1893 1193 1907 1207
rect 1753 1153 1767 1167
rect 1733 1113 1747 1127
rect 1793 1073 1807 1087
rect 1733 1053 1747 1067
rect 1753 1033 1767 1047
rect 1913 1133 1927 1147
rect 1833 693 1847 707
rect 1773 653 1787 667
rect 1113 233 1127 247
rect 1153 233 1167 247
rect 1133 173 1147 187
rect 1033 153 1047 167
rect 1053 133 1067 147
rect 1173 193 1187 207
rect 1293 313 1307 327
rect 1213 293 1227 307
rect 1193 173 1207 187
rect 1453 333 1467 347
rect 1473 353 1487 367
rect 1513 353 1527 367
rect 1553 373 1567 387
rect 1573 353 1587 367
rect 1653 373 1667 387
rect 1493 333 1507 347
rect 1413 313 1427 327
rect 1353 293 1367 307
rect 1253 273 1267 287
rect 1333 213 1347 227
rect 1373 213 1387 227
rect 1233 193 1247 207
rect 1153 133 1167 147
rect 1213 153 1227 167
rect 1273 173 1287 187
rect 1733 373 1747 387
rect 1793 633 1807 647
rect 1973 1273 1987 1287
rect 2013 1113 2027 1127
rect 1933 913 1947 927
rect 1973 913 1987 927
rect 2053 1613 2067 1627
rect 2133 1593 2147 1607
rect 2213 1733 2227 1747
rect 2433 1813 2447 1827
rect 2393 1793 2407 1807
rect 2373 1753 2387 1767
rect 2413 1773 2427 1787
rect 2193 1713 2207 1727
rect 2393 1733 2407 1747
rect 2293 1613 2307 1627
rect 2393 1613 2407 1627
rect 2233 1593 2247 1607
rect 2253 1593 2267 1607
rect 2153 1553 2167 1567
rect 2333 1593 2347 1607
rect 2273 1553 2287 1567
rect 2373 1593 2387 1607
rect 2313 1553 2327 1567
rect 2353 1433 2367 1447
rect 2393 1433 2407 1447
rect 2293 1373 2307 1387
rect 2313 1373 2327 1387
rect 2053 1313 2067 1327
rect 2093 1313 2107 1327
rect 2153 1313 2167 1327
rect 2193 1313 2207 1327
rect 2273 1313 2287 1327
rect 2433 1353 2447 1367
rect 2553 1993 2567 2007
rect 2533 1813 2547 1827
rect 2513 1773 2527 1787
rect 2733 2313 2747 2327
rect 2693 2293 2707 2307
rect 2713 2273 2727 2287
rect 2753 2173 2767 2187
rect 2673 2093 2687 2107
rect 2753 2093 2767 2107
rect 2593 2073 2607 2087
rect 2713 2073 2727 2087
rect 2693 2053 2707 2067
rect 2753 2013 2767 2027
rect 2673 1993 2687 2007
rect 2733 1993 2747 2007
rect 2633 1973 2647 1987
rect 2673 1953 2687 1967
rect 2593 1773 2607 1787
rect 2633 1773 2647 1787
rect 2633 1753 2647 1767
rect 2573 1713 2587 1727
rect 2593 1673 2607 1687
rect 2493 1393 2507 1407
rect 2453 1333 2467 1347
rect 2173 1293 2187 1307
rect 2133 1273 2147 1287
rect 2073 1213 2087 1227
rect 2453 1293 2467 1307
rect 2493 1293 2507 1307
rect 2433 1253 2447 1267
rect 2353 1173 2367 1187
rect 2153 1153 2167 1167
rect 2313 1153 2327 1167
rect 2333 1153 2347 1167
rect 2133 1133 2147 1147
rect 2053 1093 2067 1107
rect 2073 1093 2087 1107
rect 2113 1113 2127 1127
rect 2173 1133 2187 1147
rect 2213 1133 2227 1147
rect 2153 893 2167 907
rect 2033 873 2047 887
rect 1993 853 2007 867
rect 1913 813 1927 827
rect 1933 733 1947 747
rect 1873 673 1887 687
rect 1893 673 1907 687
rect 1853 653 1867 667
rect 2053 813 2067 827
rect 2093 833 2107 847
rect 2113 813 2127 827
rect 2033 793 2047 807
rect 2093 793 2107 807
rect 1993 773 2007 787
rect 2073 773 2087 787
rect 1953 693 1967 707
rect 1973 653 1987 667
rect 1913 633 1927 647
rect 2193 1113 2207 1127
rect 2253 1093 2267 1107
rect 2293 1093 2307 1107
rect 2293 1073 2307 1087
rect 2473 1233 2487 1247
rect 2533 1613 2547 1627
rect 2573 1593 2587 1607
rect 2593 1533 2607 1547
rect 2593 1513 2607 1527
rect 2633 1613 2647 1627
rect 2653 1613 2667 1627
rect 2553 1293 2567 1307
rect 2513 1273 2527 1287
rect 2493 1213 2507 1227
rect 2573 1213 2587 1227
rect 2493 1193 2507 1207
rect 2473 1113 2487 1127
rect 2253 913 2267 927
rect 2373 913 2387 927
rect 2173 853 2187 867
rect 2153 813 2167 827
rect 2193 833 2207 847
rect 2233 833 2247 847
rect 2233 813 2247 827
rect 2413 873 2427 887
rect 2553 1173 2567 1187
rect 2733 1693 2747 1707
rect 2693 1573 2707 1587
rect 2673 1453 2687 1467
rect 2793 2333 2807 2347
rect 2993 2693 3007 2707
rect 2933 2593 2947 2607
rect 3153 2953 3167 2967
rect 3113 2853 3127 2867
rect 3093 2793 3107 2807
rect 3133 2833 3147 2847
rect 3193 2913 3207 2927
rect 3213 2913 3227 2927
rect 3193 2833 3207 2847
rect 3133 2793 3147 2807
rect 3153 2793 3167 2807
rect 3193 2793 3207 2807
rect 3053 2753 3067 2767
rect 3093 2753 3107 2767
rect 3093 2733 3107 2747
rect 3153 2753 3167 2767
rect 3173 2773 3187 2787
rect 3153 2733 3167 2747
rect 3173 2733 3187 2747
rect 3053 2693 3067 2707
rect 3073 2693 3087 2707
rect 3033 2673 3047 2687
rect 3053 2613 3067 2627
rect 2833 2533 2847 2547
rect 2913 2553 2927 2567
rect 2873 2513 2887 2527
rect 2973 2553 2987 2567
rect 2973 2513 2987 2527
rect 2953 2433 2967 2447
rect 2833 2313 2847 2327
rect 2933 2313 2947 2327
rect 2813 2293 2827 2307
rect 2793 2273 2807 2287
rect 2853 2253 2867 2267
rect 2913 2253 2927 2267
rect 2873 2233 2887 2247
rect 2893 2233 2907 2247
rect 2933 2213 2947 2227
rect 2893 2193 2907 2207
rect 2913 2173 2927 2187
rect 2853 2073 2867 2087
rect 2853 1833 2867 1847
rect 2833 1813 2847 1827
rect 2813 1713 2827 1727
rect 2793 1633 2807 1647
rect 2873 1773 2887 1787
rect 2893 1693 2907 1707
rect 2873 1633 2887 1647
rect 2873 1593 2887 1607
rect 3013 2573 3027 2587
rect 3033 2533 3047 2547
rect 3073 2553 3087 2567
rect 3133 2713 3147 2727
rect 3093 2533 3107 2547
rect 2993 2493 3007 2507
rect 3033 2493 3047 2507
rect 2993 2293 3007 2307
rect 2953 2193 2967 2207
rect 2973 2193 2987 2207
rect 2973 2073 2987 2087
rect 2933 1953 2947 1967
rect 3013 2113 3027 2127
rect 3013 2073 3027 2087
rect 3013 2033 3027 2047
rect 3073 2333 3087 2347
rect 3133 2553 3147 2567
rect 3173 2693 3187 2707
rect 3193 2573 3207 2587
rect 3193 2553 3207 2567
rect 3133 2513 3147 2527
rect 3113 2473 3127 2487
rect 3173 2473 3187 2487
rect 3113 2433 3127 2447
rect 3093 2293 3107 2307
rect 3053 2253 3067 2267
rect 3073 2253 3087 2267
rect 3093 2233 3107 2247
rect 3313 3253 3327 3267
rect 3413 3273 3427 3287
rect 3293 3193 3307 3207
rect 3273 3133 3287 3147
rect 3253 3013 3267 3027
rect 3273 3033 3287 3047
rect 3253 2933 3267 2947
rect 3273 2893 3287 2907
rect 3233 2793 3247 2807
rect 3333 3233 3347 3247
rect 3353 3213 3367 3227
rect 3453 3293 3467 3307
rect 3433 3253 3447 3267
rect 3413 3193 3427 3207
rect 3373 3153 3387 3167
rect 3313 3113 3327 3127
rect 3333 3113 3347 3127
rect 3573 3453 3587 3467
rect 3553 3393 3567 3407
rect 3493 3313 3507 3327
rect 3553 3293 3567 3307
rect 3513 3273 3527 3287
rect 3493 3253 3507 3267
rect 3533 3233 3547 3247
rect 3593 3413 3607 3427
rect 3573 3233 3587 3247
rect 3493 3213 3507 3227
rect 3573 3213 3587 3227
rect 3453 3173 3467 3187
rect 3473 3173 3487 3187
rect 3433 3113 3447 3127
rect 3433 3073 3447 3087
rect 3413 3053 3427 3067
rect 3313 2993 3327 3007
rect 3373 2993 3387 3007
rect 3353 2953 3367 2967
rect 3313 2873 3327 2887
rect 3373 2853 3387 2867
rect 3473 3073 3487 3087
rect 3533 3133 3547 3147
rect 3553 3053 3567 3067
rect 3653 3413 3667 3427
rect 3653 3393 3667 3407
rect 3613 3373 3627 3387
rect 3653 3333 3667 3347
rect 3633 3293 3647 3307
rect 3613 3253 3627 3267
rect 3613 3213 3627 3227
rect 3733 3913 3747 3927
rect 3793 3993 3807 4007
rect 3773 3953 3787 3967
rect 3813 3973 3827 3987
rect 3793 3913 3807 3927
rect 3873 3953 3887 3967
rect 3893 3973 3907 3987
rect 4113 4433 4127 4447
rect 4393 4513 4407 4527
rect 4433 4493 4447 4507
rect 4173 4453 4187 4467
rect 4193 4453 4207 4467
rect 4273 4453 4287 4467
rect 4153 4433 4167 4447
rect 4113 4413 4127 4427
rect 4093 4373 4107 4387
rect 4093 4353 4107 4367
rect 4013 4233 4027 4247
rect 3973 4193 3987 4207
rect 4053 4193 4067 4207
rect 3953 4153 3967 4167
rect 4073 4153 4087 4167
rect 4033 4093 4047 4107
rect 4073 4093 4087 4107
rect 4033 4033 4047 4047
rect 3973 3973 3987 3987
rect 3953 3933 3967 3947
rect 3813 3893 3827 3907
rect 3853 3893 3867 3907
rect 3913 3893 3927 3907
rect 3753 3753 3767 3767
rect 3733 3733 3747 3747
rect 3753 3713 3767 3727
rect 3773 3713 3787 3727
rect 3713 3613 3727 3627
rect 3773 3693 3787 3707
rect 3793 3693 3807 3707
rect 3833 3713 3847 3727
rect 3873 3713 3887 3727
rect 3913 3713 3927 3727
rect 3793 3673 3807 3687
rect 3813 3673 3827 3687
rect 3853 3673 3867 3687
rect 3933 3693 3947 3707
rect 3893 3673 3907 3687
rect 3913 3673 3927 3687
rect 3773 3653 3787 3667
rect 3753 3573 3767 3587
rect 3713 3553 3727 3567
rect 3753 3513 3767 3527
rect 3733 3473 3747 3487
rect 3673 3253 3687 3267
rect 3593 3133 3607 3147
rect 3613 3093 3627 3107
rect 3433 2873 3447 2887
rect 3433 2833 3447 2847
rect 3453 2833 3467 2847
rect 3293 2813 3307 2827
rect 3313 2813 3327 2827
rect 3393 2813 3407 2827
rect 3233 2753 3247 2767
rect 3253 2693 3267 2707
rect 3273 2673 3287 2687
rect 3293 2653 3307 2667
rect 3293 2593 3307 2607
rect 3273 2573 3287 2587
rect 3233 2513 3247 2527
rect 3213 2453 3227 2467
rect 3233 2433 3247 2447
rect 3253 2433 3267 2447
rect 3173 2393 3187 2407
rect 3193 2373 3207 2387
rect 3133 2293 3147 2307
rect 3113 2213 3127 2227
rect 3133 2213 3147 2227
rect 3173 2293 3187 2307
rect 3333 2773 3347 2787
rect 3353 2753 3367 2767
rect 3393 2673 3407 2687
rect 3333 2633 3347 2647
rect 3293 2553 3307 2567
rect 3313 2553 3327 2567
rect 3353 2613 3367 2627
rect 3313 2513 3327 2527
rect 3433 2753 3447 2767
rect 3493 2993 3507 3007
rect 3493 2933 3507 2947
rect 3513 2933 3527 2947
rect 3513 2853 3527 2867
rect 3513 2813 3527 2827
rect 3493 2793 3507 2807
rect 3433 2733 3447 2747
rect 3473 2733 3487 2747
rect 3413 2573 3427 2587
rect 3413 2533 3427 2547
rect 3573 3033 3587 3047
rect 3573 2993 3587 3007
rect 3593 3013 3607 3027
rect 3733 3393 3747 3407
rect 3813 3633 3827 3647
rect 4073 3933 4087 3947
rect 4053 3893 4067 3907
rect 4013 3873 4027 3887
rect 4233 4433 4247 4447
rect 4233 4413 4247 4427
rect 4213 4393 4227 4407
rect 4133 4273 4147 4287
rect 4193 4273 4207 4287
rect 4313 4453 4327 4467
rect 4453 4453 4467 4467
rect 4553 4493 4567 4507
rect 4413 4433 4427 4447
rect 4393 4413 4407 4427
rect 4293 4393 4307 4407
rect 4333 4393 4347 4407
rect 4293 4253 4307 4267
rect 4213 4233 4227 4247
rect 4273 4233 4287 4247
rect 4133 4173 4147 4187
rect 4113 4053 4127 4067
rect 4193 4193 4207 4207
rect 4233 4213 4247 4227
rect 4273 4213 4287 4227
rect 4193 4173 4207 4187
rect 4153 4153 4167 4167
rect 4173 4153 4187 4167
rect 4153 4113 4167 4127
rect 4133 4033 4147 4047
rect 4173 4013 4187 4027
rect 4133 3993 4147 4007
rect 4113 3953 4127 3967
rect 4133 3973 4147 3987
rect 4173 3973 4187 3987
rect 4153 3953 4167 3967
rect 4133 3933 4147 3947
rect 4093 3813 4107 3827
rect 4153 3833 4167 3847
rect 4133 3793 4147 3807
rect 3973 3713 3987 3727
rect 3813 3613 3827 3627
rect 3853 3613 3867 3627
rect 3793 3513 3807 3527
rect 3853 3553 3867 3567
rect 3953 3653 3967 3667
rect 3953 3633 3967 3647
rect 3913 3513 3927 3527
rect 3993 3693 4007 3707
rect 4033 3713 4047 3727
rect 4093 3713 4107 3727
rect 4113 3693 4127 3707
rect 4053 3673 4067 3687
rect 4013 3653 4027 3667
rect 3993 3593 4007 3607
rect 3793 3413 3807 3427
rect 3753 3333 3767 3347
rect 3773 3293 3787 3307
rect 3733 3273 3747 3287
rect 3933 3473 3947 3487
rect 3893 3333 3907 3347
rect 3853 3273 3867 3287
rect 3913 3313 3927 3327
rect 3793 3253 3807 3267
rect 3753 3213 3767 3227
rect 3773 3233 3787 3247
rect 3813 3233 3827 3247
rect 3853 3233 3867 3247
rect 3873 3253 3887 3267
rect 3893 3253 3907 3267
rect 4033 3573 4047 3587
rect 4033 3553 4047 3567
rect 4053 3513 4067 3527
rect 4013 3413 4027 3427
rect 3993 3393 4007 3407
rect 4093 3613 4107 3627
rect 4173 3793 4187 3807
rect 4253 4173 4267 4187
rect 4273 4173 4287 4187
rect 4213 4133 4227 4147
rect 4233 4133 4247 4147
rect 4233 4053 4247 4067
rect 4273 4153 4287 4167
rect 4313 4193 4327 4207
rect 4353 4193 4367 4207
rect 4373 4173 4387 4187
rect 4513 4433 4527 4447
rect 4573 4453 4587 4467
rect 4553 4433 4567 4447
rect 4493 4413 4507 4427
rect 4533 4413 4547 4427
rect 4453 4333 4467 4347
rect 4493 4333 4507 4347
rect 4413 4253 4427 4267
rect 4433 4193 4447 4207
rect 4473 4193 4487 4207
rect 4293 4093 4307 4107
rect 4353 4113 4367 4127
rect 4333 4093 4347 4107
rect 4313 4033 4327 4047
rect 4253 4013 4267 4027
rect 4273 4013 4287 4027
rect 4253 3973 4267 3987
rect 4273 3993 4287 4007
rect 4293 3993 4307 4007
rect 4313 3973 4327 3987
rect 4393 4013 4407 4027
rect 4593 4373 4607 4387
rect 4533 4213 4547 4227
rect 4593 4213 4607 4227
rect 4513 4173 4527 4187
rect 4533 4193 4547 4207
rect 4573 4193 4587 4207
rect 4533 4153 4547 4167
rect 4513 4133 4527 4147
rect 4493 4093 4507 4107
rect 4253 3953 4267 3967
rect 4213 3933 4227 3947
rect 4173 3713 4187 3727
rect 4193 3713 4207 3727
rect 4213 3713 4227 3727
rect 4313 3733 4327 3747
rect 4453 3993 4467 4007
rect 4413 3973 4427 3987
rect 4493 3973 4507 3987
rect 4593 4153 4607 4167
rect 4553 4113 4567 4127
rect 4673 4453 4687 4467
rect 4653 4433 4667 4447
rect 4713 4453 4727 4467
rect 4753 4433 4767 4447
rect 4733 4393 4747 4407
rect 4713 4353 4727 4367
rect 4693 4213 4707 4227
rect 4633 4193 4647 4207
rect 4633 4133 4647 4147
rect 4653 4113 4667 4127
rect 4553 4093 4567 4107
rect 4613 4093 4627 4107
rect 4533 3973 4547 3987
rect 4513 3953 4527 3967
rect 4453 3913 4467 3927
rect 4393 3853 4407 3867
rect 4433 3853 4447 3867
rect 4393 3733 4407 3747
rect 4273 3713 4287 3727
rect 4253 3693 4267 3707
rect 4153 3673 4167 3687
rect 4173 3673 4187 3687
rect 4233 3673 4247 3687
rect 4153 3553 4167 3567
rect 4133 3533 4147 3547
rect 4073 3433 4087 3447
rect 4073 3413 4087 3427
rect 3973 3373 3987 3387
rect 4053 3373 4067 3387
rect 4053 3333 4067 3347
rect 4033 3293 4047 3307
rect 3993 3273 4007 3287
rect 3933 3253 3947 3267
rect 3673 3193 3687 3207
rect 3693 3193 3707 3207
rect 3713 3193 3727 3207
rect 3793 3193 3807 3207
rect 3833 3213 3847 3227
rect 3873 3213 3887 3227
rect 3953 3233 3967 3247
rect 4013 3233 4027 3247
rect 4053 3253 4067 3267
rect 3933 3213 3947 3227
rect 3973 3213 3987 3227
rect 3773 3153 3787 3167
rect 3813 3153 3827 3167
rect 3713 3133 3727 3147
rect 3653 3113 3667 3127
rect 3693 3093 3707 3107
rect 3673 3013 3687 3027
rect 3753 3113 3767 3127
rect 3633 2993 3647 3007
rect 3673 2993 3687 3007
rect 3613 2953 3627 2967
rect 3553 2893 3567 2907
rect 3553 2813 3567 2827
rect 3533 2773 3547 2787
rect 3613 2753 3627 2767
rect 3653 2753 3667 2767
rect 3713 2953 3727 2967
rect 3833 3093 3847 3107
rect 3893 3173 3907 3187
rect 3873 3073 3887 3087
rect 3813 3053 3827 3067
rect 3793 3033 3807 3047
rect 3753 2973 3767 2987
rect 3833 3033 3847 3047
rect 3873 3033 3887 3047
rect 3933 3033 3947 3047
rect 3973 3193 3987 3207
rect 4013 3193 4027 3207
rect 4133 3473 4147 3487
rect 4113 3453 4127 3467
rect 4093 3333 4107 3347
rect 4193 3633 4207 3647
rect 4253 3633 4267 3647
rect 4213 3613 4227 3627
rect 4193 3533 4207 3547
rect 4173 3453 4187 3467
rect 4153 3433 4167 3447
rect 4133 3333 4147 3347
rect 4113 3253 4127 3267
rect 4113 3213 4127 3227
rect 4033 3053 4047 3067
rect 4013 3033 4027 3047
rect 3813 2993 3827 3007
rect 3813 2953 3827 2967
rect 3793 2933 3807 2947
rect 3753 2893 3767 2907
rect 3733 2833 3747 2847
rect 3773 2833 3787 2847
rect 3693 2753 3707 2767
rect 3753 2773 3767 2787
rect 3493 2673 3507 2687
rect 3533 2653 3547 2667
rect 3473 2633 3487 2647
rect 3613 2713 3627 2727
rect 3633 2673 3647 2687
rect 3613 2613 3627 2627
rect 3573 2593 3587 2607
rect 3593 2593 3607 2607
rect 3513 2573 3527 2587
rect 3433 2513 3447 2527
rect 3353 2353 3367 2367
rect 3313 2333 3327 2347
rect 3293 2313 3307 2327
rect 3253 2293 3267 2307
rect 3193 2273 3207 2287
rect 3213 2253 3227 2267
rect 3233 2273 3247 2287
rect 3273 2273 3287 2287
rect 3193 2233 3207 2247
rect 3273 2233 3287 2247
rect 2993 1893 3007 1907
rect 3013 1873 3027 1887
rect 3173 2093 3187 2107
rect 3193 2093 3207 2107
rect 3333 2273 3347 2287
rect 3453 2393 3467 2407
rect 3393 2353 3407 2367
rect 3613 2573 3627 2587
rect 3533 2553 3547 2567
rect 3613 2553 3627 2567
rect 3633 2553 3647 2567
rect 3533 2513 3547 2527
rect 3613 2513 3627 2527
rect 3513 2473 3527 2487
rect 3573 2493 3587 2507
rect 3593 2493 3607 2507
rect 3533 2413 3547 2427
rect 3373 2273 3387 2287
rect 3413 2273 3427 2287
rect 3433 2293 3447 2307
rect 3453 2293 3467 2307
rect 3493 2293 3507 2307
rect 3613 2393 3627 2407
rect 3333 2193 3347 2207
rect 3373 2193 3387 2207
rect 3453 2193 3467 2207
rect 3473 2193 3487 2207
rect 3333 2133 3347 2147
rect 3293 2113 3307 2127
rect 3413 2113 3427 2127
rect 3393 2093 3407 2107
rect 3153 2073 3167 2087
rect 3253 2073 3267 2087
rect 3113 2033 3127 2047
rect 3173 2033 3187 2047
rect 3093 2013 3107 2027
rect 3213 2013 3227 2027
rect 3113 1973 3127 1987
rect 3153 1973 3167 1987
rect 3073 1953 3087 1967
rect 3053 1853 3067 1867
rect 3053 1833 3067 1847
rect 2953 1773 2967 1787
rect 3033 1813 3047 1827
rect 2953 1633 2967 1647
rect 2933 1593 2947 1607
rect 2913 1553 2927 1567
rect 2833 1513 2847 1527
rect 2893 1533 2907 1547
rect 2813 1493 2827 1507
rect 2773 1473 2787 1487
rect 2853 1473 2867 1487
rect 2893 1473 2907 1487
rect 2693 1293 2707 1307
rect 2633 1253 2647 1267
rect 2593 1173 2607 1187
rect 2613 1153 2627 1167
rect 2753 1353 2767 1367
rect 2833 1353 2847 1367
rect 2773 1293 2787 1307
rect 2933 1353 2947 1367
rect 2973 1553 2987 1567
rect 2993 1573 3007 1587
rect 3033 1573 3047 1587
rect 2993 1533 3007 1547
rect 3013 1533 3027 1547
rect 3013 1513 3027 1527
rect 3013 1453 3027 1467
rect 2993 1413 3007 1427
rect 2953 1333 2967 1347
rect 3173 1953 3187 1967
rect 3193 1893 3207 1907
rect 3093 1793 3107 1807
rect 3113 1813 3127 1827
rect 3073 1773 3087 1787
rect 3093 1753 3107 1767
rect 3073 1673 3087 1687
rect 3093 1633 3107 1647
rect 3153 1813 3167 1827
rect 3233 1833 3247 1847
rect 3293 2033 3307 2047
rect 3333 2053 3347 2067
rect 3373 2053 3387 2067
rect 3353 2033 3367 2047
rect 3313 2013 3327 2027
rect 3293 1953 3307 1967
rect 3273 1853 3287 1867
rect 3253 1813 3267 1827
rect 3153 1773 3167 1787
rect 3213 1793 3227 1807
rect 3233 1753 3247 1767
rect 3213 1733 3227 1747
rect 3153 1713 3167 1727
rect 3233 1673 3247 1687
rect 3213 1653 3227 1667
rect 3253 1653 3267 1667
rect 3193 1633 3207 1647
rect 3133 1613 3147 1627
rect 3133 1593 3147 1607
rect 3173 1593 3187 1607
rect 3113 1553 3127 1567
rect 3053 1513 3067 1527
rect 3093 1513 3107 1527
rect 3073 1453 3087 1467
rect 3033 1373 3047 1387
rect 3033 1353 3047 1367
rect 2973 1313 2987 1327
rect 2753 1173 2767 1187
rect 2813 1153 2827 1167
rect 2793 1133 2807 1147
rect 2653 1093 2667 1107
rect 2353 853 2367 867
rect 2293 833 2307 847
rect 2333 833 2347 847
rect 2133 773 2147 787
rect 2133 753 2147 767
rect 2093 733 2107 747
rect 2053 713 2067 727
rect 2073 673 2087 687
rect 2093 673 2107 687
rect 1953 613 1967 627
rect 2053 633 2067 647
rect 1913 593 1927 607
rect 1773 333 1787 347
rect 1753 313 1767 327
rect 1613 273 1627 287
rect 1513 213 1527 227
rect 1493 193 1507 207
rect 1393 173 1407 187
rect 1433 173 1447 187
rect 1153 113 1167 127
rect 1413 133 1427 147
rect 1553 193 1567 207
rect 1533 173 1547 187
rect 1693 233 1707 247
rect 1653 193 1667 207
rect 1633 133 1647 147
rect 1693 153 1707 167
rect 1673 133 1687 147
rect 1353 113 1367 127
rect 1393 113 1407 127
rect 1673 113 1687 127
rect 973 93 987 107
rect 1293 93 1307 107
rect 1473 93 1487 107
rect 1893 373 1907 387
rect 1933 373 1947 387
rect 2053 373 2067 387
rect 1753 153 1767 167
rect 1813 153 1827 167
rect 1793 113 1807 127
rect 1893 153 1907 167
rect 1993 333 2007 347
rect 2013 353 2027 367
rect 2213 773 2227 787
rect 2173 713 2187 727
rect 2273 773 2287 787
rect 2313 773 2327 787
rect 2153 633 2167 647
rect 2233 673 2247 687
rect 2133 373 2147 387
rect 2133 333 2147 347
rect 2393 833 2407 847
rect 2493 853 2507 867
rect 2413 773 2427 787
rect 2373 733 2387 747
rect 2373 653 2387 667
rect 2753 1093 2767 1107
rect 2773 1113 2787 1127
rect 2713 1073 2727 1087
rect 2653 913 2667 927
rect 2533 693 2547 707
rect 2573 693 2587 707
rect 2493 673 2507 687
rect 2453 653 2467 667
rect 2433 613 2447 627
rect 2473 613 2487 627
rect 2513 613 2527 627
rect 2353 433 2367 447
rect 2553 673 2567 687
rect 2573 653 2587 667
rect 2653 773 2667 787
rect 2713 873 2727 887
rect 2713 773 2727 787
rect 2653 693 2667 707
rect 2653 673 2667 687
rect 2773 1073 2787 1087
rect 2773 873 2787 887
rect 2873 1273 2887 1287
rect 2913 1253 2927 1267
rect 2893 1173 2907 1187
rect 2873 1153 2887 1167
rect 2853 1113 2867 1127
rect 2933 1133 2947 1147
rect 2893 1113 2907 1127
rect 2913 1113 2927 1127
rect 2873 1093 2887 1107
rect 2833 993 2847 1007
rect 2793 853 2807 867
rect 2813 853 2827 867
rect 3013 1273 3027 1287
rect 2993 1193 3007 1207
rect 3073 1273 3087 1287
rect 3053 1173 3067 1187
rect 3073 1153 3087 1167
rect 2973 1133 2987 1147
rect 3033 1133 3047 1147
rect 2953 1113 2967 1127
rect 2973 1113 2987 1127
rect 3013 1113 3027 1127
rect 2973 1093 2987 1107
rect 3033 1093 3047 1107
rect 3013 1073 3027 1087
rect 2913 1053 2927 1067
rect 2913 933 2927 947
rect 2933 853 2947 867
rect 2793 813 2807 827
rect 2833 793 2847 807
rect 2793 753 2807 767
rect 2833 673 2847 687
rect 2693 653 2707 667
rect 2713 653 2727 667
rect 2733 653 2747 667
rect 2753 653 2767 667
rect 2613 633 2627 647
rect 2533 453 2547 467
rect 2393 393 2407 407
rect 2513 393 2527 407
rect 2173 313 2187 327
rect 2213 313 2227 327
rect 2213 293 2227 307
rect 2313 353 2327 367
rect 2353 333 2367 347
rect 2413 353 2427 367
rect 2453 353 2467 367
rect 2533 353 2547 367
rect 2553 373 2567 387
rect 2273 313 2287 327
rect 2333 313 2347 327
rect 2413 313 2427 327
rect 2273 233 2287 247
rect 2113 213 2127 227
rect 2273 213 2287 227
rect 2193 193 2207 207
rect 2233 193 2247 207
rect 2033 173 2047 187
rect 2093 173 2107 187
rect 1953 133 1967 147
rect 2213 173 2227 187
rect 2133 153 2147 167
rect 2293 193 2307 207
rect 2313 193 2327 207
rect 1933 113 1947 127
rect 2233 153 2247 167
rect 2373 213 2387 227
rect 2753 613 2767 627
rect 2773 613 2787 627
rect 2813 613 2827 627
rect 2733 553 2747 567
rect 2913 833 2927 847
rect 2893 793 2907 807
rect 2993 1033 3007 1047
rect 3053 1053 3067 1067
rect 3153 1493 3167 1507
rect 3193 1413 3207 1427
rect 3133 1373 3147 1387
rect 3113 1293 3127 1307
rect 3133 1313 3147 1327
rect 3253 1633 3267 1647
rect 3553 2233 3567 2247
rect 3573 2233 3587 2247
rect 3593 2233 3607 2247
rect 3533 2113 3547 2127
rect 3473 2093 3487 2107
rect 3493 2093 3507 2107
rect 3413 2073 3427 2087
rect 3433 2073 3447 2087
rect 3413 2053 3427 2067
rect 3513 2073 3527 2087
rect 3433 2033 3447 2047
rect 3393 1993 3407 2007
rect 3373 1973 3387 1987
rect 3353 1833 3367 1847
rect 3373 1833 3387 1847
rect 3293 1773 3307 1787
rect 3313 1653 3327 1667
rect 3293 1633 3307 1647
rect 3313 1633 3327 1647
rect 3273 1593 3287 1607
rect 3233 1553 3247 1567
rect 3273 1553 3287 1567
rect 3273 1533 3287 1547
rect 3273 1473 3287 1487
rect 3253 1453 3267 1467
rect 3313 1593 3327 1607
rect 3293 1433 3307 1447
rect 3213 1293 3227 1307
rect 3153 1273 3167 1287
rect 3173 1153 3187 1167
rect 3213 1153 3227 1167
rect 3153 1133 3167 1147
rect 3213 1133 3227 1147
rect 3273 1333 3287 1347
rect 3413 1813 3427 1827
rect 3593 2153 3607 2167
rect 3573 2113 3587 2127
rect 3553 2073 3567 2087
rect 3713 2733 3727 2747
rect 3693 2693 3707 2707
rect 3673 2613 3687 2627
rect 3673 2573 3687 2587
rect 3653 2333 3667 2347
rect 3673 2333 3687 2347
rect 3653 2313 3667 2327
rect 3633 2253 3647 2267
rect 3633 2193 3647 2207
rect 3593 2093 3607 2107
rect 3613 2093 3627 2107
rect 3713 2653 3727 2667
rect 3733 2613 3747 2627
rect 3713 2573 3727 2587
rect 3753 2573 3767 2587
rect 3753 2553 3767 2567
rect 3713 2533 3727 2547
rect 3693 2293 3707 2307
rect 3733 2473 3747 2487
rect 3753 2453 3767 2467
rect 3873 2993 3887 3007
rect 3833 2813 3847 2827
rect 3813 2773 3827 2787
rect 3953 3013 3967 3027
rect 3973 3013 3987 3027
rect 3953 2993 3967 3007
rect 4013 3013 4027 3027
rect 3993 2993 4007 3007
rect 3913 2973 3927 2987
rect 3993 2973 4007 2987
rect 3973 2953 3987 2967
rect 3933 2933 3947 2947
rect 3873 2793 3887 2807
rect 3913 2793 3927 2807
rect 3953 2873 3967 2887
rect 3953 2813 3967 2827
rect 3893 2773 3907 2787
rect 3793 2753 3807 2767
rect 3893 2753 3907 2767
rect 3953 2773 3967 2787
rect 3853 2733 3867 2747
rect 3833 2713 3847 2727
rect 3813 2673 3827 2687
rect 3793 2593 3807 2607
rect 3793 2573 3807 2587
rect 3793 2513 3807 2527
rect 3813 2493 3827 2507
rect 3813 2353 3827 2367
rect 3793 2313 3807 2327
rect 3773 2293 3787 2307
rect 3693 2273 3707 2287
rect 3713 2273 3727 2287
rect 3793 2253 3807 2267
rect 3893 2713 3907 2727
rect 3873 2693 3887 2707
rect 3933 2733 3947 2747
rect 3913 2673 3927 2687
rect 3933 2673 3947 2687
rect 3973 2753 3987 2767
rect 3993 2713 4007 2727
rect 3973 2693 3987 2707
rect 3873 2633 3887 2647
rect 3913 2533 3927 2547
rect 3933 2553 3947 2567
rect 4033 2973 4047 2987
rect 4093 3173 4107 3187
rect 4053 2953 4067 2967
rect 4093 2933 4107 2947
rect 4233 3593 4247 3607
rect 4213 3513 4227 3527
rect 4293 3693 4307 3707
rect 4333 3713 4347 3727
rect 4353 3713 4367 3727
rect 4333 3673 4347 3687
rect 4373 3673 4387 3687
rect 4373 3553 4387 3567
rect 4413 3713 4427 3727
rect 4413 3653 4427 3667
rect 4673 4073 4687 4087
rect 4613 4013 4627 4027
rect 4673 4013 4687 4027
rect 4593 3973 4607 3987
rect 4633 3993 4647 4007
rect 4653 3973 4667 3987
rect 4693 3973 4707 3987
rect 4613 3953 4627 3967
rect 4533 3933 4547 3947
rect 4553 3933 4567 3947
rect 4473 3893 4487 3907
rect 4473 3813 4487 3827
rect 4453 3633 4467 3647
rect 4453 3553 4467 3567
rect 4293 3533 4307 3547
rect 4393 3533 4407 3547
rect 4273 3513 4287 3527
rect 4313 3513 4327 3527
rect 4373 3513 4387 3527
rect 4213 3473 4227 3487
rect 4253 3493 4267 3507
rect 4273 3493 4287 3507
rect 4253 3473 4267 3487
rect 4333 3493 4347 3507
rect 4213 3453 4227 3467
rect 4353 3473 4367 3487
rect 4293 3453 4307 3467
rect 4353 3453 4367 3467
rect 4193 3293 4207 3307
rect 4173 3273 4187 3287
rect 4273 3393 4287 3407
rect 4233 3373 4247 3387
rect 4153 3253 4167 3267
rect 4213 3253 4227 3267
rect 4153 3213 4167 3227
rect 4173 3213 4187 3227
rect 4133 3173 4147 3187
rect 4193 3153 4207 3167
rect 4173 3133 4187 3147
rect 4133 3113 4147 3127
rect 4173 3053 4187 3067
rect 4213 3053 4227 3067
rect 4253 3173 4267 3187
rect 4353 3433 4367 3447
rect 4293 3273 4307 3287
rect 4333 3273 4347 3287
rect 4293 3253 4307 3267
rect 4293 3213 4307 3227
rect 4313 3213 4327 3227
rect 4273 3113 4287 3127
rect 4233 3033 4247 3047
rect 4153 2993 4167 3007
rect 4213 3013 4227 3027
rect 4253 3013 4267 3027
rect 4233 2993 4247 3007
rect 4313 3193 4327 3207
rect 4493 3713 4507 3727
rect 4553 3913 4567 3927
rect 4573 3873 4587 3887
rect 4693 3953 4707 3967
rect 4713 3953 4727 3967
rect 4653 3813 4667 3827
rect 4593 3733 4607 3747
rect 4493 3633 4507 3647
rect 4493 3533 4507 3547
rect 4393 3493 4407 3507
rect 4473 3513 4487 3527
rect 4573 3673 4587 3687
rect 4553 3533 4567 3547
rect 4373 3413 4387 3427
rect 4373 3393 4387 3407
rect 4493 3493 4507 3507
rect 4533 3493 4547 3507
rect 4433 3473 4447 3487
rect 4413 3453 4427 3467
rect 4413 3353 4427 3367
rect 4393 3293 4407 3307
rect 4513 3453 4527 3467
rect 4493 3433 4507 3447
rect 4473 3273 4487 3287
rect 4413 3253 4427 3267
rect 4433 3253 4447 3267
rect 4353 3233 4367 3247
rect 4373 3233 4387 3247
rect 4433 3233 4447 3247
rect 4413 3213 4427 3227
rect 4373 3193 4387 3207
rect 4413 3193 4427 3207
rect 4333 3173 4347 3187
rect 4333 3133 4347 3147
rect 4313 3113 4327 3127
rect 4213 2973 4227 2987
rect 4373 3053 4387 3067
rect 4373 3013 4387 3027
rect 4393 3013 4407 3027
rect 4333 2993 4347 3007
rect 4313 2973 4327 2987
rect 4173 2953 4187 2967
rect 4173 2893 4187 2907
rect 4153 2873 4167 2887
rect 4233 2873 4247 2887
rect 4113 2773 4127 2787
rect 4173 2773 4187 2787
rect 4033 2753 4047 2767
rect 4073 2753 4087 2767
rect 4093 2733 4107 2747
rect 4113 2753 4127 2767
rect 4193 2753 4207 2767
rect 4273 2813 4287 2827
rect 4133 2733 4147 2747
rect 4053 2713 4067 2727
rect 4073 2693 4087 2707
rect 4033 2653 4047 2667
rect 4013 2613 4027 2627
rect 4053 2633 4067 2647
rect 4073 2573 4087 2587
rect 4113 2573 4127 2587
rect 4033 2553 4047 2567
rect 4053 2553 4067 2567
rect 3873 2513 3887 2527
rect 4033 2533 4047 2547
rect 4053 2513 4067 2527
rect 3913 2493 3927 2507
rect 3953 2493 3967 2507
rect 3993 2493 4007 2507
rect 3873 2433 3887 2447
rect 3873 2293 3887 2307
rect 3733 2173 3747 2187
rect 3773 2173 3787 2187
rect 3713 2153 3727 2167
rect 3853 2253 3867 2267
rect 3833 2233 3847 2247
rect 3853 2233 3867 2247
rect 3833 2213 3847 2227
rect 3813 2193 3827 2207
rect 3793 2073 3807 2087
rect 3593 2053 3607 2067
rect 3633 2053 3647 2067
rect 3673 2053 3687 2067
rect 3693 2053 3707 2067
rect 3453 2013 3467 2027
rect 3513 1993 3527 2007
rect 3473 1833 3487 1847
rect 3393 1773 3407 1787
rect 3433 1773 3447 1787
rect 3453 1773 3467 1787
rect 3393 1713 3407 1727
rect 3333 1553 3347 1567
rect 3353 1573 3367 1587
rect 3313 1373 3327 1387
rect 3313 1353 3327 1367
rect 3273 1293 3287 1307
rect 3293 1293 3307 1307
rect 3493 1673 3507 1687
rect 3613 2033 3627 2047
rect 3673 2033 3687 2047
rect 3733 2053 3747 2067
rect 3713 2033 3727 2047
rect 3633 2013 3647 2027
rect 3653 2013 3667 2027
rect 3633 1953 3647 1967
rect 3613 1873 3627 1887
rect 3533 1813 3547 1827
rect 3593 1813 3607 1827
rect 3533 1773 3547 1787
rect 3573 1793 3587 1807
rect 3633 1773 3647 1787
rect 3553 1753 3567 1767
rect 3633 1733 3647 1747
rect 3593 1673 3607 1687
rect 3493 1653 3507 1667
rect 3513 1653 3527 1667
rect 3453 1613 3467 1627
rect 3493 1613 3507 1627
rect 3433 1593 3447 1607
rect 3413 1573 3427 1587
rect 3473 1593 3487 1607
rect 3533 1633 3547 1647
rect 3773 2053 3787 2067
rect 3793 2033 3807 2047
rect 3793 1993 3807 2007
rect 3733 1973 3747 1987
rect 3753 1973 3767 1987
rect 3693 1873 3707 1887
rect 3693 1853 3707 1867
rect 3713 1853 3727 1867
rect 3673 1773 3687 1787
rect 3653 1713 3667 1727
rect 3633 1673 3647 1687
rect 3653 1673 3667 1687
rect 3613 1633 3627 1647
rect 3713 1753 3727 1767
rect 3833 2033 3847 2047
rect 3833 1893 3847 1907
rect 3993 2433 4007 2447
rect 3913 2273 3927 2287
rect 3953 2273 3967 2287
rect 3893 2193 3907 2207
rect 3893 2133 3907 2147
rect 3873 2073 3887 2087
rect 3973 2233 3987 2247
rect 3953 2193 3967 2207
rect 3933 2093 3947 2107
rect 3873 2033 3887 2047
rect 3853 1873 3867 1887
rect 3853 1833 3867 1847
rect 3733 1733 3747 1747
rect 3753 1733 3767 1747
rect 3753 1713 3767 1727
rect 3693 1653 3707 1667
rect 3673 1613 3687 1627
rect 3713 1633 3727 1647
rect 3513 1573 3527 1587
rect 3393 1533 3407 1547
rect 3373 1473 3387 1487
rect 3353 1373 3367 1387
rect 3333 1333 3347 1347
rect 3513 1553 3527 1567
rect 3573 1573 3587 1587
rect 3593 1573 3607 1587
rect 3673 1573 3687 1587
rect 3713 1573 3727 1587
rect 3733 1573 3747 1587
rect 3553 1513 3567 1527
rect 3453 1493 3467 1507
rect 3553 1433 3567 1447
rect 3473 1413 3487 1427
rect 3373 1333 3387 1347
rect 3353 1313 3367 1327
rect 3393 1313 3407 1327
rect 3313 1273 3327 1287
rect 3373 1273 3387 1287
rect 3293 1153 3307 1167
rect 3133 1093 3147 1107
rect 3153 1113 3167 1127
rect 3193 1113 3207 1127
rect 3233 1113 3247 1127
rect 3173 1093 3187 1107
rect 3133 1053 3147 1067
rect 3133 1033 3147 1047
rect 3093 1013 3107 1027
rect 3053 913 3067 927
rect 3013 873 3027 887
rect 2993 853 3007 867
rect 2873 773 2887 787
rect 2913 773 2927 787
rect 2853 653 2867 667
rect 2993 833 3007 847
rect 3013 833 3027 847
rect 3033 853 3047 867
rect 2953 753 2967 767
rect 2953 733 2967 747
rect 2933 653 2947 667
rect 3033 813 3047 827
rect 3013 793 3027 807
rect 2993 713 3007 727
rect 2993 673 3007 687
rect 2873 633 2887 647
rect 2893 633 2907 647
rect 2913 613 2927 627
rect 2953 633 2967 647
rect 3113 853 3127 867
rect 3093 833 3107 847
rect 3073 793 3087 807
rect 3053 753 3067 767
rect 3033 713 3047 727
rect 2853 593 2867 607
rect 2893 593 2907 607
rect 2833 573 2847 587
rect 2773 533 2787 547
rect 2693 453 2707 467
rect 2753 453 2767 467
rect 2633 413 2647 427
rect 2593 373 2607 387
rect 2633 393 2647 407
rect 2573 293 2587 307
rect 2353 193 2367 207
rect 2373 193 2387 207
rect 2433 193 2447 207
rect 2413 173 2427 187
rect 2373 153 2387 167
rect 2493 153 2507 167
rect 2473 133 2487 147
rect 1993 113 2007 127
rect 2053 113 2067 127
rect 2153 113 2167 127
rect 2673 293 2687 307
rect 2613 193 2627 207
rect 1913 93 1927 107
rect 2773 433 2787 447
rect 2713 333 2727 347
rect 2733 133 2747 147
rect 2913 413 2927 427
rect 2793 353 2807 367
rect 2853 373 2867 387
rect 2833 333 2847 347
rect 2893 393 2907 407
rect 3053 633 3067 647
rect 3073 633 3087 647
rect 3153 913 3167 927
rect 3193 913 3207 927
rect 3213 913 3227 927
rect 3193 893 3207 907
rect 3213 833 3227 847
rect 3173 813 3187 827
rect 3173 793 3187 807
rect 3233 793 3247 807
rect 3213 753 3227 767
rect 3133 733 3147 747
rect 3233 713 3247 727
rect 3173 673 3187 687
rect 3193 653 3207 667
rect 3173 613 3187 627
rect 3193 613 3207 627
rect 3053 573 3067 587
rect 2993 393 3007 407
rect 3033 393 3047 407
rect 3073 393 3087 407
rect 2953 353 2967 367
rect 2893 313 2907 327
rect 2813 293 2827 307
rect 2873 293 2887 307
rect 2853 153 2867 167
rect 3053 333 3067 347
rect 3033 313 3047 327
rect 2973 273 2987 287
rect 3053 273 3067 287
rect 2873 133 2887 147
rect 2933 193 2947 207
rect 3033 193 3047 207
rect 2953 173 2967 187
rect 2973 133 2987 147
rect 2993 153 3007 167
rect 3013 133 3027 147
rect 3053 113 3067 127
rect 2773 53 2787 67
rect 2693 33 2707 47
rect 3153 553 3167 567
rect 3173 473 3187 487
rect 3173 453 3187 467
rect 3153 393 3167 407
rect 3113 353 3127 367
rect 3093 313 3107 327
rect 3133 313 3147 327
rect 3213 593 3227 607
rect 3233 413 3247 427
rect 3193 393 3207 407
rect 3193 333 3207 347
rect 3273 1133 3287 1147
rect 3273 1093 3287 1107
rect 3453 1333 3467 1347
rect 3353 1233 3367 1247
rect 3413 1233 3427 1247
rect 3393 1173 3407 1187
rect 3333 1153 3347 1167
rect 3333 1113 3347 1127
rect 3333 1073 3347 1087
rect 3353 1093 3367 1107
rect 3453 1293 3467 1307
rect 3533 1373 3547 1387
rect 3493 1333 3507 1347
rect 3473 1253 3487 1267
rect 3453 1233 3467 1247
rect 3533 1333 3547 1347
rect 3573 1413 3587 1427
rect 3593 1393 3607 1407
rect 3633 1553 3647 1567
rect 3673 1533 3687 1547
rect 3613 1353 3627 1367
rect 3593 1333 3607 1347
rect 3513 1313 3527 1327
rect 3593 1293 3607 1307
rect 3633 1293 3647 1307
rect 3533 1253 3547 1267
rect 3533 1233 3547 1247
rect 3493 1213 3507 1227
rect 3493 1153 3507 1167
rect 3553 1193 3567 1207
rect 3593 1273 3607 1287
rect 3653 1253 3667 1267
rect 3633 1173 3647 1187
rect 3713 1513 3727 1527
rect 3793 1733 3807 1747
rect 3773 1653 3787 1667
rect 3773 1613 3787 1627
rect 3873 1813 3887 1827
rect 3933 2053 3947 2067
rect 4013 2293 4027 2307
rect 4033 2253 4047 2267
rect 4153 2713 4167 2727
rect 4173 2713 4187 2727
rect 4153 2613 4167 2627
rect 4313 2753 4327 2767
rect 4313 2733 4327 2747
rect 4233 2673 4247 2687
rect 4193 2633 4207 2647
rect 4153 2573 4167 2587
rect 4173 2573 4187 2587
rect 4133 2553 4147 2567
rect 4193 2553 4207 2567
rect 4213 2533 4227 2547
rect 4133 2513 4147 2527
rect 4073 2473 4087 2487
rect 4073 2353 4087 2367
rect 4053 2233 4067 2247
rect 4193 2513 4207 2527
rect 4173 2493 4187 2507
rect 4153 2453 4167 2467
rect 4153 2413 4167 2427
rect 4133 2393 4147 2407
rect 4153 2373 4167 2387
rect 4093 2333 4107 2347
rect 4133 2333 4147 2347
rect 4153 2293 4167 2307
rect 4093 2253 4107 2267
rect 4133 2273 4147 2287
rect 4293 2673 4307 2687
rect 4253 2613 4267 2627
rect 4253 2513 4267 2527
rect 4273 2533 4287 2547
rect 4353 2953 4367 2967
rect 4393 2993 4407 3007
rect 4473 3233 4487 3247
rect 4513 3233 4527 3247
rect 4493 3213 4507 3227
rect 4453 3173 4467 3187
rect 4433 3133 4447 3147
rect 4613 3713 4627 3727
rect 4653 3733 4667 3747
rect 4653 3713 4667 3727
rect 4593 3613 4607 3627
rect 4613 3573 4627 3587
rect 4573 3513 4587 3527
rect 4593 3513 4607 3527
rect 4693 3693 4707 3707
rect 4673 3673 4687 3687
rect 4693 3613 4707 3627
rect 4673 3573 4687 3587
rect 4653 3533 4667 3547
rect 4633 3493 4647 3507
rect 4773 4213 4787 4227
rect 4753 3953 4767 3967
rect 4753 3933 4767 3947
rect 4733 3833 4747 3847
rect 4733 3813 4747 3827
rect 4733 3693 4747 3707
rect 4733 3673 4747 3687
rect 4693 3513 4707 3527
rect 4713 3513 4727 3527
rect 4693 3493 4707 3507
rect 4653 3453 4667 3467
rect 4693 3453 4707 3467
rect 4573 3433 4587 3447
rect 4633 3413 4647 3427
rect 4593 3333 4607 3347
rect 4553 3253 4567 3267
rect 4593 3253 4607 3267
rect 4673 3433 4687 3447
rect 4713 3433 4727 3447
rect 4773 3733 4787 3747
rect 4753 3633 4767 3647
rect 4753 3613 4767 3627
rect 4773 3573 4787 3587
rect 4753 3433 4767 3447
rect 4733 3413 4747 3427
rect 4753 3393 4767 3407
rect 4733 3373 4747 3387
rect 4733 3293 4747 3307
rect 4693 3273 4707 3287
rect 4653 3253 4667 3267
rect 4553 3213 4567 3227
rect 4573 3233 4587 3247
rect 4613 3233 4627 3247
rect 4633 3233 4647 3247
rect 4573 3173 4587 3187
rect 4533 3153 4547 3167
rect 4513 3133 4527 3147
rect 4493 3073 4507 3087
rect 4493 3053 4507 3067
rect 4453 3013 4467 3027
rect 4493 3013 4507 3027
rect 4553 3093 4567 3107
rect 4573 3053 4587 3067
rect 4613 3193 4627 3207
rect 4713 3253 4727 3267
rect 4713 3233 4727 3247
rect 4733 3233 4747 3247
rect 4693 3213 4707 3227
rect 4653 3173 4667 3187
rect 4653 3093 4667 3107
rect 4673 3073 4687 3087
rect 4653 3053 4667 3067
rect 4693 3053 4707 3067
rect 4773 3193 4787 3207
rect 4753 3113 4767 3127
rect 4733 3053 4747 3067
rect 4553 3013 4567 3027
rect 4473 2993 4487 3007
rect 4513 2993 4527 3007
rect 4533 2993 4547 3007
rect 4433 2973 4447 2987
rect 4493 2973 4507 2987
rect 4413 2913 4427 2927
rect 4373 2793 4387 2807
rect 4513 2953 4527 2967
rect 4553 2973 4567 2987
rect 4353 2713 4367 2727
rect 4493 2773 4507 2787
rect 4433 2753 4447 2767
rect 4413 2733 4427 2747
rect 4393 2713 4407 2727
rect 4373 2653 4387 2667
rect 4453 2733 4467 2747
rect 4473 2753 4487 2767
rect 4513 2753 4527 2767
rect 4533 2733 4547 2747
rect 4433 2693 4447 2707
rect 4433 2633 4447 2647
rect 4393 2613 4407 2627
rect 4413 2613 4427 2627
rect 4393 2553 4407 2567
rect 4333 2533 4347 2547
rect 4313 2513 4327 2527
rect 4333 2513 4347 2527
rect 4353 2513 4367 2527
rect 4373 2533 4387 2547
rect 4393 2513 4407 2527
rect 4293 2473 4307 2487
rect 4253 2453 4267 2467
rect 4233 2413 4247 2427
rect 4193 2393 4207 2407
rect 4193 2373 4207 2387
rect 4373 2493 4387 2507
rect 4413 2493 4427 2507
rect 4353 2413 4367 2427
rect 4253 2333 4267 2347
rect 4333 2333 4347 2347
rect 4233 2273 4247 2287
rect 4273 2273 4287 2287
rect 4153 2253 4167 2267
rect 4193 2253 4207 2267
rect 4093 2233 4107 2247
rect 4173 2233 4187 2247
rect 4093 2213 4107 2227
rect 4113 2213 4127 2227
rect 4093 2093 4107 2107
rect 3913 2033 3927 2047
rect 3933 1953 3947 1967
rect 3953 1893 3967 1907
rect 3913 1813 3927 1827
rect 3893 1773 3907 1787
rect 3913 1773 3927 1787
rect 3933 1773 3947 1787
rect 3873 1753 3887 1767
rect 3913 1713 3927 1727
rect 3893 1653 3907 1667
rect 4053 2053 4067 2067
rect 4133 2073 4147 2087
rect 4053 1833 4067 1847
rect 4013 1813 4027 1827
rect 4033 1813 4047 1827
rect 4113 2013 4127 2027
rect 4073 1813 4087 1827
rect 4153 1853 4167 1867
rect 4153 1833 4167 1847
rect 4193 2213 4207 2227
rect 4253 2253 4267 2267
rect 4313 2273 4327 2287
rect 4233 2193 4247 2207
rect 4213 2173 4227 2187
rect 4333 2253 4347 2267
rect 4373 2373 4387 2387
rect 4373 2353 4387 2367
rect 4313 2233 4327 2247
rect 4353 2233 4367 2247
rect 4213 2113 4227 2127
rect 4293 2173 4307 2187
rect 4253 2133 4267 2147
rect 4513 2673 4527 2687
rect 4533 2673 4547 2687
rect 4593 3013 4607 3027
rect 4633 3013 4647 3027
rect 4693 3013 4707 3027
rect 4613 2993 4627 3007
rect 4613 2833 4627 2847
rect 4673 2793 4687 2807
rect 4573 2773 4587 2787
rect 4613 2773 4627 2787
rect 4593 2753 4607 2767
rect 4573 2713 4587 2727
rect 4593 2693 4607 2707
rect 4553 2653 4567 2667
rect 4533 2573 4547 2587
rect 4553 2573 4567 2587
rect 4493 2553 4507 2567
rect 4513 2553 4527 2567
rect 4473 2533 4487 2547
rect 4513 2533 4527 2547
rect 4493 2513 4507 2527
rect 4573 2513 4587 2527
rect 4553 2493 4567 2507
rect 4493 2473 4507 2487
rect 4533 2473 4547 2487
rect 4453 2433 4467 2447
rect 4413 2313 4427 2327
rect 4433 2313 4447 2327
rect 4553 2413 4567 2427
rect 4513 2393 4527 2407
rect 4553 2333 4567 2347
rect 4493 2293 4507 2307
rect 4513 2293 4527 2307
rect 4393 2273 4407 2287
rect 4413 2253 4427 2267
rect 4433 2273 4447 2287
rect 4493 2273 4507 2287
rect 4533 2273 4547 2287
rect 4533 2253 4547 2267
rect 4373 2133 4387 2147
rect 4433 2213 4447 2227
rect 4233 2073 4247 2087
rect 4193 2013 4207 2027
rect 4313 2073 4327 2087
rect 4333 2053 4347 2067
rect 4353 2053 4367 2067
rect 4373 2053 4387 2067
rect 4413 2073 4427 2087
rect 4273 2013 4287 2027
rect 4233 1993 4247 2007
rect 4293 1993 4307 2007
rect 4313 1953 4327 1967
rect 4213 1873 4227 1887
rect 4253 1833 4267 1847
rect 3973 1773 3987 1787
rect 4073 1773 4087 1787
rect 4093 1773 4107 1787
rect 4213 1813 4227 1827
rect 4273 1793 4287 1807
rect 4193 1773 4207 1787
rect 3993 1753 4007 1767
rect 4013 1753 4027 1767
rect 3993 1693 4007 1707
rect 4073 1753 4087 1767
rect 4053 1733 4067 1747
rect 4033 1713 4047 1727
rect 3973 1653 3987 1667
rect 4013 1653 4027 1667
rect 3813 1633 3827 1647
rect 3853 1633 3867 1647
rect 3953 1633 3967 1647
rect 3813 1593 3827 1607
rect 3773 1573 3787 1587
rect 3793 1573 3807 1587
rect 3753 1453 3767 1467
rect 3793 1393 3807 1407
rect 3773 1353 3787 1367
rect 3753 1333 3767 1347
rect 3693 1293 3707 1307
rect 3713 1293 3727 1307
rect 3733 1293 3747 1307
rect 3833 1333 3847 1347
rect 3893 1613 3907 1627
rect 3953 1613 3967 1627
rect 3873 1573 3887 1587
rect 3893 1573 3907 1587
rect 3933 1593 3947 1607
rect 3913 1553 3927 1567
rect 3933 1473 3947 1487
rect 3893 1353 3907 1367
rect 3853 1293 3867 1307
rect 3813 1273 3827 1287
rect 3693 1213 3707 1227
rect 3713 1213 3727 1227
rect 3773 1213 3787 1227
rect 3773 1173 3787 1187
rect 3613 1133 3627 1147
rect 3673 1133 3687 1147
rect 3693 1133 3707 1147
rect 3453 1073 3467 1087
rect 3473 1073 3487 1087
rect 3573 1113 3587 1127
rect 3553 1073 3567 1087
rect 3413 1053 3427 1067
rect 3493 1053 3507 1067
rect 3533 1053 3547 1067
rect 3313 1033 3327 1047
rect 3293 973 3307 987
rect 3273 893 3287 907
rect 3273 873 3287 887
rect 3373 1013 3387 1027
rect 3273 753 3287 767
rect 3353 873 3367 887
rect 3313 853 3327 867
rect 3333 793 3347 807
rect 3473 993 3487 1007
rect 3393 853 3407 867
rect 3393 813 3407 827
rect 3413 813 3427 827
rect 3373 753 3387 767
rect 3353 713 3367 727
rect 3373 713 3387 727
rect 3313 693 3327 707
rect 3353 693 3367 707
rect 3333 673 3347 687
rect 3293 653 3307 667
rect 3313 653 3327 667
rect 3273 633 3287 647
rect 3273 593 3287 607
rect 3313 593 3327 607
rect 3413 773 3427 787
rect 3453 773 3467 787
rect 3453 693 3467 707
rect 3393 673 3407 687
rect 3433 673 3447 687
rect 3393 653 3407 667
rect 3593 1053 3607 1067
rect 3553 973 3567 987
rect 3513 933 3527 947
rect 3633 1113 3647 1127
rect 3673 1113 3687 1127
rect 3713 1113 3727 1127
rect 3653 1033 3667 1047
rect 3633 1013 3647 1027
rect 3613 913 3627 927
rect 3553 873 3567 887
rect 3613 873 3627 887
rect 3493 853 3507 867
rect 3493 813 3507 827
rect 3593 853 3607 867
rect 3533 813 3547 827
rect 3573 813 3587 827
rect 3493 793 3507 807
rect 3473 653 3487 667
rect 3513 733 3527 747
rect 3553 733 3567 747
rect 3513 693 3527 707
rect 3413 633 3427 647
rect 3453 613 3467 627
rect 3473 633 3487 647
rect 3893 1333 3907 1347
rect 3913 1173 3927 1187
rect 3813 1133 3827 1147
rect 3833 1133 3847 1147
rect 3873 1133 3887 1147
rect 3773 1093 3787 1107
rect 3833 1093 3847 1107
rect 3873 1093 3887 1107
rect 3793 1073 3807 1087
rect 3713 933 3727 947
rect 3653 873 3667 887
rect 3893 1073 3907 1087
rect 3873 1053 3887 1067
rect 3673 753 3687 767
rect 3633 733 3647 747
rect 3613 693 3627 707
rect 3713 813 3727 827
rect 3693 693 3707 707
rect 3673 653 3687 667
rect 3713 653 3727 667
rect 3573 613 3587 627
rect 3353 593 3367 607
rect 3453 593 3467 607
rect 3453 533 3467 547
rect 3533 533 3547 547
rect 3353 433 3367 447
rect 3273 393 3287 407
rect 3433 393 3447 407
rect 3273 373 3287 387
rect 3253 353 3267 367
rect 3313 373 3327 387
rect 3353 373 3367 387
rect 3233 293 3247 307
rect 3213 273 3227 287
rect 3153 173 3167 187
rect 3213 193 3227 207
rect 3173 153 3187 167
rect 3373 353 3387 367
rect 3413 353 3427 367
rect 3393 333 3407 347
rect 3333 293 3347 307
rect 3353 293 3367 307
rect 3313 193 3327 207
rect 3353 193 3367 207
rect 3253 173 3267 187
rect 3293 173 3307 187
rect 3093 113 3107 127
rect 3273 153 3287 167
rect 3413 173 3427 187
rect 3293 133 3307 147
rect 3273 113 3287 127
rect 3333 113 3347 127
rect 3393 133 3407 147
rect 3553 453 3567 467
rect 3553 393 3567 407
rect 3513 373 3527 387
rect 3473 353 3487 367
rect 3493 313 3507 327
rect 3673 613 3687 627
rect 3713 613 3727 627
rect 3633 593 3647 607
rect 3753 853 3767 867
rect 3793 853 3807 867
rect 3793 833 3807 847
rect 3813 833 3827 847
rect 3833 853 3847 867
rect 3873 853 3887 867
rect 3753 793 3767 807
rect 3773 793 3787 807
rect 3873 813 3887 827
rect 3853 793 3867 807
rect 3813 713 3827 727
rect 3873 693 3887 707
rect 3793 653 3807 667
rect 3813 653 3827 667
rect 4033 1633 4047 1647
rect 4013 1613 4027 1627
rect 3993 1573 4007 1587
rect 4133 1693 4147 1707
rect 4093 1653 4107 1667
rect 4053 1613 4067 1627
rect 4073 1613 4087 1627
rect 4033 1573 4047 1587
rect 4013 1553 4027 1567
rect 4013 1513 4027 1527
rect 4013 1413 4027 1427
rect 3993 1393 4007 1407
rect 3993 1333 4007 1347
rect 4113 1633 4127 1647
rect 4093 1593 4107 1607
rect 4213 1753 4227 1767
rect 4173 1693 4187 1707
rect 4153 1653 4167 1667
rect 4193 1653 4207 1667
rect 4273 1753 4287 1767
rect 4453 2093 4467 2107
rect 4433 1993 4447 2007
rect 4393 1893 4407 1907
rect 4333 1853 4347 1867
rect 4333 1833 4347 1847
rect 4373 1853 4387 1867
rect 4353 1813 4367 1827
rect 4493 2233 4507 2247
rect 4533 2213 4547 2227
rect 4513 2193 4527 2207
rect 4713 2813 4727 2827
rect 4693 2773 4707 2787
rect 4633 2753 4647 2767
rect 4693 2733 4707 2747
rect 4733 2793 4747 2807
rect 4633 2713 4647 2727
rect 4713 2713 4727 2727
rect 4653 2673 4667 2687
rect 4653 2653 4667 2667
rect 4773 3073 4787 3087
rect 4753 2753 4767 2767
rect 4733 2673 4747 2687
rect 4713 2633 4727 2647
rect 4693 2613 4707 2627
rect 4653 2553 4667 2567
rect 4653 2513 4667 2527
rect 4673 2533 4687 2547
rect 4693 2513 4707 2527
rect 4673 2493 4687 2507
rect 4713 2493 4727 2507
rect 4633 2453 4647 2467
rect 4653 2453 4667 2467
rect 4613 2353 4627 2367
rect 4633 2313 4647 2327
rect 4693 2473 4707 2487
rect 4673 2373 4687 2387
rect 4653 2293 4667 2307
rect 4713 2433 4727 2447
rect 4713 2393 4727 2407
rect 4733 2393 4747 2407
rect 4553 2173 4567 2187
rect 4653 2253 4667 2267
rect 4693 2273 4707 2287
rect 4733 2253 4747 2267
rect 4653 2233 4667 2247
rect 4693 2233 4707 2247
rect 4593 2173 4607 2187
rect 4613 2173 4627 2187
rect 4493 2113 4507 2127
rect 4513 2113 4527 2127
rect 4573 2113 4587 2127
rect 4553 2073 4567 2087
rect 4513 2053 4527 2067
rect 4553 2053 4567 2067
rect 4493 2033 4507 2047
rect 4453 1813 4467 1827
rect 4633 2113 4647 2127
rect 4593 2073 4607 2087
rect 4593 2053 4607 2067
rect 4613 2033 4627 2047
rect 4533 2013 4547 2027
rect 4513 1853 4527 1867
rect 4573 1993 4587 2007
rect 4553 1873 4567 1887
rect 4533 1833 4547 1847
rect 4513 1813 4527 1827
rect 4393 1773 4407 1787
rect 4413 1793 4427 1807
rect 4453 1793 4467 1807
rect 4493 1793 4507 1807
rect 4473 1773 4487 1787
rect 4353 1753 4367 1767
rect 4373 1753 4387 1767
rect 4313 1733 4327 1747
rect 4293 1693 4307 1707
rect 4333 1673 4347 1687
rect 4233 1633 4247 1647
rect 4173 1613 4187 1627
rect 4193 1613 4207 1627
rect 4213 1613 4227 1627
rect 4133 1593 4147 1607
rect 4193 1573 4207 1587
rect 4213 1593 4227 1607
rect 4233 1573 4247 1587
rect 4273 1573 4287 1587
rect 4293 1593 4307 1607
rect 4313 1573 4327 1587
rect 4133 1553 4147 1567
rect 4093 1533 4107 1547
rect 4113 1533 4127 1547
rect 4153 1513 4167 1527
rect 4213 1513 4227 1527
rect 4073 1433 4087 1447
rect 4073 1373 4087 1387
rect 4053 1333 4067 1347
rect 4113 1433 4127 1447
rect 4093 1353 4107 1367
rect 4093 1333 4107 1347
rect 3973 1313 3987 1327
rect 4013 1313 4027 1327
rect 4033 1293 4047 1307
rect 4053 1253 4067 1267
rect 3993 1233 4007 1247
rect 4013 1213 4027 1227
rect 3993 1193 4007 1207
rect 3953 1093 3967 1107
rect 3973 1093 3987 1107
rect 3933 1013 3947 1027
rect 4193 1453 4207 1467
rect 4173 1433 4187 1447
rect 4133 1373 4147 1387
rect 4153 1373 4167 1387
rect 4113 1293 4127 1307
rect 4133 1293 4147 1307
rect 4133 1253 4147 1267
rect 4133 1213 4147 1227
rect 4093 1153 4107 1167
rect 4053 1133 4067 1147
rect 4173 1293 4187 1307
rect 4153 1193 4167 1207
rect 4273 1553 4287 1567
rect 4273 1453 4287 1467
rect 4233 1413 4247 1427
rect 4213 1353 4227 1367
rect 4353 1653 4367 1667
rect 4473 1733 4487 1747
rect 4393 1633 4407 1647
rect 4433 1633 4447 1647
rect 4453 1633 4467 1647
rect 4373 1573 4387 1587
rect 4373 1553 4387 1567
rect 4353 1453 4367 1467
rect 4333 1393 4347 1407
rect 4313 1373 4327 1387
rect 4433 1613 4447 1627
rect 4413 1593 4427 1607
rect 4433 1573 4447 1587
rect 4453 1553 4467 1567
rect 4433 1533 4447 1547
rect 4393 1513 4407 1527
rect 4413 1373 4427 1387
rect 4353 1353 4367 1367
rect 4373 1353 4387 1367
rect 4313 1333 4327 1347
rect 4273 1313 4287 1327
rect 4253 1293 4267 1307
rect 4253 1253 4267 1267
rect 4293 1293 4307 1307
rect 4673 2193 4687 2207
rect 4693 2173 4707 2187
rect 4733 2233 4747 2247
rect 4773 2693 4787 2707
rect 4773 2673 4787 2687
rect 4773 2453 4787 2467
rect 4773 2313 4787 2327
rect 4773 2273 4787 2287
rect 4773 2233 4787 2247
rect 4753 2193 4767 2207
rect 4733 2133 4747 2147
rect 4713 2093 4727 2107
rect 4693 2073 4707 2087
rect 4673 2033 4687 2047
rect 4693 2013 4707 2027
rect 4633 1873 4647 1887
rect 4653 1853 4667 1867
rect 4713 1993 4727 2007
rect 4713 1933 4727 1947
rect 4633 1833 4647 1847
rect 4573 1813 4587 1827
rect 4613 1813 4627 1827
rect 4693 1833 4707 1847
rect 4533 1793 4547 1807
rect 4553 1793 4567 1807
rect 4633 1793 4647 1807
rect 4673 1793 4687 1807
rect 4613 1773 4627 1787
rect 4653 1773 4667 1787
rect 4553 1753 4567 1767
rect 4573 1753 4587 1767
rect 4613 1753 4627 1767
rect 4693 1753 4707 1767
rect 4673 1713 4687 1727
rect 4693 1713 4707 1727
rect 4653 1633 4667 1647
rect 4613 1613 4627 1627
rect 4513 1593 4527 1607
rect 4553 1593 4567 1607
rect 4633 1593 4647 1607
rect 4513 1573 4527 1587
rect 4533 1553 4547 1567
rect 4493 1533 4507 1547
rect 4533 1533 4547 1547
rect 4493 1493 4507 1507
rect 4473 1353 4487 1367
rect 4533 1333 4547 1347
rect 4353 1293 4367 1307
rect 4433 1293 4447 1307
rect 4473 1313 4487 1327
rect 4513 1313 4527 1327
rect 4533 1313 4547 1327
rect 4373 1273 4387 1287
rect 4313 1253 4327 1267
rect 4193 1213 4207 1227
rect 4193 1153 4207 1167
rect 4253 1233 4267 1247
rect 4273 1233 4287 1247
rect 4233 1213 4247 1227
rect 4013 1113 4027 1127
rect 4033 1093 4047 1107
rect 4113 1133 4127 1147
rect 4133 1133 4147 1147
rect 4173 1133 4187 1147
rect 4213 1133 4227 1147
rect 4073 1113 4087 1127
rect 4093 1093 4107 1107
rect 4053 1073 4067 1087
rect 4093 1073 4107 1087
rect 3993 913 4007 927
rect 4073 913 4087 927
rect 4013 893 4027 907
rect 4053 893 4067 907
rect 3973 853 3987 867
rect 3953 833 3967 847
rect 4013 853 4027 867
rect 4033 853 4047 867
rect 4053 833 4067 847
rect 3993 813 4007 827
rect 3933 713 3947 727
rect 3913 673 3927 687
rect 3993 673 4007 687
rect 3933 653 3947 667
rect 3773 613 3787 627
rect 3793 633 3807 647
rect 3753 593 3767 607
rect 3813 593 3827 607
rect 3733 573 3747 587
rect 3713 533 3727 547
rect 3633 433 3647 447
rect 3613 393 3627 407
rect 3693 393 3707 407
rect 3593 373 3607 387
rect 3593 333 3607 347
rect 3553 293 3567 307
rect 3573 293 3587 307
rect 3533 273 3547 287
rect 3653 333 3667 347
rect 3713 333 3727 347
rect 3673 313 3687 327
rect 3613 293 3627 307
rect 3653 293 3667 307
rect 3673 293 3687 307
rect 3573 233 3587 247
rect 3593 233 3607 247
rect 3553 213 3567 227
rect 3453 193 3467 207
rect 3493 173 3507 187
rect 3893 633 3907 647
rect 3953 633 3967 647
rect 3873 593 3887 607
rect 3893 613 3907 627
rect 3913 593 3927 607
rect 3853 553 3867 567
rect 3773 473 3787 487
rect 3753 253 3767 267
rect 3753 213 3767 227
rect 3633 193 3647 207
rect 3733 193 3747 207
rect 3433 153 3447 167
rect 3673 173 3687 187
rect 3713 173 3727 187
rect 3453 133 3467 147
rect 3473 113 3487 127
rect 3533 113 3547 127
rect 3193 93 3207 107
rect 3253 93 3267 107
rect 3373 93 3387 107
rect 3693 153 3707 167
rect 3853 413 3867 427
rect 3793 273 3807 287
rect 3813 233 3827 247
rect 3913 333 3927 347
rect 3873 313 3887 327
rect 3933 313 3947 327
rect 3833 213 3847 227
rect 3893 213 3907 227
rect 3733 153 3747 167
rect 3573 93 3587 107
rect 3773 93 3787 107
rect 3613 73 3627 87
rect 3613 53 3627 67
rect 3573 33 3587 47
rect 3073 13 3087 27
rect 3493 13 3507 27
rect 3873 173 3887 187
rect 3813 153 3827 167
rect 3853 153 3867 167
rect 3933 173 3947 187
rect 4053 793 4067 807
rect 4133 1093 4147 1107
rect 4153 1073 4167 1087
rect 4113 1053 4127 1067
rect 4153 1013 4167 1027
rect 4113 953 4127 967
rect 4093 873 4107 887
rect 4153 933 4167 947
rect 4193 1093 4207 1107
rect 4193 993 4207 1007
rect 4233 1073 4247 1087
rect 4213 913 4227 927
rect 4173 873 4187 887
rect 4113 853 4127 867
rect 4153 853 4167 867
rect 4093 833 4107 847
rect 4133 833 4147 847
rect 4273 1193 4287 1207
rect 4373 1233 4387 1247
rect 4353 1173 4367 1187
rect 4313 1153 4327 1167
rect 4353 1153 4367 1167
rect 4313 1133 4327 1147
rect 4293 1093 4307 1107
rect 4313 1093 4327 1107
rect 4453 1273 4467 1287
rect 4453 1233 4467 1247
rect 4393 1173 4407 1187
rect 4533 1273 4547 1287
rect 4513 1173 4527 1187
rect 4493 1133 4507 1147
rect 4593 1573 4607 1587
rect 4673 1573 4687 1587
rect 4593 1533 4607 1547
rect 4633 1533 4647 1547
rect 4573 1453 4587 1467
rect 4593 1333 4607 1347
rect 4673 1533 4687 1547
rect 4653 1493 4667 1507
rect 4633 1433 4647 1447
rect 4693 1513 4707 1527
rect 4633 1393 4647 1407
rect 4673 1393 4687 1407
rect 4653 1333 4667 1347
rect 4593 1313 4607 1327
rect 4613 1313 4627 1327
rect 4593 1273 4607 1287
rect 4613 1273 4627 1287
rect 4573 1233 4587 1247
rect 4573 1213 4587 1227
rect 4393 1113 4407 1127
rect 4373 1093 4387 1107
rect 4493 1113 4507 1127
rect 4513 1113 4527 1127
rect 4513 1093 4527 1107
rect 4313 1053 4327 1067
rect 4273 1013 4287 1027
rect 4413 1073 4427 1087
rect 4433 1073 4447 1087
rect 4453 1073 4467 1087
rect 4353 1053 4367 1067
rect 4333 973 4347 987
rect 4313 913 4327 927
rect 4253 853 4267 867
rect 4413 1033 4427 1047
rect 4473 1033 4487 1047
rect 4453 933 4467 947
rect 4433 913 4447 927
rect 4433 893 4447 907
rect 4393 853 4407 867
rect 4193 813 4207 827
rect 4233 833 4247 847
rect 4273 833 4287 847
rect 4313 833 4327 847
rect 4353 833 4367 847
rect 4113 773 4127 787
rect 4093 733 4107 747
rect 4173 733 4187 747
rect 4013 653 4027 667
rect 4053 653 4067 667
rect 4073 653 4087 667
rect 4013 633 4027 647
rect 3993 613 4007 627
rect 4033 613 4047 627
rect 4073 613 4087 627
rect 4013 593 4027 607
rect 4053 593 4067 607
rect 3973 533 3987 547
rect 4173 633 4187 647
rect 4113 613 4127 627
rect 4153 613 4167 627
rect 4133 593 4147 607
rect 4173 553 4187 567
rect 4093 533 4107 547
rect 4053 513 4067 527
rect 3973 393 3987 407
rect 4093 393 4107 407
rect 3973 373 3987 387
rect 3993 333 4007 347
rect 4033 333 4047 347
rect 3993 273 4007 287
rect 4033 233 4047 247
rect 3993 213 4007 227
rect 3893 133 3907 147
rect 3953 153 3967 167
rect 3833 93 3847 107
rect 3893 73 3907 87
rect 3993 153 4007 167
rect 4053 213 4067 227
rect 4113 373 4127 387
rect 4233 793 4247 807
rect 4213 753 4227 767
rect 4373 813 4387 827
rect 4413 833 4427 847
rect 4433 813 4447 827
rect 4333 793 4347 807
rect 4393 793 4407 807
rect 4413 793 4427 807
rect 4293 773 4307 787
rect 4393 773 4407 787
rect 4273 753 4287 767
rect 4373 753 4387 767
rect 4213 733 4227 747
rect 4233 733 4247 747
rect 4293 693 4307 707
rect 4353 693 4367 707
rect 4233 653 4247 667
rect 4253 613 4267 627
rect 4233 593 4247 607
rect 4313 633 4327 647
rect 4433 753 4447 767
rect 4413 733 4427 747
rect 4493 913 4507 927
rect 4633 1193 4647 1207
rect 4653 1193 4667 1207
rect 4553 1113 4567 1127
rect 4593 1113 4607 1127
rect 4573 1093 4587 1107
rect 4593 1073 4607 1087
rect 4573 913 4587 927
rect 4613 933 4627 947
rect 4533 893 4547 907
rect 4573 893 4587 907
rect 4593 893 4607 907
rect 4613 893 4627 907
rect 4493 853 4507 867
rect 4473 813 4487 827
rect 4513 813 4527 827
rect 4413 653 4427 667
rect 4453 653 4467 667
rect 4393 633 4407 647
rect 4333 593 4347 607
rect 4373 613 4387 627
rect 4373 593 4387 607
rect 4313 573 4327 587
rect 4453 633 4467 647
rect 4553 773 4567 787
rect 4553 753 4567 767
rect 4533 733 4547 747
rect 4513 653 4527 667
rect 4493 633 4507 647
rect 4513 613 4527 627
rect 4473 593 4487 607
rect 4413 573 4427 587
rect 4293 393 4307 407
rect 4393 513 4407 527
rect 4433 513 4447 527
rect 4353 453 4367 467
rect 4333 393 4347 407
rect 4233 373 4247 387
rect 4153 353 4167 367
rect 4273 373 4287 387
rect 4113 293 4127 307
rect 4093 213 4107 227
rect 4073 193 4087 207
rect 4053 173 4067 187
rect 4013 113 4027 127
rect 4073 153 4087 167
rect 4253 353 4267 367
rect 4313 373 4327 387
rect 4233 333 4247 347
rect 4273 333 4287 347
rect 4353 353 4367 367
rect 4213 293 4227 307
rect 4373 333 4387 347
rect 4313 313 4327 327
rect 4333 313 4347 327
rect 4173 273 4187 287
rect 4233 273 4247 287
rect 4533 533 4547 547
rect 4553 413 4567 427
rect 4513 393 4527 407
rect 4653 1133 4667 1147
rect 4693 1293 4707 1307
rect 4673 1113 4687 1127
rect 4653 1073 4667 1087
rect 4673 1093 4687 1107
rect 4733 1153 4747 1167
rect 4773 2153 4787 2167
rect 4773 2033 4787 2047
rect 4773 1913 4787 1927
rect 4773 1893 4787 1907
rect 4773 1473 4787 1487
rect 4773 1433 4787 1447
rect 4773 1193 4787 1207
rect 4773 1153 4787 1167
rect 4753 1093 4767 1107
rect 4733 1073 4747 1087
rect 4653 1013 4667 1027
rect 4693 973 4707 987
rect 4753 1013 4767 1027
rect 4753 993 4767 1007
rect 4773 953 4787 967
rect 4753 913 4767 927
rect 4713 893 4727 907
rect 4733 893 4747 907
rect 4733 873 4747 887
rect 4653 853 4667 867
rect 4693 853 4707 867
rect 4613 833 4627 847
rect 4633 833 4647 847
rect 4653 833 4667 847
rect 4593 793 4607 807
rect 4613 793 4627 807
rect 4653 793 4667 807
rect 4633 773 4647 787
rect 4613 753 4627 767
rect 4593 693 4607 707
rect 4613 673 4627 687
rect 4593 653 4607 667
rect 4713 833 4727 847
rect 4753 853 4767 867
rect 4693 773 4707 787
rect 4673 753 4687 767
rect 4713 733 4727 747
rect 4673 713 4687 727
rect 4653 653 4667 667
rect 4713 653 4727 667
rect 4753 653 4767 667
rect 4633 613 4647 627
rect 4693 613 4707 627
rect 4733 633 4747 647
rect 4673 593 4687 607
rect 4573 373 4587 387
rect 4613 373 4627 387
rect 4433 353 4447 367
rect 4493 353 4507 367
rect 4533 353 4547 367
rect 4553 333 4567 347
rect 4593 353 4607 367
rect 4413 293 4427 307
rect 4233 213 4247 227
rect 4253 213 4267 227
rect 4393 213 4407 227
rect 4213 193 4227 207
rect 4153 173 4167 187
rect 4073 133 4087 147
rect 4093 113 4107 127
rect 4133 113 4147 127
rect 4153 113 4167 127
rect 4193 113 4207 127
rect 4473 193 4487 207
rect 4313 173 4327 187
rect 4393 173 4407 187
rect 4353 153 4367 167
rect 4253 133 4267 147
rect 4233 113 4247 127
rect 4293 113 4307 127
rect 4333 113 4347 127
rect 4553 313 4567 327
rect 4533 293 4547 307
rect 4593 293 4607 307
rect 4553 273 4567 287
rect 4573 273 4587 287
rect 4433 133 4447 147
rect 4413 113 4427 127
rect 4453 113 4467 127
rect 4513 133 4527 147
rect 4493 113 4507 127
rect 4593 113 4607 127
rect 4493 93 4507 107
rect 3973 33 3987 47
rect 4173 33 4187 47
rect 3793 13 3807 27
rect 4133 13 4147 27
rect 4653 353 4667 367
rect 4633 313 4647 327
rect 4753 573 4767 587
rect 4733 413 4747 427
rect 4653 253 4667 267
rect 4693 173 4707 187
rect 4673 133 4687 147
rect 4753 393 4767 407
rect 4773 173 4787 187
rect 4753 133 4767 147
rect 4213 13 4227 27
rect 4613 13 4627 27
<< metal3 >>
rect 327 4576 533 4584
rect 2807 4576 2873 4584
rect 447 4556 493 4564
rect 2707 4556 3153 4564
rect 747 4536 1133 4544
rect 2947 4536 3073 4544
rect 3087 4536 3933 4544
rect 427 4516 593 4524
rect 607 4516 993 4524
rect 1087 4516 1113 4524
rect 1287 4516 1413 4524
rect 3396 4516 3793 4524
rect 407 4496 453 4504
rect 507 4496 673 4504
rect 707 4496 733 4504
rect 907 4496 1233 4504
rect 1247 4496 1333 4504
rect 1347 4496 1593 4504
rect 1607 4496 1893 4504
rect 1907 4496 1913 4504
rect 2127 4496 2433 4504
rect 2467 4496 2533 4504
rect 2547 4496 2624 4504
rect 227 4476 244 4484
rect 147 4456 193 4464
rect 236 4464 244 4476
rect 267 4476 413 4484
rect 476 4467 484 4493
rect 667 4476 813 4484
rect 836 4476 1373 4484
rect 236 4456 333 4464
rect 836 4464 844 4476
rect 1487 4476 1673 4484
rect 1787 4476 1813 4484
rect 1947 4476 2073 4484
rect 2096 4476 2293 4484
rect 2096 4467 2104 4476
rect 2616 4484 2624 4496
rect 3227 4496 3293 4504
rect 3307 4496 3373 4504
rect 3396 4504 3404 4516
rect 3987 4516 4393 4524
rect 3396 4496 3433 4504
rect 2616 4476 2893 4484
rect 2907 4476 3013 4484
rect 3396 4484 3404 4496
rect 4067 4496 4133 4504
rect 4167 4496 4213 4504
rect 4447 4496 4553 4504
rect 3267 4476 3404 4484
rect 3427 4476 3604 4484
rect 767 4456 844 4464
rect 1007 4456 1053 4464
rect 1107 4456 1733 4464
rect 2416 4464 2424 4473
rect 2407 4456 2424 4464
rect 247 4436 353 4444
rect 367 4436 753 4444
rect 1027 4436 1393 4444
rect 1407 4436 1613 4444
rect 1627 4436 1713 4444
rect 167 4416 273 4424
rect 967 4416 1113 4424
rect 1467 4416 2173 4424
rect 127 4396 153 4404
rect 1687 4396 2053 4404
rect 2196 4404 2204 4453
rect 2227 4436 2353 4444
rect 2556 4444 2564 4473
rect 2596 4447 2604 4473
rect 2627 4456 2973 4464
rect 3407 4456 3473 4464
rect 3507 4456 3533 4464
rect 3596 4464 3604 4476
rect 3716 4484 3724 4493
rect 3627 4476 3724 4484
rect 3767 4476 3824 4484
rect 3816 4467 3824 4476
rect 3847 4476 3993 4484
rect 4047 4476 4084 4484
rect 3596 4456 3664 4464
rect 2367 4436 2564 4444
rect 3007 4436 3033 4444
rect 3367 4436 3553 4444
rect 3567 4436 3613 4444
rect 2956 4424 2964 4433
rect 2407 4416 3013 4424
rect 3236 4424 3244 4433
rect 3236 4416 3453 4424
rect 3467 4416 3633 4424
rect 3656 4424 3664 4456
rect 3687 4456 3733 4464
rect 3836 4456 3853 4464
rect 3836 4444 3844 4456
rect 3967 4456 4053 4464
rect 3687 4436 3844 4444
rect 4007 4436 4053 4444
rect 4076 4444 4084 4476
rect 4147 4476 4204 4484
rect 4196 4467 4204 4476
rect 4287 4456 4313 4464
rect 4467 4456 4573 4464
rect 4687 4456 4713 4464
rect 4076 4436 4113 4444
rect 4176 4444 4184 4453
rect 4176 4436 4233 4444
rect 4427 4436 4513 4444
rect 4667 4436 4753 4444
rect 3656 4416 3893 4424
rect 4156 4424 4164 4433
rect 4127 4416 4164 4424
rect 4247 4416 4393 4424
rect 4407 4416 4493 4424
rect 4556 4424 4564 4433
rect 4547 4416 4564 4424
rect 2196 4396 2213 4404
rect 2327 4396 2513 4404
rect 2527 4396 2573 4404
rect 3167 4396 3313 4404
rect 3327 4396 3493 4404
rect 3527 4396 3573 4404
rect 3587 4396 3693 4404
rect 4227 4396 4293 4404
rect 4347 4396 4733 4404
rect 2067 4376 2253 4384
rect 2267 4376 2633 4384
rect 3227 4376 3333 4384
rect 4107 4376 4593 4384
rect 2427 4356 3193 4364
rect 4107 4356 4713 4364
rect 1807 4336 2013 4344
rect 4467 4336 4493 4344
rect 907 4316 1013 4324
rect 2447 4316 2853 4324
rect 2827 4296 2913 4304
rect 2947 4296 2993 4304
rect 3207 4296 3833 4304
rect 2727 4276 3253 4284
rect 3267 4276 3273 4284
rect 3387 4276 3513 4284
rect 3567 4276 3993 4284
rect 4147 4276 4193 4284
rect 507 4256 533 4264
rect 2347 4256 2413 4264
rect 2867 4256 3113 4264
rect 3127 4256 3733 4264
rect 4307 4256 4413 4264
rect 347 4236 533 4244
rect 547 4236 693 4244
rect 2356 4236 2393 4244
rect 167 4216 173 4224
rect 187 4216 433 4224
rect 447 4216 473 4224
rect 787 4216 833 4224
rect 936 4216 1013 4224
rect 287 4196 333 4204
rect 387 4196 473 4204
rect 487 4196 573 4204
rect 587 4196 633 4204
rect 747 4196 813 4204
rect 936 4204 944 4216
rect 1127 4216 1193 4224
rect 1367 4216 1793 4224
rect 2107 4216 2124 4224
rect 927 4196 944 4204
rect 967 4196 993 4204
rect 1207 4196 1313 4204
rect 1327 4196 1573 4204
rect 2116 4204 2124 4216
rect 2147 4216 2233 4224
rect 2356 4224 2364 4236
rect 2536 4236 2824 4244
rect 2336 4216 2364 4224
rect 1967 4196 2293 4204
rect 76 4184 84 4193
rect 76 4176 133 4184
rect 187 4176 213 4184
rect 267 4176 313 4184
rect 687 4176 793 4184
rect 927 4176 1093 4184
rect 1267 4176 1373 4184
rect 1507 4176 1633 4184
rect 2147 4176 2233 4184
rect 2247 4176 2273 4184
rect 2336 4184 2344 4216
rect 2536 4224 2544 4236
rect 2387 4216 2544 4224
rect 2567 4216 2633 4224
rect 2816 4224 2824 4236
rect 2907 4236 3033 4244
rect 3047 4236 3933 4244
rect 3947 4236 4013 4244
rect 4256 4236 4273 4244
rect 2816 4216 3033 4224
rect 3087 4216 3273 4224
rect 3427 4216 3473 4224
rect 3567 4216 3613 4224
rect 3676 4216 3793 4224
rect 2327 4176 2344 4184
rect 2376 4184 2384 4213
rect 2576 4196 2593 4204
rect 2367 4176 2384 4184
rect 207 4156 253 4164
rect 467 4156 553 4164
rect 567 4156 593 4164
rect 627 4156 713 4164
rect 827 4156 933 4164
rect 987 4156 1053 4164
rect 1067 4156 1233 4164
rect 1267 4156 1293 4164
rect 1347 4156 1453 4164
rect 1747 4156 1773 4164
rect 1787 4156 1813 4164
rect 2127 4156 2153 4164
rect 2187 4156 2393 4164
rect 2516 4164 2524 4193
rect 2576 4187 2584 4196
rect 2827 4196 2904 4204
rect 2676 4167 2684 4193
rect 2516 4156 2593 4164
rect 107 4136 233 4144
rect 667 4136 1244 4144
rect 47 4116 93 4124
rect 207 4116 273 4124
rect 287 4116 1213 4124
rect 1236 4124 1244 4136
rect 1627 4136 1973 4144
rect 2267 4136 2473 4144
rect 2607 4136 2653 4144
rect 2776 4144 2784 4193
rect 2796 4184 2804 4193
rect 2796 4176 2873 4184
rect 2896 4184 2904 4196
rect 2927 4196 2953 4204
rect 3067 4196 3133 4204
rect 3156 4196 3213 4204
rect 2896 4176 2913 4184
rect 3156 4184 3164 4196
rect 3267 4196 3293 4204
rect 3427 4196 3653 4204
rect 3676 4204 3684 4216
rect 3667 4196 3684 4204
rect 3707 4196 3753 4204
rect 3987 4196 4053 4204
rect 4176 4196 4193 4204
rect 3107 4176 3164 4184
rect 3447 4176 3473 4184
rect 3647 4176 3733 4184
rect 3747 4176 3804 4184
rect 2807 4156 2893 4164
rect 3247 4156 3433 4164
rect 3447 4156 3453 4164
rect 3527 4156 3673 4164
rect 3687 4156 3773 4164
rect 3796 4164 3804 4176
rect 3876 4184 3884 4193
rect 3827 4176 3884 4184
rect 4176 4184 4184 4196
rect 4147 4176 4184 4184
rect 4216 4184 4224 4233
rect 4207 4176 4224 4184
rect 3796 4156 3913 4164
rect 3927 4156 3953 4164
rect 4087 4156 4153 4164
rect 4236 4164 4244 4213
rect 4256 4187 4264 4236
rect 4287 4216 4533 4224
rect 4556 4216 4593 4224
rect 4487 4196 4533 4204
rect 4316 4184 4324 4193
rect 4287 4176 4324 4184
rect 4187 4156 4273 4164
rect 2776 4136 2973 4144
rect 3547 4136 3653 4144
rect 3667 4136 3693 4144
rect 3907 4136 4213 4144
rect 4227 4136 4233 4144
rect 4356 4144 4364 4193
rect 4436 4184 4444 4193
rect 4387 4176 4444 4184
rect 4556 4184 4564 4216
rect 4707 4216 4773 4224
rect 4587 4196 4633 4204
rect 4527 4176 4564 4184
rect 4547 4156 4593 4164
rect 4247 4136 4364 4144
rect 4527 4136 4633 4144
rect 1236 4116 1713 4124
rect 2547 4116 2753 4124
rect 3407 4116 3493 4124
rect 3547 4116 3633 4124
rect 4167 4116 4353 4124
rect 4567 4116 4653 4124
rect 187 4096 213 4104
rect 227 4096 353 4104
rect 367 4096 393 4104
rect 927 4096 1013 4104
rect 1047 4096 1133 4104
rect 1667 4096 2493 4104
rect 2707 4096 2733 4104
rect 2907 4096 3193 4104
rect 3607 4096 4033 4104
rect 4087 4096 4293 4104
rect 4347 4096 4493 4104
rect 4567 4096 4613 4104
rect 587 4076 753 4084
rect 767 4076 1124 4084
rect 267 4056 1093 4064
rect 1116 4064 1124 4076
rect 1287 4076 1833 4084
rect 2347 4076 2553 4084
rect 2627 4076 2893 4084
rect 2987 4076 3244 4084
rect 1116 4056 1373 4064
rect 1887 4056 2133 4064
rect 2667 4056 2784 4064
rect 307 4036 333 4044
rect 407 4036 473 4044
rect 527 4036 593 4044
rect 807 4036 853 4044
rect 987 4036 1013 4044
rect 1047 4036 1193 4044
rect 1467 4036 1473 4044
rect 1487 4036 1693 4044
rect 2187 4036 2533 4044
rect 2727 4036 2753 4044
rect 2776 4044 2784 4056
rect 2847 4056 2973 4064
rect 3236 4064 3244 4076
rect 3487 4076 3553 4084
rect 3567 4076 3853 4084
rect 3876 4076 4673 4084
rect 3876 4064 3884 4076
rect 3236 4056 3884 4064
rect 4127 4056 4233 4064
rect 2776 4036 3193 4044
rect 3627 4036 3753 4044
rect 3847 4036 4033 4044
rect 4147 4036 4313 4044
rect 27 4016 293 4024
rect 467 4016 513 4024
rect 536 4016 653 4024
rect 536 4007 544 4016
rect 727 4016 993 4024
rect 1016 4016 1033 4024
rect 16 3996 53 4004
rect 16 3947 24 3996
rect 127 3996 184 4004
rect 76 3976 133 3984
rect 56 3944 64 3973
rect 76 3967 84 3976
rect 176 3984 184 3996
rect 207 3996 284 4004
rect 276 3987 284 3996
rect 507 3996 524 4004
rect 176 3976 213 3984
rect 327 3976 373 3984
rect 516 3984 524 3996
rect 607 3996 624 4004
rect 516 3976 573 3984
rect 616 3984 624 3996
rect 707 3996 733 4004
rect 827 3996 893 4004
rect 1016 4004 1024 4016
rect 1096 4016 1273 4024
rect 1007 3996 1024 4004
rect 1096 4004 1104 4016
rect 1487 4016 1673 4024
rect 1847 4016 1893 4024
rect 2127 4016 2213 4024
rect 2287 4016 2333 4024
rect 2487 4016 2513 4024
rect 2527 4016 2744 4024
rect 1087 3996 1104 4004
rect 1127 3996 1144 4004
rect 1136 3987 1144 3996
rect 1247 3996 1573 4004
rect 1296 3987 1304 3996
rect 1667 3996 1793 4004
rect 1907 3996 2013 4004
rect 2067 3996 2353 4004
rect 2396 4004 2404 4013
rect 2396 3996 2493 4004
rect 2556 3996 2673 4004
rect 2556 3987 2564 3996
rect 2687 3996 2713 4004
rect 2736 4004 2744 4016
rect 2767 4016 2904 4024
rect 2736 3996 2873 4004
rect 616 3976 673 3984
rect 727 3976 773 3984
rect 887 3976 933 3984
rect 987 3976 1013 3984
rect 1447 3976 1493 3984
rect 1647 3976 1713 3984
rect 1827 3976 1913 3984
rect 2047 3976 2093 3984
rect 2327 3976 2373 3984
rect 2387 3976 2453 3984
rect 2647 3976 2733 3984
rect 2876 3984 2884 3993
rect 2767 3976 2884 3984
rect 127 3956 613 3964
rect 847 3956 973 3964
rect 1607 3956 1673 3964
rect 1747 3956 1933 3964
rect 1996 3947 2004 3973
rect 2307 3956 2344 3964
rect 56 3936 233 3944
rect 607 3936 773 3944
rect 927 3936 1073 3944
rect 1827 3936 1953 3944
rect 2196 3944 2204 3953
rect 2196 3936 2253 3944
rect 2336 3944 2344 3956
rect 2467 3956 2593 3964
rect 2667 3956 2773 3964
rect 2896 3964 2904 4016
rect 2967 4016 3093 4024
rect 3187 4016 3213 4024
rect 3247 4016 3273 4024
rect 3327 4016 3513 4024
rect 3527 4016 3573 4024
rect 3616 4016 3673 4024
rect 2916 3987 2924 4013
rect 2947 3996 3053 4004
rect 3167 3996 3353 4004
rect 3367 3996 3404 4004
rect 3087 3976 3104 3984
rect 2896 3956 3013 3964
rect 2336 3936 2493 3944
rect 2507 3936 2793 3944
rect 2607 3916 2873 3924
rect 3036 3924 3044 3973
rect 3096 3964 3104 3976
rect 3127 3976 3253 3984
rect 3347 3976 3373 3984
rect 3096 3956 3333 3964
rect 3396 3964 3404 3996
rect 3427 3996 3473 4004
rect 3616 3984 3624 4016
rect 4187 4016 4253 4024
rect 4287 4016 4393 4024
rect 4627 4016 4673 4024
rect 3647 3996 3673 4004
rect 3716 4004 3724 4013
rect 3716 3996 3793 4004
rect 3716 3987 3724 3996
rect 4116 3996 4133 4004
rect 3616 3976 3644 3984
rect 3387 3956 3404 3964
rect 3416 3964 3424 3973
rect 3636 3967 3644 3976
rect 3747 3976 3813 3984
rect 3836 3976 3893 3984
rect 3416 3956 3453 3964
rect 3467 3956 3593 3964
rect 3667 3956 3773 3964
rect 3836 3964 3844 3976
rect 3916 3976 3973 3984
rect 3796 3956 3844 3964
rect 3056 3944 3064 3953
rect 3056 3936 3113 3944
rect 3127 3936 3173 3944
rect 3207 3936 3293 3944
rect 3307 3936 3393 3944
rect 3796 3944 3804 3956
rect 3916 3964 3924 3976
rect 4116 3967 4124 3996
rect 4236 3996 4273 4004
rect 4187 3976 4224 3984
rect 3887 3956 3924 3964
rect 4136 3947 4144 3973
rect 4167 3956 4184 3964
rect 3427 3936 3804 3944
rect 3967 3936 4073 3944
rect 3036 3916 3453 3924
rect 3527 3916 3573 3924
rect 3587 3916 3613 3924
rect 3747 3916 3793 3924
rect 4176 3924 4184 3956
rect 4216 3947 4224 3976
rect 4236 3964 4244 3996
rect 4287 3996 4293 4004
rect 4467 3996 4633 4004
rect 4647 3996 4704 4004
rect 4696 3987 4704 3996
rect 4267 3976 4313 3984
rect 4427 3976 4493 3984
rect 4607 3976 4653 3984
rect 4236 3956 4253 3964
rect 4176 3916 4453 3924
rect 4516 3924 4524 3953
rect 4536 3947 4544 3973
rect 4627 3956 4693 3964
rect 4727 3956 4753 3964
rect 4567 3936 4753 3944
rect 4516 3916 4553 3924
rect 2347 3896 2413 3904
rect 2427 3896 2613 3904
rect 3107 3896 3413 3904
rect 3707 3896 3813 3904
rect 3827 3896 3853 3904
rect 3927 3896 4053 3904
rect 4067 3896 4473 3904
rect 3247 3876 3293 3884
rect 4027 3876 4573 3884
rect 2967 3856 2993 3864
rect 4407 3856 4433 3864
rect 2807 3836 2993 3844
rect 4167 3836 4733 3844
rect 227 3816 253 3824
rect 427 3816 913 3824
rect 4107 3816 4473 3824
rect 4667 3816 4733 3824
rect 487 3796 593 3804
rect 2867 3796 2973 3804
rect 4147 3796 4173 3804
rect 447 3776 553 3784
rect 2567 3776 2693 3784
rect 2887 3776 2973 3784
rect 487 3756 533 3764
rect 547 3756 673 3764
rect 2367 3756 2433 3764
rect 2467 3756 3093 3764
rect 3607 3756 3753 3764
rect 496 3736 553 3744
rect 87 3716 413 3724
rect 496 3707 504 3736
rect 787 3736 813 3744
rect 827 3736 1053 3744
rect 1187 3736 1373 3744
rect 1467 3736 1533 3744
rect 1556 3727 1564 3753
rect 2187 3736 2373 3744
rect 2276 3727 2284 3736
rect 2427 3736 2573 3744
rect 2636 3736 2693 3744
rect 2636 3727 2644 3736
rect 2707 3736 2833 3744
rect 2847 3736 2933 3744
rect 3047 3736 3193 3744
rect 3387 3736 3424 3744
rect 967 3716 1173 3724
rect 1427 3716 1473 3724
rect 2047 3716 2113 3724
rect 2447 3716 2493 3724
rect 2807 3716 2913 3724
rect 2967 3716 3004 3724
rect 67 3696 313 3704
rect 687 3696 813 3704
rect 1267 3696 1393 3704
rect 1527 3696 1573 3704
rect 2267 3696 2293 3704
rect 2316 3704 2324 3713
rect 2316 3696 2473 3704
rect 2656 3704 2664 3713
rect 2996 3707 3004 3716
rect 3067 3716 3113 3724
rect 3187 3716 3233 3724
rect 3267 3716 3293 3724
rect 3356 3716 3393 3724
rect 2607 3696 2664 3704
rect 2747 3696 2773 3704
rect 3156 3704 3164 3713
rect 3027 3696 3173 3704
rect 27 3676 393 3684
rect 927 3676 1213 3684
rect 1367 3676 1393 3684
rect 1407 3676 1433 3684
rect 2147 3676 2173 3684
rect 2427 3676 2513 3684
rect 2627 3676 2673 3684
rect 2687 3676 2813 3684
rect 2827 3676 2853 3684
rect 2987 3676 3013 3684
rect 3067 3676 3113 3684
rect 3356 3684 3364 3716
rect 3416 3707 3424 3736
rect 3507 3736 3533 3744
rect 3387 3696 3404 3704
rect 3356 3676 3373 3684
rect 627 3656 713 3664
rect 1607 3656 1713 3664
rect 2407 3656 2573 3664
rect 2607 3656 2973 3664
rect 3047 3656 3133 3664
rect 3396 3664 3404 3696
rect 3456 3704 3464 3733
rect 3556 3724 3564 3753
rect 3647 3736 3733 3744
rect 4327 3736 4393 3744
rect 4607 3736 4653 3744
rect 4667 3736 4773 3744
rect 3487 3716 3564 3724
rect 3456 3696 3493 3704
rect 3576 3704 3584 3733
rect 3707 3716 3753 3724
rect 3787 3716 3833 3724
rect 3847 3716 3873 3724
rect 3987 3716 4033 3724
rect 4047 3716 4093 3724
rect 4227 3716 4273 3724
rect 4367 3716 4413 3724
rect 4507 3716 4613 3724
rect 4627 3716 4653 3724
rect 3576 3696 3633 3704
rect 3656 3704 3664 3713
rect 3656 3696 3773 3704
rect 3807 3696 3884 3704
rect 3687 3676 3793 3684
rect 3827 3676 3853 3684
rect 3876 3684 3884 3696
rect 3916 3687 3924 3713
rect 3947 3696 3993 3704
rect 4176 3704 4184 3713
rect 4127 3696 4184 3704
rect 3876 3676 3893 3684
rect 4067 3676 4153 3684
rect 4196 3684 4204 3713
rect 4267 3696 4293 3704
rect 4336 3704 4344 3713
rect 4316 3696 4344 3704
rect 4187 3676 4204 3684
rect 4316 3684 4324 3696
rect 4707 3696 4733 3704
rect 4247 3676 4324 3684
rect 4347 3676 4373 3684
rect 4587 3676 4673 3684
rect 4687 3676 4733 3684
rect 3187 3656 3404 3664
rect 3427 3656 3673 3664
rect 3787 3656 3953 3664
rect 4027 3656 4413 3664
rect 1147 3636 1333 3644
rect 1347 3636 1793 3644
rect 1807 3636 1813 3644
rect 2107 3636 2153 3644
rect 2167 3636 2353 3644
rect 2367 3636 3413 3644
rect 3827 3636 3953 3644
rect 4207 3636 4253 3644
rect 4267 3636 4453 3644
rect 4507 3636 4753 3644
rect 167 3616 273 3624
rect 1767 3616 1793 3624
rect 2407 3616 2493 3624
rect 2567 3616 2613 3624
rect 2767 3616 2813 3624
rect 3027 3616 3093 3624
rect 3327 3616 3353 3624
rect 3367 3616 3473 3624
rect 3727 3616 3813 3624
rect 3867 3616 4093 3624
rect 4227 3616 4593 3624
rect 4707 3616 4753 3624
rect 807 3596 1093 3604
rect 2067 3596 2193 3604
rect 2207 3596 2653 3604
rect 2967 3596 3153 3604
rect 3187 3596 3393 3604
rect 4007 3596 4233 3604
rect 967 3576 1693 3584
rect 1987 3576 2053 3584
rect 2167 3576 2453 3584
rect 2587 3576 2933 3584
rect 2987 3576 3093 3584
rect 3107 3576 3313 3584
rect 3347 3576 3533 3584
rect 3767 3576 4033 3584
rect 4627 3576 4673 3584
rect 4687 3576 4773 3584
rect 667 3556 753 3564
rect 767 3556 853 3564
rect 867 3556 973 3564
rect 1167 3556 1433 3564
rect 2147 3556 2333 3564
rect 2347 3556 2393 3564
rect 2467 3556 2753 3564
rect 2907 3556 3213 3564
rect 3247 3556 3364 3564
rect 527 3536 813 3544
rect 887 3536 933 3544
rect 1007 3536 1253 3544
rect 1276 3536 1333 3544
rect 107 3516 373 3524
rect 587 3516 613 3524
rect 656 3516 673 3524
rect 307 3496 353 3504
rect 416 3504 424 3513
rect 656 3507 664 3516
rect 716 3516 773 3524
rect 396 3496 424 3504
rect 436 3496 473 3504
rect 227 3476 313 3484
rect 396 3464 404 3496
rect 436 3484 444 3496
rect 607 3496 633 3504
rect 427 3476 444 3484
rect 467 3476 533 3484
rect 287 3456 413 3464
rect 556 3444 564 3493
rect 716 3487 724 3516
rect 1007 3516 1033 3524
rect 1276 3524 1284 3536
rect 1847 3536 1993 3544
rect 2247 3536 2293 3544
rect 2387 3536 2413 3544
rect 2447 3536 2773 3544
rect 2807 3536 2853 3544
rect 2927 3536 2973 3544
rect 2987 3536 3013 3544
rect 3047 3536 3333 3544
rect 3356 3544 3364 3556
rect 3387 3556 3553 3564
rect 3727 3556 3853 3564
rect 4047 3556 4153 3564
rect 4387 3556 4424 3564
rect 3356 3536 3613 3544
rect 3627 3536 3633 3544
rect 4147 3536 4193 3544
rect 4207 3536 4293 3544
rect 4416 3544 4424 3556
rect 4467 3556 4784 3564
rect 4416 3536 4493 3544
rect 1056 3516 1284 3524
rect 747 3496 773 3504
rect 847 3496 933 3504
rect 1056 3504 1064 3516
rect 1407 3516 1473 3524
rect 1487 3516 1593 3524
rect 1607 3516 1964 3524
rect 947 3496 1064 3504
rect 1307 3496 1413 3504
rect 1467 3496 1513 3504
rect 1707 3496 1833 3504
rect 1956 3504 1964 3516
rect 2047 3516 2173 3524
rect 2567 3516 2633 3524
rect 2656 3516 2813 3524
rect 1956 3496 1973 3504
rect 2027 3496 2093 3504
rect 2207 3496 2333 3504
rect 2527 3496 2593 3504
rect 587 3476 673 3484
rect 827 3476 913 3484
rect 1987 3476 2073 3484
rect 2247 3476 2313 3484
rect 2327 3476 2433 3484
rect 2487 3476 2533 3484
rect 2636 3484 2644 3493
rect 2596 3476 2644 3484
rect 2656 3484 2664 3516
rect 2847 3516 2873 3524
rect 2887 3516 2993 3524
rect 3136 3516 3213 3524
rect 3136 3507 3144 3516
rect 3267 3516 3353 3524
rect 3376 3516 3393 3524
rect 2687 3496 2733 3504
rect 2967 3496 3013 3504
rect 2656 3476 2673 3484
rect 2596 3467 2604 3476
rect 2776 3484 2784 3493
rect 2767 3476 2784 3484
rect 2927 3476 2973 3484
rect 687 3456 893 3464
rect 1087 3456 1313 3464
rect 1327 3456 1613 3464
rect 2067 3456 2113 3464
rect 2127 3456 2273 3464
rect 2867 3456 2993 3464
rect 3007 3456 3193 3464
rect 3376 3464 3384 3516
rect 3427 3516 3464 3524
rect 3407 3496 3433 3504
rect 3456 3484 3464 3516
rect 3767 3516 3793 3524
rect 3927 3516 3944 3524
rect 3496 3504 3504 3513
rect 3496 3496 3553 3504
rect 3936 3504 3944 3516
rect 4136 3516 4213 3524
rect 3607 3496 3944 3504
rect 3936 3487 3944 3496
rect 3427 3476 3464 3484
rect 3507 3476 3733 3484
rect 3376 3456 3393 3464
rect 3407 3456 3453 3464
rect 3496 3456 3573 3464
rect 3496 3447 3504 3456
rect 4056 3464 4064 3513
rect 4136 3487 4144 3516
rect 4287 3516 4304 3524
rect 4236 3496 4253 3504
rect 4236 3484 4244 3496
rect 4227 3476 4244 3484
rect 4056 3456 4113 3464
rect 4187 3456 4213 3464
rect 556 3436 753 3444
rect 1387 3436 1673 3444
rect 1687 3436 1933 3444
rect 2747 3436 3033 3444
rect 3127 3436 3413 3444
rect 4087 3436 4153 3444
rect 1547 3416 1593 3424
rect 2907 3416 3473 3424
rect 3527 3416 3593 3424
rect 3667 3416 3793 3424
rect 3807 3416 4013 3424
rect 4027 3416 4073 3424
rect 4256 3424 4264 3473
rect 4276 3444 4284 3493
rect 4296 3467 4304 3516
rect 4327 3516 4373 3524
rect 4396 3507 4404 3533
rect 4336 3464 4344 3493
rect 4367 3476 4433 3484
rect 4456 3484 4464 3536
rect 4567 3536 4653 3544
rect 4516 3516 4573 3524
rect 4447 3476 4464 3484
rect 4476 3484 4484 3513
rect 4516 3504 4524 3516
rect 4607 3516 4693 3524
rect 4507 3496 4524 3504
rect 4547 3496 4633 3504
rect 4696 3484 4704 3493
rect 4476 3476 4544 3484
rect 4336 3456 4353 3464
rect 4427 3456 4513 3464
rect 4536 3464 4544 3476
rect 4676 3476 4704 3484
rect 4536 3456 4653 3464
rect 4676 3447 4684 3476
rect 4716 3464 4724 3513
rect 4707 3456 4724 3464
rect 4276 3436 4353 3444
rect 4507 3436 4573 3444
rect 4727 3436 4753 3444
rect 4256 3416 4373 3424
rect 4647 3416 4733 3424
rect 2847 3396 3553 3404
rect 3667 3396 3733 3404
rect 4007 3396 4273 3404
rect 4387 3396 4753 3404
rect 3107 3376 3293 3384
rect 3347 3376 3613 3384
rect 3987 3376 4053 3384
rect 4067 3376 4233 3384
rect 4776 3384 4784 3556
rect 4747 3376 4784 3384
rect 2827 3356 3393 3364
rect 3407 3356 3433 3364
rect 3467 3356 4413 3364
rect 1267 3336 2053 3344
rect 2067 3336 3113 3344
rect 3167 3336 3273 3344
rect 3307 3336 3653 3344
rect 3767 3336 3893 3344
rect 4067 3336 4093 3344
rect 4147 3336 4593 3344
rect 2307 3316 2413 3324
rect 2667 3316 3233 3324
rect 3407 3316 3493 3324
rect 3507 3316 3913 3324
rect 127 3296 253 3304
rect 2267 3296 3053 3304
rect 3187 3296 3373 3304
rect 3467 3296 3544 3304
rect 267 3276 333 3284
rect 447 3276 533 3284
rect 587 3276 613 3284
rect 1667 3276 1913 3284
rect 2207 3276 2213 3284
rect 2227 3276 2313 3284
rect 2816 3276 2873 3284
rect 227 3256 293 3264
rect 307 3256 373 3264
rect 487 3256 544 3264
rect 407 3236 513 3244
rect 536 3244 544 3256
rect 607 3256 633 3264
rect 1927 3256 1953 3264
rect 2456 3256 2653 3264
rect 536 3236 693 3244
rect 967 3236 1013 3244
rect 1027 3236 1053 3244
rect 1227 3236 1513 3244
rect 1736 3244 1744 3253
rect 2456 3247 2464 3256
rect 2716 3256 2753 3264
rect 1627 3236 1744 3244
rect 1767 3236 1813 3244
rect 1827 3236 1853 3244
rect 1867 3236 2013 3244
rect 2387 3236 2444 3244
rect 107 3216 493 3224
rect 1236 3216 1273 3224
rect 1236 3207 1244 3216
rect 1647 3216 1713 3224
rect 1907 3216 1973 3224
rect 2087 3216 2113 3224
rect 2436 3224 2444 3236
rect 2576 3236 2633 3244
rect 2436 3216 2493 3224
rect 2556 3207 2564 3233
rect 747 3196 773 3204
rect 1707 3196 1733 3204
rect 2007 3196 2193 3204
rect 807 3176 1353 3184
rect 1407 3176 1533 3184
rect 1567 3176 1693 3184
rect 1887 3176 2113 3184
rect 2487 3176 2533 3184
rect 2576 3184 2584 3236
rect 2667 3236 2693 3244
rect 2716 3227 2724 3256
rect 2736 3204 2744 3233
rect 2667 3196 2744 3204
rect 2796 3204 2804 3233
rect 2816 3227 2824 3276
rect 3047 3276 3113 3284
rect 3367 3276 3413 3284
rect 3427 3276 3513 3284
rect 3536 3284 3544 3296
rect 3567 3296 3633 3304
rect 3647 3296 3773 3304
rect 3796 3296 4033 3304
rect 3536 3276 3733 3284
rect 3796 3284 3804 3296
rect 4207 3296 4393 3304
rect 4747 3296 4764 3304
rect 3747 3276 3804 3284
rect 4007 3276 4173 3284
rect 4307 3276 4333 3284
rect 4487 3276 4544 3284
rect 2927 3236 2973 3244
rect 3016 3244 3024 3273
rect 3136 3256 3193 3264
rect 3016 3236 3053 3244
rect 2836 3216 2893 3224
rect 2836 3204 2844 3216
rect 3136 3224 3144 3256
rect 3227 3256 3273 3264
rect 3807 3256 3844 3264
rect 3187 3236 3213 3244
rect 3316 3244 3324 3253
rect 3267 3236 3333 3244
rect 3087 3216 3144 3224
rect 3156 3207 3164 3233
rect 3176 3216 3353 3224
rect 3176 3207 3184 3216
rect 3436 3224 3444 3253
rect 3496 3244 3504 3253
rect 3496 3236 3524 3244
rect 3436 3216 3493 3224
rect 3516 3224 3524 3236
rect 3547 3236 3573 3244
rect 3616 3227 3624 3253
rect 3516 3216 3573 3224
rect 3676 3224 3684 3253
rect 3787 3236 3813 3244
rect 3836 3227 3844 3256
rect 3856 3247 3864 3273
rect 3907 3256 3924 3264
rect 3876 3227 3884 3253
rect 3916 3244 3924 3256
rect 3947 3256 3964 3264
rect 3956 3247 3964 3256
rect 4067 3256 4113 3264
rect 4227 3256 4293 3264
rect 4447 3256 4524 3264
rect 3916 3236 3944 3244
rect 3936 3227 3944 3236
rect 3967 3236 4013 3244
rect 4156 3244 4164 3253
rect 4156 3236 4184 3244
rect 4176 3227 4184 3236
rect 3676 3216 3753 3224
rect 3987 3216 4113 3224
rect 4127 3216 4153 3224
rect 2796 3196 2844 3204
rect 2867 3196 2933 3204
rect 2967 3196 3013 3204
rect 3307 3196 3413 3204
rect 3427 3196 3673 3204
rect 3687 3196 3693 3204
rect 3707 3196 3713 3204
rect 3807 3196 3973 3204
rect 4216 3204 4224 3253
rect 4296 3236 4353 3244
rect 4296 3227 4304 3236
rect 4416 3244 4424 3253
rect 4516 3247 4524 3256
rect 4416 3236 4433 3244
rect 4376 3224 4384 3233
rect 4327 3216 4384 3224
rect 4476 3224 4484 3233
rect 4427 3216 4484 3224
rect 4536 3224 4544 3276
rect 4707 3276 4744 3284
rect 4607 3256 4624 3264
rect 4556 3227 4564 3253
rect 4616 3247 4624 3256
rect 4667 3256 4713 3264
rect 4736 3247 4744 3276
rect 4647 3236 4713 3244
rect 4507 3216 4544 3224
rect 4027 3196 4224 3204
rect 4327 3196 4373 3204
rect 4576 3204 4584 3233
rect 4756 3224 4764 3296
rect 4707 3216 4764 3224
rect 4427 3196 4584 3204
rect 4627 3196 4773 3204
rect 2547 3176 2584 3184
rect 2687 3176 2713 3184
rect 2747 3176 2773 3184
rect 2847 3176 3453 3184
rect 3487 3176 3893 3184
rect 4107 3176 4133 3184
rect 4147 3176 4253 3184
rect 4347 3176 4453 3184
rect 4587 3176 4653 3184
rect 367 3156 693 3164
rect 1187 3156 1873 3164
rect 2047 3156 2153 3164
rect 2567 3156 2573 3164
rect 2587 3156 2793 3164
rect 3067 3156 3153 3164
rect 3227 3156 3373 3164
rect 3787 3156 3813 3164
rect 4207 3156 4533 3164
rect 267 3136 333 3144
rect 407 3136 613 3144
rect 1507 3136 1773 3144
rect 2387 3136 2833 3144
rect 2847 3136 3053 3144
rect 3067 3136 3273 3144
rect 3287 3136 3533 3144
rect 3607 3136 3713 3144
rect 4187 3136 4333 3144
rect 4447 3136 4513 3144
rect 267 3116 273 3124
rect 287 3116 1833 3124
rect 2407 3116 2633 3124
rect 2647 3116 2753 3124
rect 2767 3116 3093 3124
rect 3187 3116 3313 3124
rect 3347 3116 3433 3124
rect 3667 3116 3753 3124
rect 4147 3116 4273 3124
rect 4327 3116 4753 3124
rect 147 3096 533 3104
rect 1107 3096 1433 3104
rect 1487 3096 1573 3104
rect 2427 3096 2473 3104
rect 2487 3096 2513 3104
rect 2567 3096 2673 3104
rect 3087 3096 3193 3104
rect 3227 3096 3613 3104
rect 3707 3096 3833 3104
rect 4567 3096 4653 3104
rect 767 3076 1173 3084
rect 1367 3076 1453 3084
rect 1667 3076 1953 3084
rect 2307 3076 2593 3084
rect 2667 3076 2693 3084
rect 2707 3076 2993 3084
rect 3027 3076 3173 3084
rect 3396 3076 3433 3084
rect 287 3056 313 3064
rect 987 3056 1033 3064
rect 1047 3056 1193 3064
rect 1347 3056 1613 3064
rect 1647 3056 1673 3064
rect 1687 3056 1733 3064
rect 1747 3056 1813 3064
rect 1827 3056 1933 3064
rect 2007 3056 2213 3064
rect 2247 3056 2433 3064
rect 2607 3056 2753 3064
rect 2787 3056 2924 3064
rect -24 3036 93 3044
rect -24 2996 -16 3036
rect 127 3036 293 3044
rect 296 3016 313 3024
rect 296 3004 304 3016
rect 187 2996 304 3004
rect 336 3004 344 3053
rect 547 3036 793 3044
rect 967 3036 993 3044
rect 1007 3036 1133 3044
rect 1307 3036 1413 3044
rect 1547 3036 1593 3044
rect 1736 3036 1773 3044
rect 1107 3016 1144 3024
rect 1136 3007 1144 3016
rect 1287 3016 1333 3024
rect 1736 3007 1744 3036
rect 1836 3036 1853 3044
rect 327 2996 344 3004
rect 427 2996 453 3004
rect 967 2996 1073 3004
rect 1836 3004 1844 3036
rect 1887 3036 2073 3044
rect 2347 3036 2384 3044
rect 1867 3016 1924 3024
rect 1916 3007 1924 3016
rect 2227 3016 2353 3024
rect 1787 2996 1893 3004
rect 2376 3004 2384 3036
rect 2456 3036 2593 3044
rect 2456 3027 2464 3036
rect 2696 3036 2713 3044
rect 2507 3016 2553 3024
rect 2587 3016 2673 3024
rect 2376 2996 2533 3004
rect 2696 3004 2704 3036
rect 2747 3036 2813 3044
rect 2856 3036 2893 3044
rect 2727 3016 2813 3024
rect 2836 3007 2844 3033
rect 2696 2996 2773 3004
rect 127 2976 353 2984
rect 987 2976 1113 2984
rect 1847 2976 1953 2984
rect 2147 2976 2253 2984
rect 2576 2984 2584 2993
rect 2527 2976 2584 2984
rect 2856 2984 2864 3036
rect 2916 3024 2924 3056
rect 2976 3056 3033 3064
rect 2976 3027 2984 3056
rect 3396 3064 3404 3076
rect 3487 3076 3844 3084
rect 3047 3056 3404 3064
rect 3427 3056 3464 3064
rect 3047 3036 3084 3044
rect 2907 3016 2924 3024
rect 3027 3016 3053 3024
rect 3076 3024 3084 3036
rect 3167 3036 3273 3044
rect 3076 3016 3253 3024
rect 3276 3024 3284 3033
rect 3276 3016 3304 3024
rect 2887 2996 3073 3004
rect 3296 3004 3304 3016
rect 3296 2996 3313 3004
rect 3456 3004 3464 3056
rect 3567 3056 3813 3064
rect 3836 3064 3844 3076
rect 3887 3076 4064 3084
rect 3836 3056 4033 3064
rect 3587 3036 3744 3044
rect 3607 3016 3673 3024
rect 3736 3024 3744 3036
rect 3807 3036 3833 3044
rect 3687 3016 3724 3024
rect 3736 3016 3804 3024
rect 3387 2996 3464 3004
rect 3507 2996 3573 3004
rect 3647 2996 3673 3004
rect 3716 3004 3724 3016
rect 3796 3004 3804 3016
rect 3716 2996 3784 3004
rect 3796 2996 3813 3004
rect 2856 2976 2893 2984
rect 2927 2976 2973 2984
rect 3107 2976 3753 2984
rect 3776 2984 3784 2996
rect 3856 3004 3864 3056
rect 3887 3036 3933 3044
rect 4027 3036 4044 3044
rect 3967 3016 3973 3024
rect 3987 3016 4013 3024
rect 3856 2996 3873 3004
rect 4036 3004 4044 3036
rect 4007 2996 4044 3004
rect 3776 2976 3913 2984
rect 3956 2984 3964 2993
rect 3956 2976 3993 2984
rect 4056 2984 4064 3076
rect 4507 3076 4604 3084
rect 4187 3056 4213 3064
rect 4387 3056 4493 3064
rect 4247 3036 4284 3044
rect 4276 3024 4284 3036
rect 4276 3016 4373 3024
rect 4407 3016 4453 3024
rect 4507 3016 4553 3024
rect 4216 3004 4224 3013
rect 4167 2996 4224 3004
rect 4256 3004 4264 3013
rect 4256 2996 4304 3004
rect 4047 2976 4064 2984
rect 4236 2984 4244 2993
rect 4227 2976 4244 2984
rect 1747 2956 1913 2964
rect 2427 2956 2853 2964
rect 3027 2956 3153 2964
rect 3167 2956 3353 2964
rect 3367 2956 3613 2964
rect 3727 2956 3813 2964
rect 3987 2956 4053 2964
rect 4296 2964 4304 2996
rect 4347 2996 4393 3004
rect 4487 2996 4513 3004
rect 4576 3004 4584 3053
rect 4596 3027 4604 3076
rect 4687 3076 4773 3084
rect 4707 3056 4733 3064
rect 4656 3044 4664 3053
rect 4656 3036 4804 3044
rect 4607 3016 4624 3024
rect 4616 3007 4624 3016
rect 4647 3016 4693 3024
rect 4547 2996 4584 3004
rect 4796 3004 4804 3036
rect 4796 2996 4824 3004
rect 4327 2976 4433 2984
rect 4507 2976 4553 2984
rect 4187 2956 4304 2964
rect 4367 2956 4513 2964
rect 1227 2936 2333 2944
rect 2447 2936 3253 2944
rect 3267 2936 3493 2944
rect 3527 2936 3793 2944
rect 3947 2936 4093 2944
rect 1527 2916 1673 2924
rect 1687 2916 2213 2924
rect 2647 2916 3193 2924
rect 3227 2916 4413 2924
rect 1667 2896 1753 2904
rect 1767 2896 1793 2904
rect 2407 2896 3273 2904
rect 3287 2896 3553 2904
rect 3767 2896 4173 2904
rect 47 2876 233 2884
rect 2927 2876 3313 2884
rect 3447 2876 3953 2884
rect 4167 2876 4233 2884
rect 387 2856 433 2864
rect 2227 2856 2273 2864
rect 2307 2856 2453 2864
rect 2807 2856 2933 2864
rect 2947 2856 3113 2864
rect 3387 2856 3513 2864
rect 2187 2836 2293 2844
rect 2547 2836 2913 2844
rect 2967 2836 3133 2844
rect 3207 2836 3433 2844
rect 3467 2836 3733 2844
rect 3787 2836 4613 2844
rect 607 2816 633 2824
rect 967 2816 1013 2824
rect 1387 2816 1573 2824
rect 2087 2816 2173 2824
rect 2567 2816 2713 2824
rect 2827 2816 3293 2824
rect 3307 2816 3313 2824
rect 3407 2816 3513 2824
rect 3567 2816 3833 2824
rect 3856 2816 3904 2824
rect 227 2796 333 2804
rect 647 2796 704 2804
rect 167 2776 293 2784
rect 347 2776 373 2784
rect 427 2776 553 2784
rect 316 2764 324 2773
rect 296 2756 324 2764
rect 296 2727 304 2756
rect 407 2756 473 2764
rect 527 2756 653 2764
rect 676 2747 684 2773
rect 407 2736 433 2744
rect 696 2744 704 2796
rect 1567 2796 1993 2804
rect 2627 2796 2753 2804
rect 2787 2796 2924 2804
rect 736 2776 993 2784
rect 736 2767 744 2776
rect 1007 2776 1053 2784
rect 1107 2776 1133 2784
rect 1187 2776 1513 2784
rect 1827 2776 1873 2784
rect 1887 2776 1953 2784
rect 2096 2776 2213 2784
rect 2096 2767 2104 2776
rect 2587 2776 2773 2784
rect 2787 2776 2833 2784
rect 1587 2756 1744 2764
rect 696 2736 753 2744
rect 776 2744 784 2753
rect 1736 2747 1744 2756
rect 1876 2756 1913 2764
rect 776 2736 873 2744
rect 1267 2736 1293 2744
rect 1487 2736 1613 2744
rect 1647 2736 1713 2744
rect 1756 2736 1853 2744
rect 367 2716 573 2724
rect 587 2716 693 2724
rect 867 2716 893 2724
rect 987 2716 1013 2724
rect 1507 2716 1633 2724
rect 1756 2724 1764 2736
rect 1687 2716 1764 2724
rect 1876 2724 1884 2756
rect 2556 2764 2564 2773
rect 2127 2756 2464 2764
rect 2556 2756 2593 2764
rect 1847 2716 1884 2724
rect 1936 2724 1944 2753
rect 2047 2736 2153 2744
rect 2216 2736 2433 2744
rect 2216 2727 2224 2736
rect 2456 2744 2464 2756
rect 2747 2756 2793 2764
rect 2856 2764 2864 2773
rect 2847 2756 2864 2764
rect 2456 2736 2613 2744
rect 2696 2744 2704 2753
rect 2696 2736 2753 2744
rect 1927 2716 1944 2724
rect 2267 2716 2873 2724
rect 2896 2724 2904 2773
rect 2916 2764 2924 2796
rect 3207 2796 3233 2804
rect 3856 2804 3864 2816
rect 3507 2796 3864 2804
rect 3096 2767 3104 2793
rect 2916 2756 2964 2764
rect 2956 2744 2964 2756
rect 3136 2764 3144 2793
rect 3156 2784 3164 2793
rect 3156 2776 3173 2784
rect 3547 2776 3644 2784
rect 3136 2756 3153 2764
rect 3167 2756 3233 2764
rect 3336 2764 3344 2773
rect 3256 2756 3344 2764
rect 2956 2736 2973 2744
rect 2896 2716 2913 2724
rect 107 2696 493 2704
rect 887 2696 1133 2704
rect 1787 2696 1933 2704
rect 2207 2696 2553 2704
rect 2567 2696 2573 2704
rect 2667 2696 2713 2704
rect 2936 2704 2944 2733
rect 3056 2724 3064 2753
rect 3107 2736 3153 2744
rect 3256 2744 3264 2756
rect 3367 2756 3433 2764
rect 3496 2756 3613 2764
rect 3187 2736 3264 2744
rect 3447 2736 3473 2744
rect 3056 2716 3133 2724
rect 3496 2724 3504 2756
rect 3147 2716 3504 2724
rect 3636 2724 3644 2776
rect 3667 2756 3693 2764
rect 3756 2764 3764 2773
rect 3756 2756 3793 2764
rect 3816 2744 3824 2773
rect 3876 2764 3884 2793
rect 3896 2787 3904 2816
rect 3967 2816 4273 2824
rect 4287 2816 4713 2824
rect 4096 2796 4184 2804
rect 3876 2756 3893 2764
rect 3727 2736 3853 2744
rect 3916 2744 3924 2793
rect 4096 2784 4104 2796
rect 4176 2787 4184 2796
rect 4687 2796 4733 2804
rect 3967 2776 4104 2784
rect 4047 2756 4073 2764
rect 4096 2764 4104 2776
rect 4127 2776 4144 2784
rect 4096 2756 4113 2764
rect 3916 2736 3933 2744
rect 3976 2744 3984 2753
rect 4136 2747 4144 2776
rect 4207 2756 4313 2764
rect 3976 2736 4093 2744
rect 4376 2744 4384 2793
rect 4587 2776 4613 2784
rect 4707 2776 4784 2784
rect 4447 2756 4473 2764
rect 4327 2736 4413 2744
rect 4427 2736 4453 2744
rect 4496 2744 4504 2773
rect 4527 2756 4593 2764
rect 4647 2756 4753 2764
rect 4496 2736 4533 2744
rect 4776 2744 4784 2776
rect 4707 2736 4784 2744
rect 3627 2716 3644 2724
rect 3847 2716 3893 2724
rect 4007 2716 4053 2724
rect 4067 2716 4153 2724
rect 4167 2716 4173 2724
rect 4187 2716 4353 2724
rect 4407 2716 4573 2724
rect 4647 2716 4713 2724
rect 2887 2696 2944 2704
rect 3007 2696 3053 2704
rect 3087 2696 3173 2704
rect 3267 2696 3693 2704
rect 3887 2696 3973 2704
rect 4087 2696 4433 2704
rect 4607 2696 4773 2704
rect 587 2676 973 2684
rect 987 2676 1233 2684
rect 1707 2676 1813 2684
rect 2327 2676 2513 2684
rect 2567 2676 2653 2684
rect 2667 2676 2673 2684
rect 2727 2676 3033 2684
rect 3287 2676 3393 2684
rect 3507 2676 3633 2684
rect 3827 2676 3913 2684
rect 3947 2676 4233 2684
rect 4307 2676 4513 2684
rect 4547 2676 4653 2684
rect 4747 2676 4773 2684
rect 687 2656 713 2664
rect 727 2656 933 2664
rect 1807 2656 1993 2664
rect 2047 2656 2233 2664
rect 2527 2656 2833 2664
rect 2907 2656 3293 2664
rect 3416 2656 3533 2664
rect 507 2636 593 2644
rect 747 2636 873 2644
rect 1187 2636 1213 2644
rect 1227 2636 1313 2644
rect 1447 2636 1473 2644
rect 2667 2636 2893 2644
rect 3416 2644 3424 2656
rect 3727 2656 4033 2664
rect 4047 2656 4373 2664
rect 4567 2656 4653 2664
rect 3347 2636 3424 2644
rect 3487 2636 3873 2644
rect 4067 2636 4193 2644
rect 4447 2636 4713 2644
rect 107 2616 373 2624
rect 427 2616 453 2624
rect 527 2616 533 2624
rect 547 2616 593 2624
rect 687 2616 1073 2624
rect 1167 2616 1273 2624
rect 1287 2616 1353 2624
rect 1407 2616 1493 2624
rect 1507 2616 1513 2624
rect 1527 2616 1853 2624
rect 1867 2616 2013 2624
rect 2467 2616 2853 2624
rect 3067 2616 3353 2624
rect 3627 2616 3673 2624
rect 3747 2616 4013 2624
rect 4167 2616 4253 2624
rect 4267 2616 4393 2624
rect 4427 2616 4693 2624
rect 247 2596 613 2604
rect 627 2596 2133 2604
rect 2287 2596 2613 2604
rect 2827 2596 2933 2604
rect 3307 2596 3573 2604
rect 3607 2596 3793 2604
rect 287 2576 313 2584
rect 367 2576 613 2584
rect 867 2576 1653 2584
rect -24 2544 -16 2564
rect 127 2556 333 2564
rect 387 2556 553 2564
rect 607 2556 653 2564
rect 807 2556 1084 2564
rect -24 2536 104 2544
rect 96 2527 104 2536
rect 247 2536 313 2544
rect 467 2536 533 2544
rect 587 2536 673 2544
rect 767 2536 853 2544
rect 1076 2544 1084 2556
rect 1167 2556 1213 2564
rect 1296 2547 1304 2576
rect 1727 2576 2173 2584
rect 2587 2576 2673 2584
rect 2896 2576 3013 2584
rect 1367 2556 1433 2564
rect 1567 2556 1693 2564
rect 1787 2556 1813 2564
rect 1867 2556 2313 2564
rect 2327 2556 2353 2564
rect 2367 2556 2433 2564
rect 1076 2536 1133 2544
rect 1147 2536 1193 2544
rect 1316 2536 1353 2544
rect -24 2516 73 2524
rect 227 2516 373 2524
rect 387 2516 433 2524
rect 487 2516 513 2524
rect 527 2516 593 2524
rect 647 2516 753 2524
rect 947 2516 1153 2524
rect 1236 2524 1244 2533
rect 1316 2524 1324 2536
rect 2316 2544 2324 2553
rect 2516 2547 2524 2573
rect 2896 2564 2904 2576
rect 3207 2576 3273 2584
rect 3527 2576 3613 2584
rect 3687 2576 3713 2584
rect 3736 2576 3753 2584
rect 2756 2556 2904 2564
rect 2167 2536 2324 2544
rect 2567 2536 2593 2544
rect 2647 2536 2693 2544
rect 2756 2544 2764 2556
rect 2987 2556 3073 2564
rect 3096 2556 3133 2564
rect 2707 2536 2764 2544
rect 2787 2536 2833 2544
rect 2916 2544 2924 2553
rect 3096 2547 3104 2556
rect 3207 2556 3293 2564
rect 3307 2556 3313 2564
rect 3416 2547 3424 2573
rect 3547 2556 3613 2564
rect 2856 2536 2924 2544
rect 1236 2516 1324 2524
rect 1347 2516 1673 2524
rect 1687 2516 2113 2524
rect 2227 2516 2753 2524
rect 2856 2524 2864 2536
rect 3047 2536 3093 2544
rect 3636 2544 3644 2553
rect 3636 2536 3713 2544
rect 2767 2516 2864 2524
rect 2887 2516 2973 2524
rect 3147 2516 3233 2524
rect 3327 2516 3433 2524
rect 3547 2516 3613 2524
rect 3736 2524 3744 2576
rect 3807 2576 4073 2584
rect 4127 2576 4153 2584
rect 4376 2576 4533 2584
rect 3767 2556 3933 2564
rect 3956 2556 4033 2564
rect 3956 2544 3964 2556
rect 3927 2536 3964 2544
rect 4056 2544 4064 2553
rect 4047 2536 4064 2544
rect 4136 2527 4144 2553
rect 3736 2516 3793 2524
rect 3887 2516 4053 2524
rect 4176 2507 4184 2573
rect 4376 2564 4384 2576
rect 4356 2556 4384 2564
rect 4196 2527 4204 2553
rect 4227 2536 4273 2544
rect 4287 2536 4333 2544
rect 4356 2527 4364 2556
rect 4407 2556 4493 2564
rect 4556 2564 4564 2573
rect 4527 2556 4564 2564
rect 4667 2556 4704 2564
rect 4696 2544 4704 2556
rect 4696 2536 4724 2544
rect 4267 2516 4313 2524
rect 4347 2516 4353 2524
rect 4376 2507 4384 2533
rect 4407 2516 4424 2524
rect 4416 2507 4424 2516
rect 27 2496 333 2504
rect 707 2496 773 2504
rect 3007 2496 3033 2504
rect 3047 2496 3573 2504
rect 3587 2496 3593 2504
rect 3827 2496 3913 2504
rect 3927 2496 3953 2504
rect 3967 2496 3993 2504
rect 3127 2476 3173 2484
rect 3527 2476 3733 2484
rect 4087 2476 4293 2484
rect 4476 2484 4484 2533
rect 4516 2524 4524 2533
rect 4516 2516 4573 2524
rect 4587 2516 4653 2524
rect 4496 2504 4504 2513
rect 4676 2507 4684 2533
rect 4496 2496 4553 2504
rect 4696 2487 4704 2513
rect 4716 2507 4724 2536
rect 4476 2476 4493 2484
rect 4507 2476 4533 2484
rect 87 2456 2453 2464
rect 2787 2456 3213 2464
rect 3767 2456 4153 2464
rect 4267 2456 4633 2464
rect 4667 2456 4773 2464
rect 107 2436 1153 2444
rect 2967 2436 3113 2444
rect 3127 2436 3233 2444
rect 3267 2436 3873 2444
rect 4007 2436 4453 2444
rect 4467 2436 4713 2444
rect 1387 2416 1453 2424
rect 2467 2416 2613 2424
rect 2767 2416 3533 2424
rect 4167 2416 4233 2424
rect 4367 2416 4553 2424
rect 2407 2396 2573 2404
rect 2587 2396 3173 2404
rect 3187 2396 3453 2404
rect 3627 2396 4133 2404
rect 4207 2396 4513 2404
rect 4527 2396 4713 2404
rect 4727 2396 4733 2404
rect 1447 2376 1473 2384
rect 2227 2376 2533 2384
rect 2547 2376 2713 2384
rect 3207 2376 4153 2384
rect 4207 2376 4373 2384
rect 4387 2376 4673 2384
rect 507 2356 533 2364
rect 727 2356 973 2364
rect 987 2356 1073 2364
rect 1427 2356 1533 2364
rect 2527 2356 3353 2364
rect 3367 2356 3393 2364
rect 3827 2356 4073 2364
rect 4387 2356 4613 2364
rect 427 2336 493 2344
rect 627 2336 2353 2344
rect 2507 2336 2593 2344
rect 2607 2336 2673 2344
rect 2687 2336 2793 2344
rect 2807 2336 3073 2344
rect 3087 2336 3313 2344
rect 3667 2336 3673 2344
rect 3687 2336 4093 2344
rect 4147 2336 4253 2344
rect 4347 2336 4553 2344
rect 267 2316 453 2324
rect 467 2316 1893 2324
rect 2187 2316 2653 2324
rect 2667 2316 2733 2324
rect 2747 2316 2833 2324
rect 2847 2316 2933 2324
rect 3307 2316 3653 2324
rect 3807 2316 4184 2324
rect 227 2296 413 2304
rect 427 2296 553 2304
rect 827 2296 933 2304
rect 1047 2296 1593 2304
rect 1607 2296 2013 2304
rect 2167 2296 2313 2304
rect 2367 2296 2553 2304
rect 2567 2296 2693 2304
rect 2827 2296 2993 2304
rect 3107 2296 3133 2304
rect 3187 2296 3253 2304
rect 3447 2296 3453 2304
rect 3467 2296 3493 2304
rect 3636 2296 3693 2304
rect -24 2276 13 2284
rect 47 2276 273 2284
rect 356 2276 713 2284
rect 356 2267 364 2276
rect 996 2276 1053 2284
rect 107 2256 293 2264
rect 856 2247 864 2273
rect 996 2267 1004 2276
rect 1067 2276 1304 2284
rect 1027 2256 1193 2264
rect 1296 2264 1304 2276
rect 1467 2276 1564 2284
rect 1296 2256 1333 2264
rect 1507 2256 1533 2264
rect 1556 2264 1564 2276
rect 1756 2276 1793 2284
rect 1556 2256 1693 2264
rect 27 2236 613 2244
rect 927 2236 933 2244
rect 947 2236 973 2244
rect 1247 2236 1373 2244
rect 1756 2244 1764 2276
rect 2547 2276 2573 2284
rect 2727 2276 2793 2284
rect 2856 2276 3193 2284
rect 1836 2247 1844 2273
rect 1856 2247 1864 2273
rect 2856 2267 2864 2276
rect 3287 2276 3333 2284
rect 3387 2276 3413 2284
rect 1887 2256 1933 2264
rect 1947 2256 1993 2264
rect 2247 2256 2373 2264
rect 2927 2256 3053 2264
rect 3087 2256 3213 2264
rect 1727 2236 1764 2244
rect 1907 2236 1953 2244
rect 1967 2236 2173 2244
rect 2647 2236 2873 2244
rect 2907 2236 3093 2244
rect 3236 2244 3244 2273
rect 3636 2267 3644 2296
rect 3787 2296 3804 2304
rect 3656 2276 3693 2284
rect 3207 2236 3273 2244
rect 3456 2236 3553 2244
rect 327 2216 573 2224
rect 847 2216 893 2224
rect 1167 2216 2493 2224
rect 2947 2216 3113 2224
rect 3456 2224 3464 2236
rect 3567 2236 3573 2244
rect 3656 2244 3664 2276
rect 3607 2236 3664 2244
rect 3716 2244 3724 2273
rect 3796 2267 3804 2296
rect 3887 2296 4013 2304
rect 3967 2276 4133 2284
rect 3916 2264 3924 2273
rect 4156 2267 4164 2293
rect 3867 2256 3924 2264
rect 4047 2256 4093 2264
rect 4176 2264 4184 2316
rect 4396 2316 4413 2324
rect 4396 2287 4404 2316
rect 4447 2316 4564 2324
rect 4416 2296 4493 2304
rect 4247 2276 4273 2284
rect 4176 2256 4193 2264
rect 4316 2264 4324 2273
rect 4416 2267 4424 2296
rect 4527 2296 4544 2304
rect 4536 2287 4544 2296
rect 4447 2276 4493 2284
rect 4267 2256 4324 2264
rect 4347 2256 4404 2264
rect 3716 2236 3833 2244
rect 3867 2236 3973 2244
rect 3987 2236 4053 2244
rect 4107 2236 4173 2244
rect 4327 2236 4353 2244
rect 4396 2244 4404 2256
rect 4436 2244 4444 2273
rect 4556 2264 4564 2316
rect 4647 2316 4773 2324
rect 4656 2267 4664 2293
rect 4736 2276 4773 2284
rect 4547 2256 4564 2264
rect 4696 2247 4704 2273
rect 4736 2267 4744 2276
rect 4816 2264 4824 2284
rect 4756 2256 4824 2264
rect 4396 2236 4444 2244
rect 4507 2236 4653 2244
rect 4756 2244 4764 2256
rect 4747 2236 4764 2244
rect 4787 2236 4824 2244
rect 3147 2216 3464 2224
rect 3847 2216 4093 2224
rect 4127 2216 4193 2224
rect 4447 2216 4533 2224
rect 347 2196 513 2204
rect 747 2196 1033 2204
rect 1047 2196 1093 2204
rect 1587 2196 1773 2204
rect 2127 2196 2253 2204
rect 2327 2196 2893 2204
rect 2967 2196 2973 2204
rect 2987 2196 3333 2204
rect 3387 2196 3453 2204
rect 3487 2196 3633 2204
rect 3827 2196 3893 2204
rect 3967 2196 4233 2204
rect 4527 2196 4673 2204
rect 4687 2196 4753 2204
rect 647 2176 953 2184
rect 967 2176 1153 2184
rect 1767 2176 1933 2184
rect 2667 2176 2753 2184
rect 2767 2176 2913 2184
rect 2927 2176 3733 2184
rect 3787 2176 4213 2184
rect 4227 2176 4293 2184
rect 4567 2176 4593 2184
rect 4627 2176 4693 2184
rect 167 2156 633 2164
rect 727 2156 873 2164
rect 1027 2156 1773 2164
rect 1827 2156 1893 2164
rect 1907 2156 1913 2164
rect 1927 2156 3593 2164
rect 3727 2156 4773 2164
rect 327 2136 393 2144
rect 647 2136 1193 2144
rect 1727 2136 1833 2144
rect 1847 2136 1913 2144
rect 1927 2136 1973 2144
rect 1987 2136 2193 2144
rect 3347 2136 3893 2144
rect 4196 2136 4253 2144
rect 307 2116 473 2124
rect 607 2116 1133 2124
rect 1647 2116 1653 2124
rect 1667 2116 1733 2124
rect 1767 2116 2133 2124
rect 2147 2116 2153 2124
rect 2487 2116 2613 2124
rect 3027 2116 3293 2124
rect 3427 2116 3533 2124
rect 4196 2124 4204 2136
rect 4387 2136 4733 2144
rect 3587 2116 4204 2124
rect 4227 2116 4493 2124
rect 4527 2116 4573 2124
rect 4587 2116 4633 2124
rect -24 2096 53 2104
rect 267 2096 364 2104
rect 127 2076 333 2084
rect 356 2084 364 2096
rect 867 2096 873 2104
rect 887 2096 913 2104
rect 1007 2096 1033 2104
rect 1087 2096 1273 2104
rect 1307 2096 1413 2104
rect 1487 2096 1873 2104
rect 2067 2096 2313 2104
rect 2407 2096 2573 2104
rect 2687 2096 2753 2104
rect 3116 2096 3173 2104
rect 356 2076 373 2084
rect 396 2076 433 2084
rect -24 2056 13 2064
rect 27 2056 33 2064
rect 267 2056 313 2064
rect 376 2064 384 2073
rect 356 2056 384 2064
rect 167 2036 213 2044
rect 247 2036 333 2044
rect 356 2044 364 2056
rect 347 2036 364 2044
rect 396 2044 404 2076
rect 687 2076 713 2084
rect 747 2076 793 2084
rect 1116 2076 1153 2084
rect 467 2056 493 2064
rect 776 2056 853 2064
rect 776 2047 784 2056
rect 927 2056 953 2064
rect 1016 2047 1024 2073
rect 1116 2067 1124 2076
rect 1327 2076 1373 2084
rect 1507 2076 1613 2084
rect 1787 2076 1793 2084
rect 1807 2076 1853 2084
rect 2467 2076 2593 2084
rect 2727 2076 2853 2084
rect 2987 2076 3013 2084
rect 3116 2084 3124 2096
rect 3207 2096 3393 2104
rect 3407 2096 3473 2104
rect 3507 2096 3593 2104
rect 4107 2096 4453 2104
rect 4576 2096 4713 2104
rect 3056 2076 3124 2084
rect 1167 2056 1213 2064
rect 1427 2056 1633 2064
rect 1947 2056 2033 2064
rect 2267 2056 2333 2064
rect 2356 2064 2364 2073
rect 2356 2056 2464 2064
rect 387 2036 404 2044
rect 847 2036 933 2044
rect 1087 2036 1173 2044
rect 1247 2036 1373 2044
rect 1987 2036 2133 2044
rect 2187 2036 2273 2044
rect 2287 2036 2373 2044
rect 2387 2036 2433 2044
rect 207 2016 233 2024
rect 367 2016 733 2024
rect 887 2016 973 2024
rect 1067 2016 1253 2024
rect 2107 2016 2233 2024
rect 2456 2024 2464 2056
rect 2547 2056 2693 2064
rect 2487 2036 2493 2044
rect 2507 2036 2513 2044
rect 3056 2044 3064 2076
rect 3167 2076 3244 2084
rect 3236 2064 3244 2076
rect 3267 2076 3413 2084
rect 3447 2076 3513 2084
rect 3536 2076 3553 2084
rect 3236 2056 3304 2064
rect 3296 2047 3304 2056
rect 3347 2056 3373 2064
rect 3027 2036 3064 2044
rect 3127 2036 3173 2044
rect 3416 2044 3424 2053
rect 3367 2036 3433 2044
rect 2456 2016 2753 2024
rect 3107 2016 3213 2024
rect 3227 2016 3313 2024
rect 3536 2024 3544 2076
rect 3616 2084 3624 2093
rect 3596 2076 3624 2084
rect 3596 2067 3604 2076
rect 3807 2076 3864 2084
rect 3647 2056 3673 2064
rect 3707 2056 3733 2064
rect 3856 2064 3864 2076
rect 3887 2076 3924 2084
rect 3787 2056 3844 2064
rect 3856 2056 3884 2064
rect 3836 2047 3844 2056
rect 3876 2047 3884 2056
rect 3916 2047 3924 2076
rect 3936 2067 3944 2093
rect 4147 2076 4233 2084
rect 4247 2076 4304 2084
rect 4296 2064 4304 2076
rect 4327 2076 4364 2084
rect 4356 2067 4364 2076
rect 4376 2076 4413 2084
rect 4376 2067 4384 2076
rect 4516 2076 4553 2084
rect 4516 2067 4524 2076
rect 4067 2056 4284 2064
rect 4296 2056 4333 2064
rect 3627 2036 3673 2044
rect 3727 2036 3793 2044
rect 4276 2044 4284 2056
rect 4276 2036 4484 2044
rect 3467 2016 3544 2024
rect 3647 2016 3653 2024
rect 3667 2016 4113 2024
rect 4207 2016 4273 2024
rect 4476 2024 4484 2036
rect 4556 2044 4564 2053
rect 4507 2036 4564 2044
rect 4576 2044 4584 2096
rect 4607 2076 4684 2084
rect 4607 2056 4644 2064
rect 4576 2036 4613 2044
rect 4476 2016 4533 2024
rect 4636 2024 4644 2056
rect 4676 2047 4684 2076
rect 4696 2027 4704 2073
rect 4787 2036 4824 2044
rect 4547 2016 4644 2024
rect 227 1996 273 2004
rect 287 1996 413 2004
rect 827 1996 913 2004
rect 2227 1996 2553 2004
rect 2567 1996 2673 2004
rect 2747 1996 3393 2004
rect 3407 1996 3513 2004
rect 3807 1996 4233 2004
rect 4247 1996 4293 2004
rect 4447 1996 4573 2004
rect 4587 1996 4713 2004
rect 67 1976 2093 1984
rect 2447 1976 2633 1984
rect 3127 1976 3153 1984
rect 3387 1976 3733 1984
rect 3747 1976 3753 1984
rect 147 1956 733 1964
rect 827 1956 993 1964
rect 2687 1956 2933 1964
rect 2947 1956 3073 1964
rect 3087 1956 3173 1964
rect 3307 1956 3633 1964
rect 3947 1956 4313 1964
rect 1747 1936 2173 1944
rect 2187 1936 4713 1944
rect 2327 1916 4773 1924
rect 3007 1896 3193 1904
rect 3847 1896 3953 1904
rect 4407 1896 4773 1904
rect 2427 1876 2493 1884
rect 2507 1876 3013 1884
rect 3256 1876 3613 1884
rect 1987 1856 2033 1864
rect 2896 1856 3053 1864
rect 327 1836 344 1844
rect 336 1824 344 1836
rect 367 1836 553 1844
rect 567 1836 693 1844
rect 707 1836 813 1844
rect 1267 1836 2073 1844
rect 2896 1844 2904 1856
rect 3256 1864 3264 1876
rect 3707 1876 3853 1884
rect 3867 1876 4213 1884
rect 4567 1876 4633 1884
rect 3067 1856 3264 1864
rect 3287 1856 3693 1864
rect 3727 1856 4153 1864
rect 4347 1856 4373 1864
rect 4527 1856 4653 1864
rect 2867 1836 2904 1844
rect 3067 1836 3233 1844
rect 3367 1836 3373 1844
rect 3387 1836 3473 1844
rect 3867 1836 4053 1844
rect 4067 1836 4153 1844
rect 4167 1836 4253 1844
rect 4267 1836 4333 1844
rect 4547 1836 4604 1844
rect 336 1816 484 1824
rect 147 1776 173 1784
rect 147 1756 233 1764
rect 276 1764 284 1793
rect 296 1787 304 1813
rect 476 1807 484 1816
rect 496 1816 533 1824
rect 427 1796 453 1804
rect 496 1787 504 1816
rect 627 1816 773 1824
rect 927 1816 1084 1824
rect 827 1796 893 1804
rect 1076 1804 1084 1816
rect 1107 1816 1153 1824
rect 1167 1816 1193 1824
rect 1427 1816 1893 1824
rect 2027 1816 2433 1824
rect 2547 1816 2833 1824
rect 3047 1816 3113 1824
rect 3196 1816 3253 1824
rect 1236 1804 1244 1813
rect 1076 1796 1273 1804
rect 1287 1796 1333 1804
rect 1547 1796 1573 1804
rect 1587 1796 1593 1804
rect 2047 1796 2093 1804
rect 2176 1796 2213 1804
rect 516 1784 524 1793
rect 516 1776 593 1784
rect 676 1784 684 1793
rect 647 1776 684 1784
rect 736 1784 744 1793
rect 736 1776 793 1784
rect 847 1776 873 1784
rect 1227 1776 1293 1784
rect 1667 1776 1833 1784
rect 1856 1784 1864 1793
rect 2176 1784 2184 1796
rect 2307 1796 2393 1804
rect 3156 1804 3164 1813
rect 3107 1796 3164 1804
rect 1856 1776 1944 1784
rect 1936 1767 1944 1776
rect 2136 1776 2184 1784
rect 2136 1767 2144 1776
rect 2247 1776 2413 1784
rect 2527 1776 2593 1784
rect 2647 1776 2873 1784
rect 2967 1776 3073 1784
rect 3196 1784 3204 1816
rect 3547 1816 3593 1824
rect 3887 1816 3904 1824
rect 3416 1804 3424 1813
rect 3227 1796 3573 1804
rect 3896 1804 3904 1816
rect 3927 1816 4013 1824
rect 4056 1816 4073 1824
rect 4036 1804 4044 1813
rect 3896 1796 3924 1804
rect 3916 1787 3924 1796
rect 4016 1796 4044 1804
rect 3167 1776 3204 1784
rect 3216 1776 3293 1784
rect 276 1756 393 1764
rect 447 1756 633 1764
rect 647 1756 833 1764
rect 1047 1756 1313 1764
rect 1367 1756 1733 1764
rect 1807 1756 1913 1764
rect 2167 1756 2273 1764
rect 2387 1756 2633 1764
rect 3216 1764 3224 1776
rect 3407 1776 3433 1784
rect 3467 1776 3533 1784
rect 3547 1776 3633 1784
rect 3687 1776 3893 1784
rect 3947 1776 3973 1784
rect 4016 1767 4024 1796
rect 3107 1756 3224 1764
rect 3247 1756 3553 1764
rect 3567 1756 3713 1764
rect 3887 1756 3993 1764
rect 4056 1764 4064 1816
rect 4096 1816 4213 1824
rect 4096 1787 4104 1816
rect 4236 1816 4353 1824
rect 4236 1804 4244 1816
rect 4467 1816 4513 1824
rect 4176 1796 4244 1804
rect 4087 1776 4093 1784
rect 4056 1756 4073 1764
rect 4176 1764 4184 1796
rect 4287 1796 4413 1804
rect 4467 1796 4493 1804
rect 4507 1796 4533 1804
rect 4207 1776 4393 1784
rect 4556 1784 4564 1793
rect 4487 1776 4564 1784
rect 4576 1784 4584 1813
rect 4596 1804 4604 1836
rect 4647 1836 4693 1844
rect 4627 1816 4704 1824
rect 4596 1796 4633 1804
rect 4576 1776 4604 1784
rect 4176 1756 4213 1764
rect 4287 1756 4353 1764
rect 4387 1756 4553 1764
rect 4567 1756 4573 1764
rect 4596 1764 4604 1776
rect 4627 1776 4653 1784
rect 4596 1756 4613 1764
rect 4676 1764 4684 1793
rect 4696 1767 4704 1816
rect 4636 1756 4684 1764
rect 2107 1736 2213 1744
rect 2407 1736 3213 1744
rect 3647 1736 3733 1744
rect 3767 1736 3793 1744
rect 4067 1736 4313 1744
rect 4636 1744 4644 1756
rect 4487 1736 4644 1744
rect 827 1716 1813 1724
rect 1827 1716 1873 1724
rect 1887 1716 1893 1724
rect 1907 1716 1953 1724
rect 1967 1716 2053 1724
rect 2067 1716 2113 1724
rect 2127 1716 2193 1724
rect 2587 1716 2813 1724
rect 2827 1716 3153 1724
rect 3407 1716 3653 1724
rect 3767 1716 3913 1724
rect 4047 1716 4673 1724
rect 4687 1716 4693 1724
rect 1647 1696 1693 1704
rect 2747 1696 2893 1704
rect 2907 1696 3993 1704
rect 4007 1696 4133 1704
rect 4147 1696 4173 1704
rect 4187 1696 4293 1704
rect 1947 1676 1973 1684
rect 2607 1676 3073 1684
rect 3087 1676 3233 1684
rect 3507 1676 3593 1684
rect 3607 1676 3633 1684
rect 3667 1676 4333 1684
rect 367 1656 753 1664
rect 767 1656 933 1664
rect 1927 1656 2033 1664
rect 3227 1656 3253 1664
rect 3327 1656 3493 1664
rect 3527 1656 3693 1664
rect 3707 1656 3773 1664
rect 3907 1656 3973 1664
rect 4027 1656 4093 1664
rect 4167 1656 4193 1664
rect 4207 1656 4353 1664
rect 187 1636 733 1644
rect 747 1636 953 1644
rect 967 1636 1073 1644
rect 1887 1636 1913 1644
rect 2807 1636 2873 1644
rect 2967 1636 3093 1644
rect 3207 1636 3253 1644
rect 3267 1636 3293 1644
rect 3327 1636 3533 1644
rect 3627 1636 3713 1644
rect 3827 1636 3853 1644
rect 3967 1636 4033 1644
rect 4127 1636 4233 1644
rect 4407 1636 4433 1644
rect 4467 1636 4653 1644
rect 327 1616 333 1624
rect 347 1616 533 1624
rect 607 1616 693 1624
rect 707 1616 853 1624
rect 1387 1616 1473 1624
rect 1487 1616 1633 1624
rect 1647 1616 1953 1624
rect 1967 1616 2053 1624
rect 2307 1616 2393 1624
rect 2547 1616 2633 1624
rect 2647 1616 2653 1624
rect 2876 1616 3133 1624
rect 2876 1607 2884 1616
rect 3147 1616 3453 1624
rect 3467 1616 3493 1624
rect 3516 1616 3673 1624
rect 287 1596 293 1604
rect 307 1596 453 1604
rect 467 1596 673 1604
rect 687 1596 873 1604
rect 1227 1596 1413 1604
rect 1607 1596 1773 1604
rect 1796 1596 1853 1604
rect 187 1576 393 1584
rect 407 1576 473 1584
rect 527 1576 573 1584
rect 1147 1576 1193 1584
rect 1247 1576 1273 1584
rect 1796 1584 1804 1596
rect 2147 1596 2233 1604
rect 2247 1596 2253 1604
rect 2316 1596 2333 1604
rect 1727 1576 1804 1584
rect 1847 1576 1933 1584
rect 2316 1567 2324 1596
rect 2387 1596 2573 1604
rect 2896 1596 2933 1604
rect 2896 1584 2904 1596
rect 2947 1596 3133 1604
rect 3156 1596 3173 1604
rect 2707 1576 2904 1584
rect 3007 1576 3033 1584
rect 3156 1584 3164 1596
rect 3236 1596 3273 1604
rect 3056 1576 3164 1584
rect 167 1556 233 1564
rect 1127 1556 1233 1564
rect 1807 1556 1913 1564
rect 2167 1556 2273 1564
rect 2927 1556 2973 1564
rect 3056 1564 3064 1576
rect 3236 1567 3244 1596
rect 3327 1596 3433 1604
rect 3516 1604 3524 1616
rect 3787 1616 3893 1624
rect 3967 1616 4013 1624
rect 4036 1616 4053 1624
rect 3487 1596 3584 1604
rect 3576 1587 3584 1596
rect 3716 1596 3813 1604
rect 3716 1587 3724 1596
rect 3896 1596 3933 1604
rect 3896 1587 3904 1596
rect 4036 1604 4044 1616
rect 4087 1616 4173 1624
rect 4227 1616 4404 1624
rect 3996 1596 4044 1604
rect 3996 1587 4004 1596
rect 4107 1596 4124 1604
rect 3367 1576 3413 1584
rect 3527 1576 3564 1584
rect 2996 1556 3064 1564
rect 2996 1547 3004 1556
rect 3127 1556 3233 1564
rect 3287 1556 3333 1564
rect 3347 1556 3513 1564
rect 3556 1564 3564 1576
rect 3607 1576 3673 1584
rect 3747 1576 3773 1584
rect 3807 1576 3873 1584
rect 3556 1556 3633 1564
rect 3647 1556 3913 1564
rect 4036 1564 4044 1573
rect 4027 1556 4044 1564
rect 4116 1547 4124 1596
rect 4136 1567 4144 1593
rect 4196 1587 4204 1613
rect 4216 1564 4224 1593
rect 4247 1576 4273 1584
rect 4216 1556 4264 1564
rect 1167 1536 1293 1544
rect 2607 1536 2893 1544
rect 3027 1536 3273 1544
rect 3407 1536 3673 1544
rect 3687 1536 4093 1544
rect 4256 1544 4264 1556
rect 4296 1564 4304 1593
rect 4327 1576 4373 1584
rect 4287 1556 4304 1564
rect 4396 1564 4404 1616
rect 4447 1616 4464 1624
rect 4416 1584 4424 1593
rect 4416 1576 4433 1584
rect 4456 1567 4464 1616
rect 4627 1616 4664 1624
rect 4527 1596 4553 1604
rect 4576 1596 4633 1604
rect 4576 1584 4584 1596
rect 4536 1576 4584 1584
rect 4387 1556 4404 1564
rect 4256 1536 4433 1544
rect 4447 1536 4493 1544
rect 4516 1544 4524 1573
rect 4536 1567 4544 1576
rect 4656 1584 4664 1616
rect 4636 1576 4664 1584
rect 4596 1547 4604 1573
rect 4636 1547 4644 1576
rect 4676 1547 4684 1573
rect 4516 1536 4533 1544
rect 47 1516 1593 1524
rect 2607 1516 2833 1524
rect 2847 1516 3013 1524
rect 3067 1516 3093 1524
rect 3567 1516 3713 1524
rect 4027 1516 4153 1524
rect 4227 1516 4393 1524
rect 4407 1516 4693 1524
rect 2827 1496 3153 1504
rect 3167 1496 3453 1504
rect 4507 1496 4653 1504
rect 567 1476 773 1484
rect 907 1476 1153 1484
rect 2787 1476 2853 1484
rect 2907 1476 3273 1484
rect 3287 1476 3373 1484
rect 3947 1476 4773 1484
rect 2687 1456 3013 1464
rect 3027 1456 3073 1464
rect 3087 1456 3253 1464
rect 3767 1456 4193 1464
rect 4287 1456 4353 1464
rect 4367 1456 4573 1464
rect 2367 1436 2393 1444
rect 3307 1436 3553 1444
rect 4087 1436 4113 1444
rect 4127 1436 4173 1444
rect 4647 1436 4773 1444
rect 267 1416 293 1424
rect 827 1416 913 1424
rect 927 1416 1053 1424
rect 3007 1416 3193 1424
rect 3487 1416 3573 1424
rect 4027 1416 4233 1424
rect 1207 1396 1433 1404
rect 2507 1396 3593 1404
rect 3807 1396 3993 1404
rect 4007 1396 4333 1404
rect 4647 1396 4673 1404
rect 1107 1376 1133 1384
rect 1247 1376 1353 1384
rect 1367 1376 1413 1384
rect 1427 1376 1533 1384
rect 1667 1376 2293 1384
rect 2307 1376 2313 1384
rect 3047 1376 3133 1384
rect 3327 1376 3353 1384
rect 3367 1376 3533 1384
rect 4087 1376 4133 1384
rect 4147 1376 4153 1384
rect 4327 1376 4413 1384
rect 487 1356 533 1364
rect 787 1356 993 1364
rect 1107 1356 1173 1364
rect 1187 1356 1653 1364
rect 2447 1356 2753 1364
rect 2847 1356 2933 1364
rect 2947 1356 3033 1364
rect 3047 1356 3313 1364
rect 3327 1356 3613 1364
rect 3787 1356 3893 1364
rect 4107 1356 4184 1364
rect 467 1336 493 1344
rect 696 1336 813 1344
rect 696 1327 704 1336
rect 827 1336 853 1344
rect 867 1336 1093 1344
rect 1467 1336 1713 1344
rect 3216 1336 3273 1344
rect 527 1316 593 1324
rect 747 1316 773 1324
rect 967 1316 1053 1324
rect 1267 1316 1313 1324
rect 1447 1316 1493 1324
rect 1687 1316 1753 1324
rect 1807 1316 2053 1324
rect 2107 1316 2153 1324
rect 2207 1316 2273 1324
rect 347 1296 613 1304
rect 127 1276 353 1284
rect 367 1276 373 1284
rect 636 1284 644 1313
rect 2456 1307 2464 1333
rect 847 1296 913 1304
rect 927 1296 1573 1304
rect 1627 1296 1813 1304
rect 1867 1296 1893 1304
rect 1987 1296 2173 1304
rect 2507 1296 2553 1304
rect 2707 1296 2773 1304
rect 2956 1304 2964 1333
rect 2987 1316 3133 1324
rect 3216 1307 3224 1336
rect 3387 1336 3444 1344
rect 3336 1324 3344 1333
rect 3276 1316 3344 1324
rect 3276 1307 3284 1316
rect 3367 1316 3393 1324
rect 3436 1324 3444 1336
rect 3467 1336 3493 1344
rect 3516 1336 3533 1344
rect 3516 1327 3524 1336
rect 3847 1336 3893 1344
rect 4067 1336 4093 1344
rect 3436 1316 3464 1324
rect 3456 1307 3464 1316
rect 3596 1307 3604 1333
rect 3756 1324 3764 1333
rect 3716 1316 3764 1324
rect 3836 1316 3973 1324
rect 3716 1307 3724 1316
rect 2956 1296 3113 1304
rect 3307 1296 3324 1304
rect 636 1276 673 1284
rect 756 1284 764 1293
rect 3316 1287 3324 1296
rect 3647 1296 3693 1304
rect 3836 1304 3844 1316
rect 3747 1296 3844 1304
rect 3996 1304 4004 1333
rect 4027 1316 4144 1324
rect 4136 1307 4144 1316
rect 4176 1307 4184 1356
rect 4227 1356 4353 1364
rect 4487 1356 4704 1364
rect 4256 1336 4313 1344
rect 4256 1307 4264 1336
rect 4376 1344 4384 1353
rect 4336 1336 4384 1344
rect 4516 1336 4533 1344
rect 4336 1324 4344 1336
rect 4516 1327 4524 1336
rect 4607 1336 4653 1344
rect 4287 1316 4344 1324
rect 4436 1316 4473 1324
rect 4436 1307 4444 1316
rect 4547 1316 4593 1324
rect 3867 1296 4004 1304
rect 4047 1296 4113 1304
rect 4307 1296 4353 1304
rect 4616 1304 4624 1313
rect 4596 1296 4624 1304
rect 4596 1287 4604 1296
rect 756 1276 913 1284
rect 947 1276 1153 1284
rect 1167 1276 1413 1284
rect 1827 1276 1973 1284
rect 1987 1276 2133 1284
rect 2527 1276 2873 1284
rect 2887 1276 3013 1284
rect 3087 1276 3153 1284
rect 3387 1276 3593 1284
rect 3827 1276 4373 1284
rect 4387 1276 4453 1284
rect 4467 1276 4533 1284
rect 4636 1284 4644 1336
rect 4696 1307 4704 1356
rect 4627 1276 4644 1284
rect 167 1256 213 1264
rect 567 1256 713 1264
rect 1567 1256 1833 1264
rect 2447 1256 2633 1264
rect 2927 1256 3473 1264
rect 3547 1256 3653 1264
rect 4067 1256 4133 1264
rect 4267 1256 4313 1264
rect 1027 1236 1033 1244
rect 1047 1236 2473 1244
rect 3367 1236 3413 1244
rect 3467 1236 3533 1244
rect 4007 1236 4253 1244
rect 4287 1236 4373 1244
rect 4467 1236 4573 1244
rect 147 1216 193 1224
rect 267 1216 373 1224
rect 387 1216 573 1224
rect 1747 1216 1893 1224
rect 1907 1216 2073 1224
rect 2507 1216 2573 1224
rect 3507 1216 3693 1224
rect 3707 1216 3713 1224
rect 3787 1216 4013 1224
rect 4147 1216 4193 1224
rect 4247 1216 4573 1224
rect 187 1196 293 1204
rect 527 1196 553 1204
rect 567 1196 973 1204
rect 1787 1196 1893 1204
rect 2507 1196 2993 1204
rect 3007 1196 3553 1204
rect 4007 1196 4153 1204
rect 4287 1196 4633 1204
rect 4667 1196 4773 1204
rect 187 1176 233 1184
rect 887 1176 973 1184
rect 1087 1176 1273 1184
rect 1287 1176 2353 1184
rect 2567 1176 2593 1184
rect 2767 1176 2893 1184
rect 3067 1176 3393 1184
rect 3647 1176 3773 1184
rect 3927 1176 4353 1184
rect 4407 1176 4513 1184
rect 407 1156 633 1164
rect 967 1156 1053 1164
rect 1107 1156 1113 1164
rect 1127 1156 1193 1164
rect 1247 1156 1753 1164
rect 2167 1156 2313 1164
rect 2347 1156 2613 1164
rect 2827 1156 2873 1164
rect 3087 1156 3173 1164
rect 3227 1156 3293 1164
rect 3347 1156 3493 1164
rect 4107 1156 4193 1164
rect 4327 1156 4344 1164
rect 447 1136 533 1144
rect 547 1136 893 1144
rect 1027 1136 1213 1144
rect 1227 1136 1244 1144
rect 36 1116 253 1124
rect 36 1107 44 1116
rect 347 1116 504 1124
rect 496 1107 504 1116
rect 627 1116 653 1124
rect 127 1096 173 1104
rect 287 1096 413 1104
rect 427 1096 473 1104
rect 47 1076 93 1084
rect 147 1076 373 1084
rect 467 1076 513 1084
rect 856 1084 864 1113
rect 896 1104 904 1113
rect 896 1096 993 1104
rect 1236 1104 1244 1136
rect 1307 1136 1324 1144
rect 1316 1124 1324 1136
rect 1347 1136 1433 1144
rect 1647 1136 1673 1144
rect 1927 1136 2133 1144
rect 2187 1136 2213 1144
rect 2807 1136 2933 1144
rect 2987 1136 3033 1144
rect 3167 1136 3213 1144
rect 3287 1136 3464 1144
rect 1316 1116 1553 1124
rect 1656 1116 1733 1124
rect 1236 1096 1253 1104
rect 1307 1096 1613 1104
rect 1656 1087 1664 1116
rect 2027 1116 2113 1124
rect 2136 1116 2193 1124
rect 2067 1096 2073 1104
rect 2136 1104 2144 1116
rect 2487 1116 2773 1124
rect 2927 1116 2953 1124
rect 2987 1116 3013 1124
rect 3167 1116 3193 1124
rect 3247 1116 3333 1124
rect 2087 1096 2144 1104
rect 2267 1096 2293 1104
rect 2667 1096 2753 1104
rect 2856 1104 2864 1113
rect 2856 1096 2873 1104
rect 707 1076 913 1084
rect 927 1076 933 1084
rect 1187 1076 1293 1084
rect 1707 1076 1793 1084
rect 2307 1076 2713 1084
rect 2896 1084 2904 1113
rect 2987 1096 3024 1104
rect 3016 1087 3024 1096
rect 3047 1096 3133 1104
rect 3187 1096 3273 1104
rect 3287 1096 3344 1104
rect 3336 1087 3344 1096
rect 3367 1096 3444 1104
rect 2787 1076 2904 1084
rect 327 1056 633 1064
rect 687 1056 713 1064
rect 767 1056 1253 1064
rect 1607 1056 1733 1064
rect 2927 1056 3053 1064
rect 3147 1056 3413 1064
rect 3436 1064 3444 1096
rect 3456 1087 3464 1136
rect 3627 1136 3673 1144
rect 3707 1136 3813 1144
rect 3827 1136 3833 1144
rect 3856 1136 3873 1144
rect 3587 1116 3633 1124
rect 3687 1116 3713 1124
rect 3787 1096 3833 1104
rect 3487 1076 3553 1084
rect 3856 1084 3864 1136
rect 4067 1136 4113 1144
rect 4147 1136 4164 1144
rect 3976 1116 4013 1124
rect 3976 1107 3984 1116
rect 4087 1116 4144 1124
rect 4136 1107 4144 1116
rect 3887 1096 3953 1104
rect 4047 1096 4093 1104
rect 4156 1087 4164 1136
rect 4187 1136 4204 1144
rect 4196 1107 4204 1136
rect 4227 1136 4313 1144
rect 4336 1124 4344 1156
rect 4367 1156 4564 1164
rect 4456 1136 4493 1144
rect 4296 1116 4344 1124
rect 4356 1116 4393 1124
rect 4296 1107 4304 1116
rect 4356 1104 4364 1116
rect 4327 1096 4364 1104
rect 4387 1096 4444 1104
rect 4436 1087 4444 1096
rect 4456 1087 4464 1136
rect 4556 1127 4564 1156
rect 4747 1156 4773 1164
rect 4667 1136 4764 1144
rect 4476 1116 4493 1124
rect 3856 1076 3893 1084
rect 4067 1076 4093 1084
rect 4247 1076 4413 1084
rect 3436 1056 3493 1064
rect 3547 1056 3593 1064
rect 3796 1064 3804 1073
rect 3796 1056 3873 1064
rect 4127 1056 4313 1064
rect 4476 1064 4484 1116
rect 4527 1116 4544 1124
rect 4536 1104 4544 1116
rect 4607 1116 4673 1124
rect 4536 1096 4573 1104
rect 4516 1084 4524 1093
rect 4656 1087 4664 1116
rect 4756 1107 4764 1136
rect 4687 1096 4744 1104
rect 4736 1087 4744 1096
rect 4516 1076 4593 1084
rect 4367 1056 4484 1064
rect 1587 1036 1753 1044
rect 3007 1036 3133 1044
rect 3327 1036 3653 1044
rect 4427 1036 4473 1044
rect 327 1016 373 1024
rect 3107 1016 3373 1024
rect 3647 1016 3933 1024
rect 4167 1016 4273 1024
rect 4667 1016 4753 1024
rect 2847 996 3473 1004
rect 4207 996 4753 1004
rect 3307 976 3553 984
rect 4347 976 4693 984
rect 4127 956 4773 964
rect 2927 936 3513 944
rect 3727 936 4153 944
rect 4467 936 4613 944
rect 1567 916 1933 924
rect 1987 916 2253 924
rect 2267 916 2373 924
rect 2387 916 2653 924
rect 3067 916 3153 924
rect 3167 916 3193 924
rect 3227 916 3613 924
rect 4007 916 4073 924
rect 4227 916 4313 924
rect 4447 916 4493 924
rect 4587 916 4753 924
rect 127 896 353 904
rect 367 896 533 904
rect 547 896 733 904
rect 987 896 1193 904
rect 1207 896 1353 904
rect 1407 896 1453 904
rect 1467 896 2153 904
rect 3207 896 3273 904
rect 3796 896 4013 904
rect 607 876 713 884
rect 1167 876 1493 884
rect 1507 876 1613 884
rect 2047 876 2413 884
rect 2727 876 2773 884
rect 2996 876 3013 884
rect 2996 867 3004 876
rect 3287 876 3353 884
rect 3567 876 3613 884
rect 3627 876 3653 884
rect 3796 867 3804 896
rect 4067 896 4433 904
rect 4547 896 4573 904
rect 4607 896 4613 904
rect 4627 896 4713 904
rect 4747 896 4784 904
rect 3816 876 4093 884
rect 227 856 253 864
rect 307 856 333 864
rect 647 856 673 864
rect 807 856 884 864
rect 876 847 884 856
rect 927 856 1013 864
rect 1027 856 1093 864
rect 1667 856 1993 864
rect 2007 856 2173 864
rect 2187 856 2244 864
rect 287 836 353 844
rect 407 836 453 844
rect 707 836 773 844
rect 107 816 373 824
rect 527 816 793 824
rect 816 824 824 833
rect 816 816 924 824
rect 307 796 333 804
rect 347 796 413 804
rect 427 796 533 804
rect 547 796 593 804
rect 847 796 893 804
rect 916 804 924 816
rect 1087 816 1213 824
rect 916 796 1113 804
rect 1236 804 1244 853
rect 1276 844 1284 853
rect 2236 847 2244 856
rect 2367 856 2493 864
rect 2827 856 2933 864
rect 3047 856 3113 864
rect 3507 856 3524 864
rect 1276 836 1373 844
rect 2207 836 2224 844
rect 1267 816 1433 824
rect 1927 816 2053 824
rect 2096 807 2104 833
rect 2127 816 2153 824
rect 2216 824 2224 836
rect 2347 836 2393 844
rect 2216 816 2233 824
rect 1236 796 1473 804
rect 1487 796 1533 804
rect 1607 796 1633 804
rect 1647 796 2033 804
rect 2296 804 2304 833
rect 2796 827 2804 853
rect 2927 836 2993 844
rect 3027 836 3093 844
rect 3116 836 3213 844
rect 3116 824 3124 836
rect 3047 816 3124 824
rect 3316 824 3324 853
rect 3396 827 3404 853
rect 3187 816 3324 824
rect 3427 816 3493 824
rect 2116 796 2304 804
rect 187 776 353 784
rect 1007 776 1093 784
rect 1107 776 1593 784
rect 2007 776 2073 784
rect 2116 784 2124 796
rect 2847 796 2893 804
rect 2907 796 2944 804
rect 2087 776 2124 784
rect 2147 776 2213 784
rect 2287 776 2313 784
rect 2427 776 2653 784
rect 2727 776 2873 784
rect 2887 776 2913 784
rect 2936 784 2944 796
rect 3027 796 3073 804
rect 3087 796 3173 804
rect 3247 796 3333 804
rect 3516 804 3524 856
rect 3607 856 3753 864
rect 3776 856 3793 864
rect 3776 844 3784 856
rect 3816 847 3824 876
rect 4107 876 4173 884
rect 4187 876 4733 884
rect 3987 856 4013 864
rect 4047 856 4104 864
rect 3696 836 3784 844
rect 3547 816 3573 824
rect 3507 796 3524 804
rect 3696 804 3704 836
rect 3807 836 3813 844
rect 3836 824 3844 853
rect 3876 827 3884 853
rect 4096 847 4104 856
rect 4167 856 4204 864
rect 3967 836 4053 844
rect 3727 816 3844 824
rect 4116 824 4124 853
rect 4007 816 4124 824
rect 4056 807 4064 816
rect 3696 796 3753 804
rect 3787 796 3853 804
rect 2936 776 3413 784
rect 3467 776 4113 784
rect 4136 784 4144 833
rect 4196 827 4204 856
rect 4407 856 4493 864
rect 4516 856 4653 864
rect 4236 807 4244 833
rect 4256 824 4264 853
rect 4287 836 4313 844
rect 4327 836 4344 844
rect 4336 824 4344 836
rect 4367 836 4413 844
rect 4516 844 4524 856
rect 4707 856 4753 864
rect 4436 836 4524 844
rect 4436 827 4444 836
rect 4667 836 4713 844
rect 4776 844 4784 896
rect 4727 836 4784 844
rect 4256 816 4324 824
rect 4336 816 4373 824
rect 4136 776 4293 784
rect 4316 784 4324 816
rect 4487 816 4513 824
rect 4616 807 4624 833
rect 4636 824 4644 833
rect 4636 816 4664 824
rect 4656 807 4664 816
rect 4347 796 4393 804
rect 4427 796 4593 804
rect 4316 776 4393 784
rect 4567 776 4633 784
rect 4647 776 4693 784
rect 667 756 1653 764
rect 1707 756 2133 764
rect 2807 756 2953 764
rect 3067 756 3213 764
rect 3287 756 3373 764
rect 3687 756 4213 764
rect 4287 756 4373 764
rect 4447 756 4553 764
rect 4627 756 4673 764
rect 507 736 1433 744
rect 1947 736 2093 744
rect 2107 736 2373 744
rect 2967 736 3133 744
rect 3527 736 3553 744
rect 3647 736 4093 744
rect 4187 736 4213 744
rect 4247 736 4413 744
rect 4547 736 4713 744
rect 1247 716 1373 724
rect 2067 716 2173 724
rect 3007 716 3033 724
rect 3247 716 3353 724
rect 3387 716 3813 724
rect 3947 716 4673 724
rect 947 696 1193 704
rect 1347 696 1393 704
rect 1407 696 1673 704
rect 1847 696 1953 704
rect 2547 696 2573 704
rect 2667 696 3313 704
rect 3367 696 3453 704
rect 3527 696 3613 704
rect 3707 696 3873 704
rect 3887 696 4293 704
rect 4367 696 4593 704
rect 1027 676 1133 684
rect 1327 676 1353 684
rect 1367 676 1573 684
rect 1587 676 1873 684
rect 1907 676 2073 684
rect 2107 676 2233 684
rect 2247 676 2493 684
rect 2567 676 2653 684
rect 2847 676 2993 684
rect 3187 676 3333 684
rect 3347 676 3393 684
rect 3407 676 3433 684
rect 3447 676 3913 684
rect 4007 676 4613 684
rect 887 656 953 664
rect 1007 656 1053 664
rect 1087 656 1293 664
rect 1647 656 1773 664
rect 1787 656 1853 664
rect 1956 656 1973 664
rect 147 636 173 644
rect 327 636 393 644
rect 787 636 913 644
rect 1047 636 1073 644
rect 1107 636 1173 644
rect 1216 636 1273 644
rect 1216 627 1224 636
rect 1527 636 1593 644
rect 1807 636 1913 644
rect 1956 627 1964 656
rect 2387 656 2453 664
rect 2587 656 2693 664
rect 2707 656 2713 664
rect 2767 656 2853 664
rect 2947 656 3193 664
rect 3207 656 3293 664
rect 3327 656 3393 664
rect 3487 656 3604 664
rect 2067 636 2153 644
rect 2436 636 2613 644
rect 2436 627 2444 636
rect 167 616 213 624
rect 227 616 253 624
rect 387 616 433 624
rect 607 616 853 624
rect 907 616 953 624
rect 967 616 1173 624
rect 1036 607 1044 616
rect 2487 616 2513 624
rect 2736 624 2744 653
rect 2776 636 2873 644
rect 2776 627 2784 636
rect 2907 636 2944 644
rect 2736 616 2753 624
rect 2827 616 2913 624
rect 247 596 333 604
rect 467 596 593 604
rect 1927 596 2853 604
rect 2936 604 2944 636
rect 3087 636 3204 644
rect 2907 596 2944 604
rect 2956 604 2964 633
rect 3056 624 3064 633
rect 3196 627 3204 636
rect 3487 636 3584 644
rect 3056 616 3173 624
rect 3276 607 3284 633
rect 3416 624 3424 633
rect 3576 627 3584 636
rect 3416 616 3453 624
rect 3596 624 3604 656
rect 3776 656 3793 664
rect 3676 627 3684 653
rect 3716 627 3724 653
rect 3776 627 3784 656
rect 3947 656 4013 664
rect 4027 656 4053 664
rect 4087 656 4224 664
rect 3816 644 3824 653
rect 3807 636 3824 644
rect 3907 636 3953 644
rect 4027 636 4173 644
rect 4216 644 4224 656
rect 4247 656 4413 664
rect 4467 656 4513 664
rect 4607 656 4653 664
rect 4727 656 4753 664
rect 4216 636 4313 644
rect 4407 636 4453 644
rect 4507 636 4733 644
rect 3596 616 3664 624
rect 2956 596 3213 604
rect 3327 596 3353 604
rect 3467 596 3633 604
rect 3656 604 3664 616
rect 3907 616 3993 624
rect 4047 616 4073 624
rect 4087 616 4113 624
rect 4167 616 4253 624
rect 4387 616 4513 624
rect 4647 616 4693 624
rect 3656 596 3753 604
rect 3827 596 3873 604
rect 3927 596 4013 604
rect 4027 596 4053 604
rect 4147 596 4233 604
rect 4256 604 4264 613
rect 4256 596 4333 604
rect 4387 596 4473 604
rect 4487 596 4673 604
rect 2847 576 3053 584
rect 3747 576 4313 584
rect 4376 584 4384 593
rect 4327 576 4384 584
rect 4427 576 4753 584
rect 2747 556 3153 564
rect 3867 556 4173 564
rect 2787 536 3453 544
rect 3467 536 3533 544
rect 3727 536 3973 544
rect 4107 536 4533 544
rect 4067 516 4393 524
rect 4407 516 4433 524
rect 3187 476 3773 484
rect 2547 456 2693 464
rect 2767 456 3173 464
rect 3567 456 4353 464
rect 767 436 853 444
rect 2367 436 2773 444
rect 3367 436 3633 444
rect 87 416 753 424
rect 2647 416 2913 424
rect 3247 416 3853 424
rect 4567 416 4733 424
rect 187 396 273 404
rect 507 396 553 404
rect 647 396 793 404
rect 847 396 873 404
rect 1127 396 1193 404
rect 1207 396 1373 404
rect 1507 396 1593 404
rect 1607 396 2393 404
rect 2407 396 2513 404
rect 2527 396 2633 404
rect 2907 396 2993 404
rect 3047 396 3073 404
rect 3167 396 3193 404
rect 3287 396 3433 404
rect 3567 396 3613 404
rect 3627 396 3693 404
rect 3987 396 4093 404
rect 4307 396 4333 404
rect 4527 396 4753 404
rect 547 376 573 384
rect 596 376 753 384
rect 287 356 353 364
rect 476 364 484 373
rect 596 367 604 376
rect 807 376 1093 384
rect 1127 376 1133 384
rect 1147 376 1333 384
rect 1567 376 1653 384
rect 1747 376 1893 384
rect 1947 376 2053 384
rect 2147 376 2553 384
rect 2567 376 2593 384
rect 2867 376 3273 384
rect 3327 376 3353 384
rect 3916 376 3973 384
rect 476 356 513 364
rect 747 356 804 364
rect 127 336 373 344
rect 396 344 404 353
rect 396 336 613 344
rect 696 344 704 353
rect 667 336 773 344
rect 796 344 804 356
rect 847 356 933 364
rect 947 356 993 364
rect 1167 356 1233 364
rect 1527 356 1573 364
rect 2027 356 2313 364
rect 2427 356 2453 364
rect 2547 356 2793 364
rect 3056 356 3113 364
rect 796 336 833 344
rect 967 336 1013 344
rect 1107 336 1133 344
rect 1327 336 1453 344
rect 487 316 653 324
rect 687 316 753 324
rect 767 316 953 324
rect 967 316 1293 324
rect 1476 324 1484 353
rect 1507 336 1773 344
rect 2007 336 2133 344
rect 2316 344 2324 353
rect 2316 336 2353 344
rect 2727 336 2833 344
rect 1427 316 1484 324
rect 1767 316 2173 324
rect 2187 316 2213 324
rect 2287 316 2333 324
rect 2427 316 2893 324
rect 2956 324 2964 353
rect 3056 347 3064 356
rect 3267 356 3373 364
rect 3427 356 3473 364
rect 3207 336 3393 344
rect 2956 316 3033 324
rect 3107 316 3133 324
rect 3516 324 3524 373
rect 3596 347 3604 373
rect 3916 347 3924 376
rect 3987 376 4113 384
rect 4287 376 4313 384
rect 4587 376 4613 384
rect 3667 336 3713 344
rect 4007 336 4033 344
rect 3507 316 3673 324
rect 3887 316 3933 324
rect 4156 324 4164 353
rect 4236 347 4244 373
rect 4267 356 4353 364
rect 4447 356 4493 364
rect 4547 356 4593 364
rect 4287 336 4344 344
rect 4336 327 4344 336
rect 4387 336 4553 344
rect 4156 316 4313 324
rect 4567 316 4633 324
rect 587 296 813 304
rect 847 296 1053 304
rect 1227 296 1353 304
rect 2227 296 2573 304
rect 2587 296 2673 304
rect 2687 296 2813 304
rect 2887 296 3233 304
rect 3247 296 3333 304
rect 3367 296 3553 304
rect 3567 296 3573 304
rect 3627 296 3653 304
rect 3687 296 4113 304
rect 4227 296 4413 304
rect 4427 296 4533 304
rect 4656 304 4664 353
rect 4607 296 4664 304
rect 247 276 373 284
rect 387 276 433 284
rect 447 276 453 284
rect 1027 276 1253 284
rect 1267 276 1613 284
rect 2987 276 3053 284
rect 3227 276 3533 284
rect 3807 276 3993 284
rect 4187 276 4233 284
rect 4247 276 4553 284
rect 4567 276 4573 284
rect 3767 256 4653 264
rect 1127 236 1153 244
rect 1707 236 2273 244
rect 3587 236 3593 244
rect 3607 236 3813 244
rect 3827 236 4033 244
rect 247 216 333 224
rect 447 216 513 224
rect 647 216 753 224
rect 767 216 1333 224
rect 1387 216 1513 224
rect 1527 216 2113 224
rect 2287 216 2373 224
rect 3567 216 3753 224
rect 3847 216 3893 224
rect 4007 216 4053 224
rect 4107 216 4233 224
rect 4267 216 4393 224
rect 347 196 553 204
rect 627 196 713 204
rect 727 196 1173 204
rect 1187 196 1233 204
rect 1507 196 1553 204
rect 1567 196 1653 204
rect 1667 196 2193 204
rect 2247 196 2293 204
rect 2327 196 2353 204
rect 2387 196 2433 204
rect 2627 196 2933 204
rect 3047 196 3213 204
rect 3327 196 3353 204
rect 3467 196 3633 204
rect 3656 196 3733 204
rect 327 176 353 184
rect 427 176 493 184
rect 527 176 673 184
rect 1147 176 1193 184
rect 1287 176 1393 184
rect 1447 176 1533 184
rect 1896 176 2033 184
rect 1896 167 1904 176
rect 2047 176 2093 184
rect 2116 176 2164 184
rect 187 156 253 164
rect 276 156 293 164
rect 276 144 284 156
rect 367 156 704 164
rect 696 147 704 156
rect 827 156 1033 164
rect 1636 156 1693 164
rect 127 136 284 144
rect 327 136 433 144
rect 507 136 544 144
rect 287 116 353 124
rect 536 124 544 136
rect 1067 136 1153 144
rect 1216 144 1224 153
rect 1636 147 1644 156
rect 1767 156 1813 164
rect 2116 164 2124 176
rect 1916 156 2124 164
rect 1216 136 1413 144
rect 1916 144 1924 156
rect 2156 164 2164 176
rect 2227 176 2413 184
rect 2427 176 2953 184
rect 3167 176 3253 184
rect 3307 176 3413 184
rect 3656 184 3664 196
rect 3747 196 4073 204
rect 4227 196 4473 204
rect 3507 176 3664 184
rect 3687 176 3713 184
rect 3887 176 3933 184
rect 4067 176 4153 184
rect 4327 176 4393 184
rect 4707 176 4773 184
rect 2156 156 2233 164
rect 2387 156 2493 164
rect 2867 156 2993 164
rect 3187 156 3273 164
rect 3447 156 3693 164
rect 3747 156 3813 164
rect 3867 156 3904 164
rect 1687 136 1924 144
rect 2136 144 2144 153
rect 2136 136 2473 144
rect 2487 136 2733 144
rect 2887 136 2973 144
rect 3027 136 3293 144
rect 3407 136 3453 144
rect 487 116 524 124
rect 536 116 813 124
rect 516 104 524 116
rect 1167 116 1353 124
rect 1407 116 1673 124
rect 1807 116 1933 124
rect 516 96 773 104
rect 787 96 973 104
rect 1307 96 1473 104
rect 1956 104 1964 133
rect 2007 116 2053 124
rect 2067 116 2153 124
rect 3067 116 3093 124
rect 3287 116 3333 124
rect 3487 116 3533 124
rect 3816 124 3824 153
rect 3896 147 3904 156
rect 3967 156 3993 164
rect 4087 156 4353 164
rect 4087 136 4104 144
rect 4096 127 4104 136
rect 4267 136 4344 144
rect 4336 127 4344 136
rect 4447 136 4513 144
rect 4456 127 4464 136
rect 4687 136 4753 144
rect 3816 116 4013 124
rect 4147 116 4153 124
rect 4167 116 4193 124
rect 4247 116 4293 124
rect 4507 116 4593 124
rect 1927 96 1964 104
rect 3207 96 3253 104
rect 3267 96 3373 104
rect 3387 96 3573 104
rect 3787 96 3833 104
rect 4416 104 4424 113
rect 4416 96 4493 104
rect 3627 76 3893 84
rect 2787 56 3613 64
rect 2707 36 3573 44
rect 3987 36 4173 44
rect 3087 16 3493 24
rect 3807 16 4133 24
rect 4227 16 4613 24
<< m1p >>
rect 4 4562 4736 4578
rect 4 4322 4776 4338
rect 4 4082 4756 4098
rect 4 3842 4776 3858
rect 4 3602 4756 3618
rect 4 3362 4776 3378
rect 4 3122 4776 3138
rect 4 2882 4776 2898
rect 4 2642 4736 2658
rect 4 2402 4776 2418
rect 4 2162 4776 2178
rect 4 1922 4776 1938
rect 4 1682 4736 1698
rect 4 1442 4776 1458
rect 4 1202 4776 1218
rect 4 962 4776 978
rect 4 722 4776 738
rect 4 482 4776 498
rect 4 242 4756 258
rect 4 2 4776 18
<< m2p >>
rect 393 4493 407 4507
rect 473 4493 487 4507
rect 633 4493 647 4507
rect 673 4493 687 4507
rect 733 4493 747 4507
rect 2393 4493 2407 4507
rect 2433 4493 2447 4507
rect 2533 4493 2547 4507
rect 3373 4493 3387 4507
rect 3453 4493 3467 4507
rect 3713 4493 3727 4507
rect 4213 4493 4227 4507
rect 4433 4493 4447 4507
rect 4513 4493 4527 4507
rect 33 4473 47 4487
rect 73 4473 87 4487
rect 213 4473 227 4487
rect 253 4473 267 4487
rect 273 4473 287 4487
rect 313 4473 327 4487
rect 373 4473 387 4487
rect 413 4473 427 4487
rect 453 4473 467 4487
rect 493 4473 507 4487
rect 513 4473 527 4487
rect 553 4473 567 4487
rect 653 4473 667 4487
rect 693 4473 707 4487
rect 813 4473 827 4487
rect 893 4473 907 4487
rect 933 4473 947 4487
rect 1033 4473 1047 4487
rect 1073 4473 1087 4487
rect 1153 4473 1167 4487
rect 1233 4473 1247 4487
rect 1273 4473 1287 4487
rect 1373 4473 1387 4487
rect 1413 4473 1427 4487
rect 1553 4473 1567 4487
rect 1593 4473 1607 4487
rect 1673 4473 1687 4487
rect 1813 4473 1827 4487
rect 1893 4473 1907 4487
rect 1933 4473 1947 4487
rect 2033 4473 2047 4487
rect 2073 4473 2087 4487
rect 2113 4473 2127 4487
rect 2293 4473 2307 4487
rect 2333 4473 2347 4487
rect 2413 4473 2427 4487
rect 2453 4473 2467 4487
rect 2553 4473 2567 4487
rect 2593 4473 2607 4487
rect 2653 4473 2667 4487
rect 2693 4473 2707 4487
rect 2733 4473 2747 4487
rect 2773 4473 2787 4487
rect 2833 4473 2847 4487
rect 2873 4473 2887 4487
rect 3013 4473 3027 4487
rect 3073 4473 3087 4487
rect 3113 4473 3127 4487
rect 3153 4473 3167 4487
rect 3413 4473 3427 4487
rect 3753 4473 3767 4487
rect 3793 4473 3807 4487
rect 3833 4473 3847 4487
rect 3933 4473 3947 4487
rect 3973 4473 3987 4487
rect 4253 4473 4267 4487
rect 4393 4473 4407 4487
rect 133 4453 147 4467
rect 193 4453 207 4467
rect 233 4453 247 4467
rect 613 4453 627 4467
rect 753 4453 767 4467
rect 1053 4453 1067 4467
rect 1093 4453 1107 4467
rect 1393 4453 1407 4467
rect 1433 4453 1447 4467
rect 1733 4453 1747 4467
rect 2053 4453 2067 4467
rect 2093 4453 2107 4467
rect 2193 4453 2207 4467
rect 2233 4453 2247 4467
rect 2273 4453 2287 4467
rect 2313 4453 2327 4467
rect 2373 4453 2387 4467
rect 2513 4453 2527 4467
rect 2573 4453 2587 4467
rect 2613 4453 2627 4467
rect 2933 4453 2947 4467
rect 2973 4453 2987 4467
rect 3213 4453 3227 4467
rect 3253 4453 3267 4467
rect 3293 4453 3307 4467
rect 3353 4453 3367 4467
rect 3393 4453 3407 4467
rect 3473 4453 3487 4467
rect 3533 4453 3547 4467
rect 3593 4453 3607 4467
rect 3633 4453 3647 4467
rect 3693 4453 3707 4467
rect 3733 4453 3747 4467
rect 3813 4453 3827 4467
rect 3853 4453 3867 4467
rect 3913 4453 3927 4467
rect 3953 4453 3967 4467
rect 4033 4453 4047 4467
rect 4073 4453 4087 4467
rect 4133 4453 4147 4467
rect 4173 4453 4187 4467
rect 4193 4453 4207 4467
rect 4233 4453 4247 4467
rect 4313 4453 4327 4467
rect 4413 4453 4427 4467
rect 4453 4453 4467 4467
rect 4493 4453 4507 4467
rect 4533 4453 4547 4467
rect 4573 4453 4587 4467
rect 4633 4453 4647 4467
rect 4673 4453 4687 4467
rect 113 4433 127 4447
rect 153 4433 167 4447
rect 1713 4433 1727 4447
rect 1753 4433 1767 4447
rect 2173 4433 2187 4447
rect 2213 4433 2227 4447
rect 2913 4433 2927 4447
rect 2953 4433 2967 4447
rect 3033 4433 3047 4447
rect 3193 4433 3207 4447
rect 3233 4433 3247 4447
rect 3273 4433 3287 4447
rect 3313 4433 3327 4447
rect 3513 4433 3527 4447
rect 3553 4433 3567 4447
rect 3613 4433 3627 4447
rect 3653 4433 3667 4447
rect 4013 4433 4027 4447
rect 4053 4433 4067 4447
rect 4113 4433 4127 4447
rect 4153 4433 4167 4447
rect 4293 4433 4307 4447
rect 4333 4433 4347 4447
rect 4553 4433 4567 4447
rect 4593 4433 4607 4447
rect 4653 4433 4667 4447
rect 4693 4433 4707 4447
rect 153 4213 167 4227
rect 433 4213 447 4227
rect 613 4213 627 4227
rect 653 4213 667 4227
rect 833 4213 847 4227
rect 2093 4213 2107 4227
rect 2133 4213 2147 4227
rect 2373 4213 2387 4227
rect 2413 4213 2427 4227
rect 2933 4213 2947 4227
rect 2973 4213 2987 4227
rect 3033 4213 3047 4227
rect 3073 4213 3087 4227
rect 3113 4213 3127 4227
rect 3153 4213 3167 4227
rect 3273 4213 3287 4227
rect 3313 4213 3327 4227
rect 3373 4213 3387 4227
rect 3413 4213 3427 4227
rect 3473 4213 3487 4227
rect 3513 4213 3527 4227
rect 3573 4213 3587 4227
rect 3613 4213 3627 4227
rect 3673 4213 3687 4227
rect 3713 4213 3727 4227
rect 4133 4213 4147 4227
rect 4173 4213 4187 4227
rect 4233 4213 4247 4227
rect 4273 4213 4287 4227
rect 33 4193 47 4207
rect 73 4193 87 4207
rect 333 4193 347 4207
rect 373 4193 387 4207
rect 533 4193 547 4207
rect 573 4193 587 4207
rect 593 4193 607 4207
rect 633 4193 647 4207
rect 693 4193 707 4207
rect 733 4193 747 4207
rect 913 4193 927 4207
rect 953 4193 967 4207
rect 1013 4193 1027 4207
rect 1313 4193 1327 4207
rect 1613 4193 1627 4207
rect 1653 4193 1667 4207
rect 1793 4193 1807 4207
rect 2113 4193 2127 4207
rect 2213 4193 2227 4207
rect 2293 4193 2307 4207
rect 2333 4193 2347 4207
rect 2393 4193 2407 4207
rect 2473 4193 2487 4207
rect 2513 4193 2527 4207
rect 2633 4193 2647 4207
rect 2673 4193 2687 4207
rect 2773 4193 2787 4207
rect 2813 4193 2827 4207
rect 2953 4193 2967 4207
rect 2993 4193 3007 4207
rect 3053 4193 3067 4207
rect 3093 4193 3107 4207
rect 3133 4193 3147 4207
rect 3213 4193 3227 4207
rect 3293 4193 3307 4207
rect 3333 4193 3347 4207
rect 3393 4193 3407 4207
rect 3433 4193 3447 4207
rect 3493 4193 3507 4207
rect 3533 4193 3547 4207
rect 3593 4193 3607 4207
rect 3633 4193 3647 4207
rect 3653 4193 3667 4207
rect 3693 4193 3707 4207
rect 3753 4193 3767 4207
rect 3793 4193 3807 4207
rect 3873 4193 3887 4207
rect 3913 4193 3927 4207
rect 3973 4193 3987 4207
rect 4013 4193 4027 4207
rect 4053 4193 4067 4207
rect 4153 4193 4167 4207
rect 4193 4193 4207 4207
rect 4213 4193 4227 4207
rect 4253 4193 4267 4207
rect 4313 4193 4327 4207
rect 4353 4193 4367 4207
rect 4433 4193 4447 4207
rect 4473 4193 4487 4207
rect 4533 4193 4547 4207
rect 4573 4193 4587 4207
rect 53 4173 67 4187
rect 93 4173 107 4187
rect 133 4173 147 4187
rect 193 4173 207 4187
rect 213 4173 227 4187
rect 253 4173 267 4187
rect 313 4173 327 4187
rect 393 4173 407 4187
rect 453 4173 467 4187
rect 513 4173 527 4187
rect 753 4173 767 4187
rect 793 4173 807 4187
rect 853 4173 867 4187
rect 933 4173 947 4187
rect 973 4173 987 4187
rect 1053 4173 1067 4187
rect 1093 4173 1107 4187
rect 1133 4173 1147 4187
rect 1173 4173 1187 4187
rect 1213 4173 1227 4187
rect 1253 4173 1267 4187
rect 1373 4173 1387 4187
rect 1453 4173 1467 4187
rect 1493 4173 1507 4187
rect 1593 4173 1607 4187
rect 1633 4173 1647 4187
rect 1693 4173 1707 4187
rect 1733 4173 1747 4187
rect 1853 4173 1867 4187
rect 1933 4173 1947 4187
rect 1973 4173 1987 4187
rect 2173 4173 2187 4187
rect 2273 4173 2287 4187
rect 2313 4173 2327 4187
rect 2353 4173 2367 4187
rect 2493 4173 2507 4187
rect 2533 4173 2547 4187
rect 2573 4173 2587 4187
rect 2613 4173 2627 4187
rect 2693 4173 2707 4187
rect 2753 4173 2767 4187
rect 2833 4173 2847 4187
rect 2873 4173 2887 4187
rect 3813 4173 3827 4187
rect 3853 4173 3867 4187
rect 3893 4173 3907 4187
rect 4073 4173 4087 4187
rect 4373 4173 4387 4187
rect 4413 4173 4427 4187
rect 4453 4173 4467 4187
rect 4513 4173 4527 4187
rect 4553 4173 4567 4187
rect 4593 4173 4607 4187
rect 4653 4173 4667 4187
rect 4693 4173 4707 4187
rect 233 4153 247 4167
rect 353 4153 367 4167
rect 553 4153 567 4167
rect 713 4153 727 4167
rect 1033 4153 1047 4167
rect 1073 4153 1087 4167
rect 1153 4153 1167 4167
rect 1233 4153 1247 4167
rect 1293 4153 1307 4167
rect 1713 4153 1727 4167
rect 1813 4153 1827 4167
rect 2153 4153 2167 4167
rect 2593 4153 2607 4167
rect 2653 4153 2667 4167
rect 2793 4153 2807 4167
rect 3233 4153 3247 4167
rect 3773 4153 3787 4167
rect 3953 4153 3967 4167
rect 4033 4153 4047 4167
rect 4333 4153 4347 4167
rect 4673 4153 4687 4167
rect 213 4013 227 4027
rect 393 4013 407 4027
rect 453 4013 467 4027
rect 513 4013 527 4027
rect 753 4013 767 4027
rect 1033 4013 1047 4027
rect 1093 4013 1107 4027
rect 1133 4013 1147 4027
rect 1213 4013 1227 4027
rect 1273 4013 1287 4027
rect 1373 4013 1387 4027
rect 1453 4013 1467 4027
rect 1833 4013 1847 4027
rect 2113 4013 2127 4027
rect 2393 4013 2407 4027
rect 2473 4013 2487 4027
rect 2753 4013 2767 4027
rect 3133 4013 3147 4027
rect 3273 4013 3287 4027
rect 3713 4013 3727 4027
rect 4433 4013 4447 4027
rect 4673 4013 4687 4027
rect 193 3993 207 4007
rect 233 3993 247 4007
rect 253 3993 267 4007
rect 293 3993 307 4007
rect 493 3993 507 4007
rect 533 3993 547 4007
rect 553 3993 567 4007
rect 613 3993 627 4007
rect 653 3993 667 4007
rect 693 3993 707 4007
rect 813 3993 827 4007
rect 853 3993 867 4007
rect 1073 3993 1087 4007
rect 1113 3993 1127 4007
rect 1193 3993 1207 4007
rect 1233 3993 1247 4007
rect 1353 3993 1367 4007
rect 1393 3993 1407 4007
rect 1473 3993 1487 4007
rect 1513 3993 1527 4007
rect 1573 3993 1587 4007
rect 1613 3993 1627 4007
rect 1653 3993 1667 4007
rect 1793 3993 1807 4007
rect 2013 3993 2027 4007
rect 2053 3993 2067 4007
rect 2353 3993 2367 4007
rect 2533 3993 2547 4007
rect 2573 3993 2587 4007
rect 2713 3993 2727 4007
rect 2833 3993 2847 4007
rect 2873 3993 2887 4007
rect 2893 3993 2907 4007
rect 2933 3993 2947 4007
rect 3153 3993 3167 4007
rect 3193 3993 3207 4007
rect 3313 3993 3327 4007
rect 3353 3993 3367 4007
rect 3393 3993 3407 4007
rect 3493 3993 3507 4007
rect 3533 3993 3547 4007
rect 3593 3993 3607 4007
rect 3633 3993 3647 4007
rect 3673 3993 3687 4007
rect 4233 3993 4247 4007
rect 4273 3993 4287 4007
rect 4293 3993 4307 4007
rect 4333 3993 4347 4007
rect 4713 3993 4727 4007
rect 53 3973 67 3987
rect 133 3973 147 3987
rect 273 3973 287 3987
rect 313 3973 327 3987
rect 373 3973 387 3987
rect 433 3973 447 3987
rect 673 3973 687 3987
rect 713 3973 727 3987
rect 773 3973 787 3987
rect 833 3973 847 3987
rect 873 3973 887 3987
rect 933 3973 947 3987
rect 1013 3973 1027 3987
rect 1153 3973 1167 3987
rect 1293 3973 1307 3987
rect 1433 3973 1447 3987
rect 1493 3973 1507 3987
rect 1533 3973 1547 3987
rect 1593 3973 1607 3987
rect 1633 3973 1647 3987
rect 1713 3973 1727 3987
rect 1813 3973 1827 3987
rect 1853 3973 1867 3987
rect 1873 3973 1887 3987
rect 1913 3973 1927 3987
rect 1993 3973 2007 3987
rect 2033 3973 2047 3987
rect 2093 3973 2107 3987
rect 2173 3973 2187 3987
rect 2213 3973 2227 3987
rect 2273 3973 2287 3987
rect 2313 3973 2327 3987
rect 2373 3973 2387 3987
rect 2413 3973 2427 3987
rect 2453 3973 2467 3987
rect 2513 3973 2527 3987
rect 2553 3973 2567 3987
rect 2633 3973 2647 3987
rect 2673 3973 2687 3987
rect 2733 3973 2747 3987
rect 2773 3973 2787 3987
rect 2813 3973 2827 3987
rect 2853 3973 2867 3987
rect 2913 3973 2927 3987
rect 2953 3973 2967 3987
rect 3033 3973 3047 3987
rect 3073 3973 3087 3987
rect 3113 3973 3127 3987
rect 3173 3973 3187 3987
rect 3213 3973 3227 3987
rect 3253 3973 3267 3987
rect 3293 3973 3307 3987
rect 3373 3973 3387 3987
rect 3413 3973 3427 3987
rect 3473 3973 3487 3987
rect 3513 3973 3527 3987
rect 3573 3973 3587 3987
rect 3613 3973 3627 3987
rect 3693 3973 3707 3987
rect 3733 3973 3747 3987
rect 3793 3973 3807 3987
rect 3833 3973 3847 3987
rect 3893 3973 3907 3987
rect 3973 3973 3987 3987
rect 4033 3973 4047 3987
rect 4133 3973 4147 3987
rect 4173 3973 4187 3987
rect 4213 3973 4227 3987
rect 4253 3973 4267 3987
rect 4313 3973 4327 3987
rect 4353 3973 4367 3987
rect 4413 3973 4427 3987
rect 4493 3973 4507 3987
rect 4533 3973 4547 3987
rect 4593 3973 4607 3987
rect 4633 3973 4647 3987
rect 4653 3973 4667 3987
rect 4693 3973 4707 3987
rect 33 3953 47 3967
rect 73 3953 87 3967
rect 113 3953 127 3967
rect 153 3953 167 3967
rect 593 3953 607 3967
rect 913 3953 927 3967
rect 953 3953 967 3967
rect 1693 3953 1707 3967
rect 1733 3953 1747 3967
rect 1893 3953 1907 3967
rect 1933 3953 1947 3967
rect 2153 3953 2167 3967
rect 2193 3953 2207 3967
rect 2253 3953 2267 3967
rect 2293 3953 2307 3967
rect 2613 3953 2627 3967
rect 2653 3953 2667 3967
rect 3013 3953 3027 3967
rect 3053 3953 3067 3967
rect 3773 3953 3787 3967
rect 3813 3953 3827 3967
rect 3873 3953 3887 3967
rect 3913 3953 3927 3967
rect 3953 3953 3967 3967
rect 3993 3953 4007 3967
rect 4013 3953 4027 3967
rect 4053 3953 4067 3967
rect 4113 3953 4127 3967
rect 4153 3953 4167 3967
rect 4473 3953 4487 3967
rect 4513 3953 4527 3967
rect 4573 3953 4587 3967
rect 4613 3953 4627 3967
rect 553 3733 567 3747
rect 733 3733 747 3747
rect 773 3733 787 3747
rect 1453 3733 1467 3747
rect 1493 3733 1507 3747
rect 1533 3733 1547 3747
rect 1573 3733 1587 3747
rect 2173 3733 2187 3747
rect 2213 3733 2227 3747
rect 2373 3733 2387 3747
rect 2413 3733 2427 3747
rect 2573 3733 2587 3747
rect 2613 3733 2627 3747
rect 2993 3733 3007 3747
rect 3033 3733 3047 3747
rect 3193 3733 3207 3747
rect 3233 3733 3247 3747
rect 3453 3733 3467 3747
rect 3493 3733 3507 3747
rect 3553 3733 3567 3747
rect 3733 3733 3747 3747
rect 3773 3733 3787 3747
rect 4393 3733 4407 3747
rect 4433 3733 4447 3747
rect 4553 3733 4567 3747
rect 4593 3733 4607 3747
rect 4653 3733 4667 3747
rect 4693 3733 4707 3747
rect 33 3713 47 3727
rect 73 3713 87 3727
rect 133 3713 147 3727
rect 433 3713 447 3727
rect 473 3713 487 3727
rect 633 3713 647 3727
rect 753 3713 767 3727
rect 1373 3713 1387 3727
rect 1413 3713 1427 3727
rect 1473 3713 1487 3727
rect 1553 3713 1567 3727
rect 1953 3713 1967 3727
rect 2033 3713 2047 3727
rect 2073 3713 2087 3727
rect 2113 3713 2127 3727
rect 2153 3713 2167 3727
rect 2193 3713 2207 3727
rect 2273 3713 2287 3727
rect 2313 3713 2327 3727
rect 2393 3713 2407 3727
rect 2433 3713 2447 3727
rect 2493 3713 2507 3727
rect 2533 3713 2547 3727
rect 2593 3713 2607 3727
rect 2633 3713 2647 3727
rect 2653 3713 2667 3727
rect 2693 3713 2707 3727
rect 2793 3713 2807 3727
rect 2833 3713 2847 3727
rect 2873 3713 2887 3727
rect 2933 3713 2947 3727
rect 3013 3713 3027 3727
rect 3053 3713 3067 3727
rect 3113 3713 3127 3727
rect 3153 3713 3167 3727
rect 3213 3713 3227 3727
rect 3253 3713 3267 3727
rect 3293 3713 3307 3727
rect 3353 3713 3367 3727
rect 3393 3713 3407 3727
rect 3473 3713 3487 3727
rect 3653 3713 3667 3727
rect 3693 3713 3707 3727
rect 3753 3713 3767 3727
rect 3793 3713 3807 3727
rect 3833 3713 3847 3727
rect 3873 3713 3887 3727
rect 3913 3713 3927 3727
rect 3993 3713 4007 3727
rect 4033 3713 4047 3727
rect 4093 3713 4107 3727
rect 4133 3713 4147 3727
rect 4173 3713 4187 3727
rect 4213 3713 4227 3727
rect 4313 3713 4327 3727
rect 4353 3713 4367 3727
rect 4373 3713 4387 3727
rect 4413 3713 4427 3727
rect 4493 3713 4507 3727
rect 4573 3713 4587 3727
rect 4613 3713 4627 3727
rect 4633 3713 4647 3727
rect 4673 3713 4687 3727
rect 53 3693 67 3707
rect 93 3693 107 3707
rect 193 3693 207 3707
rect 273 3693 287 3707
rect 313 3693 327 3707
rect 453 3693 467 3707
rect 493 3693 507 3707
rect 513 3693 527 3707
rect 573 3693 587 3707
rect 673 3693 687 3707
rect 873 3693 887 3707
rect 913 3693 927 3707
rect 993 3693 1007 3707
rect 1053 3693 1067 3707
rect 1093 3693 1107 3707
rect 1133 3693 1147 3707
rect 1213 3693 1227 3707
rect 1253 3693 1267 3707
rect 1353 3693 1367 3707
rect 1393 3693 1407 3707
rect 1613 3693 1627 3707
rect 1653 3693 1667 3707
rect 1713 3693 1727 3707
rect 1793 3693 1807 3707
rect 1833 3693 1847 3707
rect 2013 3693 2027 3707
rect 2293 3693 2307 3707
rect 2333 3693 2347 3707
rect 2473 3693 2487 3707
rect 2713 3693 2727 3707
rect 2773 3693 2787 3707
rect 3093 3693 3107 3707
rect 3373 3693 3387 3707
rect 3413 3693 3427 3707
rect 3513 3693 3527 3707
rect 3573 3693 3587 3707
rect 3633 3693 3647 3707
rect 3933 3693 3947 3707
rect 4013 3693 4027 3707
rect 4053 3693 4067 3707
rect 4073 3693 4087 3707
rect 4113 3693 4127 3707
rect 4233 3693 4247 3707
rect 4293 3693 4307 3707
rect 153 3673 167 3687
rect 693 3673 707 3687
rect 1973 3673 1987 3687
rect 2053 3673 2067 3687
rect 2133 3673 2147 3687
rect 2513 3673 2527 3687
rect 2673 3673 2687 3687
rect 2813 3673 2827 3687
rect 2893 3673 2907 3687
rect 2953 3673 2967 3687
rect 3133 3673 3147 3687
rect 3313 3673 3327 3687
rect 3673 3673 3687 3687
rect 3853 3673 3867 3687
rect 3893 3673 3907 3687
rect 4193 3673 4207 3687
rect 4333 3673 4347 3687
rect 4513 3673 4527 3687
rect 653 3533 667 3547
rect 873 3533 887 3547
rect 973 3533 987 3547
rect 1253 3533 1267 3547
rect 1333 3533 1347 3547
rect 1693 3533 1707 3547
rect 2213 3533 2227 3547
rect 2393 3533 2407 3547
rect 3013 3533 3027 3547
rect 3553 3533 3567 3547
rect 3893 3533 3907 3547
rect 4413 3533 4427 3547
rect 4493 3533 4507 3547
rect 93 3513 107 3527
rect 133 3513 147 3527
rect 213 3513 227 3527
rect 373 3513 387 3527
rect 413 3513 427 3527
rect 713 3513 727 3527
rect 753 3513 767 3527
rect 813 3513 827 3527
rect 853 3513 867 3527
rect 953 3513 967 3527
rect 993 3513 1007 3527
rect 1033 3513 1047 3527
rect 1113 3513 1127 3527
rect 1153 3513 1167 3527
rect 1313 3513 1327 3527
rect 1353 3513 1367 3527
rect 1393 3513 1407 3527
rect 1433 3513 1447 3527
rect 1593 3513 1607 3527
rect 1633 3513 1647 3527
rect 1733 3513 1747 3527
rect 1813 3513 1827 3527
rect 1853 3513 1867 3527
rect 1953 3513 1967 3527
rect 1993 3513 2007 3527
rect 2033 3513 2047 3527
rect 2173 3513 2187 3527
rect 2653 3513 2667 3527
rect 2693 3513 2707 3527
rect 2713 3513 2727 3527
rect 2753 3513 2767 3527
rect 2893 3513 2907 3527
rect 2933 3513 2947 3527
rect 2993 3513 3007 3527
rect 3033 3513 3047 3527
rect 3113 3513 3127 3527
rect 3153 3513 3167 3527
rect 3173 3513 3187 3527
rect 3213 3513 3227 3527
rect 3253 3513 3267 3527
rect 3533 3513 3547 3527
rect 3573 3513 3587 3527
rect 3873 3513 3887 3527
rect 3913 3513 3927 3527
rect 4093 3513 4107 3527
rect 4133 3513 4147 3527
rect 4453 3513 4467 3527
rect 293 3493 307 3507
rect 353 3493 367 3507
rect 393 3493 407 3507
rect 473 3493 487 3507
rect 553 3493 567 3507
rect 593 3493 607 3507
rect 633 3493 647 3507
rect 693 3493 707 3507
rect 733 3493 747 3507
rect 793 3493 807 3507
rect 833 3493 847 3507
rect 893 3493 907 3507
rect 1273 3493 1287 3507
rect 1413 3493 1427 3507
rect 1453 3493 1467 3507
rect 1513 3493 1527 3507
rect 1673 3493 1687 3507
rect 1973 3493 1987 3507
rect 2013 3493 2027 3507
rect 2093 3493 2107 3507
rect 2193 3493 2207 3507
rect 2233 3493 2247 3507
rect 2293 3493 2307 3507
rect 2333 3493 2347 3507
rect 2373 3493 2387 3507
rect 2453 3493 2467 3507
rect 2493 3493 2507 3507
rect 2553 3493 2567 3507
rect 2593 3493 2607 3507
rect 2633 3493 2647 3507
rect 2673 3493 2687 3507
rect 2733 3493 2747 3507
rect 2773 3493 2787 3507
rect 2833 3493 2847 3507
rect 2913 3493 2927 3507
rect 2953 3493 2967 3507
rect 3093 3493 3107 3507
rect 3133 3493 3147 3507
rect 3193 3493 3207 3507
rect 3233 3493 3247 3507
rect 3313 3493 3327 3507
rect 3393 3493 3407 3507
rect 3473 3493 3487 3507
rect 3633 3493 3647 3507
rect 3713 3493 3727 3507
rect 3813 3493 3827 3507
rect 3953 3493 3967 3507
rect 4033 3493 4047 3507
rect 4113 3493 4127 3507
rect 4153 3493 4167 3507
rect 4233 3493 4247 3507
rect 4273 3493 4287 3507
rect 4293 3493 4307 3507
rect 4333 3493 4347 3507
rect 4393 3493 4407 3507
rect 4433 3493 4447 3507
rect 4513 3493 4527 3507
rect 4593 3493 4607 3507
rect 4633 3493 4647 3507
rect 4653 3493 4667 3507
rect 4693 3493 4707 3507
rect 273 3473 287 3487
rect 313 3473 327 3487
rect 453 3473 467 3487
rect 493 3473 507 3487
rect 533 3473 547 3487
rect 573 3473 587 3487
rect 1493 3473 1507 3487
rect 1533 3473 1547 3487
rect 2073 3473 2087 3487
rect 2113 3473 2127 3487
rect 2273 3473 2287 3487
rect 2313 3473 2327 3487
rect 2433 3473 2447 3487
rect 2473 3473 2487 3487
rect 2533 3473 2547 3487
rect 2573 3473 2587 3487
rect 2813 3473 2827 3487
rect 2853 3473 2867 3487
rect 3293 3473 3307 3487
rect 3333 3473 3347 3487
rect 3373 3473 3387 3487
rect 3413 3473 3427 3487
rect 3453 3473 3467 3487
rect 3493 3473 3507 3487
rect 3613 3473 3627 3487
rect 3653 3473 3667 3487
rect 3693 3473 3707 3487
rect 3733 3473 3747 3487
rect 3793 3473 3807 3487
rect 3833 3473 3847 3487
rect 3933 3473 3947 3487
rect 3973 3473 3987 3487
rect 4013 3473 4027 3487
rect 4053 3473 4067 3487
rect 4213 3473 4227 3487
rect 4253 3473 4267 3487
rect 4313 3473 4327 3487
rect 4353 3473 4367 3487
rect 4573 3473 4587 3487
rect 4613 3473 4627 3487
rect 4673 3473 4687 3487
rect 4713 3473 4727 3487
rect 373 3253 387 3267
rect 413 3253 427 3267
rect 673 3253 687 3267
rect 713 3253 727 3267
rect 2433 3253 2447 3267
rect 2473 3253 2487 3267
rect 2953 3253 2967 3267
rect 2993 3253 3007 3267
rect 3033 3253 3047 3267
rect 3073 3253 3087 3267
rect 3233 3253 3247 3267
rect 3273 3253 3287 3267
rect 3453 3253 3467 3267
rect 3513 3253 3527 3267
rect 3553 3253 3567 3267
rect 3633 3253 3647 3267
rect 3833 3253 3847 3267
rect 3873 3253 3887 3267
rect 3993 3253 4007 3267
rect 4033 3253 4047 3267
rect 4113 3253 4127 3267
rect 4173 3253 4187 3267
rect 4213 3253 4227 3267
rect 4293 3253 4307 3267
rect 4673 3253 4687 3267
rect 4713 3253 4727 3267
rect 293 3233 307 3247
rect 333 3233 347 3247
rect 393 3233 407 3247
rect 473 3233 487 3247
rect 513 3233 527 3247
rect 573 3233 587 3247
rect 613 3233 627 3247
rect 693 3233 707 3247
rect 753 3233 767 3247
rect 813 3233 827 3247
rect 953 3233 967 3247
rect 1013 3233 1027 3247
rect 1153 3233 1167 3247
rect 1213 3233 1227 3247
rect 1513 3233 1527 3247
rect 1553 3233 1567 3247
rect 1613 3233 1627 3247
rect 1653 3233 1667 3247
rect 1713 3233 1727 3247
rect 1753 3233 1767 3247
rect 1813 3233 1827 3247
rect 1873 3233 1887 3247
rect 1913 3233 1927 3247
rect 1973 3233 1987 3247
rect 2013 3233 2027 3247
rect 2313 3233 2327 3247
rect 2373 3233 2387 3247
rect 2453 3233 2467 3247
rect 2493 3233 2507 3247
rect 2513 3233 2527 3247
rect 2553 3233 2567 3247
rect 2633 3233 2647 3247
rect 2693 3233 2707 3247
rect 2733 3233 2747 3247
rect 2873 3233 2887 3247
rect 2913 3233 2927 3247
rect 2973 3233 2987 3247
rect 3053 3233 3067 3247
rect 3153 3233 3167 3247
rect 3193 3233 3207 3247
rect 3253 3233 3267 3247
rect 3293 3233 3307 3247
rect 3333 3233 3347 3247
rect 3373 3233 3387 3247
rect 3533 3233 3547 3247
rect 3733 3233 3747 3247
rect 3773 3233 3787 3247
rect 3853 3233 3867 3247
rect 3913 3233 3927 3247
rect 3953 3233 3967 3247
rect 4013 3233 4027 3247
rect 4193 3233 4207 3247
rect 4353 3233 4367 3247
rect 4393 3233 4407 3247
rect 4473 3233 4487 3247
rect 4513 3233 4527 3247
rect 4573 3233 4587 3247
rect 4613 3233 4627 3247
rect 4693 3233 4707 3247
rect 4733 3233 4747 3247
rect 93 3213 107 3227
rect 133 3213 147 3227
rect 213 3213 227 3227
rect 273 3213 287 3227
rect 313 3213 327 3227
rect 353 3213 367 3227
rect 453 3213 467 3227
rect 493 3213 507 3227
rect 553 3213 567 3227
rect 593 3213 607 3227
rect 1273 3213 1287 3227
rect 1353 3213 1367 3227
rect 1393 3213 1407 3227
rect 1493 3213 1507 3227
rect 1533 3213 1547 3227
rect 1633 3213 1647 3227
rect 1673 3213 1687 3227
rect 1733 3213 1747 3227
rect 1773 3213 1787 3227
rect 1893 3213 1907 3227
rect 1933 3213 1947 3227
rect 1993 3213 2007 3227
rect 2033 3213 2047 3227
rect 2073 3213 2087 3227
rect 2153 3213 2167 3227
rect 2193 3213 2207 3227
rect 2573 3213 2587 3227
rect 2713 3213 2727 3227
rect 2753 3213 2767 3227
rect 2773 3213 2787 3227
rect 2813 3213 2827 3227
rect 2853 3213 2867 3227
rect 2893 3213 2907 3227
rect 3133 3213 3147 3227
rect 3353 3213 3367 3227
rect 3393 3213 3407 3227
rect 3433 3213 3447 3227
rect 3493 3213 3507 3227
rect 3613 3213 3627 3227
rect 3673 3213 3687 3227
rect 3713 3213 3727 3227
rect 3753 3213 3767 3227
rect 3793 3213 3807 3227
rect 3893 3213 3907 3227
rect 3933 3213 3947 3227
rect 4093 3213 4107 3227
rect 4153 3213 4167 3227
rect 4253 3213 4267 3227
rect 4313 3213 4327 3227
rect 4413 3213 4427 3227
rect 4453 3213 4467 3227
rect 4493 3213 4507 3227
rect 4553 3213 4567 3227
rect 4593 3213 4607 3227
rect 733 3193 747 3207
rect 1233 3193 1247 3207
rect 1833 3193 1847 3207
rect 2333 3193 2347 3207
rect 2393 3193 2407 3207
rect 2533 3193 2547 3207
rect 2653 3193 2667 3207
rect 2793 3193 2807 3207
rect 3173 3193 3187 3207
rect 4373 3193 4387 3207
rect 913 3053 927 3067
rect 1013 3053 1027 3067
rect 1253 3053 1267 3067
rect 1613 3053 1627 3067
rect 2213 3053 2227 3067
rect 2293 3053 2307 3067
rect 2473 3053 2487 3067
rect 2753 3053 2767 3067
rect 4173 3053 4187 3067
rect 4373 3053 4387 3067
rect 4553 3053 4567 3067
rect 93 3033 107 3047
rect 133 3033 147 3047
rect 213 3033 227 3047
rect 293 3033 307 3047
rect 333 3033 347 3047
rect 453 3033 467 3047
rect 533 3033 547 3047
rect 573 3033 587 3047
rect 753 3033 767 3047
rect 793 3033 807 3047
rect 873 3033 887 3047
rect 993 3033 1007 3047
rect 1033 3033 1047 3047
rect 1133 3033 1147 3047
rect 1173 3033 1187 3047
rect 1293 3033 1307 3047
rect 1413 3033 1427 3047
rect 1453 3033 1467 3047
rect 1533 3033 1547 3047
rect 1593 3033 1607 3047
rect 1633 3033 1647 3047
rect 1733 3033 1747 3047
rect 1773 3033 1787 3047
rect 1873 3033 1887 3047
rect 1913 3033 1927 3047
rect 1953 3033 1967 3047
rect 2033 3033 2047 3047
rect 2073 3033 2087 3047
rect 2193 3033 2207 3047
rect 2233 3033 2247 3047
rect 2433 3033 2447 3047
rect 2653 3033 2667 3047
rect 2693 3033 2707 3047
rect 2733 3033 2747 3047
rect 2773 3033 2787 3047
rect 2953 3033 2967 3047
rect 2993 3033 3007 3047
rect 3033 3033 3047 3047
rect 3153 3033 3167 3047
rect 3193 3033 3207 3047
rect 3273 3033 3287 3047
rect 3313 3033 3327 3047
rect 3373 3033 3387 3047
rect 3433 3033 3447 3047
rect 3473 3033 3487 3047
rect 3513 3033 3527 3047
rect 3553 3033 3567 3047
rect 3653 3033 3667 3047
rect 3693 3033 3707 3047
rect 3773 3033 3787 3047
rect 3813 3033 3827 3047
rect 3833 3033 3847 3047
rect 3873 3033 3887 3047
rect 4033 3033 4047 3047
rect 4073 3033 4087 3047
rect 4133 3033 4147 3047
rect 4333 3033 4347 3047
rect 4613 3033 4627 3047
rect 4653 3033 4667 3047
rect 4673 3033 4687 3047
rect 4713 3033 4727 3047
rect 273 3013 287 3027
rect 313 3013 327 3027
rect 393 3013 407 3027
rect 933 3013 947 3027
rect 1093 3013 1107 3027
rect 1153 3013 1167 3027
rect 1193 3013 1207 3027
rect 1233 3013 1247 3027
rect 1273 3013 1287 3027
rect 1693 3013 1707 3027
rect 1753 3013 1767 3027
rect 1793 3013 1807 3027
rect 1853 3013 1867 3027
rect 1893 3013 1907 3027
rect 2273 3013 2287 3027
rect 2353 3013 2367 3027
rect 2393 3013 2407 3027
rect 2453 3013 2467 3027
rect 2493 3013 2507 3027
rect 2553 3013 2567 3027
rect 2593 3013 2607 3027
rect 2633 3013 2647 3027
rect 2673 3013 2687 3027
rect 2813 3013 2827 3027
rect 2893 3013 2907 3027
rect 2973 3013 2987 3027
rect 3013 3013 3027 3027
rect 3093 3013 3107 3027
rect 3173 3013 3187 3027
rect 3213 3013 3227 3027
rect 3253 3013 3267 3027
rect 3593 3013 3607 3027
rect 3673 3013 3687 3027
rect 3713 3013 3727 3027
rect 3853 3013 3867 3027
rect 3893 3013 3907 3027
rect 3933 3013 3947 3027
rect 3973 3013 3987 3027
rect 4153 3013 4167 3027
rect 4193 3013 4207 3027
rect 4213 3013 4227 3027
rect 4253 3013 4267 3027
rect 4353 3013 4367 3027
rect 4393 3013 4407 3027
rect 4453 3013 4467 3027
rect 4493 3013 4507 3027
rect 4533 3013 4547 3027
rect 4593 3013 4607 3027
rect 4633 3013 4647 3027
rect 4693 3013 4707 3027
rect 4733 3013 4747 3027
rect 373 2993 387 3007
rect 413 2993 427 3007
rect 1073 2993 1087 3007
rect 1113 2993 1127 3007
rect 1673 2993 1687 3007
rect 1713 2993 1727 3007
rect 2333 2993 2347 3007
rect 2373 2993 2387 3007
rect 2533 2993 2547 3007
rect 2573 2993 2587 3007
rect 2793 2993 2807 3007
rect 2833 2993 2847 3007
rect 2873 2993 2887 3007
rect 2913 2993 2927 3007
rect 3073 2993 3087 3007
rect 3113 2993 3127 3007
rect 3353 2993 3367 3007
rect 3573 2993 3587 3007
rect 3613 2993 3627 3007
rect 3953 2993 3967 3007
rect 3993 2993 4007 3007
rect 4233 2993 4247 3007
rect 4273 2993 4287 3007
rect 4433 2993 4447 3007
rect 4473 2993 4487 3007
rect 373 2773 387 2787
rect 413 2773 427 2787
rect 633 2773 647 2787
rect 673 2773 687 2787
rect 913 2773 927 2787
rect 953 2773 967 2787
rect 1053 2773 1067 2787
rect 1093 2773 1107 2787
rect 1513 2773 1527 2787
rect 1553 2773 1567 2787
rect 2073 2773 2087 2787
rect 2113 2773 2127 2787
rect 2773 2773 2787 2787
rect 2813 2773 2827 2787
rect 2853 2773 2867 2787
rect 2893 2773 2907 2787
rect 3133 2773 3147 2787
rect 3173 2773 3187 2787
rect 3333 2773 3347 2787
rect 3373 2773 3387 2787
rect 3413 2773 3427 2787
rect 3453 2773 3467 2787
rect 3713 2773 3727 2787
rect 3753 2773 3767 2787
rect 3893 2773 3907 2787
rect 3933 2773 3947 2787
rect 4173 2773 4187 2787
rect 4213 2773 4227 2787
rect 4393 2773 4407 2787
rect 293 2753 307 2767
rect 333 2753 347 2767
rect 393 2753 407 2767
rect 473 2753 487 2767
rect 513 2753 527 2767
rect 653 2753 667 2767
rect 733 2753 747 2767
rect 773 2753 787 2767
rect 933 2753 947 2767
rect 993 2753 1007 2767
rect 1073 2753 1087 2767
rect 1533 2753 1547 2767
rect 1613 2753 1627 2767
rect 1653 2753 1667 2767
rect 1713 2753 1727 2767
rect 1753 2753 1767 2767
rect 1913 2753 1927 2767
rect 1953 2753 1967 2767
rect 2093 2753 2107 2767
rect 2133 2753 2147 2767
rect 2493 2753 2507 2767
rect 2533 2753 2547 2767
rect 2593 2753 2607 2767
rect 2633 2753 2647 2767
rect 2693 2753 2707 2767
rect 2733 2753 2747 2767
rect 2793 2753 2807 2767
rect 2873 2753 2887 2767
rect 2953 2753 2967 2767
rect 2993 2753 3007 2767
rect 3053 2753 3067 2767
rect 3093 2753 3107 2767
rect 3153 2753 3167 2767
rect 3233 2753 3247 2767
rect 3273 2753 3287 2767
rect 3353 2753 3367 2767
rect 3393 2753 3407 2767
rect 3433 2753 3447 2767
rect 3513 2753 3527 2767
rect 3553 2753 3567 2767
rect 3613 2753 3627 2767
rect 3653 2753 3667 2767
rect 3733 2753 3747 2767
rect 3793 2753 3807 2767
rect 3833 2753 3847 2767
rect 3873 2753 3887 2767
rect 3913 2753 3927 2767
rect 3993 2753 4007 2767
rect 4073 2753 4087 2767
rect 4113 2753 4127 2767
rect 4153 2753 4167 2767
rect 4193 2753 4207 2767
rect 4273 2753 4287 2767
rect 4313 2753 4327 2767
rect 4473 2753 4487 2767
rect 4513 2753 4527 2767
rect 4593 2753 4607 2767
rect 4633 2753 4647 2767
rect 4673 2753 4687 2767
rect 93 2733 107 2747
rect 133 2733 147 2747
rect 213 2733 227 2747
rect 273 2733 287 2747
rect 313 2733 327 2747
rect 353 2733 367 2747
rect 493 2733 507 2747
rect 533 2733 547 2747
rect 573 2733 587 2747
rect 613 2733 627 2747
rect 753 2733 767 2747
rect 793 2733 807 2747
rect 833 2733 847 2747
rect 873 2733 887 2747
rect 1113 2733 1127 2747
rect 1153 2733 1167 2747
rect 1213 2733 1227 2747
rect 1253 2733 1267 2747
rect 1353 2733 1367 2747
rect 1393 2733 1407 2747
rect 1473 2733 1487 2747
rect 1633 2733 1647 2747
rect 1673 2733 1687 2747
rect 1733 2733 1747 2747
rect 1773 2733 1787 2747
rect 1813 2733 1827 2747
rect 1853 2733 1867 2747
rect 1893 2733 1907 2747
rect 1993 2733 2007 2747
rect 2033 2733 2047 2747
rect 2153 2733 2167 2747
rect 2193 2733 2207 2747
rect 2313 2733 2327 2747
rect 2353 2733 2367 2747
rect 2433 2733 2447 2747
rect 2513 2733 2527 2747
rect 2553 2733 2567 2747
rect 2613 2733 2627 2747
rect 2653 2733 2667 2747
rect 2673 2733 2687 2747
rect 2713 2733 2727 2747
rect 2933 2733 2947 2747
rect 2973 2733 2987 2747
rect 3033 2733 3047 2747
rect 3073 2733 3087 2747
rect 3253 2733 3267 2747
rect 3293 2733 3307 2747
rect 3533 2733 3547 2747
rect 3573 2733 3587 2747
rect 3593 2733 3607 2747
rect 3633 2733 3647 2747
rect 3813 2733 3827 2747
rect 3853 2733 3867 2747
rect 4053 2733 4067 2747
rect 4093 2733 4107 2747
rect 4133 2733 4147 2747
rect 4253 2733 4267 2747
rect 4293 2733 4307 2747
rect 4353 2733 4367 2747
rect 4413 2733 4427 2747
rect 4453 2733 4467 2747
rect 4493 2733 4507 2747
rect 4533 2733 4547 2747
rect 4693 2733 4707 2747
rect 853 2713 867 2727
rect 973 2713 987 2727
rect 1133 2713 1147 2727
rect 1833 2713 1847 2727
rect 1933 2713 1947 2727
rect 3973 2713 3987 2727
rect 4573 2713 4587 2727
rect 4653 2713 4667 2727
rect 813 2573 827 2587
rect 1113 2573 1127 2587
rect 1273 2573 1287 2587
rect 2513 2573 2527 2587
rect 2673 2573 2687 2587
rect 3393 2573 3407 2587
rect 3713 2573 3727 2587
rect 4553 2573 4567 2587
rect 93 2553 107 2567
rect 133 2553 147 2567
rect 213 2553 227 2567
rect 293 2553 307 2567
rect 333 2553 347 2567
rect 353 2553 367 2567
rect 393 2553 407 2567
rect 553 2553 567 2567
rect 593 2553 607 2567
rect 613 2553 627 2567
rect 653 2553 667 2567
rect 733 2553 747 2567
rect 773 2553 787 2567
rect 793 2553 807 2567
rect 833 2553 847 2567
rect 953 2553 967 2567
rect 993 2553 1007 2567
rect 1073 2553 1087 2567
rect 1173 2553 1187 2567
rect 1213 2553 1227 2567
rect 1433 2553 1447 2567
rect 1513 2553 1527 2567
rect 1553 2553 1567 2567
rect 1653 2553 1667 2567
rect 1693 2553 1707 2567
rect 1773 2553 1787 2567
rect 1853 2553 1867 2567
rect 1893 2553 1907 2567
rect 2273 2553 2287 2567
rect 2313 2553 2327 2567
rect 2393 2553 2407 2567
rect 2613 2553 2627 2567
rect 2653 2553 2667 2567
rect 2853 2553 2867 2567
rect 2893 2553 2907 2567
rect 2913 2553 2927 2567
rect 2973 2553 2987 2567
rect 3013 2553 3027 2567
rect 3053 2553 3067 2567
rect 3193 2553 3207 2567
rect 3253 2553 3267 2567
rect 3533 2553 3547 2567
rect 3593 2553 3607 2567
rect 3633 2553 3647 2567
rect 3673 2553 3687 2567
rect 3793 2553 3807 2567
rect 3853 2553 3867 2567
rect 3893 2553 3907 2567
rect 3933 2553 3947 2567
rect 3973 2553 3987 2567
rect 4153 2553 4167 2567
rect 4193 2553 4207 2567
rect 4593 2553 4607 2567
rect 273 2533 287 2547
rect 313 2533 327 2547
rect 453 2533 467 2547
rect 533 2533 547 2547
rect 573 2533 587 2547
rect 713 2533 727 2547
rect 753 2533 767 2547
rect 1133 2533 1147 2547
rect 1193 2533 1207 2547
rect 1233 2533 1247 2547
rect 1293 2533 1307 2547
rect 1353 2533 1367 2547
rect 1673 2533 1687 2547
rect 1713 2533 1727 2547
rect 2013 2533 2027 2547
rect 2153 2533 2167 2547
rect 2473 2533 2487 2547
rect 2533 2533 2547 2547
rect 2593 2533 2607 2547
rect 2633 2533 2647 2547
rect 2693 2533 2707 2547
rect 2773 2533 2787 2547
rect 2833 2533 2847 2547
rect 2873 2533 2887 2547
rect 3033 2533 3047 2547
rect 3073 2533 3087 2547
rect 3153 2533 3167 2547
rect 3333 2533 3347 2547
rect 3373 2533 3387 2547
rect 3413 2533 3427 2547
rect 3473 2533 3487 2547
rect 3733 2533 3747 2547
rect 3913 2533 3927 2547
rect 3953 2533 3967 2547
rect 4033 2533 4047 2547
rect 4113 2533 4127 2547
rect 4173 2533 4187 2547
rect 4213 2533 4227 2547
rect 4273 2533 4287 2547
rect 4373 2533 4387 2547
rect 4413 2533 4427 2547
rect 4473 2533 4487 2547
rect 4513 2533 4527 2547
rect 4533 2533 4547 2547
rect 4573 2533 4587 2547
rect 4673 2533 4687 2547
rect 4713 2533 4727 2547
rect 433 2513 447 2527
rect 473 2513 487 2527
rect 1333 2513 1347 2527
rect 1373 2513 1387 2527
rect 2453 2513 2467 2527
rect 2493 2513 2507 2527
rect 2753 2513 2767 2527
rect 2793 2513 2807 2527
rect 2953 2513 2967 2527
rect 3133 2513 3147 2527
rect 3173 2513 3187 2527
rect 3233 2513 3247 2527
rect 3313 2513 3327 2527
rect 3353 2513 3367 2527
rect 3453 2513 3467 2527
rect 3493 2513 3507 2527
rect 3573 2513 3587 2527
rect 3813 2513 3827 2527
rect 4013 2513 4027 2527
rect 4053 2513 4067 2527
rect 4093 2513 4107 2527
rect 4133 2513 4147 2527
rect 4253 2513 4267 2527
rect 4293 2513 4307 2527
rect 4353 2513 4367 2527
rect 4393 2513 4407 2527
rect 4453 2513 4467 2527
rect 4493 2513 4507 2527
rect 4653 2513 4667 2527
rect 4693 2513 4707 2527
rect 553 2293 567 2307
rect 593 2293 607 2307
rect 2553 2293 2567 2307
rect 2593 2293 2607 2307
rect 2613 2293 2627 2307
rect 2653 2293 2667 2307
rect 2693 2293 2707 2307
rect 2733 2293 2747 2307
rect 3313 2293 3327 2307
rect 3353 2293 3367 2307
rect 3393 2293 3407 2307
rect 3433 2293 3447 2307
rect 3493 2293 3507 2307
rect 3533 2293 3547 2307
rect 4013 2293 4027 2307
rect 4193 2293 4207 2307
rect 4233 2293 4247 2307
rect 273 2273 287 2287
rect 313 2273 327 2287
rect 373 2273 387 2287
rect 413 2273 427 2287
rect 573 2273 587 2287
rect 653 2273 667 2287
rect 813 2273 827 2287
rect 853 2273 867 2287
rect 1053 2273 1067 2287
rect 1353 2273 1367 2287
rect 1393 2273 1407 2287
rect 1793 2273 1807 2287
rect 1833 2273 1847 2287
rect 1853 2273 1867 2287
rect 2013 2273 2027 2287
rect 2153 2273 2167 2287
rect 2213 2273 2227 2287
rect 2253 2273 2267 2287
rect 2573 2273 2587 2287
rect 2633 2273 2647 2287
rect 2713 2273 2727 2287
rect 2793 2273 2807 2287
rect 2833 2273 2847 2287
rect 2893 2273 2907 2287
rect 2933 2273 2947 2287
rect 3233 2273 3247 2287
rect 3273 2273 3287 2287
rect 3333 2273 3347 2287
rect 3413 2273 3427 2287
rect 3513 2273 3527 2287
rect 3593 2273 3607 2287
rect 3653 2273 3667 2287
rect 3693 2273 3707 2287
rect 3753 2273 3767 2287
rect 3793 2273 3807 2287
rect 3913 2273 3927 2287
rect 4093 2273 4107 2287
rect 4133 2273 4147 2287
rect 4213 2273 4227 2287
rect 4253 2273 4267 2287
rect 4273 2273 4287 2287
rect 4313 2273 4327 2287
rect 4393 2273 4407 2287
rect 4433 2273 4447 2287
rect 4493 2273 4507 2287
rect 4533 2273 4547 2287
rect 4593 2273 4607 2287
rect 4633 2273 4647 2287
rect 4673 2273 4687 2287
rect 4713 2273 4727 2287
rect 93 2253 107 2267
rect 133 2253 147 2267
rect 213 2253 227 2267
rect 253 2253 267 2267
rect 293 2253 307 2267
rect 353 2253 367 2267
rect 393 2253 407 2267
rect 433 2253 447 2267
rect 473 2253 487 2267
rect 513 2253 527 2267
rect 693 2253 707 2267
rect 733 2253 747 2267
rect 793 2253 807 2267
rect 873 2253 887 2267
rect 913 2253 927 2267
rect 953 2253 967 2267
rect 993 2253 1007 2267
rect 1113 2253 1127 2267
rect 1193 2253 1207 2267
rect 1233 2253 1247 2267
rect 1333 2253 1347 2267
rect 1373 2253 1387 2267
rect 1453 2253 1467 2267
rect 1533 2253 1547 2267
rect 1573 2253 1587 2267
rect 1693 2253 1707 2267
rect 1733 2253 1747 2267
rect 1773 2253 1787 2267
rect 1873 2253 1887 2267
rect 1933 2253 1947 2267
rect 1973 2253 1987 2267
rect 2193 2253 2207 2267
rect 2233 2253 2247 2267
rect 2373 2253 2387 2267
rect 2413 2253 2427 2267
rect 2493 2253 2507 2267
rect 2813 2253 2827 2267
rect 2853 2253 2867 2267
rect 2913 2253 2927 2267
rect 2953 2253 2967 2267
rect 3053 2253 3067 2267
rect 3093 2253 3107 2267
rect 3173 2253 3187 2267
rect 3213 2253 3227 2267
rect 3253 2253 3267 2267
rect 3573 2253 3587 2267
rect 3633 2253 3647 2267
rect 3733 2253 3747 2267
rect 3773 2253 3787 2267
rect 3853 2253 3867 2267
rect 3893 2253 3907 2267
rect 3933 2253 3947 2267
rect 3973 2253 3987 2267
rect 4033 2253 4047 2267
rect 4113 2253 4127 2267
rect 4153 2253 4167 2267
rect 4333 2253 4347 2267
rect 4413 2253 4427 2267
rect 4453 2253 4467 2267
rect 4473 2253 4487 2267
rect 4513 2253 4527 2267
rect 4613 2253 4627 2267
rect 4653 2253 4667 2267
rect 4733 2253 4747 2267
rect 673 2233 687 2247
rect 713 2233 727 2247
rect 833 2233 847 2247
rect 893 2233 907 2247
rect 973 2233 987 2247
rect 1033 2233 1047 2247
rect 1713 2233 1727 2247
rect 1813 2233 1827 2247
rect 1953 2233 1967 2247
rect 3713 2233 3727 2247
rect 4293 2233 4307 2247
rect 4693 2233 4707 2247
rect 913 2093 927 2107
rect 1033 2093 1047 2107
rect 1293 2093 1307 2107
rect 1653 2093 1667 2107
rect 2053 2093 2067 2107
rect 3593 2093 3607 2107
rect 4373 2093 4387 2107
rect 4513 2093 4527 2107
rect 333 2073 347 2087
rect 373 2073 387 2087
rect 393 2073 407 2087
rect 433 2073 447 2087
rect 473 2073 487 2087
rect 593 2073 607 2087
rect 633 2073 647 2087
rect 713 2073 727 2087
rect 893 2073 907 2087
rect 1013 2073 1027 2087
rect 1053 2073 1067 2087
rect 1093 2073 1107 2087
rect 1133 2073 1147 2087
rect 1273 2073 1287 2087
rect 1313 2073 1327 2087
rect 1373 2073 1387 2087
rect 1453 2073 1467 2087
rect 1493 2073 1507 2087
rect 1613 2073 1627 2087
rect 1713 2073 1727 2087
rect 1753 2073 1767 2087
rect 1793 2073 1807 2087
rect 1873 2073 1887 2087
rect 1913 2073 1927 2087
rect 2153 2073 2167 2087
rect 2193 2073 2207 2087
rect 2353 2073 2367 2087
rect 2393 2073 2407 2087
rect 2613 2073 2627 2087
rect 2653 2073 2667 2087
rect 2713 2073 2727 2087
rect 2753 2073 2767 2087
rect 2853 2073 2867 2087
rect 2893 2073 2907 2087
rect 2973 2073 2987 2087
rect 3013 2073 3027 2087
rect 3073 2073 3087 2087
rect 3153 2073 3167 2087
rect 3193 2073 3207 2087
rect 3253 2073 3267 2087
rect 3293 2073 3307 2087
rect 3433 2073 3447 2087
rect 3473 2073 3487 2087
rect 3833 2073 3847 2087
rect 3873 2073 3887 2087
rect 3913 2073 3927 2087
rect 3953 2073 3967 2087
rect 4253 2073 4267 2087
rect 4313 2073 4327 2087
rect 4413 2073 4427 2087
rect 4473 2073 4487 2087
rect 33 2053 47 2067
rect 173 2053 187 2067
rect 253 2053 267 2067
rect 313 2053 327 2067
rect 353 2053 367 2067
rect 413 2053 427 2067
rect 453 2053 467 2067
rect 793 2053 807 2067
rect 853 2053 867 2067
rect 953 2053 967 2067
rect 1113 2053 1127 2067
rect 1153 2053 1167 2067
rect 1213 2053 1227 2067
rect 1633 2053 1647 2067
rect 1673 2053 1687 2067
rect 2033 2053 2047 2067
rect 2113 2053 2127 2067
rect 2253 2053 2267 2067
rect 2333 2053 2347 2067
rect 2373 2053 2387 2067
rect 2453 2053 2467 2067
rect 2533 2053 2547 2067
rect 2593 2053 2607 2067
rect 2633 2053 2647 2067
rect 2693 2053 2707 2067
rect 2733 2053 2747 2067
rect 3133 2053 3147 2067
rect 3173 2053 3187 2067
rect 3233 2053 3247 2067
rect 3273 2053 3287 2067
rect 3333 2053 3347 2067
rect 3413 2053 3427 2067
rect 3453 2053 3467 2067
rect 3493 2053 3507 2067
rect 3533 2053 3547 2067
rect 3613 2053 3627 2067
rect 3653 2053 3667 2067
rect 3693 2053 3707 2067
rect 3773 2053 3787 2067
rect 3933 2053 3947 2067
rect 3973 2053 3987 2067
rect 4053 2053 4067 2067
rect 4133 2053 4147 2067
rect 4213 2053 4227 2067
rect 4353 2053 4367 2067
rect 4393 2053 4407 2067
rect 4493 2053 4507 2067
rect 4533 2053 4547 2067
rect 4553 2053 4567 2067
rect 4593 2053 4607 2067
rect 4653 2053 4667 2067
rect 4693 2053 4707 2067
rect 233 2033 247 2047
rect 273 2033 287 2047
rect 773 2033 787 2047
rect 813 2033 827 2047
rect 933 2033 947 2047
rect 973 2033 987 2047
rect 1193 2033 1207 2047
rect 1233 2033 1247 2047
rect 2093 2033 2107 2047
rect 2133 2033 2147 2047
rect 2233 2033 2247 2047
rect 2273 2033 2287 2047
rect 2433 2033 2447 2047
rect 2473 2033 2487 2047
rect 2513 2033 2527 2047
rect 2553 2033 2567 2047
rect 3053 2033 3067 2047
rect 3313 2033 3327 2047
rect 3353 2033 3367 2047
rect 3513 2033 3527 2047
rect 3553 2033 3567 2047
rect 3673 2033 3687 2047
rect 3713 2033 3727 2047
rect 3753 2033 3767 2047
rect 3793 2033 3807 2047
rect 4033 2033 4047 2047
rect 4073 2033 4087 2047
rect 4113 2033 4127 2047
rect 4153 2033 4167 2047
rect 4193 2033 4207 2047
rect 4233 2033 4247 2047
rect 4293 2033 4307 2047
rect 4573 2033 4587 2047
rect 4613 2033 4627 2047
rect 4673 2033 4687 2047
rect 4713 2033 4727 2047
rect 873 1813 887 1827
rect 913 1813 927 1827
rect 1193 1813 1207 1827
rect 1233 1813 1247 1827
rect 3073 1813 3087 1827
rect 3113 1813 3127 1827
rect 3413 1813 3427 1827
rect 3913 1813 3927 1827
rect 4213 1813 4227 1827
rect 4253 1813 4267 1827
rect 4333 1813 4347 1827
rect 273 1793 287 1807
rect 313 1793 327 1807
rect 373 1793 387 1807
rect 413 1793 427 1807
rect 473 1793 487 1807
rect 513 1793 527 1807
rect 573 1793 587 1807
rect 613 1793 627 1807
rect 673 1793 687 1807
rect 733 1793 747 1807
rect 853 1793 867 1807
rect 893 1793 907 1807
rect 1213 1793 1227 1807
rect 1293 1793 1307 1807
rect 1333 1793 1347 1807
rect 1393 1793 1407 1807
rect 1533 1793 1547 1807
rect 1853 1793 1867 1807
rect 1893 1793 1907 1807
rect 2033 1793 2047 1807
rect 2073 1793 2087 1807
rect 2173 1793 2187 1807
rect 2213 1793 2227 1807
rect 3033 1793 3047 1807
rect 3093 1793 3107 1807
rect 3173 1793 3187 1807
rect 3193 1793 3207 1807
rect 3233 1793 3247 1807
rect 3473 1793 3487 1807
rect 3573 1793 3587 1807
rect 3613 1793 3627 1807
rect 3693 1793 3707 1807
rect 4013 1793 4027 1807
rect 4053 1793 4067 1807
rect 4113 1793 4127 1807
rect 4153 1793 4167 1807
rect 4233 1793 4247 1807
rect 4413 1793 4427 1807
rect 4453 1793 4467 1807
rect 4533 1793 4547 1807
rect 4593 1793 4607 1807
rect 4633 1793 4647 1807
rect 4693 1793 4707 1807
rect 93 1773 107 1787
rect 133 1773 147 1787
rect 213 1773 227 1787
rect 253 1773 267 1787
rect 293 1773 307 1787
rect 393 1773 407 1787
rect 433 1773 447 1787
rect 493 1773 507 1787
rect 533 1773 547 1787
rect 593 1773 607 1787
rect 633 1773 647 1787
rect 793 1773 807 1787
rect 833 1773 847 1787
rect 1033 1773 1047 1787
rect 1073 1773 1087 1787
rect 1153 1773 1167 1787
rect 1313 1773 1327 1787
rect 1353 1773 1367 1787
rect 1653 1773 1667 1787
rect 1693 1773 1707 1787
rect 1773 1773 1787 1787
rect 1833 1773 1847 1787
rect 1913 1773 1927 1787
rect 1953 1773 1967 1787
rect 2013 1773 2027 1787
rect 2113 1773 2127 1787
rect 2153 1773 2167 1787
rect 2233 1773 2247 1787
rect 2293 1773 2307 1787
rect 2373 1773 2387 1787
rect 2413 1773 2427 1787
rect 2593 1773 2607 1787
rect 2633 1773 2647 1787
rect 2713 1773 2727 1787
rect 2833 1773 2847 1787
rect 2873 1773 2887 1787
rect 2953 1773 2967 1787
rect 3013 1773 3027 1787
rect 3153 1773 3167 1787
rect 3253 1773 3267 1787
rect 3293 1773 3307 1787
rect 3333 1773 3347 1787
rect 3393 1773 3407 1787
rect 3453 1773 3467 1787
rect 3493 1773 3507 1787
rect 3553 1773 3567 1787
rect 3593 1773 3607 1787
rect 3633 1773 3647 1787
rect 3673 1773 3687 1787
rect 3733 1773 3747 1787
rect 3773 1773 3787 1787
rect 3793 1773 3807 1787
rect 3833 1773 3847 1787
rect 3873 1773 3887 1787
rect 3933 1773 3947 1787
rect 3993 1773 4007 1787
rect 4033 1773 4047 1787
rect 4073 1773 4087 1787
rect 4093 1773 4107 1787
rect 4133 1773 4147 1787
rect 4173 1773 4187 1787
rect 4293 1773 4307 1787
rect 4353 1773 4367 1787
rect 4393 1773 4407 1787
rect 4433 1773 4447 1787
rect 4473 1773 4487 1787
rect 4573 1773 4587 1787
rect 4613 1773 4627 1787
rect 653 1753 667 1767
rect 713 1753 727 1767
rect 813 1753 827 1767
rect 1873 1753 1887 1767
rect 1933 1753 1947 1767
rect 2053 1753 2067 1767
rect 2133 1753 2147 1767
rect 2193 1753 2207 1767
rect 3213 1753 3227 1767
rect 3313 1753 3327 1767
rect 3753 1753 3767 1767
rect 4553 1753 4567 1767
rect 4673 1753 4687 1767
rect 253 1613 267 1627
rect 1813 1613 1827 1627
rect 1873 1613 1887 1627
rect 2213 1613 2227 1627
rect 3713 1613 3727 1627
rect 3893 1613 3907 1627
rect 4173 1613 4187 1627
rect 4353 1613 4367 1627
rect 4433 1613 4447 1627
rect 233 1593 247 1607
rect 273 1593 287 1607
rect 313 1593 327 1607
rect 353 1593 367 1607
rect 453 1593 467 1607
rect 493 1593 507 1607
rect 573 1593 587 1607
rect 693 1593 707 1607
rect 733 1593 747 1607
rect 813 1593 827 1607
rect 873 1593 887 1607
rect 953 1593 967 1607
rect 993 1593 1007 1607
rect 1213 1593 1227 1607
rect 1253 1593 1267 1607
rect 1293 1593 1307 1607
rect 1373 1593 1387 1607
rect 1413 1593 1427 1607
rect 1593 1593 1607 1607
rect 1633 1593 1647 1607
rect 1713 1593 1727 1607
rect 1773 1593 1787 1607
rect 1853 1593 1867 1607
rect 1893 1593 1907 1607
rect 2013 1593 2027 1607
rect 2053 1593 2067 1607
rect 2133 1593 2147 1607
rect 2193 1593 2207 1607
rect 2233 1593 2247 1607
rect 2333 1593 2347 1607
rect 2373 1593 2387 1607
rect 2453 1593 2467 1607
rect 2533 1593 2547 1607
rect 2573 1593 2587 1607
rect 2753 1593 2767 1607
rect 2793 1593 2807 1607
rect 2873 1593 2887 1607
rect 2933 1593 2947 1607
rect 3133 1593 3147 1607
rect 3173 1593 3187 1607
rect 3433 1593 3447 1607
rect 3473 1593 3487 1607
rect 3613 1593 3627 1607
rect 3653 1593 3667 1607
rect 3693 1593 3707 1607
rect 3933 1593 3947 1607
rect 3973 1593 3987 1607
rect 4013 1593 4027 1607
rect 4213 1593 4227 1607
rect 4253 1593 4267 1607
rect 4293 1593 4307 1607
rect 4413 1593 4427 1607
rect 4453 1593 4467 1607
rect 33 1573 47 1587
rect 173 1573 187 1587
rect 1133 1573 1147 1587
rect 1193 1573 1207 1587
rect 1233 1573 1247 1587
rect 1793 1573 1807 1587
rect 1833 1573 1847 1587
rect 2293 1573 2307 1587
rect 2353 1573 2367 1587
rect 2393 1573 2407 1587
rect 2913 1573 2927 1587
rect 2993 1573 3007 1587
rect 3093 1573 3107 1587
rect 3153 1573 3167 1587
rect 3193 1573 3207 1587
rect 3253 1573 3267 1587
rect 3353 1573 3367 1587
rect 3413 1573 3427 1587
rect 3453 1573 3467 1587
rect 3493 1573 3507 1587
rect 3533 1573 3547 1587
rect 3633 1573 3647 1587
rect 3673 1573 3687 1587
rect 3733 1573 3747 1587
rect 3773 1573 3787 1587
rect 3813 1573 3827 1587
rect 3873 1573 3887 1587
rect 3913 1573 3927 1587
rect 3993 1573 4007 1587
rect 4033 1573 4047 1587
rect 4113 1573 4127 1587
rect 4153 1573 4167 1587
rect 4193 1573 4207 1587
rect 4273 1573 4287 1587
rect 4313 1573 4327 1587
rect 4373 1573 4387 1587
rect 4513 1573 4527 1587
rect 4593 1573 4607 1587
rect 4673 1573 4687 1587
rect 1113 1553 1127 1567
rect 1153 1553 1167 1567
rect 2273 1553 2287 1567
rect 2313 1553 2327 1567
rect 2973 1553 2987 1567
rect 3013 1553 3027 1567
rect 3073 1553 3087 1567
rect 3113 1553 3127 1567
rect 3233 1553 3247 1567
rect 3273 1553 3287 1567
rect 3333 1553 3347 1567
rect 3373 1553 3387 1567
rect 3513 1553 3527 1567
rect 3553 1553 3567 1567
rect 3793 1553 3807 1567
rect 3833 1553 3847 1567
rect 4093 1553 4107 1567
rect 4133 1553 4147 1567
rect 4493 1553 4507 1567
rect 4533 1553 4547 1567
rect 4573 1553 4587 1567
rect 4613 1553 4627 1567
rect 4653 1553 4667 1567
rect 4693 1553 4707 1567
rect 493 1333 507 1347
rect 533 1333 547 1347
rect 853 1333 867 1347
rect 893 1333 907 1347
rect 1233 1333 1247 1347
rect 1273 1333 1287 1347
rect 1413 1333 1427 1347
rect 1453 1333 1467 1347
rect 1653 1333 1667 1347
rect 1693 1333 1707 1347
rect 2253 1333 2267 1347
rect 2293 1333 2307 1347
rect 3253 1333 3267 1347
rect 3413 1333 3427 1347
rect 3453 1333 3467 1347
rect 3713 1333 3727 1347
rect 3753 1333 3767 1347
rect 3793 1333 3807 1347
rect 3833 1333 3847 1347
rect 3893 1333 3907 1347
rect 4133 1333 4147 1347
rect 4173 1333 4187 1347
rect 4213 1333 4227 1347
rect 4253 1333 4267 1347
rect 4653 1333 4667 1347
rect 4693 1333 4707 1347
rect 513 1313 527 1327
rect 593 1313 607 1327
rect 633 1313 647 1327
rect 693 1313 707 1327
rect 733 1313 747 1327
rect 873 1313 887 1327
rect 953 1313 967 1327
rect 993 1313 1007 1327
rect 1053 1313 1067 1327
rect 1253 1313 1267 1327
rect 1313 1313 1327 1327
rect 1353 1313 1367 1327
rect 1433 1313 1447 1327
rect 1493 1313 1507 1327
rect 1533 1313 1547 1327
rect 1673 1313 1687 1327
rect 1753 1313 1767 1327
rect 1793 1313 1807 1327
rect 2093 1313 2107 1327
rect 2153 1313 2167 1327
rect 2193 1313 2207 1327
rect 2273 1313 2287 1327
rect 2413 1313 2427 1327
rect 2893 1313 2907 1327
rect 2933 1313 2947 1327
rect 2973 1313 2987 1327
rect 3033 1313 3047 1327
rect 3073 1313 3087 1327
rect 3133 1313 3147 1327
rect 3173 1313 3187 1327
rect 3393 1313 3407 1327
rect 3433 1313 3447 1327
rect 3513 1313 3527 1327
rect 3553 1313 3567 1327
rect 3613 1313 3627 1327
rect 3653 1313 3667 1327
rect 3733 1313 3747 1327
rect 3813 1313 3827 1327
rect 3973 1313 3987 1327
rect 4013 1313 4027 1327
rect 4073 1313 4087 1327
rect 4153 1313 4167 1327
rect 4233 1313 4247 1327
rect 4373 1313 4387 1327
rect 4413 1313 4427 1327
rect 4473 1313 4487 1327
rect 4513 1313 4527 1327
rect 4593 1313 4607 1327
rect 4633 1313 4647 1327
rect 4673 1313 4687 1327
rect 33 1293 47 1307
rect 113 1293 127 1307
rect 153 1293 167 1307
rect 333 1293 347 1307
rect 373 1293 387 1307
rect 453 1293 467 1307
rect 613 1293 627 1307
rect 653 1293 667 1307
rect 713 1293 727 1307
rect 753 1293 767 1307
rect 793 1293 807 1307
rect 833 1293 847 1307
rect 973 1293 987 1307
rect 1013 1293 1027 1307
rect 1113 1293 1127 1307
rect 1153 1293 1167 1307
rect 1333 1293 1347 1307
rect 1373 1293 1387 1307
rect 1513 1293 1527 1307
rect 1553 1293 1567 1307
rect 1573 1293 1587 1307
rect 1613 1293 1627 1307
rect 1773 1293 1787 1307
rect 1813 1293 1827 1307
rect 1853 1293 1867 1307
rect 1933 1293 1947 1307
rect 1973 1293 1987 1307
rect 2133 1293 2147 1307
rect 2173 1293 2187 1307
rect 2333 1293 2347 1307
rect 2373 1293 2387 1307
rect 2453 1293 2467 1307
rect 2493 1293 2507 1307
rect 2553 1293 2567 1307
rect 2633 1293 2647 1307
rect 2673 1293 2687 1307
rect 2773 1293 2787 1307
rect 2813 1293 2827 1307
rect 2873 1293 2887 1307
rect 2913 1293 2927 1307
rect 2953 1293 2967 1307
rect 3013 1293 3027 1307
rect 3053 1293 3067 1307
rect 3113 1293 3127 1307
rect 3153 1293 3167 1307
rect 3213 1293 3227 1307
rect 3273 1293 3287 1307
rect 3333 1293 3347 1307
rect 3373 1293 3387 1307
rect 3533 1293 3547 1307
rect 3573 1293 3587 1307
rect 3593 1293 3607 1307
rect 3633 1293 3647 1307
rect 3853 1293 3867 1307
rect 3913 1293 3927 1307
rect 3993 1293 4007 1307
rect 4033 1293 4047 1307
rect 4293 1293 4307 1307
rect 4333 1293 4347 1307
rect 4393 1293 4407 1307
rect 4433 1293 4447 1307
rect 4453 1293 4467 1307
rect 4493 1293 4507 1307
rect 4573 1293 4587 1307
rect 1073 1273 1087 1287
rect 2073 1273 2087 1287
rect 2353 1273 2367 1287
rect 2433 1273 2447 1287
rect 2473 1273 2487 1287
rect 2793 1273 2807 1287
rect 3353 1273 3367 1287
rect 4053 1273 4067 1287
rect 4313 1273 4327 1287
rect 4613 1273 4627 1287
rect 13 1133 27 1147
rect 433 1133 447 1147
rect 553 1133 567 1147
rect 593 1133 607 1147
rect 873 1133 887 1147
rect 953 1133 967 1147
rect 1013 1133 1027 1147
rect 1053 1133 1067 1147
rect 1113 1133 1127 1147
rect 1213 1133 1227 1147
rect 1273 1133 1287 1147
rect 1633 1133 1647 1147
rect 1753 1133 1767 1147
rect 2093 1133 2107 1147
rect 2133 1133 2147 1147
rect 2213 1133 2227 1147
rect 2313 1133 2327 1147
rect 2573 1133 2587 1147
rect 2873 1133 2887 1147
rect 3213 1133 3227 1147
rect 3853 1133 3867 1147
rect 3973 1133 3987 1147
rect 4113 1133 4127 1147
rect 4193 1133 4207 1147
rect 4313 1133 4327 1147
rect 4573 1133 4587 1147
rect 4753 1133 4767 1147
rect 193 1113 207 1127
rect 233 1113 247 1127
rect 253 1113 267 1127
rect 293 1113 307 1127
rect 333 1113 347 1127
rect 393 1113 407 1127
rect 533 1113 547 1127
rect 573 1113 587 1127
rect 613 1113 627 1127
rect 673 1113 687 1127
rect 733 1113 747 1127
rect 773 1113 787 1127
rect 813 1113 827 1127
rect 853 1113 867 1127
rect 893 1113 907 1127
rect 1033 1113 1047 1127
rect 1073 1113 1087 1127
rect 1193 1113 1207 1127
rect 1233 1113 1247 1127
rect 1313 1113 1327 1127
rect 1433 1113 1447 1127
rect 1473 1113 1487 1127
rect 1553 1113 1567 1127
rect 1733 1113 1747 1127
rect 1773 1113 1787 1127
rect 1893 1113 1907 1127
rect 1933 1113 1947 1127
rect 2013 1113 2027 1127
rect 2113 1113 2127 1127
rect 2153 1113 2167 1127
rect 2193 1113 2207 1127
rect 2233 1113 2247 1127
rect 2353 1113 2367 1127
rect 2433 1113 2447 1127
rect 2473 1113 2487 1127
rect 2633 1113 2647 1127
rect 2673 1113 2687 1127
rect 2733 1113 2747 1127
rect 2773 1113 2787 1127
rect 2813 1113 2827 1127
rect 2853 1113 2867 1127
rect 2893 1113 2907 1127
rect 3013 1113 3027 1127
rect 3073 1113 3087 1127
rect 3113 1113 3127 1127
rect 3153 1113 3167 1127
rect 3233 1113 3247 1127
rect 3633 1113 3647 1127
rect 3673 1113 3687 1127
rect 3893 1113 3907 1127
rect 4153 1113 4167 1127
rect 4273 1113 4287 1127
rect 4393 1113 4407 1127
rect 4433 1113 4447 1127
rect 4453 1113 4467 1127
rect 4493 1113 4507 1127
rect 4553 1113 4567 1127
rect 4593 1113 4607 1127
rect 33 1093 47 1107
rect 113 1093 127 1107
rect 173 1093 187 1107
rect 213 1093 227 1107
rect 273 1093 287 1107
rect 313 1093 327 1107
rect 413 1093 427 1107
rect 453 1093 467 1107
rect 493 1093 507 1107
rect 933 1093 947 1107
rect 993 1093 1007 1107
rect 1133 1093 1147 1107
rect 1253 1093 1267 1107
rect 1293 1093 1307 1107
rect 1613 1093 1627 1107
rect 1673 1093 1687 1107
rect 2073 1093 2087 1107
rect 2293 1093 2307 1107
rect 2593 1093 2607 1107
rect 2653 1093 2667 1107
rect 2693 1093 2707 1107
rect 2753 1093 2767 1107
rect 2793 1093 2807 1107
rect 2973 1093 2987 1107
rect 3133 1093 3147 1107
rect 3173 1093 3187 1107
rect 3273 1093 3287 1107
rect 3353 1093 3367 1107
rect 3433 1093 3447 1107
rect 3493 1093 3507 1107
rect 3573 1093 3587 1107
rect 3653 1093 3667 1107
rect 3693 1093 3707 1107
rect 3773 1093 3787 1107
rect 3813 1093 3827 1107
rect 3833 1093 3847 1107
rect 3873 1093 3887 1107
rect 3953 1093 3967 1107
rect 4033 1093 4047 1107
rect 4073 1093 4087 1107
rect 4093 1093 4107 1107
rect 4133 1093 4147 1107
rect 4213 1093 4227 1107
rect 4293 1093 4307 1107
rect 4333 1093 4347 1107
rect 4373 1093 4387 1107
rect 4413 1093 4427 1107
rect 4473 1093 4487 1107
rect 4513 1093 4527 1107
rect 4673 1093 4687 1107
rect 4733 1093 4747 1107
rect 93 1073 107 1087
rect 133 1073 147 1087
rect 693 1073 707 1087
rect 1653 1073 1667 1087
rect 1693 1073 1707 1087
rect 2953 1073 2967 1087
rect 2993 1073 3007 1087
rect 3053 1073 3067 1087
rect 3333 1073 3347 1087
rect 3373 1073 3387 1087
rect 3413 1073 3427 1087
rect 3453 1073 3467 1087
rect 3473 1073 3487 1087
rect 3513 1073 3527 1087
rect 3553 1073 3567 1087
rect 3593 1073 3607 1087
rect 3753 1073 3767 1087
rect 3793 1073 3807 1087
rect 4013 1073 4027 1087
rect 4053 1073 4067 1087
rect 4653 1073 4667 1087
rect 4693 1073 4707 1087
rect 253 853 267 867
rect 293 853 307 867
rect 673 853 687 867
rect 713 853 727 867
rect 1193 853 1207 867
rect 1233 853 1247 867
rect 1273 853 1287 867
rect 1313 853 1327 867
rect 1353 853 1367 867
rect 1393 853 1407 867
rect 1553 853 1567 867
rect 1933 853 1947 867
rect 1973 853 1987 867
rect 2373 853 2387 867
rect 2413 853 2427 867
rect 2993 853 3007 867
rect 3033 853 3047 867
rect 3153 853 3167 867
rect 3193 853 3207 867
rect 3313 853 3327 867
rect 3353 853 3367 867
rect 3393 853 3407 867
rect 3433 853 3447 867
rect 3553 853 3567 867
rect 3593 853 3607 867
rect 3653 853 3667 867
rect 3693 853 3707 867
rect 3753 853 3767 867
rect 3793 853 3807 867
rect 3833 853 3847 867
rect 3873 853 3887 867
rect 3933 853 3947 867
rect 3973 853 3987 867
rect 4393 853 4407 867
rect 4433 853 4447 867
rect 4493 853 4507 867
rect 4533 853 4547 867
rect 4693 853 4707 867
rect 4733 853 4747 867
rect 273 833 287 847
rect 353 833 367 847
rect 393 833 407 847
rect 693 833 707 847
rect 773 833 787 847
rect 813 833 827 847
rect 873 833 887 847
rect 913 833 927 847
rect 973 833 987 847
rect 1213 833 1227 847
rect 1293 833 1307 847
rect 1373 833 1387 847
rect 1453 833 1467 847
rect 1493 833 1507 847
rect 1613 833 1627 847
rect 1653 833 1667 847
rect 1733 833 1747 847
rect 1873 833 1887 847
rect 1953 833 1967 847
rect 2093 833 2107 847
rect 2133 833 2147 847
rect 2193 833 2207 847
rect 2233 833 2247 847
rect 2293 833 2307 847
rect 2333 833 2347 847
rect 2393 833 2407 847
rect 2473 833 2487 847
rect 2773 833 2787 847
rect 2813 833 2827 847
rect 2873 833 2887 847
rect 2933 833 2947 847
rect 2973 833 2987 847
rect 3013 833 3027 847
rect 3093 833 3107 847
rect 3173 833 3187 847
rect 3273 833 3287 847
rect 3333 833 3347 847
rect 3413 833 3427 847
rect 3573 833 3587 847
rect 3673 833 3687 847
rect 3713 833 3727 847
rect 3773 833 3787 847
rect 3813 833 3827 847
rect 3853 833 3867 847
rect 3953 833 3967 847
rect 3993 833 4007 847
rect 4033 833 4047 847
rect 4093 833 4107 847
rect 4133 833 4147 847
rect 4193 833 4207 847
rect 4233 833 4247 847
rect 4313 833 4327 847
rect 4353 833 4367 847
rect 4373 833 4387 847
rect 4413 833 4427 847
rect 4513 833 4527 847
rect 4553 833 4567 847
rect 4613 833 4627 847
rect 4653 833 4667 847
rect 4673 833 4687 847
rect 4713 833 4727 847
rect 93 813 107 827
rect 133 813 147 827
rect 213 813 227 827
rect 373 813 387 827
rect 413 813 427 827
rect 513 813 527 827
rect 553 813 567 827
rect 633 813 647 827
rect 793 813 807 827
rect 833 813 847 827
rect 893 813 907 827
rect 933 813 947 827
rect 1033 813 1047 827
rect 1073 813 1087 827
rect 1093 813 1107 827
rect 1133 813 1147 827
rect 1433 813 1447 827
rect 1533 813 1547 827
rect 1593 813 1607 827
rect 1673 813 1687 827
rect 2013 813 2027 827
rect 2053 813 2067 827
rect 2073 813 2087 827
rect 2113 813 2127 827
rect 2173 813 2187 827
rect 2213 813 2227 827
rect 2273 813 2287 827
rect 2313 813 2327 827
rect 2533 813 2547 827
rect 2613 813 2627 827
rect 2653 813 2667 827
rect 2793 813 2807 827
rect 2833 813 2847 827
rect 3233 813 3247 827
rect 3493 813 3507 827
rect 3533 813 3547 827
rect 4113 813 4127 827
rect 4153 813 4167 827
rect 4213 813 4227 827
rect 4253 813 4267 827
rect 4293 813 4307 827
rect 4593 813 4607 827
rect 993 793 1007 807
rect 1053 793 1067 807
rect 1113 793 1127 807
rect 1473 793 1487 807
rect 1633 793 1647 807
rect 2033 793 2047 807
rect 2493 793 2507 807
rect 2893 793 2907 807
rect 2913 793 2927 807
rect 3073 793 3087 807
rect 3213 793 3227 807
rect 3513 793 3527 807
rect 4053 793 4067 807
rect 4333 793 4347 807
rect 4633 793 4647 807
rect 253 653 267 667
rect 613 653 627 667
rect 1013 653 1027 667
rect 1053 653 1067 667
rect 1373 653 1387 667
rect 1873 653 1887 667
rect 1953 653 1967 667
rect 2033 653 2047 667
rect 2073 653 2087 667
rect 2573 653 2587 667
rect 2653 653 2667 667
rect 2753 653 2767 667
rect 2793 653 2807 667
rect 3173 653 3187 667
rect 3193 653 3207 667
rect 3393 653 3407 667
rect 3553 653 3567 667
rect 3693 653 3707 667
rect 4053 653 4067 667
rect 4513 653 4527 667
rect 93 633 107 647
rect 133 633 147 647
rect 213 633 227 647
rect 313 633 327 647
rect 353 633 367 647
rect 493 633 507 647
rect 533 633 547 647
rect 653 633 667 647
rect 733 633 747 647
rect 773 633 787 647
rect 873 633 887 647
rect 913 633 927 647
rect 993 633 1007 647
rect 1033 633 1047 647
rect 1073 633 1087 647
rect 1193 633 1207 647
rect 1233 633 1247 647
rect 1273 633 1287 647
rect 1333 633 1347 647
rect 1353 633 1367 647
rect 1393 633 1407 647
rect 1433 633 1447 647
rect 1473 633 1487 647
rect 1593 633 1607 647
rect 1633 633 1647 647
rect 1713 633 1727 647
rect 1753 633 1767 647
rect 1793 633 1807 647
rect 1853 633 1867 647
rect 1893 633 1907 647
rect 1933 633 1947 647
rect 1973 633 1987 647
rect 2053 633 2067 647
rect 2093 633 2107 647
rect 2153 633 2167 647
rect 2233 633 2247 647
rect 2273 633 2287 647
rect 2373 633 2387 647
rect 2413 633 2427 647
rect 2453 633 2467 647
rect 2553 633 2567 647
rect 2613 633 2627 647
rect 2713 633 2727 647
rect 2893 633 2907 647
rect 2933 633 2947 647
rect 2953 633 2967 647
rect 2993 633 3007 647
rect 3373 633 3387 647
rect 3413 633 3427 647
rect 3433 633 3447 647
rect 3473 633 3487 647
rect 3593 633 3607 647
rect 3653 633 3667 647
rect 3753 633 3767 647
rect 3793 633 3807 647
rect 3833 633 3847 647
rect 4613 633 4627 647
rect 4653 633 4667 647
rect 4673 633 4687 647
rect 4713 633 4727 647
rect 273 613 287 627
rect 333 613 347 627
rect 373 613 387 627
rect 433 613 447 627
rect 593 613 607 627
rect 893 613 907 627
rect 933 613 947 627
rect 1113 613 1127 627
rect 1173 613 1187 627
rect 1213 613 1227 627
rect 2013 613 2027 627
rect 2393 613 2407 627
rect 2433 613 2447 627
rect 2513 613 2527 627
rect 2633 613 2647 627
rect 2673 613 2687 627
rect 2733 613 2747 627
rect 2773 613 2787 627
rect 2813 613 2827 627
rect 2873 613 2887 627
rect 2913 613 2927 627
rect 2973 613 2987 627
rect 3013 613 3027 627
rect 3073 613 3087 627
rect 3153 613 3167 627
rect 3213 613 3227 627
rect 3293 613 3307 627
rect 3333 613 3347 627
rect 3453 613 3467 627
rect 3493 613 3507 627
rect 3533 613 3547 627
rect 3573 613 3587 627
rect 3673 613 3687 627
rect 3713 613 3727 627
rect 3773 613 3787 627
rect 3813 613 3827 627
rect 3893 613 3907 627
rect 3933 613 3947 627
rect 3993 613 4007 627
rect 4033 613 4047 627
rect 4073 613 4087 627
rect 4113 613 4127 627
rect 4153 613 4167 627
rect 4213 613 4227 627
rect 4253 613 4267 627
rect 4353 613 4367 627
rect 4393 613 4407 627
rect 4453 613 4467 627
rect 4493 613 4507 627
rect 4533 613 4547 627
rect 4593 613 4607 627
rect 4633 613 4647 627
rect 4693 613 4707 627
rect 4733 613 4747 627
rect 413 593 427 607
rect 453 593 467 607
rect 1293 593 1307 607
rect 3053 593 3067 607
rect 3093 593 3107 607
rect 3273 593 3287 607
rect 3313 593 3327 607
rect 3873 593 3887 607
rect 3913 593 3927 607
rect 3973 593 3987 607
rect 4013 593 4027 607
rect 4133 593 4147 607
rect 4173 593 4187 607
rect 4233 593 4247 607
rect 4273 593 4287 607
rect 4333 593 4347 607
rect 4373 593 4387 607
rect 4433 593 4447 607
rect 4473 593 4487 607
rect 253 373 267 387
rect 293 373 307 387
rect 493 373 507 387
rect 533 373 547 387
rect 1033 373 1047 387
rect 1073 373 1087 387
rect 1553 373 1567 387
rect 1593 373 1607 387
rect 1893 373 1907 387
rect 1933 373 1947 387
rect 2513 373 2527 387
rect 2553 373 2567 387
rect 2813 373 2827 387
rect 2853 373 2867 387
rect 3173 373 3187 387
rect 3213 373 3227 387
rect 3273 373 3287 387
rect 3313 373 3327 387
rect 3513 373 3527 387
rect 3553 373 3567 387
rect 3593 373 3607 387
rect 3633 373 3647 387
rect 3973 373 3987 387
rect 4233 373 4247 387
rect 4273 373 4287 387
rect 273 353 287 367
rect 353 353 367 367
rect 393 353 407 367
rect 453 353 467 367
rect 513 353 527 367
rect 593 353 607 367
rect 633 353 647 367
rect 693 353 707 367
rect 733 353 747 367
rect 793 353 807 367
rect 833 353 847 367
rect 893 353 907 367
rect 933 353 947 367
rect 993 353 1007 367
rect 1053 353 1067 367
rect 1153 353 1167 367
rect 1193 353 1207 367
rect 1233 353 1247 367
rect 1293 353 1307 367
rect 1333 353 1347 367
rect 1473 353 1487 367
rect 1513 353 1527 367
rect 1573 353 1587 367
rect 1913 353 1927 367
rect 1973 353 1987 367
rect 2013 353 2027 367
rect 2313 353 2327 367
rect 2453 353 2467 367
rect 2533 353 2547 367
rect 2833 353 2847 367
rect 2913 353 2927 367
rect 2953 353 2967 367
rect 3113 353 3127 367
rect 3193 353 3207 367
rect 3233 353 3247 367
rect 3293 353 3307 367
rect 3333 353 3347 367
rect 3373 353 3387 367
rect 3413 353 3427 367
rect 3473 353 3487 367
rect 3533 353 3547 367
rect 3613 353 3627 367
rect 3693 353 3707 367
rect 3733 353 3747 367
rect 4153 353 4167 367
rect 4193 353 4207 367
rect 4253 353 4267 367
rect 4293 353 4307 367
rect 4313 353 4327 367
rect 4353 353 4367 367
rect 4433 353 4447 367
rect 4493 353 4507 367
rect 4533 353 4547 367
rect 4593 353 4607 367
rect 4653 353 4667 367
rect 4713 353 4727 367
rect 93 333 107 347
rect 133 333 147 347
rect 213 333 227 347
rect 373 333 387 347
rect 413 333 427 347
rect 613 333 627 347
rect 653 333 667 347
rect 673 333 687 347
rect 713 333 727 347
rect 773 333 787 347
rect 813 333 827 347
rect 913 333 927 347
rect 953 333 967 347
rect 1133 333 1147 347
rect 1313 333 1327 347
rect 1353 333 1367 347
rect 1393 333 1407 347
rect 1433 333 1447 347
rect 1453 333 1467 347
rect 1493 333 1507 347
rect 1653 333 1667 347
rect 1733 333 1747 347
rect 1773 333 1787 347
rect 1993 333 2007 347
rect 2033 333 2047 347
rect 2133 333 2147 347
rect 2173 333 2187 347
rect 2253 333 2267 347
rect 2353 333 2367 347
rect 2393 333 2407 347
rect 2593 333 2607 347
rect 2673 333 2687 347
rect 2713 333 2727 347
rect 2893 333 2907 347
rect 2933 333 2947 347
rect 2973 333 2987 347
rect 3013 333 3027 347
rect 3053 333 3067 347
rect 3353 333 3367 347
rect 3393 333 3407 347
rect 3673 333 3687 347
rect 3713 333 3727 347
rect 3793 333 3807 347
rect 3833 333 3847 347
rect 3873 333 3887 347
rect 3913 333 3927 347
rect 3933 333 3947 347
rect 3993 333 4007 347
rect 4033 333 4047 347
rect 4073 333 4087 347
rect 4133 333 4147 347
rect 4373 333 4387 347
rect 4513 333 4527 347
rect 4553 333 4567 347
rect 433 313 447 327
rect 973 313 987 327
rect 1173 313 1187 327
rect 1253 313 1267 327
rect 1413 313 1427 327
rect 2333 313 2347 327
rect 2373 313 2387 327
rect 2433 313 2447 327
rect 3033 313 3047 327
rect 3093 313 3107 327
rect 3493 313 3507 327
rect 3813 313 3827 327
rect 3893 313 3907 327
rect 4053 313 4067 327
rect 4173 313 4187 327
rect 4333 313 4347 327
rect 4413 313 4427 327
rect 4573 313 4587 327
rect 4633 313 4647 327
rect 4693 313 4707 327
rect 393 173 407 187
rect 633 173 647 187
rect 713 173 727 187
rect 1133 173 1147 187
rect 1193 173 1207 187
rect 1273 173 1287 187
rect 1433 173 1447 187
rect 1493 173 1507 187
rect 1533 173 1547 187
rect 1653 173 1667 187
rect 2033 173 2047 187
rect 2113 173 2127 187
rect 2193 173 2207 187
rect 2293 173 2307 187
rect 2353 173 2367 187
rect 2453 173 2467 187
rect 3153 173 3167 187
rect 3313 173 3327 187
rect 3553 173 3567 187
rect 3633 173 3647 187
rect 3713 173 3727 187
rect 3753 173 3767 187
rect 3933 173 3947 187
rect 4693 173 4707 187
rect 93 153 107 167
rect 133 153 147 167
rect 213 153 227 167
rect 253 153 267 167
rect 293 153 307 167
rect 333 153 347 167
rect 373 153 387 167
rect 413 153 427 167
rect 613 153 627 167
rect 673 153 687 167
rect 773 153 787 167
rect 853 153 867 167
rect 893 153 907 167
rect 1033 153 1047 167
rect 1073 153 1087 167
rect 1173 153 1187 167
rect 1213 153 1227 167
rect 1333 153 1347 167
rect 1373 153 1387 167
rect 1513 153 1527 167
rect 1553 153 1567 167
rect 1613 153 1627 167
rect 1773 153 1787 167
rect 1813 153 1827 167
rect 1893 153 1907 167
rect 1973 153 1987 167
rect 2013 153 2027 167
rect 2093 153 2107 167
rect 2133 153 2147 167
rect 2173 153 2187 167
rect 2213 153 2227 167
rect 2273 153 2287 167
rect 2313 153 2327 167
rect 2333 153 2347 167
rect 2373 153 2387 167
rect 2493 153 2507 167
rect 2573 153 2587 167
rect 2613 153 2627 167
rect 2733 153 2747 167
rect 2813 153 2827 167
rect 2853 153 2867 167
rect 2953 153 2967 167
rect 2993 153 3007 167
rect 3033 153 3047 167
rect 3133 153 3147 167
rect 3173 153 3187 167
rect 3213 153 3227 167
rect 3593 153 3607 167
rect 3693 153 3707 167
rect 3733 153 3747 167
rect 3813 153 3827 167
rect 3853 153 3867 167
rect 3913 153 3927 167
rect 3953 153 3967 167
rect 4653 153 4667 167
rect 273 133 287 147
rect 313 133 327 147
rect 453 133 467 147
rect 493 133 507 147
rect 573 133 587 147
rect 693 133 707 147
rect 733 133 747 147
rect 1013 133 1027 147
rect 1053 133 1067 147
rect 1113 133 1127 147
rect 1253 133 1267 147
rect 1313 133 1327 147
rect 1353 133 1367 147
rect 1413 133 1427 147
rect 1473 133 1487 147
rect 1633 133 1647 147
rect 1673 133 1687 147
rect 1953 133 1967 147
rect 1993 133 2007 147
rect 2053 133 2067 147
rect 2433 133 2447 147
rect 2973 133 2987 147
rect 3013 133 3027 147
rect 3093 133 3107 147
rect 3193 133 3207 147
rect 3233 133 3247 147
rect 3293 133 3307 147
rect 3353 133 3367 147
rect 3453 133 3467 147
rect 3493 133 3507 147
rect 3533 133 3547 147
rect 3613 133 3627 147
rect 3653 133 3667 147
rect 3773 133 3787 147
rect 3833 133 3847 147
rect 3873 133 3887 147
rect 4033 133 4047 147
rect 4073 133 4087 147
rect 4113 133 4127 147
rect 4213 133 4227 147
rect 4253 133 4267 147
rect 4313 133 4327 147
rect 4393 133 4407 147
rect 4433 133 4447 147
rect 4473 133 4487 147
rect 4533 133 4547 147
rect 4573 133 4587 147
rect 4673 133 4687 147
rect 4713 133 4727 147
rect 473 113 487 127
rect 513 113 527 127
rect 3333 113 3347 127
rect 3373 113 3387 127
rect 3433 113 3447 127
rect 3473 113 3487 127
rect 4013 113 4027 127
rect 4053 113 4067 127
rect 4093 113 4107 127
rect 4133 113 4147 127
rect 4193 113 4207 127
rect 4233 113 4247 127
rect 4293 113 4307 127
rect 4333 113 4347 127
rect 4373 113 4387 127
rect 4413 113 4427 127
rect 4453 113 4467 127
rect 4493 113 4507 127
rect 4553 113 4567 127
rect 4593 113 4607 127
<< labels >>
flabel metal1 s 4782 2 4842 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 3497 -23 3503 -17 7 FreeSans 16 270 0 0 Cin[5]
port 2 nsew
flabel metal2 s 3577 -23 3583 -17 7 FreeSans 16 270 0 0 Cin[4]
port 3 nsew
flabel metal2 s 3617 -23 3623 -17 7 FreeSans 16 270 0 0 Cin[3]
port 4 nsew
flabel metal2 s 4137 -23 4143 -17 7 FreeSans 16 270 0 0 Cin[2]
port 5 nsew
flabel metal2 s 4177 -23 4183 -17 7 FreeSans 16 270 0 0 Cin[1]
port 6 nsew
flabel metal2 s 4217 -23 4223 -17 7 FreeSans 16 270 0 0 Cin[0]
port 7 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal2 s 3157 4617 3163 4623 3 FreeSans 16 90 0 0 Vld
port 9 nsew
flabel metal3 s -24 2556 -16 2564 7 FreeSans 16 0 0 0 Xin[3]
port 10 nsew
flabel metal3 s -24 2516 -16 2524 7 FreeSans 16 0 0 0 Xin[2]
port 11 nsew
flabel metal3 s -24 2276 -16 2284 7 FreeSans 16 0 0 0 Xin[1]
port 12 nsew
flabel metal3 s -24 2096 -16 2104 7 FreeSans 16 0 0 0 Xin[0]
port 13 nsew
flabel metal2 s 2757 4617 2763 4623 3 FreeSans 16 90 0 0 Xout[3]
port 14 nsew
flabel metal2 s 2837 4617 2843 4623 3 FreeSans 16 90 0 0 Xout[2]
port 15 nsew
flabel metal2 s 2877 4617 2883 4623 3 FreeSans 16 90 0 0 Xout[1]
port 16 nsew
flabel metal2 s 3117 4617 3123 4623 3 FreeSans 16 90 0 0 Xout[0]
port 17 nsew
flabel metal3 s 4816 2996 4824 3004 3 FreeSans 16 0 0 0 Yin[3]
port 18 nsew
flabel metal3 s 4816 2276 4824 2284 3 FreeSans 16 0 0 0 Yin[2]
port 19 nsew
flabel metal3 s 4816 2236 4824 2244 3 FreeSans 16 0 0 0 Yin[1]
port 20 nsew
flabel metal3 s 4816 2036 4824 2044 3 FreeSans 16 0 0 0 Yin[0]
port 21 nsew
flabel metal2 s 37 4617 43 4623 3 FreeSans 16 90 0 0 Yout[3]
port 22 nsew
flabel metal2 s 497 4617 503 4623 3 FreeSans 16 90 0 0 Yout[2]
port 23 nsew
flabel metal2 s 537 4617 543 4623 3 FreeSans 16 90 0 0 Yout[1]
port 24 nsew
flabel metal2 s 577 4617 583 4623 3 FreeSans 16 90 0 0 Yout[0]
port 25 nsew
flabel metal3 s -24 2056 -16 2064 7 FreeSans 16 0 0 0 clk
port 26 nsew
rlabel metal1 4 242 256 258 0 _1573_.gnd
rlabel metal1 4 2 256 18 0 _1573_.vdd
rlabel metal2 93 153 107 167 0 _1573_.D
rlabel metal2 133 153 147 167 0 _1573_.CLK
rlabel metal2 213 153 227 167 0 _1573_.Q
rlabel metal1 4 242 256 258 0 _1544_.gnd
rlabel metal1 4 482 256 498 0 _1544_.vdd
rlabel metal2 93 333 107 347 0 _1544_.D
rlabel metal2 133 333 147 347 0 _1544_.CLK
rlabel metal2 213 333 227 347 0 _1544_.Q
rlabel metal1 244 242 336 258 0 _1464_.gnd
rlabel metal1 244 482 336 498 0 _1464_.vdd
rlabel metal2 253 373 267 387 0 _1464_.A
rlabel metal2 293 373 307 387 0 _1464_.B
rlabel metal2 273 353 287 367 0 _1464_.Y
rlabel metal1 244 242 376 258 0 _1463_.gnd
rlabel metal1 244 2 376 18 0 _1463_.vdd
rlabel metal2 253 153 267 167 0 _1463_.A
rlabel metal2 273 133 287 147 0 _1463_.B
rlabel metal2 333 153 347 167 0 _1463_.C
rlabel metal2 313 133 327 147 0 _1463_.D
rlabel metal2 293 153 307 167 0 _1463_.Y
rlabel metal1 324 242 436 258 0 _1473_.gnd
rlabel metal1 324 482 436 498 0 _1473_.vdd
rlabel metal2 413 333 427 347 0 _1473_.A
rlabel metal2 393 353 407 367 0 _1473_.B
rlabel metal2 353 353 367 367 0 _1473_.C
rlabel metal2 373 333 387 347 0 _1473_.Y
rlabel metal1 484 242 576 258 0 _1477_.gnd
rlabel metal1 484 482 576 498 0 _1477_.vdd
rlabel metal2 493 373 507 387 0 _1477_.A
rlabel metal2 533 373 547 387 0 _1477_.B
rlabel metal2 513 353 527 367 0 _1477_.Y
rlabel metal1 364 242 456 258 0 _1469_.gnd
rlabel metal1 364 2 456 18 0 _1469_.vdd
rlabel metal2 413 153 427 167 0 _1469_.B
rlabel metal2 373 153 387 167 0 _1469_.A
rlabel metal2 393 173 407 187 0 _1469_.Y
rlabel metal1 424 242 496 258 0 _845_.gnd
rlabel metal1 424 482 496 498 0 _845_.vdd
rlabel metal2 433 313 447 327 0 _845_.A
rlabel metal2 453 353 467 367 0 _845_.Y
rlabel metal1 444 242 556 258 0 _1475_.gnd
rlabel metal1 444 2 556 18 0 _1475_.vdd
rlabel metal2 453 133 467 147 0 _1475_.A
rlabel metal2 473 113 487 127 0 _1475_.B
rlabel metal2 493 133 507 147 0 _1475_.C
rlabel metal2 513 113 527 127 0 _1475_.Y
rlabel metal1 744 242 996 258 0 _1545_.gnd
rlabel metal1 744 2 996 18 0 _1545_.vdd
rlabel metal2 893 153 907 167 0 _1545_.D
rlabel metal2 853 153 867 167 0 _1545_.CLK
rlabel metal2 773 153 787 167 0 _1545_.Q
rlabel metal1 764 242 876 258 0 _1476_.gnd
rlabel metal1 764 482 876 498 0 _1476_.vdd
rlabel metal2 773 333 787 347 0 _1476_.A
rlabel metal2 793 353 807 367 0 _1476_.B
rlabel metal2 833 353 847 367 0 _1476_.C
rlabel metal2 813 333 827 347 0 _1476_.Y
rlabel metal1 564 242 676 258 0 _1472_.gnd
rlabel metal1 564 482 676 498 0 _1472_.vdd
rlabel metal2 653 333 667 347 0 _1472_.A
rlabel metal2 633 353 647 367 0 _1472_.B
rlabel metal2 593 353 607 367 0 _1472_.C
rlabel metal2 613 333 627 347 0 _1472_.Y
rlabel metal1 664 242 776 258 0 _847_.gnd
rlabel metal1 664 482 776 498 0 _847_.vdd
rlabel metal2 673 333 687 347 0 _847_.A
rlabel metal2 693 353 707 367 0 _847_.B
rlabel metal2 733 353 747 367 0 _847_.C
rlabel metal2 713 333 727 347 0 _847_.Y
rlabel metal1 644 242 756 258 0 _1462_.gnd
rlabel metal1 644 2 756 18 0 _1462_.vdd
rlabel metal2 733 133 747 147 0 _1462_.A
rlabel metal2 713 173 727 187 0 _1462_.B
rlabel metal2 693 133 707 147 0 _1462_.C
rlabel metal2 673 153 687 167 0 _1462_.Y
rlabel metal1 544 242 656 258 0 _1461_.gnd
rlabel metal1 544 2 656 18 0 _1461_.vdd
rlabel metal2 633 173 647 187 0 _1461_.A
rlabel metal2 613 153 627 167 0 _1461_.B
rlabel metal2 573 133 587 147 0 _1461_.Y
rlabel metal1 984 242 1096 258 0 _1468_.gnd
rlabel metal1 984 2 1096 18 0 _1468_.vdd
rlabel metal2 1073 153 1087 167 0 _1468_.A
rlabel metal2 1053 133 1067 147 0 _1468_.B
rlabel metal2 1013 133 1027 147 0 _1468_.C
rlabel metal2 1033 153 1047 167 0 _1468_.Y
rlabel metal1 864 242 976 258 0 _850_.gnd
rlabel metal1 864 482 976 498 0 _850_.vdd
rlabel metal2 953 333 967 347 0 _850_.A
rlabel metal2 933 353 947 367 0 _850_.B
rlabel metal2 893 353 907 367 0 _850_.C
rlabel metal2 913 333 927 347 0 _850_.Y
rlabel metal1 1024 242 1116 258 0 _846_.gnd
rlabel metal1 1024 482 1116 498 0 _846_.vdd
rlabel metal2 1033 373 1047 387 0 _846_.A
rlabel metal2 1073 373 1087 387 0 _846_.B
rlabel metal2 1053 353 1067 367 0 _846_.Y
rlabel metal1 964 242 1036 258 0 _848_.gnd
rlabel metal1 964 482 1036 498 0 _848_.vdd
rlabel metal2 973 313 987 327 0 _848_.A
rlabel metal2 993 353 1007 367 0 _848_.Y
rlabel metal1 1284 242 1396 258 0 _1456_.gnd
rlabel metal1 1284 2 1396 18 0 _1456_.vdd
rlabel metal2 1373 153 1387 167 0 _1456_.A
rlabel metal2 1353 133 1367 147 0 _1456_.B
rlabel metal2 1313 133 1327 147 0 _1456_.C
rlabel metal2 1333 153 1347 167 0 _1456_.Y
rlabel metal1 1264 242 1376 258 0 _1452_.gnd
rlabel metal1 1264 482 1376 498 0 _1452_.vdd
rlabel metal2 1353 333 1367 347 0 _1452_.A
rlabel metal2 1333 353 1347 367 0 _1452_.B
rlabel metal2 1293 353 1307 367 0 _1452_.C
rlabel metal2 1313 333 1327 347 0 _1452_.Y
rlabel metal1 1104 242 1216 258 0 _1471_.gnd
rlabel metal1 1104 482 1216 498 0 _1471_.vdd
rlabel metal2 1193 353 1207 367 0 _1471_.A
rlabel metal2 1173 313 1187 327 0 _1471_.B
rlabel metal2 1153 353 1167 367 0 _1471_.C
rlabel metal2 1133 333 1147 347 0 _1471_.Y
rlabel metal1 1144 242 1236 258 0 _1466_.gnd
rlabel metal1 1144 2 1236 18 0 _1466_.vdd
rlabel metal2 1173 153 1187 167 0 _1466_.B
rlabel metal2 1213 153 1227 167 0 _1466_.A
rlabel metal2 1193 173 1207 187 0 _1466_.Y
rlabel metal1 1204 242 1276 258 0 _1470_.gnd
rlabel metal1 1204 482 1276 498 0 _1470_.vdd
rlabel metal2 1253 313 1267 327 0 _1470_.A
rlabel metal2 1233 353 1247 367 0 _1470_.Y
rlabel metal1 1084 242 1156 258 0 _1467_.gnd
rlabel metal1 1084 2 1156 18 0 _1467_.vdd
rlabel metal2 1133 173 1147 187 0 _1467_.A
rlabel metal2 1113 133 1127 147 0 _1467_.Y
rlabel metal1 1224 242 1296 258 0 _1460_.gnd
rlabel metal1 1224 2 1296 18 0 _1460_.vdd
rlabel metal2 1273 173 1287 187 0 _1460_.A
rlabel metal2 1253 133 1267 147 0 _1460_.Y
rlabel metal1 1444 242 1556 258 0 _1453_.gnd
rlabel metal1 1444 482 1556 498 0 _1453_.vdd
rlabel metal2 1453 333 1467 347 0 _1453_.A
rlabel metal2 1473 353 1487 367 0 _1453_.B
rlabel metal2 1513 353 1527 367 0 _1453_.C
rlabel metal2 1493 333 1507 347 0 _1453_.Y
rlabel metal1 1544 242 1636 258 0 _1438_.gnd
rlabel metal1 1544 482 1636 498 0 _1438_.vdd
rlabel metal2 1553 373 1567 387 0 _1438_.A
rlabel metal2 1593 373 1607 387 0 _1438_.B
rlabel metal2 1573 353 1587 367 0 _1438_.Y
rlabel metal1 1584 242 1696 258 0 _1465_.gnd
rlabel metal1 1584 2 1696 18 0 _1465_.vdd
rlabel metal2 1673 133 1687 147 0 _1465_.A
rlabel metal2 1653 173 1667 187 0 _1465_.B
rlabel metal2 1633 133 1647 147 0 _1465_.C
rlabel metal2 1613 153 1627 167 0 _1465_.Y
rlabel metal1 1364 242 1456 258 0 _1449_.gnd
rlabel metal1 1364 482 1456 498 0 _1449_.vdd
rlabel metal2 1393 333 1407 347 0 _1449_.B
rlabel metal2 1433 333 1447 347 0 _1449_.A
rlabel metal2 1413 313 1427 327 0 _1449_.Y
rlabel metal1 1504 242 1596 258 0 _1448_.gnd
rlabel metal1 1504 2 1596 18 0 _1448_.vdd
rlabel metal2 1553 153 1567 167 0 _1448_.B
rlabel metal2 1513 153 1527 167 0 _1448_.A
rlabel metal2 1533 173 1547 187 0 _1448_.Y
rlabel metal1 1444 242 1516 258 0 _1455_.gnd
rlabel metal1 1444 2 1516 18 0 _1455_.vdd
rlabel metal2 1493 173 1507 187 0 _1455_.A
rlabel metal2 1473 133 1487 147 0 _1455_.Y
rlabel metal1 1384 242 1456 258 0 _1451_.gnd
rlabel metal1 1384 2 1456 18 0 _1451_.vdd
rlabel metal2 1433 173 1447 187 0 _1451_.A
rlabel metal2 1413 133 1427 147 0 _1451_.Y
rlabel metal1 1624 242 1876 258 0 _1572_.gnd
rlabel metal1 1624 482 1876 498 0 _1572_.vdd
rlabel metal2 1773 333 1787 347 0 _1572_.D
rlabel metal2 1733 333 1747 347 0 _1572_.CLK
rlabel metal2 1653 333 1667 347 0 _1572_.Q
rlabel metal1 1684 242 1936 258 0 _1542_.gnd
rlabel metal1 1684 2 1936 18 0 _1542_.vdd
rlabel metal2 1773 153 1787 167 0 _1542_.D
rlabel metal2 1813 153 1827 167 0 _1542_.CLK
rlabel metal2 1893 153 1907 167 0 _1542_.Q
rlabel metal1 1864 242 1956 258 0 _840_.gnd
rlabel metal1 1864 482 1956 498 0 _840_.vdd
rlabel metal2 1933 373 1947 387 0 _840_.A
rlabel metal2 1893 373 1907 387 0 _840_.B
rlabel metal2 1913 353 1927 367 0 _840_.Y
rlabel metal1 2044 242 2296 258 0 _1543_.gnd
rlabel metal1 2044 482 2296 498 0 _1543_.vdd
rlabel metal2 2133 333 2147 347 0 _1543_.D
rlabel metal2 2173 333 2187 347 0 _1543_.CLK
rlabel metal2 2253 333 2267 347 0 _1543_.Q
rlabel metal1 1944 242 2056 258 0 _844_.gnd
rlabel metal1 1944 482 2056 498 0 _844_.vdd
rlabel metal2 2033 333 2047 347 0 _844_.A
rlabel metal2 2013 353 2027 367 0 _844_.B
rlabel metal2 1973 353 1987 367 0 _844_.C
rlabel metal2 1993 333 2007 347 0 _844_.Y
rlabel metal1 1924 242 2036 258 0 _841_.gnd
rlabel metal1 1924 2 2036 18 0 _841_.vdd
rlabel metal2 2013 153 2027 167 0 _841_.A
rlabel metal2 1993 133 2007 147 0 _841_.B
rlabel metal2 1953 133 1967 147 0 _841_.C
rlabel metal2 1973 153 1987 167 0 _841_.Y
rlabel metal1 2084 242 2176 258 0 _1446_.gnd
rlabel metal1 2084 2 2176 18 0 _1446_.vdd
rlabel metal2 2133 153 2147 167 0 _1446_.B
rlabel metal2 2093 153 2107 167 0 _1446_.A
rlabel metal2 2113 173 2127 187 0 _1446_.Y
rlabel metal1 2024 242 2096 258 0 _839_.gnd
rlabel metal1 2024 2 2096 18 0 _839_.vdd
rlabel metal2 2033 173 2047 187 0 _839_.A
rlabel metal2 2053 133 2067 147 0 _839_.Y
rlabel metal1 2244 242 2336 258 0 _1459_.gnd
rlabel metal1 2244 2 2336 18 0 _1459_.vdd
rlabel metal2 2273 153 2287 167 0 _1459_.B
rlabel metal2 2313 153 2327 167 0 _1459_.A
rlabel metal2 2293 173 2307 187 0 _1459_.Y
rlabel metal1 2344 242 2436 258 0 _1458_.gnd
rlabel metal1 2344 482 2436 498 0 _1458_.vdd
rlabel metal2 2393 333 2407 347 0 _1458_.B
rlabel metal2 2353 333 2367 347 0 _1458_.A
rlabel metal2 2373 313 2387 327 0 _1458_.Y
rlabel metal1 2324 242 2416 258 0 _1457_.gnd
rlabel metal1 2324 2 2416 18 0 _1457_.vdd
rlabel metal2 2373 153 2387 167 0 _1457_.B
rlabel metal2 2333 153 2347 167 0 _1457_.A
rlabel metal2 2353 173 2367 187 0 _1457_.Y
rlabel metal1 2164 242 2256 258 0 _1447_.gnd
rlabel metal1 2164 2 2256 18 0 _1447_.vdd
rlabel metal2 2213 153 2227 167 0 _1447_.B
rlabel metal2 2173 153 2187 167 0 _1447_.A
rlabel metal2 2193 173 2207 187 0 _1447_.Y
rlabel metal1 2404 242 2476 258 0 _1295_.gnd
rlabel metal1 2404 2 2476 18 0 _1295_.vdd
rlabel metal2 2453 173 2467 187 0 _1295_.A
rlabel metal2 2433 133 2447 147 0 _1295_.Y
rlabel metal1 2284 242 2356 258 0 _842_.gnd
rlabel metal1 2284 482 2356 498 0 _842_.vdd
rlabel metal2 2333 313 2347 327 0 _842_.A
rlabel metal2 2313 353 2327 367 0 _842_.Y
rlabel metal1 2464 242 2716 258 0 _1559_.gnd
rlabel metal1 2464 2 2716 18 0 _1559_.vdd
rlabel metal2 2613 153 2627 167 0 _1559_.D
rlabel metal2 2573 153 2587 167 0 _1559_.CLK
rlabel metal2 2493 153 2507 167 0 _1559_.Q
rlabel metal1 2564 242 2816 258 0 _1557_.gnd
rlabel metal1 2564 482 2816 498 0 _1557_.vdd
rlabel metal2 2713 333 2727 347 0 _1557_.D
rlabel metal2 2673 333 2687 347 0 _1557_.CLK
rlabel metal2 2593 333 2607 347 0 _1557_.Q
rlabel metal1 2484 242 2576 258 0 _1276_.gnd
rlabel metal1 2484 482 2576 498 0 _1276_.vdd
rlabel metal2 2553 373 2567 387 0 _1276_.A
rlabel metal2 2513 373 2527 387 0 _1276_.B
rlabel metal2 2533 353 2547 367 0 _1276_.Y
rlabel metal1 2424 242 2496 258 0 _1312_.gnd
rlabel metal1 2424 482 2496 498 0 _1312_.vdd
rlabel metal2 2433 313 2447 327 0 _1312_.A
rlabel metal2 2453 353 2467 367 0 _1312_.Y
rlabel metal1 2704 242 2956 258 0 _1558_.gnd
rlabel metal1 2704 2 2956 18 0 _1558_.vdd
rlabel metal2 2853 153 2867 167 0 _1558_.D
rlabel metal2 2813 153 2827 167 0 _1558_.CLK
rlabel metal2 2733 153 2747 167 0 _1558_.Q
rlabel metal1 2804 242 2896 258 0 _1294_.gnd
rlabel metal1 2804 482 2896 498 0 _1294_.vdd
rlabel metal2 2813 373 2827 387 0 _1294_.A
rlabel metal2 2853 373 2867 387 0 _1294_.B
rlabel metal2 2833 353 2847 367 0 _1294_.Y
rlabel metal1 2884 242 3016 258 0 _1317_.gnd
rlabel metal1 2884 482 3016 498 0 _1317_.vdd
rlabel metal2 2893 333 2907 347 0 _1317_.A
rlabel metal2 2913 353 2927 367 0 _1317_.B
rlabel metal2 2973 333 2987 347 0 _1317_.C
rlabel metal2 2953 353 2967 367 0 _1317_.D
rlabel metal2 2933 333 2947 347 0 _1317_.Y
rlabel metal1 3164 242 3276 258 0 _1310_.gnd
rlabel metal1 3164 2 3276 18 0 _1310_.vdd
rlabel metal2 3173 153 3187 167 0 _1310_.A
rlabel metal2 3193 133 3207 147 0 _1310_.B
rlabel metal2 3233 133 3247 147 0 _1310_.C
rlabel metal2 3213 153 3227 167 0 _1310_.Y
rlabel metal1 3004 242 3096 258 0 _1316_.gnd
rlabel metal1 3004 482 3096 498 0 _1316_.vdd
rlabel metal2 3053 333 3067 347 0 _1316_.B
rlabel metal2 3013 333 3027 347 0 _1316_.A
rlabel metal2 3033 313 3047 327 0 _1316_.Y
rlabel metal1 3084 242 3156 258 0 _1314_.gnd
rlabel metal1 3084 482 3156 498 0 _1314_.vdd
rlabel metal2 3093 313 3107 327 0 _1314_.A
rlabel metal2 3113 353 3127 367 0 _1314_.Y
rlabel metal1 3144 242 3256 258 0 _1274_.gnd
rlabel metal1 3144 482 3256 498 0 _1274_.vdd
rlabel metal2 3233 353 3247 367 0 _1274_.A
rlabel metal2 3213 373 3227 387 0 _1274_.B
rlabel metal2 3193 353 3207 367 0 _1274_.C
rlabel metal2 3173 373 3187 387 0 _1274_.Y
rlabel metal1 3064 242 3176 258 0 _1313_.gnd
rlabel metal1 3064 2 3176 18 0 _1313_.vdd
rlabel metal2 3153 173 3167 187 0 _1313_.A
rlabel metal2 3133 153 3147 167 0 _1313_.B
rlabel metal2 3093 133 3107 147 0 _1313_.Y
rlabel metal1 2944 242 3076 258 0 _1311_.gnd
rlabel metal1 2944 2 3076 18 0 _1311_.vdd
rlabel metal2 2953 153 2967 167 0 _1311_.A
rlabel metal2 2973 133 2987 147 0 _1311_.B
rlabel metal2 3033 153 3047 167 0 _1311_.C
rlabel metal2 2993 153 3007 167 0 _1311_.Y
rlabel metal2 3013 133 3027 147 0 _1311_.D
rlabel metal1 3344 242 3456 258 0 _1273_.gnd
rlabel metal1 3344 482 3456 498 0 _1273_.vdd
rlabel metal2 3353 333 3367 347 0 _1273_.A
rlabel metal2 3373 353 3387 367 0 _1273_.B
rlabel metal2 3413 353 3427 367 0 _1273_.C
rlabel metal2 3393 333 3407 347 0 _1273_.Y
rlabel metal1 3324 242 3416 258 0 _1308_.gnd
rlabel metal1 3324 2 3416 18 0 _1308_.vdd
rlabel metal2 3333 113 3347 127 0 _1308_.A
rlabel metal2 3373 113 3387 127 0 _1308_.B
rlabel metal2 3353 133 3367 147 0 _1308_.Y
rlabel metal1 3264 242 3336 258 0 _1309_.gnd
rlabel metal1 3264 2 3336 18 0 _1309_.vdd
rlabel metal2 3313 173 3327 187 0 _1309_.A
rlabel metal2 3293 133 3307 147 0 _1309_.Y
rlabel metal1 3444 242 3516 258 0 _1272_.gnd
rlabel metal1 3444 482 3516 498 0 _1272_.vdd
rlabel metal2 3493 313 3507 327 0 _1272_.A
rlabel metal2 3473 353 3487 367 0 _1272_.Y
rlabel metal1 3244 242 3356 258 0 _1293_.gnd
rlabel metal1 3244 482 3356 498 0 _1293_.vdd
rlabel metal2 3333 353 3347 367 0 _1293_.A
rlabel metal2 3313 373 3327 387 0 _1293_.B
rlabel metal2 3293 353 3307 367 0 _1293_.C
rlabel metal2 3273 373 3287 387 0 _1293_.Y
rlabel metal1 3404 242 3516 258 0 _1290_.gnd
rlabel metal1 3404 2 3516 18 0 _1290_.vdd
rlabel metal2 3493 133 3507 147 0 _1290_.A
rlabel metal2 3473 113 3487 127 0 _1290_.B
rlabel metal2 3453 133 3467 147 0 _1290_.C
rlabel metal2 3433 113 3447 127 0 _1290_.Y
rlabel metal1 3664 242 3776 258 0 _1291_.gnd
rlabel metal1 3664 482 3776 498 0 _1291_.vdd
rlabel metal2 3673 333 3687 347 0 _1291_.A
rlabel metal2 3693 353 3707 367 0 _1291_.B
rlabel metal2 3733 353 3747 367 0 _1291_.C
rlabel metal2 3713 333 3727 347 0 _1291_.Y
rlabel metal1 3584 242 3676 258 0 _1292_.gnd
rlabel metal1 3584 482 3676 498 0 _1292_.vdd
rlabel metal2 3593 373 3607 387 0 _1292_.A
rlabel metal2 3633 373 3647 387 0 _1292_.B
rlabel metal2 3613 353 3627 367 0 _1292_.Y
rlabel metal1 3504 242 3596 258 0 _1268_.gnd
rlabel metal1 3504 482 3596 498 0 _1268_.vdd
rlabel metal2 3513 373 3527 387 0 _1268_.A
rlabel metal2 3553 373 3567 387 0 _1268_.B
rlabel metal2 3533 353 3547 367 0 _1268_.Y
rlabel metal1 3564 242 3676 258 0 _1302_.gnd
rlabel metal1 3564 2 3676 18 0 _1302_.vdd
rlabel metal2 3653 133 3667 147 0 _1302_.A
rlabel metal2 3633 173 3647 187 0 _1302_.B
rlabel metal2 3613 133 3627 147 0 _1302_.C
rlabel metal2 3593 153 3607 167 0 _1302_.Y
rlabel metal1 3664 242 3756 258 0 _1297_.gnd
rlabel metal1 3664 2 3756 18 0 _1297_.vdd
rlabel metal2 3693 153 3707 167 0 _1297_.B
rlabel metal2 3733 153 3747 167 0 _1297_.A
rlabel metal2 3713 173 3727 187 0 _1297_.Y
rlabel metal1 3504 242 3576 258 0 _1289_.gnd
rlabel metal1 3504 2 3576 18 0 _1289_.vdd
rlabel metal2 3553 173 3567 187 0 _1289_.A
rlabel metal2 3533 133 3547 147 0 _1289_.Y
rlabel metal1 3804 242 3916 258 0 _1301_.gnd
rlabel metal1 3804 2 3916 18 0 _1301_.vdd
rlabel metal2 3813 153 3827 167 0 _1301_.A
rlabel metal2 3833 133 3847 147 0 _1301_.B
rlabel metal2 3873 133 3887 147 0 _1301_.C
rlabel metal2 3853 153 3867 167 0 _1301_.Y
rlabel metal1 3904 242 3996 258 0 _1300_.gnd
rlabel metal1 3904 2 3996 18 0 _1300_.vdd
rlabel metal2 3953 153 3967 167 0 _1300_.B
rlabel metal2 3913 153 3927 167 0 _1300_.A
rlabel metal2 3933 173 3947 187 0 _1300_.Y
rlabel metal1 3764 242 3856 258 0 _1288_.gnd
rlabel metal1 3764 482 3856 498 0 _1288_.vdd
rlabel metal2 3793 333 3807 347 0 _1288_.B
rlabel metal2 3833 333 3847 347 0 _1288_.A
rlabel metal2 3813 313 3827 327 0 _1288_.Y
rlabel metal1 3844 242 3936 258 0 _1286_.gnd
rlabel metal1 3844 482 3936 498 0 _1286_.vdd
rlabel metal2 3873 333 3887 347 0 _1286_.B
rlabel metal2 3913 333 3927 347 0 _1286_.A
rlabel metal2 3893 313 3907 327 0 _1286_.Y
rlabel metal1 3744 242 3816 258 0 _1298_.gnd
rlabel metal1 3744 2 3816 18 0 _1298_.vdd
rlabel metal2 3753 173 3767 187 0 _1298_.A
rlabel metal2 3773 133 3787 147 0 _1298_.Y
rlabel metal1 3984 242 4096 258 0 _1296_.gnd
rlabel metal1 3984 2 4096 18 0 _1296_.vdd
rlabel metal2 4073 133 4087 147 0 _1296_.A
rlabel metal2 4053 113 4067 127 0 _1296_.B
rlabel metal2 4033 133 4047 147 0 _1296_.C
rlabel metal2 4013 113 4027 127 0 _1296_.Y
rlabel metal1 3924 242 4036 258 0 _1287_.gnd
rlabel metal1 3924 482 4036 498 0 _1287_.vdd
rlabel metal2 3933 333 3947 347 0 _1287_.A
rlabel metal2 3993 333 4007 347 0 _1287_.Y
rlabel metal2 3973 373 3987 387 0 _1287_.B
rlabel metal1 4084 242 4176 258 0 _1267_.gnd
rlabel metal1 4084 2 4176 18 0 _1267_.vdd
rlabel metal2 4093 113 4107 127 0 _1267_.A
rlabel metal2 4133 113 4147 127 0 _1267_.B
rlabel metal2 4113 133 4127 147 0 _1267_.Y
rlabel metal1 4264 242 4356 258 0 _1246_.gnd
rlabel metal1 4264 2 4356 18 0 _1246_.vdd
rlabel metal2 4333 113 4347 127 0 _1246_.A
rlabel metal2 4293 113 4307 127 0 _1246_.B
rlabel metal2 4313 133 4327 147 0 _1246_.Y
rlabel metal1 4104 242 4216 258 0 _1277_.gnd
rlabel metal1 4104 482 4216 498 0 _1277_.vdd
rlabel metal2 4193 353 4207 367 0 _1277_.A
rlabel metal2 4173 313 4187 327 0 _1277_.B
rlabel metal2 4153 353 4167 367 0 _1277_.C
rlabel metal2 4133 333 4147 347 0 _1277_.Y
rlabel metal1 4024 242 4116 258 0 _1299_.gnd
rlabel metal1 4024 482 4116 498 0 _1299_.vdd
rlabel metal2 4073 333 4087 347 0 _1299_.B
rlabel metal2 4033 333 4047 347 0 _1299_.A
rlabel metal2 4053 313 4067 327 0 _1299_.Y
rlabel metal1 4164 242 4276 258 0 _1266_.gnd
rlabel metal1 4164 2 4276 18 0 _1266_.vdd
rlabel metal2 4253 133 4267 147 0 _1266_.A
rlabel metal2 4233 113 4247 127 0 _1266_.B
rlabel metal2 4213 133 4227 147 0 _1266_.C
rlabel metal2 4193 113 4207 127 0 _1266_.Y
rlabel metal1 4204 242 4316 258 0 _1259_.gnd
rlabel metal1 4204 482 4316 498 0 _1259_.vdd
rlabel metal2 4293 353 4307 367 0 _1259_.A
rlabel metal2 4273 373 4287 387 0 _1259_.B
rlabel metal2 4253 353 4267 367 0 _1259_.C
rlabel metal2 4233 373 4247 387 0 _1259_.Y
rlabel metal1 4464 242 4576 258 0 _1261_.gnd
rlabel metal1 4464 482 4576 498 0 _1261_.vdd
rlabel metal2 4553 333 4567 347 0 _1261_.A
rlabel metal2 4533 353 4547 367 0 _1261_.B
rlabel metal2 4493 353 4507 367 0 _1261_.C
rlabel metal2 4513 333 4527 347 0 _1261_.Y
rlabel metal1 4444 242 4536 258 0 _1265_.gnd
rlabel metal1 4444 2 4536 18 0 _1265_.vdd
rlabel metal2 4453 113 4467 127 0 _1265_.A
rlabel metal2 4493 113 4507 127 0 _1265_.B
rlabel metal2 4473 133 4487 147 0 _1265_.Y
rlabel metal1 4304 242 4416 258 0 _1258_.gnd
rlabel metal1 4304 482 4416 498 0 _1258_.vdd
rlabel metal2 4313 353 4327 367 0 _1258_.A
rlabel metal2 4333 313 4347 327 0 _1258_.B
rlabel metal2 4353 353 4367 367 0 _1258_.C
rlabel metal2 4373 333 4387 347 0 _1258_.Y
rlabel metal1 4404 242 4476 258 0 _1248_.gnd
rlabel metal1 4404 482 4476 498 0 _1248_.vdd
rlabel metal2 4413 313 4427 327 0 _1248_.A
rlabel metal2 4433 353 4447 367 0 _1248_.Y
rlabel metal1 4344 242 4456 258 0 _1264_.gnd
rlabel metal1 4344 2 4456 18 0 _1264_.vdd
rlabel metal2 4433 133 4447 147 0 _1264_.A
rlabel metal2 4413 113 4427 127 0 _1264_.B
rlabel metal2 4393 133 4407 147 0 _1264_.C
rlabel metal2 4373 113 4387 127 0 _1264_.Y
rlabel metal1 4524 242 4636 258 0 _1263_.gnd
rlabel metal1 4524 2 4636 18 0 _1263_.vdd
rlabel metal2 4533 133 4547 147 0 _1263_.A
rlabel metal2 4553 113 4567 127 0 _1263_.B
rlabel metal2 4573 133 4587 147 0 _1263_.C
rlabel metal2 4593 113 4607 127 0 _1263_.Y
rlabel nsubstratencontact 4756 488 4756 488 0 FILL71250x3750.vdd
rlabel metal1 4744 242 4776 258 0 FILL71250x3750.gnd
rlabel nsubstratencontact 4764 12 4764 12 0 FILL71250x150.vdd
rlabel metal1 4744 242 4776 258 0 FILL71250x150.gnd
rlabel nsubstratencontact 4744 12 4744 12 0 FILL70950x150.vdd
rlabel metal1 4724 242 4756 258 0 FILL70950x150.gnd
rlabel metal1 4624 242 4736 258 0 _1140_.gnd
rlabel metal1 4624 2 4736 18 0 _1140_.vdd
rlabel metal2 4713 133 4727 147 0 _1140_.A
rlabel metal2 4693 173 4707 187 0 _1140_.B
rlabel metal2 4673 133 4687 147 0 _1140_.C
rlabel metal2 4653 153 4667 167 0 _1140_.Y
rlabel metal1 4624 242 4696 258 0 _1262_.gnd
rlabel metal1 4624 482 4696 498 0 _1262_.vdd
rlabel metal2 4633 313 4647 327 0 _1262_.A
rlabel metal2 4653 353 4667 367 0 _1262_.Y
rlabel metal1 4564 242 4636 258 0 _1260_.gnd
rlabel metal1 4564 482 4636 498 0 _1260_.vdd
rlabel metal2 4573 313 4587 327 0 _1260_.A
rlabel metal2 4593 353 4607 367 0 _1260_.Y
rlabel metal1 4684 242 4756 258 0 _1224_.gnd
rlabel metal1 4684 482 4756 498 0 _1224_.vdd
rlabel metal2 4693 313 4707 327 0 _1224_.A
rlabel metal2 4713 353 4727 367 0 _1224_.Y
rlabel metal1 4 722 256 738 0 _1574_.gnd
rlabel metal1 4 482 256 498 0 _1574_.vdd
rlabel metal2 93 633 107 647 0 _1574_.D
rlabel metal2 133 633 147 647 0 _1574_.CLK
rlabel metal2 213 633 227 647 0 _1574_.Q
rlabel metal1 244 722 316 738 0 _1454_.gnd
rlabel metal1 244 482 316 498 0 _1454_.vdd
rlabel metal2 253 653 267 667 0 _1454_.A
rlabel metal2 273 613 287 627 0 _1454_.Y
rlabel metal1 484 722 576 738 0 BUFX2_insert17.gnd
rlabel metal1 484 482 576 498 0 BUFX2_insert17.vdd
rlabel metal2 493 633 507 647 0 BUFX2_insert17.A
rlabel metal2 533 633 547 647 0 BUFX2_insert17.Y
rlabel metal1 304 722 416 738 0 _771_.gnd
rlabel metal1 304 482 416 498 0 _771_.vdd
rlabel metal2 313 633 327 647 0 _771_.A
rlabel metal2 333 613 347 627 0 _771_.B
rlabel metal2 373 613 387 627 0 _771_.C
rlabel metal2 353 633 367 647 0 _771_.Y
rlabel metal1 404 722 496 738 0 _770_.gnd
rlabel metal1 404 482 496 498 0 _770_.vdd
rlabel metal2 413 593 427 607 0 _770_.A
rlabel metal2 453 593 467 607 0 _770_.B
rlabel metal2 433 613 447 627 0 _770_.Y
rlabel metal1 624 722 876 738 0 _1569_.gnd
rlabel metal1 624 482 876 498 0 _1569_.vdd
rlabel metal2 773 633 787 647 0 _1569_.D
rlabel metal2 733 633 747 647 0 _1569_.CLK
rlabel metal2 653 633 667 647 0 _1569_.Q
rlabel metal1 564 722 636 738 0 _769_.gnd
rlabel metal1 564 482 636 498 0 _769_.vdd
rlabel metal2 613 653 627 667 0 _769_.A
rlabel metal2 593 613 607 627 0 _769_.Y
rlabel metal1 864 722 976 738 0 _1415_.gnd
rlabel metal1 864 482 976 498 0 _1415_.vdd
rlabel metal2 873 633 887 647 0 _1415_.A
rlabel metal2 893 613 907 627 0 _1415_.B
rlabel metal2 933 613 947 627 0 _1415_.C
rlabel metal2 913 633 927 647 0 _1415_.Y
rlabel metal1 964 722 1056 738 0 _1450_.gnd
rlabel metal1 964 482 1056 498 0 _1450_.vdd
rlabel metal2 993 633 1007 647 0 _1450_.B
rlabel metal2 1033 633 1047 647 0 _1450_.A
rlabel metal2 1013 653 1027 667 0 _1450_.Y
rlabel metal1 1044 722 1156 738 0 _1445_.gnd
rlabel metal1 1044 482 1156 498 0 _1445_.vdd
rlabel metal2 1053 653 1067 667 0 _1445_.A
rlabel metal2 1073 633 1087 647 0 _1445_.B
rlabel metal2 1113 613 1127 627 0 _1445_.Y
rlabel metal1 1144 722 1256 738 0 _1414_.gnd
rlabel metal1 1144 482 1256 498 0 _1414_.vdd
rlabel metal2 1233 633 1247 647 0 _1414_.A
rlabel metal2 1213 613 1227 627 0 _1414_.B
rlabel metal2 1173 613 1187 627 0 _1414_.C
rlabel metal2 1193 633 1207 647 0 _1414_.Y
rlabel metal1 1244 722 1356 738 0 _1412_.gnd
rlabel metal1 1244 482 1356 498 0 _1412_.vdd
rlabel metal2 1333 633 1347 647 0 _1412_.A
rlabel metal2 1273 633 1287 647 0 _1412_.Y
rlabel metal2 1293 593 1307 607 0 _1412_.B
rlabel metal1 1424 722 1516 738 0 BUFX2_insert20.gnd
rlabel metal1 1424 482 1516 498 0 BUFX2_insert20.vdd
rlabel metal2 1433 633 1447 647 0 BUFX2_insert20.A
rlabel metal2 1473 633 1487 647 0 BUFX2_insert20.Y
rlabel metal1 1504 722 1756 738 0 _1576_.gnd
rlabel metal1 1504 482 1756 498 0 _1576_.vdd
rlabel metal2 1593 633 1607 647 0 _1576_.D
rlabel metal2 1633 633 1647 647 0 _1576_.CLK
rlabel metal2 1713 633 1727 647 0 _1576_.Q
rlabel metal1 1344 722 1436 738 0 _1413_.gnd
rlabel metal1 1344 482 1436 498 0 _1413_.vdd
rlabel metal2 1393 633 1407 647 0 _1413_.B
rlabel metal2 1353 633 1367 647 0 _1413_.A
rlabel metal2 1373 653 1387 667 0 _1413_.Y
rlabel metal1 1744 722 1836 738 0 BUFX2_insert7.gnd
rlabel metal1 1744 482 1836 498 0 BUFX2_insert7.vdd
rlabel metal2 1753 633 1767 647 0 BUFX2_insert7.A
rlabel metal2 1793 633 1807 647 0 BUFX2_insert7.Y
rlabel metal1 1824 722 1916 738 0 _1411_.gnd
rlabel metal1 1824 482 1916 498 0 _1411_.vdd
rlabel metal2 1853 633 1867 647 0 _1411_.B
rlabel metal2 1893 633 1907 647 0 _1411_.A
rlabel metal2 1873 653 1887 667 0 _1411_.Y
rlabel metal1 2124 722 2376 738 0 _1539_.gnd
rlabel metal1 2124 482 2376 498 0 _1539_.vdd
rlabel metal2 2273 633 2287 647 0 _1539_.D
rlabel metal2 2233 633 2247 647 0 _1539_.CLK
rlabel metal2 2153 633 2167 647 0 _1539_.Q
rlabel metal1 1904 722 1996 738 0 _1410_.gnd
rlabel metal1 1904 482 1996 498 0 _1410_.vdd
rlabel metal2 1933 633 1947 647 0 _1410_.B
rlabel metal2 1973 633 1987 647 0 _1410_.A
rlabel metal2 1953 653 1967 667 0 _1410_.Y
rlabel metal1 2044 722 2136 738 0 _1409_.gnd
rlabel metal1 2044 482 2136 498 0 _1409_.vdd
rlabel metal2 2093 633 2107 647 0 _1409_.B
rlabel metal2 2053 633 2067 647 0 _1409_.A
rlabel metal2 2073 653 2087 667 0 _1409_.Y
rlabel metal1 1984 722 2056 738 0 _830_.gnd
rlabel metal1 1984 482 2056 498 0 _830_.vdd
rlabel metal2 2033 653 2047 667 0 _830_.A
rlabel metal2 2013 613 2027 627 0 _830_.Y
rlabel metal1 2364 722 2496 738 0 _1237_.gnd
rlabel metal1 2364 482 2496 498 0 _1237_.vdd
rlabel metal2 2373 633 2387 647 0 _1237_.A
rlabel metal2 2393 613 2407 627 0 _1237_.B
rlabel metal2 2453 633 2467 647 0 _1237_.C
rlabel metal2 2433 613 2447 627 0 _1237_.D
rlabel metal2 2413 633 2427 647 0 _1237_.Y
rlabel metal1 2584 722 2696 738 0 _1236_.gnd
rlabel metal1 2584 482 2696 498 0 _1236_.vdd
rlabel metal2 2673 613 2687 627 0 _1236_.A
rlabel metal2 2653 653 2667 667 0 _1236_.B
rlabel metal2 2633 613 2647 627 0 _1236_.C
rlabel metal2 2613 633 2627 647 0 _1236_.Y
rlabel metal1 2484 722 2596 738 0 _1235_.gnd
rlabel metal1 2484 482 2596 498 0 _1235_.vdd
rlabel metal2 2573 653 2587 667 0 _1235_.A
rlabel metal2 2553 633 2567 647 0 _1235_.B
rlabel metal2 2513 613 2527 627 0 _1235_.Y
rlabel metal1 2844 722 2956 738 0 _1315_.gnd
rlabel metal1 2844 482 2956 498 0 _1315_.vdd
rlabel metal2 2933 633 2947 647 0 _1315_.A
rlabel metal2 2913 613 2927 627 0 _1315_.B
rlabel metal2 2873 613 2887 627 0 _1315_.C
rlabel metal2 2893 633 2907 647 0 _1315_.Y
rlabel metal1 2684 722 2796 738 0 _1199_.gnd
rlabel metal1 2684 482 2796 498 0 _1199_.vdd
rlabel metal2 2773 613 2787 627 0 _1199_.A
rlabel metal2 2753 653 2767 667 0 _1199_.B
rlabel metal2 2733 613 2747 627 0 _1199_.C
rlabel metal2 2713 633 2727 647 0 _1199_.Y
rlabel metal1 2784 722 2856 738 0 _1305_.gnd
rlabel metal1 2784 482 2856 498 0 _1305_.vdd
rlabel metal2 2793 653 2807 667 0 _1305_.A
rlabel metal2 2813 613 2827 627 0 _1305_.Y
rlabel metal1 2944 722 3056 738 0 _1306_.gnd
rlabel metal1 2944 482 3056 498 0 _1306_.vdd
rlabel metal2 2953 633 2967 647 0 _1306_.A
rlabel metal2 2973 613 2987 627 0 _1306_.B
rlabel metal2 3013 613 3027 627 0 _1306_.C
rlabel metal2 2993 633 3007 647 0 _1306_.Y
rlabel metal1 3044 722 3136 738 0 _1307_.gnd
rlabel metal1 3044 482 3136 498 0 _1307_.vdd
rlabel metal2 3053 593 3067 607 0 _1307_.A
rlabel metal2 3093 593 3107 607 0 _1307_.B
rlabel metal2 3073 613 3087 627 0 _1307_.Y
rlabel metal1 3184 722 3256 738 0 _1208_.gnd
rlabel metal1 3184 482 3256 498 0 _1208_.vdd
rlabel metal2 3193 653 3207 667 0 _1208_.A
rlabel metal2 3213 613 3227 627 0 _1208_.Y
rlabel metal1 3124 722 3196 738 0 _1198_.gnd
rlabel metal1 3124 482 3196 498 0 _1198_.vdd
rlabel metal2 3173 653 3187 667 0 _1198_.A
rlabel metal2 3153 613 3167 627 0 _1198_.Y
rlabel metal1 3424 722 3536 738 0 _1244_.gnd
rlabel metal1 3424 482 3536 498 0 _1244_.vdd
rlabel metal2 3433 633 3447 647 0 _1244_.A
rlabel metal2 3453 613 3467 627 0 _1244_.B
rlabel metal2 3493 613 3507 627 0 _1244_.C
rlabel metal2 3473 633 3487 647 0 _1244_.Y
rlabel metal1 3344 722 3436 738 0 _1234_.gnd
rlabel metal1 3344 482 3436 498 0 _1234_.vdd
rlabel metal2 3373 633 3387 647 0 _1234_.B
rlabel metal2 3413 633 3427 647 0 _1234_.A
rlabel metal2 3393 653 3407 667 0 _1234_.Y
rlabel metal1 3244 722 3356 738 0 _1270_.gnd
rlabel metal1 3244 482 3356 498 0 _1270_.vdd
rlabel metal2 3333 613 3347 627 0 _1270_.A
rlabel metal2 3313 593 3327 607 0 _1270_.B
rlabel metal2 3293 613 3307 627 0 _1270_.C
rlabel metal2 3273 593 3287 607 0 _1270_.Y
rlabel metal1 3524 722 3636 738 0 _1245_.gnd
rlabel metal1 3524 482 3636 498 0 _1245_.vdd
rlabel metal2 3533 613 3547 627 0 _1245_.A
rlabel metal2 3553 653 3567 667 0 _1245_.B
rlabel metal2 3573 613 3587 627 0 _1245_.C
rlabel metal2 3593 633 3607 647 0 _1245_.Y
rlabel metal1 3624 722 3736 738 0 _1230_.gnd
rlabel metal1 3624 482 3736 498 0 _1230_.vdd
rlabel metal2 3713 613 3727 627 0 _1230_.A
rlabel metal2 3693 653 3707 667 0 _1230_.B
rlabel metal2 3673 613 3687 627 0 _1230_.C
rlabel metal2 3653 633 3667 647 0 _1230_.Y
rlabel metal1 3724 722 3856 738 0 _1233_.gnd
rlabel metal1 3724 482 3856 498 0 _1233_.vdd
rlabel metal2 3833 633 3847 647 0 _1233_.A
rlabel metal2 3813 613 3827 627 0 _1233_.B
rlabel metal2 3753 633 3767 647 0 _1233_.C
rlabel metal2 3773 613 3787 627 0 _1233_.D
rlabel metal2 3793 633 3807 647 0 _1233_.Y
rlabel metal1 3844 722 3956 738 0 _1232_.gnd
rlabel metal1 3844 482 3956 498 0 _1232_.vdd
rlabel metal2 3933 613 3947 627 0 _1232_.A
rlabel metal2 3913 593 3927 607 0 _1232_.B
rlabel metal2 3893 613 3907 627 0 _1232_.C
rlabel metal2 3873 593 3887 607 0 _1232_.Y
rlabel metal1 3944 722 4056 738 0 _1226_.gnd
rlabel metal1 3944 482 4056 498 0 _1226_.vdd
rlabel metal2 4033 613 4047 627 0 _1226_.A
rlabel metal2 4013 593 4027 607 0 _1226_.B
rlabel metal2 3993 613 4007 627 0 _1226_.C
rlabel metal2 3973 593 3987 607 0 _1226_.Y
rlabel metal1 4044 722 4116 738 0 _1203_.gnd
rlabel metal1 4044 482 4116 498 0 _1203_.vdd
rlabel metal2 4053 653 4067 667 0 _1203_.A
rlabel metal2 4073 613 4087 627 0 _1203_.Y
rlabel metal1 4104 722 4216 738 0 _1231_.gnd
rlabel metal1 4104 482 4216 498 0 _1231_.vdd
rlabel metal2 4113 613 4127 627 0 _1231_.A
rlabel metal2 4133 593 4147 607 0 _1231_.B
rlabel metal2 4153 613 4167 627 0 _1231_.C
rlabel metal2 4173 593 4187 607 0 _1231_.Y
rlabel metal1 4204 722 4316 738 0 _1229_.gnd
rlabel metal1 4204 482 4316 498 0 _1229_.vdd
rlabel metal2 4213 613 4227 627 0 _1229_.A
rlabel metal2 4233 593 4247 607 0 _1229_.B
rlabel metal2 4253 613 4267 627 0 _1229_.C
rlabel metal2 4273 593 4287 607 0 _1229_.Y
rlabel metal1 4504 722 4576 738 0 _1144_.gnd
rlabel metal1 4504 482 4576 498 0 _1144_.vdd
rlabel metal2 4513 653 4527 667 0 _1144_.A
rlabel metal2 4533 613 4547 627 0 _1144_.Y
rlabel metal1 4304 722 4416 738 0 _1227_.gnd
rlabel metal1 4304 482 4416 498 0 _1227_.vdd
rlabel metal2 4393 613 4407 627 0 _1227_.A
rlabel metal2 4373 593 4387 607 0 _1227_.B
rlabel metal2 4353 613 4367 627 0 _1227_.C
rlabel metal2 4333 593 4347 607 0 _1227_.Y
rlabel metal1 4404 722 4516 738 0 _1220_.gnd
rlabel metal1 4404 482 4516 498 0 _1220_.vdd
rlabel metal2 4493 613 4507 627 0 _1220_.A
rlabel metal2 4473 593 4487 607 0 _1220_.B
rlabel metal2 4453 613 4467 627 0 _1220_.C
rlabel metal2 4433 593 4447 607 0 _1220_.Y
rlabel metal1 4664 722 4776 738 0 _1228_.gnd
rlabel metal1 4664 482 4776 498 0 _1228_.vdd
rlabel metal2 4673 633 4687 647 0 _1228_.A
rlabel metal2 4693 613 4707 627 0 _1228_.B
rlabel metal2 4733 613 4747 627 0 _1228_.C
rlabel metal2 4713 633 4727 647 0 _1228_.Y
rlabel metal1 4564 722 4676 738 0 _1225_.gnd
rlabel metal1 4564 482 4676 498 0 _1225_.vdd
rlabel metal2 4653 633 4667 647 0 _1225_.A
rlabel metal2 4633 613 4647 627 0 _1225_.B
rlabel metal2 4593 613 4607 627 0 _1225_.C
rlabel metal2 4613 633 4627 647 0 _1225_.Y
rlabel metal1 4 722 256 738 0 _1575_.gnd
rlabel metal1 4 962 256 978 0 _1575_.vdd
rlabel metal2 93 813 107 827 0 _1575_.D
rlabel metal2 133 813 147 827 0 _1575_.CLK
rlabel metal2 213 813 227 827 0 _1575_.Q
rlabel metal1 244 722 336 738 0 _1474_.gnd
rlabel metal1 244 962 336 978 0 _1474_.vdd
rlabel metal2 253 853 267 867 0 _1474_.A
rlabel metal2 293 853 307 867 0 _1474_.B
rlabel metal2 273 833 287 847 0 _1474_.Y
rlabel metal1 424 722 676 738 0 _1568_.gnd
rlabel metal1 424 962 676 978 0 _1568_.vdd
rlabel metal2 513 813 527 827 0 _1568_.D
rlabel metal2 553 813 567 827 0 _1568_.CLK
rlabel metal2 633 813 647 827 0 _1568_.Q
rlabel metal1 324 722 436 738 0 _1478_.gnd
rlabel metal1 324 962 436 978 0 _1478_.vdd
rlabel metal2 413 813 427 827 0 _1478_.A
rlabel metal2 393 833 407 847 0 _1478_.B
rlabel metal2 353 833 367 847 0 _1478_.C
rlabel metal2 373 813 387 827 0 _1478_.Y
rlabel metal1 744 722 856 738 0 _1407_.gnd
rlabel metal1 744 962 856 978 0 _1407_.vdd
rlabel metal2 833 813 847 827 0 _1407_.A
rlabel metal2 813 833 827 847 0 _1407_.B
rlabel metal2 773 833 787 847 0 _1407_.C
rlabel metal2 793 813 807 827 0 _1407_.Y
rlabel metal1 664 722 756 738 0 _1393_.gnd
rlabel metal1 664 962 756 978 0 _1393_.vdd
rlabel metal2 673 853 687 867 0 _1393_.A
rlabel metal2 713 853 727 867 0 _1393_.B
rlabel metal2 693 833 707 847 0 _1393_.Y
rlabel metal1 844 722 956 738 0 _1406_.gnd
rlabel metal1 844 962 956 978 0 _1406_.vdd
rlabel metal2 933 813 947 827 0 _1406_.A
rlabel metal2 913 833 927 847 0 _1406_.B
rlabel metal2 873 833 887 847 0 _1406_.C
rlabel metal2 893 813 907 827 0 _1406_.Y
rlabel metal1 1004 722 1096 738 0 _1444_.gnd
rlabel metal1 1004 962 1096 978 0 _1444_.vdd
rlabel metal2 1033 813 1047 827 0 _1444_.B
rlabel metal2 1073 813 1087 827 0 _1444_.A
rlabel metal2 1053 793 1067 807 0 _1444_.Y
rlabel metal1 944 722 1016 738 0 _1405_.gnd
rlabel metal1 944 962 1016 978 0 _1405_.vdd
rlabel metal2 993 793 1007 807 0 _1405_.A
rlabel metal2 973 833 987 847 0 _1405_.Y
rlabel metal1 1164 722 1256 738 0 _1443_.gnd
rlabel metal1 1164 962 1256 978 0 _1443_.vdd
rlabel metal2 1233 853 1247 867 0 _1443_.A
rlabel metal2 1193 853 1207 867 0 _1443_.B
rlabel metal2 1213 833 1227 847 0 _1443_.Y
rlabel metal1 1244 722 1336 738 0 _1442_.gnd
rlabel metal1 1244 962 1336 978 0 _1442_.vdd
rlabel metal2 1313 853 1327 867 0 _1442_.A
rlabel metal2 1273 853 1287 867 0 _1442_.B
rlabel metal2 1293 833 1307 847 0 _1442_.Y
rlabel metal1 1324 722 1416 738 0 _1441_.gnd
rlabel metal1 1324 962 1416 978 0 _1441_.vdd
rlabel metal2 1393 853 1407 867 0 _1441_.A
rlabel metal2 1353 853 1367 867 0 _1441_.B
rlabel metal2 1373 833 1387 847 0 _1441_.Y
rlabel metal1 1084 722 1176 738 0 _1404_.gnd
rlabel metal1 1084 962 1176 978 0 _1404_.vdd
rlabel metal2 1133 813 1147 827 0 _1404_.B
rlabel metal2 1093 813 1107 827 0 _1404_.A
rlabel metal2 1113 793 1127 807 0 _1404_.Y
rlabel metal1 1404 722 1516 738 0 _1420_.gnd
rlabel metal1 1404 962 1516 978 0 _1420_.vdd
rlabel metal2 1493 833 1507 847 0 _1420_.A
rlabel metal2 1473 793 1487 807 0 _1420_.B
rlabel metal2 1453 833 1467 847 0 _1420_.C
rlabel metal2 1433 813 1447 827 0 _1420_.Y
rlabel metal1 1604 722 1716 738 0 _1408_.gnd
rlabel metal1 1604 962 1716 978 0 _1408_.vdd
rlabel metal2 1613 833 1627 847 0 _1408_.A
rlabel metal2 1633 793 1647 807 0 _1408_.B
rlabel metal2 1653 833 1667 847 0 _1408_.C
rlabel metal2 1673 813 1687 827 0 _1408_.Y
rlabel metal1 1504 722 1616 738 0 _1417_.gnd
rlabel metal1 1504 962 1616 978 0 _1417_.vdd
rlabel metal2 1593 813 1607 827 0 _1417_.A
rlabel metal2 1533 813 1547 827 0 _1417_.Y
rlabel metal2 1553 853 1567 867 0 _1417_.B
rlabel metal1 1704 722 1916 738 0 CLKBUF1_insert15.gnd
rlabel metal1 1704 962 1916 978 0 CLKBUF1_insert15.vdd
rlabel metal2 1733 833 1747 847 0 CLKBUF1_insert15.A
rlabel metal2 1873 833 1887 847 0 CLKBUF1_insert15.Y
rlabel metal1 2064 722 2176 738 0 _1419_.gnd
rlabel metal1 2064 962 2176 978 0 _1419_.vdd
rlabel metal2 2073 813 2087 827 0 _1419_.A
rlabel metal2 2093 833 2107 847 0 _1419_.B
rlabel metal2 2133 833 2147 847 0 _1419_.C
rlabel metal2 2113 813 2127 827 0 _1419_.Y
rlabel metal1 1904 722 1996 738 0 _843_.gnd
rlabel metal1 1904 962 1996 978 0 _843_.vdd
rlabel metal2 1973 853 1987 867 0 _843_.A
rlabel metal2 1933 853 1947 867 0 _843_.B
rlabel metal2 1953 833 1967 847 0 _843_.Y
rlabel metal1 1984 722 2076 738 0 _1403_.gnd
rlabel metal1 1984 962 2076 978 0 _1403_.vdd
rlabel metal2 2013 813 2027 827 0 _1403_.B
rlabel metal2 2053 813 2067 827 0 _1403_.A
rlabel metal2 2033 793 2047 807 0 _1403_.Y
rlabel metal1 2164 722 2276 738 0 _1418_.gnd
rlabel metal1 2164 962 2276 978 0 _1418_.vdd
rlabel metal2 2173 813 2187 827 0 _1418_.A
rlabel metal2 2193 833 2207 847 0 _1418_.B
rlabel metal2 2233 833 2247 847 0 _1418_.C
rlabel metal2 2213 813 2227 827 0 _1418_.Y
rlabel metal1 2264 722 2376 738 0 _832_.gnd
rlabel metal1 2264 962 2376 978 0 _832_.vdd
rlabel metal2 2273 813 2287 827 0 _832_.A
rlabel metal2 2293 833 2307 847 0 _832_.B
rlabel metal2 2333 833 2347 847 0 _832_.C
rlabel metal2 2313 813 2327 827 0 _832_.Y
rlabel metal1 2364 722 2456 738 0 _831_.gnd
rlabel metal1 2364 962 2456 978 0 _831_.vdd
rlabel metal2 2373 853 2387 867 0 _831_.A
rlabel metal2 2413 853 2427 867 0 _831_.B
rlabel metal2 2393 833 2407 847 0 _831_.Y
rlabel metal1 2504 722 2756 738 0 _1555_.gnd
rlabel metal1 2504 962 2756 978 0 _1555_.vdd
rlabel metal2 2653 813 2667 827 0 _1555_.D
rlabel metal2 2613 813 2627 827 0 _1555_.CLK
rlabel metal2 2533 813 2547 827 0 _1555_.Q
rlabel metal1 2444 722 2516 738 0 _1196_.gnd
rlabel metal1 2444 962 2516 978 0 _1196_.vdd
rlabel metal2 2493 793 2507 807 0 _1196_.A
rlabel metal2 2473 833 2487 847 0 _1196_.Y
rlabel metal1 2744 722 2856 738 0 _1194_.gnd
rlabel metal1 2744 962 2856 978 0 _1194_.vdd
rlabel metal2 2833 813 2847 827 0 _1194_.A
rlabel metal2 2813 833 2827 847 0 _1194_.B
rlabel metal2 2773 833 2787 847 0 _1194_.C
rlabel metal2 2793 813 2807 827 0 _1194_.Y
rlabel metal1 2904 722 2976 738 0 _1193_.gnd
rlabel metal1 2904 962 2976 978 0 _1193_.vdd
rlabel metal2 2913 793 2927 807 0 _1193_.A
rlabel metal2 2933 833 2947 847 0 _1193_.Y
rlabel metal1 2844 722 2916 738 0 _1191_.gnd
rlabel metal1 2844 962 2916 978 0 _1191_.vdd
rlabel metal2 2893 793 2907 807 0 _1191_.A
rlabel metal2 2873 833 2887 847 0 _1191_.Y
rlabel metal1 3124 722 3216 738 0 _1284_.gnd
rlabel metal1 3124 962 3216 978 0 _1284_.vdd
rlabel metal2 3193 853 3207 867 0 _1284_.A
rlabel metal2 3153 853 3167 867 0 _1284_.B
rlabel metal2 3173 833 3187 847 0 _1284_.Y
rlabel metal1 3064 722 3136 738 0 _1303_.gnd
rlabel metal1 3064 962 3136 978 0 _1303_.vdd
rlabel metal2 3073 793 3087 807 0 _1303_.A
rlabel metal2 3093 833 3107 847 0 _1303_.Y
rlabel metal1 2964 722 3076 738 0 _1304_.gnd
rlabel metal1 2964 962 3076 978 0 _1304_.vdd
rlabel metal2 2973 833 2987 847 0 _1304_.A
rlabel metal2 2993 853 3007 867 0 _1304_.B
rlabel metal2 3013 833 3027 847 0 _1304_.C
rlabel metal2 3033 853 3047 867 0 _1304_.Y
rlabel metal1 3204 722 3316 738 0 _1283_.gnd
rlabel metal1 3204 962 3316 978 0 _1283_.vdd
rlabel metal2 3213 793 3227 807 0 _1283_.A
rlabel metal2 3233 813 3247 827 0 _1283_.B
rlabel metal2 3273 833 3287 847 0 _1283_.Y
rlabel metal1 3304 722 3396 738 0 _1285_.gnd
rlabel metal1 3304 962 3396 978 0 _1285_.vdd
rlabel metal2 3313 853 3327 867 0 _1285_.A
rlabel metal2 3353 853 3367 867 0 _1285_.B
rlabel metal2 3333 833 3347 847 0 _1285_.Y
rlabel metal1 3384 722 3476 738 0 _1190_.gnd
rlabel metal1 3384 962 3476 978 0 _1190_.vdd
rlabel metal2 3393 853 3407 867 0 _1190_.A
rlabel metal2 3433 853 3447 867 0 _1190_.B
rlabel metal2 3413 833 3427 847 0 _1190_.Y
rlabel metal1 3464 722 3556 738 0 _1243_.gnd
rlabel metal1 3464 962 3556 978 0 _1243_.vdd
rlabel metal2 3493 813 3507 827 0 _1243_.B
rlabel metal2 3533 813 3547 827 0 _1243_.A
rlabel metal2 3513 793 3527 807 0 _1243_.Y
rlabel metal1 3544 722 3636 738 0 _1242_.gnd
rlabel metal1 3544 962 3636 978 0 _1242_.vdd
rlabel metal2 3553 853 3567 867 0 _1242_.A
rlabel metal2 3593 853 3607 867 0 _1242_.B
rlabel metal2 3573 833 3587 847 0 _1242_.Y
rlabel metal1 3624 722 3736 738 0 _1241_.gnd
rlabel metal1 3624 962 3736 978 0 _1241_.vdd
rlabel metal2 3713 833 3727 847 0 _1241_.A
rlabel metal2 3693 853 3707 867 0 _1241_.B
rlabel metal2 3673 833 3687 847 0 _1241_.C
rlabel metal2 3653 853 3667 867 0 _1241_.Y
rlabel metal1 3724 722 3836 738 0 _1240_.gnd
rlabel metal1 3724 962 3836 978 0 _1240_.vdd
rlabel metal2 3813 833 3827 847 0 _1240_.A
rlabel metal2 3793 853 3807 867 0 _1240_.B
rlabel metal2 3773 833 3787 847 0 _1240_.C
rlabel metal2 3753 853 3767 867 0 _1240_.Y
rlabel metal1 3824 722 3916 738 0 _1239_.gnd
rlabel metal1 3824 962 3916 978 0 _1239_.vdd
rlabel metal2 3833 853 3847 867 0 _1239_.A
rlabel metal2 3873 853 3887 867 0 _1239_.B
rlabel metal2 3853 833 3867 847 0 _1239_.Y
rlabel metal1 4004 722 4076 738 0 _1186_.gnd
rlabel metal1 4004 962 4076 978 0 _1186_.vdd
rlabel metal2 4053 793 4067 807 0 _1186_.A
rlabel metal2 4033 833 4047 847 0 _1186_.Y
rlabel metal1 3904 722 4016 738 0 _1185_.gnd
rlabel metal1 3904 962 4016 978 0 _1185_.vdd
rlabel metal2 3993 833 4007 847 0 _1185_.A
rlabel metal2 3973 853 3987 867 0 _1185_.B
rlabel metal2 3953 833 3967 847 0 _1185_.C
rlabel metal2 3933 853 3947 867 0 _1185_.Y
rlabel metal1 4164 722 4276 738 0 _1201_.gnd
rlabel metal1 4164 962 4276 978 0 _1201_.vdd
rlabel metal2 4253 813 4267 827 0 _1201_.A
rlabel metal2 4233 833 4247 847 0 _1201_.B
rlabel metal2 4193 833 4207 847 0 _1201_.C
rlabel metal2 4213 813 4227 827 0 _1201_.Y
rlabel metal1 4064 722 4176 738 0 _1189_.gnd
rlabel metal1 4064 962 4176 978 0 _1189_.vdd
rlabel metal2 4153 813 4167 827 0 _1189_.A
rlabel metal2 4133 833 4147 847 0 _1189_.B
rlabel metal2 4093 833 4107 847 0 _1189_.C
rlabel metal2 4113 813 4127 827 0 _1189_.Y
rlabel metal1 4264 722 4376 738 0 _1188_.gnd
rlabel metal1 4264 962 4376 978 0 _1188_.vdd
rlabel metal2 4353 833 4367 847 0 _1188_.A
rlabel metal2 4333 793 4347 807 0 _1188_.B
rlabel metal2 4313 833 4327 847 0 _1188_.C
rlabel metal2 4293 813 4307 827 0 _1188_.Y
rlabel metal1 4364 722 4476 738 0 _1181_.gnd
rlabel metal1 4364 962 4476 978 0 _1181_.vdd
rlabel metal2 4373 833 4387 847 0 _1181_.A
rlabel metal2 4393 853 4407 867 0 _1181_.B
rlabel metal2 4413 833 4427 847 0 _1181_.C
rlabel metal2 4433 853 4447 867 0 _1181_.Y
rlabel metal1 4464 722 4576 738 0 _1175_.gnd
rlabel metal1 4464 962 4576 978 0 _1175_.vdd
rlabel metal2 4553 833 4567 847 0 _1175_.A
rlabel metal2 4533 853 4547 867 0 _1175_.B
rlabel metal2 4513 833 4527 847 0 _1175_.C
rlabel metal2 4493 853 4507 867 0 _1175_.Y
rlabel metal1 4564 722 4676 738 0 _1200_.gnd
rlabel metal1 4564 962 4676 978 0 _1200_.vdd
rlabel metal2 4653 833 4667 847 0 _1200_.A
rlabel metal2 4633 793 4647 807 0 _1200_.B
rlabel metal2 4613 833 4627 847 0 _1200_.C
rlabel metal2 4593 813 4607 827 0 _1200_.Y
rlabel metal1 4664 722 4776 738 0 _1182_.gnd
rlabel metal1 4664 962 4776 978 0 _1182_.vdd
rlabel metal2 4673 833 4687 847 0 _1182_.A
rlabel metal2 4693 853 4707 867 0 _1182_.B
rlabel metal2 4713 833 4727 847 0 _1182_.C
rlabel metal2 4733 853 4747 867 0 _1182_.Y
rlabel metal1 144 1202 256 1218 0 _780_.gnd
rlabel metal1 144 962 256 978 0 _780_.vdd
rlabel metal2 233 1113 247 1127 0 _780_.A
rlabel metal2 213 1093 227 1107 0 _780_.B
rlabel metal2 173 1093 187 1107 0 _780_.C
rlabel metal2 193 1113 207 1127 0 _780_.Y
rlabel metal1 64 1202 156 1218 0 _779_.gnd
rlabel metal1 64 962 156 978 0 _779_.vdd
rlabel metal2 133 1073 147 1087 0 _779_.A
rlabel metal2 93 1073 107 1087 0 _779_.B
rlabel metal2 113 1093 127 1107 0 _779_.Y
rlabel metal1 4 1202 76 1218 0 _778_.gnd
rlabel metal1 4 962 76 978 0 _778_.vdd
rlabel metal2 13 1133 27 1147 0 _778_.A
rlabel metal2 33 1093 47 1107 0 _778_.Y
rlabel metal1 244 1202 376 1218 0 _1437_.gnd
rlabel metal1 244 962 376 978 0 _1437_.vdd
rlabel metal2 253 1113 267 1127 0 _1437_.A
rlabel metal2 273 1093 287 1107 0 _1437_.B
rlabel metal2 333 1113 347 1127 0 _1437_.C
rlabel metal2 313 1093 327 1107 0 _1437_.D
rlabel metal2 293 1113 307 1127 0 _1437_.Y
rlabel metal1 364 1202 476 1218 0 _1436_.gnd
rlabel metal1 364 962 476 978 0 _1436_.vdd
rlabel metal2 453 1093 467 1107 0 _1436_.A
rlabel metal2 433 1133 447 1147 0 _1436_.B
rlabel metal2 413 1093 427 1107 0 _1436_.C
rlabel metal2 393 1113 407 1127 0 _1436_.Y
rlabel metal1 464 1202 576 1218 0 _1435_.gnd
rlabel metal1 464 962 576 978 0 _1435_.vdd
rlabel metal2 553 1133 567 1147 0 _1435_.A
rlabel metal2 533 1113 547 1127 0 _1435_.B
rlabel metal2 493 1093 507 1107 0 _1435_.Y
rlabel metal1 744 1202 836 1218 0 BUFX2_insert4.gnd
rlabel metal1 744 962 836 978 0 BUFX2_insert4.vdd
rlabel metal2 813 1113 827 1127 0 BUFX2_insert4.A
rlabel metal2 773 1113 787 1127 0 BUFX2_insert4.Y
rlabel metal1 564 1202 656 1218 0 _760_.gnd
rlabel metal1 564 962 656 978 0 _760_.vdd
rlabel metal2 613 1113 627 1127 0 _760_.B
rlabel metal2 573 1113 587 1127 0 _760_.A
rlabel metal2 593 1133 607 1147 0 _760_.Y
rlabel metal1 644 1202 756 1218 0 _1425_.gnd
rlabel metal1 644 962 756 978 0 _1425_.vdd
rlabel metal2 733 1113 747 1127 0 _1425_.A
rlabel metal2 673 1113 687 1127 0 _1425_.Y
rlabel metal2 693 1073 707 1087 0 _1425_.B
rlabel metal1 824 1202 916 1218 0 _1440_.gnd
rlabel metal1 824 962 916 978 0 _1440_.vdd
rlabel metal2 853 1113 867 1127 0 _1440_.B
rlabel metal2 893 1113 907 1127 0 _1440_.A
rlabel metal2 873 1133 887 1147 0 _1440_.Y
rlabel metal1 1024 1202 1116 1218 0 _1423_.gnd
rlabel metal1 1024 962 1116 978 0 _1423_.vdd
rlabel metal2 1073 1113 1087 1127 0 _1423_.B
rlabel metal2 1033 1113 1047 1127 0 _1423_.A
rlabel metal2 1053 1133 1067 1147 0 _1423_.Y
rlabel metal1 964 1202 1036 1218 0 _1434_.gnd
rlabel metal1 964 962 1036 978 0 _1434_.vdd
rlabel metal2 1013 1133 1027 1147 0 _1434_.A
rlabel metal2 993 1093 1007 1107 0 _1434_.Y
rlabel metal1 904 1202 976 1218 0 _1424_.gnd
rlabel metal1 904 962 976 978 0 _1424_.vdd
rlabel metal2 953 1133 967 1147 0 _1424_.A
rlabel metal2 933 1093 947 1107 0 _1424_.Y
rlabel metal1 1244 1202 1356 1218 0 _1439_.gnd
rlabel metal1 1244 962 1356 978 0 _1439_.vdd
rlabel metal2 1253 1093 1267 1107 0 _1439_.A
rlabel metal2 1273 1133 1287 1147 0 _1439_.B
rlabel metal2 1293 1093 1307 1107 0 _1439_.C
rlabel metal2 1313 1113 1327 1127 0 _1439_.Y
rlabel metal1 1164 1202 1256 1218 0 _1433_.gnd
rlabel metal1 1164 962 1256 978 0 _1433_.vdd
rlabel metal2 1193 1113 1207 1127 0 _1433_.B
rlabel metal2 1233 1113 1247 1127 0 _1433_.A
rlabel metal2 1213 1133 1227 1147 0 _1433_.Y
rlabel metal1 1104 1202 1176 1218 0 _1400_.gnd
rlabel metal1 1104 962 1176 978 0 _1400_.vdd
rlabel metal2 1113 1133 1127 1147 0 _1400_.A
rlabel metal2 1133 1093 1147 1107 0 _1400_.Y
rlabel metal1 1344 1202 1596 1218 0 _1577_.gnd
rlabel metal1 1344 962 1596 978 0 _1577_.vdd
rlabel metal2 1433 1113 1447 1127 0 _1577_.D
rlabel metal2 1473 1113 1487 1127 0 _1577_.CLK
rlabel metal2 1553 1113 1567 1127 0 _1577_.Q
rlabel metal1 1584 1202 1656 1218 0 _1432_.gnd
rlabel metal1 1584 962 1656 978 0 _1432_.vdd
rlabel metal2 1633 1133 1647 1147 0 _1432_.A
rlabel metal2 1613 1093 1627 1107 0 _1432_.Y
rlabel metal1 1804 1202 2056 1218 0 _1538_.gnd
rlabel metal1 1804 962 2056 978 0 _1538_.vdd
rlabel metal2 1893 1113 1907 1127 0 _1538_.D
rlabel metal2 1933 1113 1947 1127 0 _1538_.CLK
rlabel metal2 2013 1113 2027 1127 0 _1538_.Q
rlabel metal1 1644 1202 1736 1218 0 _1431_.gnd
rlabel metal1 1644 962 1736 978 0 _1431_.vdd
rlabel metal2 1653 1073 1667 1087 0 _1431_.A
rlabel metal2 1693 1073 1707 1087 0 _1431_.B
rlabel metal2 1673 1093 1687 1107 0 _1431_.Y
rlabel metal1 1724 1202 1816 1218 0 _1430_.gnd
rlabel metal1 1724 962 1816 978 0 _1430_.vdd
rlabel metal2 1773 1113 1787 1127 0 _1430_.B
rlabel metal2 1733 1113 1747 1127 0 _1430_.A
rlabel metal2 1753 1133 1767 1147 0 _1430_.Y
rlabel metal1 2104 1202 2196 1218 0 _1401_.gnd
rlabel metal1 2104 962 2196 978 0 _1401_.vdd
rlabel metal2 2153 1113 2167 1127 0 _1401_.B
rlabel metal2 2113 1113 2127 1127 0 _1401_.A
rlabel metal2 2133 1133 2147 1147 0 _1401_.Y
rlabel metal1 2044 1202 2116 1218 0 _827_.gnd
rlabel metal1 2044 962 2116 978 0 _827_.vdd
rlabel metal2 2093 1133 2107 1147 0 _827_.A
rlabel metal2 2073 1093 2087 1107 0 _827_.Y
rlabel metal1 2324 1202 2576 1218 0 _1554_.gnd
rlabel metal1 2324 962 2576 978 0 _1554_.vdd
rlabel metal2 2473 1113 2487 1127 0 _1554_.D
rlabel metal2 2433 1113 2447 1127 0 _1554_.CLK
rlabel metal2 2353 1113 2367 1127 0 _1554_.Q
rlabel metal1 2184 1202 2276 1218 0 _1402_.gnd
rlabel metal1 2184 962 2276 978 0 _1402_.vdd
rlabel metal2 2233 1113 2247 1127 0 _1402_.B
rlabel metal2 2193 1113 2207 1127 0 _1402_.A
rlabel metal2 2213 1133 2227 1147 0 _1402_.Y
rlabel metal1 2264 1202 2336 1218 0 _1136_.gnd
rlabel metal1 2264 962 2336 978 0 _1136_.vdd
rlabel metal2 2313 1133 2327 1147 0 _1136_.A
rlabel metal2 2293 1093 2307 1107 0 _1136_.Y
rlabel metal1 2624 1202 2736 1218 0 _1275_.gnd
rlabel metal1 2624 962 2736 978 0 _1275_.vdd
rlabel metal2 2633 1113 2647 1127 0 _1275_.A
rlabel metal2 2653 1093 2667 1107 0 _1275_.B
rlabel metal2 2693 1093 2707 1107 0 _1275_.C
rlabel metal2 2673 1113 2687 1127 0 _1275_.Y
rlabel metal1 2564 1202 2636 1218 0 _1238_.gnd
rlabel metal1 2564 962 2636 978 0 _1238_.vdd
rlabel metal2 2573 1133 2587 1147 0 _1238_.A
rlabel metal2 2593 1093 2607 1107 0 _1238_.Y
rlabel metal1 2924 1202 3016 1218 0 _1281_.gnd
rlabel metal1 2924 962 3016 978 0 _1281_.vdd
rlabel metal2 2993 1073 3007 1087 0 _1281_.A
rlabel metal2 2953 1073 2967 1087 0 _1281_.B
rlabel metal2 2973 1093 2987 1107 0 _1281_.Y
rlabel metal1 2844 1202 2936 1218 0 _1192_.gnd
rlabel metal1 2844 962 2936 978 0 _1192_.vdd
rlabel metal2 2893 1113 2907 1127 0 _1192_.B
rlabel metal2 2853 1113 2867 1127 0 _1192_.A
rlabel metal2 2873 1133 2887 1147 0 _1192_.Y
rlabel metal1 2724 1202 2856 1218 0 _1195_.gnd
rlabel metal1 2724 962 2856 978 0 _1195_.vdd
rlabel metal2 2733 1113 2747 1127 0 _1195_.A
rlabel metal2 2753 1093 2767 1107 0 _1195_.B
rlabel metal2 2813 1113 2827 1127 0 _1195_.C
rlabel metal2 2773 1113 2787 1127 0 _1195_.Y
rlabel metal2 2793 1093 2807 1107 0 _1195_.D
rlabel metal1 3104 1202 3216 1218 0 _1278_.gnd
rlabel metal1 3104 962 3216 978 0 _1278_.vdd
rlabel metal2 3113 1113 3127 1127 0 _1278_.A
rlabel metal2 3133 1093 3147 1107 0 _1278_.B
rlabel metal2 3173 1093 3187 1107 0 _1278_.C
rlabel metal2 3153 1113 3167 1127 0 _1278_.Y
rlabel metal1 3204 1202 3316 1218 0 _1255_.gnd
rlabel metal1 3204 962 3316 978 0 _1255_.vdd
rlabel metal2 3213 1133 3227 1147 0 _1255_.A
rlabel metal2 3233 1113 3247 1127 0 _1255_.B
rlabel metal2 3273 1093 3287 1107 0 _1255_.Y
rlabel metal1 3004 1202 3116 1218 0 _1282_.gnd
rlabel metal1 3004 962 3116 978 0 _1282_.vdd
rlabel metal2 3013 1113 3027 1127 0 _1282_.A
rlabel metal2 3073 1113 3087 1127 0 _1282_.Y
rlabel metal2 3053 1073 3067 1087 0 _1282_.B
rlabel metal1 3304 1202 3396 1218 0 _1257_.gnd
rlabel metal1 3304 962 3396 978 0 _1257_.vdd
rlabel metal2 3373 1073 3387 1087 0 _1257_.A
rlabel metal2 3333 1073 3347 1087 0 _1257_.B
rlabel metal2 3353 1093 3367 1107 0 _1257_.Y
rlabel metal1 3464 1202 3556 1218 0 _1250_.gnd
rlabel metal1 3464 962 3556 978 0 _1250_.vdd
rlabel metal2 3473 1073 3487 1087 0 _1250_.A
rlabel metal2 3513 1073 3527 1087 0 _1250_.B
rlabel metal2 3493 1093 3507 1107 0 _1250_.Y
rlabel metal1 3384 1202 3476 1218 0 _1209_.gnd
rlabel metal1 3384 962 3476 978 0 _1209_.vdd
rlabel metal2 3453 1073 3467 1087 0 _1209_.A
rlabel metal2 3413 1073 3427 1087 0 _1209_.B
rlabel metal2 3433 1093 3447 1107 0 _1209_.Y
rlabel metal1 3624 1202 3736 1218 0 _1247_.gnd
rlabel metal1 3624 962 3736 978 0 _1247_.vdd
rlabel metal2 3633 1113 3647 1127 0 _1247_.A
rlabel metal2 3653 1093 3667 1107 0 _1247_.B
rlabel metal2 3693 1093 3707 1107 0 _1247_.C
rlabel metal2 3673 1113 3687 1127 0 _1247_.Y
rlabel metal1 3544 1202 3636 1218 0 _1212_.gnd
rlabel metal1 3544 962 3636 978 0 _1212_.vdd
rlabel metal2 3553 1073 3567 1087 0 _1212_.A
rlabel metal2 3593 1073 3607 1087 0 _1212_.B
rlabel metal2 3573 1093 3587 1107 0 _1212_.Y
rlabel metal1 3724 1202 3836 1218 0 _1219_.gnd
rlabel metal1 3724 962 3836 978 0 _1219_.vdd
rlabel metal2 3813 1093 3827 1107 0 _1219_.A
rlabel metal2 3793 1073 3807 1087 0 _1219_.B
rlabel metal2 3773 1093 3787 1107 0 _1219_.C
rlabel metal2 3753 1073 3767 1087 0 _1219_.Y
rlabel metal1 3824 1202 3936 1218 0 _1223_.gnd
rlabel metal1 3824 962 3936 978 0 _1223_.vdd
rlabel metal2 3833 1093 3847 1107 0 _1223_.A
rlabel metal2 3853 1133 3867 1147 0 _1223_.B
rlabel metal2 3873 1093 3887 1107 0 _1223_.C
rlabel metal2 3893 1113 3907 1127 0 _1223_.Y
rlabel metal1 3924 1202 3996 1218 0 _1218_.gnd
rlabel metal1 3924 962 3996 978 0 _1218_.vdd
rlabel metal2 3973 1133 3987 1147 0 _1218_.A
rlabel metal2 3953 1093 3967 1107 0 _1218_.Y
rlabel metal1 3984 1202 4096 1218 0 _1184_.gnd
rlabel metal1 3984 962 4096 978 0 _1184_.vdd
rlabel metal2 4073 1093 4087 1107 0 _1184_.A
rlabel metal2 4053 1073 4067 1087 0 _1184_.B
rlabel metal2 4033 1093 4047 1107 0 _1184_.C
rlabel metal2 4013 1073 4027 1087 0 _1184_.Y
rlabel metal1 4244 1202 4356 1218 0 _1222_.gnd
rlabel metal1 4244 962 4356 978 0 _1222_.vdd
rlabel metal2 4333 1093 4347 1107 0 _1222_.A
rlabel metal2 4313 1133 4327 1147 0 _1222_.B
rlabel metal2 4293 1093 4307 1107 0 _1222_.C
rlabel metal2 4273 1113 4287 1127 0 _1222_.Y
rlabel metal1 4084 1202 4196 1218 0 _1187_.gnd
rlabel metal1 4084 962 4196 978 0 _1187_.vdd
rlabel metal2 4093 1093 4107 1107 0 _1187_.A
rlabel metal2 4113 1133 4127 1147 0 _1187_.B
rlabel metal2 4133 1093 4147 1107 0 _1187_.C
rlabel metal2 4153 1113 4167 1127 0 _1187_.Y
rlabel metal1 4184 1202 4256 1218 0 _1143_.gnd
rlabel metal1 4184 962 4256 978 0 _1143_.vdd
rlabel metal2 4193 1133 4207 1147 0 _1143_.A
rlabel metal2 4213 1093 4227 1107 0 _1143_.Y
rlabel metal1 4344 1202 4456 1218 0 _1183_.gnd
rlabel metal1 4344 962 4456 978 0 _1183_.vdd
rlabel metal2 4433 1113 4447 1127 0 _1183_.A
rlabel metal2 4413 1093 4427 1107 0 _1183_.B
rlabel metal2 4373 1093 4387 1107 0 _1183_.C
rlabel metal2 4393 1113 4407 1127 0 _1183_.Y
rlabel metal1 4444 1202 4556 1218 0 _1180_.gnd
rlabel metal1 4444 962 4556 978 0 _1180_.vdd
rlabel metal2 4453 1113 4467 1127 0 _1180_.A
rlabel metal2 4473 1093 4487 1107 0 _1180_.B
rlabel metal2 4513 1093 4527 1107 0 _1180_.C
rlabel metal2 4493 1113 4507 1127 0 _1180_.Y
rlabel metal1 4624 1202 4716 1218 0 _1174_.gnd
rlabel metal1 4624 962 4716 978 0 _1174_.vdd
rlabel metal2 4693 1073 4707 1087 0 _1174_.A
rlabel metal2 4653 1073 4667 1087 0 _1174_.B
rlabel metal2 4673 1093 4687 1107 0 _1174_.Y
rlabel metal1 4544 1202 4636 1218 0 _1178_.gnd
rlabel metal1 4544 962 4636 978 0 _1178_.vdd
rlabel metal2 4593 1113 4607 1127 0 _1178_.B
rlabel metal2 4553 1113 4567 1127 0 _1178_.A
rlabel metal2 4573 1133 4587 1147 0 _1178_.Y
rlabel metal1 4704 1202 4776 1218 0 _1486_.gnd
rlabel metal1 4704 962 4776 978 0 _1486_.vdd
rlabel metal2 4753 1133 4767 1147 0 _1486_.A
rlabel metal2 4733 1093 4747 1107 0 _1486_.Y
rlabel metal1 4 1202 256 1218 0 _1571_.gnd
rlabel metal1 4 1442 256 1458 0 _1571_.vdd
rlabel metal2 153 1293 167 1307 0 _1571_.D
rlabel metal2 113 1293 127 1307 0 _1571_.CLK
rlabel metal2 33 1293 47 1307 0 _1571_.Q
rlabel metal1 244 1202 496 1218 0 _1570_.gnd
rlabel metal1 244 1442 496 1458 0 _1570_.vdd
rlabel metal2 333 1293 347 1307 0 _1570_.D
rlabel metal2 373 1293 387 1307 0 _1570_.CLK
rlabel metal2 453 1293 467 1307 0 _1570_.Q
rlabel metal1 484 1202 576 1218 0 _1416_.gnd
rlabel metal1 484 1442 576 1458 0 _1416_.vdd
rlabel metal2 493 1333 507 1347 0 _1416_.A
rlabel metal2 533 1333 547 1347 0 _1416_.B
rlabel metal2 513 1313 527 1327 0 _1416_.Y
rlabel metal1 764 1202 856 1218 0 BUFX2_insert0.gnd
rlabel metal1 764 1442 856 1458 0 BUFX2_insert0.vdd
rlabel metal2 833 1293 847 1307 0 BUFX2_insert0.A
rlabel metal2 793 1293 807 1307 0 BUFX2_insert0.Y
rlabel metal1 564 1202 676 1218 0 _1427_.gnd
rlabel metal1 564 1442 676 1458 0 _1427_.vdd
rlabel metal2 653 1293 667 1307 0 _1427_.A
rlabel metal2 633 1313 647 1327 0 _1427_.B
rlabel metal2 593 1313 607 1327 0 _1427_.C
rlabel metal2 613 1293 627 1307 0 _1427_.Y
rlabel metal1 664 1202 776 1218 0 _1426_.gnd
rlabel metal1 664 1442 776 1458 0 _1426_.vdd
rlabel metal2 753 1293 767 1307 0 _1426_.A
rlabel metal2 733 1313 747 1327 0 _1426_.B
rlabel metal2 693 1313 707 1327 0 _1426_.C
rlabel metal2 713 1293 727 1307 0 _1426_.Y
rlabel metal1 924 1202 1036 1218 0 _1429_.gnd
rlabel metal1 924 1442 1036 1458 0 _1429_.vdd
rlabel metal2 1013 1293 1027 1307 0 _1429_.A
rlabel metal2 993 1313 1007 1327 0 _1429_.B
rlabel metal2 953 1313 967 1327 0 _1429_.C
rlabel metal2 973 1293 987 1307 0 _1429_.Y
rlabel metal1 844 1202 936 1218 0 _849_.gnd
rlabel metal1 844 1442 936 1458 0 _849_.vdd
rlabel metal2 853 1333 867 1347 0 _849_.A
rlabel metal2 893 1333 907 1347 0 _849_.B
rlabel metal2 873 1313 887 1327 0 _849_.Y
rlabel metal1 1024 1202 1096 1218 0 _1428_.gnd
rlabel metal1 1024 1442 1096 1458 0 _1428_.vdd
rlabel metal2 1073 1273 1087 1287 0 _1428_.A
rlabel metal2 1053 1313 1067 1327 0 _1428_.Y
rlabel metal1 1284 1202 1396 1218 0 _1485_.gnd
rlabel metal1 1284 1442 1396 1458 0 _1485_.vdd
rlabel metal2 1373 1293 1387 1307 0 _1485_.A
rlabel metal2 1353 1313 1367 1327 0 _1485_.B
rlabel metal2 1313 1313 1327 1327 0 _1485_.C
rlabel metal2 1333 1293 1347 1307 0 _1485_.Y
rlabel metal1 1204 1202 1296 1218 0 _1484_.gnd
rlabel metal1 1204 1442 1296 1458 0 _1484_.vdd
rlabel metal2 1273 1333 1287 1347 0 _1484_.A
rlabel metal2 1233 1333 1247 1347 0 _1484_.B
rlabel metal2 1253 1313 1267 1327 0 _1484_.Y
rlabel metal1 1084 1202 1216 1218 0 _1197_.gnd
rlabel metal1 1084 1442 1216 1458 0 _1197_.vdd
rlabel metal2 1113 1293 1127 1307 0 _1197_.A
rlabel metal2 1153 1293 1167 1307 0 _1197_.Y
rlabel metal1 1564 1202 1656 1218 0 BUFX2_insert6.gnd
rlabel metal1 1564 1442 1656 1458 0 BUFX2_insert6.vdd
rlabel metal2 1573 1293 1587 1307 0 BUFX2_insert6.A
rlabel metal2 1613 1293 1627 1307 0 BUFX2_insert6.Y
rlabel metal1 1464 1202 1576 1218 0 _1482_.gnd
rlabel metal1 1464 1442 1576 1458 0 _1482_.vdd
rlabel metal2 1553 1293 1567 1307 0 _1482_.A
rlabel metal2 1533 1313 1547 1327 0 _1482_.B
rlabel metal2 1493 1313 1507 1327 0 _1482_.C
rlabel metal2 1513 1293 1527 1307 0 _1482_.Y
rlabel metal1 1384 1202 1476 1218 0 _1481_.gnd
rlabel metal1 1384 1442 1476 1458 0 _1481_.vdd
rlabel metal2 1453 1333 1467 1347 0 _1481_.A
rlabel metal2 1413 1333 1427 1347 0 _1481_.B
rlabel metal2 1433 1313 1447 1327 0 _1481_.Y
rlabel metal1 1824 1202 2076 1218 0 _1541_.gnd
rlabel metal1 1824 1442 2076 1458 0 _1541_.vdd
rlabel metal2 1973 1293 1987 1307 0 _1541_.D
rlabel metal2 1933 1293 1947 1307 0 _1541_.CLK
rlabel metal2 1853 1293 1867 1307 0 _1541_.Q
rlabel metal1 1724 1202 1836 1218 0 _829_.gnd
rlabel metal1 1724 1442 1836 1458 0 _829_.vdd
rlabel metal2 1813 1293 1827 1307 0 _829_.A
rlabel metal2 1793 1313 1807 1327 0 _829_.B
rlabel metal2 1753 1313 1767 1327 0 _829_.C
rlabel metal2 1773 1293 1787 1307 0 _829_.Y
rlabel metal1 1644 1202 1736 1218 0 _828_.gnd
rlabel metal1 1644 1442 1736 1458 0 _828_.vdd
rlabel metal2 1653 1333 1667 1347 0 _828_.A
rlabel metal2 1693 1333 1707 1347 0 _828_.B
rlabel metal2 1673 1313 1687 1327 0 _828_.Y
rlabel metal1 2124 1202 2236 1218 0 _838_.gnd
rlabel metal1 2124 1442 2236 1458 0 _838_.vdd
rlabel metal2 2133 1293 2147 1307 0 _838_.A
rlabel metal2 2153 1313 2167 1327 0 _838_.B
rlabel metal2 2193 1313 2207 1327 0 _838_.C
rlabel metal2 2173 1293 2187 1307 0 _838_.Y
rlabel metal1 2064 1202 2136 1218 0 _836_.gnd
rlabel metal1 2064 1442 2136 1458 0 _836_.vdd
rlabel metal2 2073 1273 2087 1287 0 _836_.A
rlabel metal2 2093 1313 2107 1327 0 _836_.Y
rlabel metal1 2224 1202 2316 1218 0 _837_.gnd
rlabel metal1 2224 1442 2316 1458 0 _837_.vdd
rlabel metal2 2293 1333 2307 1347 0 _837_.A
rlabel metal2 2253 1333 2267 1347 0 _837_.B
rlabel metal2 2273 1313 2287 1327 0 _837_.Y
rlabel metal1 2304 1202 2396 1218 0 _1422_.gnd
rlabel metal1 2304 1442 2396 1458 0 _1422_.vdd
rlabel metal2 2333 1293 2347 1307 0 _1422_.B
rlabel metal2 2373 1293 2387 1307 0 _1422_.A
rlabel metal2 2353 1273 2367 1287 0 _1422_.Y
rlabel metal1 2384 1202 2456 1218 0 _833_.gnd
rlabel metal1 2384 1442 2456 1458 0 _833_.vdd
rlabel metal2 2433 1273 2447 1287 0 _833_.A
rlabel metal2 2413 1313 2427 1327 0 _833_.Y
rlabel metal1 2524 1202 2776 1218 0 _1556_.gnd
rlabel metal1 2524 1442 2776 1458 0 _1556_.vdd
rlabel metal2 2673 1293 2687 1307 0 _1556_.D
rlabel metal2 2633 1293 2647 1307 0 _1556_.CLK
rlabel metal2 2553 1293 2567 1307 0 _1556_.Q
rlabel metal1 2444 1202 2536 1218 0 _1421_.gnd
rlabel metal1 2444 1442 2536 1458 0 _1421_.vdd
rlabel metal2 2493 1293 2507 1307 0 _1421_.B
rlabel metal2 2453 1293 2467 1307 0 _1421_.A
rlabel metal2 2473 1273 2487 1287 0 _1421_.Y
rlabel metal1 2904 1202 3016 1218 0 _1279_.gnd
rlabel metal1 2904 1442 3016 1458 0 _1279_.vdd
rlabel metal2 2913 1293 2927 1307 0 _1279_.A
rlabel metal2 2933 1313 2947 1327 0 _1279_.B
rlabel metal2 2973 1313 2987 1327 0 _1279_.C
rlabel metal2 2953 1293 2967 1307 0 _1279_.Y
rlabel metal1 2764 1202 2856 1218 0 _1280_.gnd
rlabel metal1 2764 1442 2856 1458 0 _1280_.vdd
rlabel metal2 2813 1293 2827 1307 0 _1280_.B
rlabel metal2 2773 1293 2787 1307 0 _1280_.A
rlabel metal2 2793 1273 2807 1287 0 _1280_.Y
rlabel metal1 2844 1202 2916 1218 0 _786_.gnd
rlabel metal1 2844 1442 2916 1458 0 _786_.vdd
rlabel metal2 2893 1313 2907 1327 0 _786_.A
rlabel metal2 2873 1293 2887 1307 0 _786_.Y
rlabel metal1 3004 1202 3116 1218 0 _1256_.gnd
rlabel metal1 3004 1442 3116 1458 0 _1256_.vdd
rlabel metal2 3013 1293 3027 1307 0 _1256_.A
rlabel metal2 3033 1313 3047 1327 0 _1256_.B
rlabel metal2 3073 1313 3087 1327 0 _1256_.C
rlabel metal2 3053 1293 3067 1307 0 _1256_.Y
rlabel metal1 3104 1202 3216 1218 0 _1254_.gnd
rlabel metal1 3104 1442 3216 1458 0 _1254_.vdd
rlabel metal2 3113 1293 3127 1307 0 _1254_.A
rlabel metal2 3133 1313 3147 1327 0 _1254_.B
rlabel metal2 3173 1313 3187 1327 0 _1254_.C
rlabel metal2 3153 1293 3167 1307 0 _1254_.Y
rlabel metal1 3204 1202 3316 1218 0 _1148_.gnd
rlabel metal1 3204 1442 3316 1458 0 _1148_.vdd
rlabel metal2 3213 1293 3227 1307 0 _1148_.A
rlabel metal2 3273 1293 3287 1307 0 _1148_.Y
rlabel metal2 3253 1333 3267 1347 0 _1148_.B
rlabel metal1 3304 1202 3396 1218 0 _1206_.gnd
rlabel metal1 3304 1442 3396 1458 0 _1206_.vdd
rlabel metal2 3333 1293 3347 1307 0 _1206_.B
rlabel metal2 3373 1293 3387 1307 0 _1206_.A
rlabel metal2 3353 1273 3367 1287 0 _1206_.Y
rlabel metal1 3384 1202 3496 1218 0 _1211_.gnd
rlabel metal1 3384 1442 3496 1458 0 _1211_.vdd
rlabel metal2 3393 1313 3407 1327 0 _1211_.A
rlabel metal2 3413 1333 3427 1347 0 _1211_.B
rlabel metal2 3433 1313 3447 1327 0 _1211_.C
rlabel metal2 3453 1333 3467 1347 0 _1211_.Y
rlabel metal1 3584 1202 3696 1218 0 _1214_.gnd
rlabel metal1 3584 1442 3696 1458 0 _1214_.vdd
rlabel metal2 3593 1293 3607 1307 0 _1214_.A
rlabel metal2 3613 1313 3627 1327 0 _1214_.B
rlabel metal2 3653 1313 3667 1327 0 _1214_.C
rlabel metal2 3633 1293 3647 1307 0 _1214_.Y
rlabel metal1 3484 1202 3596 1218 0 _1213_.gnd
rlabel metal1 3484 1442 3596 1458 0 _1213_.vdd
rlabel metal2 3573 1293 3587 1307 0 _1213_.A
rlabel metal2 3553 1313 3567 1327 0 _1213_.B
rlabel metal2 3513 1313 3527 1327 0 _1213_.C
rlabel metal2 3533 1293 3547 1307 0 _1213_.Y
rlabel metal1 3684 1202 3776 1218 0 _1215_.gnd
rlabel metal1 3684 1442 3776 1458 0 _1215_.vdd
rlabel metal2 3753 1333 3767 1347 0 _1215_.A
rlabel metal2 3713 1333 3727 1347 0 _1215_.B
rlabel metal2 3733 1313 3747 1327 0 _1215_.Y
rlabel metal1 3944 1202 4056 1218 0 _1216_.gnd
rlabel metal1 3944 1442 4056 1458 0 _1216_.vdd
rlabel metal2 4033 1293 4047 1307 0 _1216_.A
rlabel metal2 4013 1313 4027 1327 0 _1216_.B
rlabel metal2 3973 1313 3987 1327 0 _1216_.C
rlabel metal2 3993 1293 4007 1307 0 _1216_.Y
rlabel metal1 3764 1202 3856 1218 0 _1156_.gnd
rlabel metal1 3764 1442 3856 1458 0 _1156_.vdd
rlabel metal2 3833 1333 3847 1347 0 _1156_.A
rlabel metal2 3793 1333 3807 1347 0 _1156_.B
rlabel metal2 3813 1313 3827 1327 0 _1156_.Y
rlabel metal1 3844 1202 3956 1218 0 _1170_.gnd
rlabel metal1 3844 1442 3956 1458 0 _1170_.vdd
rlabel metal2 3853 1293 3867 1307 0 _1170_.A
rlabel metal2 3913 1293 3927 1307 0 _1170_.Y
rlabel metal2 3893 1333 3907 1347 0 _1170_.B
rlabel metal1 4104 1202 4196 1218 0 _1249_.gnd
rlabel metal1 4104 1442 4196 1458 0 _1249_.vdd
rlabel metal2 4173 1333 4187 1347 0 _1249_.A
rlabel metal2 4133 1333 4147 1347 0 _1249_.B
rlabel metal2 4153 1313 4167 1327 0 _1249_.Y
rlabel metal1 4184 1202 4276 1218 0 _1221_.gnd
rlabel metal1 4184 1442 4276 1458 0 _1221_.vdd
rlabel metal2 4253 1333 4267 1347 0 _1221_.A
rlabel metal2 4213 1333 4227 1347 0 _1221_.B
rlabel metal2 4233 1313 4247 1327 0 _1221_.Y
rlabel metal1 4264 1202 4356 1218 0 _1164_.gnd
rlabel metal1 4264 1442 4356 1458 0 _1164_.vdd
rlabel metal2 4293 1293 4307 1307 0 _1164_.B
rlabel metal2 4333 1293 4347 1307 0 _1164_.A
rlabel metal2 4313 1273 4327 1287 0 _1164_.Y
rlabel metal1 4044 1202 4116 1218 0 _1166_.gnd
rlabel metal1 4044 1442 4116 1458 0 _1166_.vdd
rlabel metal2 4053 1273 4067 1287 0 _1166_.A
rlabel metal2 4073 1313 4087 1327 0 _1166_.Y
rlabel metal1 4444 1202 4556 1218 0 _1205_.gnd
rlabel metal1 4444 1442 4556 1458 0 _1205_.vdd
rlabel metal2 4453 1293 4467 1307 0 _1205_.A
rlabel metal2 4473 1313 4487 1327 0 _1205_.B
rlabel metal2 4513 1313 4527 1327 0 _1205_.C
rlabel metal2 4493 1293 4507 1307 0 _1205_.Y
rlabel metal1 4344 1202 4456 1218 0 _1169_.gnd
rlabel metal1 4344 1442 4456 1458 0 _1169_.vdd
rlabel metal2 4433 1293 4447 1307 0 _1169_.A
rlabel metal2 4413 1313 4427 1327 0 _1169_.B
rlabel metal2 4373 1313 4387 1327 0 _1169_.C
rlabel metal2 4393 1293 4407 1307 0 _1169_.Y
rlabel nsubstratencontact 4756 1448 4756 1448 0 FILL71250x18150.vdd
rlabel metal1 4744 1202 4776 1218 0 FILL71250x18150.gnd
rlabel nsubstratencontact 4736 1448 4736 1448 0 FILL70950x18150.vdd
rlabel metal1 4724 1202 4756 1218 0 FILL70950x18150.gnd
rlabel metal1 4644 1202 4736 1218 0 _1173_.gnd
rlabel metal1 4644 1442 4736 1458 0 _1173_.vdd
rlabel metal2 4653 1333 4667 1347 0 _1173_.A
rlabel metal2 4693 1333 4707 1347 0 _1173_.B
rlabel metal2 4673 1313 4687 1327 0 _1173_.Y
rlabel metal1 4544 1202 4656 1218 0 _1179_.gnd
rlabel metal1 4544 1442 4656 1458 0 _1179_.vdd
rlabel metal2 4633 1313 4647 1327 0 _1179_.A
rlabel metal2 4613 1273 4627 1287 0 _1179_.B
rlabel metal2 4593 1313 4607 1327 0 _1179_.C
rlabel metal2 4573 1293 4587 1307 0 _1179_.Y
rlabel metal1 4 1682 216 1698 0 CLKBUF1_insert8.gnd
rlabel metal1 4 1442 216 1458 0 CLKBUF1_insert8.vdd
rlabel metal2 33 1573 47 1587 0 CLKBUF1_insert8.A
rlabel metal2 173 1573 187 1587 0 CLKBUF1_insert8.Y
rlabel metal1 204 1682 296 1698 0 _774_.gnd
rlabel metal1 204 1442 296 1458 0 _774_.vdd
rlabel metal2 233 1593 247 1607 0 _774_.B
rlabel metal2 273 1593 287 1607 0 _774_.A
rlabel metal2 253 1613 267 1627 0 _774_.Y
rlabel metal1 284 1682 376 1698 0 BUFX2_insert16.gnd
rlabel metal1 284 1442 376 1458 0 BUFX2_insert16.vdd
rlabel metal2 353 1593 367 1607 0 BUFX2_insert16.A
rlabel metal2 313 1593 327 1607 0 BUFX2_insert16.Y
rlabel metal1 364 1682 616 1698 0 _1599_.gnd
rlabel metal1 364 1442 616 1458 0 _1599_.vdd
rlabel metal2 453 1593 467 1607 0 _1599_.D
rlabel metal2 493 1593 507 1607 0 _1599_.CLK
rlabel metal2 573 1593 587 1607 0 _1599_.Q
rlabel metal1 604 1682 856 1698 0 _1600_.gnd
rlabel metal1 604 1442 856 1458 0 _1600_.vdd
rlabel metal2 693 1593 707 1607 0 _1600_.D
rlabel metal2 733 1593 747 1607 0 _1600_.CLK
rlabel metal2 813 1593 827 1607 0 _1600_.Q
rlabel metal1 844 1682 1096 1698 0 _1598_.gnd
rlabel metal1 844 1442 1096 1458 0 _1598_.vdd
rlabel metal2 993 1593 1007 1607 0 _1598_.D
rlabel metal2 953 1593 967 1607 0 _1598_.CLK
rlabel metal2 873 1593 887 1607 0 _1598_.Q
rlabel metal1 1264 1682 1516 1698 0 _1579_.gnd
rlabel metal1 1264 1442 1516 1458 0 _1579_.vdd
rlabel metal2 1413 1593 1427 1607 0 _1579_.D
rlabel metal2 1373 1593 1387 1607 0 _1579_.CLK
rlabel metal2 1293 1593 1307 1607 0 _1579_.Q
rlabel metal1 1164 1682 1276 1698 0 _1491_.gnd
rlabel metal1 1164 1442 1276 1458 0 _1491_.vdd
rlabel metal2 1253 1593 1267 1607 0 _1491_.A
rlabel metal2 1233 1573 1247 1587 0 _1491_.B
rlabel metal2 1193 1573 1207 1587 0 _1491_.C
rlabel metal2 1213 1593 1227 1607 0 _1491_.Y
rlabel metal1 1084 1682 1176 1698 0 _1490_.gnd
rlabel metal1 1084 1442 1176 1458 0 _1490_.vdd
rlabel metal2 1153 1553 1167 1567 0 _1490_.A
rlabel metal2 1113 1553 1127 1567 0 _1490_.B
rlabel metal2 1133 1573 1147 1587 0 _1490_.Y
rlabel metal1 1504 1682 1756 1698 0 _1580_.gnd
rlabel metal1 1504 1442 1756 1458 0 _1580_.vdd
rlabel metal2 1593 1593 1607 1607 0 _1580_.D
rlabel metal2 1633 1593 1647 1607 0 _1580_.CLK
rlabel metal2 1713 1593 1727 1607 0 _1580_.Q
rlabel metal1 1744 1682 1856 1698 0 _1494_.gnd
rlabel metal1 1744 1442 1856 1458 0 _1494_.vdd
rlabel metal2 1833 1573 1847 1587 0 _1494_.A
rlabel metal2 1813 1613 1827 1627 0 _1494_.B
rlabel metal2 1793 1573 1807 1587 0 _1494_.C
rlabel metal2 1773 1593 1787 1607 0 _1494_.Y
rlabel metal1 1844 1682 1936 1698 0 _1493_.gnd
rlabel metal1 1844 1442 1936 1458 0 _1493_.vdd
rlabel metal2 1893 1593 1907 1607 0 _1493_.B
rlabel metal2 1853 1593 1867 1607 0 _1493_.A
rlabel metal2 1873 1613 1887 1627 0 _1493_.Y
rlabel metal1 1924 1682 2176 1698 0 _1583_.gnd
rlabel metal1 1924 1442 2176 1458 0 _1583_.vdd
rlabel metal2 2013 1593 2027 1607 0 _1583_.D
rlabel metal2 2053 1593 2067 1607 0 _1583_.CLK
rlabel metal2 2133 1593 2147 1607 0 _1583_.Q
rlabel metal1 2324 1682 2436 1698 0 _835_.gnd
rlabel metal1 2324 1442 2436 1458 0 _835_.vdd
rlabel metal2 2333 1593 2347 1607 0 _835_.A
rlabel metal2 2353 1573 2367 1587 0 _835_.B
rlabel metal2 2393 1573 2407 1587 0 _835_.C
rlabel metal2 2373 1593 2387 1607 0 _835_.Y
rlabel metal1 2244 1682 2336 1698 0 _834_.gnd
rlabel metal1 2244 1442 2336 1458 0 _834_.vdd
rlabel metal2 2313 1553 2327 1567 0 _834_.A
rlabel metal2 2273 1553 2287 1567 0 _834_.B
rlabel metal2 2293 1573 2307 1587 0 _834_.Y
rlabel metal1 2164 1682 2256 1698 0 _1499_.gnd
rlabel metal1 2164 1442 2256 1458 0 _1499_.vdd
rlabel metal2 2193 1593 2207 1607 0 _1499_.B
rlabel metal2 2233 1593 2247 1607 0 _1499_.A
rlabel metal2 2213 1613 2227 1627 0 _1499_.Y
rlabel metal1 2424 1682 2676 1698 0 _1540_.gnd
rlabel metal1 2424 1442 2676 1458 0 _1540_.vdd
rlabel metal2 2573 1593 2587 1607 0 _1540_.D
rlabel metal2 2533 1593 2547 1607 0 _1540_.CLK
rlabel metal2 2453 1593 2467 1607 0 _1540_.Q
rlabel metal1 2664 1682 2916 1698 0 _1526_.gnd
rlabel metal1 2664 1442 2916 1458 0 _1526_.vdd
rlabel metal2 2753 1593 2767 1607 0 _1526_.D
rlabel metal2 2793 1593 2807 1607 0 _1526_.CLK
rlabel metal2 2873 1593 2887 1607 0 _1526_.Q
rlabel metal1 2904 1682 2976 1698 0 _792_.gnd
rlabel metal1 2904 1442 2976 1458 0 _792_.vdd
rlabel metal2 2913 1573 2927 1587 0 _792_.A
rlabel metal2 2933 1593 2947 1607 0 _792_.Y
rlabel metal1 3124 1682 3236 1698 0 _1252_.gnd
rlabel metal1 3124 1442 3236 1458 0 _1252_.vdd
rlabel metal2 3133 1593 3147 1607 0 _1252_.A
rlabel metal2 3153 1573 3167 1587 0 _1252_.B
rlabel metal2 3193 1573 3207 1587 0 _1252_.C
rlabel metal2 3173 1593 3187 1607 0 _1252_.Y
rlabel metal1 2964 1682 3056 1698 0 _1253_.gnd
rlabel metal1 2964 1442 3056 1458 0 _1253_.vdd
rlabel metal2 2973 1553 2987 1567 0 _1253_.A
rlabel metal2 3013 1553 3027 1567 0 _1253_.B
rlabel metal2 2993 1573 3007 1587 0 _1253_.Y
rlabel metal1 3044 1682 3136 1698 0 _1251_.gnd
rlabel metal1 3044 1442 3136 1458 0 _1251_.vdd
rlabel metal2 3113 1553 3127 1567 0 _1251_.A
rlabel metal2 3073 1553 3087 1567 0 _1251_.B
rlabel metal2 3093 1573 3107 1587 0 _1251_.Y
rlabel metal1 3384 1682 3496 1698 0 _1210_.gnd
rlabel metal1 3384 1442 3496 1458 0 _1210_.vdd
rlabel metal2 3473 1593 3487 1607 0 _1210_.A
rlabel metal2 3453 1573 3467 1587 0 _1210_.B
rlabel metal2 3413 1573 3427 1587 0 _1210_.C
rlabel metal2 3433 1593 3447 1607 0 _1210_.Y
rlabel metal1 3224 1682 3316 1698 0 _1207_.gnd
rlabel metal1 3224 1442 3316 1458 0 _1207_.vdd
rlabel metal2 3233 1553 3247 1567 0 _1207_.A
rlabel metal2 3273 1553 3287 1567 0 _1207_.B
rlabel metal2 3253 1573 3267 1587 0 _1207_.Y
rlabel metal1 3304 1682 3396 1698 0 _1153_.gnd
rlabel metal1 3304 1442 3396 1458 0 _1153_.vdd
rlabel metal2 3373 1553 3387 1567 0 _1153_.A
rlabel metal2 3333 1553 3347 1567 0 _1153_.B
rlabel metal2 3353 1573 3367 1587 0 _1153_.Y
rlabel metal1 3704 1682 3776 1698 0 _1151_.gnd
rlabel metal1 3704 1442 3776 1458 0 _1151_.vdd
rlabel metal2 3713 1613 3727 1627 0 _1151_.A
rlabel metal2 3733 1573 3747 1587 0 _1151_.Y
rlabel metal1 3484 1682 3596 1698 0 _1149_.gnd
rlabel metal1 3484 1442 3596 1458 0 _1149_.vdd
rlabel metal2 3493 1573 3507 1587 0 _1149_.A
rlabel metal2 3513 1553 3527 1567 0 _1149_.B
rlabel metal2 3533 1573 3547 1587 0 _1149_.C
rlabel metal2 3553 1553 3567 1567 0 _1149_.Y
rlabel metal1 3584 1682 3716 1698 0 _1155_.gnd
rlabel metal1 3584 1442 3716 1458 0 _1155_.vdd
rlabel metal2 3693 1593 3707 1607 0 _1155_.A
rlabel metal2 3673 1573 3687 1587 0 _1155_.B
rlabel metal2 3613 1593 3627 1607 0 _1155_.C
rlabel metal2 3653 1593 3667 1607 0 _1155_.Y
rlabel metal2 3633 1573 3647 1587 0 _1155_.D
rlabel metal1 3964 1682 4076 1698 0 _1217_.gnd
rlabel metal1 3964 1442 4076 1458 0 _1217_.vdd
rlabel metal2 3973 1593 3987 1607 0 _1217_.A
rlabel metal2 3993 1573 4007 1587 0 _1217_.B
rlabel metal2 4033 1573 4047 1587 0 _1217_.C
rlabel metal2 4013 1593 4027 1607 0 _1217_.Y
rlabel metal1 3864 1682 3976 1698 0 _1202_.gnd
rlabel metal1 3864 1442 3976 1458 0 _1202_.vdd
rlabel metal2 3873 1573 3887 1587 0 _1202_.A
rlabel metal2 3893 1613 3907 1627 0 _1202_.B
rlabel metal2 3913 1573 3927 1587 0 _1202_.C
rlabel metal2 3933 1593 3947 1607 0 _1202_.Y
rlabel metal1 3764 1682 3876 1698 0 _1152_.gnd
rlabel metal1 3764 1442 3876 1458 0 _1152_.vdd
rlabel metal2 3773 1573 3787 1587 0 _1152_.A
rlabel metal2 3793 1553 3807 1567 0 _1152_.B
rlabel metal2 3813 1573 3827 1587 0 _1152_.C
rlabel metal2 3833 1553 3847 1567 0 _1152_.Y
rlabel metal1 4244 1682 4356 1698 0 _1163_.gnd
rlabel metal1 4244 1442 4356 1458 0 _1163_.vdd
rlabel metal2 4253 1593 4267 1607 0 _1163_.A
rlabel metal2 4273 1573 4287 1587 0 _1163_.B
rlabel metal2 4313 1573 4327 1587 0 _1163_.C
rlabel metal2 4293 1593 4307 1607 0 _1163_.Y
rlabel metal1 4064 1682 4156 1698 0 _1160_.gnd
rlabel metal1 4064 1442 4156 1458 0 _1160_.vdd
rlabel metal2 4133 1553 4147 1567 0 _1160_.A
rlabel metal2 4093 1553 4107 1567 0 _1160_.B
rlabel metal2 4113 1573 4127 1587 0 _1160_.Y
rlabel metal1 4144 1682 4256 1698 0 _1167_.gnd
rlabel metal1 4144 1442 4256 1458 0 _1167_.vdd
rlabel metal2 4153 1573 4167 1587 0 _1167_.A
rlabel metal2 4173 1613 4187 1627 0 _1167_.B
rlabel metal2 4193 1573 4207 1587 0 _1167_.C
rlabel metal2 4213 1593 4227 1607 0 _1167_.Y
rlabel metal1 4484 1682 4576 1698 0 _1204_.gnd
rlabel metal1 4484 1442 4576 1458 0 _1204_.vdd
rlabel metal2 4493 1553 4507 1567 0 _1204_.A
rlabel metal2 4533 1553 4547 1567 0 _1204_.B
rlabel metal2 4513 1573 4527 1587 0 _1204_.Y
rlabel metal1 4404 1682 4496 1698 0 _1168_.gnd
rlabel metal1 4404 1442 4496 1458 0 _1168_.vdd
rlabel metal2 4453 1593 4467 1607 0 _1168_.B
rlabel metal2 4413 1593 4427 1607 0 _1168_.A
rlabel metal2 4433 1613 4447 1627 0 _1168_.Y
rlabel metal1 4344 1682 4416 1698 0 _1162_.gnd
rlabel metal1 4344 1442 4416 1458 0 _1162_.vdd
rlabel metal2 4353 1613 4367 1627 0 _1162_.A
rlabel metal2 4373 1573 4387 1587 0 _1162_.Y
rlabel nsubstratencontact 4764 1452 4764 1452 0 FILL71250x21750.vdd
rlabel metal1 4744 1682 4776 1698 0 FILL71250x21750.gnd
rlabel nsubstratencontact 4744 1452 4744 1452 0 FILL70950x21750.vdd
rlabel metal1 4724 1682 4756 1698 0 FILL70950x21750.gnd
rlabel metal1 4564 1682 4656 1698 0 _1172_.gnd
rlabel metal1 4564 1442 4656 1458 0 _1172_.vdd
rlabel metal2 4573 1553 4587 1567 0 _1172_.A
rlabel metal2 4613 1553 4627 1567 0 _1172_.B
rlabel metal2 4593 1573 4607 1587 0 _1172_.Y
rlabel metal1 4644 1682 4736 1698 0 _1171_.gnd
rlabel metal1 4644 1442 4736 1458 0 _1171_.vdd
rlabel metal2 4653 1553 4667 1567 0 _1171_.A
rlabel metal2 4693 1553 4707 1567 0 _1171_.B
rlabel metal2 4673 1573 4687 1587 0 _1171_.Y
rlabel metal1 4 1682 256 1698 0 _1562_.gnd
rlabel metal1 4 1922 256 1938 0 _1562_.vdd
rlabel metal2 93 1773 107 1787 0 _1562_.D
rlabel metal2 133 1773 147 1787 0 _1562_.CLK
rlabel metal2 213 1773 227 1787 0 _1562_.Q
rlabel metal1 244 1682 356 1698 0 _777_.gnd
rlabel metal1 244 1922 356 1938 0 _777_.vdd
rlabel metal2 253 1773 267 1787 0 _777_.A
rlabel metal2 273 1793 287 1807 0 _777_.B
rlabel metal2 313 1793 327 1807 0 _777_.C
rlabel metal2 293 1773 307 1787 0 _777_.Y
rlabel metal1 344 1682 456 1698 0 _775_.gnd
rlabel metal1 344 1922 456 1938 0 _775_.vdd
rlabel metal2 433 1773 447 1787 0 _775_.A
rlabel metal2 413 1793 427 1807 0 _775_.B
rlabel metal2 373 1793 387 1807 0 _775_.C
rlabel metal2 393 1773 407 1787 0 _775_.Y
rlabel metal1 444 1682 556 1698 0 _767_.gnd
rlabel metal1 444 1922 556 1938 0 _767_.vdd
rlabel metal2 533 1773 547 1787 0 _767_.A
rlabel metal2 513 1793 527 1807 0 _767_.B
rlabel metal2 473 1793 487 1807 0 _767_.C
rlabel metal2 493 1773 507 1787 0 _767_.Y
rlabel metal1 544 1682 656 1698 0 _763_.gnd
rlabel metal1 544 1922 656 1938 0 _763_.vdd
rlabel metal2 633 1773 647 1787 0 _763_.A
rlabel metal2 613 1793 627 1807 0 _763_.B
rlabel metal2 573 1793 587 1807 0 _763_.C
rlabel metal2 593 1773 607 1787 0 _763_.Y
rlabel metal1 764 1682 856 1698 0 _1492_.gnd
rlabel metal1 764 1922 856 1938 0 _1492_.vdd
rlabel metal2 793 1773 807 1787 0 _1492_.B
rlabel metal2 833 1773 847 1787 0 _1492_.A
rlabel metal2 813 1753 827 1767 0 _1492_.Y
rlabel metal1 704 1682 776 1698 0 _768_.gnd
rlabel metal1 704 1922 776 1938 0 _768_.vdd
rlabel metal2 713 1753 727 1767 0 _768_.A
rlabel metal2 733 1793 747 1807 0 _768_.Y
rlabel metal1 644 1682 716 1698 0 _761_.gnd
rlabel metal1 644 1922 716 1938 0 _761_.vdd
rlabel metal2 653 1753 667 1767 0 _761_.A
rlabel metal2 673 1793 687 1807 0 _761_.Y
rlabel metal1 944 1682 1196 1698 0 _1578_.gnd
rlabel metal1 944 1922 1196 1938 0 _1578_.vdd
rlabel metal2 1033 1773 1047 1787 0 _1578_.D
rlabel metal2 1073 1773 1087 1787 0 _1578_.CLK
rlabel metal2 1153 1773 1167 1787 0 _1578_.Q
rlabel metal1 844 1682 956 1698 0 _1480_.gnd
rlabel metal1 844 1922 956 1938 0 _1480_.vdd
rlabel metal2 853 1793 867 1807 0 _1480_.A
rlabel metal2 873 1813 887 1827 0 _1480_.B
rlabel metal2 893 1793 907 1807 0 _1480_.C
rlabel metal2 913 1813 927 1827 0 _1480_.Y
rlabel metal1 1264 1682 1376 1698 0 _1488_.gnd
rlabel metal1 1264 1922 1376 1938 0 _1488_.vdd
rlabel metal2 1353 1773 1367 1787 0 _1488_.A
rlabel metal2 1333 1793 1347 1807 0 _1488_.B
rlabel metal2 1293 1793 1307 1807 0 _1488_.C
rlabel metal2 1313 1773 1327 1787 0 _1488_.Y
rlabel metal1 1184 1682 1276 1698 0 _1487_.gnd
rlabel metal1 1184 1922 1276 1938 0 _1487_.vdd
rlabel metal2 1193 1813 1207 1827 0 _1487_.A
rlabel metal2 1233 1813 1247 1827 0 _1487_.B
rlabel metal2 1213 1793 1227 1807 0 _1487_.Y
rlabel metal1 1364 1682 1576 1698 0 CLKBUF1_insert13.gnd
rlabel metal1 1364 1922 1576 1938 0 CLKBUF1_insert13.vdd
rlabel metal2 1533 1793 1547 1807 0 CLKBUF1_insert13.A
rlabel metal2 1393 1793 1407 1807 0 CLKBUF1_insert13.Y
rlabel metal1 1564 1682 1816 1698 0 _1581_.gnd
rlabel metal1 1564 1922 1816 1938 0 _1581_.vdd
rlabel metal2 1653 1773 1667 1787 0 _1581_.D
rlabel metal2 1693 1773 1707 1787 0 _1581_.CLK
rlabel metal2 1773 1773 1787 1787 0 _1581_.Q
rlabel metal1 1804 1682 1916 1698 0 _1496_.gnd
rlabel metal1 1804 1922 1916 1938 0 _1496_.vdd
rlabel metal2 1893 1793 1907 1807 0 _1496_.A
rlabel metal2 1873 1753 1887 1767 0 _1496_.B
rlabel metal2 1853 1793 1867 1807 0 _1496_.C
rlabel metal2 1833 1773 1847 1787 0 _1496_.Y
rlabel metal1 1984 1682 2096 1698 0 _1500_.gnd
rlabel metal1 1984 1922 2096 1938 0 _1500_.vdd
rlabel metal2 2073 1793 2087 1807 0 _1500_.A
rlabel metal2 2053 1753 2067 1767 0 _1500_.B
rlabel metal2 2033 1793 2047 1807 0 _1500_.C
rlabel metal2 2013 1773 2027 1787 0 _1500_.Y
rlabel metal1 2084 1682 2176 1698 0 _1497_.gnd
rlabel metal1 2084 1922 2176 1938 0 _1497_.vdd
rlabel metal2 2113 1773 2127 1787 0 _1497_.B
rlabel metal2 2153 1773 2167 1787 0 _1497_.A
rlabel metal2 2133 1753 2147 1767 0 _1497_.Y
rlabel metal1 1904 1682 1996 1698 0 _1495_.gnd
rlabel metal1 1904 1922 1996 1938 0 _1495_.vdd
rlabel metal2 1953 1773 1967 1787 0 _1495_.B
rlabel metal2 1913 1773 1927 1787 0 _1495_.A
rlabel metal2 1933 1753 1947 1767 0 _1495_.Y
rlabel metal1 2264 1682 2516 1698 0 _1582_.gnd
rlabel metal1 2264 1922 2516 1938 0 _1582_.vdd
rlabel metal2 2413 1773 2427 1787 0 _1582_.D
rlabel metal2 2373 1773 2387 1787 0 _1582_.CLK
rlabel metal2 2293 1773 2307 1787 0 _1582_.Q
rlabel metal1 2164 1682 2276 1698 0 _1498_.gnd
rlabel metal1 2164 1922 2276 1938 0 _1498_.vdd
rlabel metal2 2173 1793 2187 1807 0 _1498_.A
rlabel metal2 2193 1753 2207 1767 0 _1498_.B
rlabel metal2 2213 1793 2227 1807 0 _1498_.C
rlabel metal2 2233 1773 2247 1787 0 _1498_.Y
rlabel metal1 2504 1682 2756 1698 0 _1529_.gnd
rlabel metal1 2504 1922 2756 1938 0 _1529_.vdd
rlabel metal2 2593 1773 2607 1787 0 _1529_.D
rlabel metal2 2633 1773 2647 1787 0 _1529_.CLK
rlabel metal2 2713 1773 2727 1787 0 _1529_.Q
rlabel metal1 2744 1682 2996 1698 0 _1527_.gnd
rlabel metal1 2744 1922 2996 1938 0 _1527_.vdd
rlabel metal2 2833 1773 2847 1787 0 _1527_.D
rlabel metal2 2873 1773 2887 1787 0 _1527_.CLK
rlabel metal2 2953 1773 2967 1787 0 _1527_.Q
rlabel metal1 3044 1682 3136 1698 0 _1085_.gnd
rlabel metal1 3044 1922 3136 1938 0 _1085_.vdd
rlabel metal2 3113 1813 3127 1827 0 _1085_.A
rlabel metal2 3073 1813 3087 1827 0 _1085_.B
rlabel metal2 3093 1793 3107 1807 0 _1085_.Y
rlabel metal1 3184 1682 3296 1698 0 _1271_.gnd
rlabel metal1 3184 1922 3296 1938 0 _1271_.vdd
rlabel metal2 3193 1793 3207 1807 0 _1271_.A
rlabel metal2 3213 1753 3227 1767 0 _1271_.B
rlabel metal2 3233 1793 3247 1807 0 _1271_.C
rlabel metal2 3253 1773 3267 1787 0 _1271_.Y
rlabel metal1 3124 1682 3196 1698 0 _962_.gnd
rlabel metal1 3124 1922 3196 1938 0 _962_.vdd
rlabel metal2 3173 1793 3187 1807 0 _962_.A
rlabel metal2 3153 1773 3167 1787 0 _962_.Y
rlabel metal1 2984 1682 3056 1698 0 _783_.gnd
rlabel metal1 2984 1922 3056 1938 0 _783_.vdd
rlabel metal2 3033 1793 3047 1807 0 _783_.A
rlabel metal2 3013 1773 3027 1787 0 _783_.Y
rlabel metal1 3284 1682 3376 1698 0 _1154_.gnd
rlabel metal1 3284 1922 3376 1938 0 _1154_.vdd
rlabel metal2 3333 1773 3347 1787 0 _1154_.B
rlabel metal2 3293 1773 3307 1787 0 _1154_.A
rlabel metal2 3313 1753 3327 1767 0 _1154_.Y
rlabel metal1 3364 1682 3476 1698 0 _1078_.gnd
rlabel metal1 3364 1922 3476 1938 0 _1078_.vdd
rlabel metal2 3453 1773 3467 1787 0 _1078_.A
rlabel metal2 3393 1773 3407 1787 0 _1078_.Y
rlabel metal2 3413 1813 3427 1827 0 _1078_.B
rlabel metal1 3464 1682 3536 1698 0 _1146_.gnd
rlabel metal1 3464 1922 3536 1938 0 _1146_.vdd
rlabel metal2 3473 1793 3487 1807 0 _1146_.A
rlabel metal2 3493 1773 3507 1787 0 _1146_.Y
rlabel metal1 3704 1682 3796 1698 0 _1147_.gnd
rlabel metal1 3704 1922 3796 1938 0 _1147_.vdd
rlabel metal2 3733 1773 3747 1787 0 _1147_.B
rlabel metal2 3773 1773 3787 1787 0 _1147_.A
rlabel metal2 3753 1753 3767 1767 0 _1147_.Y
rlabel metal1 3524 1682 3656 1698 0 _1150_.gnd
rlabel metal1 3524 1922 3656 1938 0 _1150_.vdd
rlabel metal2 3633 1773 3647 1787 0 _1150_.A
rlabel metal2 3613 1793 3627 1807 0 _1150_.B
rlabel metal2 3553 1773 3567 1787 0 _1150_.C
rlabel metal2 3573 1793 3587 1807 0 _1150_.D
rlabel metal2 3593 1773 3607 1787 0 _1150_.Y
rlabel metal1 3644 1682 3716 1698 0 _789_.gnd
rlabel metal1 3644 1922 3716 1938 0 _789_.vdd
rlabel metal2 3693 1793 3707 1807 0 _789_.A
rlabel metal2 3673 1773 3687 1787 0 _789_.Y
rlabel metal1 3784 1682 3876 1698 0 BUFX2_insert33.gnd
rlabel metal1 3784 1922 3876 1938 0 BUFX2_insert33.vdd
rlabel metal2 3793 1773 3807 1787 0 BUFX2_insert33.A
rlabel metal2 3833 1773 3847 1787 0 BUFX2_insert33.Y
rlabel metal1 3964 1682 4096 1698 0 _1097_.gnd
rlabel metal1 3964 1922 4096 1938 0 _1097_.vdd
rlabel metal2 4073 1773 4087 1787 0 _1097_.A
rlabel metal2 4053 1793 4067 1807 0 _1097_.B
rlabel metal2 3993 1773 4007 1787 0 _1097_.C
rlabel metal2 4013 1793 4027 1807 0 _1097_.D
rlabel metal2 4033 1773 4047 1787 0 _1097_.Y
rlabel metal1 3864 1682 3976 1698 0 _1091_.gnd
rlabel metal1 3864 1922 3976 1938 0 _1091_.vdd
rlabel metal2 3873 1773 3887 1787 0 _1091_.A
rlabel metal2 3933 1773 3947 1787 0 _1091_.Y
rlabel metal2 3913 1813 3927 1827 0 _1091_.B
rlabel metal1 4204 1682 4296 1698 0 _1159_.gnd
rlabel metal1 4204 1922 4296 1938 0 _1159_.vdd
rlabel metal2 4213 1813 4227 1827 0 _1159_.A
rlabel metal2 4253 1813 4267 1827 0 _1159_.B
rlabel metal2 4233 1793 4247 1807 0 _1159_.Y
rlabel metal1 4084 1682 4216 1698 0 _1161_.gnd
rlabel metal1 4084 1922 4216 1938 0 _1161_.vdd
rlabel metal2 4093 1773 4107 1787 0 _1161_.A
rlabel metal2 4113 1793 4127 1807 0 _1161_.B
rlabel metal2 4173 1773 4187 1787 0 _1161_.C
rlabel metal2 4153 1793 4167 1807 0 _1161_.D
rlabel metal2 4133 1773 4147 1787 0 _1161_.Y
rlabel metal1 4504 1682 4576 1698 0 _1095_.gnd
rlabel metal1 4504 1922 4576 1938 0 _1095_.vdd
rlabel metal2 4553 1753 4567 1767 0 _1095_.A
rlabel metal2 4533 1793 4547 1807 0 _1095_.Y
rlabel metal1 4384 1682 4516 1698 0 _1158_.gnd
rlabel metal1 4384 1922 4516 1938 0 _1158_.vdd
rlabel metal2 4393 1773 4407 1787 0 _1158_.A
rlabel metal2 4413 1793 4427 1807 0 _1158_.B
rlabel metal2 4473 1773 4487 1787 0 _1158_.C
rlabel metal2 4453 1793 4467 1807 0 _1158_.D
rlabel metal2 4433 1773 4447 1787 0 _1158_.Y
rlabel metal1 4284 1682 4396 1698 0 _1157_.gnd
rlabel metal1 4284 1922 4396 1938 0 _1157_.vdd
rlabel metal2 4293 1773 4307 1787 0 _1157_.A
rlabel metal2 4353 1773 4367 1787 0 _1157_.Y
rlabel metal2 4333 1813 4347 1827 0 _1157_.B
rlabel nsubstratencontact 4756 1928 4756 1928 0 FILL71250x25350.vdd
rlabel metal1 4744 1682 4776 1698 0 FILL71250x25350.gnd
rlabel nsubstratencontact 4736 1928 4736 1928 0 FILL70950x25350.vdd
rlabel metal1 4724 1682 4756 1698 0 FILL70950x25350.gnd
rlabel metal1 4564 1682 4676 1698 0 _1165_.gnd
rlabel metal1 4564 1922 4676 1938 0 _1165_.vdd
rlabel metal2 4573 1773 4587 1787 0 _1165_.A
rlabel metal2 4593 1793 4607 1807 0 _1165_.B
rlabel metal2 4633 1793 4647 1807 0 _1165_.C
rlabel metal2 4613 1773 4627 1787 0 _1165_.Y
rlabel metal1 4664 1682 4736 1698 0 _1098_.gnd
rlabel metal1 4664 1922 4736 1938 0 _1098_.vdd
rlabel metal2 4673 1753 4687 1767 0 _1098_.A
rlabel metal2 4693 1793 4707 1807 0 _1098_.Y
rlabel metal1 4 2162 216 2178 0 CLKBUF1_insert9.gnd
rlabel metal1 4 1922 216 1938 0 CLKBUF1_insert9.vdd
rlabel metal2 33 2053 47 2067 0 CLKBUF1_insert9.A
rlabel metal2 173 2053 187 2067 0 CLKBUF1_insert9.Y
rlabel metal1 204 2162 296 2178 0 _1339_.gnd
rlabel metal1 204 1922 296 1938 0 _1339_.vdd
rlabel metal2 273 2033 287 2047 0 _1339_.A
rlabel metal2 233 2033 247 2047 0 _1339_.B
rlabel metal2 253 2053 267 2067 0 _1339_.Y
rlabel metal1 504 2162 756 2178 0 _1532_.gnd
rlabel metal1 504 1922 756 1938 0 _1532_.vdd
rlabel metal2 593 2073 607 2087 0 _1532_.D
rlabel metal2 633 2073 647 2087 0 _1532_.CLK
rlabel metal2 713 2073 727 2087 0 _1532_.Q
rlabel metal1 284 2162 396 2178 0 _1340_.gnd
rlabel metal1 284 1922 396 1938 0 _1340_.vdd
rlabel metal2 373 2073 387 2087 0 _1340_.A
rlabel metal2 353 2053 367 2067 0 _1340_.B
rlabel metal2 313 2053 327 2067 0 _1340_.C
rlabel metal2 333 2073 347 2087 0 _1340_.Y
rlabel metal1 384 2162 516 2178 0 _776_.gnd
rlabel metal1 384 1922 516 1938 0 _776_.vdd
rlabel metal2 393 2073 407 2087 0 _776_.A
rlabel metal2 413 2053 427 2067 0 _776_.B
rlabel metal2 473 2073 487 2087 0 _776_.C
rlabel metal2 453 2053 467 2067 0 _776_.D
rlabel metal2 433 2073 447 2087 0 _776_.Y
rlabel metal1 744 2162 836 2178 0 _1338_.gnd
rlabel metal1 744 1922 836 1938 0 _1338_.vdd
rlabel metal2 813 2033 827 2047 0 _1338_.A
rlabel metal2 773 2033 787 2047 0 _1338_.B
rlabel metal2 793 2053 807 2067 0 _1338_.Y
rlabel metal1 924 2162 1016 2178 0 _1336_.gnd
rlabel metal1 924 1922 1016 1938 0 _1336_.vdd
rlabel metal2 933 2033 947 2047 0 _1336_.A
rlabel metal2 973 2033 987 2047 0 _1336_.B
rlabel metal2 953 2053 967 2067 0 _1336_.Y
rlabel metal1 1004 2162 1096 2178 0 _762_.gnd
rlabel metal1 1004 1922 1096 1938 0 _762_.vdd
rlabel metal2 1053 2073 1067 2087 0 _762_.B
rlabel metal2 1013 2073 1027 2087 0 _762_.A
rlabel metal2 1033 2093 1047 2107 0 _762_.Y
rlabel metal1 824 2162 936 2178 0 _1337_.gnd
rlabel metal1 824 1922 936 1938 0 _1337_.vdd
rlabel metal2 913 2093 927 2107 0 _1337_.A
rlabel metal2 893 2073 907 2087 0 _1337_.B
rlabel metal2 853 2053 867 2067 0 _1337_.Y
rlabel metal1 1084 2162 1196 2178 0 _811_.gnd
rlabel metal1 1084 1922 1196 1938 0 _811_.vdd
rlabel metal2 1093 2073 1107 2087 0 _811_.A
rlabel metal2 1113 2053 1127 2067 0 _811_.B
rlabel metal2 1153 2053 1167 2067 0 _811_.C
rlabel metal2 1133 2073 1147 2087 0 _811_.Y
rlabel metal1 1184 2162 1276 2178 0 _810_.gnd
rlabel metal1 1184 1922 1276 1938 0 _810_.vdd
rlabel metal2 1193 2033 1207 2047 0 _810_.A
rlabel metal2 1233 2033 1247 2047 0 _810_.B
rlabel metal2 1213 2053 1227 2067 0 _810_.Y
rlabel metal1 1264 2162 1356 2178 0 _1514_.gnd
rlabel metal1 1264 1922 1356 1938 0 _1514_.vdd
rlabel metal2 1313 2073 1327 2087 0 _1514_.B
rlabel metal2 1273 2073 1287 2087 0 _1514_.A
rlabel metal2 1293 2093 1307 2107 0 _1514_.Y
rlabel metal1 1344 2162 1596 2178 0 _1590_.gnd
rlabel metal1 1344 1922 1596 1938 0 _1590_.vdd
rlabel metal2 1493 2073 1507 2087 0 _1590_.D
rlabel metal2 1453 2073 1467 2087 0 _1590_.CLK
rlabel metal2 1373 2073 1387 2087 0 _1590_.Q
rlabel metal1 1584 2162 1696 2178 0 _1515_.gnd
rlabel metal1 1584 1922 1696 1938 0 _1515_.vdd
rlabel metal2 1673 2053 1687 2067 0 _1515_.A
rlabel metal2 1653 2093 1667 2107 0 _1515_.B
rlabel metal2 1633 2053 1647 2067 0 _1515_.C
rlabel metal2 1613 2073 1627 2087 0 _1515_.Y
rlabel metal1 1684 2162 1776 2178 0 BUFX2_insert25.gnd
rlabel metal1 1684 1922 1776 1938 0 BUFX2_insert25.vdd
rlabel metal2 1753 2073 1767 2087 0 BUFX2_insert25.A
rlabel metal2 1713 2073 1727 2087 0 BUFX2_insert25.Y
rlabel metal1 1764 2162 2016 2178 0 _1597_.gnd
rlabel metal1 1764 1922 2016 1938 0 _1597_.vdd
rlabel metal2 1913 2073 1927 2087 0 _1597_.D
rlabel metal2 1873 2073 1887 2087 0 _1597_.CLK
rlabel metal2 1793 2073 1807 2087 0 _1597_.Q
rlabel metal1 2064 2162 2156 2178 0 _1518_.gnd
rlabel metal1 2064 1922 2156 1938 0 _1518_.vdd
rlabel metal2 2133 2033 2147 2047 0 _1518_.A
rlabel metal2 2093 2033 2107 2047 0 _1518_.B
rlabel metal2 2113 2053 2127 2067 0 _1518_.Y
rlabel metal1 2004 2162 2076 2178 0 _1479_.gnd
rlabel metal1 2004 1922 2076 1938 0 _1479_.vdd
rlabel metal2 2053 2093 2067 2107 0 _1479_.A
rlabel metal2 2033 2053 2047 2067 0 _1479_.Y
rlabel metal1 2144 2162 2236 2178 0 BUFX2_insert29.gnd
rlabel metal1 2144 1922 2236 1938 0 BUFX2_insert29.vdd
rlabel metal2 2153 2073 2167 2087 0 BUFX2_insert29.A
rlabel metal2 2193 2073 2207 2087 0 BUFX2_insert29.Y
rlabel metal1 2304 2162 2416 2178 0 _796_.gnd
rlabel metal1 2304 1922 2416 1938 0 _796_.vdd
rlabel metal2 2393 2073 2407 2087 0 _796_.A
rlabel metal2 2373 2053 2387 2067 0 _796_.B
rlabel metal2 2333 2053 2347 2067 0 _796_.C
rlabel metal2 2353 2073 2367 2087 0 _796_.Y
rlabel metal1 2404 2162 2496 2178 0 _801_.gnd
rlabel metal1 2404 1922 2496 1938 0 _801_.vdd
rlabel metal2 2473 2033 2487 2047 0 _801_.A
rlabel metal2 2433 2033 2447 2047 0 _801_.B
rlabel metal2 2453 2053 2467 2067 0 _801_.Y
rlabel metal1 2224 2162 2316 2178 0 _795_.gnd
rlabel metal1 2224 1922 2316 1938 0 _795_.vdd
rlabel metal2 2233 2033 2247 2047 0 _795_.A
rlabel metal2 2273 2033 2287 2047 0 _795_.B
rlabel metal2 2253 2053 2267 2067 0 _795_.Y
rlabel metal1 2664 2162 2776 2178 0 _1525_.gnd
rlabel metal1 2664 1922 2776 1938 0 _1525_.vdd
rlabel metal2 2753 2073 2767 2087 0 _1525_.A
rlabel metal2 2733 2053 2747 2067 0 _1525_.B
rlabel metal2 2693 2053 2707 2067 0 _1525_.C
rlabel metal2 2713 2073 2727 2087 0 _1525_.Y
rlabel metal1 2564 2162 2676 2178 0 _802_.gnd
rlabel metal1 2564 1922 2676 1938 0 _802_.vdd
rlabel metal2 2653 2073 2667 2087 0 _802_.A
rlabel metal2 2633 2053 2647 2067 0 _802_.B
rlabel metal2 2593 2053 2607 2067 0 _802_.C
rlabel metal2 2613 2073 2627 2087 0 _802_.Y
rlabel metal1 2484 2162 2576 2178 0 _1524_.gnd
rlabel metal1 2484 1922 2576 1938 0 _1524_.vdd
rlabel metal2 2553 2033 2567 2047 0 _1524_.A
rlabel metal2 2513 2033 2527 2047 0 _1524_.B
rlabel metal2 2533 2053 2547 2067 0 _1524_.Y
rlabel metal1 2764 2162 3016 2178 0 _1595_.gnd
rlabel metal1 2764 1922 3016 1938 0 _1595_.vdd
rlabel metal2 2853 2073 2867 2087 0 _1595_.D
rlabel metal2 2893 2073 2907 2087 0 _1595_.CLK
rlabel metal2 2973 2073 2987 2087 0 _1595_.Q
rlabel metal1 3104 2162 3216 2178 0 _1086_.gnd
rlabel metal1 3104 1922 3216 1938 0 _1086_.vdd
rlabel metal2 3193 2073 3207 2087 0 _1086_.A
rlabel metal2 3173 2053 3187 2067 0 _1086_.B
rlabel metal2 3133 2053 3147 2067 0 _1086_.C
rlabel metal2 3153 2073 3167 2087 0 _1086_.Y
rlabel metal1 3204 2162 3316 2178 0 _1081_.gnd
rlabel metal1 3204 1922 3316 1938 0 _1081_.vdd
rlabel metal2 3293 2073 3307 2087 0 _1081_.A
rlabel metal2 3273 2053 3287 2067 0 _1081_.B
rlabel metal2 3233 2053 3247 2067 0 _1081_.C
rlabel metal2 3253 2073 3267 2087 0 _1081_.Y
rlabel metal1 3004 2162 3116 2178 0 _1080_.gnd
rlabel metal1 3004 1922 3116 1938 0 _1080_.vdd
rlabel metal2 3013 2073 3027 2087 0 _1080_.A
rlabel metal2 3073 2073 3087 2087 0 _1080_.Y
rlabel metal2 3053 2033 3067 2047 0 _1080_.B
rlabel metal1 3384 2162 3496 2178 0 _1079_.gnd
rlabel metal1 3384 1922 3496 1938 0 _1079_.vdd
rlabel metal2 3473 2073 3487 2087 0 _1079_.A
rlabel metal2 3453 2053 3467 2067 0 _1079_.B
rlabel metal2 3413 2053 3427 2067 0 _1079_.C
rlabel metal2 3433 2073 3447 2087 0 _1079_.Y
rlabel metal1 3304 2162 3396 2178 0 _1084_.gnd
rlabel metal1 3304 1922 3396 1938 0 _1084_.vdd
rlabel metal2 3313 2033 3327 2047 0 _1084_.A
rlabel metal2 3353 2033 3367 2047 0 _1084_.B
rlabel metal2 3333 2053 3347 2067 0 _1084_.Y
rlabel metal1 3584 2162 3656 2178 0 _1083_.gnd
rlabel metal1 3584 1922 3656 1938 0 _1083_.vdd
rlabel metal2 3593 2093 3607 2107 0 _1083_.A
rlabel metal2 3613 2053 3627 2067 0 _1083_.Y
rlabel metal1 3644 2162 3756 2178 0 _1087_.gnd
rlabel metal1 3644 1922 3756 1938 0 _1087_.vdd
rlabel metal2 3653 2053 3667 2067 0 _1087_.A
rlabel metal2 3673 2033 3687 2047 0 _1087_.B
rlabel metal2 3693 2053 3707 2067 0 _1087_.C
rlabel metal2 3713 2033 3727 2047 0 _1087_.Y
rlabel metal1 3484 2162 3596 2178 0 _1082_.gnd
rlabel metal1 3484 1922 3596 1938 0 _1082_.vdd
rlabel metal2 3493 2053 3507 2067 0 _1082_.A
rlabel metal2 3513 2033 3527 2047 0 _1082_.B
rlabel metal2 3533 2053 3547 2067 0 _1082_.C
rlabel metal2 3553 2033 3567 2047 0 _1082_.Y
rlabel metal1 3824 2162 3916 2178 0 BUFX2_insert24.gnd
rlabel metal1 3824 1922 3916 1938 0 BUFX2_insert24.vdd
rlabel metal2 3833 2073 3847 2087 0 BUFX2_insert24.A
rlabel metal2 3873 2073 3887 2087 0 BUFX2_insert24.Y
rlabel metal1 3904 2162 4016 2178 0 _1092_.gnd
rlabel metal1 3904 1922 4016 1938 0 _1092_.vdd
rlabel metal2 3913 2073 3927 2087 0 _1092_.A
rlabel metal2 3933 2053 3947 2067 0 _1092_.B
rlabel metal2 3973 2053 3987 2067 0 _1092_.C
rlabel metal2 3953 2073 3967 2087 0 _1092_.Y
rlabel metal1 3744 2162 3836 2178 0 _1142_.gnd
rlabel metal1 3744 1922 3836 1938 0 _1142_.vdd
rlabel metal2 3753 2033 3767 2047 0 _1142_.A
rlabel metal2 3793 2033 3807 2047 0 _1142_.B
rlabel metal2 3773 2053 3787 2067 0 _1142_.Y
rlabel metal1 4004 2162 4096 2178 0 _1096_.gnd
rlabel metal1 4004 1922 4096 1938 0 _1096_.vdd
rlabel metal2 4073 2033 4087 2047 0 _1096_.A
rlabel metal2 4033 2033 4047 2047 0 _1096_.B
rlabel metal2 4053 2053 4067 2067 0 _1096_.Y
rlabel metal1 4084 2162 4176 2178 0 _1090_.gnd
rlabel metal1 4084 1922 4176 1938 0 _1090_.vdd
rlabel metal2 4153 2033 4167 2047 0 _1090_.A
rlabel metal2 4113 2033 4127 2047 0 _1090_.B
rlabel metal2 4133 2053 4147 2067 0 _1090_.Y
rlabel metal1 4164 2162 4256 2178 0 _1088_.gnd
rlabel metal1 4164 1922 4256 1938 0 _1088_.vdd
rlabel metal2 4233 2033 4247 2047 0 _1088_.A
rlabel metal2 4193 2033 4207 2047 0 _1088_.B
rlabel metal2 4213 2053 4227 2067 0 _1088_.Y
rlabel metal1 4244 2162 4356 2178 0 _1107_.gnd
rlabel metal1 4244 1922 4356 1938 0 _1107_.vdd
rlabel metal2 4253 2073 4267 2087 0 _1107_.A
rlabel metal2 4313 2073 4327 2087 0 _1107_.Y
rlabel metal2 4293 2033 4307 2047 0 _1107_.B
rlabel metal1 4344 2162 4456 2178 0 _1145_.gnd
rlabel metal1 4344 1922 4456 1938 0 _1145_.vdd
rlabel metal2 4353 2053 4367 2067 0 _1145_.A
rlabel metal2 4373 2093 4387 2107 0 _1145_.B
rlabel metal2 4393 2053 4407 2067 0 _1145_.C
rlabel metal2 4413 2073 4427 2087 0 _1145_.Y
rlabel metal1 4444 2162 4556 2178 0 _1103_.gnd
rlabel metal1 4444 1922 4556 1938 0 _1103_.vdd
rlabel metal2 4533 2053 4547 2067 0 _1103_.A
rlabel metal2 4513 2093 4527 2107 0 _1103_.B
rlabel metal2 4493 2053 4507 2067 0 _1103_.C
rlabel metal2 4473 2073 4487 2087 0 _1103_.Y
rlabel nsubstratencontact 4764 1932 4764 1932 0 FILL71250x28950.vdd
rlabel metal1 4744 2162 4776 2178 0 FILL71250x28950.gnd
rlabel metal1 4644 2162 4756 2178 0 _1106_.gnd
rlabel metal1 4644 1922 4756 1938 0 _1106_.vdd
rlabel metal2 4653 2053 4667 2067 0 _1106_.A
rlabel metal2 4673 2033 4687 2047 0 _1106_.B
rlabel metal2 4693 2053 4707 2067 0 _1106_.C
rlabel metal2 4713 2033 4727 2047 0 _1106_.Y
rlabel metal1 4544 2162 4656 2178 0 _1099_.gnd
rlabel metal1 4544 1922 4656 1938 0 _1099_.vdd
rlabel metal2 4553 2053 4567 2067 0 _1099_.A
rlabel metal2 4573 2033 4587 2047 0 _1099_.B
rlabel metal2 4593 2053 4607 2067 0 _1099_.C
rlabel metal2 4613 2033 4627 2047 0 _1099_.Y
rlabel metal1 4 2162 256 2178 0 _1564_.gnd
rlabel metal1 4 2402 256 2418 0 _1564_.vdd
rlabel metal2 93 2253 107 2267 0 _1564_.D
rlabel metal2 133 2253 147 2267 0 _1564_.CLK
rlabel metal2 213 2253 227 2267 0 _1564_.Q
rlabel metal1 244 2162 356 2178 0 _1361_.gnd
rlabel metal1 244 2402 356 2418 0 _1361_.vdd
rlabel metal2 253 2253 267 2267 0 _1361_.A
rlabel metal2 273 2273 287 2287 0 _1361_.B
rlabel metal2 313 2273 327 2287 0 _1361_.C
rlabel metal2 293 2253 307 2267 0 _1361_.Y
rlabel metal1 464 2162 556 2178 0 _1608_.gnd
rlabel metal1 464 2402 556 2418 0 _1608_.vdd
rlabel metal2 473 2253 487 2267 0 _1608_.A
rlabel metal2 513 2253 527 2267 0 _1608_.Y
rlabel metal1 344 2162 476 2178 0 _766_.gnd
rlabel metal1 344 2402 476 2418 0 _766_.vdd
rlabel metal2 353 2253 367 2267 0 _766_.A
rlabel metal2 373 2273 387 2287 0 _766_.B
rlabel metal2 433 2253 447 2267 0 _766_.C
rlabel metal2 413 2273 427 2287 0 _766_.D
rlabel metal2 393 2253 407 2267 0 _766_.Y
rlabel metal1 544 2162 636 2178 0 _1352_.gnd
rlabel metal1 544 2402 636 2418 0 _1352_.vdd
rlabel metal2 553 2293 567 2307 0 _1352_.A
rlabel metal2 593 2293 607 2307 0 _1352_.B
rlabel metal2 573 2273 587 2287 0 _1352_.Y
rlabel metal1 764 2162 876 2178 0 _1341_.gnd
rlabel metal1 764 2402 876 2418 0 _1341_.vdd
rlabel metal2 853 2273 867 2287 0 _1341_.A
rlabel metal2 833 2233 847 2247 0 _1341_.B
rlabel metal2 813 2273 827 2287 0 _1341_.C
rlabel metal2 793 2253 807 2267 0 _1341_.Y
rlabel metal1 684 2162 776 2178 0 _1333_.gnd
rlabel metal1 684 2402 776 2418 0 _1333_.vdd
rlabel metal2 733 2253 747 2267 0 _1333_.B
rlabel metal2 693 2253 707 2267 0 _1333_.A
rlabel metal2 713 2233 727 2247 0 _1333_.Y
rlabel metal1 624 2162 696 2178 0 _809_.gnd
rlabel metal1 624 2402 696 2418 0 _809_.vdd
rlabel metal2 673 2233 687 2247 0 _809_.A
rlabel metal2 653 2273 667 2287 0 _809_.Y
rlabel metal1 864 2162 956 2178 0 _1335_.gnd
rlabel metal1 864 2402 956 2418 0 _1335_.vdd
rlabel metal2 913 2253 927 2267 0 _1335_.B
rlabel metal2 873 2253 887 2267 0 _1335_.A
rlabel metal2 893 2233 907 2247 0 _1335_.Y
rlabel metal1 944 2162 1036 2178 0 _1334_.gnd
rlabel metal1 944 2402 1036 2418 0 _1334_.vdd
rlabel metal2 993 2253 1007 2267 0 _1334_.B
rlabel metal2 953 2253 967 2267 0 _1334_.A
rlabel metal2 973 2233 987 2247 0 _1334_.Y
rlabel metal1 1024 2162 1096 2178 0 _864_.gnd
rlabel metal1 1024 2402 1096 2418 0 _864_.vdd
rlabel metal2 1033 2233 1047 2247 0 _864_.A
rlabel metal2 1053 2273 1067 2287 0 _864_.Y
rlabel metal1 1084 2162 1336 2178 0 _1548_.gnd
rlabel metal1 1084 2402 1336 2418 0 _1548_.vdd
rlabel metal2 1233 2253 1247 2267 0 _1548_.D
rlabel metal2 1193 2253 1207 2267 0 _1548_.CLK
rlabel metal2 1113 2253 1127 2267 0 _1548_.Q
rlabel metal1 1324 2162 1436 2178 0 _880_.gnd
rlabel metal1 1324 2402 1436 2418 0 _880_.vdd
rlabel metal2 1333 2253 1347 2267 0 _880_.A
rlabel metal2 1353 2273 1367 2287 0 _880_.B
rlabel metal2 1393 2273 1407 2287 0 _880_.C
rlabel metal2 1373 2253 1387 2267 0 _880_.Y
rlabel metal1 1424 2162 1676 2178 0 _1589_.gnd
rlabel metal1 1424 2402 1676 2418 0 _1589_.vdd
rlabel metal2 1573 2253 1587 2267 0 _1589_.D
rlabel metal2 1533 2253 1547 2267 0 _1589_.CLK
rlabel metal2 1453 2253 1467 2267 0 _1589_.Q
rlabel metal1 1744 2162 1856 2178 0 _1513_.gnd
rlabel metal1 1744 2402 1856 2418 0 _1513_.vdd
rlabel metal2 1833 2273 1847 2287 0 _1513_.A
rlabel metal2 1813 2233 1827 2247 0 _1513_.B
rlabel metal2 1793 2273 1807 2287 0 _1513_.C
rlabel metal2 1773 2253 1787 2267 0 _1513_.Y
rlabel metal1 1664 2162 1756 2178 0 _1512_.gnd
rlabel metal1 1664 2402 1756 2418 0 _1512_.vdd
rlabel metal2 1693 2253 1707 2267 0 _1512_.B
rlabel metal2 1733 2253 1747 2267 0 _1512_.A
rlabel metal2 1713 2233 1727 2247 0 _1512_.Y
rlabel metal1 1844 2162 1916 2178 0 _764_.gnd
rlabel metal1 1844 2402 1916 2418 0 _764_.vdd
rlabel metal2 1853 2273 1867 2287 0 _764_.A
rlabel metal2 1873 2253 1887 2267 0 _764_.Y
rlabel metal1 1984 2162 2196 2178 0 CLKBUF1_insert12.gnd
rlabel metal1 1984 2402 2196 2418 0 CLKBUF1_insert12.vdd
rlabel metal2 2013 2273 2027 2287 0 CLKBUF1_insert12.A
rlabel metal2 2153 2273 2167 2287 0 CLKBUF1_insert12.Y
rlabel metal1 1904 2162 1996 2178 0 _765_.gnd
rlabel metal1 1904 2402 1996 2418 0 _765_.vdd
rlabel metal2 1933 2253 1947 2267 0 _765_.B
rlabel metal2 1973 2253 1987 2267 0 _765_.A
rlabel metal2 1953 2233 1967 2247 0 _765_.Y
rlabel metal1 2284 2162 2536 2178 0 _1592_.gnd
rlabel metal1 2284 2402 2536 2418 0 _1592_.vdd
rlabel metal2 2373 2253 2387 2267 0 _1592_.D
rlabel metal2 2413 2253 2427 2267 0 _1592_.CLK
rlabel metal2 2493 2253 2507 2267 0 _1592_.Q
rlabel metal1 2184 2162 2296 2178 0 _1519_.gnd
rlabel metal1 2184 2402 2296 2418 0 _1519_.vdd
rlabel metal2 2193 2253 2207 2267 0 _1519_.A
rlabel metal2 2213 2273 2227 2287 0 _1519_.B
rlabel metal2 2253 2273 2267 2287 0 _1519_.C
rlabel metal2 2233 2253 2247 2267 0 _1519_.Y
rlabel metal1 2524 2162 2616 2178 0 _1520_.gnd
rlabel metal1 2524 2402 2616 2418 0 _1520_.vdd
rlabel metal2 2593 2293 2607 2307 0 _1520_.A
rlabel metal2 2553 2293 2567 2307 0 _1520_.B
rlabel metal2 2573 2273 2587 2287 0 _1520_.Y
rlabel metal1 2604 2162 2696 2178 0 _799_.gnd
rlabel metal1 2604 2402 2696 2418 0 _799_.vdd
rlabel metal2 2613 2293 2627 2307 0 _799_.A
rlabel metal2 2653 2293 2667 2307 0 _799_.B
rlabel metal2 2633 2273 2647 2287 0 _799_.Y
rlabel metal1 2864 2162 2976 2178 0 _800_.gnd
rlabel metal1 2864 2402 2976 2418 0 _800_.vdd
rlabel metal2 2953 2253 2967 2267 0 _800_.A
rlabel metal2 2933 2273 2947 2287 0 _800_.B
rlabel metal2 2893 2273 2907 2287 0 _800_.C
rlabel metal2 2913 2253 2927 2267 0 _800_.Y
rlabel metal1 2764 2162 2876 2178 0 _798_.gnd
rlabel metal1 2764 2402 2876 2418 0 _798_.vdd
rlabel metal2 2853 2253 2867 2267 0 _798_.A
rlabel metal2 2833 2273 2847 2287 0 _798_.B
rlabel metal2 2793 2273 2807 2287 0 _798_.C
rlabel metal2 2813 2253 2827 2267 0 _798_.Y
rlabel metal1 2684 2162 2776 2178 0 _797_.gnd
rlabel metal1 2684 2402 2776 2418 0 _797_.vdd
rlabel metal2 2693 2293 2707 2307 0 _797_.A
rlabel metal2 2733 2293 2747 2307 0 _797_.B
rlabel metal2 2713 2273 2727 2287 0 _797_.Y
rlabel metal1 2964 2162 3216 2178 0 _1528_.gnd
rlabel metal1 2964 2402 3216 2418 0 _1528_.vdd
rlabel metal2 3053 2253 3067 2267 0 _1528_.D
rlabel metal2 3093 2253 3107 2267 0 _1528_.CLK
rlabel metal2 3173 2253 3187 2267 0 _1528_.Q
rlabel metal1 3204 2162 3316 2178 0 _785_.gnd
rlabel metal1 3204 2402 3316 2418 0 _785_.vdd
rlabel metal2 3213 2253 3227 2267 0 _785_.A
rlabel metal2 3233 2273 3247 2287 0 _785_.B
rlabel metal2 3273 2273 3287 2287 0 _785_.C
rlabel metal2 3253 2253 3267 2267 0 _785_.Y
rlabel metal1 3464 2162 3556 2178 0 _1077_.gnd
rlabel metal1 3464 2402 3556 2418 0 _1077_.vdd
rlabel metal2 3533 2293 3547 2307 0 _1077_.A
rlabel metal2 3493 2293 3507 2307 0 _1077_.B
rlabel metal2 3513 2273 3527 2287 0 _1077_.Y
rlabel metal1 3384 2162 3476 2178 0 _958_.gnd
rlabel metal1 3384 2402 3476 2418 0 _958_.vdd
rlabel metal2 3393 2293 3407 2307 0 _958_.A
rlabel metal2 3433 2293 3447 2307 0 _958_.B
rlabel metal2 3413 2273 3427 2287 0 _958_.Y
rlabel metal1 3304 2162 3396 2178 0 _784_.gnd
rlabel metal1 3304 2402 3396 2418 0 _784_.vdd
rlabel metal2 3313 2293 3327 2307 0 _784_.A
rlabel metal2 3353 2293 3367 2307 0 _784_.B
rlabel metal2 3333 2273 3347 2287 0 _784_.Y
rlabel metal1 3724 2162 3836 2178 0 _1093_.gnd
rlabel metal1 3724 2402 3836 2418 0 _1093_.vdd
rlabel metal2 3733 2253 3747 2267 0 _1093_.A
rlabel metal2 3753 2273 3767 2287 0 _1093_.B
rlabel metal2 3793 2273 3807 2287 0 _1093_.C
rlabel metal2 3773 2253 3787 2267 0 _1093_.Y
rlabel metal1 3664 2162 3736 2178 0 _1483_.gnd
rlabel metal1 3664 2402 3736 2418 0 _1483_.vdd
rlabel metal2 3713 2233 3727 2247 0 _1483_.A
rlabel metal2 3693 2273 3707 2287 0 _1483_.Y
rlabel metal1 3544 2162 3616 2178 0 _934_.gnd
rlabel metal1 3544 2402 3616 2418 0 _934_.vdd
rlabel metal2 3593 2273 3607 2287 0 _934_.A
rlabel metal2 3573 2253 3587 2267 0 _934_.Y
rlabel metal1 3604 2162 3676 2178 0 _899_.gnd
rlabel metal1 3604 2402 3676 2418 0 _899_.vdd
rlabel metal2 3653 2273 3667 2287 0 _899_.A
rlabel metal2 3633 2253 3647 2267 0 _899_.Y
rlabel metal1 3824 2162 3916 2178 0 BUFX2_insert30.gnd
rlabel metal1 3824 2402 3916 2418 0 BUFX2_insert30.vdd
rlabel metal2 3893 2253 3907 2267 0 BUFX2_insert30.A
rlabel metal2 3853 2253 3867 2267 0 BUFX2_insert30.Y
rlabel metal1 3964 2162 4076 2178 0 _1028_.gnd
rlabel metal1 3964 2402 4076 2418 0 _1028_.vdd
rlabel metal2 3973 2253 3987 2267 0 _1028_.A
rlabel metal2 4033 2253 4047 2267 0 _1028_.Y
rlabel metal2 4013 2293 4027 2307 0 _1028_.B
rlabel metal1 3904 2162 3976 2178 0 _860_.gnd
rlabel metal1 3904 2402 3976 2418 0 _860_.vdd
rlabel metal2 3913 2273 3927 2287 0 _860_.A
rlabel metal2 3933 2253 3947 2267 0 _860_.Y
rlabel metal1 4064 2162 4176 2178 0 _1029_.gnd
rlabel metal1 4064 2402 4176 2418 0 _1029_.vdd
rlabel metal2 4153 2253 4167 2267 0 _1029_.A
rlabel metal2 4133 2273 4147 2287 0 _1029_.B
rlabel metal2 4093 2273 4107 2287 0 _1029_.C
rlabel metal2 4113 2253 4127 2267 0 _1029_.Y
rlabel metal1 4264 2162 4376 2178 0 _1104_.gnd
rlabel metal1 4264 2402 4376 2418 0 _1104_.vdd
rlabel metal2 4273 2273 4287 2287 0 _1104_.A
rlabel metal2 4293 2233 4307 2247 0 _1104_.B
rlabel metal2 4313 2273 4327 2287 0 _1104_.C
rlabel metal2 4333 2253 4347 2267 0 _1104_.Y
rlabel metal1 4164 2162 4276 2178 0 _1094_.gnd
rlabel metal1 4164 2402 4276 2418 0 _1094_.vdd
rlabel metal2 4253 2273 4267 2287 0 _1094_.A
rlabel metal2 4233 2293 4247 2307 0 _1094_.B
rlabel metal2 4213 2273 4227 2287 0 _1094_.C
rlabel metal2 4193 2293 4207 2307 0 _1094_.Y
rlabel metal1 4364 2162 4476 2178 0 _1109_.gnd
rlabel metal1 4364 2402 4476 2418 0 _1109_.vdd
rlabel metal2 4453 2253 4467 2267 0 _1109_.A
rlabel metal2 4433 2273 4447 2287 0 _1109_.B
rlabel metal2 4393 2273 4407 2287 0 _1109_.C
rlabel metal2 4413 2253 4427 2267 0 _1109_.Y
rlabel metal1 4464 2162 4576 2178 0 _1105_.gnd
rlabel metal1 4464 2402 4576 2418 0 _1105_.vdd
rlabel metal2 4473 2253 4487 2267 0 _1105_.A
rlabel metal2 4493 2273 4507 2287 0 _1105_.B
rlabel metal2 4533 2273 4547 2287 0 _1105_.C
rlabel metal2 4513 2253 4527 2267 0 _1105_.Y
rlabel metal1 4564 2162 4676 2178 0 _1177_.gnd
rlabel metal1 4564 2402 4676 2418 0 _1177_.vdd
rlabel metal2 4653 2253 4667 2267 0 _1177_.A
rlabel metal2 4633 2273 4647 2287 0 _1177_.B
rlabel metal2 4593 2273 4607 2287 0 _1177_.C
rlabel metal2 4613 2253 4627 2267 0 _1177_.Y
rlabel metal1 4664 2162 4776 2178 0 _1176_.gnd
rlabel metal1 4664 2402 4776 2418 0 _1176_.vdd
rlabel metal2 4673 2273 4687 2287 0 _1176_.A
rlabel metal2 4693 2233 4707 2247 0 _1176_.B
rlabel metal2 4713 2273 4727 2287 0 _1176_.C
rlabel metal2 4733 2253 4747 2267 0 _1176_.Y
rlabel metal1 4 2642 256 2658 0 _1560_.gnd
rlabel metal1 4 2402 256 2418 0 _1560_.vdd
rlabel metal2 93 2553 107 2567 0 _1560_.D
rlabel metal2 133 2553 147 2567 0 _1560_.CLK
rlabel metal2 213 2553 227 2567 0 _1560_.Q
rlabel metal1 244 2642 356 2658 0 _773_.gnd
rlabel metal1 244 2402 356 2418 0 _773_.vdd
rlabel metal2 333 2553 347 2567 0 _773_.A
rlabel metal2 313 2533 327 2547 0 _773_.B
rlabel metal2 273 2533 287 2547 0 _773_.C
rlabel metal2 293 2553 307 2567 0 _773_.Y
rlabel metal1 344 2642 436 2658 0 BUFX2_insert18.gnd
rlabel metal1 344 2402 436 2418 0 BUFX2_insert18.vdd
rlabel metal2 353 2553 367 2567 0 BUFX2_insert18.A
rlabel metal2 393 2553 407 2567 0 BUFX2_insert18.Y
rlabel metal1 504 2642 616 2658 0 _1323_.gnd
rlabel metal1 504 2402 616 2418 0 _1323_.vdd
rlabel metal2 593 2553 607 2567 0 _1323_.A
rlabel metal2 573 2533 587 2547 0 _1323_.B
rlabel metal2 533 2533 547 2547 0 _1323_.C
rlabel metal2 553 2553 567 2567 0 _1323_.Y
rlabel metal1 424 2642 516 2658 0 _1322_.gnd
rlabel metal1 424 2402 516 2418 0 _1322_.vdd
rlabel metal2 433 2513 447 2527 0 _1322_.A
rlabel metal2 473 2513 487 2527 0 _1322_.B
rlabel metal2 453 2533 467 2547 0 _1322_.Y
rlabel metal1 604 2642 696 2658 0 BUFX2_insert19.gnd
rlabel metal1 604 2402 696 2418 0 BUFX2_insert19.vdd
rlabel metal2 613 2553 627 2567 0 BUFX2_insert19.A
rlabel metal2 653 2553 667 2567 0 BUFX2_insert19.Y
rlabel metal1 684 2642 796 2658 0 _1332_.gnd
rlabel metal1 684 2402 796 2418 0 _1332_.vdd
rlabel metal2 773 2553 787 2567 0 _1332_.A
rlabel metal2 753 2533 767 2547 0 _1332_.B
rlabel metal2 713 2533 727 2547 0 _1332_.C
rlabel metal2 733 2553 747 2567 0 _1332_.Y
rlabel metal1 784 2642 876 2658 0 _1324_.gnd
rlabel metal1 784 2402 876 2418 0 _1324_.vdd
rlabel metal2 833 2553 847 2567 0 _1324_.B
rlabel metal2 793 2553 807 2567 0 _1324_.A
rlabel metal2 813 2573 827 2587 0 _1324_.Y
rlabel metal1 864 2642 1116 2658 0 _1531_.gnd
rlabel metal1 864 2402 1116 2418 0 _1531_.vdd
rlabel metal2 953 2553 967 2567 0 _1531_.D
rlabel metal2 993 2553 1007 2567 0 _1531_.CLK
rlabel metal2 1073 2553 1087 2567 0 _1531_.Q
rlabel metal1 1164 2642 1276 2658 0 _808_.gnd
rlabel metal1 1164 2402 1276 2418 0 _808_.vdd
rlabel metal2 1173 2553 1187 2567 0 _808_.A
rlabel metal2 1193 2533 1207 2547 0 _808_.B
rlabel metal2 1233 2533 1247 2547 0 _808_.C
rlabel metal2 1213 2553 1227 2567 0 _808_.Y
rlabel metal1 1324 2642 1416 2658 0 _807_.gnd
rlabel metal1 1324 2402 1416 2418 0 _807_.vdd
rlabel metal2 1333 2513 1347 2527 0 _807_.A
rlabel metal2 1373 2513 1387 2527 0 _807_.B
rlabel metal2 1353 2533 1367 2547 0 _807_.Y
rlabel metal1 1264 2642 1336 2658 0 _854_.gnd
rlabel metal1 1264 2402 1336 2418 0 _854_.vdd
rlabel metal2 1273 2573 1287 2587 0 _854_.A
rlabel metal2 1293 2533 1307 2547 0 _854_.Y
rlabel metal1 1104 2642 1176 2658 0 _806_.gnd
rlabel metal1 1104 2402 1176 2418 0 _806_.vdd
rlabel metal2 1113 2573 1127 2587 0 _806_.A
rlabel metal2 1133 2533 1147 2547 0 _806_.Y
rlabel metal1 1404 2642 1656 2658 0 _1547_.gnd
rlabel metal1 1404 2402 1656 2418 0 _1547_.vdd
rlabel metal2 1553 2553 1567 2567 0 _1547_.D
rlabel metal2 1513 2553 1527 2567 0 _1547_.CLK
rlabel metal2 1433 2553 1447 2567 0 _1547_.Q
rlabel metal1 1744 2642 1996 2658 0 _1588_.gnd
rlabel metal1 1744 2402 1996 2418 0 _1588_.vdd
rlabel metal2 1893 2553 1907 2567 0 _1588_.D
rlabel metal2 1853 2553 1867 2567 0 _1588_.CLK
rlabel metal2 1773 2553 1787 2567 0 _1588_.Q
rlabel metal1 1644 2642 1756 2658 0 _863_.gnd
rlabel metal1 1644 2402 1756 2418 0 _863_.vdd
rlabel metal2 1653 2553 1667 2567 0 _863_.A
rlabel metal2 1673 2533 1687 2547 0 _863_.B
rlabel metal2 1713 2533 1727 2547 0 _863_.C
rlabel metal2 1693 2553 1707 2567 0 _863_.Y
rlabel metal1 1984 2642 2196 2658 0 CLKBUF1_insert14.gnd
rlabel metal1 1984 2402 2196 2418 0 CLKBUF1_insert14.vdd
rlabel metal2 2013 2533 2027 2547 0 CLKBUF1_insert14.A
rlabel metal2 2153 2533 2167 2547 0 CLKBUF1_insert14.Y
rlabel metal1 2184 2642 2436 2658 0 _1593_.gnd
rlabel metal1 2184 2402 2436 2418 0 _1593_.vdd
rlabel metal2 2273 2553 2287 2567 0 _1593_.D
rlabel metal2 2313 2553 2327 2567 0 _1593_.CLK
rlabel metal2 2393 2553 2407 2567 0 _1593_.Q
rlabel metal1 2564 2642 2676 2658 0 _1521_.gnd
rlabel metal1 2564 2402 2676 2418 0 _1521_.vdd
rlabel metal2 2653 2553 2667 2567 0 _1521_.A
rlabel metal2 2633 2533 2647 2547 0 _1521_.B
rlabel metal2 2593 2533 2607 2547 0 _1521_.C
rlabel metal2 2613 2553 2627 2567 0 _1521_.Y
rlabel metal1 2424 2642 2516 2658 0 _1522_.gnd
rlabel metal1 2424 2402 2516 2418 0 _1522_.vdd
rlabel metal2 2493 2513 2507 2527 0 _1522_.A
rlabel metal2 2453 2513 2467 2527 0 _1522_.B
rlabel metal2 2473 2533 2487 2547 0 _1522_.Y
rlabel metal1 2664 2642 2736 2658 0 _959_.gnd
rlabel metal1 2664 2402 2736 2418 0 _959_.vdd
rlabel metal2 2673 2573 2687 2587 0 _959_.A
rlabel metal2 2693 2533 2707 2547 0 _959_.Y
rlabel metal1 2504 2642 2576 2658 0 _859_.gnd
rlabel metal1 2504 2402 2576 2418 0 _859_.vdd
rlabel metal2 2513 2573 2527 2587 0 _859_.A
rlabel metal2 2533 2533 2547 2547 0 _859_.Y
rlabel metal1 2804 2642 2916 2658 0 _791_.gnd
rlabel metal1 2804 2402 2916 2418 0 _791_.vdd
rlabel metal2 2893 2553 2907 2567 0 _791_.A
rlabel metal2 2873 2533 2887 2547 0 _791_.B
rlabel metal2 2833 2533 2847 2547 0 _791_.C
rlabel metal2 2853 2553 2867 2567 0 _791_.Y
rlabel metal1 2724 2642 2816 2658 0 _790_.gnd
rlabel metal1 2724 2402 2816 2418 0 _790_.vdd
rlabel metal2 2793 2513 2807 2527 0 _790_.A
rlabel metal2 2753 2513 2767 2527 0 _790_.B
rlabel metal2 2773 2533 2787 2547 0 _790_.Y
rlabel metal1 2904 2642 3016 2658 0 _960_.gnd
rlabel metal1 2904 2402 3016 2418 0 _960_.vdd
rlabel metal2 2913 2553 2927 2567 0 _960_.A
rlabel metal2 2973 2553 2987 2567 0 _960_.Y
rlabel metal2 2953 2513 2967 2527 0 _960_.B
rlabel metal1 3004 2642 3116 2658 0 _961_.gnd
rlabel metal1 3004 2402 3116 2418 0 _961_.vdd
rlabel metal2 3013 2553 3027 2567 0 _961_.A
rlabel metal2 3033 2533 3047 2547 0 _961_.B
rlabel metal2 3073 2533 3087 2547 0 _961_.C
rlabel metal2 3053 2553 3067 2567 0 _961_.Y
rlabel metal1 3104 2642 3196 2658 0 _935_.gnd
rlabel metal1 3104 2402 3196 2418 0 _935_.vdd
rlabel metal2 3173 2513 3187 2527 0 _935_.A
rlabel metal2 3133 2513 3147 2527 0 _935_.B
rlabel metal2 3153 2533 3167 2547 0 _935_.Y
rlabel metal1 3184 2642 3296 2658 0 _1015_.gnd
rlabel metal1 3184 2402 3296 2418 0 _1015_.vdd
rlabel metal2 3193 2553 3207 2567 0 _1015_.A
rlabel metal2 3253 2553 3267 2567 0 _1015_.Y
rlabel metal2 3233 2513 3247 2527 0 _1015_.B
rlabel metal1 3444 2642 3536 2658 0 _1014_.gnd
rlabel metal1 3444 2402 3536 2418 0 _1014_.vdd
rlabel metal2 3453 2513 3467 2527 0 _1014_.A
rlabel metal2 3493 2513 3507 2527 0 _1014_.B
rlabel metal2 3473 2533 3487 2547 0 _1014_.Y
rlabel metal1 3384 2642 3456 2658 0 _965_.gnd
rlabel metal1 3384 2402 3456 2418 0 _965_.vdd
rlabel metal2 3393 2573 3407 2587 0 _965_.A
rlabel metal2 3413 2533 3427 2547 0 _965_.Y
rlabel metal1 3284 2642 3396 2658 0 _964_.gnd
rlabel metal1 3284 2402 3396 2418 0 _964_.vdd
rlabel metal2 3373 2533 3387 2547 0 _964_.A
rlabel metal2 3353 2513 3367 2527 0 _964_.B
rlabel metal2 3333 2533 3347 2547 0 _964_.C
rlabel metal2 3313 2513 3327 2527 0 _964_.Y
rlabel metal1 3624 2642 3716 2658 0 BUFX2_insert23.gnd
rlabel metal1 3624 2402 3716 2418 0 BUFX2_insert23.vdd
rlabel metal2 3633 2553 3647 2567 0 BUFX2_insert23.A
rlabel metal2 3673 2553 3687 2567 0 BUFX2_insert23.Y
rlabel metal1 3704 2642 3776 2658 0 _900_.gnd
rlabel metal1 3704 2402 3776 2418 0 _900_.vdd
rlabel metal2 3713 2573 3727 2587 0 _900_.A
rlabel metal2 3733 2533 3747 2547 0 _900_.Y
rlabel metal1 3524 2642 3636 2658 0 _1017_.gnd
rlabel metal1 3524 2402 3636 2418 0 _1017_.vdd
rlabel metal2 3533 2553 3547 2567 0 _1017_.A
rlabel metal2 3593 2553 3607 2567 0 _1017_.Y
rlabel metal2 3573 2513 3587 2527 0 _1017_.B
rlabel metal1 3984 2642 4076 2658 0 _1030_.gnd
rlabel metal1 3984 2402 4076 2418 0 _1030_.vdd
rlabel metal2 4053 2513 4067 2527 0 _1030_.A
rlabel metal2 4013 2513 4027 2527 0 _1030_.B
rlabel metal2 4033 2533 4047 2547 0 _1030_.Y
rlabel metal1 3864 2642 3996 2658 0 _1101_.gnd
rlabel metal1 3864 2402 3996 2418 0 _1101_.vdd
rlabel metal2 3973 2553 3987 2567 0 _1101_.A
rlabel metal2 3953 2533 3967 2547 0 _1101_.B
rlabel metal2 3893 2553 3907 2567 0 _1101_.C
rlabel metal2 3913 2533 3927 2547 0 _1101_.D
rlabel metal2 3933 2553 3947 2567 0 _1101_.Y
rlabel metal1 3764 2642 3876 2658 0 _1034_.gnd
rlabel metal1 3764 2402 3876 2418 0 _1034_.vdd
rlabel metal2 3853 2553 3867 2567 0 _1034_.A
rlabel metal2 3793 2553 3807 2567 0 _1034_.Y
rlabel metal2 3813 2513 3827 2527 0 _1034_.B
rlabel metal1 4144 2642 4256 2658 0 _1102_.gnd
rlabel metal1 4144 2402 4256 2418 0 _1102_.vdd
rlabel metal2 4153 2553 4167 2567 0 _1102_.A
rlabel metal2 4173 2533 4187 2547 0 _1102_.B
rlabel metal2 4213 2533 4227 2547 0 _1102_.C
rlabel metal2 4193 2553 4207 2567 0 _1102_.Y
rlabel metal1 4244 2642 4336 2658 0 _1035_.gnd
rlabel metal1 4244 2402 4336 2418 0 _1035_.vdd
rlabel metal2 4253 2513 4267 2527 0 _1035_.A
rlabel metal2 4293 2513 4307 2527 0 _1035_.B
rlabel metal2 4273 2533 4287 2547 0 _1035_.Y
rlabel metal1 4064 2642 4156 2658 0 _1027_.gnd
rlabel metal1 4064 2402 4156 2418 0 _1027_.vdd
rlabel metal2 4133 2513 4147 2527 0 _1027_.A
rlabel metal2 4093 2513 4107 2527 0 _1027_.B
rlabel metal2 4113 2533 4127 2547 0 _1027_.Y
rlabel metal1 4524 2642 4636 2658 0 _1114_.gnd
rlabel metal1 4524 2402 4636 2418 0 _1114_.vdd
rlabel metal2 4533 2533 4547 2547 0 _1114_.A
rlabel metal2 4553 2573 4567 2587 0 _1114_.B
rlabel metal2 4573 2533 4587 2547 0 _1114_.C
rlabel metal2 4593 2553 4607 2567 0 _1114_.Y
rlabel metal1 4424 2642 4536 2658 0 _1110_.gnd
rlabel metal1 4424 2402 4536 2418 0 _1110_.vdd
rlabel metal2 4513 2533 4527 2547 0 _1110_.A
rlabel metal2 4493 2513 4507 2527 0 _1110_.B
rlabel metal2 4473 2533 4487 2547 0 _1110_.C
rlabel metal2 4453 2513 4467 2527 0 _1110_.Y
rlabel metal1 4324 2642 4436 2658 0 _1100_.gnd
rlabel metal1 4324 2402 4436 2418 0 _1100_.vdd
rlabel metal2 4413 2533 4427 2547 0 _1100_.A
rlabel metal2 4393 2513 4407 2527 0 _1100_.B
rlabel metal2 4373 2533 4387 2547 0 _1100_.C
rlabel metal2 4353 2513 4367 2527 0 _1100_.Y
rlabel nsubstratencontact 4764 2412 4764 2412 0 FILL71250x36150.vdd
rlabel metal1 4744 2642 4776 2658 0 FILL71250x36150.gnd
rlabel nsubstratencontact 4744 2412 4744 2412 0 FILL70950x36150.vdd
rlabel metal1 4724 2642 4756 2658 0 FILL70950x36150.gnd
rlabel metal1 4624 2642 4736 2658 0 _1108_.gnd
rlabel metal1 4624 2402 4736 2418 0 _1108_.vdd
rlabel metal2 4713 2533 4727 2547 0 _1108_.A
rlabel metal2 4693 2513 4707 2527 0 _1108_.B
rlabel metal2 4673 2533 4687 2547 0 _1108_.C
rlabel metal2 4653 2513 4667 2527 0 _1108_.Y
rlabel metal1 4 2642 256 2658 0 _1561_.gnd
rlabel metal1 4 2882 256 2898 0 _1561_.vdd
rlabel metal2 93 2733 107 2747 0 _1561_.D
rlabel metal2 133 2733 147 2747 0 _1561_.CLK
rlabel metal2 213 2733 227 2747 0 _1561_.Q
rlabel metal1 244 2642 376 2658 0 _772_.gnd
rlabel metal1 244 2882 376 2898 0 _772_.vdd
rlabel metal2 353 2733 367 2747 0 _772_.A
rlabel metal2 333 2753 347 2767 0 _772_.B
rlabel metal2 273 2733 287 2747 0 _772_.C
rlabel metal2 293 2753 307 2767 0 _772_.D
rlabel metal2 313 2733 327 2747 0 _772_.Y
rlabel metal1 444 2642 556 2658 0 _1331_.gnd
rlabel metal1 444 2882 556 2898 0 _1331_.vdd
rlabel metal2 533 2733 547 2747 0 _1331_.A
rlabel metal2 513 2753 527 2767 0 _1331_.B
rlabel metal2 473 2753 487 2767 0 _1331_.C
rlabel metal2 493 2733 507 2747 0 _1331_.Y
rlabel metal1 364 2642 456 2658 0 _1330_.gnd
rlabel metal1 364 2882 456 2898 0 _1330_.vdd
rlabel metal2 373 2773 387 2787 0 _1330_.A
rlabel metal2 413 2773 427 2787 0 _1330_.B
rlabel metal2 393 2753 407 2767 0 _1330_.Y
rlabel metal1 544 2642 636 2658 0 BUFX2_insert26.gnd
rlabel metal1 544 2882 636 2898 0 BUFX2_insert26.vdd
rlabel metal2 613 2733 627 2747 0 BUFX2_insert26.A
rlabel metal2 573 2733 587 2747 0 BUFX2_insert26.Y
rlabel metal1 704 2642 816 2658 0 _1328_.gnd
rlabel metal1 704 2882 816 2898 0 _1328_.vdd
rlabel metal2 793 2733 807 2747 0 _1328_.A
rlabel metal2 773 2753 787 2767 0 _1328_.B
rlabel metal2 733 2753 747 2767 0 _1328_.C
rlabel metal2 753 2733 767 2747 0 _1328_.Y
rlabel metal1 624 2642 716 2658 0 _1329_.gnd
rlabel metal1 624 2882 716 2898 0 _1329_.vdd
rlabel metal2 633 2773 647 2787 0 _1329_.A
rlabel metal2 673 2773 687 2787 0 _1329_.B
rlabel metal2 653 2753 667 2767 0 _1329_.Y
rlabel metal1 884 2642 976 2658 0 _1327_.gnd
rlabel metal1 884 2882 976 2898 0 _1327_.vdd
rlabel metal2 953 2773 967 2787 0 _1327_.A
rlabel metal2 913 2773 927 2787 0 _1327_.B
rlabel metal2 933 2753 947 2767 0 _1327_.Y
rlabel metal1 1024 2642 1116 2658 0 _1321_.gnd
rlabel metal1 1024 2882 1116 2898 0 _1321_.vdd
rlabel metal2 1093 2773 1107 2787 0 _1321_.A
rlabel metal2 1053 2773 1067 2787 0 _1321_.B
rlabel metal2 1073 2753 1087 2767 0 _1321_.Y
rlabel metal1 804 2642 896 2658 0 _1326_.gnd
rlabel metal1 804 2882 896 2898 0 _1326_.vdd
rlabel metal2 833 2733 847 2747 0 _1326_.B
rlabel metal2 873 2733 887 2747 0 _1326_.A
rlabel metal2 853 2713 867 2727 0 _1326_.Y
rlabel metal1 964 2642 1036 2658 0 _1319_.gnd
rlabel metal1 964 2882 1036 2898 0 _1319_.vdd
rlabel metal2 973 2713 987 2727 0 _1319_.A
rlabel metal2 993 2753 1007 2767 0 _1319_.Y
rlabel metal1 1184 2642 1276 2658 0 BUFX2_insert2.gnd
rlabel metal1 1184 2882 1276 2898 0 BUFX2_insert2.vdd
rlabel metal2 1253 2733 1267 2747 0 BUFX2_insert2.A
rlabel metal2 1213 2733 1227 2747 0 BUFX2_insert2.Y
rlabel metal1 1264 2642 1516 2658 0 _1584_.gnd
rlabel metal1 1264 2882 1516 2898 0 _1584_.vdd
rlabel metal2 1353 2733 1367 2747 0 _1584_.D
rlabel metal2 1393 2733 1407 2747 0 _1584_.CLK
rlabel metal2 1473 2733 1487 2747 0 _1584_.Q
rlabel metal1 1104 2642 1196 2658 0 _1325_.gnd
rlabel metal1 1104 2882 1196 2898 0 _1325_.vdd
rlabel metal2 1153 2733 1167 2747 0 _1325_.B
rlabel metal2 1113 2733 1127 2747 0 _1325_.A
rlabel metal2 1133 2713 1147 2727 0 _1325_.Y
rlabel metal1 1584 2642 1696 2658 0 _1502_.gnd
rlabel metal1 1584 2882 1696 2898 0 _1502_.vdd
rlabel metal2 1673 2733 1687 2747 0 _1502_.A
rlabel metal2 1653 2753 1667 2767 0 _1502_.B
rlabel metal2 1613 2753 1627 2767 0 _1502_.C
rlabel metal2 1633 2733 1647 2747 0 _1502_.Y
rlabel metal1 1504 2642 1596 2658 0 _879_.gnd
rlabel metal1 1504 2882 1596 2898 0 _879_.vdd
rlabel metal2 1513 2773 1527 2787 0 _879_.A
rlabel metal2 1553 2773 1567 2787 0 _879_.B
rlabel metal2 1533 2753 1547 2767 0 _879_.Y
rlabel metal1 1684 2642 1796 2658 0 _1503_.gnd
rlabel metal1 1684 2882 1796 2898 0 _1503_.vdd
rlabel metal2 1773 2733 1787 2747 0 _1503_.A
rlabel metal2 1753 2753 1767 2767 0 _1503_.B
rlabel metal2 1713 2753 1727 2767 0 _1503_.C
rlabel metal2 1733 2733 1747 2747 0 _1503_.Y
rlabel metal1 1864 2642 1976 2658 0 _1511_.gnd
rlabel metal1 1864 2882 1976 2898 0 _1511_.vdd
rlabel metal2 1953 2753 1967 2767 0 _1511_.A
rlabel metal2 1933 2713 1947 2727 0 _1511_.B
rlabel metal2 1913 2753 1927 2767 0 _1511_.C
rlabel metal2 1893 2733 1907 2747 0 _1511_.Y
rlabel metal1 1784 2642 1876 2658 0 _1510_.gnd
rlabel metal1 1784 2882 1876 2898 0 _1510_.vdd
rlabel metal2 1813 2733 1827 2747 0 _1510_.B
rlabel metal2 1853 2733 1867 2747 0 _1510_.A
rlabel metal2 1833 2713 1847 2727 0 _1510_.Y
rlabel metal1 1964 2642 2056 2658 0 BUFX2_insert28.gnd
rlabel metal1 1964 2882 2056 2898 0 BUFX2_insert28.vdd
rlabel metal2 2033 2733 2047 2747 0 BUFX2_insert28.A
rlabel metal2 1993 2733 2007 2747 0 BUFX2_insert28.Y
rlabel metal1 2044 2642 2156 2658 0 _862_.gnd
rlabel metal1 2044 2882 2156 2898 0 _862_.vdd
rlabel metal2 2133 2753 2147 2767 0 _862_.A
rlabel metal2 2113 2773 2127 2787 0 _862_.B
rlabel metal2 2093 2753 2107 2767 0 _862_.C
rlabel metal2 2073 2773 2087 2787 0 _862_.Y
rlabel metal1 2144 2642 2236 2658 0 BUFX2_insert27.gnd
rlabel metal1 2144 2882 2236 2898 0 BUFX2_insert27.vdd
rlabel metal2 2153 2733 2167 2747 0 BUFX2_insert27.A
rlabel metal2 2193 2733 2207 2747 0 BUFX2_insert27.Y
rlabel metal1 2224 2642 2476 2658 0 _1594_.gnd
rlabel metal1 2224 2882 2476 2898 0 _1594_.vdd
rlabel metal2 2313 2733 2327 2747 0 _1594_.D
rlabel metal2 2353 2733 2367 2747 0 _1594_.CLK
rlabel metal2 2433 2733 2447 2747 0 _1594_.Q
rlabel metal1 2464 2642 2576 2658 0 _1523_.gnd
rlabel metal1 2464 2882 2576 2898 0 _1523_.vdd
rlabel metal2 2553 2733 2567 2747 0 _1523_.A
rlabel metal2 2533 2753 2547 2767 0 _1523_.B
rlabel metal2 2493 2753 2507 2767 0 _1523_.C
rlabel metal2 2513 2733 2527 2747 0 _1523_.Y
rlabel metal1 2564 2642 2676 2658 0 _861_.gnd
rlabel metal1 2564 2882 2676 2898 0 _861_.vdd
rlabel metal2 2653 2733 2667 2747 0 _861_.A
rlabel metal2 2633 2753 2647 2767 0 _861_.B
rlabel metal2 2593 2753 2607 2767 0 _861_.C
rlabel metal2 2613 2733 2627 2747 0 _861_.Y
rlabel metal1 2664 2642 2776 2658 0 _794_.gnd
rlabel metal1 2664 2882 2776 2898 0 _794_.vdd
rlabel metal2 2673 2733 2687 2747 0 _794_.A
rlabel metal2 2693 2753 2707 2767 0 _794_.B
rlabel metal2 2733 2753 2747 2767 0 _794_.C
rlabel metal2 2713 2733 2727 2747 0 _794_.Y
rlabel metal1 2924 2642 3036 2658 0 _937_.gnd
rlabel metal1 2924 2882 3036 2898 0 _937_.vdd
rlabel metal2 2933 2733 2947 2747 0 _937_.A
rlabel metal2 2953 2753 2967 2767 0 _937_.B
rlabel metal2 2993 2753 3007 2767 0 _937_.C
rlabel metal2 2973 2733 2987 2747 0 _937_.Y
rlabel metal1 2844 2642 2936 2658 0 _882_.gnd
rlabel metal1 2844 2882 2936 2898 0 _882_.vdd
rlabel metal2 2853 2773 2867 2787 0 _882_.A
rlabel metal2 2893 2773 2907 2787 0 _882_.B
rlabel metal2 2873 2753 2887 2767 0 _882_.Y
rlabel metal1 2764 2642 2856 2658 0 _793_.gnd
rlabel metal1 2764 2882 2856 2898 0 _793_.vdd
rlabel metal2 2773 2773 2787 2787 0 _793_.A
rlabel metal2 2813 2773 2827 2787 0 _793_.B
rlabel metal2 2793 2753 2807 2767 0 _793_.Y
rlabel metal1 3204 2642 3316 2658 0 _967_.gnd
rlabel metal1 3204 2882 3316 2898 0 _967_.vdd
rlabel metal2 3293 2733 3307 2747 0 _967_.A
rlabel metal2 3273 2753 3287 2767 0 _967_.B
rlabel metal2 3233 2753 3247 2767 0 _967_.C
rlabel metal2 3253 2733 3267 2747 0 _967_.Y
rlabel metal1 3024 2642 3136 2658 0 _936_.gnd
rlabel metal1 3024 2882 3136 2898 0 _936_.vdd
rlabel metal2 3033 2733 3047 2747 0 _936_.A
rlabel metal2 3053 2753 3067 2767 0 _936_.B
rlabel metal2 3093 2753 3107 2767 0 _936_.C
rlabel metal2 3073 2733 3087 2747 0 _936_.Y
rlabel metal1 3124 2642 3216 2658 0 _933_.gnd
rlabel metal1 3124 2882 3216 2898 0 _933_.vdd
rlabel metal2 3133 2773 3147 2787 0 _933_.A
rlabel metal2 3173 2773 3187 2787 0 _933_.B
rlabel metal2 3153 2753 3167 2767 0 _933_.Y
rlabel metal1 3304 2642 3396 2658 0 _966_.gnd
rlabel metal1 3304 2882 3396 2898 0 _966_.vdd
rlabel metal2 3373 2773 3387 2787 0 _966_.A
rlabel metal2 3333 2773 3347 2787 0 _966_.B
rlabel metal2 3353 2753 3367 2767 0 _966_.Y
rlabel metal1 3384 2642 3496 2658 0 _968_.gnd
rlabel metal1 3384 2882 3496 2898 0 _968_.vdd
rlabel metal2 3393 2753 3407 2767 0 _968_.A
rlabel metal2 3413 2773 3427 2787 0 _968_.B
rlabel metal2 3433 2753 3447 2767 0 _968_.C
rlabel metal2 3453 2773 3467 2787 0 _968_.Y
rlabel metal1 3584 2642 3696 2658 0 _1016_.gnd
rlabel metal1 3584 2882 3696 2898 0 _1016_.vdd
rlabel metal2 3593 2733 3607 2747 0 _1016_.A
rlabel metal2 3613 2753 3627 2767 0 _1016_.B
rlabel metal2 3653 2753 3667 2767 0 _1016_.C
rlabel metal2 3633 2733 3647 2747 0 _1016_.Y
rlabel metal1 3484 2642 3596 2658 0 _963_.gnd
rlabel metal1 3484 2882 3596 2898 0 _963_.vdd
rlabel metal2 3573 2733 3587 2747 0 _963_.A
rlabel metal2 3553 2753 3567 2767 0 _963_.B
rlabel metal2 3513 2753 3527 2767 0 _963_.C
rlabel metal2 3533 2733 3547 2747 0 _963_.Y
rlabel metal1 3684 2642 3776 2658 0 _1021_.gnd
rlabel metal1 3684 2882 3776 2898 0 _1021_.vdd
rlabel metal2 3753 2773 3767 2787 0 _1021_.A
rlabel metal2 3713 2773 3727 2787 0 _1021_.B
rlabel metal2 3733 2753 3747 2767 0 _1021_.Y
rlabel metal1 3764 2642 3876 2658 0 _1018_.gnd
rlabel metal1 3764 2882 3876 2898 0 _1018_.vdd
rlabel metal2 3853 2733 3867 2747 0 _1018_.A
rlabel metal2 3833 2753 3847 2767 0 _1018_.B
rlabel metal2 3793 2753 3807 2767 0 _1018_.C
rlabel metal2 3813 2733 3827 2747 0 _1018_.Y
rlabel metal1 3964 2642 4036 2658 0 _1020_.gnd
rlabel metal1 3964 2882 4036 2898 0 _1020_.vdd
rlabel metal2 3973 2713 3987 2727 0 _1020_.A
rlabel metal2 3993 2753 4007 2767 0 _1020_.Y
rlabel metal1 3864 2642 3976 2658 0 _1019_.gnd
rlabel metal1 3864 2882 3976 2898 0 _1019_.vdd
rlabel metal2 3873 2753 3887 2767 0 _1019_.A
rlabel metal2 3893 2773 3907 2787 0 _1019_.B
rlabel metal2 3913 2753 3927 2767 0 _1019_.C
rlabel metal2 3933 2773 3947 2787 0 _1019_.Y
rlabel metal1 4244 2642 4356 2658 0 _1036_.gnd
rlabel metal1 4244 2882 4356 2898 0 _1036_.vdd
rlabel metal2 4253 2733 4267 2747 0 _1036_.A
rlabel metal2 4273 2753 4287 2767 0 _1036_.B
rlabel metal2 4313 2753 4327 2767 0 _1036_.C
rlabel metal2 4293 2733 4307 2747 0 _1036_.Y
rlabel metal1 4144 2642 4256 2658 0 _1031_.gnd
rlabel metal1 4144 2882 4256 2898 0 _1031_.vdd
rlabel metal2 4153 2753 4167 2767 0 _1031_.A
rlabel metal2 4173 2773 4187 2787 0 _1031_.B
rlabel metal2 4193 2753 4207 2767 0 _1031_.C
rlabel metal2 4213 2773 4227 2787 0 _1031_.Y
rlabel metal1 4024 2642 4156 2658 0 _1039_.gnd
rlabel metal1 4024 2882 4156 2898 0 _1039_.vdd
rlabel metal2 4133 2733 4147 2747 0 _1039_.A
rlabel metal2 4113 2753 4127 2767 0 _1039_.B
rlabel metal2 4053 2733 4067 2747 0 _1039_.C
rlabel metal2 4073 2753 4087 2767 0 _1039_.D
rlabel metal2 4093 2733 4107 2747 0 _1039_.Y
rlabel metal1 4444 2642 4576 2658 0 _1089_.gnd
rlabel metal1 4444 2882 4576 2898 0 _1089_.vdd
rlabel metal2 4453 2733 4467 2747 0 _1089_.A
rlabel metal2 4473 2753 4487 2767 0 _1089_.B
rlabel metal2 4533 2733 4547 2747 0 _1089_.C
rlabel metal2 4513 2753 4527 2767 0 _1089_.D
rlabel metal2 4493 2733 4507 2747 0 _1089_.Y
rlabel metal1 4344 2642 4456 2658 0 _972_.gnd
rlabel metal1 4344 2882 4456 2898 0 _972_.vdd
rlabel metal2 4353 2733 4367 2747 0 _972_.A
rlabel metal2 4413 2733 4427 2747 0 _972_.Y
rlabel metal2 4393 2773 4407 2787 0 _972_.B
rlabel nsubstratencontact 4756 2888 4756 2888 0 FILL71250x39750.vdd
rlabel metal1 4744 2642 4776 2658 0 FILL71250x39750.gnd
rlabel nsubstratencontact 4736 2888 4736 2888 0 FILL70950x39750.vdd
rlabel metal1 4724 2642 4756 2658 0 FILL70950x39750.gnd
rlabel metal1 4624 2642 4736 2658 0 _1115_.gnd
rlabel metal1 4624 2882 4736 2898 0 _1115_.vdd
rlabel metal2 4633 2753 4647 2767 0 _1115_.A
rlabel metal2 4653 2713 4667 2727 0 _1115_.B
rlabel metal2 4673 2753 4687 2767 0 _1115_.C
rlabel metal2 4693 2733 4707 2747 0 _1115_.Y
rlabel metal1 4564 2642 4636 2658 0 _1033_.gnd
rlabel metal1 4564 2882 4636 2898 0 _1033_.vdd
rlabel metal2 4573 2713 4587 2727 0 _1033_.A
rlabel metal2 4593 2753 4607 2767 0 _1033_.Y
rlabel metal1 4 3122 256 3138 0 _1596_.gnd
rlabel metal1 4 2882 256 2898 0 _1596_.vdd
rlabel metal2 93 3033 107 3047 0 _1596_.D
rlabel metal2 133 3033 147 3047 0 _1596_.CLK
rlabel metal2 213 3033 227 3047 0 _1596_.Q
rlabel metal1 4 3122 256 3138 0 _1567_.gnd
rlabel metal1 4 3362 256 3378 0 _1567_.vdd
rlabel metal2 93 3213 107 3227 0 _1567_.D
rlabel metal2 133 3213 147 3227 0 _1567_.CLK
rlabel metal2 213 3213 227 3227 0 _1567_.Q
rlabel metal1 244 3122 356 3138 0 _782_.gnd
rlabel metal1 244 2882 356 2898 0 _782_.vdd
rlabel metal2 333 3033 347 3047 0 _782_.A
rlabel metal2 313 3013 327 3027 0 _782_.B
rlabel metal2 273 3013 287 3027 0 _782_.C
rlabel metal2 293 3033 307 3047 0 _782_.Y
rlabel metal1 244 3122 376 3138 0 _781_.gnd
rlabel metal1 244 3362 376 3378 0 _781_.vdd
rlabel metal2 353 3213 367 3227 0 _781_.A
rlabel metal2 333 3233 347 3247 0 _781_.B
rlabel metal2 273 3213 287 3227 0 _781_.C
rlabel metal2 293 3233 307 3247 0 _781_.D
rlabel metal2 313 3213 327 3227 0 _781_.Y
rlabel metal1 424 3122 676 3138 0 _1566_.gnd
rlabel metal1 424 2882 676 2898 0 _1566_.vdd
rlabel metal2 573 3033 587 3047 0 _1566_.D
rlabel metal2 533 3033 547 3047 0 _1566_.CLK
rlabel metal2 453 3033 467 3047 0 _1566_.Q
rlabel metal1 444 3122 556 3138 0 _1392_.gnd
rlabel metal1 444 3362 556 3378 0 _1392_.vdd
rlabel metal2 453 3213 467 3227 0 _1392_.A
rlabel metal2 473 3233 487 3247 0 _1392_.B
rlabel metal2 513 3233 527 3247 0 _1392_.C
rlabel metal2 493 3213 507 3227 0 _1392_.Y
rlabel metal1 364 3122 456 3138 0 _1391_.gnd
rlabel metal1 364 3362 456 3378 0 _1391_.vdd
rlabel metal2 373 3253 387 3267 0 _1391_.A
rlabel metal2 413 3253 427 3267 0 _1391_.B
rlabel metal2 393 3233 407 3247 0 _1391_.Y
rlabel metal1 344 3122 436 3138 0 _1371_.gnd
rlabel metal1 344 2882 436 2898 0 _1371_.vdd
rlabel metal2 413 2993 427 3007 0 _1371_.A
rlabel metal2 373 2993 387 3007 0 _1371_.B
rlabel metal2 393 3013 407 3027 0 _1371_.Y
rlabel metal1 784 3122 996 3138 0 CLKBUF1_insert10.gnd
rlabel metal1 784 3362 996 3378 0 CLKBUF1_insert10.vdd
rlabel metal2 953 3233 967 3247 0 CLKBUF1_insert10.A
rlabel metal2 813 3233 827 3247 0 CLKBUF1_insert10.Y
rlabel metal1 664 3122 916 3138 0 _1546_.gnd
rlabel metal1 664 2882 916 2898 0 _1546_.vdd
rlabel metal2 753 3033 767 3047 0 _1546_.D
rlabel metal2 793 3033 807 3047 0 _1546_.CLK
rlabel metal2 873 3033 887 3047 0 _1546_.Q
rlabel metal1 544 3122 656 3138 0 _1382_.gnd
rlabel metal1 544 3362 656 3378 0 _1382_.vdd
rlabel metal2 553 3213 567 3227 0 _1382_.A
rlabel metal2 573 3233 587 3247 0 _1382_.B
rlabel metal2 613 3233 627 3247 0 _1382_.C
rlabel metal2 593 3213 607 3227 0 _1382_.Y
rlabel metal1 644 3122 736 3138 0 _1390_.gnd
rlabel metal1 644 3362 736 3378 0 _1390_.vdd
rlabel metal2 713 3253 727 3267 0 _1390_.A
rlabel metal2 673 3253 687 3267 0 _1390_.B
rlabel metal2 693 3233 707 3247 0 _1390_.Y
rlabel metal1 724 3122 796 3138 0 _1345_.gnd
rlabel metal1 724 3362 796 3378 0 _1345_.vdd
rlabel metal2 733 3193 747 3207 0 _1345_.A
rlabel metal2 753 3233 767 3247 0 _1345_.Y
rlabel metal1 984 3122 1196 3138 0 CLKBUF1_insert11.gnd
rlabel metal1 984 3362 1196 3378 0 CLKBUF1_insert11.vdd
rlabel metal2 1013 3233 1027 3247 0 CLKBUF1_insert11.A
rlabel metal2 1153 3233 1167 3247 0 CLKBUF1_insert11.Y
rlabel metal1 1044 3122 1136 3138 0 _1320_.gnd
rlabel metal1 1044 2882 1136 2898 0 _1320_.vdd
rlabel metal2 1113 2993 1127 3007 0 _1320_.A
rlabel metal2 1073 2993 1087 3007 0 _1320_.B
rlabel metal2 1093 3013 1107 3027 0 _1320_.Y
rlabel metal1 964 3122 1056 3138 0 _1318_.gnd
rlabel metal1 964 2882 1056 2898 0 _1318_.vdd
rlabel metal2 993 3033 1007 3047 0 _1318_.B
rlabel metal2 1033 3033 1047 3047 0 _1318_.A
rlabel metal2 1013 3053 1027 3067 0 _1318_.Y
rlabel metal1 904 3122 976 3138 0 _851_.gnd
rlabel metal1 904 2882 976 2898 0 _851_.vdd
rlabel metal2 913 3053 927 3067 0 _851_.A
rlabel metal2 933 3013 947 3027 0 _851_.Y
rlabel metal1 1324 3122 1576 3138 0 _1591_.gnd
rlabel metal1 1324 2882 1576 2898 0 _1591_.vdd
rlabel metal2 1413 3033 1427 3047 0 _1591_.D
rlabel metal2 1453 3033 1467 3047 0 _1591_.CLK
rlabel metal2 1533 3033 1547 3047 0 _1591_.Q
rlabel metal1 1244 3122 1496 3138 0 _1530_.gnd
rlabel metal1 1244 3362 1496 3378 0 _1530_.vdd
rlabel metal2 1393 3213 1407 3227 0 _1530_.D
rlabel metal2 1353 3213 1367 3227 0 _1530_.CLK
rlabel metal2 1273 3213 1287 3227 0 _1530_.Q
rlabel metal1 1124 3122 1236 3138 0 _853_.gnd
rlabel metal1 1124 2882 1236 2898 0 _853_.vdd
rlabel metal2 1133 3033 1147 3047 0 _853_.A
rlabel metal2 1153 3013 1167 3027 0 _853_.B
rlabel metal2 1193 3013 1207 3027 0 _853_.C
rlabel metal2 1173 3033 1187 3047 0 _853_.Y
rlabel metal1 1224 3122 1336 3138 0 _1517_.gnd
rlabel metal1 1224 2882 1336 2898 0 _1517_.vdd
rlabel metal2 1233 3013 1247 3027 0 _1517_.A
rlabel metal2 1253 3053 1267 3067 0 _1517_.B
rlabel metal2 1273 3013 1287 3027 0 _1517_.C
rlabel metal2 1293 3033 1307 3047 0 _1517_.Y
rlabel metal1 1184 3122 1256 3138 0 _803_.gnd
rlabel metal1 1184 3362 1256 3378 0 _803_.vdd
rlabel metal2 1233 3193 1247 3207 0 _803_.A
rlabel metal2 1213 3233 1227 3247 0 _803_.Y
rlabel metal1 1584 3122 1696 3138 0 _1506_.gnd
rlabel metal1 1584 3362 1696 3378 0 _1506_.vdd
rlabel metal2 1673 3213 1687 3227 0 _1506_.A
rlabel metal2 1653 3233 1667 3247 0 _1506_.B
rlabel metal2 1613 3233 1627 3247 0 _1506_.C
rlabel metal2 1633 3213 1647 3227 0 _1506_.Y
rlabel metal1 1484 3122 1596 3138 0 _805_.gnd
rlabel metal1 1484 3362 1596 3378 0 _805_.vdd
rlabel metal2 1493 3213 1507 3227 0 _805_.A
rlabel metal2 1513 3233 1527 3247 0 _805_.B
rlabel metal2 1553 3233 1567 3247 0 _805_.C
rlabel metal2 1533 3213 1547 3227 0 _805_.Y
rlabel metal1 1564 3122 1656 3138 0 _1516_.gnd
rlabel metal1 1564 2882 1656 2898 0 _1516_.vdd
rlabel metal2 1593 3033 1607 3047 0 _1516_.B
rlabel metal2 1633 3033 1647 3047 0 _1516_.A
rlabel metal2 1613 3053 1627 3067 0 _1516_.Y
rlabel metal1 1844 3122 1956 3138 0 _1508_.gnd
rlabel metal1 1844 3362 1956 3378 0 _1508_.vdd
rlabel metal2 1933 3213 1947 3227 0 _1508_.A
rlabel metal2 1913 3233 1927 3247 0 _1508_.B
rlabel metal2 1873 3233 1887 3247 0 _1508_.C
rlabel metal2 1893 3213 1907 3227 0 _1508_.Y
rlabel metal1 1684 3122 1796 3138 0 _1507_.gnd
rlabel metal1 1684 3362 1796 3378 0 _1507_.vdd
rlabel metal2 1773 3213 1787 3227 0 _1507_.A
rlabel metal2 1753 3233 1767 3247 0 _1507_.B
rlabel metal2 1713 3233 1727 3247 0 _1507_.C
rlabel metal2 1733 3213 1747 3227 0 _1507_.Y
rlabel metal1 1824 3122 1936 3138 0 _1505_.gnd
rlabel metal1 1824 2882 1936 2898 0 _1505_.vdd
rlabel metal2 1913 3033 1927 3047 0 _1505_.A
rlabel metal2 1893 3013 1907 3027 0 _1505_.B
rlabel metal2 1853 3013 1867 3027 0 _1505_.C
rlabel metal2 1873 3033 1887 3047 0 _1505_.Y
rlabel metal1 1724 3122 1836 3138 0 _1504_.gnd
rlabel metal1 1724 2882 1836 2898 0 _1504_.vdd
rlabel metal2 1733 3033 1747 3047 0 _1504_.A
rlabel metal2 1753 3013 1767 3027 0 _1504_.B
rlabel metal2 1793 3013 1807 3027 0 _1504_.C
rlabel metal2 1773 3033 1787 3047 0 _1504_.Y
rlabel metal1 1644 3122 1736 3138 0 _804_.gnd
rlabel metal1 1644 2882 1736 2898 0 _804_.vdd
rlabel metal2 1713 2993 1727 3007 0 _804_.A
rlabel metal2 1673 2993 1687 3007 0 _804_.B
rlabel metal2 1693 3013 1707 3027 0 _804_.Y
rlabel metal1 1784 3122 1856 3138 0 _1501_.gnd
rlabel metal1 1784 3362 1856 3378 0 _1501_.vdd
rlabel metal2 1833 3193 1847 3207 0 _1501_.A
rlabel metal2 1813 3233 1827 3247 0 _1501_.Y
rlabel metal1 2044 3122 2296 3138 0 _1587_.gnd
rlabel metal1 2044 3362 2296 3378 0 _1587_.vdd
rlabel metal2 2193 3213 2207 3227 0 _1587_.D
rlabel metal2 2153 3213 2167 3227 0 _1587_.CLK
rlabel metal2 2073 3213 2087 3227 0 _1587_.Q
rlabel metal1 1924 3122 2176 3138 0 _1585_.gnd
rlabel metal1 1924 2882 2176 2898 0 _1585_.vdd
rlabel metal2 2073 3033 2087 3047 0 _1585_.D
rlabel metal2 2033 3033 2047 3047 0 _1585_.CLK
rlabel metal2 1953 3033 1967 3047 0 _1585_.Q
rlabel metal1 1944 3122 2056 3138 0 _1509_.gnd
rlabel metal1 1944 3362 2056 3378 0 _1509_.vdd
rlabel metal2 2033 3213 2047 3227 0 _1509_.A
rlabel metal2 2013 3233 2027 3247 0 _1509_.B
rlabel metal2 1973 3233 1987 3247 0 _1509_.C
rlabel metal2 1993 3213 2007 3227 0 _1509_.Y
rlabel metal1 2404 3122 2516 3138 0 _877_.gnd
rlabel metal1 2404 2882 2516 2898 0 _877_.vdd
rlabel metal2 2493 3013 2507 3027 0 _877_.A
rlabel metal2 2473 3053 2487 3067 0 _877_.B
rlabel metal2 2453 3013 2467 3027 0 _877_.C
rlabel metal2 2433 3033 2447 3047 0 _877_.Y
rlabel metal1 2164 3122 2256 3138 0 _878_.gnd
rlabel metal1 2164 2882 2256 2898 0 _878_.vdd
rlabel metal2 2193 3033 2207 3047 0 _878_.B
rlabel metal2 2233 3033 2247 3047 0 _878_.A
rlabel metal2 2213 3053 2227 3067 0 _878_.Y
rlabel metal1 2284 3122 2356 3138 0 _876_.gnd
rlabel metal1 2284 3362 2356 3378 0 _876_.vdd
rlabel metal2 2333 3193 2347 3207 0 _876_.A
rlabel metal2 2313 3233 2327 3247 0 _876_.Y
rlabel metal1 2344 3122 2416 3138 0 _870_.gnd
rlabel metal1 2344 3362 2416 3378 0 _870_.vdd
rlabel metal2 2393 3193 2407 3207 0 _870_.A
rlabel metal2 2373 3233 2387 3247 0 _870_.Y
rlabel metal1 2244 3122 2316 3138 0 _858_.gnd
rlabel metal1 2244 2882 2316 2898 0 _858_.vdd
rlabel metal2 2293 3053 2307 3067 0 _858_.A
rlabel metal2 2273 3013 2287 3027 0 _858_.Y
rlabel metal1 2404 3122 2516 3138 0 _874_.gnd
rlabel metal1 2404 3362 2516 3378 0 _874_.vdd
rlabel metal2 2493 3233 2507 3247 0 _874_.A
rlabel metal2 2473 3253 2487 3267 0 _874_.B
rlabel metal2 2453 3233 2467 3247 0 _874_.C
rlabel metal2 2433 3253 2447 3267 0 _874_.Y
rlabel metal1 2304 3122 2416 3138 0 _852_.gnd
rlabel metal1 2304 2882 2416 2898 0 _852_.vdd
rlabel metal2 2393 3013 2407 3027 0 _852_.A
rlabel metal2 2373 2993 2387 3007 0 _852_.B
rlabel metal2 2353 3013 2367 3027 0 _852_.C
rlabel metal2 2333 2993 2347 3007 0 _852_.Y
rlabel metal1 2664 3122 2776 3138 0 _895_.gnd
rlabel metal1 2664 3362 2776 3378 0 _895_.vdd
rlabel metal2 2753 3213 2767 3227 0 _895_.A
rlabel metal2 2733 3233 2747 3247 0 _895_.B
rlabel metal2 2693 3233 2707 3247 0 _895_.C
rlabel metal2 2713 3213 2727 3227 0 _895_.Y
rlabel metal1 2604 3122 2716 3138 0 _869_.gnd
rlabel metal1 2604 2882 2716 2898 0 _869_.vdd
rlabel metal2 2693 3033 2707 3047 0 _869_.A
rlabel metal2 2673 3013 2687 3027 0 _869_.B
rlabel metal2 2633 3013 2647 3027 0 _869_.C
rlabel metal2 2653 3033 2667 3047 0 _869_.Y
rlabel metal1 2504 3122 2616 3138 0 _883_.gnd
rlabel metal1 2504 3362 2616 3378 0 _883_.vdd
rlabel metal2 2513 3233 2527 3247 0 _883_.A
rlabel metal2 2533 3193 2547 3207 0 _883_.B
rlabel metal2 2553 3233 2567 3247 0 _883_.C
rlabel metal2 2573 3213 2587 3227 0 _883_.Y
rlabel metal1 2604 3122 2676 3138 0 _873_.gnd
rlabel metal1 2604 3362 2676 3378 0 _873_.vdd
rlabel metal2 2653 3193 2667 3207 0 _873_.A
rlabel metal2 2633 3233 2647 3247 0 _873_.Y
rlabel metal1 2504 3122 2616 3138 0 _875_.gnd
rlabel metal1 2504 2882 2616 2898 0 _875_.vdd
rlabel metal2 2593 3013 2607 3027 0 _875_.A
rlabel metal2 2573 2993 2587 3007 0 _875_.B
rlabel metal2 2553 3013 2567 3027 0 _875_.C
rlabel metal2 2533 2993 2547 3007 0 _875_.Y
rlabel metal1 2844 3122 2956 3138 0 _788_.gnd
rlabel metal1 2844 3362 2956 3378 0 _788_.vdd
rlabel metal2 2853 3213 2867 3227 0 _788_.A
rlabel metal2 2873 3233 2887 3247 0 _788_.B
rlabel metal2 2913 3233 2927 3247 0 _788_.C
rlabel metal2 2893 3213 2907 3227 0 _788_.Y
rlabel metal1 2784 3122 2876 3138 0 _856_.gnd
rlabel metal1 2784 2882 2876 2898 0 _856_.vdd
rlabel metal2 2793 2993 2807 3007 0 _856_.A
rlabel metal2 2833 2993 2847 3007 0 _856_.B
rlabel metal2 2813 3013 2827 3027 0 _856_.Y
rlabel metal1 2864 3122 2956 3138 0 _855_.gnd
rlabel metal1 2864 2882 2956 2898 0 _855_.vdd
rlabel metal2 2873 2993 2887 3007 0 _855_.A
rlabel metal2 2913 2993 2927 3007 0 _855_.B
rlabel metal2 2893 3013 2907 3027 0 _855_.Y
rlabel metal1 2764 3122 2856 3138 0 _867_.gnd
rlabel metal1 2764 3362 2856 3378 0 _867_.vdd
rlabel metal2 2813 3213 2827 3227 0 _867_.B
rlabel metal2 2773 3213 2787 3227 0 _867_.A
rlabel metal2 2793 3193 2807 3207 0 _867_.Y
rlabel metal1 2704 3122 2796 3138 0 _857_.gnd
rlabel metal1 2704 2882 2796 2898 0 _857_.vdd
rlabel metal2 2733 3033 2747 3047 0 _857_.B
rlabel metal2 2773 3033 2787 3047 0 _857_.A
rlabel metal2 2753 3053 2767 3067 0 _857_.Y
rlabel metal1 3144 3122 3256 3138 0 _898_.gnd
rlabel metal1 3144 2882 3256 2898 0 _898_.vdd
rlabel metal2 3153 3033 3167 3047 0 _898_.A
rlabel metal2 3173 3013 3187 3027 0 _898_.B
rlabel metal2 3213 3013 3227 3027 0 _898_.C
rlabel metal2 3193 3033 3207 3047 0 _898_.Y
rlabel metal1 3024 3122 3116 3138 0 _884_.gnd
rlabel metal1 3024 3362 3116 3378 0 _884_.vdd
rlabel metal2 3033 3253 3047 3267 0 _884_.A
rlabel metal2 3073 3253 3087 3267 0 _884_.B
rlabel metal2 3053 3233 3067 3247 0 _884_.Y
rlabel metal1 3064 3122 3156 3138 0 _865_.gnd
rlabel metal1 3064 2882 3156 2898 0 _865_.vdd
rlabel metal2 3073 2993 3087 3007 0 _865_.A
rlabel metal2 3113 2993 3127 3007 0 _865_.B
rlabel metal2 3093 3013 3107 3027 0 _865_.Y
rlabel metal1 2944 3122 3036 3138 0 _787_.gnd
rlabel metal1 2944 3362 3036 3378 0 _787_.vdd
rlabel metal2 2953 3253 2967 3267 0 _787_.A
rlabel metal2 2993 3253 3007 3267 0 _787_.B
rlabel metal2 2973 3233 2987 3247 0 _787_.Y
rlabel metal1 3104 3122 3216 3138 0 _902_.gnd
rlabel metal1 3104 3362 3216 3378 0 _902_.vdd
rlabel metal2 3193 3233 3207 3247 0 _902_.A
rlabel metal2 3173 3193 3187 3207 0 _902_.B
rlabel metal2 3153 3233 3167 3247 0 _902_.C
rlabel metal2 3133 3213 3147 3227 0 _902_.Y
rlabel metal1 3204 3122 3316 3138 0 _872_.gnd
rlabel metal1 3204 3362 3316 3378 0 _872_.vdd
rlabel metal2 3293 3233 3307 3247 0 _872_.A
rlabel metal2 3273 3253 3287 3267 0 _872_.B
rlabel metal2 3253 3233 3267 3247 0 _872_.C
rlabel metal2 3233 3253 3247 3267 0 _872_.Y
rlabel metal1 2944 3122 3076 3138 0 _868_.gnd
rlabel metal1 2944 2882 3076 2898 0 _868_.vdd
rlabel metal2 2953 3033 2967 3047 0 _868_.A
rlabel metal2 2973 3013 2987 3027 0 _868_.B
rlabel metal2 3033 3033 3047 3047 0 _868_.C
rlabel metal2 3013 3013 3027 3027 0 _868_.D
rlabel metal2 2993 3033 3007 3047 0 _868_.Y
rlabel metal1 3404 3122 3496 3138 0 BUFX2_insert31.gnd
rlabel metal1 3404 2882 3496 2898 0 BUFX2_insert31.vdd
rlabel metal2 3473 3033 3487 3047 0 BUFX2_insert31.A
rlabel metal2 3433 3033 3447 3047 0 BUFX2_insert31.Y
rlabel metal1 3304 3122 3416 3138 0 _901_.gnd
rlabel metal1 3304 3362 3416 3378 0 _901_.vdd
rlabel metal2 3393 3213 3407 3227 0 _901_.A
rlabel metal2 3373 3233 3387 3247 0 _901_.B
rlabel metal2 3333 3233 3347 3247 0 _901_.C
rlabel metal2 3353 3213 3367 3227 0 _901_.Y
rlabel metal1 3304 3122 3416 3138 0 _954_.gnd
rlabel metal1 3304 2882 3416 2898 0 _954_.vdd
rlabel metal2 3313 3033 3327 3047 0 _954_.A
rlabel metal2 3373 3033 3387 3047 0 _954_.Y
rlabel metal2 3353 2993 3367 3007 0 _954_.B
rlabel metal1 3404 3122 3516 3138 0 _871_.gnd
rlabel metal1 3404 3362 3516 3378 0 _871_.vdd
rlabel metal2 3493 3213 3507 3227 0 _871_.A
rlabel metal2 3433 3213 3447 3227 0 _871_.Y
rlabel metal2 3453 3253 3467 3267 0 _871_.B
rlabel metal1 3244 3122 3316 3138 0 _897_.gnd
rlabel metal1 3244 2882 3316 2898 0 _897_.vdd
rlabel metal2 3253 3013 3267 3027 0 _897_.A
rlabel metal2 3273 3033 3287 3047 0 _897_.Y
rlabel metal1 3484 3122 3576 3138 0 BUFX2_insert21.gnd
rlabel metal1 3484 2882 3576 2898 0 BUFX2_insert21.vdd
rlabel metal2 3553 3033 3567 3047 0 BUFX2_insert21.A
rlabel metal2 3513 3033 3527 3047 0 BUFX2_insert21.Y
rlabel metal1 3644 3122 3756 3138 0 _1010_.gnd
rlabel metal1 3644 2882 3756 2898 0 _1010_.vdd
rlabel metal2 3653 3033 3667 3047 0 _1010_.A
rlabel metal2 3673 3013 3687 3027 0 _1010_.B
rlabel metal2 3713 3013 3727 3027 0 _1010_.C
rlabel metal2 3693 3033 3707 3047 0 _1010_.Y
rlabel metal1 3564 3122 3656 3138 0 _1009_.gnd
rlabel metal1 3564 2882 3656 2898 0 _1009_.vdd
rlabel metal2 3573 2993 3587 3007 0 _1009_.A
rlabel metal2 3613 2993 3627 3007 0 _1009_.B
rlabel metal2 3593 3013 3607 3027 0 _1009_.Y
rlabel metal1 3504 3122 3596 3138 0 _885_.gnd
rlabel metal1 3504 3362 3596 3378 0 _885_.vdd
rlabel metal2 3513 3253 3527 3267 0 _885_.A
rlabel metal2 3553 3253 3567 3267 0 _885_.B
rlabel metal2 3533 3233 3547 3247 0 _885_.Y
rlabel metal1 3684 3122 3816 3138 0 _920_.gnd
rlabel metal1 3684 3362 3816 3378 0 _920_.vdd
rlabel metal2 3793 3213 3807 3227 0 _920_.A
rlabel metal2 3773 3233 3787 3247 0 _920_.B
rlabel metal2 3713 3213 3727 3227 0 _920_.C
rlabel metal2 3733 3233 3747 3247 0 _920_.D
rlabel metal2 3753 3213 3767 3227 0 _920_.Y
rlabel metal1 3584 3122 3696 3138 0 _890_.gnd
rlabel metal1 3584 3362 3696 3378 0 _890_.vdd
rlabel metal2 3673 3213 3687 3227 0 _890_.A
rlabel metal2 3613 3213 3627 3227 0 _890_.Y
rlabel metal2 3633 3253 3647 3267 0 _890_.B
rlabel metal1 3744 3122 3836 3138 0 BUFX2_insert22.gnd
rlabel metal1 3744 2882 3836 2898 0 BUFX2_insert22.vdd
rlabel metal2 3813 3033 3827 3047 0 BUFX2_insert22.A
rlabel metal2 3773 3033 3787 3047 0 BUFX2_insert22.Y
rlabel metal1 3824 3122 3936 3138 0 _1022_.gnd
rlabel metal1 3824 2882 3936 2898 0 _1022_.vdd
rlabel metal2 3833 3033 3847 3047 0 _1022_.A
rlabel metal2 3853 3013 3867 3027 0 _1022_.B
rlabel metal2 3893 3013 3907 3027 0 _1022_.C
rlabel metal2 3873 3033 3887 3047 0 _1022_.Y
rlabel metal1 3884 3122 3996 3138 0 _979_.gnd
rlabel metal1 3884 3362 3996 3378 0 _979_.vdd
rlabel metal2 3893 3213 3907 3227 0 _979_.A
rlabel metal2 3913 3233 3927 3247 0 _979_.B
rlabel metal2 3953 3233 3967 3247 0 _979_.C
rlabel metal2 3933 3213 3947 3227 0 _979_.Y
rlabel metal1 3804 3122 3896 3138 0 _974_.gnd
rlabel metal1 3804 3362 3896 3378 0 _974_.vdd
rlabel metal2 3873 3253 3887 3267 0 _974_.A
rlabel metal2 3833 3253 3847 3267 0 _974_.B
rlabel metal2 3853 3233 3867 3247 0 _974_.Y
rlabel metal1 3984 3122 4076 3138 0 _925_.gnd
rlabel metal1 3984 3362 4076 3378 0 _925_.vdd
rlabel metal2 3993 3253 4007 3267 0 _925_.A
rlabel metal2 4033 3253 4047 3267 0 _925_.B
rlabel metal2 4013 3233 4027 3247 0 _925_.Y
rlabel metal1 3924 3122 4036 3138 0 _1023_.gnd
rlabel metal1 3924 2882 4036 2898 0 _1023_.vdd
rlabel metal2 3933 3013 3947 3027 0 _1023_.A
rlabel metal2 3953 2993 3967 3007 0 _1023_.B
rlabel metal2 3973 3013 3987 3027 0 _1023_.C
rlabel metal2 3993 2993 4007 3007 0 _1023_.Y
rlabel metal1 4024 3122 4116 3138 0 BUFX2_insert32.gnd
rlabel metal1 4024 2882 4116 2898 0 BUFX2_insert32.vdd
rlabel metal2 4033 3033 4047 3047 0 BUFX2_insert32.A
rlabel metal2 4073 3033 4087 3047 0 BUFX2_insert32.Y
rlabel metal1 4164 3122 4256 3138 0 _1074_.gnd
rlabel metal1 4164 3362 4256 3378 0 _1074_.vdd
rlabel metal2 4173 3253 4187 3267 0 _1074_.A
rlabel metal2 4213 3253 4227 3267 0 _1074_.B
rlabel metal2 4193 3233 4207 3247 0 _1074_.Y
rlabel metal1 4104 3122 4216 3138 0 _1042_.gnd
rlabel metal1 4104 2882 4216 2898 0 _1042_.vdd
rlabel metal2 4193 3013 4207 3027 0 _1042_.A
rlabel metal2 4173 3053 4187 3067 0 _1042_.B
rlabel metal2 4153 3013 4167 3027 0 _1042_.C
rlabel metal2 4133 3033 4147 3047 0 _1042_.Y
rlabel metal1 4204 3122 4316 3138 0 _1032_.gnd
rlabel metal1 4204 2882 4316 2898 0 _1032_.vdd
rlabel metal2 4213 3013 4227 3027 0 _1032_.A
rlabel metal2 4233 2993 4247 3007 0 _1032_.B
rlabel metal2 4253 3013 4267 3027 0 _1032_.C
rlabel metal2 4273 2993 4287 3007 0 _1032_.Y
rlabel metal1 4244 3122 4356 3138 0 _1045_.gnd
rlabel metal1 4244 3362 4356 3378 0 _1045_.vdd
rlabel metal2 4253 3213 4267 3227 0 _1045_.A
rlabel metal2 4313 3213 4327 3227 0 _1045_.Y
rlabel metal2 4293 3253 4307 3267 0 _1045_.B
rlabel metal1 4064 3122 4176 3138 0 _918_.gnd
rlabel metal1 4064 3362 4176 3378 0 _918_.vdd
rlabel metal2 4153 3213 4167 3227 0 _918_.A
rlabel metal2 4093 3213 4107 3227 0 _918_.Y
rlabel metal2 4113 3253 4127 3267 0 _918_.B
rlabel metal1 4444 3122 4556 3138 0 _1076_.gnd
rlabel metal1 4444 3362 4556 3378 0 _1076_.vdd
rlabel metal2 4453 3213 4467 3227 0 _1076_.A
rlabel metal2 4473 3233 4487 3247 0 _1076_.B
rlabel metal2 4513 3233 4527 3247 0 _1076_.C
rlabel metal2 4493 3213 4507 3227 0 _1076_.Y
rlabel metal1 4344 3122 4456 3138 0 _1075_.gnd
rlabel metal1 4344 3362 4456 3378 0 _1075_.vdd
rlabel metal2 4353 3233 4367 3247 0 _1075_.A
rlabel metal2 4373 3193 4387 3207 0 _1075_.B
rlabel metal2 4393 3233 4407 3247 0 _1075_.C
rlabel metal2 4413 3213 4427 3227 0 _1075_.Y
rlabel metal1 4304 3122 4416 3138 0 _1041_.gnd
rlabel metal1 4304 2882 4416 2898 0 _1041_.vdd
rlabel metal2 4393 3013 4407 3027 0 _1041_.A
rlabel metal2 4373 3053 4387 3067 0 _1041_.B
rlabel metal2 4353 3013 4367 3027 0 _1041_.C
rlabel metal2 4333 3033 4347 3047 0 _1041_.Y
rlabel metal1 4504 3122 4576 3138 0 _1489_.gnd
rlabel metal1 4504 2882 4576 2898 0 _1489_.vdd
rlabel metal2 4553 3053 4567 3067 0 _1489_.A
rlabel metal2 4533 3013 4547 3027 0 _1489_.Y
rlabel metal1 4404 3122 4516 3138 0 _1037_.gnd
rlabel metal1 4404 2882 4516 2898 0 _1037_.vdd
rlabel metal2 4493 3013 4507 3027 0 _1037_.A
rlabel metal2 4473 2993 4487 3007 0 _1037_.B
rlabel metal2 4453 3013 4467 3027 0 _1037_.C
rlabel metal2 4433 2993 4447 3007 0 _1037_.Y
rlabel nsubstratencontact 4756 3368 4756 3368 0 FILL71250x46950.vdd
rlabel metal1 4744 3122 4776 3138 0 FILL71250x46950.gnd
rlabel metal1 4544 3122 4656 3138 0 _1141_.gnd
rlabel metal1 4544 3362 4656 3378 0 _1141_.vdd
rlabel metal2 4553 3213 4567 3227 0 _1141_.A
rlabel metal2 4573 3233 4587 3247 0 _1141_.B
rlabel metal2 4613 3233 4627 3247 0 _1141_.C
rlabel metal2 4593 3213 4607 3227 0 _1141_.Y
rlabel metal1 4564 3122 4676 3138 0 _1120_.gnd
rlabel metal1 4564 2882 4676 2898 0 _1120_.vdd
rlabel metal2 4653 3033 4667 3047 0 _1120_.A
rlabel metal2 4633 3013 4647 3027 0 _1120_.B
rlabel metal2 4593 3013 4607 3027 0 _1120_.C
rlabel metal2 4613 3033 4627 3047 0 _1120_.Y
rlabel metal1 4664 3122 4776 3138 0 _1116_.gnd
rlabel metal1 4664 2882 4776 2898 0 _1116_.vdd
rlabel metal2 4673 3033 4687 3047 0 _1116_.A
rlabel metal2 4693 3013 4707 3027 0 _1116_.B
rlabel metal2 4733 3013 4747 3027 0 _1116_.C
rlabel metal2 4713 3033 4727 3047 0 _1116_.Y
rlabel metal1 4644 3122 4756 3138 0 _1119_.gnd
rlabel metal1 4644 3362 4756 3378 0 _1119_.vdd
rlabel metal2 4733 3233 4747 3247 0 _1119_.A
rlabel metal2 4713 3253 4727 3267 0 _1119_.B
rlabel metal2 4693 3233 4707 3247 0 _1119_.C
rlabel metal2 4673 3253 4687 3267 0 _1119_.Y
rlabel metal1 4 3602 256 3618 0 _1563_.gnd
rlabel metal1 4 3362 256 3378 0 _1563_.vdd
rlabel metal2 93 3513 107 3527 0 _1563_.D
rlabel metal2 133 3513 147 3527 0 _1563_.CLK
rlabel metal2 213 3513 227 3527 0 _1563_.Q
rlabel metal1 244 3602 336 3618 0 _1350_.gnd
rlabel metal1 244 3362 336 3378 0 _1350_.vdd
rlabel metal2 313 3473 327 3487 0 _1350_.A
rlabel metal2 273 3473 287 3487 0 _1350_.B
rlabel metal2 293 3493 307 3507 0 _1350_.Y
rlabel metal1 324 3602 436 3618 0 _1351_.gnd
rlabel metal1 324 3362 436 3378 0 _1351_.vdd
rlabel metal2 413 3513 427 3527 0 _1351_.A
rlabel metal2 393 3493 407 3507 0 _1351_.B
rlabel metal2 353 3493 367 3507 0 _1351_.C
rlabel metal2 373 3513 387 3527 0 _1351_.Y
rlabel metal1 424 3602 516 3618 0 _1349_.gnd
rlabel metal1 424 3362 516 3378 0 _1349_.vdd
rlabel metal2 493 3473 507 3487 0 _1349_.A
rlabel metal2 453 3473 467 3487 0 _1349_.B
rlabel metal2 473 3493 487 3507 0 _1349_.Y
rlabel metal1 504 3602 616 3618 0 _1348_.gnd
rlabel metal1 504 3362 616 3378 0 _1348_.vdd
rlabel metal2 593 3493 607 3507 0 _1348_.A
rlabel metal2 573 3473 587 3487 0 _1348_.B
rlabel metal2 553 3493 567 3507 0 _1348_.C
rlabel metal2 533 3473 547 3487 0 _1348_.Y
rlabel metal1 664 3602 776 3618 0 _1355_.gnd
rlabel metal1 664 3362 776 3378 0 _1355_.vdd
rlabel metal2 753 3513 767 3527 0 _1355_.A
rlabel metal2 733 3493 747 3507 0 _1355_.B
rlabel metal2 693 3493 707 3507 0 _1355_.C
rlabel metal2 713 3513 727 3527 0 _1355_.Y
rlabel metal1 764 3602 876 3618 0 _1344_.gnd
rlabel metal1 764 3362 876 3378 0 _1344_.vdd
rlabel metal2 853 3513 867 3527 0 _1344_.A
rlabel metal2 833 3493 847 3507 0 _1344_.B
rlabel metal2 793 3493 807 3507 0 _1344_.C
rlabel metal2 813 3513 827 3527 0 _1344_.Y
rlabel metal1 604 3602 676 3618 0 _1346_.gnd
rlabel metal1 604 3362 676 3378 0 _1346_.vdd
rlabel metal2 653 3533 667 3547 0 _1346_.A
rlabel metal2 633 3493 647 3507 0 _1346_.Y
rlabel metal1 1004 3602 1256 3618 0 _1533_.gnd
rlabel metal1 1004 3362 1256 3378 0 _1533_.vdd
rlabel metal2 1153 3513 1167 3527 0 _1533_.D
rlabel metal2 1113 3513 1127 3527 0 _1533_.CLK
rlabel metal2 1033 3513 1047 3527 0 _1533_.Q
rlabel metal1 924 3602 1016 3618 0 _1342_.gnd
rlabel metal1 924 3362 1016 3378 0 _1342_.vdd
rlabel metal2 953 3513 967 3527 0 _1342_.B
rlabel metal2 993 3513 1007 3527 0 _1342_.A
rlabel metal2 973 3533 987 3547 0 _1342_.Y
rlabel metal1 864 3602 936 3618 0 _1347_.gnd
rlabel metal1 864 3362 936 3378 0 _1347_.vdd
rlabel metal2 873 3533 887 3547 0 _1347_.A
rlabel metal2 893 3493 907 3507 0 _1347_.Y
rlabel metal1 1304 3602 1396 3618 0 _1343_.gnd
rlabel metal1 1304 3362 1396 3378 0 _1343_.vdd
rlabel metal2 1353 3513 1367 3527 0 _1343_.B
rlabel metal2 1313 3513 1327 3527 0 _1343_.A
rlabel metal2 1333 3533 1347 3547 0 _1343_.Y
rlabel metal1 1244 3602 1316 3618 0 _812_.gnd
rlabel metal1 1244 3362 1316 3378 0 _812_.vdd
rlabel metal2 1253 3533 1267 3547 0 _812_.A
rlabel metal2 1273 3493 1287 3507 0 _812_.Y
rlabel metal1 1564 3602 1656 3618 0 BUFX2_insert3.gnd
rlabel metal1 1564 3362 1656 3378 0 BUFX2_insert3.vdd
rlabel metal2 1633 3513 1647 3527 0 BUFX2_insert3.A
rlabel metal2 1593 3513 1607 3527 0 BUFX2_insert3.Y
rlabel metal1 1384 3602 1496 3618 0 _814_.gnd
rlabel metal1 1384 3362 1496 3378 0 _814_.vdd
rlabel metal2 1393 3513 1407 3527 0 _814_.A
rlabel metal2 1413 3493 1427 3507 0 _814_.B
rlabel metal2 1453 3493 1467 3507 0 _814_.C
rlabel metal2 1433 3513 1447 3527 0 _814_.Y
rlabel metal1 1484 3602 1576 3618 0 _813_.gnd
rlabel metal1 1484 3362 1576 3378 0 _813_.vdd
rlabel metal2 1493 3473 1507 3487 0 _813_.A
rlabel metal2 1533 3473 1547 3487 0 _813_.B
rlabel metal2 1513 3493 1527 3507 0 _813_.Y
rlabel metal1 1704 3602 1956 3618 0 _1586_.gnd
rlabel metal1 1704 3362 1956 3378 0 _1586_.vdd
rlabel metal2 1853 3513 1867 3527 0 _1586_.D
rlabel metal2 1813 3513 1827 3527 0 _1586_.CLK
rlabel metal2 1733 3513 1747 3527 0 _1586_.Q
rlabel metal1 1644 3602 1716 3618 0 _881_.gnd
rlabel metal1 1644 3362 1716 3378 0 _881_.vdd
rlabel metal2 1693 3533 1707 3547 0 _881_.A
rlabel metal2 1673 3493 1687 3507 0 _881_.Y
rlabel metal1 2064 3602 2156 3618 0 _911_.gnd
rlabel metal1 2064 3362 2156 3378 0 _911_.vdd
rlabel metal2 2073 3473 2087 3487 0 _911_.A
rlabel metal2 2113 3473 2127 3487 0 _911_.B
rlabel metal2 2093 3493 2107 3507 0 _911_.Y
rlabel metal1 1944 3602 2076 3618 0 _912_.gnd
rlabel metal1 1944 3362 2076 3378 0 _912_.vdd
rlabel metal2 1953 3513 1967 3527 0 _912_.A
rlabel metal2 1973 3493 1987 3507 0 _912_.B
rlabel metal2 2033 3513 2047 3527 0 _912_.C
rlabel metal2 1993 3513 2007 3527 0 _912_.Y
rlabel metal2 2013 3493 2027 3507 0 _912_.D
rlabel metal1 2144 3602 2256 3618 0 _909_.gnd
rlabel metal1 2144 3362 2256 3378 0 _909_.vdd
rlabel metal2 2233 3493 2247 3507 0 _909_.A
rlabel metal2 2213 3533 2227 3547 0 _909_.B
rlabel metal2 2193 3493 2207 3507 0 _909_.C
rlabel metal2 2173 3513 2187 3527 0 _909_.Y
rlabel metal1 2344 3602 2416 3618 0 _905_.gnd
rlabel metal1 2344 3362 2416 3378 0 _905_.vdd
rlabel metal2 2393 3533 2407 3547 0 _905_.A
rlabel metal2 2373 3493 2387 3507 0 _905_.Y
rlabel metal1 2244 3602 2356 3618 0 _910_.gnd
rlabel metal1 2244 3362 2356 3378 0 _910_.vdd
rlabel metal2 2333 3493 2347 3507 0 _910_.A
rlabel metal2 2313 3473 2327 3487 0 _910_.B
rlabel metal2 2293 3493 2307 3507 0 _910_.C
rlabel metal2 2273 3473 2287 3487 0 _910_.Y
rlabel metal1 2404 3602 2516 3618 0 _904_.gnd
rlabel metal1 2404 3362 2516 3378 0 _904_.vdd
rlabel metal2 2493 3493 2507 3507 0 _904_.A
rlabel metal2 2473 3473 2487 3487 0 _904_.B
rlabel metal2 2453 3493 2467 3507 0 _904_.C
rlabel metal2 2433 3473 2447 3487 0 _904_.Y
rlabel metal1 2604 3602 2716 3618 0 _907_.gnd
rlabel metal1 2604 3362 2716 3378 0 _907_.vdd
rlabel metal2 2693 3513 2707 3527 0 _907_.A
rlabel metal2 2673 3493 2687 3507 0 _907_.B
rlabel metal2 2633 3493 2647 3507 0 _907_.C
rlabel metal2 2653 3513 2667 3527 0 _907_.Y
rlabel metal1 2504 3602 2616 3618 0 _894_.gnd
rlabel metal1 2504 3362 2616 3378 0 _894_.vdd
rlabel metal2 2593 3493 2607 3507 0 _894_.A
rlabel metal2 2573 3473 2587 3487 0 _894_.B
rlabel metal2 2553 3493 2567 3507 0 _894_.C
rlabel metal2 2533 3473 2547 3487 0 _894_.Y
rlabel metal1 2704 3602 2816 3618 0 _903_.gnd
rlabel metal1 2704 3362 2816 3378 0 _903_.vdd
rlabel metal2 2713 3513 2727 3527 0 _903_.A
rlabel metal2 2733 3493 2747 3507 0 _903_.B
rlabel metal2 2773 3493 2787 3507 0 _903_.C
rlabel metal2 2753 3513 2767 3527 0 _903_.Y
rlabel metal1 2884 3602 2996 3618 0 _888_.gnd
rlabel metal1 2884 3362 2996 3378 0 _888_.vdd
rlabel metal2 2893 3513 2907 3527 0 _888_.A
rlabel metal2 2913 3493 2927 3507 0 _888_.B
rlabel metal2 2953 3493 2967 3507 0 _888_.C
rlabel metal2 2933 3513 2947 3527 0 _888_.Y
rlabel metal1 2804 3602 2896 3618 0 _866_.gnd
rlabel metal1 2804 3362 2896 3378 0 _866_.vdd
rlabel metal2 2813 3473 2827 3487 0 _866_.A
rlabel metal2 2853 3473 2867 3487 0 _866_.B
rlabel metal2 2833 3493 2847 3507 0 _866_.Y
rlabel metal1 3064 3602 3176 3618 0 _917_.gnd
rlabel metal1 3064 3362 3176 3378 0 _917_.vdd
rlabel metal2 3153 3513 3167 3527 0 _917_.A
rlabel metal2 3133 3493 3147 3507 0 _917_.B
rlabel metal2 3093 3493 3107 3507 0 _917_.C
rlabel metal2 3113 3513 3127 3527 0 _917_.Y
rlabel metal1 2984 3602 3076 3618 0 _886_.gnd
rlabel metal1 2984 3362 3076 3378 0 _886_.vdd
rlabel metal2 3033 3513 3047 3527 0 _886_.B
rlabel metal2 2993 3513 3007 3527 0 _886_.A
rlabel metal2 3013 3533 3027 3547 0 _886_.Y
rlabel metal1 3164 3602 3296 3618 0 _887_.gnd
rlabel metal1 3164 3362 3296 3378 0 _887_.vdd
rlabel metal2 3173 3513 3187 3527 0 _887_.A
rlabel metal2 3193 3493 3207 3507 0 _887_.B
rlabel metal2 3253 3513 3267 3527 0 _887_.C
rlabel metal2 3233 3493 3247 3507 0 _887_.D
rlabel metal2 3213 3513 3227 3527 0 _887_.Y
rlabel metal1 3364 3602 3456 3618 0 _955_.gnd
rlabel metal1 3364 3362 3456 3378 0 _955_.vdd
rlabel metal2 3373 3473 3387 3487 0 _955_.A
rlabel metal2 3413 3473 3427 3487 0 _955_.B
rlabel metal2 3393 3493 3407 3507 0 _955_.Y
rlabel metal1 3444 3602 3536 3618 0 _922_.gnd
rlabel metal1 3444 3362 3536 3378 0 _922_.vdd
rlabel metal2 3453 3473 3467 3487 0 _922_.A
rlabel metal2 3493 3473 3507 3487 0 _922_.B
rlabel metal2 3473 3493 3487 3507 0 _922_.Y
rlabel metal1 3284 3602 3376 3618 0 _891_.gnd
rlabel metal1 3284 3362 3376 3378 0 _891_.vdd
rlabel metal2 3293 3473 3307 3487 0 _891_.A
rlabel metal2 3333 3473 3347 3487 0 _891_.B
rlabel metal2 3313 3493 3327 3507 0 _891_.Y
rlabel metal1 3684 3602 3776 3618 0 _971_.gnd
rlabel metal1 3684 3362 3776 3378 0 _971_.vdd
rlabel metal2 3693 3473 3707 3487 0 _971_.A
rlabel metal2 3733 3473 3747 3487 0 _971_.B
rlabel metal2 3713 3493 3727 3507 0 _971_.Y
rlabel metal1 3604 3602 3696 3618 0 _919_.gnd
rlabel metal1 3604 3362 3696 3378 0 _919_.vdd
rlabel metal2 3613 3473 3627 3487 0 _919_.A
rlabel metal2 3653 3473 3667 3487 0 _919_.B
rlabel metal2 3633 3493 3647 3507 0 _919_.Y
rlabel metal1 3524 3602 3616 3618 0 _926_.gnd
rlabel metal1 3524 3362 3616 3378 0 _926_.vdd
rlabel metal2 3573 3513 3587 3527 0 _926_.B
rlabel metal2 3533 3513 3547 3527 0 _926_.A
rlabel metal2 3553 3533 3567 3547 0 _926_.Y
rlabel metal1 4004 3602 4096 3618 0 _978_.gnd
rlabel metal1 4004 3362 4096 3378 0 _978_.vdd
rlabel metal2 4013 3473 4027 3487 0 _978_.A
rlabel metal2 4053 3473 4067 3487 0 _978_.B
rlabel metal2 4033 3493 4047 3507 0 _978_.Y
rlabel metal1 3764 3602 3856 3618 0 _975_.gnd
rlabel metal1 3764 3362 3856 3378 0 _975_.vdd
rlabel metal2 3833 3473 3847 3487 0 _975_.A
rlabel metal2 3793 3473 3807 3487 0 _975_.B
rlabel metal2 3813 3493 3827 3507 0 _975_.Y
rlabel metal1 3924 3602 4016 3618 0 _973_.gnd
rlabel metal1 3924 3362 4016 3378 0 _973_.vdd
rlabel metal2 3933 3473 3947 3487 0 _973_.A
rlabel metal2 3973 3473 3987 3487 0 _973_.B
rlabel metal2 3953 3493 3967 3507 0 _973_.Y
rlabel metal1 3844 3602 3936 3618 0 _1025_.gnd
rlabel metal1 3844 3362 3936 3378 0 _1025_.vdd
rlabel metal2 3873 3513 3887 3527 0 _1025_.B
rlabel metal2 3913 3513 3927 3527 0 _1025_.A
rlabel metal2 3893 3533 3907 3547 0 _1025_.Y
rlabel metal1 4084 3602 4196 3618 0 _1040_.gnd
rlabel metal1 4084 3362 4196 3378 0 _1040_.vdd
rlabel metal2 4093 3513 4107 3527 0 _1040_.A
rlabel metal2 4113 3493 4127 3507 0 _1040_.B
rlabel metal2 4153 3493 4167 3507 0 _1040_.C
rlabel metal2 4133 3513 4147 3527 0 _1040_.Y
rlabel metal1 4184 3602 4296 3618 0 _1038_.gnd
rlabel metal1 4184 3362 4296 3378 0 _1038_.vdd
rlabel metal2 4273 3493 4287 3507 0 _1038_.A
rlabel metal2 4253 3473 4267 3487 0 _1038_.B
rlabel metal2 4233 3493 4247 3507 0 _1038_.C
rlabel metal2 4213 3473 4227 3487 0 _1038_.Y
rlabel metal1 4384 3602 4496 3618 0 _1113_.gnd
rlabel metal1 4384 3362 4496 3378 0 _1113_.vdd
rlabel metal2 4393 3493 4407 3507 0 _1113_.A
rlabel metal2 4413 3533 4427 3547 0 _1113_.B
rlabel metal2 4433 3493 4447 3507 0 _1113_.C
rlabel metal2 4453 3513 4467 3527 0 _1113_.Y
rlabel metal1 4484 3602 4556 3618 0 _1112_.gnd
rlabel metal1 4484 3362 4556 3378 0 _1112_.vdd
rlabel metal2 4493 3533 4507 3547 0 _1112_.A
rlabel metal2 4513 3493 4527 3507 0 _1112_.Y
rlabel metal1 4284 3602 4396 3618 0 _1046_.gnd
rlabel metal1 4284 3362 4396 3378 0 _1046_.vdd
rlabel metal2 4293 3493 4307 3507 0 _1046_.A
rlabel metal2 4313 3473 4327 3487 0 _1046_.B
rlabel metal2 4333 3493 4347 3507 0 _1046_.C
rlabel metal2 4353 3473 4367 3487 0 _1046_.Y
rlabel nsubstratencontact 4764 3372 4764 3372 0 FILL71250x50550.vdd
rlabel metal1 4744 3602 4776 3618 0 FILL71250x50550.gnd
rlabel metal1 4544 3602 4656 3618 0 _1123_.gnd
rlabel metal1 4544 3362 4656 3378 0 _1123_.vdd
rlabel metal2 4633 3493 4647 3507 0 _1123_.A
rlabel metal2 4613 3473 4627 3487 0 _1123_.B
rlabel metal2 4593 3493 4607 3507 0 _1123_.C
rlabel metal2 4573 3473 4587 3487 0 _1123_.Y
rlabel metal1 4644 3602 4756 3618 0 _1121_.gnd
rlabel metal1 4644 3362 4756 3378 0 _1121_.vdd
rlabel metal2 4653 3493 4667 3507 0 _1121_.A
rlabel metal2 4673 3473 4687 3487 0 _1121_.B
rlabel metal2 4693 3493 4707 3507 0 _1121_.C
rlabel metal2 4713 3473 4727 3487 0 _1121_.Y
rlabel metal1 164 3602 416 3618 0 _1565_.gnd
rlabel metal1 164 3842 416 3858 0 _1565_.vdd
rlabel metal2 313 3693 327 3707 0 _1565_.D
rlabel metal2 273 3693 287 3707 0 _1565_.CLK
rlabel metal2 193 3693 207 3707 0 _1565_.Q
rlabel metal1 4 3602 116 3618 0 _1370_.gnd
rlabel metal1 4 3842 116 3858 0 _1370_.vdd
rlabel metal2 93 3693 107 3707 0 _1370_.A
rlabel metal2 73 3713 87 3727 0 _1370_.B
rlabel metal2 33 3713 47 3727 0 _1370_.C
rlabel metal2 53 3693 67 3707 0 _1370_.Y
rlabel metal1 104 3602 176 3618 0 _1362_.gnd
rlabel metal1 104 3842 176 3858 0 _1362_.vdd
rlabel metal2 153 3673 167 3687 0 _1362_.A
rlabel metal2 133 3713 147 3727 0 _1362_.Y
rlabel metal1 404 3602 516 3618 0 _1381_.gnd
rlabel metal1 404 3842 516 3858 0 _1381_.vdd
rlabel metal2 493 3693 507 3707 0 _1381_.A
rlabel metal2 473 3713 487 3727 0 _1381_.B
rlabel metal2 433 3713 447 3727 0 _1381_.C
rlabel metal2 453 3693 467 3707 0 _1381_.Y
rlabel metal1 504 3602 616 3618 0 _1380_.gnd
rlabel metal1 504 3842 616 3858 0 _1380_.vdd
rlabel metal2 513 3693 527 3707 0 _1380_.A
rlabel metal2 573 3693 587 3707 0 _1380_.Y
rlabel metal2 553 3733 567 3747 0 _1380_.B
rlabel metal1 784 3602 1036 3618 0 _1537_.gnd
rlabel metal1 784 3842 1036 3858 0 _1537_.vdd
rlabel metal2 873 3693 887 3707 0 _1537_.D
rlabel metal2 913 3693 927 3707 0 _1537_.CLK
rlabel metal2 993 3693 1007 3707 0 _1537_.Q
rlabel metal1 704 3602 796 3618 0 _1389_.gnd
rlabel metal1 704 3842 796 3858 0 _1389_.vdd
rlabel metal2 773 3733 787 3747 0 _1389_.A
rlabel metal2 733 3733 747 3747 0 _1389_.B
rlabel metal2 753 3713 767 3727 0 _1389_.Y
rlabel metal1 604 3602 716 3618 0 _1388_.gnd
rlabel metal1 604 3842 716 3858 0 _1388_.vdd
rlabel metal2 693 3673 707 3687 0 _1388_.A
rlabel metal2 673 3693 687 3707 0 _1388_.B
rlabel metal2 633 3713 647 3727 0 _1388_.Y
rlabel metal1 1024 3602 1116 3618 0 BUFX2_insert1.gnd
rlabel metal1 1024 3842 1116 3858 0 BUFX2_insert1.vdd
rlabel metal2 1093 3693 1107 3707 0 BUFX2_insert1.A
rlabel metal2 1053 3693 1067 3707 0 BUFX2_insert1.Y
rlabel metal1 1104 3602 1356 3618 0 _1534_.gnd
rlabel metal1 1104 3842 1356 3858 0 _1534_.vdd
rlabel metal2 1253 3693 1267 3707 0 _1534_.D
rlabel metal2 1213 3693 1227 3707 0 _1534_.CLK
rlabel metal2 1133 3693 1147 3707 0 _1534_.Q
rlabel metal1 1604 3602 1696 3618 0 BUFX2_insert5.gnd
rlabel metal1 1604 3842 1696 3858 0 BUFX2_insert5.vdd
rlabel metal2 1613 3693 1627 3707 0 BUFX2_insert5.A
rlabel metal2 1653 3693 1667 3707 0 BUFX2_insert5.Y
rlabel metal1 1344 3602 1456 3618 0 _817_.gnd
rlabel metal1 1344 3842 1456 3858 0 _817_.vdd
rlabel metal2 1353 3693 1367 3707 0 _817_.A
rlabel metal2 1373 3713 1387 3727 0 _817_.B
rlabel metal2 1413 3713 1427 3727 0 _817_.C
rlabel metal2 1393 3693 1407 3707 0 _817_.Y
rlabel metal1 1524 3602 1616 3618 0 _822_.gnd
rlabel metal1 1524 3842 1616 3858 0 _822_.vdd
rlabel metal2 1533 3733 1547 3747 0 _822_.A
rlabel metal2 1573 3733 1587 3747 0 _822_.B
rlabel metal2 1553 3713 1567 3727 0 _822_.Y
rlabel metal1 1444 3602 1536 3618 0 _816_.gnd
rlabel metal1 1444 3842 1536 3858 0 _816_.vdd
rlabel metal2 1453 3733 1467 3747 0 _816_.A
rlabel metal2 1493 3733 1507 3747 0 _816_.B
rlabel metal2 1473 3713 1487 3727 0 _816_.Y
rlabel metal1 1684 3602 1936 3618 0 _1549_.gnd
rlabel metal1 1684 3842 1936 3858 0 _1549_.vdd
rlabel metal2 1833 3693 1847 3707 0 _1549_.D
rlabel metal2 1793 3693 1807 3707 0 _1549_.CLK
rlabel metal2 1713 3693 1727 3707 0 _1549_.Q
rlabel metal1 1984 3602 2096 3618 0 _945_.gnd
rlabel metal1 1984 3842 2096 3858 0 _945_.vdd
rlabel metal2 2073 3713 2087 3727 0 _945_.A
rlabel metal2 2053 3673 2067 3687 0 _945_.B
rlabel metal2 2033 3713 2047 3727 0 _945_.C
rlabel metal2 2013 3693 2027 3707 0 _945_.Y
rlabel metal1 2084 3602 2156 3618 0 _944_.gnd
rlabel metal1 2084 3842 2156 3858 0 _944_.vdd
rlabel metal2 2133 3673 2147 3687 0 _944_.A
rlabel metal2 2113 3713 2127 3727 0 _944_.Y
rlabel metal1 1924 3602 1996 3618 0 _914_.gnd
rlabel metal1 1924 3842 1996 3858 0 _914_.vdd
rlabel metal2 1973 3673 1987 3687 0 _914_.A
rlabel metal2 1953 3713 1967 3727 0 _914_.Y
rlabel metal1 2244 3602 2356 3618 0 _916_.gnd
rlabel metal1 2244 3842 2356 3858 0 _916_.vdd
rlabel metal2 2333 3693 2347 3707 0 _916_.A
rlabel metal2 2313 3713 2327 3727 0 _916_.B
rlabel metal2 2273 3713 2287 3727 0 _916_.C
rlabel metal2 2293 3693 2307 3707 0 _916_.Y
rlabel metal1 2144 3602 2256 3618 0 _908_.gnd
rlabel metal1 2144 3842 2256 3858 0 _908_.vdd
rlabel metal2 2153 3713 2167 3727 0 _908_.A
rlabel metal2 2173 3733 2187 3747 0 _908_.B
rlabel metal2 2193 3713 2207 3727 0 _908_.C
rlabel metal2 2213 3733 2227 3747 0 _908_.Y
rlabel metal1 2344 3602 2456 3618 0 _906_.gnd
rlabel metal1 2344 3842 2456 3858 0 _906_.vdd
rlabel metal2 2433 3713 2447 3727 0 _906_.A
rlabel metal2 2413 3733 2427 3747 0 _906_.B
rlabel metal2 2393 3713 2407 3727 0 _906_.C
rlabel metal2 2373 3733 2387 3747 0 _906_.Y
rlabel metal1 2444 3602 2556 3618 0 _915_.gnd
rlabel metal1 2444 3842 2556 3858 0 _915_.vdd
rlabel metal2 2533 3713 2547 3727 0 _915_.A
rlabel metal2 2513 3673 2527 3687 0 _915_.B
rlabel metal2 2493 3713 2507 3727 0 _915_.C
rlabel metal2 2473 3693 2487 3707 0 _915_.Y
rlabel metal1 2644 3602 2756 3618 0 _896_.gnd
rlabel metal1 2644 3842 2756 3858 0 _896_.vdd
rlabel metal2 2653 3713 2667 3727 0 _896_.A
rlabel metal2 2673 3673 2687 3687 0 _896_.B
rlabel metal2 2693 3713 2707 3727 0 _896_.C
rlabel metal2 2713 3693 2727 3707 0 _896_.Y
rlabel metal1 2544 3602 2656 3618 0 _893_.gnd
rlabel metal1 2544 3842 2656 3858 0 _893_.vdd
rlabel metal2 2633 3713 2647 3727 0 _893_.A
rlabel metal2 2613 3733 2627 3747 0 _893_.B
rlabel metal2 2593 3713 2607 3727 0 _893_.C
rlabel metal2 2573 3733 2587 3747 0 _893_.Y
rlabel metal1 2744 3602 2856 3618 0 _929_.gnd
rlabel metal1 2744 3842 2856 3858 0 _929_.vdd
rlabel metal2 2833 3713 2847 3727 0 _929_.A
rlabel metal2 2813 3673 2827 3687 0 _929_.B
rlabel metal2 2793 3713 2807 3727 0 _929_.C
rlabel metal2 2773 3693 2787 3707 0 _929_.Y
rlabel metal1 2844 3602 2916 3618 0 _892_.gnd
rlabel metal1 2844 3842 2916 3858 0 _892_.vdd
rlabel metal2 2893 3673 2907 3687 0 _892_.A
rlabel metal2 2873 3713 2887 3727 0 _892_.Y
rlabel metal1 2904 3602 2976 3618 0 _889_.gnd
rlabel metal1 2904 3842 2976 3858 0 _889_.vdd
rlabel metal2 2953 3673 2967 3687 0 _889_.A
rlabel metal2 2933 3713 2947 3727 0 _889_.Y
rlabel metal1 3064 3602 3176 3618 0 _928_.gnd
rlabel metal1 3064 3842 3176 3858 0 _928_.vdd
rlabel metal2 3153 3713 3167 3727 0 _928_.A
rlabel metal2 3133 3673 3147 3687 0 _928_.B
rlabel metal2 3113 3713 3127 3727 0 _928_.C
rlabel metal2 3093 3693 3107 3707 0 _928_.Y
rlabel metal1 2964 3602 3076 3618 0 _940_.gnd
rlabel metal1 2964 3842 3076 3858 0 _940_.vdd
rlabel metal2 3053 3713 3067 3727 0 _940_.A
rlabel metal2 3033 3733 3047 3747 0 _940_.B
rlabel metal2 3013 3713 3027 3727 0 _940_.C
rlabel metal2 2993 3733 3007 3747 0 _940_.Y
rlabel metal1 3164 3602 3276 3618 0 _924_.gnd
rlabel metal1 3164 3842 3276 3858 0 _924_.vdd
rlabel metal2 3253 3713 3267 3727 0 _924_.A
rlabel metal2 3233 3733 3247 3747 0 _924_.B
rlabel metal2 3213 3713 3227 3727 0 _924_.C
rlabel metal2 3193 3733 3207 3747 0 _924_.Y
rlabel metal1 3324 3602 3436 3618 0 _927_.gnd
rlabel metal1 3324 3842 3436 3858 0 _927_.vdd
rlabel metal2 3413 3693 3427 3707 0 _927_.A
rlabel metal2 3393 3713 3407 3727 0 _927_.B
rlabel metal2 3353 3713 3367 3727 0 _927_.C
rlabel metal2 3373 3693 3387 3707 0 _927_.Y
rlabel metal1 3424 3602 3516 3618 0 _969_.gnd
rlabel metal1 3424 3842 3516 3858 0 _969_.vdd
rlabel metal2 3493 3733 3507 3747 0 _969_.A
rlabel metal2 3453 3733 3467 3747 0 _969_.B
rlabel metal2 3473 3713 3487 3727 0 _969_.Y
rlabel metal1 3264 3602 3336 3618 0 _923_.gnd
rlabel metal1 3264 3842 3336 3858 0 _923_.vdd
rlabel metal2 3313 3673 3327 3687 0 _923_.A
rlabel metal2 3293 3713 3307 3727 0 _923_.Y
rlabel metal1 3604 3602 3716 3618 0 _983_.gnd
rlabel metal1 3604 3842 3716 3858 0 _983_.vdd
rlabel metal2 3693 3713 3707 3727 0 _983_.A
rlabel metal2 3673 3673 3687 3687 0 _983_.B
rlabel metal2 3653 3713 3667 3727 0 _983_.C
rlabel metal2 3633 3693 3647 3707 0 _983_.Y
rlabel metal1 3704 3602 3816 3618 0 _980_.gnd
rlabel metal1 3704 3842 3816 3858 0 _980_.vdd
rlabel metal2 3793 3713 3807 3727 0 _980_.A
rlabel metal2 3773 3733 3787 3747 0 _980_.B
rlabel metal2 3753 3713 3767 3727 0 _980_.C
rlabel metal2 3733 3733 3747 3747 0 _980_.Y
rlabel metal1 3504 3602 3616 3618 0 _987_.gnd
rlabel metal1 3504 3842 3616 3858 0 _987_.vdd
rlabel metal2 3513 3693 3527 3707 0 _987_.A
rlabel metal2 3573 3693 3587 3707 0 _987_.Y
rlabel metal2 3553 3733 3567 3747 0 _987_.B
rlabel metal1 3964 3602 4076 3618 0 _1047_.gnd
rlabel metal1 3964 3842 4076 3858 0 _1047_.vdd
rlabel metal2 4053 3693 4067 3707 0 _1047_.A
rlabel metal2 4033 3713 4047 3727 0 _1047_.B
rlabel metal2 3993 3713 4007 3727 0 _1047_.C
rlabel metal2 4013 3693 4027 3707 0 _1047_.Y
rlabel metal1 3864 3602 3976 3618 0 _1026_.gnd
rlabel metal1 3864 3842 3976 3858 0 _1026_.vdd
rlabel metal2 3873 3713 3887 3727 0 _1026_.A
rlabel metal2 3893 3673 3907 3687 0 _1026_.B
rlabel metal2 3913 3713 3927 3727 0 _1026_.C
rlabel metal2 3933 3693 3947 3707 0 _1026_.Y
rlabel metal1 3804 3602 3876 3618 0 _977_.gnd
rlabel metal1 3804 3842 3876 3858 0 _977_.vdd
rlabel metal2 3853 3673 3867 3687 0 _977_.A
rlabel metal2 3833 3713 3847 3727 0 _977_.Y
rlabel metal1 4064 3602 4176 3618 0 _1043_.gnd
rlabel metal1 4064 3842 4176 3858 0 _1043_.vdd
rlabel metal2 4073 3693 4087 3707 0 _1043_.A
rlabel metal2 4093 3713 4107 3727 0 _1043_.B
rlabel metal2 4133 3713 4147 3727 0 _1043_.C
rlabel metal2 4113 3693 4127 3707 0 _1043_.Y
rlabel metal1 4164 3602 4276 3618 0 _1053_.gnd
rlabel metal1 4164 3842 4276 3858 0 _1053_.vdd
rlabel metal2 4173 3713 4187 3727 0 _1053_.A
rlabel metal2 4193 3673 4207 3687 0 _1053_.B
rlabel metal2 4213 3713 4227 3727 0 _1053_.C
rlabel metal2 4233 3693 4247 3707 0 _1053_.Y
rlabel metal1 4264 3602 4376 3618 0 _1052_.gnd
rlabel metal1 4264 3842 4376 3858 0 _1052_.vdd
rlabel metal2 4353 3713 4367 3727 0 _1052_.A
rlabel metal2 4333 3673 4347 3687 0 _1052_.B
rlabel metal2 4313 3713 4327 3727 0 _1052_.C
rlabel metal2 4293 3693 4307 3707 0 _1052_.Y
rlabel metal1 4464 3602 4536 3618 0 _1118_.gnd
rlabel metal1 4464 3842 4536 3858 0 _1118_.vdd
rlabel metal2 4513 3673 4527 3687 0 _1118_.A
rlabel metal2 4493 3713 4507 3727 0 _1118_.Y
rlabel metal1 4524 3602 4636 3618 0 _1124_.gnd
rlabel metal1 4524 3842 4636 3858 0 _1124_.vdd
rlabel metal2 4613 3713 4627 3727 0 _1124_.A
rlabel metal2 4593 3733 4607 3747 0 _1124_.B
rlabel metal2 4573 3713 4587 3727 0 _1124_.C
rlabel metal2 4553 3733 4567 3747 0 _1124_.Y
rlabel metal1 4364 3602 4476 3618 0 _1048_.gnd
rlabel metal1 4364 3842 4476 3858 0 _1048_.vdd
rlabel metal2 4373 3713 4387 3727 0 _1048_.A
rlabel metal2 4393 3733 4407 3747 0 _1048_.B
rlabel metal2 4413 3713 4427 3727 0 _1048_.C
rlabel metal2 4433 3733 4447 3747 0 _1048_.Y
rlabel nsubstratencontact 4756 3848 4756 3848 0 FILL71250x54150.vdd
rlabel metal1 4744 3602 4776 3618 0 FILL71250x54150.gnd
rlabel nsubstratencontact 4736 3848 4736 3848 0 FILL70950x54150.vdd
rlabel metal1 4724 3602 4756 3618 0 FILL70950x54150.gnd
rlabel metal1 4624 3602 4736 3618 0 _1117_.gnd
rlabel metal1 4624 3842 4736 3858 0 _1117_.vdd
rlabel metal2 4633 3713 4647 3727 0 _1117_.A
rlabel metal2 4653 3733 4667 3747 0 _1117_.B
rlabel metal2 4673 3713 4687 3727 0 _1117_.C
rlabel metal2 4693 3733 4707 3747 0 _1117_.Y
rlabel metal1 244 4082 356 4098 0 _1357_.gnd
rlabel metal1 244 3842 356 3858 0 _1357_.vdd
rlabel metal2 253 3993 267 4007 0 _1357_.A
rlabel metal2 273 3973 287 3987 0 _1357_.B
rlabel metal2 313 3973 327 3987 0 _1357_.C
rlabel metal2 293 3993 307 4007 0 _1357_.Y
rlabel metal1 4 4082 96 4098 0 _1360_.gnd
rlabel metal1 4 3842 96 3858 0 _1360_.vdd
rlabel metal2 73 3953 87 3967 0 _1360_.A
rlabel metal2 33 3953 47 3967 0 _1360_.B
rlabel metal2 53 3973 67 3987 0 _1360_.Y
rlabel metal1 84 4082 176 4098 0 _1359_.gnd
rlabel metal1 84 3842 176 3858 0 _1359_.vdd
rlabel metal2 153 3953 167 3967 0 _1359_.A
rlabel metal2 113 3953 127 3967 0 _1359_.B
rlabel metal2 133 3973 147 3987 0 _1359_.Y
rlabel metal1 164 4082 256 4098 0 _1358_.gnd
rlabel metal1 164 3842 256 3858 0 _1358_.vdd
rlabel metal2 193 3993 207 4007 0 _1358_.B
rlabel metal2 233 3993 247 4007 0 _1358_.A
rlabel metal2 213 4013 227 4027 0 _1358_.Y
rlabel metal1 464 4082 556 4098 0 _1378_.gnd
rlabel metal1 464 3842 556 3858 0 _1378_.vdd
rlabel metal2 493 3993 507 4007 0 _1378_.B
rlabel metal2 533 3993 547 4007 0 _1378_.A
rlabel metal2 513 4013 527 4027 0 _1378_.Y
rlabel metal1 404 4082 476 4098 0 _1379_.gnd
rlabel metal1 404 3842 476 3858 0 _1379_.vdd
rlabel metal2 453 4013 467 4027 0 _1379_.A
rlabel metal2 433 3973 447 3987 0 _1379_.Y
rlabel metal1 344 4082 416 4098 0 _1356_.gnd
rlabel metal1 344 3842 416 3858 0 _1356_.vdd
rlabel metal2 393 4013 407 4027 0 _1356_.A
rlabel metal2 373 3973 387 3987 0 _1356_.Y
rlabel metal1 644 4082 756 4098 0 _1384_.gnd
rlabel metal1 644 3842 756 3858 0 _1384_.vdd
rlabel metal2 653 3993 667 4007 0 _1384_.A
rlabel metal2 673 3973 687 3987 0 _1384_.B
rlabel metal2 713 3973 727 3987 0 _1384_.C
rlabel metal2 693 3993 707 4007 0 _1384_.Y
rlabel metal1 744 4082 816 4098 0 _1383_.gnd
rlabel metal1 744 3842 816 3858 0 _1383_.vdd
rlabel metal2 753 4013 767 4027 0 _1383_.A
rlabel metal2 773 3973 787 3987 0 _1383_.Y
rlabel metal1 544 4082 656 4098 0 _1396_.gnd
rlabel metal1 544 3842 656 3858 0 _1396_.vdd
rlabel metal2 553 3993 567 4007 0 _1396_.A
rlabel metal2 613 3993 627 4007 0 _1396_.Y
rlabel metal2 593 3953 607 3967 0 _1396_.B
rlabel metal1 804 4082 916 4098 0 _826_.gnd
rlabel metal1 804 3842 916 3858 0 _826_.vdd
rlabel metal2 813 3993 827 4007 0 _826_.A
rlabel metal2 833 3973 847 3987 0 _826_.B
rlabel metal2 873 3973 887 3987 0 _826_.C
rlabel metal2 853 3993 867 4007 0 _826_.Y
rlabel metal1 904 4082 996 4098 0 _825_.gnd
rlabel metal1 904 3842 996 3858 0 _825_.vdd
rlabel metal2 913 3953 927 3967 0 _825_.A
rlabel metal2 953 3953 967 3967 0 _825_.B
rlabel metal2 933 3973 947 3987 0 _825_.Y
rlabel metal1 1044 4082 1136 4098 0 _1353_.gnd
rlabel metal1 1044 3842 1136 3858 0 _1353_.vdd
rlabel metal2 1073 3993 1087 4007 0 _1353_.B
rlabel metal2 1113 3993 1127 4007 0 _1353_.A
rlabel metal2 1093 4013 1107 4027 0 _1353_.Y
rlabel metal1 984 4082 1056 4098 0 _824_.gnd
rlabel metal1 984 3842 1056 3858 0 _824_.vdd
rlabel metal2 1033 4013 1047 4027 0 _824_.A
rlabel metal2 1013 3973 1027 3987 0 _824_.Y
rlabel metal1 1324 4082 1416 4098 0 _1377_.gnd
rlabel metal1 1324 3842 1416 3858 0 _1377_.vdd
rlabel metal2 1353 3993 1367 4007 0 _1377_.B
rlabel metal2 1393 3993 1407 4007 0 _1377_.A
rlabel metal2 1373 4013 1387 4027 0 _1377_.Y
rlabel metal1 1184 4082 1276 4098 0 _1354_.gnd
rlabel metal1 1184 3842 1276 3858 0 _1354_.vdd
rlabel metal2 1233 3993 1247 4007 0 _1354_.B
rlabel metal2 1193 3993 1207 4007 0 _1354_.A
rlabel metal2 1213 4013 1227 4027 0 _1354_.Y
rlabel metal1 1264 4082 1336 4098 0 _913_.gnd
rlabel metal1 1264 3842 1336 3858 0 _913_.vdd
rlabel metal2 1273 4013 1287 4027 0 _913_.A
rlabel metal2 1293 3973 1307 3987 0 _913_.Y
rlabel metal1 1124 4082 1196 4098 0 _815_.gnd
rlabel metal1 1124 3842 1196 3858 0 _815_.vdd
rlabel metal2 1133 4013 1147 4027 0 _815_.A
rlabel metal2 1153 3973 1167 3987 0 _815_.Y
rlabel metal1 1464 4082 1576 4098 0 _823_.gnd
rlabel metal1 1464 3842 1576 3858 0 _823_.vdd
rlabel metal2 1473 3993 1487 4007 0 _823_.A
rlabel metal2 1493 3973 1507 3987 0 _823_.B
rlabel metal2 1533 3973 1547 3987 0 _823_.C
rlabel metal2 1513 3993 1527 4007 0 _823_.Y
rlabel metal1 1404 4082 1476 4098 0 _821_.gnd
rlabel metal1 1404 3842 1476 3858 0 _821_.vdd
rlabel metal2 1453 4013 1467 4027 0 _821_.A
rlabel metal2 1433 3973 1447 3987 0 _821_.Y
rlabel metal1 1564 4082 1696 4098 0 _952_.gnd
rlabel metal1 1564 3842 1696 3858 0 _952_.vdd
rlabel metal2 1573 3993 1587 4007 0 _952_.A
rlabel metal2 1593 3973 1607 3987 0 _952_.B
rlabel metal2 1653 3993 1667 4007 0 _952_.C
rlabel metal2 1613 3993 1627 4007 0 _952_.Y
rlabel metal2 1633 3973 1647 3987 0 _952_.D
rlabel metal1 1684 4082 1776 4098 0 _951_.gnd
rlabel metal1 1684 3842 1776 3858 0 _951_.vdd
rlabel metal2 1693 3953 1707 3967 0 _951_.A
rlabel metal2 1733 3953 1747 3967 0 _951_.B
rlabel metal2 1713 3973 1727 3987 0 _951_.Y
rlabel metal1 1764 4082 1876 4098 0 _949_.gnd
rlabel metal1 1764 3842 1876 3858 0 _949_.vdd
rlabel metal2 1853 3973 1867 3987 0 _949_.A
rlabel metal2 1833 4013 1847 4027 0 _949_.B
rlabel metal2 1813 3973 1827 3987 0 _949_.C
rlabel metal2 1793 3993 1807 4007 0 _949_.Y
rlabel metal1 1864 4082 1976 4098 0 _950_.gnd
rlabel metal1 1864 3842 1976 3858 0 _950_.vdd
rlabel metal2 1873 3973 1887 3987 0 _950_.A
rlabel metal2 1893 3953 1907 3967 0 _950_.B
rlabel metal2 1913 3973 1927 3987 0 _950_.C
rlabel metal2 1933 3953 1947 3967 0 _950_.Y
rlabel metal1 1964 4082 2076 4098 0 _948_.gnd
rlabel metal1 1964 3842 2076 3858 0 _948_.vdd
rlabel metal2 2053 3993 2067 4007 0 _948_.A
rlabel metal2 2033 3973 2047 3987 0 _948_.B
rlabel metal2 1993 3973 2007 3987 0 _948_.C
rlabel metal2 2013 3993 2027 4007 0 _948_.Y
rlabel metal1 2064 4082 2136 4098 0 _947_.gnd
rlabel metal1 2064 3842 2136 3858 0 _947_.vdd
rlabel metal2 2113 4013 2127 4027 0 _947_.A
rlabel metal2 2093 3973 2107 3987 0 _947_.Y
rlabel metal1 2124 4082 2236 4098 0 _943_.gnd
rlabel metal1 2124 3842 2236 3858 0 _943_.vdd
rlabel metal2 2213 3973 2227 3987 0 _943_.A
rlabel metal2 2193 3953 2207 3967 0 _943_.B
rlabel metal2 2173 3973 2187 3987 0 _943_.C
rlabel metal2 2153 3953 2167 3967 0 _943_.Y
rlabel metal1 2324 4082 2436 4098 0 _946_.gnd
rlabel metal1 2324 3842 2436 3858 0 _946_.vdd
rlabel metal2 2413 3973 2427 3987 0 _946_.A
rlabel metal2 2393 4013 2407 4027 0 _946_.B
rlabel metal2 2373 3973 2387 3987 0 _946_.C
rlabel metal2 2353 3993 2367 4007 0 _946_.Y
rlabel metal1 2224 4082 2336 4098 0 _942_.gnd
rlabel metal1 2224 3842 2336 3858 0 _942_.vdd
rlabel metal2 2313 3973 2327 3987 0 _942_.A
rlabel metal2 2293 3953 2307 3967 0 _942_.B
rlabel metal2 2273 3973 2287 3987 0 _942_.C
rlabel metal2 2253 3953 2267 3967 0 _942_.Y
rlabel metal1 2484 4082 2596 4098 0 _938_.gnd
rlabel metal1 2484 3842 2596 3858 0 _938_.vdd
rlabel metal2 2573 3993 2587 4007 0 _938_.A
rlabel metal2 2553 3973 2567 3987 0 _938_.B
rlabel metal2 2513 3973 2527 3987 0 _938_.C
rlabel metal2 2533 3993 2547 4007 0 _938_.Y
rlabel metal1 2424 4082 2496 4098 0 _941_.gnd
rlabel metal1 2424 3842 2496 3858 0 _941_.vdd
rlabel metal2 2473 4013 2487 4027 0 _941_.A
rlabel metal2 2453 3973 2467 3987 0 _941_.Y
rlabel metal1 2584 4082 2696 4098 0 _939_.gnd
rlabel metal1 2584 3842 2696 3858 0 _939_.vdd
rlabel metal2 2673 3973 2687 3987 0 _939_.A
rlabel metal2 2653 3953 2667 3967 0 _939_.B
rlabel metal2 2633 3973 2647 3987 0 _939_.C
rlabel metal2 2613 3953 2627 3967 0 _939_.Y
rlabel metal1 2884 4082 2996 4098 0 _1139_.gnd
rlabel metal1 2884 3842 2996 3858 0 _1139_.vdd
rlabel metal2 2893 3993 2907 4007 0 _1139_.A
rlabel metal2 2913 3973 2927 3987 0 _1139_.B
rlabel metal2 2953 3973 2967 3987 0 _1139_.C
rlabel metal2 2933 3993 2947 4007 0 _1139_.Y
rlabel metal1 2784 4082 2896 4098 0 _992_.gnd
rlabel metal1 2784 3842 2896 3858 0 _992_.vdd
rlabel metal2 2873 3993 2887 4007 0 _992_.A
rlabel metal2 2853 3973 2867 3987 0 _992_.B
rlabel metal2 2813 3973 2827 3987 0 _992_.C
rlabel metal2 2833 3993 2847 4007 0 _992_.Y
rlabel metal1 2684 4082 2796 4098 0 _932_.gnd
rlabel metal1 2684 3842 2796 3858 0 _932_.vdd
rlabel metal2 2773 3973 2787 3987 0 _932_.A
rlabel metal2 2753 4013 2767 4027 0 _932_.B
rlabel metal2 2733 3973 2747 3987 0 _932_.C
rlabel metal2 2713 3993 2727 4007 0 _932_.Y
rlabel metal1 3144 4082 3256 4098 0 _931_.gnd
rlabel metal1 3144 3842 3256 3858 0 _931_.vdd
rlabel metal2 3153 3993 3167 4007 0 _931_.A
rlabel metal2 3173 3973 3187 3987 0 _931_.B
rlabel metal2 3213 3973 3227 3987 0 _931_.C
rlabel metal2 3193 3993 3207 4007 0 _931_.Y
rlabel metal1 3084 4082 3156 4098 0 _921_.gnd
rlabel metal1 3084 3842 3156 3858 0 _921_.vdd
rlabel metal2 3133 4013 3147 4027 0 _921_.A
rlabel metal2 3113 3973 3127 3987 0 _921_.Y
rlabel metal1 2984 4082 3096 4098 0 _930_.gnd
rlabel metal1 2984 3842 3096 3858 0 _930_.vdd
rlabel metal2 3073 3973 3087 3987 0 _930_.A
rlabel metal2 3053 3953 3067 3967 0 _930_.B
rlabel metal2 3033 3973 3047 3987 0 _930_.C
rlabel metal2 3013 3953 3027 3967 0 _930_.Y
rlabel metal1 3444 4082 3556 4098 0 _985_.gnd
rlabel metal1 3444 3842 3556 3858 0 _985_.vdd
rlabel metal2 3533 3993 3547 4007 0 _985_.A
rlabel metal2 3513 3973 3527 3987 0 _985_.B
rlabel metal2 3473 3973 3487 3987 0 _985_.C
rlabel metal2 3493 3993 3507 4007 0 _985_.Y
rlabel metal1 3344 4082 3456 4098 0 _982_.gnd
rlabel metal1 3344 3842 3456 3858 0 _982_.vdd
rlabel metal2 3353 3993 3367 4007 0 _982_.A
rlabel metal2 3373 3973 3387 3987 0 _982_.B
rlabel metal2 3413 3973 3427 3987 0 _982_.C
rlabel metal2 3393 3993 3407 4007 0 _982_.Y
rlabel metal1 3244 4082 3356 4098 0 _970_.gnd
rlabel metal1 3244 3842 3356 3858 0 _970_.vdd
rlabel metal2 3253 3973 3267 3987 0 _970_.A
rlabel metal2 3273 4013 3287 4027 0 _970_.B
rlabel metal2 3293 3973 3307 3987 0 _970_.C
rlabel metal2 3313 3993 3327 4007 0 _970_.Y
rlabel metal1 3544 4082 3656 4098 0 _989_.gnd
rlabel metal1 3544 3842 3656 3858 0 _989_.vdd
rlabel metal2 3633 3993 3647 4007 0 _989_.A
rlabel metal2 3613 3973 3627 3987 0 _989_.B
rlabel metal2 3573 3973 3587 3987 0 _989_.C
rlabel metal2 3593 3993 3607 4007 0 _989_.Y
rlabel metal1 3644 4082 3756 4098 0 _984_.gnd
rlabel metal1 3644 3842 3756 3858 0 _984_.vdd
rlabel metal2 3733 3973 3747 3987 0 _984_.A
rlabel metal2 3713 4013 3727 4027 0 _984_.B
rlabel metal2 3693 3973 3707 3987 0 _984_.C
rlabel metal2 3673 3993 3687 4007 0 _984_.Y
rlabel metal1 3844 4082 3936 4098 0 _1138_.gnd
rlabel metal1 3844 3842 3936 3858 0 _1138_.vdd
rlabel metal2 3913 3953 3927 3967 0 _1138_.A
rlabel metal2 3873 3953 3887 3967 0 _1138_.B
rlabel metal2 3893 3973 3907 3987 0 _1138_.Y
rlabel metal1 3924 4082 4016 4098 0 _1137_.gnd
rlabel metal1 3924 3842 4016 3858 0 _1137_.vdd
rlabel metal2 3993 3953 4007 3967 0 _1137_.A
rlabel metal2 3953 3953 3967 3967 0 _1137_.B
rlabel metal2 3973 3973 3987 3987 0 _1137_.Y
rlabel metal1 4004 4082 4096 4098 0 _1132_.gnd
rlabel metal1 4004 3842 4096 3858 0 _1132_.vdd
rlabel metal2 4013 3953 4027 3967 0 _1132_.A
rlabel metal2 4053 3953 4067 3967 0 _1132_.B
rlabel metal2 4033 3973 4047 3987 0 _1132_.Y
rlabel metal1 3744 4082 3856 4098 0 _976_.gnd
rlabel metal1 3744 3842 3856 3858 0 _976_.vdd
rlabel metal2 3833 3973 3847 3987 0 _976_.A
rlabel metal2 3813 3953 3827 3967 0 _976_.B
rlabel metal2 3793 3973 3807 3987 0 _976_.C
rlabel metal2 3773 3953 3787 3967 0 _976_.Y
rlabel metal1 4184 4082 4296 4098 0 _1054_.gnd
rlabel metal1 4184 3842 4296 3858 0 _1054_.vdd
rlabel metal2 4273 3993 4287 4007 0 _1054_.A
rlabel metal2 4253 3973 4267 3987 0 _1054_.B
rlabel metal2 4213 3973 4227 3987 0 _1054_.C
rlabel metal2 4233 3993 4247 4007 0 _1054_.Y
rlabel metal1 4084 4082 4196 4098 0 _1044_.gnd
rlabel metal1 4084 3842 4196 3858 0 _1044_.vdd
rlabel metal2 4173 3973 4187 3987 0 _1044_.A
rlabel metal2 4153 3953 4167 3967 0 _1044_.B
rlabel metal2 4133 3973 4147 3987 0 _1044_.C
rlabel metal2 4113 3953 4127 3967 0 _1044_.Y
rlabel metal1 4284 4082 4396 4098 0 _1057_.gnd
rlabel metal1 4284 3842 4396 3858 0 _1057_.vdd
rlabel metal2 4293 3993 4307 4007 0 _1057_.A
rlabel metal2 4313 3973 4327 3987 0 _1057_.B
rlabel metal2 4353 3973 4367 3987 0 _1057_.C
rlabel metal2 4333 3993 4347 4007 0 _1057_.Y
rlabel metal1 4384 4082 4456 4098 0 _1129_.gnd
rlabel metal1 4384 3842 4456 3858 0 _1129_.vdd
rlabel metal2 4433 4013 4447 4027 0 _1129_.A
rlabel metal2 4413 3973 4427 3987 0 _1129_.Y
rlabel metal1 4444 4082 4556 4098 0 _1130_.gnd
rlabel metal1 4444 3842 4556 3858 0 _1130_.vdd
rlabel metal2 4533 3973 4547 3987 0 _1130_.A
rlabel metal2 4513 3953 4527 3967 0 _1130_.B
rlabel metal2 4493 3973 4507 3987 0 _1130_.C
rlabel metal2 4473 3953 4487 3967 0 _1130_.Y
rlabel nsubstratencontact 4764 3852 4764 3852 0 FILL71250x57750.vdd
rlabel metal1 4744 4082 4776 4098 0 FILL71250x57750.gnd
rlabel metal1 4644 4082 4756 4098 0 _1122_.gnd
rlabel metal1 4644 3842 4756 3858 0 _1122_.vdd
rlabel metal2 4653 3973 4667 3987 0 _1122_.A
rlabel metal2 4673 4013 4687 4027 0 _1122_.B
rlabel metal2 4693 3973 4707 3987 0 _1122_.C
rlabel metal2 4713 3993 4727 4007 0 _1122_.Y
rlabel metal1 4544 4082 4656 4098 0 _1131_.gnd
rlabel metal1 4544 3842 4656 3858 0 _1131_.vdd
rlabel metal2 4633 3973 4647 3987 0 _1131_.A
rlabel metal2 4613 3953 4627 3967 0 _1131_.B
rlabel metal2 4593 3973 4607 3987 0 _1131_.C
rlabel metal2 4573 3953 4587 3967 0 _1131_.Y
rlabel metal1 4 4082 116 4098 0 _1369_.gnd
rlabel metal1 4 4322 116 4338 0 _1369_.vdd
rlabel metal2 93 4173 107 4187 0 _1369_.A
rlabel metal2 73 4193 87 4207 0 _1369_.B
rlabel metal2 33 4193 47 4207 0 _1369_.C
rlabel metal2 53 4173 67 4187 0 _1369_.Y
rlabel metal1 204 4082 296 4098 0 _1368_.gnd
rlabel metal1 204 4322 296 4338 0 _1368_.vdd
rlabel metal2 253 4173 267 4187 0 _1368_.B
rlabel metal2 213 4173 227 4187 0 _1368_.A
rlabel metal2 233 4153 247 4167 0 _1368_.Y
rlabel metal1 104 4082 216 4098 0 _1367_.gnd
rlabel metal1 104 4322 216 4338 0 _1367_.vdd
rlabel metal2 193 4173 207 4187 0 _1367_.A
rlabel metal2 133 4173 147 4187 0 _1367_.Y
rlabel metal2 153 4213 167 4227 0 _1367_.B
rlabel metal1 484 4082 596 4098 0 _1375_.gnd
rlabel metal1 484 4322 596 4338 0 _1375_.vdd
rlabel metal2 573 4193 587 4207 0 _1375_.A
rlabel metal2 553 4153 567 4167 0 _1375_.B
rlabel metal2 533 4193 547 4207 0 _1375_.C
rlabel metal2 513 4173 527 4187 0 _1375_.Y
rlabel metal1 284 4082 396 4098 0 _1363_.gnd
rlabel metal1 284 4322 396 4338 0 _1363_.vdd
rlabel metal2 373 4193 387 4207 0 _1363_.A
rlabel metal2 353 4153 367 4167 0 _1363_.B
rlabel metal2 333 4193 347 4207 0 _1363_.C
rlabel metal2 313 4173 327 4187 0 _1363_.Y
rlabel metal1 384 4082 496 4098 0 _1374_.gnd
rlabel metal1 384 4322 496 4338 0 _1374_.vdd
rlabel metal2 393 4173 407 4187 0 _1374_.A
rlabel metal2 453 4173 467 4187 0 _1374_.Y
rlabel metal2 433 4213 447 4227 0 _1374_.B
rlabel metal1 684 4082 796 4098 0 _1397_.gnd
rlabel metal1 684 4322 796 4338 0 _1397_.vdd
rlabel metal2 693 4193 707 4207 0 _1397_.A
rlabel metal2 713 4153 727 4167 0 _1397_.B
rlabel metal2 733 4193 747 4207 0 _1397_.C
rlabel metal2 753 4173 767 4187 0 _1397_.Y
rlabel metal1 584 4082 696 4098 0 _1398_.gnd
rlabel metal1 584 4322 696 4338 0 _1398_.vdd
rlabel metal2 593 4193 607 4207 0 _1398_.A
rlabel metal2 613 4213 627 4227 0 _1398_.B
rlabel metal2 633 4193 647 4207 0 _1398_.C
rlabel metal2 653 4213 667 4227 0 _1398_.Y
rlabel metal1 784 4082 896 4098 0 _1399_.gnd
rlabel metal1 784 4322 896 4338 0 _1399_.vdd
rlabel metal2 793 4173 807 4187 0 _1399_.A
rlabel metal2 853 4173 867 4187 0 _1399_.Y
rlabel metal2 833 4213 847 4227 0 _1399_.B
rlabel metal1 884 4082 996 4098 0 _1395_.gnd
rlabel metal1 884 4322 996 4338 0 _1395_.vdd
rlabel metal2 973 4173 987 4187 0 _1395_.A
rlabel metal2 953 4193 967 4207 0 _1395_.B
rlabel metal2 913 4193 927 4207 0 _1395_.C
rlabel metal2 933 4173 947 4187 0 _1395_.Y
rlabel metal1 1044 4082 1136 4098 0 _1387_.gnd
rlabel metal1 1044 4322 1136 4338 0 _1387_.vdd
rlabel metal2 1093 4173 1107 4187 0 _1387_.B
rlabel metal2 1053 4173 1067 4187 0 _1387_.A
rlabel metal2 1073 4153 1087 4167 0 _1387_.Y
rlabel metal1 984 4082 1056 4098 0 _1394_.gnd
rlabel metal1 984 4322 1056 4338 0 _1394_.vdd
rlabel metal2 1033 4153 1047 4167 0 _1394_.A
rlabel metal2 1013 4193 1027 4207 0 _1394_.Y
rlabel metal1 1124 4082 1216 4098 0 _1386_.gnd
rlabel metal1 1124 4322 1216 4338 0 _1386_.vdd
rlabel metal2 1173 4173 1187 4187 0 _1386_.B
rlabel metal2 1133 4173 1147 4187 0 _1386_.A
rlabel metal2 1153 4153 1167 4167 0 _1386_.Y
rlabel metal1 1204 4082 1296 4098 0 _1385_.gnd
rlabel metal1 1204 4322 1296 4338 0 _1385_.vdd
rlabel metal2 1253 4173 1267 4187 0 _1385_.B
rlabel metal2 1213 4173 1227 4187 0 _1385_.A
rlabel metal2 1233 4153 1247 4167 0 _1385_.Y
rlabel metal1 1284 4082 1356 4098 0 _1070_.gnd
rlabel metal1 1284 4322 1356 4338 0 _1070_.vdd
rlabel metal2 1293 4153 1307 4167 0 _1070_.A
rlabel metal2 1313 4193 1327 4207 0 _1070_.Y
rlabel metal1 1344 4082 1596 4098 0 _1553_.gnd
rlabel metal1 1344 4322 1596 4338 0 _1553_.vdd
rlabel metal2 1493 4173 1507 4187 0 _1553_.D
rlabel metal2 1453 4173 1467 4187 0 _1553_.CLK
rlabel metal2 1373 4173 1387 4187 0 _1553_.Q
rlabel metal1 1584 4082 1696 4098 0 _1135_.gnd
rlabel metal1 1584 4322 1696 4338 0 _1135_.vdd
rlabel metal2 1593 4173 1607 4187 0 _1135_.A
rlabel metal2 1613 4193 1627 4207 0 _1135_.B
rlabel metal2 1653 4193 1667 4207 0 _1135_.C
rlabel metal2 1633 4173 1647 4187 0 _1135_.Y
rlabel metal1 1824 4082 2076 4098 0 _1550_.gnd
rlabel metal1 1824 4322 2076 4338 0 _1550_.vdd
rlabel metal2 1973 4173 1987 4187 0 _1550_.D
rlabel metal2 1933 4173 1947 4187 0 _1550_.CLK
rlabel metal2 1853 4173 1867 4187 0 _1550_.Q
rlabel metal1 1684 4082 1776 4098 0 _1376_.gnd
rlabel metal1 1684 4322 1776 4338 0 _1376_.vdd
rlabel metal2 1733 4173 1747 4187 0 _1376_.B
rlabel metal2 1693 4173 1707 4187 0 _1376_.A
rlabel metal2 1713 4153 1727 4167 0 _1376_.Y
rlabel metal1 1764 4082 1836 4098 0 _1006_.gnd
rlabel metal1 1764 4322 1836 4338 0 _1006_.vdd
rlabel metal2 1813 4153 1827 4167 0 _1006_.A
rlabel metal2 1793 4193 1807 4207 0 _1006_.Y
rlabel metal1 2064 4082 2156 4098 0 _1000_.gnd
rlabel metal1 2064 4322 2156 4338 0 _1000_.vdd
rlabel metal2 2133 4213 2147 4227 0 _1000_.A
rlabel metal2 2093 4213 2107 4227 0 _1000_.B
rlabel metal2 2113 4193 2127 4207 0 _1000_.Y
rlabel metal1 2364 4082 2456 4098 0 _999_.gnd
rlabel metal1 2364 4322 2456 4338 0 _999_.vdd
rlabel metal2 2373 4213 2387 4227 0 _999_.A
rlabel metal2 2413 4213 2427 4227 0 _999_.B
rlabel metal2 2393 4193 2407 4207 0 _999_.Y
rlabel metal1 2244 4082 2376 4098 0 _1002_.gnd
rlabel metal1 2244 4322 2376 4338 0 _1002_.vdd
rlabel metal2 2353 4173 2367 4187 0 _1002_.A
rlabel metal2 2333 4193 2347 4207 0 _1002_.B
rlabel metal2 2273 4173 2287 4187 0 _1002_.C
rlabel metal2 2293 4193 2307 4207 0 _1002_.D
rlabel metal2 2313 4173 2327 4187 0 _1002_.Y
rlabel metal1 2144 4082 2256 4098 0 _1001_.gnd
rlabel metal1 2144 4322 2256 4338 0 _1001_.vdd
rlabel metal2 2153 4153 2167 4167 0 _1001_.A
rlabel metal2 2173 4173 2187 4187 0 _1001_.B
rlabel metal2 2213 4193 2227 4207 0 _1001_.Y
rlabel metal1 2444 4082 2556 4098 0 _1134_.gnd
rlabel metal1 2444 4322 2556 4338 0 _1134_.vdd
rlabel metal2 2533 4173 2547 4187 0 _1134_.A
rlabel metal2 2513 4193 2527 4207 0 _1134_.B
rlabel metal2 2473 4193 2487 4207 0 _1134_.C
rlabel metal2 2493 4173 2507 4187 0 _1134_.Y
rlabel metal1 2624 4082 2736 4098 0 _957_.gnd
rlabel metal1 2624 4322 2736 4338 0 _957_.vdd
rlabel metal2 2633 4193 2647 4207 0 _957_.A
rlabel metal2 2653 4153 2667 4167 0 _957_.B
rlabel metal2 2673 4193 2687 4207 0 _957_.C
rlabel metal2 2693 4173 2707 4187 0 _957_.Y
rlabel metal1 2544 4082 2636 4098 0 _1133_.gnd
rlabel metal1 2544 4322 2636 4338 0 _1133_.vdd
rlabel metal2 2573 4173 2587 4187 0 _1133_.B
rlabel metal2 2613 4173 2627 4187 0 _1133_.A
rlabel metal2 2593 4153 2607 4167 0 _1133_.Y
rlabel metal1 2824 4082 2916 4098 0 _1603_.gnd
rlabel metal1 2824 4322 2916 4338 0 _1603_.vdd
rlabel metal2 2833 4173 2847 4187 0 _1603_.A
rlabel metal2 2873 4173 2887 4187 0 _1603_.Y
rlabel metal1 2724 4082 2836 4098 0 _1127_.gnd
rlabel metal1 2724 4322 2836 4338 0 _1127_.vdd
rlabel metal2 2813 4193 2827 4207 0 _1127_.A
rlabel metal2 2793 4153 2807 4167 0 _1127_.B
rlabel metal2 2773 4193 2787 4207 0 _1127_.C
rlabel metal2 2753 4173 2767 4187 0 _1127_.Y
rlabel metal1 2904 4082 3016 4098 0 _1269_.gnd
rlabel metal1 2904 4322 3016 4338 0 _1269_.vdd
rlabel metal2 2993 4193 3007 4207 0 _1269_.A
rlabel metal2 2973 4213 2987 4227 0 _1269_.B
rlabel metal2 2953 4193 2967 4207 0 _1269_.C
rlabel metal2 2933 4213 2947 4227 0 _1269_.Y
rlabel metal1 3104 4082 3196 4098 0 _994_.gnd
rlabel metal1 3104 4322 3196 4338 0 _994_.vdd
rlabel metal2 3113 4213 3127 4227 0 _994_.A
rlabel metal2 3153 4213 3167 4227 0 _994_.B
rlabel metal2 3133 4193 3147 4207 0 _994_.Y
rlabel metal1 3184 4082 3256 4098 0 _956_.gnd
rlabel metal1 3184 4322 3256 4338 0 _956_.vdd
rlabel metal2 3233 4153 3247 4167 0 _956_.A
rlabel metal2 3213 4193 3227 4207 0 _956_.Y
rlabel metal1 3004 4082 3116 4098 0 _995_.gnd
rlabel metal1 3004 4322 3116 4338 0 _995_.vdd
rlabel metal2 3093 4193 3107 4207 0 _995_.A
rlabel metal2 3073 4213 3087 4227 0 _995_.B
rlabel metal2 3053 4193 3067 4207 0 _995_.C
rlabel metal2 3033 4213 3047 4227 0 _995_.Y
rlabel metal1 3244 4082 3356 4098 0 _991_.gnd
rlabel metal1 3244 4322 3356 4338 0 _991_.vdd
rlabel metal2 3333 4193 3347 4207 0 _991_.A
rlabel metal2 3313 4213 3327 4227 0 _991_.B
rlabel metal2 3293 4193 3307 4207 0 _991_.C
rlabel metal2 3273 4213 3287 4227 0 _991_.Y
rlabel metal1 3344 4082 3456 4098 0 _986_.gnd
rlabel metal1 3344 4322 3456 4338 0 _986_.vdd
rlabel metal2 3433 4193 3447 4207 0 _986_.A
rlabel metal2 3413 4213 3427 4227 0 _986_.B
rlabel metal2 3393 4193 3407 4207 0 _986_.C
rlabel metal2 3373 4213 3387 4227 0 _986_.Y
rlabel metal1 3444 4082 3556 4098 0 _981_.gnd
rlabel metal1 3444 4322 3556 4338 0 _981_.vdd
rlabel metal2 3533 4193 3547 4207 0 _981_.A
rlabel metal2 3513 4213 3527 4227 0 _981_.B
rlabel metal2 3493 4193 3507 4207 0 _981_.C
rlabel metal2 3473 4213 3487 4227 0 _981_.Y
rlabel metal1 3544 4082 3656 4098 0 _990_.gnd
rlabel metal1 3544 4322 3656 4338 0 _990_.vdd
rlabel metal2 3633 4193 3647 4207 0 _990_.A
rlabel metal2 3613 4213 3627 4227 0 _990_.B
rlabel metal2 3593 4193 3607 4207 0 _990_.C
rlabel metal2 3573 4213 3587 4227 0 _990_.Y
rlabel metal1 3644 4082 3756 4098 0 _988_.gnd
rlabel metal1 3644 4322 3756 4338 0 _988_.vdd
rlabel metal2 3653 4193 3667 4207 0 _988_.A
rlabel metal2 3673 4213 3687 4227 0 _988_.B
rlabel metal2 3693 4193 3707 4207 0 _988_.C
rlabel metal2 3713 4213 3727 4227 0 _988_.Y
rlabel metal1 3844 4082 3956 4098 0 _1051_.gnd
rlabel metal1 3844 4322 3956 4338 0 _1051_.vdd
rlabel metal2 3853 4173 3867 4187 0 _1051_.A
rlabel metal2 3873 4193 3887 4207 0 _1051_.B
rlabel metal2 3913 4193 3927 4207 0 _1051_.C
rlabel metal2 3893 4173 3907 4187 0 _1051_.Y
rlabel metal1 3744 4082 3856 4098 0 _1050_.gnd
rlabel metal1 3744 4322 3856 4338 0 _1050_.vdd
rlabel metal2 3753 4193 3767 4207 0 _1050_.A
rlabel metal2 3773 4153 3787 4167 0 _1050_.B
rlabel metal2 3793 4193 3807 4207 0 _1050_.C
rlabel metal2 3813 4173 3827 4187 0 _1050_.Y
rlabel metal1 4004 4082 4116 4098 0 _1013_.gnd
rlabel metal1 4004 4322 4116 4338 0 _1013_.vdd
rlabel metal2 4013 4193 4027 4207 0 _1013_.A
rlabel metal2 4033 4153 4047 4167 0 _1013_.B
rlabel metal2 4053 4193 4067 4207 0 _1013_.C
rlabel metal2 4073 4173 4087 4187 0 _1013_.Y
rlabel metal1 3944 4082 4016 4098 0 _1012_.gnd
rlabel metal1 3944 4322 4016 4338 0 _1012_.vdd
rlabel metal2 3953 4153 3967 4167 0 _1012_.A
rlabel metal2 3973 4193 3987 4207 0 _1012_.Y
rlabel metal1 4204 4082 4316 4098 0 _1056_.gnd
rlabel metal1 4204 4322 4316 4338 0 _1056_.vdd
rlabel metal2 4213 4193 4227 4207 0 _1056_.A
rlabel metal2 4233 4213 4247 4227 0 _1056_.B
rlabel metal2 4253 4193 4267 4207 0 _1056_.C
rlabel metal2 4273 4213 4287 4227 0 _1056_.Y
rlabel metal1 4104 4082 4216 4098 0 _1049_.gnd
rlabel metal1 4104 4322 4216 4338 0 _1049_.vdd
rlabel metal2 4193 4193 4207 4207 0 _1049_.A
rlabel metal2 4173 4213 4187 4227 0 _1049_.B
rlabel metal2 4153 4193 4167 4207 0 _1049_.C
rlabel metal2 4133 4213 4147 4227 0 _1049_.Y
rlabel metal1 4404 4082 4516 4098 0 _1073_.gnd
rlabel metal1 4404 4322 4516 4338 0 _1073_.vdd
rlabel metal2 4413 4173 4427 4187 0 _1073_.A
rlabel metal2 4433 4193 4447 4207 0 _1073_.B
rlabel metal2 4473 4193 4487 4207 0 _1073_.C
rlabel metal2 4453 4173 4467 4187 0 _1073_.Y
rlabel metal1 4304 4082 4416 4098 0 _1072_.gnd
rlabel metal1 4304 4322 4416 4338 0 _1072_.vdd
rlabel metal2 4313 4193 4327 4207 0 _1072_.A
rlabel metal2 4333 4153 4347 4167 0 _1072_.B
rlabel metal2 4353 4193 4367 4207 0 _1072_.C
rlabel metal2 4373 4173 4387 4187 0 _1072_.Y
rlabel metal1 4504 4082 4636 4098 0 _1125_.gnd
rlabel metal1 4504 4322 4636 4338 0 _1125_.vdd
rlabel metal2 4513 4173 4527 4187 0 _1125_.A
rlabel metal2 4533 4193 4547 4207 0 _1125_.B
rlabel metal2 4593 4173 4607 4187 0 _1125_.C
rlabel metal2 4573 4193 4587 4207 0 _1125_.D
rlabel metal2 4553 4173 4567 4187 0 _1125_.Y
rlabel nsubstratencontact 4756 4328 4756 4328 0 FILL71250x61350.vdd
rlabel metal1 4744 4082 4776 4098 0 FILL71250x61350.gnd
rlabel nsubstratencontact 4736 4328 4736 4328 0 FILL70950x61350.vdd
rlabel metal1 4724 4082 4756 4098 0 FILL70950x61350.gnd
rlabel nsubstratencontact 4716 4328 4716 4328 0 FILL70650x61350.vdd
rlabel metal1 4704 4082 4736 4098 0 FILL70650x61350.gnd
rlabel metal1 4624 4082 4716 4098 0 _1126_.gnd
rlabel metal1 4624 4322 4716 4338 0 _1126_.vdd
rlabel metal2 4653 4173 4667 4187 0 _1126_.B
rlabel metal2 4693 4173 4707 4187 0 _1126_.A
rlabel metal2 4673 4153 4687 4167 0 _1126_.Y
rlabel metal1 4 4562 96 4578 0 _1609_.gnd
rlabel metal1 4 4322 96 4338 0 _1609_.vdd
rlabel metal2 73 4473 87 4487 0 _1609_.A
rlabel metal2 33 4473 47 4487 0 _1609_.Y
rlabel metal1 264 4562 356 4578 0 _1607_.gnd
rlabel metal1 264 4322 356 4338 0 _1607_.vdd
rlabel metal2 273 4473 287 4487 0 _1607_.A
rlabel metal2 313 4473 327 4487 0 _1607_.Y
rlabel metal1 164 4562 276 4578 0 _1373_.gnd
rlabel metal1 164 4322 276 4338 0 _1373_.vdd
rlabel metal2 253 4473 267 4487 0 _1373_.A
rlabel metal2 233 4453 247 4467 0 _1373_.B
rlabel metal2 193 4453 207 4467 0 _1373_.C
rlabel metal2 213 4473 227 4487 0 _1373_.Y
rlabel metal1 84 4562 176 4578 0 _1372_.gnd
rlabel metal1 84 4322 176 4338 0 _1372_.vdd
rlabel metal2 153 4433 167 4447 0 _1372_.A
rlabel metal2 113 4433 127 4447 0 _1372_.B
rlabel metal2 133 4453 147 4467 0 _1372_.Y
rlabel metal1 504 4562 596 4578 0 _1606_.gnd
rlabel metal1 504 4322 596 4338 0 _1606_.vdd
rlabel metal2 513 4473 527 4487 0 _1606_.A
rlabel metal2 553 4473 567 4487 0 _1606_.Y
rlabel metal1 424 4562 516 4578 0 _1366_.gnd
rlabel metal1 424 4322 516 4338 0 _1366_.vdd
rlabel metal2 453 4473 467 4487 0 _1366_.B
rlabel metal2 493 4473 507 4487 0 _1366_.A
rlabel metal2 473 4493 487 4507 0 _1366_.Y
rlabel metal1 344 4562 436 4578 0 _1365_.gnd
rlabel metal1 344 4322 436 4338 0 _1365_.vdd
rlabel metal2 373 4473 387 4487 0 _1365_.B
rlabel metal2 413 4473 427 4487 0 _1365_.A
rlabel metal2 393 4493 407 4507 0 _1365_.Y
rlabel metal1 784 4562 1036 4578 0 _1535_.gnd
rlabel metal1 784 4322 1036 4338 0 _1535_.vdd
rlabel metal2 933 4473 947 4487 0 _1535_.D
rlabel metal2 893 4473 907 4487 0 _1535_.CLK
rlabel metal2 813 4473 827 4487 0 _1535_.Q
rlabel metal1 644 4562 736 4578 0 _1364_.gnd
rlabel metal1 644 4322 736 4338 0 _1364_.vdd
rlabel metal2 693 4473 707 4487 0 _1364_.B
rlabel metal2 653 4473 667 4487 0 _1364_.A
rlabel metal2 673 4493 687 4507 0 _1364_.Y
rlabel metal1 724 4562 796 4578 0 _953_.gnd
rlabel metal1 724 4322 796 4338 0 _953_.vdd
rlabel metal2 733 4493 747 4507 0 _953_.A
rlabel metal2 753 4453 767 4467 0 _953_.Y
rlabel metal1 584 4562 656 4578 0 _818_.gnd
rlabel metal1 584 4322 656 4338 0 _818_.vdd
rlabel metal2 633 4493 647 4507 0 _818_.A
rlabel metal2 613 4453 627 4467 0 _818_.Y
rlabel metal1 1024 4562 1136 4578 0 _820_.gnd
rlabel metal1 1024 4322 1136 4338 0 _820_.vdd
rlabel metal2 1033 4473 1047 4487 0 _820_.A
rlabel metal2 1053 4453 1067 4467 0 _820_.B
rlabel metal2 1093 4453 1107 4467 0 _820_.C
rlabel metal2 1073 4473 1087 4487 0 _820_.Y
rlabel metal1 1124 4562 1376 4578 0 _1551_.gnd
rlabel metal1 1124 4322 1376 4338 0 _1551_.vdd
rlabel metal2 1273 4473 1287 4487 0 _1551_.D
rlabel metal2 1233 4473 1247 4487 0 _1551_.CLK
rlabel metal2 1153 4473 1167 4487 0 _1551_.Q
rlabel metal1 1464 4562 1716 4578 0 _1536_.gnd
rlabel metal1 1464 4322 1716 4338 0 _1536_.vdd
rlabel metal2 1553 4473 1567 4487 0 _1536_.D
rlabel metal2 1593 4473 1607 4487 0 _1536_.CLK
rlabel metal2 1673 4473 1687 4487 0 _1536_.Q
rlabel metal1 1364 4562 1476 4578 0 _1005_.gnd
rlabel metal1 1364 4322 1476 4338 0 _1005_.vdd
rlabel metal2 1373 4473 1387 4487 0 _1005_.A
rlabel metal2 1393 4453 1407 4467 0 _1005_.B
rlabel metal2 1433 4453 1447 4467 0 _1005_.C
rlabel metal2 1413 4473 1427 4487 0 _1005_.Y
rlabel metal1 1784 4562 2036 4578 0 _1552_.gnd
rlabel metal1 1784 4322 2036 4338 0 _1552_.vdd
rlabel metal2 1933 4473 1947 4487 0 _1552_.D
rlabel metal2 1893 4473 1907 4487 0 _1552_.CLK
rlabel metal2 1813 4473 1827 4487 0 _1552_.Q
rlabel metal1 1704 4562 1796 4578 0 _819_.gnd
rlabel metal1 1704 4322 1796 4338 0 _819_.vdd
rlabel metal2 1713 4433 1727 4447 0 _819_.A
rlabel metal2 1753 4433 1767 4447 0 _819_.B
rlabel metal2 1733 4453 1747 4467 0 _819_.Y
rlabel metal1 2024 4562 2156 4578 0 _1069_.gnd
rlabel metal1 2024 4322 2156 4338 0 _1069_.vdd
rlabel metal2 2033 4473 2047 4487 0 _1069_.A
rlabel metal2 2053 4453 2067 4467 0 _1069_.B
rlabel metal2 2113 4473 2127 4487 0 _1069_.C
rlabel metal2 2073 4473 2087 4487 0 _1069_.Y
rlabel metal2 2093 4453 2107 4467 0 _1069_.D
rlabel metal1 2244 4562 2356 4578 0 _1068_.gnd
rlabel metal1 2244 4322 2356 4338 0 _1068_.vdd
rlabel metal2 2333 4473 2347 4487 0 _1068_.A
rlabel metal2 2313 4453 2327 4467 0 _1068_.B
rlabel metal2 2273 4453 2287 4467 0 _1068_.C
rlabel metal2 2293 4473 2307 4487 0 _1068_.Y
rlabel metal1 2404 4562 2496 4578 0 _1066_.gnd
rlabel metal1 2404 4322 2496 4338 0 _1066_.vdd
rlabel metal2 2453 4473 2467 4487 0 _1066_.B
rlabel metal2 2413 4473 2427 4487 0 _1066_.A
rlabel metal2 2433 4493 2447 4507 0 _1066_.Y
rlabel metal1 2344 4562 2416 4578 0 _1003_.gnd
rlabel metal1 2344 4322 2416 4338 0 _1003_.vdd
rlabel metal2 2393 4493 2407 4507 0 _1003_.A
rlabel metal2 2373 4453 2387 4467 0 _1003_.Y
rlabel metal1 2144 4562 2256 4578 0 _1004_.gnd
rlabel metal1 2144 4322 2256 4338 0 _1004_.vdd
rlabel metal2 2233 4453 2247 4467 0 _1004_.A
rlabel metal2 2213 4433 2227 4447 0 _1004_.B
rlabel metal2 2193 4453 2207 4467 0 _1004_.C
rlabel metal2 2173 4433 2187 4447 0 _1004_.Y
rlabel metal1 2644 4562 2736 4578 0 _1601_.gnd
rlabel metal1 2644 4322 2736 4338 0 _1601_.vdd
rlabel metal2 2653 4473 2667 4487 0 _1601_.A
rlabel metal2 2693 4473 2707 4487 0 _1601_.Y
rlabel metal1 2544 4562 2656 4578 0 _1128_.gnd
rlabel metal1 2544 4322 2656 4338 0 _1128_.vdd
rlabel metal2 2553 4473 2567 4487 0 _1128_.A
rlabel metal2 2573 4453 2587 4467 0 _1128_.B
rlabel metal2 2613 4453 2627 4467 0 _1128_.C
rlabel metal2 2593 4473 2607 4487 0 _1128_.Y
rlabel metal1 2484 4562 2556 4578 0 _1067_.gnd
rlabel metal1 2484 4322 2556 4338 0 _1067_.vdd
rlabel metal2 2533 4493 2547 4507 0 _1067_.A
rlabel metal2 2513 4453 2527 4467 0 _1067_.Y
rlabel metal1 2724 4562 2816 4578 0 _1605_.gnd
rlabel metal1 2724 4322 2816 4338 0 _1605_.vdd
rlabel metal2 2733 4473 2747 4487 0 _1605_.A
rlabel metal2 2773 4473 2787 4487 0 _1605_.Y
rlabel metal1 2804 4562 2896 4578 0 _1604_.gnd
rlabel metal1 2804 4322 2896 4338 0 _1604_.vdd
rlabel metal2 2873 4473 2887 4487 0 _1604_.A
rlabel metal2 2833 4473 2847 4487 0 _1604_.Y
rlabel metal1 2884 4562 2996 4578 0 _1071_.gnd
rlabel metal1 2884 4322 2996 4338 0 _1071_.vdd
rlabel metal2 2973 4453 2987 4467 0 _1071_.A
rlabel metal2 2953 4433 2967 4447 0 _1071_.B
rlabel metal2 2933 4453 2947 4467 0 _1071_.C
rlabel metal2 2913 4433 2927 4447 0 _1071_.Y
rlabel metal1 3084 4562 3176 4578 0 _1602_.gnd
rlabel metal1 3084 4322 3176 4338 0 _1602_.vdd
rlabel metal2 3153 4473 3167 4487 0 _1602_.A
rlabel metal2 3113 4473 3127 4487 0 _1602_.Y
rlabel metal1 3164 4562 3276 4578 0 _998_.gnd
rlabel metal1 3164 4322 3276 4338 0 _998_.vdd
rlabel metal2 3253 4453 3267 4467 0 _998_.A
rlabel metal2 3233 4433 3247 4447 0 _998_.B
rlabel metal2 3213 4453 3227 4467 0 _998_.C
rlabel metal2 3193 4433 3207 4447 0 _998_.Y
rlabel metal1 2984 4562 3096 4578 0 _1065_.gnd
rlabel metal1 2984 4322 3096 4338 0 _1065_.vdd
rlabel metal2 3073 4473 3087 4487 0 _1065_.A
rlabel metal2 3013 4473 3027 4487 0 _1065_.Y
rlabel metal2 3033 4433 3047 4447 0 _1065_.B
rlabel metal1 3264 4562 3356 4578 0 _997_.gnd
rlabel metal1 3264 4322 3356 4338 0 _997_.vdd
rlabel metal2 3273 4433 3287 4447 0 _997_.A
rlabel metal2 3313 4433 3327 4447 0 _997_.B
rlabel metal2 3293 4453 3307 4467 0 _997_.Y
rlabel metal1 3344 4562 3456 4578 0 _1061_.gnd
rlabel metal1 3344 4322 3456 4338 0 _1061_.vdd
rlabel metal2 3353 4453 3367 4467 0 _1061_.A
rlabel metal2 3373 4493 3387 4507 0 _1061_.B
rlabel metal2 3393 4453 3407 4467 0 _1061_.C
rlabel metal2 3413 4473 3427 4487 0 _1061_.Y
rlabel metal1 3444 4562 3516 4578 0 _1060_.gnd
rlabel metal1 3444 4322 3516 4338 0 _1060_.vdd
rlabel metal2 3453 4493 3467 4507 0 _1060_.A
rlabel metal2 3473 4453 3487 4467 0 _1060_.Y
rlabel metal1 3504 4562 3596 4578 0 _993_.gnd
rlabel metal1 3504 4322 3596 4338 0 _993_.vdd
rlabel metal2 3513 4433 3527 4447 0 _993_.A
rlabel metal2 3553 4433 3567 4447 0 _993_.B
rlabel metal2 3533 4453 3547 4467 0 _993_.Y
rlabel metal1 3684 4562 3796 4578 0 _1007_.gnd
rlabel metal1 3684 4322 3796 4338 0 _1007_.vdd
rlabel metal2 3693 4453 3707 4467 0 _1007_.A
rlabel metal2 3713 4493 3727 4507 0 _1007_.B
rlabel metal2 3733 4453 3747 4467 0 _1007_.C
rlabel metal2 3753 4473 3767 4487 0 _1007_.Y
rlabel metal1 3584 4562 3696 4578 0 _996_.gnd
rlabel metal1 3584 4322 3696 4338 0 _996_.vdd
rlabel metal2 3593 4453 3607 4467 0 _996_.A
rlabel metal2 3613 4433 3627 4447 0 _996_.B
rlabel metal2 3633 4453 3647 4467 0 _996_.C
rlabel metal2 3653 4433 3667 4447 0 _996_.Y
rlabel metal1 3884 4562 3996 4578 0 _1064_.gnd
rlabel metal1 3884 4322 3996 4338 0 _1064_.vdd
rlabel metal2 3973 4473 3987 4487 0 _1064_.A
rlabel metal2 3953 4453 3967 4467 0 _1064_.B
rlabel metal2 3913 4453 3927 4467 0 _1064_.C
rlabel metal2 3933 4473 3947 4487 0 _1064_.Y
rlabel metal1 3784 4562 3896 4578 0 _1008_.gnd
rlabel metal1 3784 4322 3896 4338 0 _1008_.vdd
rlabel metal2 3793 4473 3807 4487 0 _1008_.A
rlabel metal2 3813 4453 3827 4467 0 _1008_.B
rlabel metal2 3853 4453 3867 4467 0 _1008_.C
rlabel metal2 3833 4473 3847 4487 0 _1008_.Y
rlabel metal1 3984 4562 4096 4578 0 _1059_.gnd
rlabel metal1 3984 4322 4096 4338 0 _1059_.vdd
rlabel metal2 4073 4453 4087 4467 0 _1059_.A
rlabel metal2 4053 4433 4067 4447 0 _1059_.B
rlabel metal2 4033 4453 4047 4467 0 _1059_.C
rlabel metal2 4013 4433 4027 4447 0 _1059_.Y
rlabel metal1 4184 4562 4296 4578 0 _1063_.gnd
rlabel metal1 4184 4322 4296 4338 0 _1063_.vdd
rlabel metal2 4193 4453 4207 4467 0 _1063_.A
rlabel metal2 4213 4493 4227 4507 0 _1063_.B
rlabel metal2 4233 4453 4247 4467 0 _1063_.C
rlabel metal2 4253 4473 4267 4487 0 _1063_.Y
rlabel metal1 4084 4562 4196 4578 0 _1055_.gnd
rlabel metal1 4084 4322 4196 4338 0 _1055_.vdd
rlabel metal2 4173 4453 4187 4467 0 _1055_.A
rlabel metal2 4153 4433 4167 4447 0 _1055_.B
rlabel metal2 4133 4453 4147 4467 0 _1055_.C
rlabel metal2 4113 4433 4127 4447 0 _1055_.Y
rlabel metal1 4284 4562 4376 4578 0 _1024_.gnd
rlabel metal1 4284 4322 4376 4338 0 _1024_.vdd
rlabel metal2 4293 4433 4307 4447 0 _1024_.A
rlabel metal2 4333 4433 4347 4447 0 _1024_.B
rlabel metal2 4313 4453 4327 4467 0 _1024_.Y
rlabel metal1 4364 4562 4476 4578 0 _1062_.gnd
rlabel metal1 4364 4322 4476 4338 0 _1062_.vdd
rlabel metal2 4453 4453 4467 4467 0 _1062_.A
rlabel metal2 4433 4493 4447 4507 0 _1062_.B
rlabel metal2 4413 4453 4427 4467 0 _1062_.C
rlabel metal2 4393 4473 4407 4487 0 _1062_.Y
rlabel metal1 4464 4562 4536 4578 0 _1011_.gnd
rlabel metal1 4464 4322 4536 4338 0 _1011_.vdd
rlabel metal2 4513 4493 4527 4507 0 _1011_.A
rlabel metal2 4493 4453 4507 4467 0 _1011_.Y
rlabel metal1 4524 4562 4636 4578 0 _1058_.gnd
rlabel metal1 4524 4322 4636 4338 0 _1058_.vdd
rlabel metal2 4533 4453 4547 4467 0 _1058_.A
rlabel metal2 4553 4433 4567 4447 0 _1058_.B
rlabel metal2 4573 4453 4587 4467 0 _1058_.C
rlabel metal2 4593 4433 4607 4447 0 _1058_.Y
rlabel nsubstratencontact 4764 4332 4764 4332 0 FILL71250x64950.vdd
rlabel metal1 4744 4562 4776 4578 0 FILL71250x64950.gnd
rlabel nsubstratencontact 4744 4332 4744 4332 0 FILL70950x64950.vdd
rlabel metal1 4724 4562 4756 4578 0 FILL70950x64950.gnd
rlabel metal1 4624 4562 4736 4578 0 _1111_.gnd
rlabel metal1 4624 4322 4736 4338 0 _1111_.vdd
rlabel metal2 4633 4453 4647 4467 0 _1111_.A
rlabel metal2 4653 4433 4667 4447 0 _1111_.B
rlabel metal2 4673 4453 4687 4467 0 _1111_.C
rlabel metal2 4693 4433 4707 4447 0 _1111_.Y
<< end >>
