magic
tech scmos
magscale 1 2
timestamp 1727155535
<< error_s >>
rect 4 6244 6136 6256
rect 4 5984 6136 5996
rect 4 5724 6136 5736
rect 4 5464 6136 5476
rect 4 5204 6136 5216
rect 4 4944 6136 4956
rect 4 4684 6136 4696
rect 4 4424 6136 4436
rect 4 4164 6136 4176
rect 4 3904 6136 3916
rect 4 3644 6136 3656
rect 4 3384 6136 3396
rect 4 3124 6136 3136
rect 4 2864 6136 2876
rect 4 2604 6136 2616
rect 4 2344 6136 2356
rect 4 2084 6136 2096
rect 4 1824 6136 1836
rect 4 1564 6136 1576
rect 4 1304 6136 1316
rect 4 1044 6136 1056
rect 4 784 6136 796
rect 4 524 6136 536
rect 4 264 6136 276
rect 4 4 6136 16
<< nwell >>
rect 2200 3751 2215 3756
<< metal1 >>
rect -63 6242 30 6258
rect -63 5738 -3 6242
rect 2287 6137 2333 6143
rect 2547 6137 2653 6143
rect 5607 6137 5693 6143
rect 3913 6123 3927 6133
rect 3897 6120 3927 6123
rect 3897 6117 3923 6120
rect 3897 6087 3903 6117
rect 4027 6123 4040 6127
rect 5900 6123 5913 6127
rect 4027 6113 4043 6123
rect 4037 6087 4043 6113
rect 5897 6113 5913 6123
rect 4587 6103 4600 6107
rect 4587 6097 4614 6103
rect 4587 6093 4600 6097
rect 5897 6087 5903 6113
rect 3897 6077 3913 6087
rect 3900 6073 3913 6077
rect 4037 6077 4053 6087
rect 4040 6073 4053 6077
rect 4720 6083 4733 6087
rect 4717 6077 4733 6083
rect 4720 6073 4733 6077
rect 5897 6077 5913 6087
rect 5900 6073 5913 6077
rect 5187 6057 5253 6063
rect 6143 5998 6203 6258
rect 6110 5982 6203 5998
rect 2861 5937 2893 5943
rect 2147 5917 2193 5923
rect 2807 5917 2853 5923
rect 4287 5917 4353 5923
rect 207 5903 220 5907
rect 3700 5903 3713 5907
rect 207 5893 223 5903
rect 217 5867 223 5893
rect 3697 5893 3713 5903
rect 5307 5903 5320 5907
rect 5620 5903 5633 5907
rect 5307 5893 5323 5903
rect 3697 5867 3703 5893
rect 5317 5867 5323 5893
rect 207 5857 223 5867
rect 207 5853 220 5857
rect 2987 5857 3013 5863
rect 3680 5866 3703 5867
rect 3687 5857 3703 5866
rect 3687 5853 3700 5857
rect 5307 5857 5323 5867
rect 5617 5893 5633 5903
rect 5617 5867 5623 5893
rect 5617 5857 5633 5867
rect 5307 5853 5320 5857
rect 5620 5853 5633 5857
rect 2587 5837 2653 5843
rect 4187 5837 4233 5843
rect 5447 5837 5513 5843
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 387 5617 433 5623
rect 2267 5617 2293 5623
rect 3007 5617 3053 5623
rect 4887 5617 4913 5623
rect 2213 5603 2227 5613
rect 527 5597 583 5603
rect 2213 5600 2243 5603
rect 2217 5597 2243 5600
rect 527 5557 553 5563
rect 577 5547 583 5597
rect 2237 5563 2243 5597
rect 4387 5597 4443 5603
rect 4437 5567 4443 5597
rect 4827 5597 4883 5603
rect 4877 5567 4883 5597
rect 5480 5583 5493 5587
rect 5327 5577 5374 5583
rect 5477 5577 5493 5583
rect 5480 5573 5493 5577
rect 2237 5557 2273 5563
rect 4437 5557 4453 5567
rect 4440 5553 4453 5557
rect 4877 5557 4893 5567
rect 4880 5553 4893 5557
rect 560 5546 583 5547
rect 567 5537 583 5546
rect 567 5533 580 5537
rect 1107 5537 1153 5543
rect 3461 5537 3493 5543
rect 5147 5537 5193 5543
rect 5207 5537 5233 5543
rect 1647 5517 1713 5523
rect 1927 5497 1973 5503
rect 6143 5478 6203 5982
rect 6110 5462 6203 5478
rect 1077 5343 1083 5393
rect 2600 5383 2613 5387
rect 2597 5373 2613 5383
rect 2707 5383 2720 5387
rect 2707 5373 2723 5383
rect 2847 5383 2860 5387
rect 2960 5383 2973 5387
rect 2847 5373 2863 5383
rect 2597 5347 2603 5373
rect 2717 5347 2723 5373
rect 2857 5347 2863 5373
rect 1077 5337 1133 5343
rect 1517 5337 1553 5343
rect 2597 5337 2613 5347
rect 2600 5333 2613 5337
rect 2707 5337 2723 5347
rect 2707 5333 2720 5337
rect 2847 5337 2863 5347
rect 2957 5373 2973 5383
rect 3187 5383 3200 5387
rect 3380 5383 3393 5387
rect 3187 5373 3203 5383
rect 2957 5347 2963 5373
rect 3197 5347 3203 5373
rect 2957 5337 2973 5347
rect 2847 5333 2860 5337
rect 2960 5333 2973 5337
rect 3187 5337 3203 5347
rect 3377 5373 3393 5383
rect 3647 5383 3660 5387
rect 3647 5373 3663 5383
rect 4367 5383 4380 5387
rect 4367 5373 4383 5383
rect 3377 5347 3383 5373
rect 3657 5347 3663 5373
rect 4377 5347 4383 5373
rect 5597 5377 5633 5383
rect 5597 5347 5603 5377
rect 3377 5337 3393 5347
rect 3187 5333 3200 5337
rect 3380 5333 3393 5337
rect 3647 5337 3663 5347
rect 3647 5333 3660 5337
rect 4247 5337 4273 5343
rect 4367 5337 4383 5347
rect 4367 5333 4380 5337
rect 5587 5337 5603 5347
rect 5587 5333 5600 5337
rect 1127 5317 1153 5323
rect 1987 5317 2053 5323
rect 2387 5317 2513 5323
rect 3207 5317 3273 5323
rect 3327 5317 3373 5323
rect 4707 5317 4773 5323
rect 2567 5297 2633 5303
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 4167 5177 4193 5183
rect 3997 5097 4053 5103
rect 1680 5083 1693 5087
rect 1677 5073 1693 5083
rect 2447 5083 2460 5087
rect 2447 5073 2463 5083
rect 2607 5077 2643 5083
rect 1677 5047 1683 5073
rect 2457 5047 2463 5073
rect 2637 5047 2643 5077
rect 3207 5077 3233 5083
rect 3527 5077 3553 5083
rect 3667 5083 3680 5087
rect 3667 5073 3683 5083
rect 3677 5047 3683 5073
rect 3997 5047 4003 5097
rect 5057 5097 5113 5103
rect 4180 5083 4193 5087
rect 1167 5037 1193 5043
rect 1677 5037 1693 5047
rect 1680 5033 1693 5037
rect 2457 5037 2473 5047
rect 2460 5033 2473 5037
rect 2637 5037 2653 5047
rect 2640 5033 2653 5037
rect 2747 5037 2773 5043
rect 3667 5037 3683 5047
rect 3667 5033 3680 5037
rect 3987 5037 4003 5047
rect 4177 5073 4193 5083
rect 4640 5083 4653 5087
rect 4637 5073 4653 5083
rect 4767 5083 4780 5087
rect 4767 5073 4783 5083
rect 4177 5047 4183 5073
rect 4637 5047 4643 5073
rect 4777 5047 4783 5073
rect 5057 5047 5063 5097
rect 5207 5083 5220 5087
rect 5380 5083 5393 5087
rect 5207 5073 5223 5083
rect 4177 5037 4193 5047
rect 3987 5033 4000 5037
rect 4180 5033 4193 5037
rect 4637 5037 4653 5047
rect 4640 5033 4653 5037
rect 4777 5037 4793 5047
rect 4780 5033 4793 5037
rect 5047 5037 5063 5047
rect 5047 5033 5060 5037
rect 1407 5017 1553 5023
rect 3227 5017 3253 5023
rect 5217 5023 5223 5073
rect 5377 5073 5393 5083
rect 5377 5043 5383 5073
rect 5347 5037 5383 5043
rect 5217 5017 5253 5023
rect 6143 4958 6203 5462
rect 6110 4942 6203 4958
rect 5727 4917 5753 4923
rect 2107 4877 2133 4883
rect 2627 4877 2673 4883
rect 4077 4877 4153 4883
rect 2747 4863 2760 4867
rect 2800 4863 2813 4867
rect 2747 4853 2763 4863
rect 2757 4827 2763 4853
rect 2577 4817 2613 4823
rect 2747 4817 2763 4827
rect 2797 4853 2813 4863
rect 3360 4863 3373 4867
rect 3067 4857 3103 4863
rect 2747 4813 2760 4817
rect 927 4797 1013 4803
rect 2287 4797 2333 4803
rect 2797 4806 2803 4853
rect 3097 4823 3103 4857
rect 3357 4853 3373 4863
rect 3607 4863 3620 4867
rect 3607 4853 3623 4863
rect 3097 4817 3123 4823
rect 3117 4807 3123 4817
rect 3117 4797 3133 4807
rect 3120 4793 3133 4797
rect 3357 4803 3363 4853
rect 3617 4827 3623 4853
rect 3607 4817 3623 4827
rect 4077 4827 4083 4877
rect 4647 4877 4693 4883
rect 5277 4877 5333 4883
rect 4347 4863 4360 4867
rect 4520 4863 4533 4867
rect 4347 4853 4363 4863
rect 4357 4827 4363 4853
rect 4517 4853 4533 4863
rect 4660 4863 4673 4867
rect 4657 4853 4673 4863
rect 4827 4863 4840 4867
rect 4827 4853 4843 4863
rect 5140 4863 5153 4867
rect 4927 4857 4963 4863
rect 4517 4827 4523 4853
rect 4657 4827 4663 4853
rect 4837 4827 4843 4853
rect 4077 4817 4093 4827
rect 3607 4813 3620 4817
rect 4080 4813 4093 4817
rect 4347 4817 4363 4827
rect 4347 4813 4360 4817
rect 4507 4817 4523 4827
rect 4507 4813 4520 4817
rect 4647 4817 4663 4827
rect 4647 4813 4660 4817
rect 4827 4817 4843 4827
rect 4957 4827 4963 4857
rect 5137 4853 5153 4863
rect 5137 4827 5143 4853
rect 5277 4827 5283 4877
rect 5440 4863 5453 4867
rect 4957 4817 4973 4827
rect 4827 4813 4840 4817
rect 4960 4813 4973 4817
rect 5137 4817 5153 4827
rect 5140 4813 5153 4817
rect 5267 4817 5283 4827
rect 5437 4853 5453 4863
rect 5867 4857 5943 4863
rect 5437 4827 5443 4853
rect 6060 4843 6073 4847
rect 6046 4837 6073 4843
rect 6060 4833 6073 4837
rect 5437 4817 5453 4827
rect 5267 4813 5280 4817
rect 5440 4813 5453 4817
rect 5867 4817 5893 4823
rect 3327 4797 3363 4803
rect 5067 4797 5113 4803
rect 5687 4797 5753 4803
rect 4487 4757 4513 4763
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 5187 4657 5253 4663
rect 4667 4617 4733 4623
rect 407 4577 473 4583
rect 2900 4583 2913 4587
rect 2897 4573 2913 4583
rect 5040 4583 5053 4587
rect 5037 4573 5053 4583
rect 1307 4563 1320 4567
rect 1307 4553 1323 4563
rect 2447 4563 2460 4567
rect 2780 4563 2793 4567
rect 2447 4553 2463 4563
rect 946 4537 993 4543
rect 613 4523 627 4533
rect 1317 4527 1323 4553
rect 2457 4543 2463 4553
rect 2777 4553 2793 4563
rect 2897 4563 2903 4573
rect 2877 4557 2903 4563
rect 2600 4543 2613 4547
rect 2457 4537 2494 4543
rect 2597 4537 2613 4543
rect 2600 4533 2613 4537
rect 2777 4527 2783 4553
rect 613 4520 653 4523
rect 617 4517 653 4520
rect 827 4523 840 4527
rect 827 4517 843 4523
rect 1317 4517 1333 4527
rect 827 4513 840 4517
rect 1320 4513 1333 4517
rect 1427 4517 1453 4523
rect 2767 4517 2783 4527
rect 2877 4527 2883 4557
rect 4687 4563 4700 4567
rect 4687 4553 4703 4563
rect 3347 4543 3360 4547
rect 3480 4543 3493 4547
rect 3347 4537 3363 4543
rect 3466 4537 3493 4543
rect 3347 4533 3360 4537
rect 3480 4533 3493 4537
rect 2877 4517 2893 4527
rect 2767 4513 2780 4517
rect 2880 4513 2893 4517
rect 3517 4507 3523 4553
rect 4697 4527 4703 4553
rect 4747 4543 4760 4547
rect 4747 4537 4763 4543
rect 4866 4537 4903 4543
rect 4747 4533 4760 4537
rect 4687 4517 4703 4527
rect 4897 4527 4903 4537
rect 5037 4527 5043 4573
rect 5060 4563 5073 4567
rect 4897 4517 4913 4527
rect 4687 4513 4700 4517
rect 4900 4513 4913 4517
rect 5027 4517 5043 4527
rect 5057 4553 5073 4563
rect 5487 4557 5523 4563
rect 5057 4527 5063 4553
rect 5057 4517 5073 4527
rect 5027 4513 5040 4517
rect 5060 4513 5073 4517
rect 5517 4523 5523 4557
rect 5647 4557 5703 4563
rect 5697 4543 5703 4557
rect 5697 4537 5734 4543
rect 5997 4527 6003 4573
rect 5517 4517 5543 4523
rect 5837 4517 5893 4523
rect 1707 4497 1773 4503
rect 2007 4497 2053 4503
rect 3507 4497 3523 4507
rect 5537 4507 5543 4517
rect 5987 4517 6003 4527
rect 5987 4513 6000 4517
rect 5537 4497 5553 4507
rect 3507 4493 3520 4497
rect 5540 4493 5553 4497
rect 6143 4438 6203 4942
rect 6110 4422 6203 4438
rect 1247 4397 1273 4403
rect 447 4343 460 4347
rect 447 4333 463 4343
rect 2467 4343 2480 4347
rect 2467 4333 2483 4343
rect 2637 4337 2673 4343
rect 4397 4337 4433 4343
rect 457 4303 463 4333
rect 1560 4323 1573 4327
rect 1557 4317 1573 4323
rect 1560 4313 1573 4317
rect 457 4297 483 4303
rect 917 4297 953 4303
rect 477 4287 483 4297
rect 1440 4306 1460 4307
rect 1447 4303 1460 4306
rect 2477 4303 2483 4333
rect 2507 4323 2520 4327
rect 2507 4317 2534 4323
rect 2507 4313 2520 4317
rect 4397 4303 4403 4337
rect 4597 4343 4603 4373
rect 4687 4357 4773 4363
rect 5227 4357 5293 4363
rect 4567 4337 4603 4343
rect 4727 4337 4763 4343
rect 1447 4297 1463 4303
rect 2477 4297 2503 4303
rect 4357 4297 4403 4303
rect 4757 4307 4763 4337
rect 4977 4337 5013 4343
rect 4977 4307 4983 4337
rect 5127 4337 5163 4343
rect 4757 4297 4773 4307
rect 1447 4293 1460 4297
rect 477 4277 493 4287
rect 480 4273 493 4277
rect 1437 4283 1443 4292
rect 2497 4287 2503 4297
rect 4760 4293 4773 4297
rect 4967 4297 4983 4307
rect 5157 4307 5163 4337
rect 5367 4343 5380 4347
rect 5367 4333 5383 4343
rect 5527 4337 5553 4343
rect 5700 4343 5713 4347
rect 5697 4333 5713 4343
rect 5827 4343 5840 4347
rect 5827 4333 5843 4343
rect 5377 4307 5383 4333
rect 5157 4297 5173 4307
rect 4967 4293 4980 4297
rect 5160 4293 5173 4297
rect 5367 4297 5383 4307
rect 5697 4303 5703 4333
rect 5837 4303 5843 4333
rect 5697 4297 5723 4303
rect 5367 4293 5380 4297
rect 5717 4287 5723 4297
rect 5817 4297 5843 4303
rect 5817 4287 5823 4297
rect 1367 4277 1443 4283
rect 2027 4277 2113 4283
rect 2497 4277 2513 4287
rect 2500 4273 2513 4277
rect 4527 4277 4593 4283
rect 4667 4277 4753 4283
rect 5717 4277 5733 4287
rect 5720 4273 5733 4277
rect 5807 4277 5823 4287
rect 5807 4273 5820 4277
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 2667 4093 2673 4107
rect 207 4057 273 4063
rect 1787 4057 1853 4063
rect 1967 4057 2013 4063
rect 2367 4057 2393 4063
rect 4087 4057 4153 4063
rect 4327 4057 4413 4063
rect 5207 4057 5293 4063
rect 5707 4057 5753 4063
rect 5927 4057 5993 4063
rect 6017 4057 6073 4063
rect 880 4043 893 4047
rect 877 4037 893 4043
rect 880 4033 893 4037
rect 1580 4043 1593 4047
rect 1577 4033 1593 4043
rect 1667 4043 1680 4047
rect 1860 4043 1873 4047
rect 1667 4033 1683 4043
rect 1080 4023 1093 4027
rect 1066 4017 1093 4023
rect 1080 4013 1093 4017
rect 1577 4007 1583 4033
rect 467 3997 513 4003
rect 1577 3997 1593 4007
rect 1580 3993 1593 3997
rect 1677 4003 1683 4033
rect 1857 4033 1873 4043
rect 1980 4043 1993 4047
rect 1977 4033 1993 4043
rect 2097 4037 2133 4043
rect 1857 4007 1863 4033
rect 1677 3997 1733 4003
rect 1847 3997 1863 4007
rect 1847 3993 1860 3997
rect 1977 3987 1983 4033
rect 2097 4007 2103 4037
rect 2787 4043 2800 4047
rect 2940 4043 2953 4047
rect 2787 4033 2803 4043
rect 2797 4007 2803 4033
rect 2087 3997 2103 4007
rect 2087 3993 2100 3997
rect 2787 3997 2803 4007
rect 2937 4033 2953 4043
rect 4247 4043 4260 4047
rect 4247 4033 4263 4043
rect 4627 4043 4640 4047
rect 5100 4043 5113 4047
rect 4627 4033 4643 4043
rect 2937 4007 2943 4033
rect 2937 3997 2953 4007
rect 2787 3993 2800 3997
rect 2940 3993 2953 3997
rect 4257 3987 4263 4033
rect 1967 3977 1983 3987
rect 1967 3973 1980 3977
rect 2347 3977 2373 3983
rect 4507 3977 4553 3983
rect 4637 3966 4643 4033
rect 5097 4033 5113 4043
rect 5407 4043 5420 4047
rect 6017 4043 6023 4057
rect 5407 4033 5427 4043
rect 5097 4023 5103 4033
rect 5413 4027 5427 4033
rect 5997 4037 6023 4043
rect 5540 4023 5553 4027
rect 5046 4017 5103 4023
rect 5526 4017 5553 4023
rect 5097 4007 5103 4017
rect 5540 4013 5553 4017
rect 5997 4007 6003 4037
rect 4927 4003 4940 4007
rect 4927 3997 4943 4003
rect 5097 3997 5113 4007
rect 4927 3993 4940 3997
rect 5100 3993 5113 3997
rect 5347 3997 5423 4003
rect 5997 3997 6013 4007
rect 6000 3993 6013 3997
rect 6143 3918 6203 4422
rect 6110 3902 6203 3918
rect 2627 3877 2653 3883
rect 2647 3857 2713 3863
rect 5687 3857 5713 3863
rect 1507 3837 1543 3843
rect 760 3823 773 3827
rect 757 3813 773 3823
rect 867 3817 893 3823
rect 1220 3823 1233 3827
rect 1217 3813 1233 3823
rect 757 3787 763 3813
rect 1217 3787 1223 3813
rect 1357 3787 1363 3813
rect 1537 3787 1543 3837
rect 1920 3843 1933 3847
rect 1627 3837 1663 3843
rect 1657 3787 1663 3837
rect 1917 3833 1933 3843
rect 4967 3837 4993 3843
rect 5007 3837 5033 3843
rect 5807 3837 5873 3843
rect 1917 3787 1923 3833
rect 1940 3823 1953 3827
rect 757 3777 773 3787
rect 760 3773 773 3777
rect 1217 3777 1233 3787
rect 1220 3773 1233 3777
rect 1357 3777 1373 3787
rect 1360 3773 1373 3777
rect 1537 3777 1553 3787
rect 1540 3773 1553 3777
rect 1647 3777 1663 3787
rect 1647 3773 1660 3777
rect 1907 3777 1923 3787
rect 1937 3813 1953 3823
rect 2077 3817 2133 3823
rect 1937 3787 1943 3813
rect 2077 3787 2083 3817
rect 2800 3823 2813 3827
rect 2797 3813 2813 3823
rect 3987 3823 4000 3827
rect 3987 3813 4003 3823
rect 5687 3817 5723 3823
rect 1937 3777 1953 3787
rect 1907 3773 1920 3777
rect 1940 3773 1953 3777
rect 2067 3777 2083 3787
rect 2067 3773 2080 3777
rect 927 3757 973 3763
rect 1727 3757 1753 3763
rect 2087 3757 2133 3763
rect 2797 3766 2803 3813
rect 3997 3786 4003 3813
rect 5717 3787 5723 3817
rect 5827 3823 5840 3827
rect 5827 3813 5843 3823
rect 5947 3823 5960 3827
rect 5947 3813 5963 3823
rect 5837 3787 5843 3813
rect 5957 3787 5963 3813
rect 5717 3777 5733 3787
rect 5720 3773 5733 3777
rect 5837 3777 5853 3787
rect 5840 3773 5853 3777
rect 5947 3777 5963 3787
rect 5947 3773 5960 3777
rect 3067 3757 3133 3763
rect 5627 3757 5753 3763
rect 5807 3757 5873 3763
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 2687 3617 2713 3623
rect 1867 3577 1933 3583
rect 1567 3557 1653 3563
rect 67 3537 133 3543
rect 507 3537 593 3543
rect 1917 3537 1953 3543
rect 1620 3523 1633 3527
rect 1617 3513 1633 3523
rect 1917 3523 1923 3537
rect 2807 3537 2853 3543
rect 5487 3537 5533 3543
rect 5657 3537 5713 3543
rect 2040 3523 2053 3527
rect 1897 3520 1923 3523
rect 1893 3517 1923 3520
rect 1617 3487 1623 3513
rect 1893 3506 1907 3517
rect 2037 3513 2053 3523
rect 3787 3517 3813 3523
rect 4460 3523 4473 3527
rect 4457 3513 4473 3523
rect 5320 3523 5333 3527
rect 5317 3513 5333 3523
rect 2037 3487 2043 3513
rect 4457 3487 4463 3513
rect 1617 3477 1633 3487
rect 1620 3473 1633 3477
rect 2037 3477 2053 3487
rect 2040 3473 2053 3477
rect 4447 3477 4463 3487
rect 5317 3487 5323 3513
rect 5657 3487 5663 3537
rect 5977 3517 6013 3523
rect 5977 3487 5983 3517
rect 5317 3477 5333 3487
rect 4447 3473 4460 3477
rect 5320 3473 5333 3477
rect 5647 3477 5663 3487
rect 5647 3473 5660 3477
rect 5967 3477 5983 3487
rect 5967 3473 5980 3477
rect 2267 3457 2353 3463
rect 6143 3398 6203 3902
rect 6110 3382 6203 3398
rect 2507 3357 2553 3363
rect 3037 3327 3043 3353
rect 2360 3323 2373 3327
rect 2357 3313 2373 3323
rect 607 3303 620 3307
rect 640 3303 653 3307
rect 607 3293 623 3303
rect 617 3267 623 3293
rect 607 3257 623 3267
rect 637 3293 653 3303
rect 767 3303 780 3307
rect 1540 3303 1553 3307
rect 767 3293 783 3303
rect 607 3253 620 3257
rect 637 3247 643 3293
rect 777 3267 783 3293
rect 767 3257 783 3267
rect 1537 3293 1553 3303
rect 1627 3303 1640 3307
rect 1627 3293 1643 3303
rect 1947 3303 1960 3307
rect 1947 3293 1963 3303
rect 1537 3267 1543 3293
rect 1537 3257 1553 3267
rect 767 3253 780 3257
rect 1540 3253 1553 3257
rect 467 3237 513 3243
rect 1207 3237 1273 3243
rect 1637 3243 1643 3293
rect 1957 3267 1963 3293
rect 1947 3257 1963 3267
rect 2357 3263 2363 3313
rect 2380 3303 2393 3307
rect 2337 3257 2363 3263
rect 2377 3293 2393 3303
rect 2647 3303 2660 3307
rect 2647 3293 2663 3303
rect 2887 3303 2900 3307
rect 3360 3303 3373 3307
rect 2887 3293 2903 3303
rect 2377 3267 2383 3293
rect 2657 3267 2663 3293
rect 2897 3283 2903 3293
rect 3357 3293 3373 3303
rect 4067 3303 4080 3307
rect 4067 3293 4083 3303
rect 2897 3277 2923 3283
rect 2377 3257 2393 3267
rect 1947 3253 1960 3257
rect 2337 3247 2343 3257
rect 2380 3253 2393 3257
rect 2647 3257 2663 3267
rect 2917 3267 2923 3277
rect 3357 3267 3363 3293
rect 4077 3267 4083 3293
rect 4837 3297 4873 3303
rect 4837 3267 4843 3297
rect 2917 3257 2933 3267
rect 2647 3253 2660 3257
rect 2920 3253 2933 3257
rect 3357 3257 3373 3267
rect 3360 3253 3373 3257
rect 4067 3257 4083 3267
rect 4400 3263 4413 3267
rect 4067 3253 4080 3257
rect 4397 3253 4413 3263
rect 4827 3257 4843 3267
rect 4827 3253 4840 3257
rect 5157 3263 5163 3313
rect 5547 3303 5560 3307
rect 5547 3293 5563 3303
rect 5557 3267 5563 3293
rect 5967 3297 6003 3303
rect 5107 3257 5163 3263
rect 5547 3257 5563 3267
rect 5997 3263 6003 3297
rect 5997 3257 6023 3263
rect 5547 3253 5560 3257
rect 1637 3237 1693 3243
rect 2347 3237 2413 3243
rect 2507 3237 2553 3243
rect 3887 3237 3993 3243
rect 4397 3226 4403 3253
rect 4427 3237 4453 3243
rect 4947 3237 5013 3243
rect 6017 3243 6023 3257
rect 6017 3240 6043 3243
rect 6017 3237 6047 3240
rect 6033 3226 6047 3237
rect 5647 3197 5673 3203
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 2107 3097 2153 3103
rect 287 3017 393 3023
rect 1667 3017 1713 3023
rect 1947 3017 2033 3023
rect 2727 3017 2753 3023
rect 2827 3017 2893 3023
rect 1087 3003 1100 3007
rect 1087 2993 1103 3003
rect 1097 2967 1103 2993
rect 1357 2997 1413 3003
rect 1357 2967 1363 2997
rect 1827 2997 1853 3003
rect 1967 3003 1980 3007
rect 2160 3003 2173 3007
rect 1967 2993 1983 3003
rect 807 2957 853 2963
rect 1087 2957 1103 2967
rect 1087 2953 1100 2957
rect 1347 2957 1363 2967
rect 1347 2953 1360 2957
rect 1977 2947 1983 2993
rect 2157 2993 2173 3003
rect 2560 3003 2573 3007
rect 2557 2993 2573 3003
rect 3040 3003 3053 3007
rect 3037 2993 3053 3003
rect 3160 3003 3173 3007
rect 3157 2993 3173 3003
rect 3287 3003 3300 3007
rect 4000 3003 4013 3007
rect 3287 2993 3303 3003
rect 2157 2967 2163 2993
rect 2157 2957 2173 2967
rect 2160 2953 2173 2957
rect 2247 2937 2333 2943
rect 2557 2943 2563 2993
rect 2557 2937 2593 2943
rect 3037 2946 3043 2993
rect 3157 2967 3163 2993
rect 3297 2967 3303 2993
rect 3157 2957 3173 2967
rect 3160 2953 3173 2957
rect 3287 2957 3303 2967
rect 3997 2993 4013 3003
rect 4107 2997 4163 3003
rect 3997 2967 4003 2993
rect 4157 2967 4163 2997
rect 4287 3003 4300 3007
rect 5320 3003 5333 3007
rect 4287 2993 4303 3003
rect 4297 2967 4303 2993
rect 5317 2993 5333 3003
rect 5640 3003 5653 3007
rect 5637 2993 5653 3003
rect 5317 2967 5323 2993
rect 3997 2957 4013 2967
rect 3287 2953 3300 2957
rect 4000 2953 4013 2957
rect 4157 2957 4173 2967
rect 4160 2953 4173 2957
rect 4297 2957 4313 2967
rect 4300 2953 4313 2957
rect 4947 2957 4973 2963
rect 5317 2957 5333 2967
rect 5320 2953 5333 2957
rect 5637 2963 5643 2993
rect 5607 2957 5643 2963
rect 5167 2937 5213 2943
rect 5827 2917 5873 2923
rect 6143 2878 6203 3382
rect 6110 2862 6203 2878
rect 1647 2817 1713 2823
rect 5537 2807 5543 2833
rect 5673 2827 5687 2833
rect 5667 2820 5687 2827
rect 5667 2817 5683 2820
rect 5667 2813 5680 2817
rect 1487 2797 1513 2803
rect 1537 2797 1593 2803
rect 960 2783 973 2787
rect 957 2773 973 2783
rect 957 2747 963 2773
rect 957 2737 973 2747
rect 960 2733 973 2737
rect 427 2717 533 2723
rect 887 2717 953 2723
rect 1537 2726 1543 2797
rect 1927 2797 1993 2803
rect 2467 2797 2533 2803
rect 5367 2797 5433 2803
rect 5527 2797 5543 2807
rect 5527 2793 5540 2797
rect 1657 2777 1713 2783
rect 1657 2747 1663 2777
rect 2100 2783 2113 2787
rect 2097 2780 2113 2783
rect 2093 2773 2113 2780
rect 2240 2783 2253 2787
rect 2237 2773 2253 2783
rect 2477 2777 2513 2783
rect 2093 2766 2107 2773
rect 1647 2737 1663 2747
rect 2237 2747 2243 2773
rect 2477 2747 2483 2777
rect 2780 2783 2793 2787
rect 2777 2773 2793 2783
rect 3047 2783 3060 2787
rect 3280 2783 3293 2787
rect 3047 2773 3063 2783
rect 2593 2747 2607 2753
rect 2777 2747 2783 2773
rect 3057 2747 3063 2773
rect 3277 2773 3293 2783
rect 5100 2783 5113 2787
rect 5097 2773 5113 2783
rect 5227 2783 5240 2787
rect 5227 2773 5243 2783
rect 5347 2783 5360 2787
rect 5347 2773 5363 2783
rect 5377 2780 5413 2783
rect 3107 2763 3120 2767
rect 3240 2763 3253 2767
rect 3107 2757 3134 2763
rect 3237 2757 3253 2763
rect 3107 2753 3120 2757
rect 3240 2753 3253 2757
rect 2237 2737 2253 2747
rect 1647 2733 1660 2737
rect 2240 2733 2253 2737
rect 2467 2737 2483 2747
rect 2467 2733 2480 2737
rect 2587 2740 2607 2747
rect 2587 2737 2603 2740
rect 2587 2733 2600 2737
rect 2767 2737 2783 2747
rect 2767 2733 2780 2737
rect 3047 2737 3063 2747
rect 3277 2747 3283 2773
rect 5097 2767 5103 2773
rect 5080 2766 5103 2767
rect 5087 2757 5103 2766
rect 5087 2753 5100 2757
rect 5237 2747 5243 2773
rect 5357 2747 5363 2773
rect 5373 2777 5413 2780
rect 5373 2767 5387 2777
rect 5557 2747 5563 2813
rect 5767 2797 5813 2803
rect 5907 2797 5943 2803
rect 5660 2783 5673 2787
rect 3277 2737 3293 2747
rect 3047 2733 3060 2737
rect 3280 2733 3293 2737
rect 5107 2743 5120 2747
rect 5107 2740 5123 2743
rect 5107 2733 5127 2740
rect 5237 2737 5253 2747
rect 5240 2733 5253 2737
rect 5347 2737 5363 2747
rect 5347 2733 5360 2737
rect 5547 2737 5563 2747
rect 5657 2773 5673 2783
rect 5807 2783 5820 2787
rect 5807 2773 5823 2783
rect 5657 2747 5663 2773
rect 5817 2747 5823 2773
rect 5937 2747 5943 2797
rect 5657 2737 5673 2747
rect 5547 2733 5560 2737
rect 5660 2733 5673 2737
rect 5807 2737 5823 2747
rect 5807 2733 5820 2737
rect 5927 2737 5943 2747
rect 5927 2733 5940 2737
rect 5113 2727 5127 2733
rect 2187 2717 2213 2723
rect 2487 2717 2533 2723
rect 2627 2717 2653 2723
rect 5327 2717 5373 2723
rect 947 2677 973 2683
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 1967 2537 2033 2543
rect 1107 2517 1173 2523
rect 1367 2497 1433 2503
rect 1981 2497 2053 2503
rect 2707 2497 2853 2503
rect 3667 2497 3733 2503
rect 4387 2497 4423 2503
rect 167 2483 180 2487
rect 1020 2483 1033 2487
rect 167 2473 183 2483
rect 177 2447 183 2473
rect 1017 2473 1033 2483
rect 1227 2483 1240 2487
rect 1227 2480 1243 2483
rect 1227 2473 1247 2480
rect 2760 2483 2773 2487
rect 2427 2477 2463 2483
rect 177 2437 193 2447
rect 180 2433 193 2437
rect 1017 2423 1023 2473
rect 1233 2466 1247 2473
rect 1257 2447 1263 2473
rect 2457 2447 2463 2477
rect 2757 2473 2773 2483
rect 2927 2483 2940 2487
rect 2927 2473 2943 2483
rect 3107 2483 3120 2487
rect 3107 2473 3123 2483
rect 3367 2483 3380 2487
rect 3367 2473 3383 2483
rect 1257 2437 1273 2447
rect 1260 2433 1273 2437
rect 2457 2437 2473 2447
rect 2460 2433 2473 2437
rect 2757 2443 2763 2473
rect 2937 2447 2943 2473
rect 2727 2437 2763 2443
rect 2927 2437 2943 2447
rect 3117 2447 3123 2473
rect 3377 2447 3383 2473
rect 4417 2447 4423 2497
rect 5977 2497 6013 2503
rect 4687 2483 4700 2487
rect 4687 2473 4703 2483
rect 4827 2483 4840 2487
rect 4827 2473 4843 2483
rect 5107 2483 5120 2487
rect 5107 2473 5123 2483
rect 5687 2483 5700 2487
rect 5687 2473 5703 2483
rect 3117 2437 3133 2447
rect 2927 2433 2940 2437
rect 3120 2433 3133 2437
rect 3377 2437 3393 2447
rect 3380 2433 3393 2437
rect 4407 2437 4423 2447
rect 4697 2443 4703 2473
rect 4837 2447 4843 2473
rect 4697 2437 4733 2443
rect 4407 2433 4420 2437
rect 4827 2437 4843 2447
rect 5117 2447 5123 2473
rect 5697 2447 5703 2473
rect 5837 2477 5873 2483
rect 5837 2447 5843 2477
rect 5977 2447 5983 2497
rect 5117 2437 5133 2447
rect 4827 2433 4840 2437
rect 5120 2433 5133 2437
rect 5697 2437 5713 2447
rect 5700 2433 5713 2437
rect 5827 2437 5843 2447
rect 5827 2433 5840 2437
rect 5967 2437 5983 2447
rect 5967 2433 5980 2437
rect 987 2417 1023 2423
rect 2727 2417 2813 2423
rect 6143 2358 6203 2862
rect 6110 2342 6203 2358
rect 5087 2317 5113 2323
rect 1687 2297 1733 2303
rect 2407 2277 2453 2283
rect 60 2263 73 2267
rect 57 2253 73 2263
rect 507 2263 520 2267
rect 1120 2263 1133 2267
rect 507 2253 523 2263
rect 57 2223 63 2253
rect 200 2243 213 2247
rect 197 2233 213 2243
rect 197 2227 203 2233
rect 57 2217 83 2223
rect 77 2207 83 2217
rect 187 2217 203 2227
rect 517 2227 523 2253
rect 1117 2253 1133 2263
rect 1707 2263 1720 2267
rect 1707 2253 1723 2263
rect 2040 2263 2053 2267
rect 2037 2253 2053 2263
rect 517 2217 533 2227
rect 187 2213 200 2217
rect 520 2213 533 2217
rect 847 2217 873 2223
rect 1117 2223 1123 2253
rect 1717 2227 1723 2253
rect 1097 2217 1123 2223
rect 77 2205 100 2207
rect 77 2197 93 2205
rect 80 2193 93 2197
rect 1097 2203 1103 2217
rect 1567 2217 1613 2223
rect 1717 2217 1733 2227
rect 1720 2213 1733 2217
rect 1877 2223 1883 2253
rect 1857 2217 1883 2223
rect 2037 2227 2043 2253
rect 2177 2227 2183 2273
rect 2387 2263 2400 2267
rect 2387 2253 2403 2263
rect 2707 2263 2720 2267
rect 2707 2253 2723 2263
rect 3227 2263 3240 2267
rect 3227 2253 3243 2263
rect 4027 2263 4040 2267
rect 4060 2263 4073 2267
rect 4027 2253 4043 2263
rect 2037 2217 2053 2227
rect 1047 2197 1103 2203
rect 1857 2203 1863 2217
rect 2040 2213 2053 2217
rect 2177 2217 2193 2227
rect 2180 2213 2193 2217
rect 2397 2223 2403 2253
rect 2717 2226 2723 2253
rect 3237 2227 3243 2253
rect 2397 2217 2433 2223
rect 3227 2217 3243 2227
rect 3877 2223 3883 2253
rect 4037 2227 4043 2253
rect 3877 2217 3903 2223
rect 3227 2213 3240 2217
rect 1827 2197 1893 2203
rect 3897 2203 3903 2217
rect 4027 2217 4043 2227
rect 4057 2253 4073 2263
rect 4867 2257 4893 2263
rect 5067 2257 5123 2263
rect 4057 2227 4063 2253
rect 5117 2227 5123 2257
rect 4057 2217 4073 2227
rect 4027 2213 4040 2217
rect 4060 2213 4073 2217
rect 5117 2217 5133 2227
rect 5120 2213 5133 2217
rect 3897 2197 3933 2203
rect 5347 2177 5413 2183
rect 1987 2157 2073 2163
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 1587 2017 1653 2023
rect 2167 2017 2213 2023
rect 4487 2017 4533 2023
rect 2487 1997 2513 2003
rect 3427 1997 3453 2003
rect 5707 1997 5773 2003
rect 647 1977 673 1983
rect 887 1983 900 1987
rect 887 1973 903 1983
rect 1047 1977 1073 1983
rect 1847 1977 1933 1983
rect 2287 1977 2333 1983
rect 2447 1977 2513 1983
rect 897 1963 903 1973
rect 4187 1977 4233 1983
rect 4587 1977 4623 1983
rect 1740 1963 1753 1967
rect 897 1957 923 1963
rect 917 1927 923 1957
rect 1737 1953 1753 1963
rect 2007 1963 2020 1967
rect 2007 1953 2023 1963
rect 2747 1963 2760 1967
rect 2780 1963 2793 1967
rect 2747 1953 2763 1963
rect 1737 1927 1743 1953
rect 2017 1927 2023 1953
rect 907 1917 923 1927
rect 907 1913 920 1917
rect 1727 1917 1743 1927
rect 1727 1913 1740 1917
rect 2007 1917 2023 1927
rect 2007 1913 2020 1917
rect 2757 1907 2763 1953
rect 2777 1953 2793 1963
rect 4327 1963 4340 1967
rect 4327 1953 4343 1963
rect 2777 1927 2783 1953
rect 2777 1917 2793 1927
rect 2780 1913 2793 1917
rect 4337 1926 4343 1953
rect 4617 1927 4623 1977
rect 5277 1977 5313 1983
rect 5277 1963 5283 1977
rect 5567 1977 5633 1983
rect 5707 1977 5753 1983
rect 4607 1917 4623 1927
rect 5257 1957 5283 1963
rect 4607 1913 4620 1917
rect 2757 1897 2773 1907
rect 2760 1893 2773 1897
rect 2977 1900 3033 1903
rect 2973 1897 3033 1900
rect 2973 1887 2987 1897
rect 4507 1897 4533 1903
rect 5257 1903 5263 1957
rect 5387 1963 5400 1967
rect 5600 1963 5613 1967
rect 5387 1953 5403 1963
rect 5397 1927 5403 1953
rect 5387 1917 5403 1927
rect 5597 1953 5613 1963
rect 5867 1957 5903 1963
rect 5597 1923 5603 1953
rect 5897 1927 5903 1957
rect 5597 1920 5623 1923
rect 5597 1917 5627 1920
rect 5897 1917 5913 1927
rect 5387 1913 5400 1917
rect 5613 1907 5627 1917
rect 5900 1913 5913 1917
rect 5257 1897 5313 1903
rect 5727 1897 5773 1903
rect 6143 1838 6203 2342
rect 6110 1822 6203 1838
rect 5367 1777 5393 1783
rect 187 1743 200 1747
rect 187 1733 203 1743
rect 347 1737 373 1743
rect 197 1707 203 1733
rect 1617 1707 1623 1773
rect 3587 1757 3653 1763
rect 1937 1737 1973 1743
rect 1757 1707 1763 1733
rect 197 1697 213 1707
rect 200 1693 213 1697
rect 1617 1697 1633 1707
rect 1620 1693 1633 1697
rect 1747 1697 1763 1707
rect 1937 1703 1943 1737
rect 2100 1743 2113 1747
rect 2097 1733 2113 1743
rect 2240 1743 2253 1747
rect 2237 1733 2253 1743
rect 3493 1743 3507 1753
rect 5247 1757 5273 1763
rect 3780 1743 3793 1747
rect 3477 1740 3507 1743
rect 3477 1737 3503 1740
rect 2097 1707 2103 1733
rect 1917 1697 1943 1703
rect 1747 1693 1760 1697
rect 1917 1683 1923 1697
rect 2087 1697 2103 1707
rect 2237 1707 2243 1733
rect 3477 1707 3483 1737
rect 3777 1733 3793 1743
rect 4140 1743 4153 1747
rect 4137 1733 4153 1743
rect 4547 1743 4560 1747
rect 4547 1733 4563 1743
rect 5227 1733 5243 1745
rect 3777 1707 3783 1733
rect 4137 1707 4143 1733
rect 2237 1697 2253 1707
rect 2087 1693 2100 1697
rect 2240 1693 2253 1697
rect 3477 1697 3493 1707
rect 3480 1693 3493 1697
rect 3777 1697 3793 1707
rect 3780 1693 3793 1697
rect 4137 1697 4153 1707
rect 4140 1693 4153 1697
rect 1887 1677 1923 1683
rect 2067 1677 2133 1683
rect 2747 1677 2773 1683
rect 4447 1677 4473 1683
rect 4557 1683 4563 1733
rect 5237 1707 5243 1733
rect 5457 1737 5493 1743
rect 5457 1707 5463 1737
rect 5237 1697 5253 1707
rect 5240 1693 5253 1697
rect 5447 1697 5463 1707
rect 5447 1693 5460 1697
rect 4557 1677 4593 1683
rect 1687 1657 1773 1663
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 3447 1537 3493 1543
rect 1887 1477 1973 1483
rect 1147 1457 1233 1463
rect 1627 1457 1653 1463
rect 1747 1457 1813 1463
rect 4267 1457 4373 1463
rect 4747 1457 4793 1463
rect 6047 1457 6073 1463
rect 1960 1443 1973 1447
rect 1957 1433 1973 1443
rect 2207 1443 2220 1447
rect 2900 1443 2913 1447
rect 2207 1433 2223 1443
rect 1957 1407 1963 1433
rect 2217 1407 2223 1433
rect 587 1397 613 1403
rect 1957 1397 1973 1407
rect 1960 1393 1973 1397
rect 2207 1397 2223 1407
rect 2897 1433 2913 1443
rect 3287 1443 3300 1447
rect 3287 1433 3303 1443
rect 3427 1443 3440 1447
rect 3427 1433 3443 1443
rect 2897 1407 2903 1433
rect 2897 1397 2913 1407
rect 2207 1393 2220 1397
rect 2900 1393 2913 1397
rect 3297 1403 3303 1433
rect 3437 1407 3443 1433
rect 4617 1437 4653 1443
rect 4617 1407 4623 1437
rect 5207 1437 5243 1443
rect 3277 1400 3303 1403
rect 3273 1397 3303 1400
rect 3273 1387 3287 1397
rect 3427 1397 3443 1407
rect 3427 1393 3440 1397
rect 4607 1397 4623 1407
rect 5237 1407 5243 1437
rect 5327 1443 5340 1447
rect 5327 1433 5343 1443
rect 5337 1407 5343 1433
rect 5237 1397 5253 1407
rect 4607 1393 4620 1397
rect 5240 1393 5253 1397
rect 5337 1397 5353 1407
rect 5340 1393 5353 1397
rect 6067 1397 6113 1403
rect 1487 1377 1533 1383
rect 3447 1377 3493 1383
rect 5947 1357 5993 1363
rect 6143 1318 6203 1822
rect 6110 1302 6203 1318
rect 4447 1237 4473 1243
rect 2287 1223 2300 1227
rect 3020 1223 3033 1227
rect 2287 1213 2303 1223
rect 47 1203 60 1207
rect 47 1193 63 1203
rect 57 1187 63 1193
rect 57 1177 73 1187
rect 60 1173 73 1177
rect 2297 1183 2303 1213
rect 3017 1213 3033 1223
rect 3627 1223 3640 1227
rect 3627 1213 3643 1223
rect 3727 1223 3740 1227
rect 3760 1223 3773 1227
rect 3727 1213 3743 1223
rect 3017 1187 3023 1213
rect 3637 1187 3643 1213
rect 2297 1177 2353 1183
rect 3017 1177 3033 1187
rect 3020 1173 3033 1177
rect 3637 1177 3653 1187
rect 3640 1173 3653 1177
rect 587 1157 613 1163
rect 1207 1157 1233 1163
rect 3737 1163 3743 1213
rect 3757 1213 3773 1223
rect 5513 1223 5527 1233
rect 5497 1220 5527 1223
rect 5497 1217 5523 1220
rect 3757 1187 3763 1213
rect 3757 1177 3773 1187
rect 3760 1173 3773 1177
rect 5497 1183 5503 1217
rect 5467 1177 5503 1183
rect 3737 1157 3793 1163
rect 3907 1157 3953 1163
rect 5227 1157 5293 1163
rect 6077 1147 6083 1193
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 3167 1017 3193 1023
rect 2173 963 2187 973
rect 2127 960 2187 963
rect 2127 957 2183 960
rect 5067 957 5093 963
rect 127 937 253 943
rect 1027 937 1073 943
rect 1207 937 1313 943
rect 1507 937 1553 943
rect 2547 937 2633 943
rect 4181 937 4213 943
rect 4307 937 4393 943
rect 5667 937 5693 943
rect 1587 917 1613 923
rect 1987 917 2013 923
rect 4047 923 4060 927
rect 5080 923 5093 927
rect 4047 913 4063 923
rect 4057 883 4063 913
rect 5077 913 5093 923
rect 5220 923 5233 927
rect 5217 913 5233 923
rect 5467 923 5480 927
rect 5467 913 5483 923
rect 5077 887 5083 913
rect 5217 887 5223 913
rect 5477 887 5483 913
rect 4057 880 4083 883
rect 4057 877 4087 880
rect 5077 877 5093 887
rect 4073 867 4087 877
rect 5080 873 5093 877
rect 5207 877 5223 887
rect 5207 873 5220 877
rect 5467 877 5483 887
rect 5467 873 5480 877
rect 3287 857 3333 863
rect 6143 798 6203 1302
rect 6110 782 6203 798
rect 1867 717 1893 723
rect 2987 717 3053 723
rect 3927 717 3973 723
rect 4267 717 4333 723
rect 4900 723 4913 727
rect 4897 713 4913 723
rect 1287 703 1300 707
rect 1287 693 1303 703
rect 1727 703 1740 707
rect 1727 693 1743 703
rect 1297 667 1303 693
rect 1297 657 1313 667
rect 1300 653 1313 657
rect 1737 663 1743 693
rect 2037 697 2073 703
rect 2037 667 2043 697
rect 2220 703 2233 707
rect 2217 693 2233 703
rect 2967 697 3013 703
rect 4897 703 4903 713
rect 5820 703 5833 707
rect 4877 697 4903 703
rect 2217 683 2223 693
rect 2197 677 2223 683
rect 2197 667 2203 677
rect 3153 667 3167 673
rect 3177 667 3183 693
rect 1737 660 1783 663
rect 1737 657 1787 660
rect 1773 647 1787 657
rect 2027 657 2043 667
rect 2027 653 2040 657
rect 2187 657 2203 667
rect 2187 653 2200 657
rect 3147 660 3167 667
rect 3147 657 3163 660
rect 3147 653 3160 657
rect 3727 657 3753 663
rect 3777 647 3783 673
rect 4877 667 4883 697
rect 5817 693 5833 703
rect 5817 667 5823 693
rect 4867 657 4883 667
rect 4867 653 4880 657
rect 5807 657 5823 667
rect 5807 653 5820 657
rect 1547 637 1673 643
rect 3847 637 3953 643
rect -63 522 30 538
rect -63 18 -3 522
rect 467 417 493 423
rect 2127 417 2273 423
rect 2727 417 2793 423
rect 2807 417 2873 423
rect 5867 417 5913 423
rect 1517 397 1593 403
rect 2200 403 2213 407
rect 2197 393 2213 403
rect 3227 403 3240 407
rect 3260 403 3273 407
rect 3227 393 3243 403
rect 2197 363 2203 393
rect 3237 367 3243 393
rect 2177 360 2203 363
rect 2173 357 2203 360
rect 2173 347 2187 357
rect 3227 357 3243 367
rect 3257 393 3273 403
rect 3227 353 3240 357
rect 3257 347 3263 393
rect 887 337 933 343
rect 1707 337 1793 343
rect 3240 346 3263 347
rect 3247 337 3263 346
rect 3247 333 3260 337
rect 3627 337 3673 343
rect 2027 317 2053 323
rect 1687 297 1753 303
rect 6143 278 6203 782
rect 6110 262 6203 278
rect 1627 237 1673 243
rect 2847 197 2913 203
rect 1487 177 1533 183
rect 2540 183 2553 187
rect 2537 173 2553 183
rect 2967 183 2980 187
rect 2967 173 2983 183
rect 4147 183 4160 187
rect 4440 183 4453 187
rect 4147 173 4163 183
rect 2537 147 2543 173
rect 2107 137 2133 143
rect 2527 137 2543 147
rect 2977 147 2983 173
rect 4000 163 4013 167
rect 3997 157 4013 163
rect 4000 153 4013 157
rect 2977 137 2993 147
rect 2527 133 2540 137
rect 2980 133 2993 137
rect 4157 143 4163 173
rect 4437 173 4453 183
rect 4437 147 4443 173
rect 3847 137 3903 143
rect 4157 137 4183 143
rect 587 117 673 123
rect 1007 117 1093 123
rect 1166 113 1167 120
rect 1187 117 1253 123
rect 2087 117 2193 123
rect 4177 123 4183 137
rect 4427 137 4443 147
rect 4427 133 4440 137
rect 4177 117 4213 123
rect 5987 117 6073 123
rect 1153 103 1167 113
rect 1153 100 1233 103
rect 1157 97 1233 100
rect 2807 37 2833 43
rect -63 2 30 18
rect 6143 2 6203 262
<< m2contact >>
rect 2273 6134 2287 6148
rect 2333 6133 2347 6147
rect 2533 6133 2547 6147
rect 2653 6133 2667 6147
rect 3913 6133 3927 6147
rect 5593 6133 5607 6147
rect 5693 6133 5707 6147
rect 4013 6113 4027 6127
rect 5913 6113 5927 6127
rect 4573 6093 4587 6107
rect 3913 6073 3927 6087
rect 4053 6073 4067 6087
rect 4733 6073 4747 6087
rect 5913 6073 5927 6087
rect 5173 6053 5187 6067
rect 5253 6053 5267 6067
rect 2847 5933 2861 5947
rect 2893 5933 2907 5947
rect 2133 5913 2147 5927
rect 2193 5913 2207 5927
rect 2793 5913 2807 5927
rect 2853 5913 2867 5927
rect 4273 5913 4287 5927
rect 4353 5913 4367 5927
rect 193 5893 207 5907
rect 3713 5893 3727 5907
rect 5293 5893 5307 5907
rect 193 5853 207 5867
rect 2973 5853 2987 5867
rect 3013 5853 3027 5867
rect 3673 5852 3687 5866
rect 5293 5853 5307 5867
rect 5633 5893 5647 5907
rect 5633 5853 5647 5867
rect 2573 5833 2587 5847
rect 2653 5833 2667 5847
rect 4173 5833 4187 5847
rect 4233 5833 4247 5847
rect 5433 5833 5447 5847
rect 5513 5833 5527 5847
rect 373 5613 387 5627
rect 433 5613 447 5627
rect 2213 5613 2227 5627
rect 2253 5613 2267 5627
rect 2293 5613 2307 5627
rect 2993 5613 3007 5627
rect 3053 5613 3067 5627
rect 4873 5613 4887 5627
rect 4913 5614 4927 5628
rect 513 5593 527 5607
rect 513 5553 527 5567
rect 553 5553 567 5567
rect 4373 5593 4387 5607
rect 4813 5593 4827 5607
rect 5313 5573 5327 5587
rect 5493 5573 5507 5587
rect 2273 5553 2287 5567
rect 4453 5553 4467 5567
rect 4893 5553 4907 5567
rect 553 5532 567 5546
rect 1093 5533 1107 5547
rect 1153 5533 1167 5547
rect 3447 5533 3461 5547
rect 3493 5533 3507 5547
rect 5133 5533 5147 5547
rect 5193 5533 5207 5547
rect 5233 5533 5247 5547
rect 1633 5513 1647 5527
rect 1713 5513 1727 5527
rect 1913 5493 1927 5507
rect 1973 5493 1987 5507
rect 1073 5393 1087 5407
rect 2613 5373 2627 5387
rect 2693 5373 2707 5387
rect 2833 5373 2847 5387
rect 1133 5333 1147 5347
rect 1553 5333 1567 5347
rect 2613 5333 2627 5347
rect 2693 5333 2707 5347
rect 2833 5333 2847 5347
rect 2973 5373 2987 5387
rect 3173 5373 3187 5387
rect 2973 5333 2987 5347
rect 3173 5333 3187 5347
rect 3393 5373 3407 5387
rect 3633 5373 3647 5387
rect 4353 5373 4367 5387
rect 5633 5373 5647 5387
rect 3393 5333 3407 5347
rect 3633 5333 3647 5347
rect 4233 5333 4247 5347
rect 4273 5333 4287 5347
rect 4353 5333 4367 5347
rect 5573 5333 5587 5347
rect 1113 5313 1127 5327
rect 1153 5313 1167 5327
rect 1973 5313 1987 5327
rect 2053 5313 2067 5327
rect 2373 5313 2387 5327
rect 2513 5313 2527 5327
rect 3193 5313 3207 5327
rect 3273 5313 3287 5327
rect 3313 5313 3327 5327
rect 3373 5312 3387 5326
rect 4693 5313 4707 5327
rect 4773 5313 4787 5327
rect 2553 5293 2567 5307
rect 2633 5293 2647 5307
rect 4153 5173 4167 5187
rect 4193 5173 4207 5187
rect 1693 5073 1707 5087
rect 2433 5073 2447 5087
rect 2593 5073 2607 5087
rect 3193 5073 3207 5087
rect 3233 5073 3247 5087
rect 3513 5073 3527 5087
rect 3553 5072 3567 5086
rect 3653 5073 3667 5087
rect 4053 5093 4067 5107
rect 1153 5033 1167 5047
rect 1193 5033 1207 5047
rect 1693 5033 1707 5047
rect 2473 5033 2487 5047
rect 2653 5033 2667 5047
rect 2733 5033 2747 5047
rect 2773 5033 2787 5047
rect 3653 5033 3667 5047
rect 3973 5033 3987 5047
rect 4193 5073 4207 5087
rect 4653 5073 4667 5087
rect 4753 5073 4767 5087
rect 5113 5093 5127 5107
rect 5193 5073 5207 5087
rect 4193 5033 4207 5047
rect 4653 5033 4667 5047
rect 4793 5033 4807 5047
rect 5033 5033 5047 5047
rect 1393 5013 1407 5027
rect 1553 5013 1567 5027
rect 3213 5013 3227 5027
rect 3253 5013 3267 5027
rect 5393 5073 5407 5087
rect 5333 5033 5347 5047
rect 5253 5013 5267 5027
rect 5713 4913 5727 4927
rect 5753 4913 5767 4927
rect 2093 4873 2107 4887
rect 2133 4873 2147 4887
rect 2613 4872 2627 4886
rect 2673 4873 2687 4887
rect 2733 4853 2747 4867
rect 2613 4813 2627 4827
rect 2733 4813 2747 4827
rect 2813 4853 2827 4867
rect 3053 4853 3067 4867
rect 913 4793 927 4807
rect 1013 4793 1027 4807
rect 2273 4793 2287 4807
rect 2333 4793 2347 4807
rect 3373 4853 3387 4867
rect 3593 4853 3607 4867
rect 2793 4792 2807 4806
rect 3133 4793 3147 4807
rect 3313 4793 3327 4807
rect 3593 4813 3607 4827
rect 4153 4873 4167 4887
rect 4633 4873 4647 4887
rect 4693 4873 4707 4887
rect 4333 4853 4347 4867
rect 4533 4853 4547 4867
rect 4673 4853 4687 4867
rect 4813 4853 4827 4867
rect 4913 4853 4927 4867
rect 4093 4813 4107 4827
rect 4333 4813 4347 4827
rect 4493 4813 4507 4827
rect 4633 4813 4647 4827
rect 4813 4813 4827 4827
rect 5153 4853 5167 4867
rect 5333 4873 5347 4887
rect 4973 4813 4987 4827
rect 5153 4813 5167 4827
rect 5253 4813 5267 4827
rect 5453 4853 5467 4867
rect 5853 4853 5867 4867
rect 6073 4833 6087 4847
rect 5453 4813 5467 4827
rect 5853 4813 5867 4827
rect 5893 4813 5907 4827
rect 5053 4793 5067 4807
rect 5113 4793 5127 4807
rect 5673 4793 5687 4807
rect 5753 4793 5767 4807
rect 4473 4753 4487 4767
rect 4513 4753 4527 4767
rect 5993 4713 6007 4727
rect 5173 4653 5187 4667
rect 5253 4653 5267 4667
rect 4653 4613 4667 4627
rect 4733 4613 4747 4627
rect 393 4574 407 4588
rect 473 4573 487 4587
rect 2913 4573 2927 4587
rect 5053 4573 5067 4587
rect 5993 4573 6007 4587
rect 1293 4553 1307 4567
rect 2433 4553 2447 4567
rect 613 4533 627 4547
rect 993 4533 1007 4547
rect 2793 4553 2807 4567
rect 2613 4533 2627 4547
rect 653 4513 667 4527
rect 813 4513 827 4527
rect 1333 4513 1347 4527
rect 1413 4513 1427 4527
rect 1453 4513 1467 4527
rect 2753 4513 2767 4527
rect 3513 4553 3527 4567
rect 4673 4553 4687 4567
rect 3333 4533 3347 4547
rect 3493 4533 3507 4547
rect 2893 4513 2907 4527
rect 4733 4533 4747 4547
rect 4673 4513 4687 4527
rect 4913 4513 4927 4527
rect 5013 4513 5027 4527
rect 5073 4553 5087 4567
rect 5473 4553 5487 4567
rect 5073 4513 5087 4527
rect 5633 4553 5647 4567
rect 1693 4493 1707 4507
rect 1773 4493 1787 4507
rect 1993 4493 2007 4507
rect 2053 4493 2067 4507
rect 3493 4493 3507 4507
rect 5893 4513 5907 4527
rect 5973 4513 5987 4527
rect 5553 4493 5567 4507
rect 1233 4393 1247 4407
rect 1273 4393 1287 4407
rect 4593 4373 4607 4387
rect 433 4333 447 4347
rect 2453 4333 2467 4347
rect 2673 4333 2687 4347
rect 1573 4313 1587 4327
rect 953 4293 967 4307
rect 1433 4292 1447 4306
rect 2493 4313 2507 4327
rect 4433 4333 4447 4347
rect 4553 4332 4567 4346
rect 4673 4353 4687 4367
rect 4773 4353 4787 4367
rect 5213 4353 5227 4367
rect 5293 4353 5307 4367
rect 4713 4333 4727 4347
rect 5013 4333 5027 4347
rect 5113 4333 5127 4347
rect 493 4273 507 4287
rect 1353 4273 1367 4287
rect 4773 4293 4787 4307
rect 4953 4293 4967 4307
rect 5353 4333 5367 4347
rect 5513 4333 5527 4347
rect 5553 4333 5567 4347
rect 5713 4333 5727 4347
rect 5813 4333 5827 4347
rect 5173 4293 5187 4307
rect 5353 4293 5367 4307
rect 2013 4273 2027 4287
rect 2113 4273 2127 4287
rect 2513 4273 2527 4287
rect 4513 4273 4527 4287
rect 4593 4273 4607 4287
rect 4653 4273 4667 4287
rect 4753 4273 4767 4287
rect 5733 4273 5747 4287
rect 5793 4273 5807 4287
rect 2573 4193 2587 4207
rect 2653 4093 2667 4107
rect 2673 4093 2687 4107
rect 193 4053 207 4067
rect 273 4053 287 4067
rect 1773 4053 1787 4067
rect 1853 4053 1867 4067
rect 1953 4053 1967 4067
rect 2013 4053 2027 4067
rect 2353 4053 2367 4067
rect 2393 4053 2407 4067
rect 4073 4053 4087 4067
rect 4153 4053 4167 4067
rect 4313 4053 4327 4067
rect 4413 4052 4427 4066
rect 5193 4053 5207 4067
rect 5293 4053 5307 4067
rect 5693 4053 5707 4067
rect 5753 4052 5767 4066
rect 5913 4054 5927 4068
rect 5993 4053 6007 4067
rect 893 4033 907 4047
rect 1593 4033 1607 4047
rect 1653 4033 1667 4047
rect 1093 4013 1107 4027
rect 453 3993 467 4007
rect 513 3993 527 4007
rect 1593 3993 1607 4007
rect 1873 4033 1887 4047
rect 1993 4033 2007 4047
rect 1733 3993 1747 4007
rect 1833 3993 1847 4007
rect 2133 4033 2147 4047
rect 2773 4033 2787 4047
rect 2073 3993 2087 4007
rect 2773 3993 2787 4007
rect 2953 4033 2967 4047
rect 4233 4033 4247 4047
rect 4613 4033 4627 4047
rect 2953 3993 2967 4007
rect 1953 3973 1967 3987
rect 2333 3973 2347 3987
rect 2373 3973 2387 3987
rect 4253 3973 4267 3987
rect 4493 3973 4507 3987
rect 4553 3973 4567 3987
rect 5113 4033 5127 4047
rect 5393 4033 5407 4047
rect 6073 4054 6087 4068
rect 5553 4013 5567 4027
rect 4913 3993 4927 4007
rect 5113 3993 5127 4007
rect 5333 3993 5347 4007
rect 6013 3993 6027 4007
rect 4633 3952 4647 3966
rect 2613 3873 2627 3887
rect 2653 3872 2667 3886
rect 2633 3852 2647 3866
rect 2713 3853 2727 3867
rect 5673 3853 5687 3867
rect 5713 3853 5727 3867
rect 1493 3833 1507 3847
rect 773 3813 787 3827
rect 853 3813 867 3827
rect 893 3813 907 3827
rect 1233 3813 1247 3827
rect 1353 3813 1367 3827
rect 1613 3833 1627 3847
rect 1933 3833 1947 3847
rect 4953 3833 4967 3847
rect 4993 3833 5007 3847
rect 5033 3833 5047 3847
rect 5793 3833 5807 3847
rect 5873 3833 5887 3847
rect 773 3773 787 3787
rect 1233 3773 1247 3787
rect 1373 3773 1387 3787
rect 1553 3773 1567 3787
rect 1633 3773 1647 3787
rect 1893 3773 1907 3787
rect 1953 3813 1967 3827
rect 2133 3813 2147 3827
rect 2813 3813 2827 3827
rect 3973 3813 3987 3827
rect 5673 3813 5687 3827
rect 1953 3773 1967 3787
rect 2053 3773 2067 3787
rect 913 3753 927 3767
rect 973 3753 987 3767
rect 1713 3751 1727 3765
rect 1753 3753 1767 3767
rect 2073 3753 2087 3767
rect 2133 3753 2147 3767
rect 5813 3813 5827 3827
rect 5933 3813 5947 3827
rect 3993 3772 4007 3786
rect 5733 3773 5747 3787
rect 5853 3773 5867 3787
rect 5933 3773 5947 3787
rect 2793 3752 2807 3766
rect 3053 3753 3067 3767
rect 3133 3753 3147 3767
rect 5613 3753 5627 3767
rect 5753 3753 5767 3767
rect 5793 3751 5807 3765
rect 5873 3753 5887 3767
rect 2673 3613 2687 3627
rect 2713 3613 2727 3627
rect 1853 3573 1867 3587
rect 1933 3573 1947 3587
rect 1553 3553 1567 3567
rect 1653 3553 1667 3567
rect 53 3533 67 3547
rect 133 3533 147 3547
rect 493 3533 507 3547
rect 593 3533 607 3547
rect 1633 3513 1647 3527
rect 1953 3533 1967 3547
rect 2793 3533 2807 3547
rect 2853 3533 2867 3547
rect 5473 3533 5487 3547
rect 5533 3533 5547 3547
rect 1893 3492 1907 3506
rect 2053 3513 2067 3527
rect 3773 3513 3787 3527
rect 3813 3513 3827 3527
rect 4473 3513 4487 3527
rect 5333 3513 5347 3527
rect 1633 3473 1647 3487
rect 2053 3473 2067 3487
rect 4433 3473 4447 3487
rect 5713 3533 5727 3547
rect 6013 3513 6027 3527
rect 5333 3473 5347 3487
rect 5633 3473 5647 3487
rect 5953 3473 5967 3487
rect 2253 3453 2267 3467
rect 2353 3453 2367 3467
rect 2493 3353 2507 3367
rect 2553 3353 2567 3367
rect 3033 3353 3047 3367
rect 2373 3313 2387 3327
rect 3033 3313 3047 3327
rect 5153 3313 5167 3327
rect 593 3293 607 3307
rect 593 3253 607 3267
rect 653 3293 667 3307
rect 753 3293 767 3307
rect 753 3253 767 3267
rect 1553 3293 1567 3307
rect 1613 3293 1627 3307
rect 1933 3293 1947 3307
rect 1553 3253 1567 3267
rect 453 3233 467 3247
rect 513 3233 527 3247
rect 633 3233 647 3247
rect 1193 3233 1207 3247
rect 1273 3233 1287 3247
rect 1933 3253 1947 3267
rect 2393 3293 2407 3307
rect 2633 3293 2647 3307
rect 2873 3293 2887 3307
rect 3373 3293 3387 3307
rect 4053 3293 4067 3307
rect 2393 3253 2407 3267
rect 2633 3253 2647 3267
rect 4873 3293 4887 3307
rect 2933 3253 2947 3267
rect 3373 3253 3387 3267
rect 4053 3253 4067 3267
rect 4413 3253 4427 3267
rect 4813 3253 4827 3267
rect 5093 3253 5107 3267
rect 5533 3293 5547 3307
rect 5953 3292 5967 3306
rect 5533 3253 5547 3267
rect 1693 3233 1707 3247
rect 2333 3233 2347 3247
rect 2413 3233 2427 3247
rect 2493 3233 2507 3247
rect 2553 3231 2567 3245
rect 3873 3233 3887 3247
rect 3993 3233 4007 3247
rect 4413 3232 4427 3246
rect 4453 3233 4467 3247
rect 4933 3233 4947 3247
rect 5013 3233 5027 3247
rect 4393 3212 4407 3226
rect 6033 3212 6047 3226
rect 5633 3192 5647 3206
rect 5673 3193 5687 3207
rect 2093 3093 2107 3107
rect 2153 3093 2167 3107
rect 273 3013 287 3027
rect 393 3013 407 3027
rect 1653 3013 1667 3027
rect 1713 3013 1727 3027
rect 1933 3013 1947 3027
rect 2033 3013 2047 3027
rect 2713 3013 2727 3027
rect 2753 3013 2767 3027
rect 2813 3014 2827 3028
rect 2893 3012 2907 3026
rect 1073 2993 1087 3007
rect 1413 2993 1427 3007
rect 1813 2992 1827 3006
rect 1853 2993 1867 3007
rect 1953 2993 1967 3007
rect 793 2953 807 2967
rect 853 2953 867 2967
rect 1073 2953 1087 2967
rect 1333 2953 1347 2967
rect 2173 2993 2187 3007
rect 2573 2993 2587 3007
rect 3053 2993 3067 3007
rect 3173 2993 3187 3007
rect 3273 2993 3287 3007
rect 2173 2953 2187 2967
rect 1973 2933 1987 2947
rect 2233 2933 2247 2947
rect 2333 2933 2347 2947
rect 2593 2933 2607 2947
rect 3173 2953 3187 2967
rect 3273 2953 3287 2967
rect 4013 2993 4027 3007
rect 4093 2993 4107 3007
rect 4273 2993 4287 3007
rect 5333 2993 5347 3007
rect 5653 2993 5667 3007
rect 4013 2953 4027 2967
rect 4173 2953 4187 2967
rect 4313 2953 4327 2967
rect 4933 2953 4947 2967
rect 4973 2953 4987 2967
rect 5333 2953 5347 2967
rect 5593 2953 5607 2967
rect 3033 2932 3047 2946
rect 5153 2933 5167 2947
rect 5213 2933 5227 2947
rect 5813 2913 5827 2927
rect 5873 2913 5887 2927
rect 5533 2833 5547 2847
rect 5673 2833 5687 2847
rect 1633 2813 1647 2827
rect 1713 2813 1727 2827
rect 5553 2813 5567 2827
rect 5653 2813 5667 2827
rect 1473 2793 1487 2807
rect 1513 2793 1527 2807
rect 973 2773 987 2787
rect 973 2733 987 2747
rect 413 2713 427 2727
rect 533 2713 547 2727
rect 873 2713 887 2727
rect 953 2713 967 2727
rect 1593 2792 1607 2806
rect 1913 2793 1927 2807
rect 1993 2793 2007 2807
rect 2453 2793 2467 2807
rect 2533 2793 2547 2807
rect 5353 2793 5367 2807
rect 5433 2792 5447 2806
rect 5513 2793 5527 2807
rect 1713 2773 1727 2787
rect 2113 2773 2127 2787
rect 2253 2773 2267 2787
rect 2093 2752 2107 2766
rect 1633 2733 1647 2747
rect 2513 2773 2527 2787
rect 2793 2773 2807 2787
rect 3033 2773 3047 2787
rect 2593 2753 2607 2767
rect 3293 2773 3307 2787
rect 5113 2773 5127 2787
rect 5213 2773 5227 2787
rect 5333 2773 5347 2787
rect 3093 2753 3107 2767
rect 3253 2753 3267 2767
rect 2253 2733 2267 2747
rect 2453 2733 2467 2747
rect 2573 2733 2587 2747
rect 2753 2733 2767 2747
rect 3033 2733 3047 2747
rect 5073 2752 5087 2766
rect 5413 2773 5427 2787
rect 5373 2753 5387 2767
rect 5753 2793 5767 2807
rect 5813 2793 5827 2807
rect 5893 2794 5907 2808
rect 3293 2733 3307 2747
rect 5093 2733 5107 2747
rect 5253 2733 5267 2747
rect 5333 2733 5347 2747
rect 5533 2733 5547 2747
rect 5673 2773 5687 2787
rect 5793 2773 5807 2787
rect 5673 2733 5687 2747
rect 5793 2733 5807 2747
rect 5913 2733 5927 2747
rect 1533 2712 1547 2726
rect 2173 2713 2187 2727
rect 2213 2713 2227 2727
rect 2473 2713 2487 2727
rect 2533 2713 2547 2727
rect 2613 2713 2627 2727
rect 2653 2713 2667 2727
rect 5113 2713 5127 2727
rect 5313 2711 5327 2725
rect 5373 2713 5387 2727
rect 933 2673 947 2687
rect 973 2673 987 2687
rect 1953 2533 1967 2547
rect 2033 2533 2047 2547
rect 1093 2513 1107 2527
rect 1173 2513 1187 2527
rect 1353 2493 1367 2507
rect 1433 2493 1447 2507
rect 1967 2493 1981 2507
rect 2053 2493 2067 2507
rect 2693 2493 2707 2507
rect 2853 2493 2867 2507
rect 3653 2493 3667 2507
rect 3733 2494 3747 2508
rect 4373 2493 4387 2507
rect 153 2473 167 2487
rect 1033 2473 1047 2487
rect 1213 2473 1227 2487
rect 1253 2473 1267 2487
rect 2413 2473 2427 2487
rect 193 2433 207 2447
rect 973 2413 987 2427
rect 1233 2452 1247 2466
rect 2773 2473 2787 2487
rect 2913 2473 2927 2487
rect 3093 2473 3107 2487
rect 3353 2473 3367 2487
rect 1273 2433 1287 2447
rect 2473 2433 2487 2447
rect 2713 2433 2727 2447
rect 2913 2433 2927 2447
rect 4673 2473 4687 2487
rect 4813 2473 4827 2487
rect 5093 2473 5107 2487
rect 5673 2473 5687 2487
rect 3133 2433 3147 2447
rect 3393 2433 3407 2447
rect 4393 2433 4407 2447
rect 4733 2433 4747 2447
rect 4813 2433 4827 2447
rect 5873 2473 5887 2487
rect 6013 2493 6027 2507
rect 5133 2433 5147 2447
rect 5713 2433 5727 2447
rect 5813 2433 5827 2447
rect 5953 2433 5967 2447
rect 2713 2412 2727 2426
rect 2813 2413 2827 2427
rect 5073 2313 5087 2327
rect 5113 2313 5127 2327
rect 1673 2293 1687 2307
rect 1733 2293 1747 2307
rect 2173 2273 2187 2287
rect 2393 2273 2407 2287
rect 2453 2273 2467 2287
rect 73 2253 87 2267
rect 493 2253 507 2267
rect 213 2233 227 2247
rect 173 2213 187 2227
rect 1133 2253 1147 2267
rect 1693 2253 1707 2267
rect 1873 2253 1887 2267
rect 2053 2253 2067 2267
rect 533 2213 547 2227
rect 833 2213 847 2227
rect 873 2213 887 2227
rect 93 2191 107 2205
rect 1033 2193 1047 2207
rect 1553 2213 1567 2227
rect 1613 2213 1627 2227
rect 1733 2213 1747 2227
rect 2373 2253 2387 2267
rect 2693 2253 2707 2267
rect 3213 2253 3227 2267
rect 3873 2253 3887 2267
rect 4013 2253 4027 2267
rect 1813 2193 1827 2207
rect 2053 2213 2067 2227
rect 2193 2213 2207 2227
rect 2433 2212 2447 2226
rect 2713 2212 2727 2226
rect 3213 2213 3227 2227
rect 1893 2193 1907 2207
rect 4013 2213 4027 2227
rect 4073 2253 4087 2267
rect 4853 2253 4867 2267
rect 4893 2253 4907 2267
rect 5053 2253 5067 2267
rect 4073 2213 4087 2227
rect 5133 2213 5147 2227
rect 3933 2193 3947 2207
rect 5333 2173 5347 2187
rect 5413 2173 5427 2187
rect 1973 2153 1987 2167
rect 2073 2153 2087 2167
rect 1573 2013 1587 2027
rect 1653 2013 1667 2027
rect 2153 2013 2167 2027
rect 2213 2013 2227 2027
rect 4473 2013 4487 2027
rect 4533 2013 4547 2027
rect 2473 1993 2487 2007
rect 2513 1993 2527 2007
rect 3413 1993 3427 2007
rect 3453 1993 3467 2007
rect 5693 1993 5707 2007
rect 5773 1992 5787 2006
rect 633 1973 647 1987
rect 673 1973 687 1987
rect 873 1973 887 1987
rect 1033 1973 1047 1987
rect 1073 1973 1087 1987
rect 1833 1973 1847 1987
rect 1933 1973 1947 1987
rect 2273 1973 2287 1987
rect 2333 1973 2347 1987
rect 2433 1973 2447 1987
rect 2513 1972 2527 1986
rect 4173 1973 4187 1987
rect 4233 1973 4247 1987
rect 4573 1973 4587 1987
rect 1753 1953 1767 1967
rect 1993 1953 2007 1967
rect 2733 1953 2747 1967
rect 893 1913 907 1927
rect 1713 1913 1727 1927
rect 1993 1913 2007 1927
rect 2793 1953 2807 1967
rect 4313 1953 4327 1967
rect 2793 1913 2807 1927
rect 5313 1973 5327 1987
rect 5553 1973 5567 1987
rect 5633 1973 5647 1987
rect 5693 1972 5707 1986
rect 5753 1973 5767 1987
rect 4333 1912 4347 1926
rect 4593 1913 4607 1927
rect 2773 1893 2787 1907
rect 3033 1893 3047 1907
rect 4493 1893 4507 1907
rect 4533 1893 4547 1907
rect 5373 1953 5387 1967
rect 5373 1913 5387 1927
rect 5613 1953 5627 1967
rect 5853 1953 5867 1967
rect 5913 1913 5927 1927
rect 5313 1893 5327 1907
rect 5613 1893 5627 1907
rect 5713 1893 5727 1907
rect 5773 1893 5787 1907
rect 2973 1873 2987 1887
rect 1613 1773 1627 1787
rect 5353 1773 5367 1787
rect 5393 1773 5407 1787
rect 173 1733 187 1747
rect 333 1733 347 1747
rect 373 1733 387 1747
rect 3493 1753 3507 1767
rect 3573 1753 3587 1767
rect 3653 1753 3667 1767
rect 1753 1733 1767 1747
rect 213 1693 227 1707
rect 1633 1693 1647 1707
rect 1733 1693 1747 1707
rect 1973 1733 1987 1747
rect 2113 1733 2127 1747
rect 2253 1733 2267 1747
rect 5233 1752 5247 1766
rect 5273 1753 5287 1767
rect 1873 1673 1887 1687
rect 2073 1693 2087 1707
rect 3793 1733 3807 1747
rect 4153 1733 4167 1747
rect 4533 1733 4547 1747
rect 5213 1733 5227 1747
rect 2253 1693 2267 1707
rect 3493 1693 3507 1707
rect 3793 1693 3807 1707
rect 4153 1693 4167 1707
rect 2053 1673 2067 1687
rect 2133 1673 2147 1687
rect 2733 1671 2747 1685
rect 2773 1673 2787 1687
rect 4433 1673 4447 1687
rect 4473 1673 4487 1687
rect 5493 1733 5507 1747
rect 5253 1693 5267 1707
rect 5433 1693 5447 1707
rect 4593 1671 4607 1685
rect 1673 1653 1687 1667
rect 1773 1653 1787 1667
rect 5671 1593 5685 1607
rect 3433 1533 3447 1547
rect 3493 1533 3507 1547
rect 5913 1517 5927 1531
rect 1873 1473 1887 1487
rect 1973 1473 1987 1487
rect 1133 1453 1147 1467
rect 1233 1453 1247 1467
rect 1613 1453 1627 1467
rect 1653 1453 1667 1467
rect 1733 1453 1747 1467
rect 1813 1453 1827 1467
rect 4253 1453 4267 1467
rect 4373 1453 4387 1467
rect 4733 1453 4747 1467
rect 4793 1453 4807 1467
rect 6033 1453 6047 1467
rect 6073 1453 6087 1467
rect 1973 1433 1987 1447
rect 2193 1433 2207 1447
rect 573 1393 587 1407
rect 613 1393 627 1407
rect 1973 1393 1987 1407
rect 2193 1393 2207 1407
rect 2913 1433 2927 1447
rect 3273 1433 3287 1447
rect 3413 1433 3427 1447
rect 2913 1393 2927 1407
rect 4653 1433 4667 1447
rect 5193 1433 5207 1447
rect 3413 1393 3427 1407
rect 4593 1393 4607 1407
rect 5313 1433 5327 1447
rect 5253 1393 5267 1407
rect 5353 1393 5367 1407
rect 6053 1393 6067 1407
rect 6113 1393 6127 1407
rect 1473 1373 1487 1387
rect 1533 1373 1547 1387
rect 3273 1373 3287 1387
rect 3433 1372 3447 1386
rect 3493 1373 3507 1387
rect 5933 1353 5947 1367
rect 5993 1353 6007 1367
rect 4433 1233 4447 1247
rect 4473 1233 4487 1247
rect 5513 1233 5527 1247
rect 2273 1213 2287 1227
rect 33 1193 47 1207
rect 73 1173 87 1187
rect 3033 1213 3047 1227
rect 3613 1213 3627 1227
rect 3713 1213 3727 1227
rect 2353 1173 2367 1187
rect 3033 1173 3047 1187
rect 3653 1173 3667 1187
rect 573 1153 587 1167
rect 613 1151 627 1165
rect 1193 1153 1207 1167
rect 1233 1153 1247 1167
rect 3773 1213 3787 1227
rect 3773 1173 3787 1187
rect 5453 1173 5467 1187
rect 6073 1193 6087 1207
rect 3793 1153 3807 1167
rect 3893 1153 3907 1167
rect 3953 1153 3967 1167
rect 5213 1153 5227 1167
rect 5293 1153 5307 1167
rect 6073 1133 6087 1147
rect 6009 1093 6023 1107
rect 3153 1012 3167 1026
rect 3193 1013 3207 1027
rect 2173 973 2187 987
rect 2113 953 2127 967
rect 5053 953 5067 967
rect 5093 953 5107 967
rect 113 933 127 947
rect 253 933 267 947
rect 1013 933 1027 947
rect 1073 933 1087 947
rect 1193 933 1207 947
rect 1313 933 1327 947
rect 1493 933 1507 947
rect 1553 933 1567 947
rect 2533 933 2547 947
rect 2633 933 2647 947
rect 4167 933 4181 947
rect 4213 933 4227 947
rect 4293 934 4307 948
rect 4393 933 4407 947
rect 5653 933 5667 947
rect 5693 934 5707 948
rect 1573 912 1587 926
rect 1613 913 1627 927
rect 1973 913 1987 927
rect 2013 913 2027 927
rect 4033 913 4047 927
rect 5093 913 5107 927
rect 5233 913 5247 927
rect 5453 913 5467 927
rect 5093 873 5107 887
rect 5193 873 5207 887
rect 5453 873 5467 887
rect 3273 853 3287 867
rect 3333 853 3347 867
rect 4073 853 4087 867
rect 1853 713 1867 727
rect 1893 713 1907 727
rect 2973 713 2987 727
rect 3053 713 3067 727
rect 3913 713 3927 727
rect 3973 713 3987 727
rect 4253 713 4267 727
rect 4333 713 4347 727
rect 4913 713 4927 727
rect 1273 693 1287 707
rect 1713 693 1727 707
rect 1313 653 1327 667
rect 2073 693 2087 707
rect 2233 693 2247 707
rect 2953 693 2967 707
rect 3013 693 3027 707
rect 3173 693 3187 707
rect 3153 673 3167 687
rect 3773 673 3787 687
rect 2013 653 2027 667
rect 2173 653 2187 667
rect 3133 653 3147 667
rect 3173 653 3187 667
rect 3713 653 3727 667
rect 3753 653 3767 667
rect 5833 693 5847 707
rect 4853 653 4867 667
rect 5793 653 5807 667
rect 1533 633 1547 647
rect 1673 633 1687 647
rect 1773 633 1787 647
rect 3773 633 3787 647
rect 3833 633 3847 647
rect 3953 633 3967 647
rect 453 413 467 427
rect 493 413 507 427
rect 2113 413 2127 427
rect 2273 413 2287 427
rect 2713 413 2727 427
rect 2793 413 2807 427
rect 2873 413 2887 427
rect 5853 413 5867 427
rect 5913 413 5927 427
rect 1593 393 1607 407
rect 2213 393 2227 407
rect 3213 393 3227 407
rect 3213 353 3227 367
rect 3273 393 3287 407
rect 873 333 887 347
rect 933 333 947 347
rect 1693 333 1707 347
rect 1793 333 1807 347
rect 2173 333 2187 347
rect 3233 332 3247 346
rect 3613 333 3627 347
rect 3673 331 3687 345
rect 2013 313 2027 327
rect 2053 313 2067 327
rect 1673 293 1687 307
rect 1753 293 1767 307
rect 1613 233 1627 247
rect 1673 233 1687 247
rect 2833 193 2847 207
rect 2913 193 2927 207
rect 1473 173 1487 187
rect 1533 173 1547 187
rect 2553 173 2567 187
rect 2953 173 2967 187
rect 4133 173 4147 187
rect 2093 133 2107 147
rect 2133 133 2147 147
rect 2513 133 2527 147
rect 4013 153 4027 167
rect 2993 133 3007 147
rect 3833 133 3847 147
rect 4453 173 4467 187
rect 573 113 587 127
rect 673 113 687 127
rect 993 113 1007 127
rect 1093 113 1107 127
rect 1152 113 1166 127
rect 1173 113 1187 127
rect 1253 113 1267 127
rect 2073 113 2087 127
rect 2193 113 2207 127
rect 4413 133 4427 147
rect 4213 113 4227 127
rect 5973 113 5987 127
rect 6073 113 6087 127
rect 1233 92 1247 106
rect 2793 33 2807 47
rect 2833 33 2847 47
<< metal2 >>
rect 3336 6267 3344 6304
rect 4856 6267 4864 6304
rect 96 6116 104 6153
rect 256 6116 264 6153
rect 296 6127 304 6213
rect 176 6084 184 6114
rect 396 6116 404 6153
rect 516 6128 524 6173
rect 316 6087 324 6114
rect 596 6087 604 6133
rect 656 6116 664 6213
rect 736 6124 744 6173
rect 756 6147 764 6193
rect 736 6116 764 6124
rect 793 6120 807 6133
rect 796 6116 804 6120
rect 116 5927 124 6084
rect 176 6076 204 6084
rect 113 5900 127 5913
rect 116 5896 124 5900
rect 196 5907 204 6076
rect 276 5908 284 6072
rect 376 5967 384 6084
rect 393 5908 407 5914
rect 96 5827 104 5864
rect 96 5627 104 5813
rect 16 5247 24 5374
rect 36 5046 44 5513
rect 96 5487 104 5564
rect 136 5527 144 5864
rect 176 5787 184 5864
rect 196 5827 204 5853
rect 156 5484 164 5713
rect 216 5667 224 5893
rect 256 5787 264 5864
rect 296 5707 304 5852
rect 336 5847 344 5894
rect 376 5827 384 5864
rect 187 5604 200 5607
rect 187 5596 204 5604
rect 187 5593 200 5596
rect 147 5476 164 5484
rect 56 5088 64 5433
rect 136 5388 144 5473
rect 96 5287 104 5344
rect 156 5340 164 5344
rect 153 5327 167 5340
rect 196 5327 204 5453
rect 216 5346 224 5393
rect 256 5376 264 5433
rect 276 5407 284 5653
rect 373 5600 387 5613
rect 396 5607 404 5833
rect 476 5827 484 6072
rect 536 6047 544 6084
rect 776 6047 784 6072
rect 856 6067 864 6133
rect 876 6107 884 6153
rect 916 6116 924 6213
rect 3536 6207 3544 6233
rect 1096 6116 1104 6153
rect 553 5900 567 5913
rect 556 5896 564 5900
rect 596 5896 604 5993
rect 636 5987 644 6033
rect 796 5987 804 6013
rect 856 6007 864 6053
rect 976 6027 984 6084
rect 1016 5987 1024 6114
rect 636 5976 653 5987
rect 640 5973 653 5976
rect 433 5608 447 5613
rect 376 5596 384 5600
rect 296 5567 304 5594
rect 476 5596 484 5713
rect 496 5624 504 5893
rect 616 5827 624 5852
rect 496 5620 524 5624
rect 496 5616 527 5620
rect 513 5607 527 5616
rect 296 5467 304 5553
rect 500 5564 513 5567
rect 396 5487 404 5553
rect 456 5487 464 5564
rect 496 5556 513 5564
rect 500 5553 513 5556
rect 536 5547 544 5594
rect 556 5567 564 5813
rect 296 5376 304 5413
rect 316 5287 324 5344
rect 96 5076 104 5133
rect 116 5040 124 5044
rect 113 5027 127 5040
rect 196 4884 204 5213
rect 336 5147 344 5273
rect 356 5227 364 5473
rect 416 5376 424 5413
rect 476 5344 484 5533
rect 556 5427 564 5532
rect 556 5376 564 5413
rect 576 5407 584 5633
rect 616 5624 624 5713
rect 636 5647 644 5953
rect 1076 5947 1084 6084
rect 1196 5987 1204 6153
rect 1376 6116 1384 6153
rect 1436 6086 1444 6193
rect 1656 6116 1664 6153
rect 1696 6116 1733 6124
rect 1776 6116 1784 6153
rect 1256 6080 1264 6084
rect 1253 6067 1267 6080
rect 716 5860 724 5864
rect 713 5847 727 5860
rect 776 5807 784 5864
rect 616 5616 644 5624
rect 636 5596 644 5616
rect 716 5567 724 5793
rect 816 5707 824 5893
rect 793 5624 807 5633
rect 776 5620 807 5624
rect 776 5616 804 5620
rect 776 5596 784 5616
rect 856 5587 864 5653
rect 656 5487 664 5564
rect 876 5527 884 5864
rect 916 5860 924 5864
rect 913 5847 927 5860
rect 936 5527 944 5564
rect 996 5447 1004 5933
rect 1156 5896 1204 5904
rect 1233 5900 1247 5913
rect 1236 5896 1244 5900
rect 1036 5860 1044 5864
rect 1033 5847 1047 5860
rect 1096 5687 1104 5864
rect 1036 5596 1044 5633
rect 1096 5596 1104 5673
rect 1136 5627 1144 5894
rect 1156 5687 1164 5896
rect 1336 5896 1344 6053
rect 1356 6007 1364 6084
rect 1396 6027 1404 6084
rect 1396 5947 1404 6013
rect 1356 5827 1364 5864
rect 1136 5567 1144 5613
rect 1156 5608 1164 5673
rect 1256 5667 1264 5813
rect 1233 5600 1247 5613
rect 1256 5607 1264 5653
rect 1236 5596 1244 5600
rect 616 5346 624 5393
rect 673 5380 687 5393
rect 676 5376 684 5380
rect 756 5346 764 5413
rect 836 5376 844 5413
rect 396 5307 404 5344
rect 276 4987 284 5044
rect 187 4876 204 4884
rect 96 4747 104 4824
rect 136 4820 144 4824
rect 133 4807 147 4820
rect 16 4324 24 4653
rect 76 4568 84 4593
rect 156 4568 164 4813
rect 176 4807 184 4873
rect 233 4860 247 4873
rect 236 4856 244 4860
rect 316 4826 324 4853
rect 176 4567 184 4793
rect 216 4747 224 4824
rect 256 4787 264 4824
rect 336 4804 344 5133
rect 356 5027 364 5093
rect 416 5076 424 5313
rect 436 5267 444 5344
rect 476 5336 504 5344
rect 456 5076 464 5133
rect 396 4907 404 5044
rect 436 4987 444 5044
rect 496 5007 504 5336
rect 536 5287 544 5344
rect 696 5307 704 5344
rect 516 5088 524 5193
rect 556 5147 564 5233
rect 696 5207 704 5293
rect 776 5167 784 5373
rect 816 5340 824 5344
rect 813 5327 827 5340
rect 856 5307 864 5344
rect 556 5076 564 5133
rect 673 5080 687 5093
rect 676 5076 684 5080
rect 516 4967 524 5074
rect 576 4967 584 5044
rect 416 4856 424 4953
rect 316 4796 344 4804
rect 36 4344 44 4554
rect 96 4467 104 4524
rect 36 4336 53 4344
rect 156 4347 164 4554
rect 196 4556 204 4733
rect 236 4556 244 4593
rect 136 4336 153 4344
rect 16 4316 44 4324
rect 16 3627 24 3933
rect 16 2687 24 3613
rect 36 3447 44 4316
rect 56 4007 64 4334
rect 176 4307 184 4473
rect 236 4336 244 4373
rect 256 4367 264 4524
rect 296 4487 304 4553
rect 316 4527 324 4796
rect 336 4727 344 4773
rect 296 4367 304 4473
rect 336 4347 344 4713
rect 396 4588 404 4812
rect 476 4687 484 4854
rect 496 4627 504 4893
rect 553 4860 567 4873
rect 556 4856 564 4860
rect 536 4747 544 4824
rect 416 4467 424 4524
rect 116 4036 124 4073
rect 256 4067 264 4304
rect 316 4087 324 4334
rect 376 4336 384 4373
rect 420 4344 433 4347
rect 416 4336 433 4344
rect 420 4333 433 4336
rect 396 4300 404 4304
rect 393 4287 407 4300
rect 436 4244 444 4293
rect 456 4267 464 4353
rect 476 4344 484 4573
rect 556 4568 564 4793
rect 576 4727 584 4824
rect 616 4547 624 4673
rect 536 4467 544 4512
rect 576 4467 584 4524
rect 636 4507 644 4993
rect 656 4827 664 5044
rect 696 5040 704 5044
rect 693 5027 707 5040
rect 756 4967 764 5074
rect 776 5027 784 5153
rect 916 5104 924 5413
rect 1076 5407 1084 5552
rect 1156 5547 1164 5594
rect 936 5247 944 5374
rect 1036 5307 1044 5344
rect 1076 5307 1084 5372
rect 976 5167 984 5293
rect 1096 5207 1104 5533
rect 1116 5327 1124 5433
rect 1176 5376 1184 5413
rect 1276 5388 1284 5773
rect 1376 5604 1384 5833
rect 1356 5596 1384 5604
rect 1336 5527 1344 5564
rect 1396 5527 1404 5894
rect 1416 5867 1424 5973
rect 1496 5896 1504 6033
rect 1536 5787 1544 6084
rect 1576 6007 1584 6114
rect 1636 5947 1644 6084
rect 1716 5896 1724 6072
rect 1736 6027 1744 6114
rect 1836 6047 1844 6084
rect 1876 5967 1884 6153
rect 1996 6116 2004 6193
rect 1916 6086 1924 6114
rect 1976 6080 1984 6084
rect 1556 5827 1564 5894
rect 1736 5856 1764 5864
rect 1556 5724 1564 5813
rect 1536 5716 1564 5724
rect 1536 5567 1544 5716
rect 1613 5600 1627 5613
rect 1616 5596 1624 5600
rect 1736 5596 1744 5733
rect 1756 5727 1764 5856
rect 1776 5687 1784 5953
rect 1796 5747 1804 5853
rect 1876 5827 1884 5894
rect 1896 5724 1904 5933
rect 1916 5787 1924 6072
rect 1973 6067 1987 6080
rect 2036 6067 2044 6173
rect 2076 6116 2084 6193
rect 2236 6116 2244 6193
rect 2256 6147 2264 6173
rect 2256 6137 2273 6147
rect 2260 6134 2273 6137
rect 2260 6133 2280 6134
rect 2176 6087 2184 6114
rect 2333 6120 2347 6133
rect 2336 6116 2344 6120
rect 2376 6116 2384 6173
rect 1956 5896 1964 6013
rect 2056 5847 2064 5993
rect 2136 5967 2144 6084
rect 2113 5924 2127 5933
rect 2113 5920 2133 5924
rect 2116 5916 2133 5920
rect 2136 5896 2144 5913
rect 2193 5904 2207 5913
rect 2193 5900 2224 5904
rect 2196 5896 2224 5900
rect 2396 5904 2404 6084
rect 2396 5896 2424 5904
rect 2236 5747 2244 5864
rect 2276 5827 2284 5864
rect 2416 5727 2424 5896
rect 1896 5716 1913 5724
rect 1456 5507 1464 5564
rect 1496 5527 1504 5564
rect 1656 5566 1664 5593
rect 1633 5507 1647 5513
rect 1456 5467 1464 5493
rect 1696 5487 1704 5513
rect 1713 5507 1727 5513
rect 1156 5340 1164 5344
rect 1136 5247 1144 5333
rect 1153 5327 1167 5340
rect 1156 5287 1164 5313
rect 1256 5287 1264 5344
rect 1296 5307 1304 5344
rect 916 5096 944 5104
rect 936 5076 944 5096
rect 976 5076 984 5153
rect 1096 5088 1104 5153
rect 1016 5076 1064 5084
rect 876 5027 884 5073
rect 693 4860 707 4873
rect 696 4856 704 4860
rect 716 4787 724 4824
rect 736 4587 744 4733
rect 756 4727 764 4824
rect 776 4667 784 4693
rect 476 4336 504 4344
rect 436 4236 464 4244
rect 193 4048 207 4053
rect 273 4040 287 4053
rect 276 4036 284 4040
rect 136 4000 144 4004
rect 133 3987 147 4000
rect 56 3786 64 3833
rect 116 3816 124 3913
rect 156 3816 164 3893
rect 196 3827 204 4034
rect 396 4036 404 4073
rect 136 3547 144 3784
rect 176 3747 184 3784
rect 56 3485 64 3533
rect 196 3516 204 3593
rect 216 3524 224 3993
rect 256 3987 264 4004
rect 256 3847 264 3973
rect 276 3816 284 3893
rect 296 3827 304 4004
rect 336 3927 344 4033
rect 456 4007 464 4236
rect 376 3887 384 4004
rect 416 3947 424 4004
rect 476 3967 484 4293
rect 496 4087 504 4273
rect 516 4267 524 4304
rect 556 4300 564 4304
rect 553 4287 567 4300
rect 596 4247 604 4493
rect 656 4407 664 4513
rect 616 4287 624 4393
rect 736 4367 744 4524
rect 776 4504 784 4553
rect 796 4527 804 4953
rect 816 4827 824 4953
rect 876 4884 884 5013
rect 916 4987 924 5044
rect 956 4967 964 5044
rect 876 4876 904 4884
rect 896 4856 904 4876
rect 996 4856 1004 5013
rect 1016 4947 1024 5076
rect 1156 5047 1164 5113
rect 1076 4987 1084 5044
rect 1016 4887 1024 4933
rect 1036 4856 1084 4864
rect 816 4567 824 4813
rect 916 4820 924 4824
rect 913 4807 927 4820
rect 1013 4807 1027 4812
rect 876 4647 884 4773
rect 756 4496 784 4504
rect 656 4207 664 4304
rect 696 4147 704 4293
rect 716 4247 724 4304
rect 756 4247 764 4496
rect 816 4487 824 4513
rect 776 4287 784 4453
rect 856 4387 864 4473
rect 976 4427 984 4613
rect 1036 4567 1044 4593
rect 1056 4584 1064 4713
rect 1076 4607 1084 4856
rect 1116 4867 1124 5044
rect 1176 4987 1184 5193
rect 1236 5076 1244 5233
rect 1356 5127 1364 5453
rect 1473 5444 1487 5453
rect 1456 5440 1487 5444
rect 1456 5436 1484 5440
rect 1456 5376 1464 5436
rect 1396 5187 1404 5373
rect 1556 5347 1564 5373
rect 1696 5344 1704 5473
rect 1756 5427 1764 5564
rect 1796 5427 1804 5613
rect 1916 5567 1924 5713
rect 1936 5608 1944 5693
rect 1936 5507 1944 5594
rect 1956 5547 1964 5613
rect 1996 5596 2004 5673
rect 2436 5667 2444 5953
rect 2456 5907 2464 6114
rect 2476 6084 2484 6173
rect 2667 6144 2680 6147
rect 2667 6133 2684 6144
rect 2533 6120 2547 6133
rect 2536 6116 2544 6120
rect 2676 6116 2684 6133
rect 2776 6128 2784 6153
rect 2856 6116 2864 6153
rect 2476 6076 2504 6084
rect 2496 5896 2504 6076
rect 2556 5947 2564 6084
rect 2776 6084 2784 6114
rect 3096 6116 3104 6173
rect 3196 6116 3204 6193
rect 3036 6086 3044 6113
rect 2776 6076 2804 6084
rect 2716 6047 2724 6072
rect 2636 5896 2644 5933
rect 2516 5827 2524 5864
rect 2576 5847 2584 5894
rect 2756 5896 2764 6033
rect 2796 5927 2804 6076
rect 2836 5947 2844 6084
rect 2793 5900 2807 5913
rect 2796 5896 2804 5900
rect 2653 5847 2667 5852
rect 2213 5608 2227 5613
rect 1907 5493 1913 5507
rect 1976 5467 1984 5493
rect 1796 5376 1804 5413
rect 1956 5376 1964 5453
rect 2016 5447 2024 5564
rect 1476 5267 1484 5324
rect 1207 5044 1220 5047
rect 1207 5036 1224 5044
rect 1256 5040 1264 5044
rect 1207 5033 1220 5036
rect 1253 5027 1267 5040
rect 1296 5027 1304 5093
rect 1333 5080 1347 5093
rect 1336 5076 1344 5080
rect 1376 5076 1384 5153
rect 1456 5088 1464 5153
rect 1396 5040 1404 5044
rect 1096 4767 1104 4854
rect 1196 4707 1204 4853
rect 1216 4667 1224 5013
rect 1276 4856 1284 4933
rect 1316 4867 1324 4913
rect 1256 4787 1264 4824
rect 1296 4707 1304 4824
rect 1336 4807 1344 5013
rect 1356 4868 1364 5032
rect 1393 5027 1407 5040
rect 1456 4947 1464 5074
rect 1476 5027 1484 5093
rect 1356 4747 1364 4854
rect 1396 4787 1404 4824
rect 1456 4807 1464 4824
rect 1396 4727 1404 4773
rect 1056 4576 1084 4584
rect 1076 4556 1084 4576
rect 996 4407 1004 4533
rect 873 4380 887 4393
rect 876 4376 884 4380
rect 496 3947 504 4034
rect 513 3987 527 3993
rect 413 3820 427 3833
rect 416 3816 424 3820
rect 316 3747 324 3784
rect 216 3516 233 3524
rect 76 3308 84 3473
rect 156 3476 184 3484
rect 116 3296 124 3393
rect 156 3307 164 3453
rect 36 2966 44 3293
rect 96 2996 104 3252
rect 136 3227 144 3264
rect 176 3224 184 3476
rect 236 3467 244 3513
rect 196 3244 204 3313
rect 233 3300 247 3313
rect 276 3308 284 3573
rect 336 3516 344 3613
rect 356 3587 364 3813
rect 516 3786 524 3873
rect 596 3847 604 4004
rect 376 3516 384 3753
rect 436 3627 444 3784
rect 596 3727 604 3784
rect 616 3547 624 3773
rect 493 3528 507 3533
rect 533 3520 547 3533
rect 593 3520 607 3533
rect 636 3528 644 3833
rect 656 3827 664 4004
rect 696 4000 724 4004
rect 696 3996 727 4000
rect 713 3987 727 3996
rect 727 3976 744 3984
rect 676 3927 684 3953
rect 696 3816 704 3933
rect 736 3827 744 3976
rect 756 3924 764 4073
rect 776 4036 784 4193
rect 796 4187 804 4353
rect 856 4336 864 4373
rect 956 4307 964 4393
rect 996 4336 1004 4393
rect 1036 4336 1044 4513
rect 1056 4487 1064 4524
rect 1136 4427 1144 4573
rect 1156 4467 1164 4633
rect 1213 4560 1227 4573
rect 1216 4556 1224 4560
rect 1296 4567 1304 4653
rect 1356 4556 1364 4712
rect 1396 4556 1404 4633
rect 1316 4527 1324 4554
rect 1456 4527 1464 4793
rect 1496 4687 1504 5233
rect 1536 5107 1544 5193
rect 1533 5080 1547 5093
rect 1536 5076 1544 5080
rect 1576 5076 1584 5253
rect 1616 5167 1624 5344
rect 1656 5247 1664 5344
rect 1676 5336 1704 5344
rect 1556 5027 1564 5044
rect 1556 4907 1564 5013
rect 1576 4884 1584 4993
rect 1596 4987 1604 5032
rect 1656 4927 1664 5074
rect 1676 5007 1684 5336
rect 1776 5267 1784 5344
rect 1756 5088 1764 5113
rect 1707 5084 1720 5087
rect 1707 5076 1724 5084
rect 1707 5073 1720 5076
rect 1696 4907 1704 5033
rect 1556 4876 1584 4884
rect 1556 4856 1564 4876
rect 1596 4767 1604 4853
rect 1716 4827 1724 4933
rect 1636 4787 1644 4824
rect 1556 4568 1564 4753
rect 1676 4687 1684 4824
rect 1176 4447 1184 4512
rect 1096 4306 1104 4353
rect 896 4047 904 4133
rect 816 3947 824 4004
rect 756 3916 784 3924
rect 756 3786 764 3893
rect 776 3827 784 3916
rect 836 3887 844 3964
rect 813 3820 827 3833
rect 856 3827 864 3913
rect 816 3816 824 3820
rect 676 3727 684 3772
rect 536 3516 544 3520
rect 596 3516 604 3520
rect 676 3527 684 3553
rect 436 3487 444 3514
rect 476 3364 484 3484
rect 616 3464 624 3484
rect 656 3480 664 3484
rect 653 3467 667 3480
rect 616 3456 644 3464
rect 636 3444 644 3456
rect 676 3444 684 3473
rect 636 3436 684 3444
rect 456 3356 484 3364
rect 376 3308 384 3353
rect 236 3296 244 3300
rect 416 3296 424 3333
rect 456 3287 464 3356
rect 196 3236 224 3244
rect 176 3216 193 3224
rect 176 3008 184 3113
rect 136 2776 144 2893
rect 176 2827 184 2994
rect 56 2607 64 2773
rect 116 2740 124 2744
rect 113 2727 127 2740
rect 196 2744 204 3213
rect 216 3008 224 3236
rect 256 3227 264 3264
rect 273 3008 287 3013
rect 316 2996 324 3153
rect 396 3127 404 3252
rect 456 3247 464 3273
rect 476 3187 484 3333
rect 536 3296 544 3353
rect 596 3307 604 3433
rect 696 3427 704 3653
rect 756 3544 764 3593
rect 776 3567 784 3773
rect 836 3747 844 3784
rect 756 3536 784 3544
rect 776 3516 784 3536
rect 836 3487 844 3514
rect 516 3260 524 3264
rect 513 3247 527 3260
rect 616 3266 624 3333
rect 596 3227 604 3253
rect 636 3264 644 3413
rect 716 3347 724 3413
rect 756 3407 764 3484
rect 856 3467 864 3773
rect 876 3667 884 3933
rect 896 3827 904 3853
rect 916 3827 924 4173
rect 936 3844 944 4273
rect 1076 4107 1084 4233
rect 1116 4187 1124 4413
rect 1236 4407 1244 4473
rect 1276 4407 1284 4524
rect 1316 4447 1324 4513
rect 1336 4447 1344 4513
rect 1413 4504 1427 4513
rect 1396 4500 1427 4504
rect 1396 4496 1424 4500
rect 1167 4356 1193 4364
rect 1136 4296 1164 4304
rect 1136 4227 1144 4296
rect 1136 4164 1144 4213
rect 1116 4156 1144 4164
rect 1096 4027 1104 4133
rect 936 3836 964 3844
rect 956 3828 964 3836
rect 996 3816 1004 3933
rect 1116 3907 1124 4156
rect 1156 4036 1164 4253
rect 1196 4207 1204 4304
rect 1216 4147 1224 4293
rect 1236 4247 1244 4393
rect 1333 4340 1347 4353
rect 1336 4336 1344 4340
rect 1396 4327 1404 4496
rect 1476 4487 1484 4513
rect 1496 4464 1504 4524
rect 1467 4456 1504 4464
rect 1416 4327 1424 4433
rect 1576 4327 1584 4373
rect 1276 4204 1284 4313
rect 1316 4300 1324 4304
rect 1356 4300 1364 4304
rect 1313 4287 1327 4300
rect 1353 4287 1367 4300
rect 1556 4300 1564 4305
rect 1276 4196 1293 4204
rect 1176 3984 1184 4004
rect 1156 3976 1184 3984
rect 896 3786 904 3813
rect 976 3780 984 3784
rect 973 3767 987 3780
rect 896 3644 904 3713
rect 876 3636 904 3644
rect 876 3447 884 3636
rect 916 3528 924 3753
rect 1036 3727 1044 3893
rect 1156 3867 1164 3976
rect 1067 3784 1080 3787
rect 1067 3776 1084 3784
rect 1067 3773 1080 3776
rect 1116 3767 1124 3784
rect 1176 3767 1184 3893
rect 956 3567 964 3593
rect 956 3516 964 3553
rect 996 3527 1004 3673
rect 896 3427 904 3473
rect 976 3480 984 3484
rect 973 3467 987 3480
rect 756 3367 764 3393
rect 667 3304 680 3307
rect 667 3296 684 3304
rect 667 3293 680 3296
rect 756 3307 764 3353
rect 856 3296 864 3393
rect 896 3307 904 3413
rect 636 3256 664 3264
rect 256 2867 264 2964
rect 216 2787 224 2853
rect 276 2804 284 2893
rect 256 2796 284 2804
rect 256 2776 264 2796
rect 176 2736 204 2744
rect 16 247 24 2573
rect 36 2387 44 2513
rect 156 2487 164 2673
rect 36 2107 44 2253
rect 36 1207 44 1853
rect 56 1807 64 2413
rect 96 2387 104 2444
rect 116 2347 124 2433
rect 176 2427 184 2736
rect 216 2527 224 2633
rect 276 2567 284 2744
rect 216 2476 224 2513
rect 256 2488 264 2533
rect 193 2427 207 2433
rect 76 2267 84 2333
rect 116 2256 124 2293
rect 76 2087 84 2193
rect 96 2027 104 2191
rect 136 2127 144 2224
rect 196 2224 204 2333
rect 236 2268 244 2444
rect 296 2387 304 2673
rect 256 2307 264 2373
rect 260 2284 273 2287
rect 256 2273 273 2284
rect 216 2260 233 2264
rect 213 2256 233 2260
rect 213 2247 227 2256
rect 256 2256 264 2273
rect 296 2256 304 2333
rect 316 2287 324 2713
rect 336 2687 344 2813
rect 356 2727 364 3013
rect 393 3000 407 3013
rect 396 2996 404 3000
rect 436 2996 444 3153
rect 496 2967 504 3053
rect 593 3000 607 3013
rect 636 3007 644 3233
rect 596 2996 604 3000
rect 396 2776 404 2873
rect 516 2867 524 2994
rect 576 2907 584 2952
rect 616 2927 624 2964
rect 496 2746 504 2813
rect 556 2788 564 2833
rect 456 2736 493 2744
rect 536 2740 544 2744
rect 413 2727 427 2732
rect 533 2727 547 2740
rect 516 2607 524 2693
rect 636 2567 644 2933
rect 656 2627 664 3256
rect 740 3264 753 3267
rect 736 3256 753 3264
rect 740 3253 753 3256
rect 716 3187 724 3233
rect 776 3167 784 3294
rect 836 3260 844 3264
rect 833 3247 847 3260
rect 916 3207 924 3433
rect 1016 3407 1024 3553
rect 1076 3516 1084 3593
rect 1116 3567 1124 3753
rect 1116 3516 1124 3553
rect 1036 3480 1064 3484
rect 1033 3476 1064 3480
rect 1033 3467 1047 3476
rect 1096 3447 1104 3484
rect 1156 3407 1164 3713
rect 996 3296 1004 3353
rect 1036 3296 1044 3353
rect 1116 3327 1124 3353
rect 1156 3327 1164 3353
rect 1156 3296 1164 3313
rect 1176 3307 1184 3593
rect 1196 3567 1204 3933
rect 1216 3786 1224 4004
rect 1256 3967 1264 4093
rect 1236 3827 1244 3933
rect 1276 3907 1284 4034
rect 1296 4007 1304 4193
rect 1336 4067 1344 4173
rect 1436 4107 1444 4292
rect 1553 4287 1567 4300
rect 1336 4036 1344 4053
rect 1376 4036 1384 4093
rect 1276 3816 1284 3853
rect 1356 3827 1364 4004
rect 1396 3844 1404 3953
rect 1416 3947 1424 4033
rect 1436 3887 1444 4053
rect 1476 4048 1484 4233
rect 1596 4227 1604 4633
rect 1616 4227 1624 4673
rect 1736 4667 1744 4953
rect 1716 4568 1724 4613
rect 1656 4427 1664 4524
rect 1696 4520 1704 4524
rect 1693 4507 1707 4520
rect 1693 4487 1707 4493
rect 1676 4336 1684 4393
rect 1536 4036 1544 4153
rect 1396 3836 1424 3844
rect 1416 3816 1424 3836
rect 1456 3816 1464 3953
rect 1496 3847 1504 3992
rect 1236 3607 1244 3773
rect 1256 3647 1264 3772
rect 1336 3567 1344 3773
rect 1356 3747 1364 3792
rect 1376 3587 1384 3773
rect 1396 3747 1404 3784
rect 1256 3528 1264 3553
rect 1296 3516 1304 3553
rect 1496 3524 1504 3812
rect 1516 3786 1524 3853
rect 1536 3747 1544 3873
rect 1556 3827 1564 3993
rect 1576 3967 1584 4173
rect 1596 4047 1604 4192
rect 1636 4104 1644 4293
rect 1656 4127 1664 4304
rect 1636 4096 1664 4104
rect 1656 4047 1664 4096
rect 1676 4004 1684 4253
rect 1696 4247 1704 4304
rect 1716 4224 1724 4293
rect 1736 4267 1744 4493
rect 1756 4487 1764 4993
rect 1776 4987 1784 5033
rect 1796 5027 1804 5313
rect 1816 5307 1824 5344
rect 1876 5327 1884 5374
rect 1936 5307 1944 5344
rect 1976 5340 1984 5344
rect 1973 5327 1987 5340
rect 1816 5087 1824 5293
rect 1936 5247 1944 5293
rect 2016 5267 2024 5374
rect 2076 5327 2084 5344
rect 2067 5316 2084 5327
rect 2067 5313 2080 5316
rect 1916 5207 1924 5233
rect 1876 5076 1884 5193
rect 2016 5076 2024 5213
rect 1856 5040 1864 5044
rect 1853 5027 1867 5040
rect 1816 4868 1824 4893
rect 1796 4744 1804 4824
rect 1896 4784 1904 5033
rect 1916 5027 1924 5074
rect 2056 5047 2064 5253
rect 2076 5227 2084 5293
rect 2116 5267 2124 5533
rect 2136 5187 2144 5493
rect 2156 5307 2164 5513
rect 2196 5507 2204 5564
rect 2236 5527 2244 5613
rect 2256 5567 2264 5613
rect 2293 5600 2307 5613
rect 2296 5596 2304 5600
rect 2316 5560 2324 5564
rect 2276 5527 2284 5553
rect 2313 5547 2327 5560
rect 2356 5527 2364 5564
rect 2396 5547 2404 5613
rect 2493 5600 2507 5613
rect 2496 5596 2504 5600
rect 2216 5376 2224 5433
rect 2256 5376 2264 5493
rect 2316 5467 2324 5512
rect 2276 5387 2284 5413
rect 2316 5388 2324 5453
rect 2396 5444 2404 5493
rect 2436 5487 2444 5564
rect 2396 5436 2424 5444
rect 2356 5376 2364 5413
rect 2416 5347 2424 5436
rect 2476 5404 2484 5564
rect 2536 5407 2544 5594
rect 2476 5396 2504 5404
rect 2496 5388 2504 5396
rect 2556 5384 2564 5613
rect 2596 5596 2604 5633
rect 2616 5507 2624 5564
rect 2536 5376 2584 5384
rect 2196 5247 2204 5344
rect 2236 5267 2244 5344
rect 1956 4856 1964 5013
rect 1976 4987 1984 5044
rect 1936 4820 1944 4824
rect 1887 4776 1904 4784
rect 1796 4736 1824 4744
rect 1796 4556 1804 4713
rect 1816 4707 1824 4736
rect 1876 4567 1884 4773
rect 1916 4627 1924 4812
rect 1933 4807 1947 4820
rect 1987 4816 2004 4824
rect 1936 4687 1944 4793
rect 1996 4787 2004 4816
rect 1896 4527 1904 4613
rect 1996 4556 2004 4733
rect 1773 4507 1787 4513
rect 1856 4487 1864 4524
rect 1816 4336 1824 4373
rect 1856 4336 1864 4413
rect 1876 4347 1884 4393
rect 1596 3947 1604 3993
rect 1616 3984 1624 4004
rect 1656 3996 1684 4004
rect 1696 4216 1724 4224
rect 1616 3976 1644 3984
rect 1596 3816 1604 3893
rect 1616 3847 1624 3953
rect 1636 3907 1644 3976
rect 1636 3827 1644 3853
rect 1476 3516 1504 3524
rect 1536 3516 1544 3673
rect 1556 3607 1564 3773
rect 1616 3707 1624 3784
rect 1553 3567 1567 3572
rect 1576 3528 1584 3553
rect 1236 3384 1244 3484
rect 1276 3447 1284 3484
rect 1376 3424 1384 3484
rect 1416 3447 1424 3484
rect 1456 3447 1464 3473
rect 1376 3416 1404 3424
rect 1236 3376 1264 3384
rect 713 3000 727 3013
rect 716 2996 724 3000
rect 756 2996 764 3053
rect 796 3007 804 3073
rect 676 2927 684 2993
rect 780 2964 793 2967
rect 736 2847 744 2964
rect 776 2956 793 2964
rect 780 2953 793 2956
rect 816 2947 824 2994
rect 773 2780 787 2793
rect 776 2776 784 2780
rect 676 2667 684 2773
rect 716 2587 724 2744
rect 816 2627 824 2873
rect 836 2787 844 3193
rect 1016 3127 1024 3264
rect 1056 3227 1064 3264
rect 1196 3260 1204 3264
rect 1193 3247 1207 3260
rect 1236 3264 1244 3353
rect 1256 3347 1264 3376
rect 1236 3256 1284 3264
rect 1193 3227 1207 3233
rect 916 2996 924 3033
rect 956 3007 964 3113
rect 1016 2996 1024 3073
rect 1060 3004 1073 3007
rect 1056 2996 1073 3004
rect 1060 2993 1073 2996
rect 1096 2967 1104 3013
rect 1216 3004 1224 3253
rect 1287 3233 1293 3247
rect 1216 2996 1244 3004
rect 853 2947 867 2953
rect 896 2887 904 2964
rect 976 2956 1004 2964
rect 853 2780 867 2793
rect 856 2776 864 2780
rect 896 2776 904 2873
rect 976 2827 984 2956
rect 1076 2927 1084 2953
rect 976 2787 984 2813
rect 876 2740 884 2744
rect 396 2476 404 2513
rect 376 2424 384 2444
rect 416 2440 424 2444
rect 356 2416 384 2424
rect 413 2427 427 2440
rect 356 2347 364 2416
rect 196 2216 224 2224
rect 176 1967 184 2213
rect 216 2147 224 2216
rect 236 2187 244 2212
rect 276 2127 284 2224
rect 156 1956 173 1964
rect 96 1867 104 1924
rect 116 1847 124 1893
rect 136 1867 144 1924
rect 176 1747 184 1913
rect 196 1907 204 2113
rect 296 2067 304 2193
rect 296 1968 304 2013
rect 36 1107 44 1172
rect 36 727 44 1013
rect 56 1007 64 1733
rect 196 1706 204 1893
rect 216 1747 224 1913
rect 236 1807 244 1924
rect 276 1847 284 1924
rect 256 1736 264 1773
rect 316 1767 324 1913
rect 336 1867 344 2173
rect 356 1967 364 2273
rect 376 2226 384 2293
rect 396 2267 404 2333
rect 456 2287 464 2473
rect 476 2444 484 2553
rect 476 2436 504 2444
rect 476 2256 484 2373
rect 496 2267 504 2436
rect 536 2387 544 2444
rect 576 2347 584 2453
rect 616 2387 624 2444
rect 656 2427 664 2444
rect 656 2416 673 2427
rect 660 2413 673 2416
rect 516 2226 524 2273
rect 576 2256 584 2333
rect 393 1960 407 1973
rect 436 1968 444 2193
rect 456 2167 464 2224
rect 536 2027 544 2213
rect 596 2187 604 2224
rect 596 2127 604 2173
rect 396 1956 404 1960
rect 493 1960 507 1973
rect 496 1956 504 1960
rect 596 1926 604 2053
rect 376 1920 384 1924
rect 96 1587 104 1704
rect 227 1704 240 1707
rect 227 1696 244 1704
rect 227 1693 240 1696
rect 336 1567 344 1733
rect 116 1436 124 1513
rect 156 1436 164 1553
rect 216 1436 224 1513
rect 256 1436 264 1493
rect 96 1247 104 1404
rect 136 1367 144 1404
rect 116 1216 124 1313
rect 276 1267 284 1404
rect 316 1367 324 1493
rect 336 1406 344 1553
rect 196 1186 204 1253
rect 76 947 84 1173
rect 316 1184 324 1332
rect 356 1327 364 1913
rect 373 1907 387 1920
rect 556 1887 564 1924
rect 387 1744 400 1747
rect 387 1736 404 1744
rect 436 1736 444 1833
rect 556 1767 564 1873
rect 387 1733 400 1736
rect 496 1706 504 1753
rect 376 1647 384 1693
rect 396 1436 404 1593
rect 416 1587 424 1692
rect 436 1527 444 1673
rect 416 1228 424 1404
rect 476 1347 484 1553
rect 556 1467 564 1704
rect 596 1607 604 1693
rect 556 1436 564 1453
rect 616 1407 624 2013
rect 633 1967 647 1973
rect 656 1968 664 2253
rect 676 1987 684 2273
rect 696 2267 704 2433
rect 716 2427 724 2552
rect 716 2256 724 2373
rect 736 2367 744 2613
rect 836 2567 844 2733
rect 873 2727 887 2740
rect 916 2707 924 2744
rect 956 2727 964 2773
rect 973 2727 987 2733
rect 916 2687 924 2693
rect 916 2676 933 2687
rect 920 2673 933 2676
rect 987 2673 993 2687
rect 756 2407 764 2513
rect 816 2476 824 2513
rect 796 2367 804 2444
rect 836 2307 844 2444
rect 753 2260 767 2273
rect 756 2256 764 2260
rect 836 2227 844 2272
rect 696 2187 704 2213
rect 736 2187 744 2224
rect 776 2147 784 2212
rect 856 2187 864 2393
rect 876 2287 884 2593
rect 896 2407 904 2533
rect 936 2476 944 2513
rect 976 2476 984 2553
rect 1036 2487 1044 2533
rect 1056 2488 1064 2833
rect 1076 2687 1084 2913
rect 1096 2787 1104 2932
rect 1156 2887 1164 2964
rect 1236 2904 1244 2996
rect 1216 2896 1244 2904
rect 1136 2776 1144 2873
rect 1173 2780 1187 2793
rect 1176 2776 1184 2780
rect 1116 2547 1124 2732
rect 1156 2687 1164 2744
rect 1173 2527 1187 2533
rect 956 2347 964 2444
rect 1016 2427 1024 2474
rect 1096 2476 1104 2513
rect 916 2256 924 2333
rect 787 2024 800 2027
rect 787 2020 804 2024
rect 787 2013 807 2020
rect 646 1960 647 1967
rect 696 1956 704 2013
rect 793 2007 807 2013
rect 876 1987 884 2213
rect 636 1747 644 1913
rect 716 1847 724 1924
rect 716 1736 724 1793
rect 756 1748 764 1953
rect 776 1887 784 1973
rect 896 1967 904 2033
rect 916 1927 924 1993
rect 796 1767 804 1913
rect 836 1887 844 1924
rect 856 1827 864 1893
rect 876 1706 884 1753
rect 696 1647 704 1704
rect 796 1700 804 1704
rect 793 1687 807 1700
rect 636 1476 713 1484
rect 636 1448 644 1476
rect 653 1440 667 1453
rect 693 1440 707 1453
rect 656 1436 664 1440
rect 696 1436 704 1440
rect 496 1216 504 1293
rect 536 1287 544 1404
rect 276 1176 324 1184
rect 96 1067 104 1172
rect 56 936 73 944
rect 56 867 64 936
rect 113 920 127 933
rect 116 916 124 920
rect 156 916 164 993
rect 196 927 204 1172
rect 253 947 267 953
rect 213 920 227 933
rect 216 916 224 920
rect 256 916 264 933
rect 36 627 44 713
rect 56 666 64 753
rect 96 727 104 884
rect 136 880 144 884
rect 133 867 147 880
rect 316 886 324 993
rect 116 696 124 733
rect 176 708 184 873
rect 276 787 284 884
rect 156 696 173 704
rect 136 627 144 664
rect 116 396 124 473
rect 153 400 167 413
rect 196 407 204 733
rect 276 724 284 773
rect 276 716 304 724
rect 216 696 264 704
rect 296 696 304 716
rect 336 704 344 1213
rect 396 1147 404 1184
rect 436 1087 444 1184
rect 396 947 404 1053
rect 416 916 424 1013
rect 476 886 484 1173
rect 516 916 524 1172
rect 556 1147 564 1233
rect 576 1167 584 1393
rect 676 1384 684 1404
rect 656 1376 684 1384
rect 636 1216 644 1253
rect 656 1247 664 1376
rect 693 1367 707 1373
rect 716 1367 724 1404
rect 687 1360 707 1367
rect 687 1356 704 1360
rect 687 1353 700 1356
rect 676 1216 684 1332
rect 756 1287 764 1673
rect 836 1567 844 1704
rect 816 1436 824 1473
rect 876 1406 884 1453
rect 796 1367 804 1404
rect 896 1384 904 1913
rect 916 1487 924 1793
rect 936 1747 944 2213
rect 956 1968 964 2312
rect 976 2227 984 2413
rect 1036 2327 1044 2433
rect 1056 2268 1064 2413
rect 1076 2367 1084 2444
rect 1136 2407 1144 2513
rect 1193 2480 1207 2493
rect 1216 2487 1224 2896
rect 1236 2487 1244 2873
rect 1256 2847 1264 3193
rect 1356 3167 1364 3293
rect 1376 3144 1384 3393
rect 1356 3136 1384 3144
rect 1296 2927 1304 2964
rect 1336 2887 1344 2953
rect 1356 2944 1364 3136
rect 1376 2967 1384 3053
rect 1356 2936 1384 2944
rect 1336 2776 1344 2813
rect 1276 2627 1284 2744
rect 1316 2607 1324 2744
rect 1376 2567 1384 2936
rect 1396 2927 1404 3416
rect 1476 3407 1484 3516
rect 1516 3307 1524 3484
rect 1616 3387 1624 3593
rect 1636 3527 1644 3773
rect 1656 3667 1664 3996
rect 1696 3907 1704 4216
rect 1676 3896 1693 3904
rect 1676 3827 1684 3896
rect 1696 3816 1704 3853
rect 1716 3847 1724 4093
rect 1736 4067 1744 4232
rect 1796 4087 1804 4304
rect 1896 4247 1904 4492
rect 1916 4068 1924 4473
rect 1976 4427 1984 4524
rect 1996 4367 2004 4493
rect 2036 4484 2044 4993
rect 2076 4907 2084 5173
rect 2116 5076 2124 5113
rect 2156 5088 2164 5193
rect 2136 4987 2144 5044
rect 2196 5007 2204 5173
rect 2276 5076 2284 5273
rect 2296 5247 2304 5333
rect 2256 4987 2264 5044
rect 2296 4967 2304 5033
rect 2093 4860 2107 4873
rect 2096 4856 2104 4860
rect 2116 4727 2124 4773
rect 2136 4767 2144 4873
rect 2096 4556 2104 4693
rect 2156 4587 2164 4893
rect 2316 4884 2324 5313
rect 2336 5307 2344 5344
rect 2376 5340 2384 5344
rect 2373 5327 2387 5340
rect 2336 5067 2344 5233
rect 2336 4887 2344 5053
rect 2356 5027 2364 5093
rect 2393 5080 2407 5093
rect 2436 5087 2444 5293
rect 2396 5076 2404 5080
rect 2456 5046 2464 5333
rect 2476 5287 2484 5344
rect 2516 5327 2524 5344
rect 2516 5167 2524 5313
rect 2576 5307 2584 5376
rect 2556 5267 2564 5293
rect 2576 5127 2584 5253
rect 2596 5187 2604 5413
rect 2613 5387 2627 5393
rect 2656 5376 2664 5453
rect 2676 5407 2684 5553
rect 2696 5387 2704 5653
rect 2716 5427 2724 5893
rect 2856 5807 2864 5913
rect 2896 5896 2904 5933
rect 2976 5927 2984 6084
rect 2976 5867 2984 5913
rect 2996 5887 3004 6033
rect 3116 5984 3124 6084
rect 3227 6076 3244 6084
rect 3096 5976 3124 5984
rect 2736 5607 2744 5793
rect 2756 5596 2764 5633
rect 2796 5376 2804 5533
rect 2836 5387 2844 5713
rect 2856 5467 2864 5693
rect 2876 5547 2884 5852
rect 2916 5827 2924 5864
rect 3016 5707 3024 5853
rect 3056 5767 3064 5864
rect 3096 5767 3104 5976
rect 3153 5900 3167 5913
rect 3156 5896 3164 5900
rect 2916 5596 2924 5693
rect 2993 5608 3007 5613
rect 2936 5507 2944 5564
rect 2856 5456 2873 5467
rect 2860 5453 2873 5456
rect 2616 5267 2624 5333
rect 2647 5293 2653 5307
rect 2587 5116 2604 5124
rect 2516 5076 2524 5113
rect 2596 5087 2604 5116
rect 2616 5107 2624 5193
rect 2676 5167 2684 5332
rect 2696 5127 2704 5333
rect 2716 5207 2724 5374
rect 2776 5340 2784 5344
rect 2773 5327 2787 5340
rect 2856 5346 2864 5433
rect 2956 5347 2964 5533
rect 2996 5524 3004 5594
rect 3016 5527 3024 5693
rect 3053 5600 3067 5613
rect 3056 5596 3064 5600
rect 3096 5596 3104 5633
rect 2976 5516 3004 5524
rect 2976 5387 2984 5516
rect 2996 5376 3004 5453
rect 3036 5387 3044 5453
rect 2416 5040 2424 5044
rect 2413 5027 2427 5040
rect 2416 4987 2424 5013
rect 2296 4876 2324 4884
rect 2276 4807 2284 4853
rect 2296 4826 2304 4876
rect 2356 4856 2364 4893
rect 2396 4856 2404 4913
rect 2336 4820 2344 4824
rect 2376 4820 2384 4824
rect 2056 4507 2064 4554
rect 2036 4476 2064 4484
rect 1993 4344 2007 4353
rect 1976 4340 2007 4344
rect 1976 4336 2004 4340
rect 1956 4067 1964 4304
rect 2016 4300 2024 4304
rect 2013 4287 2027 4300
rect 1976 4207 1984 4273
rect 1773 4040 1787 4053
rect 1776 4036 1784 4040
rect 1736 3904 1744 3993
rect 1756 3927 1764 4004
rect 1787 3984 1800 3986
rect 1787 3980 1804 3984
rect 1787 3973 1807 3980
rect 1793 3967 1807 3973
rect 1836 3967 1844 3993
rect 1736 3900 1764 3904
rect 1736 3896 1767 3900
rect 1753 3887 1767 3896
rect 1736 3816 1744 3853
rect 1776 3827 1784 3933
rect 1836 3844 1844 3953
rect 1856 3947 1864 4053
rect 1873 4047 1887 4053
rect 1956 4004 1964 4053
rect 1996 4047 2004 4213
rect 2056 4127 2064 4476
rect 2076 4287 2084 4473
rect 2156 4467 2164 4524
rect 2176 4487 2184 4513
rect 2196 4507 2204 4673
rect 2136 4336 2144 4393
rect 2116 4287 2124 4304
rect 2116 4244 2124 4273
rect 2116 4236 2144 4244
rect 1936 3996 1964 4004
rect 1816 3836 1844 3844
rect 1816 3816 1824 3836
rect 1856 3816 1864 3853
rect 1896 3827 1904 3873
rect 1756 3780 1764 3784
rect 1676 3747 1684 3772
rect 1753 3767 1767 3780
rect 1707 3753 1713 3765
rect 1656 3567 1664 3632
rect 1716 3547 1724 3653
rect 1736 3587 1744 3613
rect 1756 3607 1764 3732
rect 1776 3727 1784 3773
rect 1880 3784 1893 3787
rect 1876 3776 1893 3784
rect 1880 3773 1893 3776
rect 1836 3764 1844 3772
rect 1916 3767 1924 3853
rect 1936 3847 1944 3996
rect 1956 3827 1964 3973
rect 1976 3967 1984 4034
rect 2013 4040 2027 4053
rect 2016 4036 2024 4040
rect 2096 4007 2104 4233
rect 2136 4184 2144 4236
rect 2156 4204 2164 4304
rect 2196 4247 2204 4472
rect 2156 4196 2184 4204
rect 2136 4176 2164 4184
rect 2036 3947 2044 4004
rect 2016 3816 2024 3853
rect 1836 3756 1864 3764
rect 1796 3707 1804 3733
rect 1836 3707 1844 3733
rect 1856 3724 1864 3756
rect 1856 3716 1884 3724
rect 1416 3007 1424 3133
rect 1456 3127 1464 3264
rect 1496 3008 1504 3193
rect 1476 2927 1484 2964
rect 1487 2916 1504 2924
rect 1496 2807 1504 2916
rect 1516 2807 1524 2953
rect 1536 2804 1544 3373
rect 1556 3307 1564 3333
rect 1616 3307 1624 3333
rect 1600 3304 1613 3307
rect 1596 3296 1613 3304
rect 1600 3293 1613 3296
rect 1556 2947 1564 3253
rect 1636 3147 1644 3473
rect 1656 3447 1664 3472
rect 1716 3467 1724 3533
rect 1736 3507 1744 3573
rect 1816 3516 1824 3673
rect 1876 3667 1884 3716
rect 1853 3567 1867 3573
rect 1736 3447 1744 3493
rect 1656 3327 1664 3433
rect 1713 3300 1727 3313
rect 1716 3296 1724 3300
rect 1756 3296 1764 3333
rect 1776 3307 1784 3453
rect 1796 3447 1804 3484
rect 1836 3464 1844 3472
rect 1816 3456 1844 3464
rect 1656 3207 1664 3292
rect 1687 3256 1704 3264
rect 1676 3187 1684 3253
rect 1696 3147 1704 3233
rect 1716 3127 1724 3213
rect 1736 3207 1744 3264
rect 1616 3047 1624 3073
rect 1676 3067 1684 3093
rect 1616 2996 1624 3033
rect 1653 3000 1667 3013
rect 1696 3007 1704 3053
rect 1656 2996 1664 3000
rect 1713 3000 1727 3013
rect 1716 2996 1724 3000
rect 1756 2996 1764 3073
rect 1776 3067 1784 3253
rect 1796 3207 1804 3313
rect 1816 3027 1824 3456
rect 1876 3447 1884 3653
rect 1896 3527 1904 3593
rect 1936 3587 1944 3812
rect 1956 3707 1964 3773
rect 2036 3780 2044 3784
rect 2033 3767 2047 3780
rect 1916 3524 1924 3573
rect 1956 3547 1964 3613
rect 1916 3516 1944 3524
rect 1976 3516 1984 3633
rect 2056 3527 2064 3773
rect 2076 3767 2084 3993
rect 2096 3767 2104 3953
rect 2116 3727 2124 4113
rect 2133 4047 2147 4053
rect 2156 4048 2164 4176
rect 2176 4127 2184 4196
rect 2216 4067 2224 4573
rect 2256 4556 2264 4733
rect 2296 4627 2304 4812
rect 2333 4807 2347 4820
rect 2373 4807 2387 4820
rect 2296 4487 2304 4524
rect 2296 4336 2304 4413
rect 2256 4147 2264 4304
rect 2256 4036 2264 4112
rect 2336 4087 2344 4653
rect 2356 4568 2364 4693
rect 2396 4667 2404 4733
rect 2416 4707 2424 4813
rect 2436 4727 2444 4893
rect 2376 4556 2384 4593
rect 2436 4567 2444 4613
rect 2456 4547 2464 5032
rect 2476 4927 2484 5033
rect 2536 4927 2544 5044
rect 2516 4856 2524 4913
rect 2596 4887 2604 4913
rect 2616 4907 2624 5072
rect 2616 4827 2624 4872
rect 2613 4807 2627 4813
rect 2536 4767 2544 4804
rect 2536 4607 2544 4753
rect 2616 4547 2624 4593
rect 2416 4516 2444 4524
rect 2356 4347 2364 4493
rect 2436 4444 2444 4516
rect 2456 4467 2464 4533
rect 2436 4436 2473 4444
rect 2536 4427 2544 4484
rect 2416 4347 2424 4393
rect 2436 4367 2444 4413
rect 2456 4347 2464 4373
rect 2436 4336 2453 4344
rect 2356 4304 2364 4333
rect 2496 4327 2504 4413
rect 2636 4407 2644 5113
rect 2667 5044 2680 5047
rect 2667 5036 2684 5044
rect 2667 5033 2680 5036
rect 2687 4884 2700 4887
rect 2687 4873 2704 4884
rect 2696 4856 2704 4873
rect 2736 4867 2744 5033
rect 2756 4884 2764 5173
rect 2776 5047 2784 5213
rect 2836 5107 2844 5333
rect 2916 5340 2924 5344
rect 2873 5324 2887 5333
rect 2913 5327 2927 5340
rect 2873 5320 2904 5324
rect 2876 5316 2904 5320
rect 2876 5076 2884 5273
rect 2896 5267 2904 5316
rect 2916 5047 2924 5193
rect 2756 4876 2784 4884
rect 2756 4826 2764 4853
rect 2656 4447 2664 4593
rect 2696 4556 2704 4653
rect 2736 4647 2744 4813
rect 2356 4296 2384 4304
rect 2376 4227 2384 4296
rect 2296 4036 2304 4073
rect 2353 4044 2367 4053
rect 2347 4040 2367 4044
rect 2347 4036 2364 4040
rect 2176 3996 2204 4004
rect 2136 3827 2144 3953
rect 2176 3816 2184 3873
rect 2196 3827 2204 3996
rect 2216 3847 2224 4032
rect 2236 3827 2244 3913
rect 2276 3887 2284 4004
rect 2316 3984 2324 4004
rect 2316 3976 2333 3984
rect 2156 3780 2164 3784
rect 2153 3767 2167 3780
rect 2206 3772 2207 3780
rect 2193 3765 2207 3772
rect 2193 3760 2213 3765
rect 2196 3756 2213 3760
rect 2096 3516 2104 3713
rect 2136 3707 2144 3753
rect 2200 3751 2213 3756
rect 1836 3307 1844 3433
rect 1896 3387 1904 3492
rect 1876 3296 1884 3353
rect 1936 3307 1944 3413
rect 1996 3387 2004 3484
rect 2036 3427 2044 3513
rect 2053 3467 2067 3473
rect 2016 3367 2024 3393
rect 2016 3308 2024 3332
rect 2056 3327 2064 3453
rect 2076 3407 2084 3484
rect 2116 3480 2124 3484
rect 2113 3467 2127 3480
rect 2136 3447 2144 3473
rect 2156 3327 2164 3653
rect 2196 3516 2204 3573
rect 2256 3544 2264 3833
rect 2276 3787 2284 3873
rect 2336 3827 2344 3973
rect 2356 3828 2364 3993
rect 2376 3987 2384 4213
rect 2396 4067 2404 4304
rect 2416 4044 2424 4293
rect 2496 4267 2504 4313
rect 2656 4287 2664 4433
rect 2676 4347 2684 4393
rect 2696 4367 2704 4433
rect 2736 4427 2744 4524
rect 2716 4336 2724 4393
rect 2736 4387 2744 4413
rect 2756 4364 2764 4513
rect 2776 4407 2784 4876
rect 2796 4827 2804 4893
rect 2816 4867 2824 5013
rect 2836 4967 2844 5044
rect 2936 5044 2944 5253
rect 2976 5187 2984 5333
rect 3016 5247 3024 5344
rect 3036 5204 3044 5333
rect 3056 5227 3064 5513
rect 3076 5467 3084 5564
rect 3136 5487 3144 5633
rect 3176 5608 3184 5852
rect 3196 5596 3204 5813
rect 3236 5807 3244 6076
rect 3236 5687 3244 5753
rect 3236 5596 3244 5673
rect 3256 5647 3264 6193
rect 3296 6087 3304 6133
rect 3333 6120 3347 6133
rect 3336 6116 3344 6120
rect 3376 6116 3384 6173
rect 3536 6116 3544 6193
rect 3356 5947 3364 6084
rect 3396 6047 3404 6084
rect 3456 6047 3464 6114
rect 3276 5787 3284 5933
rect 3496 5896 3504 5973
rect 3516 5927 3524 6084
rect 3556 5867 3564 5993
rect 3576 5987 3584 6114
rect 3636 6047 3644 6084
rect 3716 6047 3724 6153
rect 3816 6116 3824 6153
rect 3756 5987 3764 6084
rect 3613 5900 3627 5913
rect 3616 5896 3624 5900
rect 3676 5887 3684 5913
rect 3727 5904 3740 5907
rect 3727 5896 3744 5904
rect 3776 5896 3784 6013
rect 3796 6007 3804 6084
rect 3727 5893 3740 5896
rect 3336 5608 3344 5733
rect 3356 5667 3364 5831
rect 3396 5827 3404 5864
rect 3376 5596 3384 5713
rect 3176 5407 3184 5493
rect 3133 5380 3147 5393
rect 3173 5387 3187 5393
rect 3136 5376 3144 5380
rect 3196 5347 3204 5413
rect 3096 5287 3104 5344
rect 3176 5247 3184 5333
rect 3193 5327 3207 5333
rect 3216 5287 3224 5433
rect 3036 5196 3064 5204
rect 2976 5088 2984 5152
rect 3016 5088 3024 5173
rect 2936 5036 2964 5044
rect 2836 4868 2844 4893
rect 2796 4567 2804 4792
rect 2896 4747 2904 4824
rect 2796 4387 2804 4433
rect 2756 4360 2804 4364
rect 2756 4356 2807 4360
rect 2793 4347 2807 4356
rect 2816 4344 2824 4493
rect 2876 4467 2884 4633
rect 2896 4567 2904 4733
rect 2916 4587 2924 4693
rect 2936 4647 2944 4973
rect 2956 4967 2964 5036
rect 3056 5044 3064 5196
rect 3116 5076 3124 5153
rect 3156 5076 3164 5153
rect 3056 5036 3084 5044
rect 3056 4967 3064 5013
rect 2996 4856 3004 4893
rect 3056 4867 3064 4893
rect 2976 4820 2984 4824
rect 2973 4807 2987 4820
rect 2947 4604 2960 4607
rect 2947 4600 2964 4604
rect 2947 4593 2967 4600
rect 2953 4587 2967 4593
rect 2927 4584 2940 4587
rect 2927 4573 2944 4584
rect 2936 4556 2944 4573
rect 2976 4556 2984 4793
rect 3016 4727 3024 4824
rect 3036 4707 3044 4793
rect 3016 4526 3024 4573
rect 2896 4364 2904 4513
rect 2916 4387 2924 4473
rect 3036 4447 3044 4693
rect 3076 4667 3084 5036
rect 3096 4824 3104 5032
rect 3136 4927 3144 5044
rect 3176 4947 3184 5032
rect 3196 4907 3204 5073
rect 3216 5027 3224 5233
rect 3236 5087 3244 5473
rect 3276 5447 3284 5593
rect 3293 5380 3307 5393
rect 3336 5387 3344 5513
rect 3356 5487 3364 5564
rect 3296 5376 3304 5380
rect 3276 5340 3284 5344
rect 3256 5224 3264 5333
rect 3273 5327 3287 5340
rect 3313 5327 3327 5332
rect 3256 5216 3284 5224
rect 3256 5076 3264 5193
rect 3276 5147 3284 5216
rect 3336 5076 3344 5233
rect 3356 5227 3364 5452
rect 3376 5347 3384 5393
rect 3396 5387 3404 5473
rect 3416 5407 3424 5793
rect 3476 5787 3484 5864
rect 3696 5866 3704 5893
rect 3436 5547 3444 5653
rect 3516 5596 3524 5653
rect 3556 5608 3564 5813
rect 3596 5787 3604 5864
rect 3636 5784 3644 5852
rect 3616 5776 3644 5784
rect 3496 5560 3504 5564
rect 3493 5547 3507 5560
rect 3436 5376 3444 5533
rect 3496 5507 3504 5533
rect 3476 5376 3484 5493
rect 3496 5407 3504 5472
rect 3536 5467 3544 5564
rect 3536 5387 3544 5413
rect 3556 5376 3564 5533
rect 3576 5487 3584 5553
rect 3596 5467 3604 5752
rect 3616 5424 3624 5776
rect 3656 5596 3664 5773
rect 3676 5667 3684 5852
rect 3756 5844 3764 5864
rect 3736 5836 3764 5844
rect 3696 5608 3704 5713
rect 3636 5524 3644 5553
rect 3636 5516 3653 5524
rect 3636 5447 3644 5492
rect 3616 5416 3644 5424
rect 3636 5387 3644 5416
rect 3316 5040 3324 5044
rect 3313 5027 3327 5040
rect 3096 4816 3124 4824
rect 3136 4820 3144 4824
rect 3176 4820 3184 4824
rect 3096 4567 3104 4593
rect 3116 4556 3124 4816
rect 3133 4807 3147 4820
rect 3173 4807 3187 4820
rect 3196 4784 3204 4812
rect 3216 4787 3224 4953
rect 3176 4776 3204 4784
rect 2896 4356 2924 4364
rect 2816 4336 2844 4344
rect 2396 4036 2424 4044
rect 2436 4036 2444 4133
rect 2476 4067 2484 4093
rect 2473 4040 2487 4053
rect 2476 4036 2484 4040
rect 2276 3587 2284 3773
rect 2336 3747 2344 3773
rect 2256 3536 2284 3544
rect 2276 3516 2284 3536
rect 2296 3527 2304 3733
rect 2216 3464 2224 3484
rect 2256 3480 2264 3484
rect 2253 3467 2267 3480
rect 2216 3456 2244 3464
rect 2236 3424 2244 3456
rect 2253 3447 2267 3453
rect 2236 3416 2273 3424
rect 2296 3424 2304 3473
rect 2287 3416 2304 3424
rect 1556 2827 1564 2873
rect 1536 2796 1564 2804
rect 1473 2780 1487 2793
rect 1476 2776 1484 2780
rect 1536 2747 1544 2773
rect 1416 2687 1424 2744
rect 1456 2707 1464 2744
rect 1253 2487 1267 2493
rect 1196 2476 1204 2480
rect 1353 2480 1367 2493
rect 1356 2476 1364 2480
rect 1096 2367 1104 2393
rect 1036 2220 1044 2224
rect 1033 2207 1047 2220
rect 1036 2067 1044 2193
rect 1076 2187 1084 2224
rect 1116 2167 1124 2373
rect 1156 2324 1164 2373
rect 1176 2327 1184 2444
rect 1236 2387 1244 2452
rect 1287 2444 1300 2447
rect 1287 2436 1304 2444
rect 1287 2433 1300 2436
rect 1376 2407 1384 2433
rect 1136 2316 1164 2324
rect 1136 2267 1144 2316
rect 1167 2296 1193 2304
rect 1276 2226 1284 2313
rect 1336 2268 1344 2333
rect 1376 2256 1384 2393
rect 1396 2347 1404 2573
rect 1416 2327 1424 2513
rect 1436 2287 1444 2493
rect 1493 2480 1507 2493
rect 1496 2476 1504 2480
rect 1536 2476 1544 2712
rect 1556 2587 1564 2796
rect 1576 2787 1584 2953
rect 1596 2827 1604 2964
rect 1636 2960 1644 2964
rect 1633 2947 1647 2960
rect 1616 2804 1624 2853
rect 1636 2827 1644 2873
rect 1607 2796 1624 2804
rect 1596 2776 1604 2792
rect 1573 2724 1587 2733
rect 1573 2720 1604 2724
rect 1576 2716 1604 2720
rect 1476 2367 1484 2444
rect 1516 2440 1524 2444
rect 1513 2427 1527 2440
rect 1456 2264 1464 2333
rect 1436 2256 1464 2264
rect 1493 2260 1507 2273
rect 1496 2256 1504 2260
rect 1156 2187 1164 2224
rect 1196 2167 1204 2224
rect 1276 2167 1284 2212
rect 1316 2187 1324 2212
rect 996 1956 1004 1993
rect 1316 1987 1324 2113
rect 1356 2047 1364 2224
rect 1033 1968 1047 1973
rect 1016 1904 1024 1912
rect 996 1896 1024 1904
rect 956 1736 964 1793
rect 996 1748 1004 1896
rect 1076 1887 1084 1973
rect 1153 1960 1167 1973
rect 1156 1956 1164 1960
rect 1316 1956 1324 1973
rect 1356 1967 1364 2033
rect 1136 1904 1144 1924
rect 1136 1896 1164 1904
rect 1076 1736 1084 1813
rect 1016 1700 1024 1704
rect 1013 1687 1027 1700
rect 1136 1687 1144 1873
rect 1156 1804 1164 1896
rect 1236 1824 1244 1954
rect 1236 1816 1253 1824
rect 1156 1796 1184 1804
rect 996 1567 1004 1593
rect 953 1440 967 1453
rect 956 1436 964 1440
rect 996 1436 1004 1553
rect 876 1376 904 1384
rect 716 1186 724 1273
rect 816 1216 824 1253
rect 856 1227 864 1293
rect 556 916 564 1133
rect 356 787 364 873
rect 396 767 404 884
rect 436 847 444 884
rect 616 847 624 1151
rect 516 776 564 784
rect 336 696 364 704
rect 216 427 224 696
rect 356 666 364 696
rect 276 587 284 664
rect 416 660 424 664
rect 356 627 364 652
rect 413 647 427 660
rect 456 627 464 664
rect 156 396 164 400
rect 207 396 224 404
rect 256 396 264 473
rect 96 287 104 364
rect 236 327 244 364
rect 96 176 104 233
rect 136 176 144 273
rect 276 247 284 364
rect 316 327 324 413
rect 416 396 424 493
rect 496 447 504 693
rect 493 427 507 433
rect 453 400 467 413
rect 516 408 524 776
rect 536 707 544 753
rect 556 747 564 776
rect 576 696 584 773
rect 616 696 624 733
rect 636 707 644 933
rect 596 660 604 664
rect 593 647 607 660
rect 596 587 604 633
rect 456 396 464 400
rect 556 396 564 493
rect 396 327 404 364
rect 256 176 264 213
rect 276 187 284 233
rect 396 207 404 313
rect 536 307 544 364
rect 416 188 424 233
rect 496 176 504 273
rect 536 176 544 253
rect 316 67 324 173
rect 476 140 484 144
rect 516 140 524 144
rect 473 127 487 140
rect 513 127 527 140
rect 576 127 584 352
rect 616 307 624 433
rect 636 367 644 394
rect 656 347 664 1133
rect 736 916 744 1213
rect 836 1087 844 1172
rect 876 1147 884 1376
rect 936 1367 944 1404
rect 956 1216 964 1373
rect 976 1267 984 1404
rect 936 1180 944 1184
rect 933 1167 947 1180
rect 856 1067 864 1093
rect 776 887 784 953
rect 853 920 867 933
rect 856 916 864 920
rect 716 767 724 884
rect 936 886 944 1153
rect 976 1047 984 1184
rect 956 1036 973 1044
rect 876 847 884 884
rect 756 696 764 733
rect 796 696 804 773
rect 816 707 824 833
rect 936 787 944 872
rect 956 867 964 1036
rect 996 1007 1004 1173
rect 1016 1167 1024 1333
rect 1036 1307 1044 1593
rect 1056 1387 1064 1473
rect 1076 1327 1084 1513
rect 1156 1487 1164 1773
rect 1176 1527 1184 1796
rect 1216 1736 1224 1773
rect 1256 1736 1264 1813
rect 1296 1747 1304 1924
rect 1376 1887 1384 2193
rect 1396 2167 1404 2224
rect 1436 2207 1444 2256
rect 1556 2227 1564 2353
rect 1396 1967 1404 2073
rect 1416 1956 1424 2053
rect 1456 1956 1464 2033
rect 1476 2007 1484 2212
rect 1536 2147 1544 2213
rect 1576 2067 1584 2553
rect 1596 2547 1604 2716
rect 1636 2647 1644 2733
rect 1656 2707 1664 2833
rect 1676 2727 1684 2893
rect 1696 2747 1704 2953
rect 1716 2827 1724 2933
rect 1736 2927 1744 2964
rect 1776 2807 1784 2964
rect 1816 2947 1824 2992
rect 1836 2907 1844 3253
rect 1856 3147 1864 3264
rect 1956 3264 1964 3294
rect 1956 3256 1984 3264
rect 1856 3007 1864 3093
rect 1896 2996 1904 3033
rect 1916 3027 1924 3093
rect 1936 3047 1944 3253
rect 1916 3015 1933 3027
rect 1920 3013 1933 3015
rect 1956 3007 1964 3113
rect 1876 2887 1884 2964
rect 1976 2964 1984 3256
rect 2056 3260 2064 3264
rect 2053 3247 2067 3260
rect 2073 3244 2087 3253
rect 2116 3247 2124 3264
rect 2073 3240 2104 3244
rect 2076 3236 2104 3240
rect 2116 3236 2133 3247
rect 2016 3167 2024 3233
rect 1956 2956 1984 2964
rect 1956 2947 1964 2956
rect 1776 2796 1793 2807
rect 1780 2794 1793 2796
rect 1727 2784 1740 2787
rect 1727 2776 1744 2784
rect 1727 2773 1740 2776
rect 1913 2780 1927 2793
rect 1916 2776 1924 2780
rect 1656 2476 1664 2573
rect 1696 2488 1704 2593
rect 1636 2440 1644 2444
rect 1633 2427 1647 2440
rect 1676 2387 1684 2444
rect 1596 2167 1604 2373
rect 1696 2347 1704 2433
rect 1716 2427 1724 2493
rect 1736 2407 1744 2713
rect 1836 2707 1844 2774
rect 1856 2667 1864 2753
rect 1827 2596 1853 2604
rect 1807 2576 1844 2584
rect 1756 2487 1764 2533
rect 1816 2527 1824 2553
rect 1836 2547 1844 2576
rect 1773 2480 1787 2493
rect 1776 2476 1784 2480
rect 1796 2440 1804 2444
rect 1656 2307 1664 2333
rect 1633 2260 1647 2273
rect 1636 2256 1644 2260
rect 1676 2256 1684 2293
rect 1696 2267 1704 2312
rect 1736 2307 1744 2372
rect 1756 2307 1764 2432
rect 1793 2427 1807 2440
rect 1876 2407 1884 2713
rect 1896 2707 1904 2744
rect 1896 2487 1904 2653
rect 1916 2488 1924 2593
rect 1956 2547 1964 2933
rect 1976 2787 1984 2933
rect 1996 2807 2004 3033
rect 2016 3007 2024 3153
rect 2033 3027 2047 3033
rect 2056 2996 2064 3193
rect 2076 3067 2084 3213
rect 2096 3107 2104 3236
rect 2120 3233 2133 3236
rect 2116 3007 2124 3193
rect 2156 3167 2164 3264
rect 2176 3187 2184 3253
rect 2196 3247 2204 3333
rect 2216 3127 2224 3393
rect 2256 3367 2264 3393
rect 2316 3387 2324 3713
rect 2336 3347 2344 3693
rect 2376 3647 2384 3753
rect 2396 3747 2404 4036
rect 2456 3827 2464 4004
rect 2516 3847 2524 4273
rect 2696 4227 2704 4293
rect 2736 4267 2744 4304
rect 2536 3907 2544 4173
rect 2576 4167 2584 4193
rect 2613 4040 2627 4053
rect 2636 4047 2644 4113
rect 2656 4107 2664 4213
rect 2687 4093 2693 4107
rect 2616 4036 2624 4040
rect 2656 3907 2664 4053
rect 2613 3887 2627 3893
rect 2620 3866 2640 3867
rect 2473 3820 2487 3833
rect 2476 3816 2484 3820
rect 2556 3816 2564 3853
rect 2627 3853 2633 3866
rect 2356 3527 2364 3633
rect 2376 3516 2384 3573
rect 2416 3527 2424 3673
rect 2436 3667 2444 3784
rect 2276 3296 2284 3333
rect 2236 3207 2244 3253
rect 2256 3167 2264 3264
rect 2316 3207 2324 3264
rect 2136 2984 2144 3093
rect 2116 2976 2144 2984
rect 2036 2960 2044 2964
rect 2033 2947 2047 2960
rect 2016 2776 2024 2873
rect 2096 2864 2104 2953
rect 2076 2856 2104 2864
rect 2056 2827 2064 2853
rect 2016 2687 2024 2713
rect 1953 2480 1967 2493
rect 1956 2476 1964 2480
rect 1780 2304 1793 2307
rect 1776 2293 1793 2304
rect 1776 2268 1784 2293
rect 1816 2256 1824 2313
rect 1856 2287 1864 2373
rect 1876 2267 1884 2333
rect 1896 2267 1904 2433
rect 1916 2347 1924 2413
rect 1936 2407 1944 2444
rect 1616 2147 1624 2213
rect 1716 2187 1724 2254
rect 1933 2260 1947 2273
rect 1956 2267 1964 2373
rect 1976 2367 1984 2433
rect 1996 2284 2004 2453
rect 2016 2447 2024 2673
rect 2036 2627 2044 2744
rect 2076 2607 2084 2856
rect 2096 2787 2104 2833
rect 2116 2787 2124 2976
rect 2136 2827 2144 2953
rect 2156 2887 2164 3093
rect 2176 3007 2184 3033
rect 2196 2996 2204 3073
rect 2276 3067 2284 3193
rect 2316 3107 2324 3172
rect 2336 3084 2344 3233
rect 2356 3187 2364 3453
rect 2436 3387 2444 3593
rect 2376 3327 2384 3373
rect 2396 3307 2404 3373
rect 2456 3367 2464 3753
rect 2476 3564 2484 3613
rect 2496 3607 2504 3773
rect 2536 3707 2544 3784
rect 2476 3556 2504 3564
rect 2496 3516 2504 3556
rect 2556 3527 2564 3753
rect 2576 3747 2584 3784
rect 2576 3547 2584 3733
rect 2636 3664 2644 3813
rect 2656 3767 2664 3872
rect 2636 3656 2664 3664
rect 2536 3516 2553 3524
rect 2636 3524 2644 3633
rect 2656 3607 2664 3656
rect 2676 3627 2684 4072
rect 2716 4036 2724 4153
rect 2776 4047 2784 4304
rect 2696 3867 2704 3992
rect 2773 3987 2787 3993
rect 2696 3827 2704 3853
rect 2713 3847 2727 3853
rect 2713 3820 2727 3833
rect 2716 3816 2724 3820
rect 2756 3816 2764 3873
rect 2796 3867 2804 4273
rect 2816 4067 2824 4293
rect 2833 4087 2847 4093
rect 2833 4080 2853 4087
rect 2836 4076 2853 4080
rect 2840 4073 2853 4076
rect 2876 4044 2884 4173
rect 2896 4167 2904 4333
rect 2876 4036 2904 4044
rect 2816 3996 2833 4004
rect 2796 3787 2804 3832
rect 2816 3827 2824 3996
rect 2876 3967 2884 3993
rect 2896 3847 2904 4036
rect 2916 4007 2924 4356
rect 2936 4347 2944 4433
rect 3056 4344 3064 4413
rect 3056 4336 3084 4344
rect 2960 4304 2973 4307
rect 2956 4296 2973 4304
rect 2960 4293 2973 4296
rect 3016 4267 3024 4304
rect 3136 4204 3144 4493
rect 3116 4196 3144 4204
rect 2956 4047 2964 4193
rect 3016 4036 3024 4153
rect 2936 3964 2944 4033
rect 2916 3956 2944 3964
rect 2916 3887 2924 3956
rect 2916 3824 2924 3873
rect 2896 3816 2924 3824
rect 2636 3516 2684 3524
rect 2516 3480 2524 3484
rect 2476 3307 2484 3473
rect 2513 3467 2527 3480
rect 2576 3447 2584 3493
rect 2676 3484 2684 3516
rect 2493 3347 2507 3353
rect 2376 3147 2384 3292
rect 2416 3260 2424 3264
rect 2396 3227 2404 3253
rect 2413 3247 2427 3260
rect 2316 3076 2344 3084
rect 2296 2996 2304 3033
rect 2316 3027 2324 3076
rect 2176 2927 2184 2953
rect 2176 2807 2184 2853
rect 2196 2824 2204 2933
rect 2216 2847 2224 2964
rect 2233 2927 2247 2933
rect 2196 2816 2224 2824
rect 2176 2776 2184 2793
rect 2016 2307 2024 2353
rect 1996 2276 2013 2284
rect 1936 2256 1944 2260
rect 1747 2224 1760 2227
rect 1747 2216 1764 2224
rect 1796 2220 1804 2224
rect 1747 2213 1760 2216
rect 1793 2207 1807 2220
rect 1536 1968 1544 2053
rect 1596 2047 1604 2073
rect 1616 2047 1624 2112
rect 1656 2067 1664 2173
rect 1656 2027 1664 2053
rect 1576 1956 1584 2013
rect 1676 2004 1684 2133
rect 1716 2007 1724 2093
rect 1656 1996 1684 2004
rect 1656 1956 1664 1996
rect 1096 1447 1104 1473
rect 1133 1440 1147 1453
rect 1196 1448 1204 1693
rect 1276 1667 1284 1704
rect 1316 1547 1324 1873
rect 1336 1727 1344 1753
rect 1396 1736 1404 1793
rect 1436 1767 1444 1924
rect 1496 1787 1504 1953
rect 1376 1667 1384 1704
rect 1233 1467 1247 1473
rect 1136 1436 1144 1440
rect 1176 1436 1193 1444
rect 1236 1436 1244 1453
rect 1056 1316 1073 1324
rect 1036 947 1044 1213
rect 1056 1167 1064 1316
rect 1096 1287 1104 1393
rect 1116 1347 1124 1404
rect 1156 1400 1164 1404
rect 1256 1400 1264 1404
rect 1153 1387 1167 1400
rect 1253 1387 1267 1400
rect 1136 1216 1144 1273
rect 1013 928 1027 933
rect 1056 916 1064 993
rect 1076 987 1084 1173
rect 1116 1087 1124 1184
rect 1156 1180 1164 1184
rect 1153 1167 1167 1180
rect 1196 1167 1204 1273
rect 1256 1216 1264 1313
rect 1296 1267 1304 1404
rect 1336 1387 1344 1473
rect 1236 1180 1244 1184
rect 1233 1167 1247 1180
rect 1276 1127 1284 1184
rect 1276 1087 1284 1113
rect 1076 947 1084 973
rect 1196 947 1204 993
rect 676 647 684 693
rect 776 627 784 664
rect 836 587 844 733
rect 796 367 804 473
rect 856 467 864 733
rect 996 708 1004 884
rect 1036 880 1044 884
rect 1033 867 1047 880
rect 1096 807 1104 933
rect 1153 920 1167 933
rect 1193 920 1207 933
rect 1156 916 1164 920
rect 1196 916 1204 920
rect 1236 886 1244 973
rect 1296 916 1304 953
rect 1316 947 1324 1173
rect 1336 1047 1344 1253
rect 1356 1167 1364 1293
rect 1376 1186 1384 1473
rect 1416 1436 1424 1593
rect 1436 1487 1444 1713
rect 1456 1487 1464 1773
rect 1536 1736 1544 1873
rect 1556 1827 1564 1924
rect 1576 1747 1584 1793
rect 1516 1647 1524 1704
rect 1596 1587 1604 1813
rect 1616 1787 1624 1954
rect 1616 1667 1624 1752
rect 1636 1747 1644 1913
rect 1656 1736 1664 1813
rect 1676 1807 1684 1924
rect 1736 1924 1744 2153
rect 1756 1967 1764 2193
rect 1816 1984 1824 2193
rect 1836 2107 1844 2224
rect 1796 1976 1824 1984
rect 1796 1956 1804 1976
rect 1833 1960 1847 1973
rect 1856 1967 1864 2213
rect 1836 1956 1844 1960
rect 1736 1916 1784 1924
rect 1696 1827 1704 1873
rect 1716 1867 1724 1913
rect 1776 1904 1784 1916
rect 1776 1896 1804 1904
rect 1693 1740 1707 1753
rect 1756 1747 1764 1893
rect 1796 1867 1804 1896
rect 1696 1736 1704 1740
rect 1456 1473 1473 1487
rect 1456 1436 1464 1473
rect 1496 1467 1504 1533
rect 1636 1527 1644 1693
rect 1716 1700 1724 1704
rect 1713 1687 1727 1700
rect 1516 1406 1524 1493
rect 1556 1436 1564 1513
rect 1596 1436 1604 1493
rect 1616 1467 1624 1513
rect 1576 1400 1584 1404
rect 1467 1373 1473 1387
rect 1516 1267 1524 1392
rect 1573 1387 1587 1400
rect 1547 1373 1553 1387
rect 1556 1216 1564 1293
rect 1616 1264 1624 1392
rect 1616 1256 1644 1264
rect 1616 1207 1624 1233
rect 1456 1180 1464 1184
rect 1416 1107 1424 1172
rect 1453 1167 1467 1180
rect 1476 1127 1484 1173
rect 1516 1107 1524 1184
rect 1336 967 1344 1033
rect 1576 987 1584 1184
rect 1387 976 1404 984
rect 1376 928 1384 973
rect 1096 696 1104 733
rect 876 547 884 653
rect 996 664 1004 694
rect 916 607 924 652
rect 956 587 964 664
rect 996 656 1044 664
rect 1076 587 1084 664
rect 876 424 884 533
rect 1136 527 1144 693
rect 1156 627 1164 793
rect 1176 747 1184 884
rect 1236 708 1244 733
rect 1273 707 1287 713
rect 1296 666 1304 733
rect 1356 708 1364 884
rect 1396 847 1404 976
rect 1567 933 1573 947
rect 1493 920 1507 933
rect 1496 916 1504 920
rect 1616 927 1624 1073
rect 1636 1027 1644 1256
rect 1636 928 1644 953
rect 1656 947 1664 1453
rect 1676 1407 1684 1653
rect 1736 1627 1744 1693
rect 1756 1647 1764 1712
rect 1776 1667 1784 1853
rect 1816 1827 1824 1924
rect 1833 1740 1847 1753
rect 1836 1736 1844 1740
rect 1876 1736 1884 2213
rect 1967 2224 1980 2227
rect 1967 2213 1984 2224
rect 1893 2187 1907 2193
rect 1976 2167 1984 2213
rect 1896 1947 1904 2113
rect 1976 2087 1984 2132
rect 1996 2107 2004 2213
rect 2016 2107 2024 2272
rect 2036 2167 2044 2533
rect 2096 2507 2104 2752
rect 2156 2740 2164 2744
rect 2116 2584 2124 2733
rect 2153 2727 2167 2740
rect 2216 2727 2224 2816
rect 2116 2576 2133 2584
rect 2136 2547 2144 2573
rect 2067 2504 2080 2507
rect 2067 2493 2084 2504
rect 2076 2476 2084 2493
rect 2133 2480 2147 2493
rect 2156 2487 2164 2653
rect 2136 2476 2144 2480
rect 2056 2267 2064 2393
rect 2096 2367 2104 2432
rect 2116 2327 2124 2353
rect 2176 2287 2184 2713
rect 2196 2307 2204 2493
rect 2216 2487 2224 2613
rect 2236 2584 2244 2873
rect 2256 2787 2264 2833
rect 2276 2807 2284 2953
rect 2316 2847 2324 2964
rect 2356 2960 2364 2964
rect 2353 2947 2367 2960
rect 2336 2867 2344 2933
rect 2376 2924 2384 2953
rect 2396 2947 2404 3053
rect 2356 2916 2384 2924
rect 2296 2776 2304 2813
rect 2356 2787 2364 2916
rect 2416 2907 2424 3093
rect 2436 2927 2444 3213
rect 2456 3147 2464 3264
rect 2476 3107 2484 3253
rect 2496 3247 2504 3333
rect 2516 3187 2524 3393
rect 2553 3367 2567 3373
rect 2476 2996 2484 3033
rect 2536 3004 2544 3353
rect 2596 3347 2604 3473
rect 2616 3464 2624 3484
rect 2656 3476 2684 3484
rect 2616 3456 2644 3464
rect 2636 3427 2644 3456
rect 2556 3307 2564 3332
rect 2636 3307 2644 3413
rect 2616 3260 2624 3264
rect 2613 3247 2627 3260
rect 2567 3233 2573 3245
rect 2576 3007 2584 3113
rect 2536 2996 2564 3004
rect 2396 2784 2404 2853
rect 2456 2807 2464 2933
rect 2396 2776 2413 2784
rect 2256 2707 2264 2733
rect 2276 2647 2284 2744
rect 2316 2724 2324 2744
rect 2296 2716 2324 2724
rect 2236 2576 2264 2584
rect 2236 2476 2244 2553
rect 2256 2487 2264 2576
rect 2296 2547 2304 2716
rect 2276 2436 2304 2444
rect 1933 1968 1947 1973
rect 1980 1964 1993 1967
rect 1976 1956 1993 1964
rect 1980 1953 1993 1956
rect 1936 1706 1944 1813
rect 1816 1700 1824 1704
rect 1813 1687 1827 1700
rect 1720 1464 1733 1467
rect 1716 1453 1733 1464
rect 1716 1448 1727 1453
rect 1776 1307 1784 1573
rect 1796 1527 1804 1573
rect 1856 1567 1864 1704
rect 1796 1447 1804 1513
rect 1856 1467 1864 1513
rect 1876 1487 1884 1673
rect 1896 1467 1904 1704
rect 1916 1547 1924 1633
rect 1956 1607 1964 1753
rect 1976 1747 1984 1873
rect 1996 1827 2004 1913
rect 2016 1768 2024 2093
rect 2036 2047 2044 2073
rect 2056 1984 2064 2213
rect 2116 2184 2124 2224
rect 2116 2176 2144 2184
rect 2076 2027 2084 2153
rect 2096 2047 2104 2073
rect 2116 1987 2124 2073
rect 2036 1976 2064 1984
rect 2036 1887 2044 1976
rect 2073 1964 2087 1973
rect 2136 1968 2144 2176
rect 2156 2087 2164 2253
rect 2216 2256 2224 2413
rect 2256 2287 2264 2433
rect 2296 2287 2304 2436
rect 2316 2387 2324 2593
rect 2336 2487 2344 2733
rect 2376 2647 2384 2744
rect 2416 2607 2424 2713
rect 2456 2704 2464 2733
rect 2476 2727 2484 2913
rect 2456 2696 2484 2704
rect 2353 2480 2367 2493
rect 2416 2487 2424 2572
rect 2436 2567 2444 2693
rect 2356 2476 2364 2480
rect 2436 2446 2444 2473
rect 2336 2407 2344 2433
rect 2256 2256 2304 2264
rect 2356 2256 2364 2333
rect 2373 2267 2387 2273
rect 2176 2184 2184 2252
rect 2193 2207 2207 2213
rect 2206 2200 2207 2207
rect 2176 2176 2204 2184
rect 2153 2027 2167 2033
rect 2056 1960 2087 1964
rect 2056 1956 2084 1960
rect 2056 1907 2064 1956
rect 2156 1956 2164 1992
rect 2096 1748 2104 1853
rect 2116 1847 2124 1924
rect 2196 1847 2204 2176
rect 2216 2127 2224 2193
rect 2236 2167 2244 2224
rect 2213 2027 2227 2033
rect 2236 2007 2244 2053
rect 2276 1987 2284 2173
rect 2296 2167 2304 2256
rect 2336 2207 2344 2224
rect 2336 2196 2353 2207
rect 2340 2193 2353 2196
rect 2367 2196 2384 2204
rect 2336 2027 2344 2173
rect 2296 1964 2304 1993
rect 2276 1956 2304 1964
rect 2116 1747 2124 1773
rect 2036 1687 2044 1704
rect 2073 1687 2087 1693
rect 2036 1676 2053 1687
rect 2040 1673 2053 1676
rect 2096 1607 2104 1734
rect 2176 1736 2184 1773
rect 2216 1747 2224 1853
rect 2116 1524 2124 1693
rect 2136 1604 2144 1673
rect 2156 1627 2164 1692
rect 2136 1596 2164 1604
rect 2156 1547 2164 1596
rect 2116 1516 2132 1524
rect 1827 1464 1840 1467
rect 1827 1453 1844 1464
rect 1836 1436 1844 1453
rect 1873 1440 1887 1452
rect 1876 1436 1884 1440
rect 1856 1400 1864 1404
rect 1853 1387 1867 1400
rect 1916 1387 1924 1434
rect 1936 1407 1944 1513
rect 1976 1447 1984 1473
rect 2056 1436 2064 1493
rect 2136 1436 2144 1513
rect 2156 1467 2164 1512
rect 2196 1447 2204 1692
rect 2236 1647 2244 1893
rect 2256 1747 2264 1924
rect 2316 1787 2324 1933
rect 2336 1867 2344 1973
rect 2256 1507 2264 1693
rect 2276 1667 2284 1704
rect 2296 1567 2304 1633
rect 2216 1407 2224 1493
rect 1816 1327 1824 1353
rect 1976 1327 1984 1393
rect 1996 1384 2004 1404
rect 1996 1376 2024 1384
rect 1693 1220 1707 1233
rect 1856 1228 1864 1253
rect 1976 1244 1984 1313
rect 1956 1236 1984 1244
rect 1696 1216 1704 1220
rect 1956 1216 1964 1236
rect 1996 1216 2004 1353
rect 2016 1227 2024 1376
rect 2053 1220 2067 1233
rect 2056 1216 2064 1220
rect 2096 1216 2104 1392
rect 2116 1367 2124 1404
rect 2156 1367 2164 1404
rect 2116 1327 2124 1353
rect 2116 1296 2153 1304
rect 2116 1247 2124 1296
rect 1796 1186 1804 1213
rect 1576 886 1584 912
rect 1696 886 1704 1013
rect 1716 1007 1724 1184
rect 1716 928 1724 993
rect 1756 967 1764 1184
rect 1796 916 1804 1172
rect 1836 886 1844 1172
rect 1476 707 1484 884
rect 1516 696 1524 793
rect 1656 708 1664 773
rect 1700 704 1713 707
rect 1696 696 1713 704
rect 1700 693 1713 696
rect 1216 660 1224 664
rect 1213 647 1227 660
rect 1327 664 1340 667
rect 1327 656 1344 664
rect 1327 653 1340 656
rect 856 416 884 424
rect 856 396 864 416
rect 896 396 904 453
rect 716 360 724 364
rect 676 327 684 353
rect 713 347 727 360
rect 596 146 604 213
rect 656 176 664 273
rect 736 204 744 253
rect 756 227 764 364
rect 936 364 944 453
rect 956 367 964 493
rect 996 396 1004 513
rect 1036 396 1044 493
rect 876 360 884 364
rect 873 347 887 360
rect 916 356 944 364
rect 816 207 824 313
rect 916 287 924 356
rect 933 327 947 333
rect 736 196 764 204
rect 696 176 744 184
rect 676 140 684 144
rect 673 127 687 140
rect 736 87 744 176
rect 756 47 764 196
rect 836 176 844 253
rect 876 187 884 213
rect 896 107 904 253
rect 916 167 924 273
rect 936 147 944 313
rect 1056 267 1064 364
rect 996 188 1004 253
rect 1096 247 1104 513
rect 1176 467 1184 493
rect 1127 404 1140 407
rect 1127 396 1144 404
rect 1176 396 1184 453
rect 1216 407 1224 533
rect 1127 393 1140 396
rect 1276 396 1284 453
rect 1116 327 1124 353
rect 1096 204 1104 233
rect 1076 196 1104 204
rect 1076 176 1084 196
rect 1096 140 1104 144
rect 976 127 987 132
rect 1093 127 1107 140
rect 1156 127 1164 173
rect 1176 127 1184 233
rect 1236 176 1244 273
rect 1276 176 1284 313
rect 1296 247 1304 364
rect 1376 327 1384 493
rect 1416 467 1424 653
rect 1476 627 1484 693
rect 1736 667 1744 813
rect 1776 787 1784 884
rect 1816 747 1824 773
rect 1856 727 1864 1093
rect 1916 1087 1924 1213
rect 1916 1047 1924 1073
rect 1896 916 1904 973
rect 1933 920 1947 933
rect 1976 927 1984 1184
rect 2156 1186 2164 1253
rect 2196 1244 2204 1393
rect 2216 1247 2224 1372
rect 2316 1367 2324 1593
rect 2356 1564 2364 2153
rect 2376 2107 2384 2196
rect 2396 2007 2404 2273
rect 2416 2167 2424 2293
rect 2436 2247 2444 2293
rect 2456 2287 2464 2673
rect 2476 2487 2484 2696
rect 2496 2687 2504 2893
rect 2516 2787 2524 2813
rect 2536 2807 2544 2873
rect 2556 2827 2564 2996
rect 2596 2996 2604 3153
rect 2636 3127 2644 3253
rect 2636 2996 2644 3053
rect 2656 3027 2664 3476
rect 2676 3304 2684 3333
rect 2696 3327 2704 3773
rect 2736 3647 2744 3784
rect 2936 3786 2944 3893
rect 2956 3827 2964 3993
rect 3036 3996 3064 4004
rect 3036 3867 3044 3996
rect 3116 3907 3124 4196
rect 3156 4044 3164 4553
rect 3176 4507 3184 4776
rect 3236 4567 3244 4853
rect 3256 4647 3264 5013
rect 3296 4947 3304 4973
rect 3316 4868 3324 4893
rect 3276 4667 3284 4693
rect 3256 4556 3264 4633
rect 3216 4427 3224 4524
rect 3296 4427 3304 4753
rect 3316 4567 3324 4793
rect 3356 4767 3364 5032
rect 3376 4867 3384 5312
rect 3396 5207 3404 5333
rect 3436 5167 3444 5313
rect 3456 5267 3464 5344
rect 3496 5247 3504 5332
rect 3616 5307 3624 5332
rect 3436 5076 3444 5153
rect 3516 5087 3524 5193
rect 3636 5187 3644 5333
rect 3396 4967 3404 5073
rect 3536 5047 3544 5173
rect 3556 5107 3564 5133
rect 3596 5088 3604 5133
rect 3636 5076 3644 5173
rect 3656 5087 3664 5513
rect 3456 4927 3464 5044
rect 3476 4947 3484 4973
rect 3396 4856 3404 4913
rect 3436 4856 3444 4893
rect 3496 4824 3504 4993
rect 3556 4987 3564 5072
rect 3596 4867 3604 4973
rect 3416 4787 3424 4824
rect 3456 4787 3464 4824
rect 3496 4816 3524 4824
rect 3316 4524 3324 4553
rect 3336 4547 3344 4713
rect 3496 4547 3504 4593
rect 3516 4567 3524 4816
rect 3576 4747 3584 4824
rect 3556 4647 3564 4673
rect 3576 4647 3584 4733
rect 3596 4556 3604 4813
rect 3616 4787 3624 4853
rect 3616 4567 3624 4693
rect 3316 4516 3344 4524
rect 3196 4247 3204 4304
rect 3256 4296 3284 4304
rect 3276 4267 3284 4296
rect 3256 4127 3264 4193
rect 3136 4036 3164 4044
rect 3136 3867 3144 4036
rect 3276 4024 3284 4253
rect 3296 4087 3304 4373
rect 3316 4107 3324 4473
rect 3336 4387 3344 4516
rect 3416 4407 3424 4484
rect 3336 4036 3344 4073
rect 3356 4067 3364 4304
rect 3396 4044 3404 4304
rect 3456 4247 3464 4373
rect 3496 4348 3504 4493
rect 3556 4487 3564 4524
rect 3536 4336 3544 4373
rect 3576 4347 3584 4433
rect 3516 4127 3524 4304
rect 3576 4207 3584 4273
rect 3596 4147 3604 4393
rect 3616 4267 3624 4473
rect 3636 4367 3644 5013
rect 3656 4987 3664 5033
rect 3676 5027 3684 5493
rect 3736 5467 3744 5836
rect 3796 5767 3804 5793
rect 3856 5787 3864 6233
rect 3776 5487 3784 5564
rect 3836 5387 3844 5593
rect 3856 5567 3864 5713
rect 3876 5607 3884 6253
rect 3896 6128 3904 6153
rect 3913 6128 3927 6133
rect 4016 6127 4024 6153
rect 3896 6087 3904 6114
rect 3913 6064 3927 6073
rect 3976 6080 3984 6084
rect 3973 6067 3987 6080
rect 3913 6060 3944 6064
rect 3916 6056 3944 6060
rect 3936 5896 3944 6056
rect 3976 5896 3984 5933
rect 3956 5847 3964 5864
rect 4016 5847 4024 6053
rect 4036 5947 4044 6114
rect 4067 6084 4080 6087
rect 4067 6076 4084 6084
rect 4067 6073 4080 6076
rect 4136 6067 4144 6113
rect 4156 6027 4164 6114
rect 4216 6047 4224 6084
rect 4296 6084 4304 6153
rect 4356 6128 4364 6213
rect 4376 6207 4384 6233
rect 4396 6116 4404 6153
rect 4276 6076 4304 6084
rect 4236 6007 4244 6053
rect 4256 6024 4264 6072
rect 4276 6047 4284 6076
rect 4256 6016 4284 6024
rect 4196 5967 4204 5993
rect 4136 5908 4144 5933
rect 4276 5927 4284 6016
rect 4296 5927 4304 6053
rect 4336 6027 4344 6084
rect 4253 5900 4267 5913
rect 4256 5896 4264 5900
rect 3896 5596 3904 5733
rect 3936 5687 3944 5753
rect 3956 5707 3964 5833
rect 4076 5827 4084 5852
rect 4116 5807 4124 5864
rect 4186 5853 4187 5860
rect 4173 5847 4187 5853
rect 4236 5860 4244 5864
rect 4233 5847 4247 5860
rect 4336 5866 4344 5992
rect 4356 5927 4364 5993
rect 4376 5927 4384 6084
rect 4396 5896 4404 6033
rect 4436 6007 4444 6233
rect 4796 6116 4804 6153
rect 4556 6086 4564 6113
rect 4456 5967 4464 6072
rect 4516 6047 4524 6072
rect 4433 5900 4447 5913
rect 4436 5896 4444 5900
rect 4476 5866 4484 5973
rect 4496 5947 4504 6033
rect 4536 5896 4544 5933
rect 4556 5924 4564 6072
rect 4576 6047 4584 6093
rect 4556 5916 4584 5924
rect 4576 5896 4584 5916
rect 4616 5907 4624 5933
rect 4636 5866 4644 5973
rect 4276 5807 4284 5853
rect 4416 5827 4424 5864
rect 4396 5816 4413 5824
rect 3856 5376 3864 5513
rect 3876 5507 3884 5553
rect 3916 5487 3924 5564
rect 3956 5504 3964 5553
rect 3996 5527 4004 5693
rect 4016 5607 4024 5653
rect 4036 5647 4044 5753
rect 4056 5596 4064 5773
rect 4236 5596 4244 5713
rect 4376 5647 4384 5793
rect 4376 5607 4384 5633
rect 3956 5496 3984 5504
rect 3896 5376 3904 5453
rect 3976 5447 3984 5496
rect 3936 5387 3944 5433
rect 4016 5404 4024 5553
rect 4036 5527 4044 5564
rect 4076 5527 4084 5564
rect 4136 5484 4144 5594
rect 4176 5560 4184 5564
rect 4173 5547 4187 5560
rect 4216 5487 4224 5564
rect 4136 5476 4153 5484
rect 4016 5396 4044 5404
rect 3947 5376 3964 5384
rect 4036 5376 4044 5396
rect 3736 5267 3744 5344
rect 3716 5167 3724 5233
rect 3776 5227 3784 5344
rect 3816 5307 3824 5373
rect 3876 5324 3884 5344
rect 3856 5316 3884 5324
rect 3827 5156 3844 5164
rect 3696 4887 3704 5113
rect 3776 5076 3784 5113
rect 3816 5076 3824 5153
rect 3836 5127 3844 5156
rect 3716 5007 3724 5033
rect 3756 5024 3764 5044
rect 3756 5016 3784 5024
rect 3756 4867 3764 4973
rect 3776 4947 3784 5016
rect 3796 5007 3804 5044
rect 3856 5027 3864 5316
rect 3916 5267 3924 5332
rect 3936 5247 3944 5332
rect 3876 5087 3884 5233
rect 3956 5204 3964 5376
rect 4076 5307 4084 5433
rect 3976 5247 3984 5273
rect 3936 5196 3964 5204
rect 3896 5076 3904 5133
rect 3936 5087 3944 5196
rect 3956 5127 3964 5173
rect 3976 5084 3984 5233
rect 3956 5076 3984 5084
rect 3916 5040 3924 5044
rect 3913 5027 3927 5040
rect 3816 4947 3824 4973
rect 3796 4856 3804 4913
rect 3656 4787 3664 4853
rect 3696 4707 3704 4824
rect 3656 4344 3664 4673
rect 3696 4556 3704 4672
rect 3776 4527 3784 4713
rect 3716 4447 3724 4524
rect 3716 4364 3724 4393
rect 3716 4356 3744 4364
rect 3736 4350 3744 4356
rect 3636 4336 3664 4344
rect 3636 4187 3644 4336
rect 3656 4207 3664 4293
rect 3676 4267 3684 4304
rect 3387 4036 3404 4044
rect 3276 4016 3293 4024
rect 2993 3820 3007 3833
rect 2996 3816 3004 3820
rect 2796 3707 2804 3752
rect 2716 3367 2724 3613
rect 2796 3547 2804 3693
rect 2856 3587 2864 3753
rect 2876 3627 2884 3784
rect 3056 3767 3064 3833
rect 2896 3687 2904 3753
rect 2753 3520 2767 3533
rect 2756 3516 2764 3520
rect 2796 3516 2804 3533
rect 2853 3527 2867 3533
rect 2873 3520 2887 3533
rect 2876 3516 2884 3520
rect 2916 3516 2924 3653
rect 2996 3528 3004 3693
rect 2776 3427 2784 3484
rect 2736 3307 2744 3373
rect 2676 3296 2704 3304
rect 2676 3127 2684 3253
rect 2716 3227 2724 3264
rect 2676 3004 2684 3113
rect 2696 3047 2704 3193
rect 2676 2996 2704 3004
rect 2696 2967 2704 2996
rect 2616 2960 2624 2964
rect 2613 2947 2627 2960
rect 2533 2780 2547 2793
rect 2536 2776 2544 2780
rect 2596 2767 2604 2933
rect 2656 2867 2664 2964
rect 2716 2927 2724 3013
rect 2736 3007 2744 3253
rect 2756 3107 2764 3313
rect 2776 3247 2784 3353
rect 2816 3327 2824 3433
rect 2836 3367 2844 3493
rect 2936 3407 2944 3484
rect 2873 3307 2887 3313
rect 2896 3247 2904 3373
rect 2976 3347 2984 3453
rect 2996 3447 3004 3514
rect 3016 3387 3024 3573
rect 3036 3367 3044 3673
rect 3056 3524 3064 3633
rect 3076 3567 3084 3853
rect 3156 3816 3164 3993
rect 3296 3967 3304 4013
rect 3496 4004 3504 4093
rect 3396 3927 3404 3993
rect 3196 3867 3204 3893
rect 3196 3816 3204 3853
rect 3216 3827 3224 3873
rect 3227 3824 3240 3827
rect 3227 3816 3244 3824
rect 3227 3813 3240 3816
rect 3096 3767 3104 3813
rect 3136 3780 3144 3784
rect 3133 3767 3147 3780
rect 3176 3747 3184 3772
rect 3176 3607 3184 3633
rect 3196 3607 3204 3693
rect 3216 3567 3224 3753
rect 3296 3744 3304 3913
rect 3416 3907 3424 3953
rect 3496 3947 3504 3990
rect 3516 3927 3524 4033
rect 3636 3967 3644 3993
rect 3316 3787 3324 3833
rect 3436 3827 3444 3913
rect 3456 3784 3464 3893
rect 3296 3736 3313 3744
rect 3376 3744 3384 3773
rect 3476 3767 3484 3873
rect 3507 3836 3564 3844
rect 3556 3816 3564 3836
rect 3356 3736 3384 3744
rect 3316 3667 3324 3733
rect 3356 3687 3364 3736
rect 3056 3516 3084 3524
rect 3156 3527 3164 3553
rect 3236 3516 3244 3593
rect 3256 3527 3264 3633
rect 2776 3167 2784 3233
rect 2756 3027 2764 3093
rect 2816 3028 2824 3153
rect 2836 3087 2844 3113
rect 2756 2944 2764 2964
rect 2756 2936 2784 2944
rect 2736 2807 2744 2833
rect 2733 2780 2747 2793
rect 2736 2776 2744 2780
rect 2516 2547 2524 2713
rect 2533 2707 2547 2713
rect 2556 2687 2564 2744
rect 2576 2667 2584 2733
rect 2616 2727 2624 2773
rect 2636 2704 2644 2753
rect 2776 2746 2784 2936
rect 2796 2927 2804 2964
rect 2796 2787 2804 2892
rect 2836 2788 2844 2953
rect 2856 2907 2864 3193
rect 2876 3127 2884 3213
rect 2896 3047 2904 3173
rect 2916 3067 2924 3333
rect 2936 3227 2944 3253
rect 2893 3000 2907 3012
rect 2896 2996 2904 3000
rect 2936 2996 2944 3153
rect 2996 3087 3004 3264
rect 2973 3000 2987 3013
rect 2996 3007 3004 3073
rect 2976 2996 2984 3000
rect 2876 2867 2884 2953
rect 2956 2887 2964 2964
rect 3016 2927 3024 3213
rect 3036 3207 3044 3313
rect 3076 3296 3084 3333
rect 3096 3327 3104 3484
rect 3136 3427 3144 3484
rect 3156 3447 3164 3473
rect 3116 3296 3124 3393
rect 3136 3347 3144 3413
rect 3096 3227 3104 3264
rect 3047 3136 3073 3144
rect 3036 2967 3044 3053
rect 3056 3007 3064 3113
rect 3136 3107 3144 3173
rect 3176 3107 3184 3473
rect 3196 3407 3204 3453
rect 3216 3447 3224 3484
rect 3256 3427 3264 3473
rect 3276 3467 3284 3653
rect 3496 3627 3504 3773
rect 3536 3627 3544 3784
rect 3576 3747 3584 3784
rect 3616 3627 3624 3893
rect 3656 3847 3664 4133
rect 3676 3907 3684 4113
rect 3696 4047 3704 4253
rect 3716 4167 3724 4293
rect 3716 4036 3724 4153
rect 3776 4144 3784 4193
rect 3796 4167 3804 4793
rect 3856 4787 3864 4824
rect 3816 4568 3824 4613
rect 3876 4607 3884 4813
rect 3896 4584 3904 5013
rect 3916 4687 3924 4893
rect 3936 4727 3944 4913
rect 3976 4887 3984 5033
rect 3996 4927 4004 5293
rect 4036 5187 4044 5213
rect 4016 5127 4024 5153
rect 4036 5076 4044 5173
rect 4066 5113 4067 5120
rect 4053 5107 4067 5113
rect 4076 5076 4084 5113
rect 4096 5107 4104 5413
rect 4156 5376 4164 5473
rect 4256 5347 4264 5533
rect 4276 5347 4284 5594
rect 4340 5384 4353 5387
rect 4336 5376 4353 5384
rect 4340 5373 4353 5376
rect 4376 5347 4384 5513
rect 4396 5447 4404 5816
rect 4556 5687 4564 5864
rect 4416 5427 4424 5673
rect 4516 5596 4524 5633
rect 4596 5596 4604 5693
rect 4656 5604 4664 6044
rect 4676 5907 4684 6033
rect 4736 5987 4744 6073
rect 4856 6007 4864 6084
rect 4896 6007 4904 6114
rect 4936 6047 4944 6213
rect 4956 6207 4964 6304
rect 5116 6247 5124 6304
rect 4976 6116 4984 6153
rect 5013 6120 5027 6133
rect 5016 6116 5024 6120
rect 4747 5976 4764 5984
rect 4716 5896 4724 5953
rect 4756 5907 4764 5976
rect 4776 5866 4784 5953
rect 4796 5907 4804 5993
rect 4996 5987 5004 6084
rect 4836 5896 4844 5933
rect 4816 5747 4824 5813
rect 4656 5596 4684 5604
rect 4436 5527 4444 5594
rect 4456 5507 4464 5553
rect 4536 5507 4544 5564
rect 4616 5560 4624 5564
rect 4613 5547 4627 5560
rect 4536 5447 4544 5493
rect 4596 5388 4604 5513
rect 4636 5487 4644 5513
rect 4656 5464 4664 5553
rect 4676 5487 4684 5596
rect 4696 5507 4704 5633
rect 4736 5596 4744 5713
rect 4816 5607 4824 5673
rect 4656 5456 4684 5464
rect 4116 5147 4124 5333
rect 4216 5307 4224 5344
rect 4287 5340 4304 5344
rect 4287 5336 4307 5340
rect 4216 5244 4224 5293
rect 4236 5267 4244 5333
rect 4293 5327 4307 5336
rect 4496 5346 4504 5373
rect 4356 5307 4364 5333
rect 4216 5236 4244 5244
rect 4156 5187 4164 5213
rect 4136 5107 4144 5153
rect 4016 4987 4024 5033
rect 4056 4927 4064 5044
rect 4033 4860 4047 4873
rect 4076 4868 4084 5013
rect 4096 4987 4104 5044
rect 4116 4927 4124 4993
rect 4136 4947 4144 5033
rect 4156 4887 4164 5133
rect 4176 4907 4184 5193
rect 4207 5184 4220 5187
rect 4207 5173 4224 5184
rect 4196 5087 4204 5152
rect 4216 5076 4224 5173
rect 4236 5107 4244 5236
rect 4336 5207 4344 5233
rect 4256 5076 4264 5173
rect 4296 5076 4304 5193
rect 4356 5084 4364 5293
rect 4416 5287 4424 5344
rect 4456 5307 4464 5344
rect 4336 5076 4364 5084
rect 4376 5076 4384 5213
rect 4416 5147 4424 5273
rect 4413 5080 4427 5093
rect 4416 5076 4424 5080
rect 4196 4967 4204 5033
rect 4196 4887 4204 4913
rect 4036 4856 4044 4860
rect 4180 4866 4200 4867
rect 4180 4863 4193 4866
rect 4176 4855 4193 4863
rect 4076 4827 4084 4854
rect 4180 4853 4193 4855
rect 4216 4847 4224 4993
rect 4276 4987 4284 5044
rect 4316 4967 4324 5033
rect 4116 4820 4124 4824
rect 3956 4704 3964 4753
rect 3936 4696 3964 4704
rect 3876 4576 3904 4584
rect 3876 4556 3884 4576
rect 3776 4136 3804 4144
rect 3756 4036 3764 4073
rect 3796 4004 3804 4136
rect 3816 4127 3824 4554
rect 3836 4347 3844 4513
rect 3856 4487 3864 4524
rect 3896 4487 3904 4524
rect 3936 4467 3944 4696
rect 3996 4667 4004 4693
rect 4016 4568 4024 4812
rect 3956 4516 3984 4524
rect 3956 4407 3964 4516
rect 3860 4304 3873 4307
rect 3856 4296 3873 4304
rect 3860 4293 3873 4296
rect 3836 4104 3844 4293
rect 3916 4267 3924 4304
rect 3776 3996 3804 4004
rect 3816 4096 3844 4104
rect 3656 3780 3664 3784
rect 3653 3767 3667 3780
rect 3336 3528 3344 3613
rect 3376 3528 3384 3613
rect 3656 3607 3664 3753
rect 3696 3707 3704 3784
rect 3316 3480 3324 3484
rect 3296 3387 3304 3473
rect 3313 3467 3327 3480
rect 3196 3047 3204 3313
rect 3216 3266 3224 3333
rect 3256 3296 3264 3373
rect 3236 3067 3244 3233
rect 3256 3127 3264 3173
rect 3176 3007 3184 3033
rect 3047 2956 3064 2964
rect 2896 2747 2904 2813
rect 2976 2776 2984 2813
rect 3036 2787 3044 2932
rect 2616 2696 2644 2704
rect 2753 2724 2767 2733
rect 2653 2704 2667 2713
rect 2736 2720 2767 2724
rect 2736 2716 2764 2720
rect 2653 2700 2684 2704
rect 2656 2696 2684 2700
rect 2516 2476 2524 2512
rect 2556 2476 2564 2613
rect 2476 2327 2484 2433
rect 2496 2387 2504 2444
rect 2596 2367 2604 2633
rect 2616 2488 2624 2696
rect 2636 2507 2644 2673
rect 2676 2644 2684 2696
rect 2736 2684 2744 2716
rect 2716 2676 2744 2684
rect 2716 2667 2724 2676
rect 2707 2656 2724 2667
rect 2707 2653 2720 2656
rect 2676 2636 2713 2644
rect 2696 2587 2704 2613
rect 2756 2604 2764 2693
rect 2736 2596 2764 2604
rect 2676 2507 2684 2553
rect 2676 2494 2693 2507
rect 2636 2476 2644 2493
rect 2716 2487 2724 2513
rect 2700 2444 2713 2447
rect 2656 2367 2664 2444
rect 2696 2433 2713 2444
rect 2496 2256 2504 2352
rect 2436 2147 2444 2212
rect 2476 2127 2484 2224
rect 2416 1956 2424 2113
rect 2516 2067 2524 2113
rect 2536 2087 2544 2224
rect 2556 2107 2564 2193
rect 2547 2076 2564 2084
rect 2453 2047 2467 2053
rect 2447 2040 2467 2047
rect 2447 2036 2464 2040
rect 2447 2033 2460 2036
rect 2433 1987 2447 1993
rect 2456 1956 2464 2013
rect 2527 1993 2533 2007
rect 2476 1967 2484 1993
rect 2556 1984 2564 2076
rect 2596 1987 2604 2313
rect 2676 2256 2684 2333
rect 2696 2267 2704 2433
rect 2713 2407 2727 2412
rect 2716 2247 2724 2293
rect 2716 2184 2724 2212
rect 2736 2207 2744 2596
rect 2756 2445 2764 2493
rect 2776 2487 2784 2732
rect 2816 2707 2824 2744
rect 2796 2587 2804 2653
rect 2856 2607 2864 2732
rect 2916 2724 2924 2773
rect 2896 2716 2924 2724
rect 2896 2667 2904 2716
rect 2956 2707 2964 2744
rect 2836 2476 2844 2513
rect 2856 2507 2864 2553
rect 2916 2487 2924 2693
rect 2956 2667 2964 2693
rect 2936 2467 2944 2573
rect 2976 2504 2984 2673
rect 3036 2507 3044 2733
rect 3056 2587 3064 2956
rect 3116 2927 3124 2964
rect 3156 2947 3164 2994
rect 3276 3007 3284 3193
rect 3296 2967 3304 3233
rect 3316 3167 3324 3264
rect 3356 3027 3364 3484
rect 3436 3484 3444 3514
rect 3576 3486 3584 3553
rect 3736 3547 3744 3833
rect 3776 3827 3784 3996
rect 3816 3827 3824 4096
rect 3916 4036 3924 4073
rect 3956 4047 3964 4353
rect 3976 4267 3984 4413
rect 3996 4306 4004 4493
rect 4016 4447 4024 4473
rect 4056 4427 4064 4713
rect 4076 4367 4084 4773
rect 4096 4667 4104 4813
rect 4113 4807 4127 4820
rect 4156 4556 4164 4613
rect 4176 4567 4184 4793
rect 4196 4727 4204 4813
rect 4216 4707 4224 4833
rect 4236 4747 4244 4953
rect 4296 4856 4304 4933
rect 4336 4867 4344 5076
rect 4276 4747 4284 4824
rect 4336 4787 4344 4813
rect 4196 4526 4204 4653
rect 4276 4627 4284 4733
rect 4356 4707 4364 5033
rect 4376 4767 4384 4973
rect 4396 4907 4404 5044
rect 4436 4868 4444 5013
rect 4456 4987 4464 5213
rect 4476 4887 4484 5253
rect 4496 5087 4504 5233
rect 4516 5088 4524 5193
rect 4556 5127 4564 5173
rect 4576 5167 4584 5344
rect 4496 4867 4504 5033
rect 4480 4824 4493 4827
rect 4476 4816 4493 4824
rect 4480 4813 4493 4816
rect 4456 4787 4464 4813
rect 4516 4767 4524 4873
rect 4536 4867 4544 5033
rect 4556 4967 4564 5044
rect 4556 4907 4564 4953
rect 4616 4947 4624 5413
rect 4676 5376 4684 5456
rect 4756 5444 4764 5564
rect 4796 5507 4804 5564
rect 4776 5467 4784 5493
rect 4816 5444 4824 5553
rect 4836 5527 4844 5633
rect 4856 5507 4864 5693
rect 4916 5628 4924 5933
rect 4936 5687 4944 5893
rect 4956 5864 4964 5913
rect 4956 5856 5004 5864
rect 4876 5467 4884 5613
rect 4956 5596 4964 5733
rect 4756 5436 4824 5444
rect 4716 5384 4724 5433
rect 4856 5427 4864 5453
rect 4716 5376 4744 5384
rect 4696 5340 4704 5344
rect 4693 5327 4707 5340
rect 4636 5027 4644 5153
rect 4656 5087 4664 5213
rect 4716 5104 4724 5313
rect 4736 5227 4744 5376
rect 4756 5327 4764 5413
rect 4836 5376 4844 5413
rect 4787 5313 4793 5327
rect 4716 5096 4744 5104
rect 4736 5087 4744 5096
rect 4736 5076 4753 5087
rect 4740 5073 4753 5076
rect 4656 4924 4664 5033
rect 4676 4987 4684 5044
rect 4776 5027 4784 5173
rect 4816 5107 4824 5344
rect 4876 5307 4884 5374
rect 4896 5267 4904 5553
rect 4916 5207 4924 5473
rect 4976 5464 4984 5564
rect 5016 5507 5024 5853
rect 5076 5687 5084 6233
rect 5096 5847 5104 6053
rect 5116 6047 5124 6072
rect 5156 6027 5164 6084
rect 5173 6067 5187 6073
rect 5196 6067 5204 6253
rect 5216 6087 5224 6133
rect 5276 6116 5284 6153
rect 5256 6080 5264 6084
rect 5253 6067 5267 6080
rect 5216 6007 5224 6033
rect 5116 5907 5124 5953
rect 5216 5907 5224 5993
rect 5256 5896 5264 5933
rect 5296 5907 5304 6073
rect 5176 5856 5204 5864
rect 5053 5600 5067 5613
rect 5056 5596 5064 5600
rect 5096 5596 5104 5753
rect 5116 5647 5124 5773
rect 5156 5747 5164 5773
rect 5136 5596 5144 5693
rect 5156 5607 5164 5653
rect 4976 5456 5004 5464
rect 4996 5387 5004 5456
rect 5013 5404 5027 5413
rect 5036 5404 5044 5513
rect 5013 5400 5044 5404
rect 5016 5396 5044 5400
rect 5016 5376 5024 5396
rect 4976 5340 4984 5344
rect 4973 5327 4987 5340
rect 5036 5336 5064 5344
rect 4976 5227 4984 5253
rect 4996 5167 5004 5333
rect 4836 5076 4844 5113
rect 4733 5004 4747 5013
rect 4716 5000 4747 5004
rect 4716 4996 4744 5000
rect 4716 4984 4724 4996
rect 4696 4976 4724 4984
rect 4656 4916 4684 4924
rect 4636 4887 4644 4913
rect 4536 4767 4544 4813
rect 4336 4647 4344 4673
rect 4316 4556 4364 4564
rect 4136 4520 4144 4524
rect 4133 4507 4147 4520
rect 4146 4500 4147 4507
rect 4156 4336 4164 4493
rect 4296 4487 4304 4554
rect 4316 4487 4324 4556
rect 4016 4087 4024 4153
rect 4076 4127 4084 4304
rect 3836 4007 3844 4034
rect 3836 3816 3844 3933
rect 3856 3827 3864 3973
rect 3896 3927 3904 4004
rect 3936 3927 3944 4004
rect 3756 3747 3764 3813
rect 3796 3764 3804 3772
rect 3776 3756 3804 3764
rect 3696 3486 3704 3533
rect 3776 3527 3784 3756
rect 3856 3724 3864 3773
rect 3836 3716 3864 3724
rect 3436 3476 3464 3484
rect 3376 3307 3384 3453
rect 3396 3347 3404 3473
rect 3436 3327 3444 3413
rect 3456 3296 3464 3476
rect 3476 3307 3484 3393
rect 3496 3266 3504 3313
rect 3376 3207 3384 3253
rect 3396 3167 3404 3264
rect 3516 3227 3524 3484
rect 3576 3447 3584 3472
rect 3736 3447 3744 3484
rect 3553 3300 3567 3313
rect 3556 3296 3564 3300
rect 3616 3267 3624 3313
rect 3693 3300 3707 3313
rect 3733 3300 3747 3313
rect 3696 3296 3704 3300
rect 3736 3296 3744 3300
rect 3776 3266 3784 3473
rect 3796 3347 3804 3513
rect 3816 3304 3824 3513
rect 3836 3427 3844 3716
rect 3876 3547 3884 3853
rect 3976 3827 3984 4073
rect 4016 4036 4024 4073
rect 4053 4040 4067 4053
rect 4073 4047 4087 4053
rect 4056 4036 4064 4040
rect 4096 3987 4104 4253
rect 4136 4207 4144 4293
rect 3996 3807 4004 3973
rect 4076 3816 4084 3853
rect 4116 3847 4124 4073
rect 4136 4047 4144 4193
rect 4176 4127 4184 4304
rect 4196 4187 4204 4293
rect 4216 4067 4224 4473
rect 4376 4447 4384 4512
rect 4236 4167 4244 4413
rect 4296 4336 4304 4373
rect 4256 4247 4264 4304
rect 4316 4127 4324 4284
rect 4153 4040 4167 4053
rect 4156 4036 4164 4040
rect 4236 4047 4244 4113
rect 4300 4064 4313 4067
rect 4296 4053 4313 4064
rect 4296 4036 4304 4053
rect 4136 3824 4144 3993
rect 4176 3907 4184 4004
rect 4256 4004 4264 4034
rect 4356 4006 4364 4093
rect 4236 3996 4264 4004
rect 4216 3927 4224 3992
rect 4116 3816 4144 3824
rect 3896 3687 3904 3773
rect 3916 3664 3924 3784
rect 4016 3784 4024 3816
rect 4216 3787 4224 3892
rect 4016 3776 4044 3784
rect 3956 3764 3964 3772
rect 3896 3656 3924 3664
rect 3936 3756 3964 3764
rect 3896 3647 3904 3656
rect 3896 3524 3904 3633
rect 3936 3527 3944 3756
rect 3996 3704 4004 3772
rect 3996 3696 4013 3704
rect 3876 3516 3904 3524
rect 4016 3507 4024 3693
rect 3916 3407 3924 3484
rect 4036 3467 4044 3776
rect 4056 3687 4064 3784
rect 4096 3727 4104 3784
rect 4073 3520 4087 3533
rect 4156 3524 4164 3653
rect 4076 3516 4084 3520
rect 4136 3516 4164 3524
rect 3796 3296 3824 3304
rect 3076 2527 3084 2913
rect 3176 2907 3184 2953
rect 3173 2820 3187 2833
rect 3176 2816 3184 2820
rect 3236 2759 3244 2933
rect 3096 2667 3104 2753
rect 3233 2746 3247 2753
rect 3256 2684 3264 2753
rect 3276 2687 3284 2953
rect 3296 2787 3304 2893
rect 3316 2807 3324 3013
rect 3356 2867 3364 2964
rect 3396 2867 3404 2964
rect 3396 2787 3404 2853
rect 3236 2676 3264 2684
rect 3087 2516 3104 2524
rect 2956 2496 2984 2504
rect 2813 2427 2827 2433
rect 2856 2387 2864 2444
rect 2913 2427 2927 2433
rect 2836 2327 2844 2353
rect 2816 2256 2824 2293
rect 2936 2268 2944 2453
rect 2767 2224 2780 2227
rect 2767 2216 2784 2224
rect 2767 2213 2780 2216
rect 2716 2176 2744 2184
rect 2513 1968 2527 1972
rect 2496 1956 2513 1964
rect 2496 1926 2504 1956
rect 2536 1976 2564 1984
rect 2536 1956 2544 1976
rect 2396 1920 2404 1924
rect 2393 1907 2407 1920
rect 2556 1867 2564 1924
rect 2376 1706 2384 1833
rect 2396 1767 2404 1813
rect 2416 1787 2424 1813
rect 2416 1736 2424 1773
rect 2456 1736 2464 1853
rect 2436 1684 2444 1704
rect 2436 1676 2464 1684
rect 2347 1556 2364 1564
rect 2176 1240 2204 1244
rect 2173 1236 2204 1240
rect 2173 1227 2187 1236
rect 2186 1220 2187 1227
rect 2233 1220 2247 1233
rect 2276 1227 2284 1353
rect 2316 1307 2324 1353
rect 2336 1264 2344 1553
rect 2416 1436 2424 1533
rect 2436 1487 2444 1513
rect 2316 1256 2344 1264
rect 2236 1216 2244 1220
rect 2296 1186 2304 1213
rect 2076 1180 2084 1184
rect 2036 1087 2044 1173
rect 2073 1167 2087 1180
rect 1936 916 1944 920
rect 1996 886 2004 953
rect 2036 928 2044 1073
rect 2076 916 2084 993
rect 2096 944 2104 1033
rect 2127 953 2133 967
rect 2096 936 2124 944
rect 2116 916 2124 936
rect 1956 787 1964 813
rect 1946 773 1947 780
rect 1933 764 1947 773
rect 1933 760 1964 764
rect 1936 756 1964 760
rect 1833 700 1847 713
rect 1836 696 1844 700
rect 1536 660 1544 664
rect 1533 647 1547 660
rect 1496 607 1504 633
rect 1636 627 1644 664
rect 1673 647 1687 652
rect 1756 647 1764 693
rect 1773 647 1787 653
rect 1396 347 1404 413
rect 1476 267 1484 324
rect 1256 140 1264 144
rect 1253 127 1267 140
rect 976 116 993 127
rect 980 113 993 116
rect 1240 106 1260 107
rect 1213 84 1227 93
rect 1247 93 1253 106
rect 1276 84 1284 113
rect 1213 80 1284 84
rect 1216 76 1284 80
rect 1336 47 1344 174
rect 1476 146 1484 173
rect 1376 140 1384 144
rect 1373 127 1387 140
rect 1496 87 1504 293
rect 1516 146 1524 233
rect 1536 187 1544 273
rect 1576 176 1584 433
rect 1616 407 1624 553
rect 1656 408 1664 573
rect 1816 547 1824 664
rect 1607 396 1624 407
rect 1607 393 1620 396
rect 1616 187 1624 233
rect 1636 227 1644 364
rect 1696 347 1704 493
rect 1856 487 1864 652
rect 1896 587 1904 713
rect 1916 707 1924 753
rect 1956 696 1964 756
rect 1996 696 2004 733
rect 2016 704 2024 913
rect 2156 886 2164 973
rect 2173 967 2187 973
rect 2056 880 2064 884
rect 2053 867 2067 880
rect 2076 707 2084 793
rect 2016 696 2044 704
rect 1976 607 1984 664
rect 2016 547 2024 653
rect 2036 567 2044 696
rect 2156 696 2164 793
rect 2196 787 2204 993
rect 2296 927 2304 1172
rect 2316 1167 2324 1256
rect 2396 1247 2404 1404
rect 2336 1107 2344 1233
rect 2416 1216 2424 1373
rect 2456 1244 2464 1676
rect 2476 1467 2484 1693
rect 2496 1667 2504 1793
rect 2616 1706 2624 2153
rect 2636 1807 2644 2173
rect 2676 1968 2684 2093
rect 2716 1956 2724 2013
rect 2736 1967 2744 2176
rect 2756 1947 2764 2073
rect 2776 1924 2784 2193
rect 2956 2147 2964 2496
rect 3047 2496 3064 2504
rect 3056 2476 3064 2496
rect 3096 2487 3104 2516
rect 2976 2407 2984 2473
rect 3036 2440 3044 2444
rect 2976 2167 2984 2353
rect 2996 2327 3004 2433
rect 3033 2427 3047 2440
rect 3036 2256 3044 2313
rect 3076 2268 3084 2411
rect 3116 2367 3124 2593
rect 3147 2444 3160 2447
rect 3147 2436 3164 2444
rect 3147 2433 3160 2436
rect 3136 2256 3144 2373
rect 3216 2267 3224 2573
rect 2996 2227 3004 2254
rect 3200 2224 3213 2227
rect 3056 2220 3064 2224
rect 3156 2220 3164 2224
rect 3053 2207 3067 2220
rect 3153 2207 3167 2220
rect 3196 2216 3213 2224
rect 3200 2213 3213 2216
rect 2807 1964 2820 1967
rect 2807 1956 2824 1964
rect 2853 1960 2867 1973
rect 2856 1956 2864 1960
rect 2807 1953 2820 1956
rect 3116 1956 3164 1964
rect 2636 1707 2644 1753
rect 2656 1747 2664 1913
rect 2696 1807 2704 1924
rect 2756 1916 2784 1924
rect 2716 1787 2724 1833
rect 2756 1827 2764 1916
rect 2496 1467 2504 1653
rect 2576 1647 2584 1704
rect 2616 1647 2624 1692
rect 2776 1687 2784 1893
rect 2796 1807 2804 1913
rect 2836 1867 2844 1924
rect 2876 1920 2884 1924
rect 2873 1907 2887 1920
rect 2916 1907 2924 1954
rect 2986 1891 2987 1900
rect 2973 1887 2987 1891
rect 2856 1736 2864 1773
rect 2573 1440 2587 1453
rect 2633 1440 2647 1453
rect 2676 1448 2684 1653
rect 2576 1436 2584 1440
rect 2636 1436 2644 1440
rect 2476 1267 2484 1432
rect 2516 1247 2524 1353
rect 2456 1236 2484 1244
rect 2276 916 2293 924
rect 2336 916 2344 1072
rect 2356 1047 2364 1173
rect 2476 1184 2484 1236
rect 2513 1220 2527 1233
rect 2516 1216 2524 1220
rect 2616 1184 2624 1353
rect 2656 1307 2664 1404
rect 2736 1367 2744 1671
rect 2816 1647 2824 1692
rect 2876 1547 2884 1704
rect 2833 1440 2847 1453
rect 2836 1436 2844 1440
rect 2756 1387 2764 1434
rect 2740 1344 2753 1347
rect 2736 1333 2753 1344
rect 2676 1216 2684 1313
rect 2713 1220 2727 1233
rect 2736 1227 2744 1333
rect 2796 1307 2804 1373
rect 2816 1347 2824 1404
rect 2856 1347 2864 1404
rect 2716 1216 2724 1220
rect 2456 1176 2484 1184
rect 2536 1180 2544 1184
rect 2576 1180 2584 1184
rect 2376 1067 2384 1093
rect 2456 1027 2464 1176
rect 2533 1167 2547 1180
rect 2573 1167 2587 1180
rect 2596 1176 2624 1184
rect 2256 827 2264 884
rect 2256 747 2264 813
rect 1676 247 1684 293
rect 1716 287 1724 453
rect 1816 396 1824 453
rect 1976 396 1984 433
rect 1736 347 1744 394
rect 1796 360 1804 364
rect 1793 347 1807 360
rect 1996 327 2004 364
rect 2036 347 2044 513
rect 2056 408 2064 693
rect 2096 660 2104 664
rect 2093 647 2107 660
rect 2136 607 2144 664
rect 2113 400 2127 413
rect 2176 404 2184 653
rect 2196 647 2204 733
rect 2216 666 2224 713
rect 2247 704 2260 707
rect 2247 696 2264 704
rect 2296 696 2304 733
rect 2247 693 2260 696
rect 2276 427 2284 553
rect 2356 547 2364 733
rect 2376 707 2384 753
rect 2396 696 2404 793
rect 2436 784 2444 913
rect 2456 887 2464 953
rect 2516 916 2524 1053
rect 2533 947 2547 953
rect 2556 928 2564 973
rect 2416 776 2444 784
rect 2416 727 2424 776
rect 2436 696 2444 733
rect 2476 707 2484 813
rect 2416 627 2424 664
rect 2496 627 2504 884
rect 2596 867 2604 1176
rect 2636 1067 2644 1213
rect 2633 920 2647 933
rect 2636 916 2644 920
rect 2676 916 2684 1053
rect 2696 987 2704 1184
rect 2756 1167 2764 1293
rect 2756 886 2764 1153
rect 2776 924 2784 1273
rect 2876 1264 2884 1393
rect 2896 1387 2904 1692
rect 2916 1607 2924 1833
rect 2996 1787 3004 1893
rect 3016 1847 3024 1954
rect 3156 1927 3164 1956
rect 3056 1907 3064 1924
rect 3047 1896 3064 1907
rect 3047 1893 3060 1896
rect 2996 1736 3004 1773
rect 2936 1647 2944 1733
rect 2976 1567 2984 1704
rect 2927 1444 2940 1447
rect 2927 1436 2944 1444
rect 2973 1440 2987 1453
rect 3036 1447 3044 1853
rect 3076 1736 3084 1793
rect 3096 1767 3104 1924
rect 3116 1787 3124 1873
rect 3116 1736 3124 1773
rect 3156 1667 3164 1873
rect 3076 1467 3084 1613
rect 2976 1436 2984 1440
rect 2927 1433 2940 1436
rect 3073 1440 3087 1453
rect 3076 1436 3084 1440
rect 3176 1447 3184 2173
rect 3216 2107 3224 2213
rect 3236 2187 3244 2676
rect 3276 2547 3284 2673
rect 3296 2607 3304 2733
rect 3316 2727 3324 2744
rect 3316 2647 3324 2713
rect 3316 2544 3324 2573
rect 3336 2567 3344 2733
rect 3376 2647 3384 2744
rect 3316 2536 3344 2544
rect 3293 2480 3307 2493
rect 3336 2488 3344 2536
rect 3296 2476 3304 2480
rect 3356 2487 3364 2533
rect 3316 2440 3324 2444
rect 3313 2427 3327 2440
rect 3376 2327 3384 2593
rect 3396 2488 3404 2733
rect 3416 2547 3424 2793
rect 3436 2787 3444 3193
rect 3456 2966 3464 3033
rect 3536 2996 3544 3053
rect 3596 2966 3604 3093
rect 3656 2996 3664 3233
rect 3716 3127 3724 3264
rect 3796 3107 3804 3296
rect 3876 3296 3884 3333
rect 3936 3266 3944 3313
rect 3996 3296 4004 3353
rect 4056 3307 4064 3413
rect 3976 3260 3984 3264
rect 3973 3247 3987 3260
rect 3873 3224 3887 3233
rect 3847 3220 3887 3224
rect 3993 3227 4007 3233
rect 3847 3216 3884 3220
rect 3836 3147 3844 3173
rect 3816 3008 3824 3073
rect 3456 2776 3464 2853
rect 3476 2740 3484 2744
rect 3473 2727 3487 2740
rect 3556 2507 3564 2964
rect 3576 2607 3584 2933
rect 3676 2867 3684 2964
rect 3736 2956 3753 2964
rect 3736 2907 3744 2956
rect 3816 2887 3824 2994
rect 3836 2964 3844 3133
rect 4056 3127 4064 3253
rect 4076 3187 4084 3453
rect 4176 3327 4184 3573
rect 4216 3387 4224 3752
rect 4236 3727 4244 3996
rect 4256 3827 4264 3973
rect 4336 3776 4364 3784
rect 4236 3527 4244 3713
rect 4356 3667 4364 3776
rect 4256 3516 4264 3613
rect 4336 3484 4344 3633
rect 4376 3587 4384 4073
rect 4396 4047 4404 4353
rect 4416 4087 4424 4753
rect 4476 4607 4484 4753
rect 4496 4667 4504 4713
rect 4456 4568 4464 4593
rect 4496 4556 4504 4653
rect 4516 4587 4524 4713
rect 4536 4627 4544 4753
rect 4476 4427 4484 4524
rect 4516 4516 4544 4524
rect 4456 4347 4464 4393
rect 4447 4336 4464 4347
rect 4496 4336 4504 4453
rect 4516 4387 4524 4433
rect 4536 4387 4544 4516
rect 4556 4367 4564 4793
rect 4576 4787 4584 4824
rect 4616 4687 4624 4824
rect 4636 4727 4644 4813
rect 4656 4767 4664 4893
rect 4676 4867 4684 4916
rect 4696 4887 4704 4976
rect 4716 4887 4724 4953
rect 4736 4947 4744 4973
rect 4776 4947 4784 5013
rect 4716 4874 4733 4887
rect 4796 4867 4804 5033
rect 4856 5007 4864 5044
rect 4796 4856 4813 4867
rect 4800 4853 4813 4856
rect 4676 4787 4684 4832
rect 4736 4804 4744 4824
rect 4716 4796 4744 4804
rect 4576 4567 4584 4593
rect 4616 4556 4624 4652
rect 4653 4627 4667 4633
rect 4636 4587 4644 4613
rect 4660 4564 4673 4567
rect 4656 4556 4673 4564
rect 4660 4553 4673 4556
rect 4587 4524 4600 4527
rect 4587 4516 4604 4524
rect 4587 4513 4600 4516
rect 4447 4333 4460 4336
rect 4556 4307 4564 4332
rect 4576 4307 4584 4473
rect 4596 4447 4604 4493
rect 4616 4427 4624 4473
rect 4636 4447 4644 4524
rect 4696 4526 4704 4713
rect 4716 4707 4724 4796
rect 4736 4627 4744 4693
rect 4816 4687 4824 4813
rect 4836 4624 4844 4973
rect 4853 4864 4867 4873
rect 4916 4867 4924 5093
rect 4936 4907 4944 5153
rect 4993 5104 5007 5113
rect 4976 5100 5007 5104
rect 4976 5096 5004 5100
rect 4976 5076 4984 5096
rect 5016 5076 5024 5313
rect 5036 5187 5044 5293
rect 5056 5267 5064 5336
rect 5076 5287 5084 5453
rect 5136 5387 5144 5533
rect 5156 5447 5164 5493
rect 5156 5376 5164 5433
rect 5176 5387 5184 5833
rect 5196 5827 5204 5856
rect 5296 5827 5304 5853
rect 5196 5767 5204 5813
rect 5196 5547 5204 5673
rect 5236 5627 5244 5713
rect 5256 5596 5264 5693
rect 5276 5607 5284 5653
rect 5296 5647 5304 5733
rect 5316 5707 5324 5894
rect 5316 5587 5324 5693
rect 5227 5556 5244 5564
rect 5196 5487 5204 5512
rect 4853 4860 4884 4864
rect 4856 4856 4884 4860
rect 4876 4687 4884 4773
rect 4896 4767 4904 4812
rect 4816 4620 4844 4624
rect 4813 4616 4844 4620
rect 4813 4607 4827 4616
rect 4593 4367 4607 4373
rect 4616 4344 4624 4413
rect 4636 4407 4644 4433
rect 4656 4427 4664 4493
rect 4676 4487 4684 4513
rect 4696 4367 4704 4512
rect 4673 4348 4687 4353
rect 4596 4336 4624 4344
rect 4476 4247 4484 4304
rect 4516 4300 4524 4304
rect 4513 4287 4527 4300
rect 4596 4287 4604 4336
rect 4716 4347 4724 4573
rect 4736 4547 4744 4592
rect 4736 4427 4744 4533
rect 4796 4476 4824 4484
rect 4656 4300 4664 4304
rect 4413 4040 4427 4052
rect 4416 4036 4424 4040
rect 4456 4036 4464 4113
rect 4516 4004 4524 4213
rect 4556 4036 4564 4113
rect 4616 4047 4624 4293
rect 4653 4287 4667 4300
rect 4636 4147 4644 4273
rect 4396 3767 4404 3993
rect 4416 3828 4424 3933
rect 4436 3907 4444 4004
rect 4476 4000 4504 4004
rect 4476 3996 4507 4000
rect 4516 3996 4544 4004
rect 4493 3987 4507 3996
rect 4416 3727 4424 3814
rect 4536 3784 4544 3996
rect 4567 3980 4604 3984
rect 4567 3976 4607 3980
rect 4593 3967 4607 3976
rect 4556 3827 4564 3952
rect 4616 3887 4624 3993
rect 4636 3987 4644 4112
rect 4656 4107 4664 4273
rect 4676 4127 4684 4273
rect 4736 4167 4744 4392
rect 4756 4287 4764 4453
rect 4776 4407 4784 4473
rect 4796 4384 4804 4476
rect 4816 4387 4824 4453
rect 4776 4380 4804 4384
rect 4773 4376 4804 4380
rect 4773 4367 4787 4376
rect 4896 4348 4904 4573
rect 4936 4556 4944 4853
rect 4956 4587 4964 4973
rect 4996 4868 5004 4933
rect 5036 4927 5044 5033
rect 5056 5027 5064 5213
rect 5076 4867 5084 5193
rect 5096 5087 5104 5333
rect 5116 5167 5124 5344
rect 5136 5104 5144 5233
rect 5196 5127 5204 5393
rect 5216 5387 5224 5552
rect 5247 5544 5260 5547
rect 5247 5533 5264 5544
rect 5236 5407 5244 5453
rect 5256 5427 5264 5533
rect 5233 5380 5247 5393
rect 5273 5380 5287 5393
rect 5236 5376 5244 5380
rect 5276 5376 5284 5380
rect 5187 5116 5204 5127
rect 5187 5113 5200 5116
rect 5127 5096 5144 5104
rect 5116 5076 5124 5093
rect 5153 5080 5167 5093
rect 5193 5087 5207 5093
rect 5156 5076 5164 5080
rect 4976 4607 4984 4813
rect 4996 4584 5004 4793
rect 5016 4727 5024 4824
rect 5056 4820 5064 4824
rect 5053 4807 5067 4820
rect 5076 4664 5084 4813
rect 5056 4656 5084 4664
rect 5056 4587 5064 4656
rect 4976 4576 5004 4584
rect 4976 4556 4984 4576
rect 5076 4567 5084 4633
rect 5096 4627 5104 5033
rect 5136 4967 5144 5044
rect 5116 4826 5124 4913
rect 5156 4867 5164 5013
rect 5176 4887 5184 5032
rect 5216 4987 5224 5273
rect 5316 5227 5324 5493
rect 5336 5467 5344 6193
rect 5593 6147 5607 6153
rect 5487 6136 5513 6144
rect 5433 6120 5447 6133
rect 5436 6116 5444 6120
rect 5553 6120 5567 6133
rect 5593 6127 5607 6133
rect 5556 6116 5564 6120
rect 5376 6007 5384 6073
rect 5416 6047 5424 6084
rect 5476 6027 5484 6073
rect 5416 5896 5424 5993
rect 5436 5860 5444 5864
rect 5433 5847 5447 5860
rect 5476 5827 5484 5894
rect 5456 5707 5464 5773
rect 5476 5727 5484 5813
rect 5496 5587 5504 5933
rect 5536 5908 5544 5953
rect 5516 5767 5524 5833
rect 5616 5704 5624 6173
rect 5636 5907 5644 6153
rect 5656 6047 5664 6233
rect 5816 6147 5824 6304
rect 5856 6267 5864 6304
rect 5896 6296 5924 6304
rect 5693 6120 5707 6133
rect 5696 6116 5704 6120
rect 5836 6116 5844 6173
rect 5756 6080 5764 6084
rect 5753 6067 5767 6080
rect 5736 5987 5744 6033
rect 5796 6007 5804 6093
rect 5656 5896 5664 5953
rect 5696 5896 5704 5933
rect 5636 5724 5644 5853
rect 5676 5807 5684 5852
rect 5636 5716 5664 5724
rect 5616 5696 5644 5704
rect 5416 5520 5424 5524
rect 5413 5507 5427 5520
rect 5336 5347 5344 5413
rect 5356 5387 5364 5413
rect 5393 5380 5407 5393
rect 5436 5388 5444 5513
rect 5496 5504 5504 5552
rect 5516 5547 5524 5593
rect 5496 5496 5524 5504
rect 5396 5376 5404 5380
rect 5496 5376 5504 5453
rect 5516 5404 5524 5496
rect 5536 5427 5544 5693
rect 5616 5607 5624 5673
rect 5516 5396 5544 5404
rect 5536 5376 5544 5396
rect 5576 5387 5584 5533
rect 5416 5287 5424 5332
rect 5416 5247 5424 5273
rect 5256 5088 5264 5193
rect 5376 5187 5384 5213
rect 5396 5087 5404 5173
rect 5276 5024 5284 5044
rect 5267 5016 5284 5024
rect 5233 4860 5247 4873
rect 5256 4867 5264 5013
rect 5316 5007 5324 5044
rect 5336 4987 5344 5033
rect 5356 4967 5364 5074
rect 5376 4987 5384 5074
rect 5456 5087 5464 5153
rect 5333 4887 5347 4893
rect 5236 4856 5244 4860
rect 5113 4807 5127 4812
rect 5136 4787 5144 4853
rect 5156 4647 5164 4813
rect 5216 4747 5224 4824
rect 5276 4826 5284 4873
rect 5336 4856 5344 4873
rect 5376 4856 5384 4933
rect 5416 4826 5424 4993
rect 5176 4667 5184 4733
rect 5216 4647 5224 4693
rect 4916 4447 4924 4513
rect 4996 4520 5004 4524
rect 4993 4507 5007 4520
rect 4916 4336 4924 4393
rect 4756 4006 4764 4033
rect 4656 3996 4684 4004
rect 4456 3780 4464 3784
rect 4453 3767 4467 3780
rect 4516 3776 4544 3784
rect 3876 2996 3884 3033
rect 3836 2956 3864 2964
rect 3407 2444 3420 2447
rect 3407 2436 3424 2444
rect 3407 2433 3420 2436
rect 3276 2207 3284 2253
rect 3216 1956 3224 2013
rect 3256 1968 3264 2153
rect 3316 2127 3324 2224
rect 3396 2067 3404 2254
rect 3416 2007 3424 2273
rect 3476 2267 3484 2433
rect 3496 2287 3504 2493
rect 3616 2476 3624 2673
rect 3636 2647 3644 2744
rect 3516 2427 3524 2453
rect 3556 2407 3564 2444
rect 3516 2264 3524 2313
rect 3496 2256 3524 2264
rect 3456 2087 3464 2224
rect 3456 2024 3464 2073
rect 3456 2016 3484 2024
rect 3356 1968 3364 1993
rect 3376 1956 3384 1993
rect 3196 1467 3204 1912
rect 3296 1907 3304 1954
rect 3296 1867 3304 1893
rect 3396 1827 3404 1924
rect 3256 1748 3264 1773
rect 3336 1707 3344 1793
rect 3456 1747 3464 1993
rect 3236 1627 3244 1704
rect 3476 1706 3484 2016
rect 3516 2007 3524 2213
rect 3536 2207 3544 2293
rect 3596 2287 3604 2444
rect 3656 2347 3664 2493
rect 3676 2447 3684 2744
rect 3696 2647 3704 2732
rect 3716 2484 3724 2773
rect 3736 2508 3744 2853
rect 3756 2687 3764 2813
rect 3776 2787 3784 2873
rect 3756 2547 3764 2593
rect 3696 2476 3724 2484
rect 3696 2344 3704 2476
rect 3776 2476 3784 2553
rect 3836 2487 3844 2732
rect 3856 2707 3864 2956
rect 3936 2776 3944 2813
rect 3976 2807 3984 2996
rect 3996 2967 4004 3053
rect 4016 3007 4024 3093
rect 4096 3007 4104 3313
rect 4296 3308 4304 3484
rect 4336 3476 4364 3484
rect 4356 3307 4364 3476
rect 4416 3480 4424 3484
rect 4116 3227 4124 3252
rect 3996 2784 4004 2893
rect 3976 2776 4004 2784
rect 3876 2747 3884 2774
rect 3836 2347 3844 2473
rect 3696 2336 3724 2344
rect 3556 2047 3564 2273
rect 3616 2268 3624 2333
rect 3576 2107 3584 2193
rect 3596 2187 3604 2224
rect 3716 2167 3724 2336
rect 3516 1956 3524 1993
rect 3553 1960 3567 1973
rect 3556 1956 3564 1960
rect 3596 1956 3604 2073
rect 3636 1926 3644 1973
rect 3536 1887 3544 1912
rect 3576 1867 3584 1924
rect 3587 1856 3604 1864
rect 3493 1748 3507 1753
rect 3573 1747 3587 1753
rect 3256 1507 3264 1593
rect 2867 1256 2884 1264
rect 2856 1216 2864 1253
rect 2916 1228 2924 1393
rect 3007 1396 3024 1404
rect 2956 1216 2964 1333
rect 2916 1186 2924 1214
rect 2836 1180 2844 1184
rect 2796 1027 2804 1173
rect 2833 1167 2847 1180
rect 3016 1167 3024 1396
rect 3096 1367 3104 1404
rect 3036 1227 3044 1253
rect 3096 1247 3104 1293
rect 3136 1224 3144 1353
rect 3156 1347 3164 1434
rect 3193 1440 3207 1453
rect 3196 1436 3204 1440
rect 3276 1447 3284 1513
rect 3296 1407 3304 1453
rect 3336 1447 3344 1672
rect 3416 1567 3424 1693
rect 3436 1644 3444 1704
rect 3596 1706 3604 1856
rect 3656 1807 3664 2033
rect 3736 1964 3744 2333
rect 3856 2267 3864 2653
rect 3936 2544 3944 2693
rect 3956 2567 3964 2744
rect 3996 2667 4004 2733
rect 4016 2547 4024 2953
rect 4096 2887 4104 2953
rect 4116 2907 4124 3153
rect 4136 3087 4144 3264
rect 4136 2987 4144 3033
rect 4156 2947 4164 3213
rect 4216 3107 4224 3173
rect 4176 3004 4184 3053
rect 4236 3047 4244 3293
rect 4256 3267 4264 3294
rect 4336 3260 4344 3264
rect 4316 3087 4324 3253
rect 4333 3247 4347 3260
rect 4356 3147 4364 3253
rect 4376 3227 4384 3313
rect 4396 3247 4404 3473
rect 4413 3467 4427 3480
rect 4416 3407 4424 3453
rect 4436 3447 4444 3473
rect 4416 3267 4424 3333
rect 4456 3327 4464 3713
rect 4496 3647 4504 3733
rect 4516 3607 4524 3776
rect 4636 3727 4644 3952
rect 4656 3947 4664 3996
rect 4656 3747 4664 3933
rect 4536 3567 4544 3633
rect 4476 3527 4484 3553
rect 4536 3516 4544 3553
rect 4556 3527 4564 3713
rect 4476 3347 4484 3473
rect 4516 3407 4524 3484
rect 4556 3476 4584 3484
rect 4456 3260 4464 3264
rect 4453 3247 4467 3260
rect 4407 3246 4420 3247
rect 4407 3233 4413 3246
rect 4396 3067 4404 3212
rect 4176 2996 4204 3004
rect 4276 3007 4284 3033
rect 4036 2707 4044 2833
rect 4096 2787 4104 2873
rect 4176 2867 4184 2953
rect 4256 2960 4264 2964
rect 4253 2947 4267 2960
rect 4276 2887 4284 2953
rect 4296 2927 4304 3053
rect 4416 3027 4424 3113
rect 4436 3007 4444 3233
rect 4496 3127 4504 3264
rect 4256 2827 4264 2853
rect 4113 2780 4127 2793
rect 4116 2776 4124 2780
rect 4276 2787 4284 2873
rect 4316 2844 4324 2953
rect 4336 2927 4344 2964
rect 4376 2927 4384 2964
rect 4413 2944 4427 2953
rect 4396 2940 4427 2944
rect 4436 2956 4453 2964
rect 4396 2936 4424 2940
rect 4296 2836 4324 2844
rect 3936 2536 3964 2544
rect 3916 2407 3924 2444
rect 3956 2387 3964 2536
rect 4016 2504 4024 2533
rect 3996 2496 4024 2504
rect 3996 2476 4004 2496
rect 4033 2480 4047 2493
rect 4076 2487 4084 2573
rect 4036 2476 4044 2480
rect 4056 2440 4064 2444
rect 4053 2427 4067 2440
rect 3876 2267 3884 2293
rect 3933 2260 3947 2273
rect 3936 2256 3944 2260
rect 4016 2267 4024 2373
rect 3776 2147 3784 2224
rect 3876 2167 3884 2232
rect 3896 2144 3904 2213
rect 3916 2187 3924 2224
rect 3936 2167 3944 2193
rect 4016 2187 4024 2213
rect 3867 2136 3904 2144
rect 3916 1987 3924 2113
rect 3736 1956 3764 1964
rect 3716 1847 3724 1912
rect 3436 1636 3464 1644
rect 3433 1527 3447 1533
rect 3136 1216 3164 1224
rect 3047 1184 3060 1187
rect 3047 1176 3064 1184
rect 3047 1173 3060 1176
rect 2776 916 2804 924
rect 2836 916 2844 973
rect 2896 967 2904 1033
rect 3136 1007 3144 1173
rect 3156 1047 3164 1216
rect 2556 696 2564 753
rect 2576 547 2584 664
rect 2356 487 2364 533
rect 2213 407 2227 413
rect 2116 396 2124 400
rect 2156 396 2204 404
rect 2196 366 2204 396
rect 2273 400 2287 413
rect 2276 396 2284 400
rect 2376 367 2384 433
rect 2456 396 2464 433
rect 2616 367 2624 433
rect 2186 352 2187 360
rect 2173 347 2187 352
rect 1996 316 2013 327
rect 2000 313 2013 316
rect 2067 313 2073 327
rect 1767 293 1773 307
rect 1596 107 1604 144
rect 1656 107 1664 193
rect 1696 176 1704 213
rect 1736 188 1744 293
rect 1996 227 2004 273
rect 1756 140 1764 144
rect 1716 67 1724 132
rect 1753 127 1767 140
rect 1796 87 1804 213
rect 1936 107 1944 173
rect 1956 146 1964 193
rect 2016 176 2024 253
rect 2096 147 2104 213
rect 2116 146 2124 253
rect 2436 247 2444 364
rect 2173 180 2187 193
rect 2176 176 2184 180
rect 2216 176 2224 213
rect 2256 146 2264 233
rect 2427 216 2453 224
rect 2433 180 2447 193
rect 2436 176 2444 180
rect 2556 187 2564 253
rect 2073 127 2087 132
rect 2136 47 2144 133
rect 2193 127 2207 132
rect 2356 107 2364 174
rect 2500 144 2513 147
rect 2416 67 2424 113
rect 2456 107 2464 144
rect 2496 136 2513 144
rect 2500 133 2513 136
rect 2536 127 2544 174
rect 2596 176 2604 273
rect 2636 207 2644 853
rect 2656 567 2664 793
rect 2696 767 2704 884
rect 2693 724 2707 732
rect 2693 720 2713 724
rect 2696 716 2713 720
rect 2716 696 2724 713
rect 2756 696 2804 704
rect 2736 587 2744 664
rect 2656 367 2664 513
rect 2713 400 2727 413
rect 2756 408 2764 453
rect 2796 427 2804 696
rect 2816 667 2824 884
rect 2896 696 2904 953
rect 2996 916 3004 953
rect 3056 886 3064 973
rect 3116 928 3124 953
rect 2976 827 2984 884
rect 3136 807 3144 833
rect 2973 707 2987 713
rect 2856 447 2864 652
rect 2916 627 2924 664
rect 2956 587 2964 693
rect 2996 666 3004 713
rect 3016 707 3024 733
rect 3053 700 3067 713
rect 3056 696 3064 700
rect 3156 687 3164 1012
rect 3176 886 3184 1393
rect 3196 1227 3204 1333
rect 3216 1247 3224 1393
rect 3286 1392 3287 1400
rect 3273 1387 3287 1392
rect 3316 1367 3324 1434
rect 3413 1447 3427 1453
rect 3436 1407 3444 1513
rect 3236 1216 3244 1253
rect 3276 1216 3324 1224
rect 3196 1027 3204 1153
rect 3253 920 3267 933
rect 3316 928 3324 1216
rect 3336 1207 3344 1273
rect 3416 1247 3424 1393
rect 3436 1216 3444 1372
rect 3456 1287 3464 1636
rect 3496 1547 3504 1693
rect 3556 1647 3564 1704
rect 3616 1704 3624 1773
rect 3667 1764 3680 1767
rect 3667 1753 3684 1764
rect 3676 1736 3684 1753
rect 3616 1696 3664 1704
rect 3716 1696 3744 1704
rect 3516 1436 3524 1493
rect 3476 1367 3484 1434
rect 3616 1407 3624 1553
rect 3636 1487 3644 1696
rect 3656 1436 3664 1593
rect 3736 1507 3744 1696
rect 3493 1387 3507 1393
rect 3476 1227 3484 1353
rect 3536 1307 3544 1404
rect 3576 1367 3584 1404
rect 3676 1367 3684 1404
rect 3356 947 3364 1213
rect 3496 1186 3504 1233
rect 3533 1220 3547 1233
rect 3536 1216 3544 1220
rect 3576 1216 3584 1253
rect 3616 1227 3624 1293
rect 3636 1186 3644 1353
rect 3676 1216 3684 1353
rect 3716 1227 3724 1393
rect 3456 1147 3464 1184
rect 3256 916 3264 920
rect 3296 916 3313 924
rect 3356 916 3364 933
rect 3556 916 3564 993
rect 3596 916 3604 1033
rect 3656 947 3664 1173
rect 3696 1147 3704 1172
rect 3736 1167 3744 1493
rect 3756 1064 3764 1956
rect 3776 1448 3784 1873
rect 3816 1867 3824 1924
rect 3796 1747 3804 1793
rect 3856 1787 3864 1924
rect 3896 1887 3904 1954
rect 3916 1764 3924 1973
rect 3956 1968 3964 2173
rect 3996 1956 4004 2073
rect 4036 1927 4044 2254
rect 3976 1887 3984 1924
rect 4056 1867 4064 2333
rect 4076 2267 4084 2432
rect 4096 2287 4104 2533
rect 4156 2507 4164 2773
rect 4216 2707 4224 2744
rect 4256 2687 4264 2744
rect 4116 2447 4124 2493
rect 4176 2476 4184 2613
rect 4276 2488 4284 2733
rect 4156 2440 4164 2444
rect 4153 2427 4167 2440
rect 4196 2367 4204 2444
rect 4296 2347 4304 2836
rect 4316 2547 4324 2813
rect 4336 2587 4344 2873
rect 4396 2776 4404 2936
rect 4436 2887 4444 2956
rect 4516 2827 4524 3133
rect 4536 2907 4544 3453
rect 4556 3327 4564 3476
rect 4636 3467 4644 3593
rect 4656 3484 4664 3693
rect 4676 3527 4684 3973
rect 4776 3647 4784 4293
rect 4856 4267 4864 4304
rect 4956 4267 4964 4293
rect 4796 4187 4804 4213
rect 4796 3947 4804 4152
rect 4836 4048 4844 4213
rect 4876 4036 4884 4093
rect 4896 4047 4904 4253
rect 4936 4127 4944 4153
rect 4976 4087 4984 4333
rect 4996 4227 5004 4353
rect 5016 4347 5024 4513
rect 5036 4367 5044 4533
rect 5056 4507 5064 4552
rect 5056 4336 5064 4373
rect 5076 4367 5084 4513
rect 5096 4487 5104 4524
rect 5136 4447 5144 4524
rect 5096 4348 5104 4433
rect 5116 4347 5124 4373
rect 5016 4127 5024 4293
rect 5036 4247 5044 4304
rect 5056 4187 5064 4253
rect 5076 4147 5084 4304
rect 4836 3816 4844 3973
rect 4856 3967 4864 4004
rect 4796 3776 4824 3784
rect 4796 3607 4804 3776
rect 4696 3516 4704 3553
rect 4656 3476 4684 3484
rect 4576 3308 4584 3373
rect 4613 3300 4627 3313
rect 4616 3296 4624 3300
rect 4556 3227 4564 3253
rect 4636 3227 4644 3264
rect 4676 3207 4684 3476
rect 4796 3476 4824 3484
rect 4696 3227 4704 3453
rect 4796 3447 4804 3476
rect 4876 3404 4884 3933
rect 4916 3927 4924 3993
rect 4896 3824 4904 3873
rect 4996 3847 5004 3964
rect 5016 3867 5024 3913
rect 5076 3887 5084 4073
rect 5096 4006 5104 4273
rect 5136 4107 5144 4393
rect 5176 4344 5184 4513
rect 5196 4407 5204 4613
rect 5216 4447 5224 4633
rect 5167 4336 5184 4344
rect 5213 4348 5227 4353
rect 5236 4344 5244 4793
rect 5256 4747 5264 4813
rect 5356 4787 5364 4824
rect 5256 4667 5264 4693
rect 5356 4607 5364 4653
rect 5313 4560 5327 4573
rect 5376 4567 5384 4733
rect 5416 4607 5424 4812
rect 5316 4556 5324 4560
rect 5416 4556 5424 4593
rect 5436 4587 5444 4973
rect 5453 4867 5467 4873
rect 5476 4856 5484 5113
rect 5496 5087 5504 5293
rect 5516 5076 5524 5193
rect 5576 5104 5584 5333
rect 5596 5167 5604 5473
rect 5636 5444 5644 5696
rect 5656 5487 5664 5716
rect 5676 5607 5684 5793
rect 5716 5767 5724 5852
rect 5756 5707 5764 5993
rect 5796 5896 5804 5972
rect 5856 5967 5864 6084
rect 5816 5807 5824 5864
rect 5856 5827 5864 5864
rect 5716 5596 5724 5673
rect 5836 5608 5844 5633
rect 5856 5624 5864 5693
rect 5876 5647 5884 5853
rect 5896 5847 5904 6213
rect 5916 6127 5924 6296
rect 5936 6227 5944 6304
rect 5933 6120 5947 6133
rect 5936 6116 5944 6120
rect 5856 5616 5884 5624
rect 5876 5596 5884 5616
rect 5687 5564 5700 5567
rect 5687 5556 5704 5564
rect 5736 5560 5744 5564
rect 5687 5553 5700 5556
rect 5733 5547 5747 5560
rect 5807 5556 5824 5564
rect 5616 5436 5644 5444
rect 5616 5144 5624 5436
rect 5736 5427 5744 5533
rect 5636 5387 5644 5413
rect 5696 5376 5704 5413
rect 5796 5407 5804 5553
rect 5916 5564 5924 6073
rect 5936 5947 5944 5973
rect 5956 5908 5964 6053
rect 5976 6007 5984 6084
rect 5976 5924 5984 5993
rect 5976 5916 6004 5924
rect 5996 5896 6004 5916
rect 6036 5867 6044 5933
rect 5936 5567 5944 5673
rect 5896 5556 5924 5564
rect 5836 5484 5844 5513
rect 5836 5476 5864 5484
rect 5813 5444 5827 5453
rect 5813 5440 5844 5444
rect 5816 5436 5844 5440
rect 5676 5307 5684 5344
rect 5716 5287 5724 5344
rect 5736 5207 5744 5333
rect 5756 5267 5764 5393
rect 5793 5380 5807 5393
rect 5836 5387 5844 5436
rect 5796 5376 5804 5380
rect 5856 5347 5864 5476
rect 5676 5147 5684 5173
rect 5616 5136 5644 5144
rect 5556 5096 5584 5104
rect 5556 5076 5564 5096
rect 5616 5046 5624 5113
rect 5536 4984 5544 5032
rect 5536 4976 5564 4984
rect 5556 4867 5564 4976
rect 5456 4568 5464 4813
rect 5476 4567 5484 4693
rect 5536 4647 5544 4824
rect 5556 4707 5564 4813
rect 5576 4627 5584 4873
rect 5596 4867 5604 4933
rect 5616 4887 5624 5032
rect 5636 4907 5644 5136
rect 5676 5076 5684 5133
rect 5776 5044 5784 5233
rect 5736 5007 5744 5044
rect 5756 5036 5784 5044
rect 5616 4856 5624 4873
rect 5656 4856 5664 4973
rect 5696 4867 5704 4953
rect 5716 4927 5724 4973
rect 5756 4967 5764 5036
rect 5796 4947 5804 5273
rect 5816 4967 5824 5293
rect 5876 5247 5884 5513
rect 5896 5307 5904 5556
rect 5956 5527 5964 5833
rect 5996 5596 6004 5633
rect 6076 5567 6084 6253
rect 5956 5376 5964 5413
rect 5856 5088 5864 5133
rect 5996 5127 6004 5473
rect 6016 5287 6024 5553
rect 6036 5447 6044 5564
rect 6096 5487 6104 5853
rect 6096 5376 6104 5433
rect 6116 5387 6124 5953
rect 6136 5407 6144 5693
rect 6056 5304 6064 5344
rect 6036 5296 6064 5304
rect 6036 5207 6044 5296
rect 6056 5227 6064 5273
rect 5987 5104 6000 5107
rect 5987 5093 6004 5104
rect 5893 5080 5907 5093
rect 5896 5076 5904 5080
rect 5996 5076 6004 5093
rect 5876 5007 5884 5044
rect 5916 5040 5944 5044
rect 5916 5036 5947 5040
rect 5933 5027 5947 5036
rect 5636 4787 5644 4812
rect 5676 4807 5684 4824
rect 5656 4796 5673 4804
rect 5656 4687 5664 4796
rect 5696 4784 5704 4813
rect 5676 4776 5704 4784
rect 5256 4487 5264 4513
rect 5236 4336 5264 4344
rect 5156 4247 5164 4333
rect 5176 4227 5184 4293
rect 5113 4047 5127 4053
rect 5153 4040 5167 4053
rect 5176 4044 5184 4093
rect 5196 4067 5204 4304
rect 5256 4287 5264 4336
rect 5276 4307 5284 4373
rect 5296 4367 5304 4524
rect 5336 4467 5344 4524
rect 5356 4347 5364 4513
rect 5396 4507 5404 4524
rect 5436 4504 5444 4524
rect 5416 4496 5444 4504
rect 5316 4247 5324 4292
rect 5356 4127 5364 4293
rect 5376 4207 5384 4473
rect 5396 4447 5404 4493
rect 5416 4348 5424 4496
rect 5476 4487 5484 4513
rect 5496 4347 5504 4553
rect 5516 4467 5524 4613
rect 5556 4556 5564 4593
rect 5636 4567 5644 4653
rect 5436 4147 5444 4304
rect 5156 4036 5164 4040
rect 5176 4036 5204 4044
rect 5116 3967 5124 3993
rect 5096 3907 5104 3933
rect 4896 3816 4924 3824
rect 4953 3820 4967 3833
rect 4956 3816 4964 3820
rect 4896 3607 4904 3772
rect 4856 3396 4884 3404
rect 4736 3296 4744 3333
rect 4776 3296 4784 3353
rect 4816 3307 4824 3393
rect 4800 3264 4813 3267
rect 4796 3256 4813 3264
rect 4800 3253 4813 3256
rect 4836 3244 4844 3313
rect 4816 3236 4844 3244
rect 4636 2996 4644 3033
rect 4656 3007 4664 3073
rect 4676 2956 4693 2964
rect 4556 2927 4564 2953
rect 4536 2847 4544 2893
rect 4556 2776 4564 2813
rect 4416 2724 4424 2744
rect 4396 2716 4424 2724
rect 4396 2587 4404 2716
rect 4360 2504 4373 2507
rect 4356 2493 4373 2504
rect 4356 2476 4364 2493
rect 4396 2487 4404 2552
rect 4287 2336 4304 2347
rect 4316 2436 4333 2444
rect 4287 2333 4300 2336
rect 4116 2256 4124 2313
rect 4156 2256 4164 2313
rect 4096 2220 4104 2224
rect 4076 2127 4084 2213
rect 4093 2207 4107 2220
rect 4096 1987 4104 2193
rect 4136 2004 4144 2212
rect 4116 1996 4144 2004
rect 4116 1956 4124 1996
rect 4156 1956 4164 2013
rect 4173 1987 4187 1993
rect 3916 1756 3944 1764
rect 3936 1748 3944 1756
rect 3976 1747 3984 1852
rect 3796 1527 3804 1693
rect 3816 1607 3824 1704
rect 3896 1664 3904 1734
rect 3876 1656 3904 1664
rect 3776 1227 3784 1373
rect 3796 1367 3804 1404
rect 3856 1367 3864 1593
rect 3876 1347 3884 1656
rect 3916 1627 3924 1693
rect 3956 1467 3964 1704
rect 3976 1448 3984 1693
rect 3996 1444 4004 1793
rect 4056 1767 4064 1832
rect 4136 1804 4144 1924
rect 4136 1796 4164 1804
rect 4076 1736 4084 1793
rect 4136 1706 4144 1773
rect 4156 1747 4164 1796
rect 4196 1767 4204 2313
rect 4216 2087 4224 2273
rect 4296 2256 4304 2313
rect 4316 2267 4324 2436
rect 4416 2446 4424 2693
rect 4436 2647 4444 2733
rect 4456 2627 4464 2773
rect 4496 2567 4504 2744
rect 4536 2587 4544 2732
rect 4576 2707 4584 2733
rect 4456 2488 4464 2533
rect 4496 2476 4504 2513
rect 4596 2508 4604 2853
rect 4656 2827 4664 2953
rect 4676 2884 4684 2956
rect 4676 2876 4704 2884
rect 4676 2776 4684 2853
rect 4696 2787 4704 2876
rect 4756 2867 4764 3193
rect 4776 2847 4784 3213
rect 4796 3007 4804 3113
rect 4816 2996 4824 3236
rect 4856 3107 4864 3396
rect 4896 3367 4904 3553
rect 4936 3516 4944 3751
rect 5016 3747 5024 3853
rect 5036 3687 5044 3833
rect 5196 3824 5204 4036
rect 5216 3927 5224 4113
rect 5293 4040 5307 4053
rect 5296 4036 5304 4040
rect 5320 4004 5333 4007
rect 5236 3867 5244 3993
rect 5276 3967 5284 4004
rect 5316 3996 5333 4004
rect 5320 3993 5333 3996
rect 5176 3816 5204 3824
rect 5016 3627 5024 3653
rect 5056 3624 5064 3773
rect 5076 3707 5084 3784
rect 5136 3776 5164 3784
rect 5036 3616 5064 3624
rect 5016 3564 5024 3613
rect 4996 3556 5024 3564
rect 4996 3530 5004 3556
rect 5036 3527 5044 3616
rect 5036 3476 5053 3484
rect 5016 3404 5024 3473
rect 4996 3396 5024 3404
rect 4873 3307 4887 3313
rect 4913 3300 4927 3313
rect 4916 3296 4924 3300
rect 4876 3256 4904 3264
rect 4876 3187 4884 3256
rect 4976 3264 4984 3293
rect 4933 3247 4947 3252
rect 4956 3256 4984 3264
rect 4956 3187 4964 3256
rect 4876 3010 4884 3033
rect 4896 3027 4904 3153
rect 4896 2907 4904 2952
rect 4696 2644 4704 2733
rect 4716 2647 4724 2813
rect 4676 2636 4704 2644
rect 4616 2547 4624 2593
rect 4636 2527 4644 2613
rect 4356 2387 4364 2413
rect 4336 2107 4344 2353
rect 4356 2267 4364 2373
rect 4396 2256 4404 2433
rect 4536 2347 4544 2453
rect 4476 2264 4484 2333
rect 4476 2256 4504 2264
rect 4376 2167 4384 2224
rect 4416 2087 4424 2224
rect 4456 2127 4464 2224
rect 4476 2027 4484 2213
rect 4216 1996 4253 2004
rect 4216 1967 4224 1996
rect 4233 1960 4247 1973
rect 4236 1956 4244 1960
rect 4316 1967 4324 1993
rect 4336 1947 4344 1973
rect 4296 1887 4304 1924
rect 4216 1744 4224 1873
rect 4196 1736 4224 1744
rect 4096 1700 4104 1704
rect 4093 1687 4107 1700
rect 3996 1436 4024 1444
rect 3916 1327 3924 1392
rect 3956 1367 3964 1404
rect 4016 1267 4024 1436
rect 4036 1406 4044 1673
rect 4156 1667 4164 1693
rect 4236 1700 4244 1704
rect 4233 1687 4247 1700
rect 4176 1287 4184 1513
rect 4276 1487 4284 1853
rect 4316 1827 4324 1913
rect 4376 1920 4384 1924
rect 4333 1907 4347 1912
rect 4356 1787 4364 1913
rect 4373 1907 4387 1920
rect 4416 1867 4424 1924
rect 4296 1567 4304 1753
rect 4416 1704 4424 1773
rect 4336 1627 4344 1704
rect 4356 1587 4364 1653
rect 4376 1607 4384 1704
rect 4396 1696 4424 1704
rect 4027 1256 4044 1264
rect 3787 1184 3800 1187
rect 3787 1176 3804 1184
rect 3836 1180 3844 1184
rect 3787 1173 3800 1176
rect 3833 1167 3847 1180
rect 3896 1167 3904 1253
rect 3956 1216 3964 1253
rect 4036 1186 4044 1256
rect 4116 1216 4124 1253
rect 3756 1056 3784 1064
rect 3636 936 3653 944
rect 3636 907 3644 936
rect 3676 916 3684 993
rect 3713 920 3727 933
rect 3756 927 3764 1033
rect 3716 916 3724 920
rect 3236 787 3244 884
rect 3273 867 3287 872
rect 3333 867 3347 872
rect 3176 707 3184 773
rect 3416 747 3424 884
rect 3216 696 3224 733
rect 3256 696 3264 733
rect 3356 696 3364 733
rect 2716 396 2724 400
rect 2836 396 2844 433
rect 2873 400 2887 413
rect 2876 396 2884 400
rect 2976 387 2984 593
rect 3076 447 3084 664
rect 3116 567 3124 664
rect 3187 666 3200 667
rect 3187 653 3193 666
rect 3136 607 3144 653
rect 3276 627 3284 664
rect 3336 627 3344 664
rect 3376 607 3384 664
rect 3436 647 3444 693
rect 3456 607 3464 872
rect 3516 696 3524 833
rect 3736 827 3744 884
rect 3556 747 3564 813
rect 3556 696 3564 733
rect 3596 667 3604 813
rect 3616 707 3624 733
rect 3636 696 3644 773
rect 3673 700 3687 713
rect 3676 696 3684 700
rect 3496 607 3504 664
rect 3736 666 3744 713
rect 3756 667 3764 693
rect 3776 687 3784 1056
rect 3796 787 3804 1153
rect 3953 1147 3967 1153
rect 3836 916 3844 973
rect 3956 887 3964 1073
rect 4036 927 4044 953
rect 4056 928 4064 1213
rect 4096 1147 4104 1184
rect 4136 1180 4144 1184
rect 4133 1167 4147 1180
rect 4196 1147 4204 1473
rect 4253 1448 4267 1453
rect 4316 1444 4324 1493
rect 4396 1467 4404 1696
rect 4436 1687 4444 1893
rect 4476 1867 4484 1992
rect 4496 1907 4504 2113
rect 4556 2027 4564 2493
rect 4636 2476 4644 2513
rect 4676 2487 4684 2636
rect 4736 2624 4744 2833
rect 4816 2776 4824 2813
rect 4836 2787 4844 2853
rect 4916 2827 4924 3113
rect 4936 2967 4944 3153
rect 4976 3087 4984 3233
rect 4996 3227 5004 3396
rect 5036 3367 5044 3476
rect 5076 3296 5084 3393
rect 5013 3247 5027 3253
rect 4976 3047 4984 3073
rect 5016 3007 5024 3033
rect 4716 2616 4744 2624
rect 4696 2446 4704 2573
rect 4616 2284 4624 2444
rect 4656 2387 4664 2432
rect 4716 2427 4724 2616
rect 4756 2567 4764 2733
rect 4796 2707 4804 2744
rect 4856 2740 4864 2744
rect 4816 2687 4824 2713
rect 4816 2487 4824 2673
rect 4836 2507 4844 2733
rect 4853 2727 4867 2740
rect 4956 2727 4964 2993
rect 4976 2704 4984 2953
rect 5036 2947 5044 3213
rect 5056 3127 5064 3264
rect 5096 3167 5104 3253
rect 5116 3144 5124 3553
rect 5136 3407 5144 3733
rect 5156 3727 5164 3776
rect 5156 3527 5164 3673
rect 5176 3547 5184 3816
rect 5256 3787 5264 3913
rect 5276 3847 5284 3893
rect 5216 3627 5224 3784
rect 5276 3764 5284 3833
rect 5256 3756 5284 3764
rect 5256 3667 5264 3756
rect 5180 3524 5193 3527
rect 5176 3516 5193 3524
rect 5180 3513 5193 3516
rect 5256 3524 5264 3613
rect 5276 3607 5284 3733
rect 5236 3516 5264 3524
rect 5136 3207 5144 3353
rect 5156 3327 5164 3473
rect 5256 3407 5264 3473
rect 5276 3427 5284 3593
rect 5296 3567 5304 3873
rect 5376 3827 5384 4053
rect 5396 4047 5404 4133
rect 5476 4107 5484 4271
rect 5516 4187 5524 4333
rect 5536 4306 5544 4493
rect 5556 4347 5564 4493
rect 5576 4467 5584 4524
rect 5636 4427 5644 4513
rect 5596 4336 5604 4413
rect 5636 4336 5644 4373
rect 5656 4367 5664 4613
rect 5676 4347 5684 4776
rect 5716 4664 5724 4892
rect 5756 4887 5764 4913
rect 5836 4884 5844 4993
rect 5836 4880 5864 4884
rect 5836 4876 5867 4880
rect 5853 4867 5867 4876
rect 5753 4807 5767 4813
rect 5796 4787 5804 4824
rect 5696 4656 5724 4664
rect 5616 4300 5624 4304
rect 5613 4287 5627 4300
rect 5536 4067 5544 4133
rect 5556 4027 5564 4233
rect 5296 3486 5304 3532
rect 5216 3296 5224 3333
rect 5256 3296 5264 3372
rect 5316 3347 5324 3753
rect 5356 3747 5364 3784
rect 5396 3527 5404 4012
rect 5476 3867 5484 3964
rect 5416 3747 5424 3853
rect 5493 3820 5507 3833
rect 5496 3816 5504 3820
rect 5536 3827 5544 3853
rect 5527 3814 5544 3827
rect 5576 3824 5584 4173
rect 5596 4007 5604 4233
rect 5616 4047 5624 4073
rect 5636 4036 5644 4273
rect 5656 4227 5664 4304
rect 5676 4247 5684 4293
rect 5696 4067 5704 4656
rect 5836 4647 5844 4812
rect 5716 4587 5724 4633
rect 5716 4447 5724 4493
rect 5776 4407 5784 4484
rect 5716 4347 5724 4393
rect 5733 4340 5747 4353
rect 5736 4336 5744 4340
rect 5816 4347 5824 4433
rect 5836 4304 5844 4493
rect 5756 4300 5764 4304
rect 5796 4300 5804 4304
rect 5696 4044 5704 4053
rect 5676 4036 5704 4044
rect 5520 3813 5544 3814
rect 5476 3727 5484 3784
rect 5347 3524 5360 3527
rect 5347 3516 5364 3524
rect 5347 3513 5360 3516
rect 5433 3520 5447 3533
rect 5473 3520 5487 3533
rect 5436 3516 5444 3520
rect 5476 3516 5484 3520
rect 5336 3387 5344 3473
rect 5096 3136 5124 3144
rect 5056 2807 5064 3053
rect 5076 2927 5084 3093
rect 5047 2796 5064 2807
rect 5047 2793 5060 2796
rect 5036 2776 5073 2784
rect 4956 2700 4984 2704
rect 4953 2696 4984 2700
rect 4953 2687 4967 2696
rect 4873 2480 4887 2493
rect 4876 2476 4884 2480
rect 4916 2476 4924 2673
rect 4936 2484 4944 2593
rect 4956 2504 4964 2633
rect 4976 2576 5024 2584
rect 4976 2547 4984 2576
rect 4956 2496 4984 2504
rect 4936 2476 4964 2484
rect 4756 2440 4764 2444
rect 4616 2280 4644 2284
rect 4616 2276 4647 2280
rect 4633 2267 4647 2276
rect 4576 2224 4584 2254
rect 4716 2224 4724 2333
rect 4576 2216 4604 2224
rect 4596 2167 4604 2216
rect 4676 2216 4724 2224
rect 4616 2107 4624 2133
rect 4533 2004 4547 2013
rect 4533 2000 4564 2004
rect 4536 1996 4564 2000
rect 4556 1984 4564 1996
rect 4556 1976 4573 1984
rect 4533 1960 4547 1973
rect 4536 1956 4544 1960
rect 4576 1956 4584 1973
rect 4596 1967 4604 2073
rect 4716 2047 4724 2093
rect 4476 1736 4484 1813
rect 4516 1748 4524 1873
rect 4536 1747 4544 1893
rect 4496 1700 4504 1704
rect 4493 1687 4507 1700
rect 4416 1507 4424 1673
rect 4473 1664 4487 1673
rect 4473 1660 4513 1664
rect 4476 1656 4513 1660
rect 4556 1607 4564 1873
rect 4596 1767 4604 1913
rect 4616 1867 4624 2013
rect 4736 1987 4744 2433
rect 4753 2427 4767 2440
rect 4816 2347 4824 2433
rect 4816 2256 4824 2312
rect 4836 2268 4844 2453
rect 4796 2167 4804 2224
rect 4856 2187 4864 2253
rect 4636 1887 4644 1973
rect 4636 1736 4644 1813
rect 4656 1767 4664 1953
rect 4296 1436 4324 1444
rect 4236 1247 4244 1404
rect 4276 1367 4284 1404
rect 4336 1304 4344 1453
rect 4373 1440 4387 1453
rect 4376 1436 4384 1440
rect 4416 1436 4424 1493
rect 4573 1440 4587 1453
rect 4596 1447 4604 1671
rect 4576 1436 4584 1440
rect 4396 1367 4404 1404
rect 4487 1396 4524 1404
rect 4336 1296 4364 1304
rect 4216 987 4224 1213
rect 4216 947 4224 973
rect 4256 967 4264 1184
rect 4296 1087 4304 1184
rect 4336 1127 4344 1273
rect 4356 1087 4364 1296
rect 4420 1244 4433 1247
rect 4416 1233 4433 1244
rect 4416 1216 4424 1233
rect 4296 1027 4304 1073
rect 4336 967 4344 1053
rect 4256 936 4293 944
rect 4153 920 4167 933
rect 4156 916 4164 920
rect 4056 886 4064 914
rect 4256 916 4264 936
rect 4196 887 4204 913
rect 4336 887 4344 953
rect 4076 880 4093 884
rect 4073 876 4093 880
rect 4073 867 4087 876
rect 3856 696 3864 733
rect 3376 567 3384 593
rect 3016 396 3024 433
rect 3053 400 3067 413
rect 3153 400 3167 413
rect 3056 396 3064 400
rect 3156 396 3164 400
rect 3196 396 3204 453
rect 3216 407 3224 433
rect 2796 347 2804 373
rect 3236 367 3244 394
rect 2676 146 2684 213
rect 2716 176 2724 293
rect 2756 176 2764 333
rect 2576 140 2584 144
rect 2573 127 2587 140
rect 2776 140 2784 144
rect 2773 127 2787 140
rect 2816 67 2824 273
rect 2836 207 2844 313
rect 2896 287 2904 364
rect 3076 360 3084 364
rect 3136 360 3144 364
rect 3073 347 3087 360
rect 3133 347 3147 360
rect 3176 327 3184 364
rect 3213 347 3227 353
rect 3233 327 3247 332
rect 3256 307 3264 413
rect 3276 407 3284 453
rect 3293 400 3307 413
rect 3296 396 3304 400
rect 3376 396 3384 513
rect 3696 487 3704 513
rect 3476 366 3484 473
rect 3533 400 3547 413
rect 3536 396 3544 400
rect 3576 396 3584 453
rect 3636 366 3644 413
rect 3696 396 3704 473
rect 3716 427 3724 653
rect 3833 647 3847 652
rect 3776 467 3784 633
rect 3876 627 3884 664
rect 3916 627 3924 713
rect 3973 700 3987 713
rect 3976 696 3984 700
rect 4016 696 4024 753
rect 3956 660 3964 664
rect 3953 647 3967 660
rect 3816 396 3824 433
rect 3976 396 3984 433
rect 3316 327 3324 364
rect 3436 327 3444 364
rect 2927 193 2933 207
rect 2836 146 2844 193
rect 3036 188 3044 293
rect 3247 276 3273 284
rect 2940 184 2953 187
rect 2936 176 2953 184
rect 2940 173 2953 176
rect 3216 176 3224 253
rect 3256 176 3264 253
rect 3356 176 3364 313
rect 3376 187 3384 213
rect 3416 176 3424 233
rect 2976 146 2984 173
rect 3136 146 3144 173
rect 2996 107 3004 133
rect 3156 107 3164 153
rect 3516 147 3524 293
rect 3556 287 3564 364
rect 3596 347 3604 364
rect 3596 336 3613 347
rect 3600 333 3613 336
rect 3687 333 3693 345
rect 3756 327 3764 394
rect 3196 87 3204 132
rect 3396 47 3404 133
rect 3456 47 3464 144
rect 3536 127 3544 233
rect 3556 187 3564 213
rect 3576 176 3584 293
rect 3656 187 3664 313
rect 3796 267 3804 364
rect 3836 360 3844 364
rect 3956 360 3964 364
rect 3833 347 3847 360
rect 3953 347 3967 360
rect 3936 216 3944 313
rect 4036 227 4044 393
rect 4056 327 4064 813
rect 4076 666 4084 733
rect 4096 607 4104 773
rect 4136 747 4144 884
rect 4236 880 4244 884
rect 4233 867 4247 880
rect 4256 727 4264 753
rect 4256 696 4264 713
rect 4116 527 4124 673
rect 4220 664 4233 667
rect 4156 587 4164 664
rect 4216 656 4233 664
rect 4220 653 4233 656
rect 4156 447 4164 573
rect 4296 408 4304 713
rect 4316 666 4324 773
rect 4356 727 4364 1073
rect 4376 927 4384 973
rect 4407 944 4420 947
rect 4407 933 4424 944
rect 4416 916 4424 933
rect 4436 924 4444 1133
rect 4476 1127 4484 1233
rect 4496 1227 4504 1373
rect 4513 1220 4527 1233
rect 4516 1216 4524 1220
rect 4456 1064 4464 1113
rect 4456 1056 4484 1064
rect 4436 916 4464 924
rect 4456 807 4464 916
rect 4476 747 4484 1056
rect 4496 927 4504 1013
rect 4536 944 4544 1172
rect 4516 936 4544 944
rect 4516 916 4524 936
rect 4556 916 4564 1053
rect 4596 1047 4604 1393
rect 4616 1367 4624 1693
rect 4656 1667 4664 1704
rect 4636 1406 4644 1473
rect 4656 1447 4664 1573
rect 4676 1464 4684 1693
rect 4696 1487 4704 1773
rect 4716 1767 4724 1924
rect 4736 1736 4744 1913
rect 4756 1767 4764 2053
rect 4836 1956 4844 2133
rect 4876 2027 4884 2273
rect 4896 2267 4904 2444
rect 4956 2407 4964 2476
rect 4916 2256 4924 2373
rect 4976 2367 4984 2496
rect 4996 2487 5004 2553
rect 5016 2504 5024 2576
rect 5056 2507 5064 2733
rect 5076 2607 5084 2752
rect 5096 2747 5104 3136
rect 5116 3027 5124 3093
rect 5156 3087 5164 3292
rect 5196 3187 5204 3264
rect 5236 3227 5244 3264
rect 5167 3076 5184 3084
rect 5147 2933 5153 2947
rect 5116 2787 5124 2913
rect 5136 2776 5144 2853
rect 5156 2807 5164 2893
rect 5176 2847 5184 3076
rect 5276 3027 5284 3213
rect 5196 2887 5204 3013
rect 5276 2996 5284 3013
rect 5316 3008 5324 3173
rect 5376 3164 5384 3213
rect 5396 3187 5404 3413
rect 5376 3156 5404 3164
rect 5336 3007 5344 3153
rect 5356 3024 5364 3133
rect 5396 3047 5404 3156
rect 5416 3087 5424 3433
rect 5456 3427 5464 3484
rect 5436 3307 5444 3393
rect 5456 3296 5464 3373
rect 5496 3328 5504 3453
rect 5516 3407 5524 3733
rect 5536 3547 5544 3813
rect 5556 3816 5584 3824
rect 5596 3816 5604 3853
rect 5636 3816 5644 3873
rect 5656 3847 5664 4004
rect 5676 3827 5684 3853
rect 5556 3607 5564 3816
rect 5576 3587 5584 3773
rect 5696 3784 5704 3993
rect 5716 3867 5724 4293
rect 5753 4287 5767 4300
rect 5793 4287 5807 4300
rect 5816 4296 5844 4304
rect 5736 4047 5744 4273
rect 5796 4127 5804 4273
rect 5816 4267 5824 4296
rect 5856 4284 5864 4813
rect 5876 4507 5884 4953
rect 5896 4827 5904 4933
rect 5896 4567 5904 4653
rect 5916 4627 5924 4993
rect 6016 4927 6024 5044
rect 6076 5007 6084 5074
rect 6096 5027 6104 5113
rect 6116 4864 6124 5333
rect 6136 5287 6144 5353
rect 6107 4856 6124 4864
rect 6076 4804 6084 4833
rect 6056 4796 6084 4804
rect 6056 4767 6064 4796
rect 5996 4587 6004 4713
rect 6096 4667 6104 4853
rect 6136 4587 6144 4893
rect 5996 4556 6044 4564
rect 5896 4487 5904 4513
rect 5916 4367 5924 4512
rect 5956 4427 5964 4524
rect 5936 4336 5944 4373
rect 5976 4347 5984 4513
rect 5996 4467 6004 4556
rect 6096 4487 6104 4524
rect 6016 4336 6024 4413
rect 5876 4287 5884 4333
rect 5916 4300 5924 4304
rect 5836 4276 5864 4284
rect 5756 4087 5764 4113
rect 5753 4040 5767 4052
rect 5796 4048 5804 4092
rect 5756 4036 5764 4040
rect 5613 3767 5627 3772
rect 5656 3747 5664 3784
rect 5676 3776 5704 3784
rect 5533 3527 5547 3533
rect 5553 3520 5567 3533
rect 5556 3516 5564 3520
rect 5596 3516 5604 3653
rect 5536 3307 5544 3473
rect 5356 3020 5384 3024
rect 5356 3016 5387 3020
rect 5373 3007 5387 3016
rect 5176 2776 5184 2812
rect 5216 2787 5224 2933
rect 5016 2496 5044 2504
rect 5036 2476 5044 2496
rect 5096 2487 5104 2712
rect 4996 2347 5004 2433
rect 4936 2107 4944 2224
rect 4776 1736 4784 1833
rect 4836 1747 4844 1893
rect 4876 1827 4884 2013
rect 4976 1987 4984 2273
rect 4996 2264 5004 2333
rect 5016 2287 5024 2444
rect 5056 2267 5064 2333
rect 5076 2327 5084 2393
rect 5096 2327 5104 2433
rect 5116 2387 5124 2713
rect 5196 2707 5204 2744
rect 5236 2627 5244 2873
rect 5316 2867 5324 2994
rect 5396 2996 5404 3033
rect 5256 2787 5264 2813
rect 5336 2787 5344 2953
rect 5416 2907 5424 2953
rect 5356 2807 5364 2873
rect 5136 2487 5144 2613
rect 5256 2604 5264 2733
rect 5276 2724 5284 2744
rect 5276 2716 5313 2724
rect 5236 2596 5264 2604
rect 5176 2476 5184 2513
rect 5113 2327 5127 2333
rect 4996 2256 5024 2264
rect 5076 2224 5084 2273
rect 5096 2247 5104 2313
rect 5136 2264 5144 2433
rect 5216 2384 5224 2553
rect 5196 2376 5224 2384
rect 5116 2256 5144 2264
rect 5156 2256 5164 2313
rect 5196 2256 5204 2376
rect 5236 2364 5244 2596
rect 5336 2567 5344 2733
rect 5356 2707 5364 2772
rect 5376 2727 5384 2753
rect 5256 2427 5264 2533
rect 5376 2487 5384 2553
rect 5316 2440 5324 2444
rect 5216 2356 5244 2364
rect 5216 2287 5224 2356
rect 5256 2347 5264 2373
rect 5236 2336 5253 2344
rect 5056 2216 5084 2224
rect 4896 1824 4904 1973
rect 4896 1816 4924 1824
rect 4853 1740 4867 1753
rect 4856 1736 4864 1740
rect 4756 1527 4764 1704
rect 4836 1567 4844 1693
rect 4676 1456 4704 1464
rect 4696 1436 4704 1456
rect 4733 1440 4747 1453
rect 4736 1436 4744 1440
rect 4676 1347 4684 1392
rect 4716 1307 4724 1404
rect 4776 1230 4784 1433
rect 4796 1407 4804 1453
rect 4896 1436 4904 1493
rect 4916 1467 4924 1816
rect 4936 1704 4944 1893
rect 4956 1747 4964 1913
rect 4976 1827 4984 1924
rect 5016 1827 5024 1973
rect 5036 1824 5044 2173
rect 5056 1907 5064 2216
rect 5116 2107 5124 2256
rect 5133 2207 5147 2213
rect 5076 1967 5084 2053
rect 5176 2007 5184 2224
rect 5093 1960 5107 1973
rect 5096 1956 5104 1960
rect 5176 1904 5184 1924
rect 5176 1896 5204 1904
rect 5036 1816 5064 1824
rect 4976 1787 4984 1813
rect 5056 1747 5064 1816
rect 4936 1696 4964 1704
rect 4936 1447 4944 1673
rect 4956 1527 4964 1696
rect 4976 1647 4984 1704
rect 5036 1700 5044 1704
rect 5033 1687 5047 1700
rect 4916 1367 4924 1404
rect 4636 1107 4644 1184
rect 4796 1147 4804 1333
rect 4816 1227 4824 1293
rect 4827 1184 4840 1187
rect 4936 1184 4944 1393
rect 4956 1387 4964 1492
rect 4827 1176 4844 1184
rect 4827 1173 4840 1176
rect 4907 1176 4944 1184
rect 4576 787 4584 872
rect 4616 827 4624 993
rect 4676 967 4684 1113
rect 4696 1087 4704 1113
rect 4716 916 4724 953
rect 4636 887 4644 914
rect 4756 887 4764 1073
rect 4776 847 4784 973
rect 4836 916 4844 993
rect 4816 847 4824 884
rect 4333 704 4347 713
rect 4333 700 4364 704
rect 4336 696 4364 700
rect 4376 527 4384 664
rect 4456 627 4464 693
rect 4516 660 4524 664
rect 4476 587 4484 653
rect 4513 647 4527 660
rect 4576 547 4584 733
rect 4636 696 4644 833
rect 4616 627 4624 664
rect 4656 660 4664 664
rect 4653 647 4667 660
rect 4596 567 4604 593
rect 4096 267 4104 364
rect 3736 176 3744 213
rect 3596 140 3604 144
rect 3593 127 3607 140
rect 3696 107 3704 153
rect 3836 147 3844 213
rect 3756 47 3764 144
rect 4016 67 4024 153
rect 4036 146 4044 213
rect 4133 187 4147 193
rect 4076 87 4084 132
rect 4116 107 4124 144
rect 4156 107 4164 174
rect 4213 107 4227 113
rect 4296 67 4304 394
rect 4316 367 4324 473
rect 4356 396 4364 453
rect 4393 400 4407 413
rect 4396 396 4404 400
rect 4496 364 4504 493
rect 4696 404 4704 713
rect 4736 587 4744 793
rect 4773 700 4787 713
rect 4776 696 4784 700
rect 4816 696 4824 773
rect 4856 707 4864 884
rect 4916 727 4924 1176
rect 4956 1167 4964 1333
rect 4956 1067 4964 1153
rect 4953 987 4967 993
rect 4947 980 4967 987
rect 4947 976 4964 980
rect 4947 973 4960 976
rect 4956 916 4964 953
rect 4976 947 4984 1453
rect 5036 1436 5044 1513
rect 5056 1467 5064 1693
rect 5076 1647 5084 1833
rect 5016 1400 5024 1404
rect 5013 1387 5027 1400
rect 5056 1367 5064 1404
rect 4996 928 5004 1053
rect 5056 967 5064 1213
rect 5076 947 5084 1393
rect 5096 1007 5104 1893
rect 5116 1487 5124 1793
rect 5176 1736 5184 1853
rect 5196 1847 5204 1896
rect 5216 1747 5224 1913
rect 5236 1787 5244 2336
rect 5276 2327 5284 2433
rect 5313 2427 5327 2440
rect 5396 2444 5404 2853
rect 5416 2787 5424 2893
rect 5436 2827 5444 3173
rect 5456 2807 5464 3033
rect 5516 2996 5524 3053
rect 5536 3007 5544 3253
rect 5556 3187 5564 3393
rect 5576 3307 5584 3353
rect 5596 3324 5604 3453
rect 5616 3347 5624 3484
rect 5636 3367 5644 3473
rect 5596 3316 5624 3324
rect 5616 3296 5624 3316
rect 5656 3308 5664 3433
rect 5576 3147 5584 3253
rect 5596 3207 5604 3264
rect 5636 3227 5644 3264
rect 5676 3207 5684 3776
rect 5716 3764 5724 3832
rect 5736 3827 5744 3993
rect 5776 3967 5784 4004
rect 5776 3816 5784 3853
rect 5796 3847 5804 3873
rect 5816 3827 5824 3993
rect 5836 3947 5844 4276
rect 5756 3780 5764 3784
rect 5696 3756 5724 3764
rect 5696 3527 5704 3756
rect 5736 3627 5744 3773
rect 5753 3767 5767 3780
rect 5716 3547 5724 3593
rect 5776 3528 5784 3753
rect 5796 3587 5804 3751
rect 5696 3247 5704 3473
rect 5716 3427 5724 3484
rect 5716 3347 5724 3373
rect 5756 3327 5764 3373
rect 5776 3296 5784 3413
rect 5796 3307 5804 3472
rect 5556 3067 5564 3093
rect 5576 2996 5584 3073
rect 5476 2847 5484 2993
rect 5593 2947 5607 2953
rect 5616 2887 5624 2993
rect 5636 2967 5644 3192
rect 5656 3007 5664 3173
rect 5756 3167 5764 3264
rect 5536 2847 5544 2873
rect 5616 2847 5624 2873
rect 5676 2847 5684 2964
rect 5716 2944 5724 2952
rect 5696 2936 5724 2944
rect 5553 2827 5567 2833
rect 5433 2780 5447 2792
rect 5436 2776 5444 2780
rect 5513 2780 5527 2793
rect 5516 2776 5524 2780
rect 5416 2487 5424 2733
rect 5456 2647 5464 2744
rect 5556 2746 5564 2792
rect 5613 2780 5627 2793
rect 5616 2776 5624 2780
rect 5536 2624 5544 2733
rect 5596 2740 5604 2744
rect 5593 2727 5607 2740
rect 5516 2616 5544 2624
rect 5436 2476 5444 2533
rect 5493 2480 5507 2493
rect 5516 2487 5524 2616
rect 5496 2476 5504 2480
rect 5536 2447 5544 2553
rect 5376 2436 5404 2444
rect 5326 2420 5327 2427
rect 5296 2256 5304 2353
rect 5336 2267 5344 2413
rect 5276 2204 5284 2224
rect 5276 2196 5304 2204
rect 5156 1667 5164 1704
rect 5136 1436 5144 1513
rect 5176 1448 5184 1553
rect 5196 1547 5204 1704
rect 5196 1447 5204 1473
rect 5116 1087 5124 1393
rect 5156 1267 5164 1404
rect 5216 1244 5224 1693
rect 5236 1607 5244 1752
rect 5256 1747 5264 2073
rect 5276 1967 5284 2173
rect 5296 2067 5304 2196
rect 5316 1987 5324 2224
rect 5336 2187 5344 2213
rect 5356 2087 5364 2333
rect 5376 2187 5384 2436
rect 5476 2347 5484 2433
rect 5556 2427 5564 2493
rect 5596 2476 5604 2653
rect 5636 2507 5644 2733
rect 5656 2667 5664 2813
rect 5696 2804 5704 2936
rect 5756 2907 5764 3093
rect 5776 3007 5784 3233
rect 5796 3187 5804 3253
rect 5816 3247 5824 3513
rect 5836 3427 5844 3853
rect 5856 3847 5864 4253
rect 5896 4167 5904 4293
rect 5913 4287 5927 4300
rect 5916 4068 5924 4273
rect 5956 4247 5964 4304
rect 5956 4036 5964 4113
rect 5976 4047 5984 4293
rect 6036 4247 6044 4304
rect 6016 4236 6033 4244
rect 5876 3967 5884 3993
rect 5896 3867 5904 4004
rect 5936 3967 5944 4004
rect 5887 3844 5900 3847
rect 5887 3833 5904 3844
rect 5893 3828 5904 3833
rect 5936 3827 5944 3853
rect 5876 3780 5884 3784
rect 5856 3747 5864 3773
rect 5873 3767 5887 3780
rect 5916 3747 5924 3784
rect 5856 3387 5864 3613
rect 5876 3527 5884 3653
rect 5936 3607 5944 3773
rect 5896 3516 5904 3553
rect 5936 3516 5944 3593
rect 5956 3527 5964 3813
rect 5876 3347 5884 3473
rect 5916 3447 5924 3484
rect 5796 2996 5804 3053
rect 5836 3007 5844 3333
rect 5936 3327 5944 3453
rect 5956 3327 5964 3473
rect 5893 3300 5907 3313
rect 5940 3306 5960 3307
rect 5940 3303 5953 3306
rect 5896 3296 5904 3300
rect 5936 3295 5953 3303
rect 5940 3293 5953 3295
rect 5876 3260 5884 3264
rect 5873 3247 5887 3260
rect 5676 2800 5704 2804
rect 5673 2796 5704 2800
rect 5673 2787 5687 2796
rect 5716 2776 5724 2833
rect 5776 2807 5784 2953
rect 5816 2927 5824 2964
rect 5836 2827 5844 2953
rect 5856 2927 5864 3113
rect 5876 3047 5884 3173
rect 5896 3127 5904 3213
rect 5916 3207 5924 3264
rect 5896 2996 5904 3092
rect 5936 3084 5944 3233
rect 5916 3076 5944 3084
rect 5916 3027 5924 3076
rect 5936 2996 5944 3053
rect 5956 3007 5964 3253
rect 5876 2867 5884 2913
rect 5753 2780 5767 2793
rect 5796 2787 5804 2813
rect 5896 2808 5904 2933
rect 5916 2867 5924 2964
rect 5756 2776 5764 2780
rect 5816 2747 5824 2793
rect 5696 2740 5704 2744
rect 5633 2480 5647 2493
rect 5676 2487 5684 2733
rect 5693 2727 5707 2740
rect 5736 2524 5744 2744
rect 5716 2516 5744 2524
rect 5636 2476 5644 2480
rect 5496 2324 5504 2353
rect 5596 2347 5604 2413
rect 5656 2407 5664 2444
rect 5476 2316 5504 2324
rect 5476 2256 5484 2316
rect 5576 2287 5584 2313
rect 5416 2204 5424 2224
rect 5396 2196 5424 2204
rect 5376 1967 5384 2093
rect 5396 2067 5404 2196
rect 5516 2187 5524 2254
rect 5416 2127 5424 2173
rect 5316 1907 5324 1924
rect 5276 1767 5284 1893
rect 5316 1807 5324 1893
rect 5376 1847 5384 1913
rect 5396 1787 5404 1993
rect 5416 1927 5424 2113
rect 5436 1967 5444 2153
rect 5576 2067 5584 2093
rect 5456 1956 5464 2013
rect 5533 1960 5547 1973
rect 5553 1967 5567 1973
rect 5536 1956 5544 1960
rect 5576 1926 5584 2053
rect 5596 1987 5604 2193
rect 5616 1967 5624 2224
rect 5656 2167 5664 2333
rect 5676 2067 5684 2433
rect 5696 2427 5704 2493
rect 5716 2487 5724 2516
rect 5756 2504 5764 2573
rect 5776 2547 5784 2744
rect 5796 2507 5804 2733
rect 5816 2647 5824 2733
rect 5916 2627 5924 2733
rect 5756 2496 5784 2504
rect 5733 2480 5747 2493
rect 5736 2476 5744 2480
rect 5776 2476 5784 2496
rect 5716 2407 5724 2433
rect 5736 2284 5744 2413
rect 5756 2304 5764 2444
rect 5836 2446 5844 2553
rect 5756 2296 5784 2304
rect 5736 2276 5764 2284
rect 5756 2256 5764 2276
rect 5776 2267 5784 2296
rect 5816 2264 5824 2433
rect 5796 2256 5824 2264
rect 5836 2256 5844 2393
rect 5856 2327 5864 2493
rect 5876 2487 5884 2593
rect 5916 2476 5924 2573
rect 5936 2507 5944 2913
rect 5956 2867 5964 2953
rect 5976 2804 5984 3933
rect 5996 3827 6004 4053
rect 6016 4047 6024 4236
rect 6036 4036 6044 4113
rect 6076 4068 6084 4373
rect 6096 4087 6104 4452
rect 6116 4427 6124 4513
rect 6116 4044 6124 4413
rect 6136 4067 6144 4552
rect 6116 4036 6144 4044
rect 6016 3887 6024 3993
rect 6036 3847 6044 3973
rect 6096 3927 6104 4004
rect 6136 3967 6144 4036
rect 6116 3956 6133 3964
rect 6016 3836 6033 3844
rect 6016 3816 6024 3836
rect 6056 3827 6064 3913
rect 6016 3527 6024 3673
rect 6036 3647 6044 3784
rect 6056 3564 6064 3773
rect 6076 3567 6084 3873
rect 6096 3667 6104 3833
rect 6116 3687 6124 3956
rect 6036 3560 6064 3564
rect 6033 3556 6064 3560
rect 6033 3547 6047 3556
rect 6076 3544 6084 3553
rect 6056 3536 6084 3544
rect 6056 3516 6064 3536
rect 6096 3516 6104 3593
rect 6116 3527 6124 3633
rect 5996 3227 6004 3513
rect 6016 3307 6024 3373
rect 6036 3327 6044 3484
rect 6056 3296 6064 3333
rect 6036 3260 6044 3264
rect 5996 2947 6004 3153
rect 6016 3007 6024 3253
rect 6033 3247 6047 3260
rect 6036 3067 6044 3212
rect 6076 3167 6084 3264
rect 6056 2996 6064 3033
rect 6096 3027 6104 3233
rect 6116 3207 6124 3333
rect 6116 3004 6124 3153
rect 6136 3067 6144 3913
rect 6096 2996 6124 3004
rect 6136 2966 6144 3013
rect 6016 2827 6024 2953
rect 6036 2907 6044 2964
rect 5967 2796 5984 2804
rect 5956 2744 5964 2793
rect 5993 2780 6007 2793
rect 5996 2776 6004 2780
rect 5956 2736 5984 2744
rect 5976 2447 5984 2736
rect 6016 2667 6024 2732
rect 5996 2487 6004 2573
rect 6016 2507 6024 2613
rect 6056 2587 6064 2813
rect 6016 2476 6024 2493
rect 6056 2476 6064 2533
rect 6076 2487 6084 2653
rect 5876 2264 5884 2433
rect 5896 2407 5904 2444
rect 5956 2327 5964 2433
rect 5916 2267 5924 2313
rect 5876 2256 5904 2264
rect 5736 2187 5744 2224
rect 5776 2027 5784 2113
rect 5687 1993 5693 2007
rect 5633 1987 5647 1993
rect 5693 1960 5707 1972
rect 5696 1956 5704 1960
rect 5273 1740 5287 1753
rect 5313 1740 5327 1753
rect 5276 1736 5284 1740
rect 5316 1736 5324 1740
rect 5356 1704 5364 1773
rect 5393 1740 5407 1752
rect 5436 1747 5444 1912
rect 5456 1867 5464 1893
rect 5596 1887 5604 1933
rect 5613 1907 5627 1913
rect 5396 1736 5404 1740
rect 5256 1447 5264 1693
rect 5296 1667 5304 1704
rect 5336 1696 5364 1704
rect 5276 1547 5284 1613
rect 5276 1436 5284 1533
rect 5316 1447 5324 1533
rect 5196 1236 5224 1244
rect 5036 886 5044 913
rect 5036 847 5044 872
rect 4973 700 4987 713
rect 4976 696 4984 700
rect 4796 624 4804 664
rect 4813 624 4827 633
rect 4796 620 4827 624
rect 4796 616 4824 620
rect 4676 396 4704 404
rect 4713 400 4727 413
rect 4716 396 4724 400
rect 4376 327 4384 364
rect 4416 360 4424 364
rect 4413 347 4427 360
rect 4496 356 4524 364
rect 4356 176 4364 253
rect 4316 127 4324 173
rect 4413 127 4427 133
rect 4436 107 4444 174
rect 4467 184 4480 187
rect 4467 176 4484 184
rect 4516 176 4524 356
rect 4556 188 4564 352
rect 4676 327 4684 396
rect 4816 347 4824 616
rect 4856 410 4864 653
rect 4876 647 4884 694
rect 4896 656 4924 664
rect 4896 396 4904 656
rect 4467 173 4480 176
rect 4836 144 4844 213
rect 4856 144 4864 396
rect 4916 267 4924 364
rect 4956 227 4964 664
rect 4976 487 4984 613
rect 4996 587 5004 664
rect 5016 396 5024 553
rect 5036 427 5044 693
rect 5056 647 5064 932
rect 5096 927 5104 953
rect 5136 947 5144 1173
rect 5156 1087 5164 1184
rect 5126 933 5127 940
rect 5113 920 5127 933
rect 5116 916 5124 920
rect 5156 916 5164 973
rect 5196 967 5204 1236
rect 5236 1224 5244 1433
rect 5256 1244 5264 1393
rect 5296 1367 5304 1404
rect 5256 1236 5284 1244
rect 5216 1216 5244 1224
rect 5276 1216 5284 1236
rect 5216 1167 5224 1216
rect 5336 1227 5344 1696
rect 5356 1447 5364 1673
rect 5376 1524 5384 1693
rect 5376 1516 5404 1524
rect 5376 1436 5384 1493
rect 5396 1467 5404 1516
rect 5416 1507 5424 1704
rect 5436 1547 5444 1693
rect 5456 1487 5464 1853
rect 5476 1704 5484 1873
rect 5616 1787 5624 1872
rect 5636 1847 5644 1924
rect 5713 1887 5727 1893
rect 5736 1867 5744 1954
rect 5756 1927 5764 1973
rect 5776 1964 5784 1992
rect 5796 1987 5804 2256
rect 5816 1984 5824 2213
rect 5856 2107 5864 2224
rect 5816 1976 5844 1984
rect 5776 1956 5804 1964
rect 5836 1956 5844 1976
rect 5853 1967 5867 1973
rect 5787 1893 5793 1907
rect 5636 1807 5644 1833
rect 5496 1747 5504 1773
rect 5593 1720 5607 1734
rect 5596 1716 5604 1720
rect 5476 1696 5504 1704
rect 5476 1627 5484 1673
rect 5496 1467 5504 1696
rect 5536 1647 5544 1704
rect 5576 1426 5584 1673
rect 5674 1607 5682 1673
rect 5696 1647 5704 1833
rect 5816 1827 5824 1924
rect 5876 1907 5884 1953
rect 5856 1827 5864 1873
rect 5896 1827 5904 2256
rect 5976 2256 5984 2353
rect 5996 2287 6004 2433
rect 6016 2364 6024 2393
rect 6036 2387 6044 2444
rect 6016 2356 6044 2364
rect 6016 2267 6024 2313
rect 5916 1967 5924 2213
rect 5936 2067 5944 2224
rect 5956 1956 5964 2013
rect 5996 1956 6004 2224
rect 6016 1964 6024 2213
rect 6036 2027 6044 2356
rect 6056 2327 6064 2393
rect 6016 1956 6044 1964
rect 5916 1847 5924 1913
rect 5976 1887 5984 1924
rect 5967 1836 6004 1844
rect 5716 1687 5724 1753
rect 5976 1747 5984 1813
rect 5996 1727 6004 1836
rect 5967 1724 5980 1727
rect 5967 1716 5984 1724
rect 5967 1713 5980 1716
rect 6036 1724 6044 1956
rect 6056 1744 6064 2273
rect 6076 1926 6084 2433
rect 6096 2407 6104 2933
rect 6056 1736 6084 1744
rect 6036 1716 6064 1724
rect 5716 1527 5724 1573
rect 5896 1517 5913 1524
rect 5896 1516 5924 1517
rect 5896 1456 5904 1516
rect 5256 1180 5264 1184
rect 5296 1180 5304 1184
rect 5253 1167 5267 1180
rect 5293 1167 5307 1180
rect 5076 747 5084 912
rect 5096 807 5104 873
rect 5136 844 5144 884
rect 5216 886 5224 1033
rect 5276 944 5284 1133
rect 5356 1127 5364 1393
rect 5436 1264 5444 1404
rect 5476 1367 5484 1412
rect 5436 1256 5464 1264
rect 5416 1216 5424 1253
rect 5456 1227 5464 1256
rect 5376 1187 5384 1213
rect 5476 1187 5484 1273
rect 5296 967 5304 1113
rect 5436 1007 5444 1172
rect 5456 1047 5464 1173
rect 5496 1047 5504 1393
rect 5536 1307 5544 1373
rect 5556 1287 5564 1353
rect 5576 1327 5584 1412
rect 5596 1387 5604 1453
rect 5513 1228 5527 1233
rect 5676 1208 5684 1313
rect 5696 1227 5704 1293
rect 5716 1224 5724 1313
rect 5856 1307 5864 1412
rect 5936 1367 5944 1473
rect 5956 1347 5964 1513
rect 5976 1327 5984 1653
rect 6016 1448 6024 1684
rect 6036 1467 6044 1673
rect 6056 1487 6064 1716
rect 6076 1527 6084 1736
rect 5996 1227 6004 1353
rect 5716 1216 5744 1224
rect 5516 1180 5533 1184
rect 5513 1176 5533 1180
rect 5513 1167 5527 1176
rect 5716 1164 5724 1194
rect 5736 1167 5744 1216
rect 6016 1207 6024 1333
rect 6056 1227 6064 1393
rect 6076 1207 6084 1453
rect 6096 1304 6104 2353
rect 6116 2344 6124 2913
rect 6136 2607 6144 2853
rect 6136 2367 6144 2533
rect 6116 2336 6144 2344
rect 6116 1407 6124 2313
rect 6096 1296 6124 1304
rect 5987 1204 6000 1207
rect 5987 1196 6004 1204
rect 5987 1193 6000 1196
rect 6096 1184 6104 1273
rect 6076 1176 6104 1184
rect 5696 1156 5724 1164
rect 5276 936 5304 944
rect 5296 928 5304 936
rect 5247 924 5260 927
rect 5247 916 5264 924
rect 5247 913 5260 916
rect 5336 927 5344 953
rect 5356 887 5364 933
rect 5396 916 5404 993
rect 5440 924 5453 927
rect 5436 916 5453 924
rect 5440 913 5453 916
rect 5196 844 5204 873
rect 5136 836 5204 844
rect 5093 700 5107 713
rect 5096 696 5104 700
rect 5136 696 5144 733
rect 5236 696 5244 793
rect 5276 787 5284 872
rect 5276 747 5284 773
rect 5316 708 5324 884
rect 5453 867 5467 873
rect 5476 708 5484 893
rect 5056 396 5064 433
rect 5116 404 5124 652
rect 5156 507 5164 664
rect 5216 627 5224 664
rect 5376 660 5384 664
rect 5256 607 5264 652
rect 5373 647 5387 660
rect 5416 507 5424 664
rect 5456 587 5464 664
rect 5496 567 5504 993
rect 5516 807 5524 1113
rect 5553 920 5567 933
rect 5556 916 5564 920
rect 5596 916 5604 1093
rect 5696 984 5704 1156
rect 6076 1164 6084 1176
rect 6036 1156 6084 1164
rect 5716 1007 5724 1133
rect 6012 1107 6020 1133
rect 5856 1007 5864 1073
rect 5696 980 5724 984
rect 5696 976 5727 980
rect 5696 948 5704 976
rect 5713 967 5727 976
rect 5576 747 5584 884
rect 5616 880 5624 884
rect 5613 867 5627 880
rect 5596 756 5633 764
rect 5556 696 5564 733
rect 5596 696 5604 756
rect 5656 744 5664 933
rect 5736 880 5744 884
rect 5733 867 5747 880
rect 5636 736 5664 744
rect 5616 707 5624 733
rect 5576 607 5584 664
rect 5636 504 5644 736
rect 5656 607 5664 713
rect 5716 696 5724 753
rect 5753 700 5767 713
rect 5756 696 5764 700
rect 5616 496 5644 504
rect 5676 504 5684 653
rect 5696 547 5704 664
rect 5676 496 5704 504
rect 5116 396 5144 404
rect 5076 360 5084 364
rect 5073 347 5087 360
rect 5136 347 5144 396
rect 5156 267 5164 433
rect 5376 396 5384 493
rect 5433 400 5447 413
rect 5493 400 5507 413
rect 5436 396 5444 400
rect 5496 396 5504 400
rect 5556 396 5564 453
rect 5596 387 5604 473
rect 5616 427 5624 496
rect 5696 407 5704 496
rect 5016 188 5024 253
rect 5196 184 5204 253
rect 5216 227 5224 364
rect 5196 176 5224 184
rect 5376 188 5384 213
rect 5596 188 5604 373
rect 5687 356 5704 364
rect 5216 144 5224 176
rect 5696 184 5704 356
rect 5716 307 5724 553
rect 5736 467 5744 664
rect 5776 660 5784 664
rect 5773 647 5787 660
rect 5773 524 5787 533
rect 5756 520 5787 524
rect 5756 516 5784 520
rect 5756 396 5764 516
rect 5776 424 5784 493
rect 5796 487 5804 653
rect 5816 427 5824 993
rect 5856 916 5864 953
rect 5847 704 5860 707
rect 5847 696 5864 704
rect 5847 693 5860 696
rect 5876 587 5884 664
rect 5916 427 5924 793
rect 5936 547 5944 1073
rect 5996 928 6004 993
rect 5996 660 6004 664
rect 5993 647 6007 660
rect 5776 416 5804 424
rect 5796 396 5804 416
rect 5816 307 5824 364
rect 5696 176 5724 184
rect 5776 176 5784 293
rect 5856 146 5864 413
rect 5876 366 5884 413
rect 5936 396 5944 433
rect 5956 344 5964 364
rect 5956 336 5984 344
rect 5956 176 5964 313
rect 5976 287 5984 336
rect 6016 327 6024 493
rect 6036 366 6044 1033
rect 6056 287 6064 1113
rect 6076 447 6084 1133
rect 4536 67 4544 144
rect 2787 33 2793 47
rect 2847 33 2853 47
rect 4676 -16 4684 144
rect 5056 -16 5064 144
rect 5416 -16 5424 144
rect 5556 -16 5564 144
rect 4656 -24 4684 -16
rect 5036 -24 5064 -16
rect 5396 -24 5424 -16
rect 5536 -24 5564 -16
rect 5676 -24 5684 144
rect 5816 -16 5824 144
rect 5976 140 5984 144
rect 5973 127 5987 140
rect 6076 127 6084 433
rect 6096 408 6104 1153
rect 6116 507 6124 1296
rect 6136 1127 6144 2336
rect 6136 307 6144 1073
rect 5796 -24 5824 -16
<< m3contact >>
rect 3333 6253 3347 6267
rect 3873 6253 3887 6267
rect 4853 6253 4867 6267
rect 3533 6233 3547 6247
rect 3853 6233 3867 6247
rect 293 6213 307 6227
rect 653 6213 667 6227
rect 913 6213 927 6227
rect 93 6153 107 6167
rect 253 6153 267 6167
rect 173 6114 187 6128
rect 213 6114 227 6128
rect 513 6173 527 6187
rect 393 6153 407 6167
rect 292 6113 306 6127
rect 313 6114 327 6128
rect 353 6114 367 6128
rect 593 6133 607 6147
rect 513 6114 527 6128
rect 753 6193 767 6207
rect 733 6173 747 6187
rect 693 6114 707 6128
rect 873 6153 887 6167
rect 753 6133 767 6147
rect 793 6133 807 6147
rect 853 6133 867 6147
rect 113 5913 127 5927
rect 153 5894 167 5908
rect 233 6072 247 6086
rect 273 6072 287 6086
rect 313 6073 327 6087
rect 413 6072 427 6086
rect 473 6072 487 6086
rect 373 5953 387 5967
rect 393 5914 407 5928
rect 213 5893 227 5907
rect 273 5894 287 5908
rect 333 5894 347 5908
rect 393 5894 407 5908
rect 433 5894 447 5908
rect 93 5813 107 5827
rect 93 5613 107 5627
rect 73 5594 87 5608
rect 33 5513 47 5527
rect 13 5374 27 5388
rect 13 5233 27 5247
rect 193 5813 207 5827
rect 173 5773 187 5787
rect 153 5713 167 5727
rect 133 5513 147 5527
rect 93 5473 107 5487
rect 133 5473 147 5487
rect 293 5852 307 5866
rect 253 5773 267 5787
rect 333 5833 347 5847
rect 413 5852 427 5866
rect 393 5833 407 5847
rect 373 5813 387 5827
rect 293 5693 307 5707
rect 213 5653 227 5667
rect 273 5653 287 5667
rect 173 5593 187 5607
rect 233 5594 247 5608
rect 213 5552 227 5566
rect 53 5433 67 5447
rect 193 5453 207 5467
rect 133 5374 147 5388
rect 253 5433 267 5447
rect 213 5393 227 5407
rect 293 5594 307 5608
rect 333 5594 347 5608
rect 593 6073 607 6087
rect 633 6072 647 6086
rect 673 6072 687 6086
rect 773 6072 787 6086
rect 813 6072 827 6086
rect 1433 6193 1447 6207
rect 1993 6193 2007 6207
rect 2073 6193 2087 6207
rect 2233 6193 2247 6207
rect 3193 6193 3207 6207
rect 3253 6193 3267 6207
rect 3533 6193 3547 6207
rect 1093 6153 1107 6167
rect 1193 6153 1207 6167
rect 1373 6153 1387 6167
rect 953 6114 967 6128
rect 1013 6114 1027 6128
rect 1133 6114 1147 6128
rect 873 6093 887 6107
rect 933 6072 947 6086
rect 853 6053 867 6067
rect 533 6033 547 6047
rect 633 6033 647 6047
rect 773 6033 787 6047
rect 593 5993 607 6007
rect 553 5913 567 5927
rect 493 5893 507 5907
rect 793 6013 807 6027
rect 973 6013 987 6027
rect 853 5993 867 6007
rect 653 5973 667 5987
rect 793 5973 807 5987
rect 1013 5973 1027 5987
rect 633 5953 647 5967
rect 473 5813 487 5827
rect 473 5713 487 5727
rect 393 5593 407 5607
rect 433 5594 447 5608
rect 533 5852 547 5866
rect 573 5852 587 5866
rect 613 5852 627 5866
rect 553 5813 567 5827
rect 613 5813 627 5827
rect 533 5594 547 5608
rect 293 5553 307 5567
rect 353 5552 367 5566
rect 393 5553 407 5567
rect 613 5713 627 5727
rect 573 5633 587 5647
rect 473 5533 487 5547
rect 533 5533 547 5547
rect 353 5473 367 5487
rect 393 5473 407 5487
rect 453 5473 467 5487
rect 293 5453 307 5467
rect 293 5413 307 5427
rect 273 5393 287 5407
rect 213 5332 227 5346
rect 273 5332 287 5346
rect 153 5313 167 5327
rect 193 5313 207 5327
rect 93 5273 107 5287
rect 312 5273 326 5287
rect 333 5273 347 5287
rect 193 5213 207 5227
rect 93 5133 107 5147
rect 53 5074 67 5088
rect 133 5074 147 5088
rect 33 5032 47 5046
rect 153 5032 167 5046
rect 113 5013 127 5027
rect 173 4873 187 4887
rect 413 5413 427 5427
rect 553 5413 567 5427
rect 513 5374 527 5388
rect 1113 6072 1127 6086
rect 1233 6114 1247 6128
rect 1333 6114 1347 6128
rect 1653 6153 1667 6167
rect 1773 6153 1787 6167
rect 1873 6153 1887 6167
rect 1473 6114 1487 6128
rect 1513 6114 1527 6128
rect 1573 6114 1587 6128
rect 1733 6114 1747 6128
rect 1813 6114 1827 6128
rect 1253 6053 1267 6067
rect 1333 6053 1347 6067
rect 1193 5973 1207 5987
rect 993 5933 1007 5947
rect 1073 5933 1087 5947
rect 733 5894 747 5908
rect 813 5893 827 5907
rect 893 5894 907 5908
rect 933 5894 947 5908
rect 713 5833 727 5847
rect 713 5793 727 5807
rect 773 5793 787 5807
rect 633 5633 647 5647
rect 673 5594 687 5608
rect 813 5693 827 5707
rect 853 5653 867 5667
rect 793 5633 807 5647
rect 813 5594 827 5608
rect 853 5573 867 5587
rect 613 5552 627 5566
rect 713 5553 727 5567
rect 753 5552 767 5566
rect 793 5552 807 5566
rect 913 5833 927 5847
rect 913 5594 927 5608
rect 873 5513 887 5527
rect 933 5513 947 5527
rect 653 5473 667 5487
rect 1233 5913 1247 5927
rect 1053 5894 1067 5908
rect 1133 5894 1147 5908
rect 1033 5833 1047 5847
rect 1093 5673 1107 5687
rect 1033 5633 1047 5647
rect 1293 5894 1307 5908
rect 1433 6072 1447 6086
rect 1493 6072 1507 6086
rect 1493 6033 1507 6047
rect 1393 6013 1407 6027
rect 1353 5993 1367 6007
rect 1413 5973 1427 5987
rect 1393 5933 1407 5947
rect 1393 5894 1407 5908
rect 1213 5852 1227 5866
rect 1313 5852 1327 5866
rect 1373 5833 1387 5847
rect 1253 5813 1267 5827
rect 1353 5813 1367 5827
rect 1153 5673 1167 5687
rect 1133 5613 1147 5627
rect 1273 5773 1287 5787
rect 1253 5653 1267 5667
rect 1233 5613 1247 5627
rect 1153 5594 1167 5608
rect 1193 5594 1207 5608
rect 1073 5552 1087 5566
rect 1133 5553 1147 5567
rect 993 5433 1007 5447
rect 753 5413 767 5427
rect 833 5413 847 5427
rect 913 5413 927 5427
rect 573 5393 587 5407
rect 613 5393 627 5407
rect 673 5393 687 5407
rect 713 5374 727 5388
rect 773 5373 787 5387
rect 873 5374 887 5388
rect 413 5313 427 5327
rect 393 5293 407 5307
rect 353 5213 367 5227
rect 333 5133 347 5147
rect 253 5074 267 5088
rect 293 5074 307 5088
rect 233 5032 247 5046
rect 273 4973 287 4987
rect 233 4873 247 4887
rect 113 4854 127 4868
rect 153 4813 167 4827
rect 133 4793 147 4807
rect 93 4733 107 4747
rect 13 4653 27 4667
rect 73 4593 87 4607
rect 273 4854 287 4868
rect 313 4853 327 4867
rect 173 4793 187 4807
rect 33 4554 47 4568
rect 73 4554 87 4568
rect 113 4554 127 4568
rect 152 4554 166 4568
rect 313 4812 327 4826
rect 353 5093 367 5107
rect 433 5253 447 5267
rect 453 5133 467 5147
rect 353 5013 367 5027
rect 573 5332 587 5346
rect 613 5332 627 5346
rect 653 5332 667 5346
rect 753 5332 767 5346
rect 693 5293 707 5307
rect 533 5273 547 5287
rect 553 5233 567 5247
rect 513 5193 527 5207
rect 693 5193 707 5207
rect 813 5313 827 5327
rect 853 5293 867 5307
rect 773 5153 787 5167
rect 553 5133 567 5147
rect 513 5074 527 5088
rect 673 5093 687 5107
rect 713 5074 727 5088
rect 753 5074 767 5088
rect 493 4993 507 5007
rect 433 4973 447 4987
rect 633 4993 647 5007
rect 413 4953 427 4967
rect 513 4953 527 4967
rect 573 4953 587 4967
rect 393 4893 407 4907
rect 373 4854 387 4868
rect 493 4893 507 4907
rect 473 4854 487 4868
rect 393 4812 407 4826
rect 433 4812 447 4826
rect 253 4773 267 4787
rect 193 4733 207 4747
rect 213 4733 227 4747
rect 93 4453 107 4467
rect 53 4334 67 4348
rect 93 4334 107 4348
rect 173 4553 187 4567
rect 233 4593 247 4607
rect 293 4553 307 4567
rect 213 4512 227 4526
rect 173 4473 187 4487
rect 13 3933 27 3947
rect 13 3613 27 3627
rect 153 4333 167 4347
rect 233 4373 247 4387
rect 333 4773 347 4787
rect 333 4713 347 4727
rect 313 4513 327 4527
rect 293 4473 307 4487
rect 253 4353 267 4367
rect 293 4353 307 4367
rect 273 4334 287 4348
rect 312 4334 326 4348
rect 473 4673 487 4687
rect 553 4873 567 4887
rect 593 4854 607 4868
rect 553 4793 567 4807
rect 533 4733 547 4747
rect 493 4613 507 4627
rect 393 4553 407 4567
rect 433 4554 447 4568
rect 373 4512 387 4526
rect 413 4453 427 4467
rect 373 4373 387 4387
rect 113 4292 127 4306
rect 173 4293 187 4307
rect 213 4292 227 4306
rect 113 4073 127 4087
rect 333 4333 347 4347
rect 453 4353 467 4367
rect 353 4292 367 4306
rect 433 4293 447 4307
rect 393 4273 407 4287
rect 573 4713 587 4727
rect 613 4673 627 4687
rect 513 4554 527 4568
rect 553 4554 567 4568
rect 533 4512 547 4526
rect 693 5013 707 5027
rect 1253 5593 1267 5607
rect 1213 5552 1227 5566
rect 933 5374 947 5388
rect 973 5374 987 5388
rect 1013 5374 1027 5388
rect 1073 5372 1087 5386
rect 993 5332 1007 5346
rect 973 5293 987 5307
rect 1033 5293 1047 5307
rect 1073 5293 1087 5307
rect 933 5233 947 5247
rect 1113 5433 1127 5447
rect 1173 5413 1187 5427
rect 1313 5594 1327 5608
rect 1413 5853 1427 5867
rect 1473 5852 1487 5866
rect 1573 5993 1587 6007
rect 1673 6072 1687 6086
rect 1713 6072 1727 6086
rect 1633 5933 1647 5947
rect 1553 5894 1567 5908
rect 1613 5894 1627 5908
rect 1673 5894 1687 5908
rect 1793 6072 1807 6086
rect 1833 6033 1847 6047
rect 1733 6013 1747 6027
rect 1913 6114 1927 6128
rect 1953 6114 1967 6128
rect 2033 6173 2047 6187
rect 1913 6072 1927 6086
rect 1773 5953 1787 5967
rect 1873 5953 1887 5967
rect 1593 5852 1607 5866
rect 1693 5852 1707 5866
rect 1553 5813 1567 5827
rect 1533 5773 1547 5787
rect 1733 5733 1747 5747
rect 1473 5594 1487 5608
rect 1613 5613 1627 5627
rect 1573 5594 1587 5608
rect 1653 5593 1667 5607
rect 1753 5713 1767 5727
rect 1893 5933 1907 5947
rect 1813 5894 1827 5908
rect 1873 5894 1887 5908
rect 1793 5853 1807 5867
rect 1833 5852 1847 5866
rect 1873 5813 1887 5827
rect 1793 5733 1807 5747
rect 2113 6114 2127 6128
rect 2173 6114 2187 6128
rect 2253 6173 2267 6187
rect 2373 6173 2387 6187
rect 2473 6173 2487 6187
rect 3093 6173 3107 6187
rect 2273 6113 2287 6127
rect 2453 6114 2467 6128
rect 2093 6072 2107 6086
rect 1973 6053 1987 6067
rect 2033 6053 2047 6067
rect 1953 6013 1967 6027
rect 2053 5993 2067 6007
rect 1993 5894 2007 5908
rect 1973 5852 1987 5866
rect 2013 5852 2027 5866
rect 2173 6073 2187 6087
rect 2253 6072 2267 6086
rect 2353 6072 2367 6086
rect 2133 5953 2147 5967
rect 2113 5933 2127 5947
rect 2253 5894 2267 5908
rect 2353 5894 2367 5908
rect 2433 5953 2447 5967
rect 2113 5852 2127 5866
rect 2053 5833 2067 5847
rect 1913 5773 1927 5787
rect 2373 5852 2387 5866
rect 2273 5813 2287 5827
rect 2233 5733 2247 5747
rect 1913 5713 1927 5727
rect 2413 5713 2427 5727
rect 1773 5673 1787 5687
rect 1793 5613 1807 5627
rect 1333 5513 1347 5527
rect 1393 5513 1407 5527
rect 1533 5553 1547 5567
rect 1593 5552 1607 5566
rect 1653 5552 1667 5566
rect 1713 5552 1727 5566
rect 1493 5513 1507 5527
rect 1693 5513 1707 5527
rect 1453 5493 1467 5507
rect 1633 5493 1647 5507
rect 1713 5493 1727 5507
rect 1693 5473 1707 5487
rect 1353 5453 1367 5467
rect 1452 5453 1466 5467
rect 1473 5453 1487 5467
rect 1273 5374 1287 5388
rect 1313 5374 1327 5388
rect 1193 5332 1207 5346
rect 1293 5293 1307 5307
rect 1153 5273 1167 5287
rect 1253 5273 1267 5287
rect 1133 5233 1147 5247
rect 1233 5233 1247 5247
rect 1093 5193 1107 5207
rect 1173 5193 1187 5207
rect 973 5153 987 5167
rect 1093 5153 1107 5167
rect 813 5074 827 5088
rect 873 5073 887 5087
rect 1153 5113 1167 5127
rect 833 5032 847 5046
rect 773 5013 787 5027
rect 873 5013 887 5027
rect 753 4953 767 4967
rect 792 4953 806 4967
rect 813 4953 827 4967
rect 693 4873 707 4887
rect 733 4854 747 4868
rect 653 4813 667 4827
rect 713 4773 727 4787
rect 733 4733 747 4747
rect 753 4713 767 4727
rect 773 4693 787 4707
rect 773 4653 787 4667
rect 733 4573 747 4587
rect 673 4554 687 4568
rect 713 4554 727 4568
rect 773 4553 787 4567
rect 593 4493 607 4507
rect 633 4493 647 4507
rect 533 4453 547 4467
rect 573 4453 587 4467
rect 533 4334 547 4348
rect 473 4293 487 4307
rect 453 4253 467 4267
rect 313 4073 327 4087
rect 393 4073 407 4087
rect 253 4053 267 4067
rect 153 4034 167 4048
rect 193 4034 207 4048
rect 233 4034 247 4048
rect 53 3993 67 4007
rect 93 3992 107 4006
rect 133 3973 147 3987
rect 113 3913 127 3927
rect 53 3833 67 3847
rect 153 3893 167 3907
rect 333 4033 347 4047
rect 213 3993 227 4007
rect 193 3813 207 3827
rect 53 3772 67 3786
rect 93 3772 107 3786
rect 173 3733 187 3747
rect 193 3593 207 3607
rect 133 3512 147 3526
rect 253 3973 267 3987
rect 273 3893 287 3907
rect 253 3833 267 3847
rect 333 3913 347 3927
rect 553 4273 567 4287
rect 513 4253 527 4267
rect 693 4512 707 4526
rect 613 4393 627 4407
rect 653 4393 667 4407
rect 913 4973 927 4987
rect 993 5013 1007 5027
rect 953 4953 967 4967
rect 853 4854 867 4868
rect 1093 5074 1107 5088
rect 1073 4973 1087 4987
rect 1013 4933 1027 4947
rect 1013 4873 1027 4887
rect 813 4813 827 4827
rect 873 4812 887 4826
rect 973 4812 987 4826
rect 1013 4812 1027 4826
rect 873 4773 887 4787
rect 1053 4713 1067 4727
rect 873 4633 887 4647
rect 973 4613 987 4627
rect 813 4553 827 4567
rect 793 4513 807 4527
rect 733 4353 747 4367
rect 673 4334 687 4348
rect 613 4273 627 4287
rect 593 4233 607 4247
rect 693 4293 707 4307
rect 653 4193 667 4207
rect 893 4493 907 4507
rect 813 4473 827 4487
rect 853 4473 867 4487
rect 773 4453 787 4467
rect 1033 4593 1047 4607
rect 1093 4854 1107 4868
rect 1393 5373 1407 5387
rect 1553 5373 1567 5387
rect 1633 5374 1647 5388
rect 1833 5594 1847 5608
rect 1873 5594 1887 5608
rect 1933 5693 1947 5707
rect 1993 5673 2007 5687
rect 1953 5613 1967 5627
rect 1933 5594 1947 5608
rect 1853 5552 1867 5566
rect 1913 5553 1927 5567
rect 2773 6153 2787 6167
rect 2853 6153 2867 6167
rect 2573 6114 2587 6128
rect 2733 6114 2747 6128
rect 2773 6114 2787 6128
rect 2813 6114 2827 6128
rect 2953 6114 2967 6128
rect 2453 5893 2467 5907
rect 2513 6072 2527 6086
rect 2713 6072 2727 6086
rect 3033 6113 3047 6127
rect 2713 6033 2727 6047
rect 2753 6033 2767 6047
rect 2553 5933 2567 5947
rect 2633 5933 2647 5947
rect 2533 5894 2547 5908
rect 2573 5894 2587 5908
rect 2673 5894 2687 5908
rect 2473 5852 2487 5866
rect 2713 5893 2727 5907
rect 2833 5933 2847 5947
rect 2613 5852 2627 5866
rect 2653 5852 2667 5866
rect 2513 5813 2527 5827
rect 2433 5653 2447 5667
rect 2693 5653 2707 5667
rect 2593 5633 2607 5647
rect 2233 5613 2247 5627
rect 2393 5613 2407 5627
rect 2493 5613 2507 5627
rect 2553 5613 2567 5627
rect 2053 5594 2067 5608
rect 2133 5594 2147 5608
rect 2173 5594 2187 5608
rect 2213 5594 2227 5608
rect 1953 5533 1967 5547
rect 1893 5493 1907 5507
rect 1933 5493 1947 5507
rect 1952 5453 1966 5467
rect 1973 5453 1987 5467
rect 1753 5413 1767 5427
rect 1793 5413 1807 5427
rect 1753 5374 1767 5388
rect 1833 5374 1847 5388
rect 1873 5374 1887 5388
rect 1913 5374 1927 5388
rect 2153 5552 2167 5566
rect 2113 5533 2127 5547
rect 2013 5433 2027 5447
rect 2013 5374 2027 5388
rect 2053 5374 2067 5388
rect 1473 5253 1487 5267
rect 1573 5253 1587 5267
rect 1493 5233 1507 5247
rect 1393 5173 1407 5187
rect 1373 5153 1387 5167
rect 1453 5153 1467 5167
rect 1353 5113 1367 5127
rect 1293 5093 1307 5107
rect 1333 5093 1347 5107
rect 1473 5093 1487 5107
rect 1413 5074 1427 5088
rect 1453 5074 1467 5088
rect 1353 5032 1367 5046
rect 1213 5013 1227 5027
rect 1253 5013 1267 5027
rect 1293 5013 1307 5027
rect 1333 5013 1347 5027
rect 1173 4973 1187 4987
rect 1113 4853 1127 4867
rect 1133 4854 1147 4868
rect 1193 4853 1207 4867
rect 1153 4812 1167 4826
rect 1093 4753 1107 4767
rect 1193 4693 1207 4707
rect 1273 4933 1287 4947
rect 1313 4913 1327 4927
rect 1313 4853 1327 4867
rect 1253 4773 1267 4787
rect 1473 5013 1487 5027
rect 1453 4933 1467 4947
rect 1353 4854 1367 4868
rect 1413 4854 1427 4868
rect 1333 4793 1347 4807
rect 1453 4793 1467 4807
rect 1393 4773 1407 4787
rect 1353 4733 1367 4747
rect 1353 4712 1367 4726
rect 1393 4713 1407 4727
rect 1293 4693 1307 4707
rect 1213 4653 1227 4667
rect 1293 4653 1307 4667
rect 1153 4633 1167 4647
rect 1073 4593 1087 4607
rect 1033 4553 1047 4567
rect 1133 4573 1147 4587
rect 973 4413 987 4427
rect 1033 4513 1047 4527
rect 873 4393 887 4407
rect 953 4393 967 4407
rect 993 4393 1007 4407
rect 853 4373 867 4387
rect 793 4353 807 4367
rect 773 4273 787 4287
rect 713 4233 727 4247
rect 753 4233 767 4247
rect 773 4193 787 4207
rect 693 4133 707 4147
rect 493 4073 507 4087
rect 753 4073 767 4087
rect 493 4034 507 4048
rect 533 4034 547 4048
rect 573 4034 587 4048
rect 673 4034 687 4048
rect 473 3953 487 3967
rect 553 3992 567 4006
rect 513 3973 527 3987
rect 413 3933 427 3947
rect 493 3933 507 3947
rect 373 3873 387 3887
rect 513 3873 527 3887
rect 413 3833 427 3847
rect 293 3813 307 3827
rect 353 3813 367 3827
rect 253 3772 267 3786
rect 313 3733 327 3747
rect 333 3613 347 3627
rect 273 3573 287 3587
rect 233 3513 247 3527
rect 53 3471 67 3485
rect 73 3473 87 3487
rect 33 3433 47 3447
rect 93 3471 107 3485
rect 153 3453 167 3467
rect 113 3393 127 3407
rect 33 3293 47 3307
rect 73 3294 87 3308
rect 153 3293 167 3307
rect 93 3252 107 3266
rect 133 3213 147 3227
rect 233 3453 247 3467
rect 193 3313 207 3327
rect 233 3313 247 3327
rect 593 3833 607 3847
rect 633 3833 647 3847
rect 573 3814 587 3828
rect 393 3772 407 3786
rect 373 3753 387 3767
rect 353 3573 367 3587
rect 513 3772 527 3786
rect 553 3772 567 3786
rect 613 3773 627 3787
rect 593 3713 607 3727
rect 433 3613 447 3627
rect 433 3514 447 3528
rect 493 3514 507 3528
rect 533 3533 547 3547
rect 613 3533 627 3547
rect 713 3973 727 3987
rect 673 3953 687 3967
rect 693 3933 707 3947
rect 673 3913 687 3927
rect 653 3813 667 3827
rect 1093 4512 1107 4526
rect 1053 4473 1067 4487
rect 1213 4573 1227 4587
rect 1253 4554 1267 4568
rect 1313 4554 1327 4568
rect 1393 4633 1407 4647
rect 1533 5193 1547 5207
rect 1533 5093 1547 5107
rect 1653 5233 1667 5247
rect 1613 5153 1627 5167
rect 1613 5074 1627 5088
rect 1653 5074 1667 5088
rect 1593 5032 1607 5046
rect 1573 4993 1587 5007
rect 1553 4893 1567 4907
rect 1593 4973 1607 4987
rect 1793 5313 1807 5327
rect 1773 5253 1787 5267
rect 1753 5113 1767 5127
rect 1753 5074 1767 5088
rect 1673 4993 1687 5007
rect 1653 4913 1667 4927
rect 1733 5032 1747 5046
rect 1773 5033 1787 5047
rect 1753 4993 1767 5007
rect 1733 4953 1747 4967
rect 1713 4933 1727 4947
rect 1693 4893 1707 4907
rect 1593 4853 1607 4867
rect 1653 4854 1667 4868
rect 1533 4812 1547 4826
rect 1633 4773 1647 4787
rect 1553 4753 1567 4767
rect 1593 4753 1607 4767
rect 1493 4673 1507 4687
rect 1713 4813 1727 4827
rect 1613 4673 1627 4687
rect 1673 4673 1687 4687
rect 1593 4633 1607 4647
rect 1513 4554 1527 4568
rect 1553 4554 1567 4568
rect 1172 4512 1186 4526
rect 1193 4512 1207 4526
rect 1233 4512 1247 4526
rect 1153 4453 1167 4467
rect 1233 4473 1247 4487
rect 1173 4433 1187 4447
rect 1112 4413 1126 4427
rect 1133 4413 1147 4427
rect 1093 4353 1107 4367
rect 813 4292 827 4306
rect 1013 4292 1027 4306
rect 1053 4292 1067 4306
rect 1093 4292 1107 4306
rect 933 4273 947 4287
rect 793 4173 807 4187
rect 913 4173 927 4187
rect 893 4133 907 4147
rect 773 4013 787 4027
rect 813 3933 827 3947
rect 753 3893 767 3907
rect 733 3813 747 3827
rect 873 3933 887 3947
rect 853 3913 867 3927
rect 833 3873 847 3887
rect 813 3833 827 3847
rect 673 3772 687 3786
rect 713 3772 727 3786
rect 753 3772 767 3786
rect 673 3713 687 3727
rect 693 3653 707 3667
rect 673 3553 687 3567
rect 633 3514 647 3528
rect 673 3513 687 3527
rect 353 3472 367 3486
rect 433 3473 447 3487
rect 373 3353 387 3367
rect 513 3472 527 3486
rect 673 3473 687 3487
rect 593 3433 607 3447
rect 653 3453 667 3467
rect 413 3333 427 3347
rect 273 3294 287 3308
rect 373 3294 387 3308
rect 533 3353 547 3367
rect 473 3333 487 3347
rect 453 3273 467 3287
rect 193 3213 207 3227
rect 173 3113 187 3127
rect 133 2994 147 3008
rect 173 2994 187 3008
rect 33 2952 47 2966
rect 73 2952 87 2966
rect 113 2952 127 2966
rect 133 2893 147 2907
rect 53 2773 67 2787
rect 93 2774 107 2788
rect 173 2813 187 2827
rect 13 2673 27 2687
rect 153 2732 167 2746
rect 293 3252 307 3266
rect 353 3252 367 3266
rect 393 3252 407 3266
rect 253 3213 267 3227
rect 313 3153 327 3167
rect 213 2994 227 3008
rect 273 2994 287 3008
rect 573 3294 587 3308
rect 753 3593 767 3607
rect 793 3772 807 3786
rect 853 3773 867 3787
rect 833 3733 847 3747
rect 773 3553 787 3567
rect 733 3514 747 3528
rect 833 3514 847 3528
rect 633 3413 647 3427
rect 692 3413 706 3427
rect 713 3413 727 3427
rect 613 3333 627 3347
rect 553 3252 567 3266
rect 613 3252 627 3266
rect 793 3472 807 3486
rect 833 3473 847 3487
rect 893 3853 907 3867
rect 1073 4233 1087 4247
rect 1313 4513 1327 4527
rect 1373 4512 1387 4526
rect 1473 4513 1487 4527
rect 1312 4433 1326 4447
rect 1333 4433 1347 4447
rect 1153 4353 1167 4367
rect 1193 4353 1207 4367
rect 1173 4334 1187 4348
rect 1153 4253 1167 4267
rect 1133 4213 1147 4227
rect 1113 4173 1127 4187
rect 1093 4133 1107 4147
rect 1073 4093 1087 4107
rect 953 4012 967 4026
rect 1013 3973 1027 3987
rect 993 3933 1007 3947
rect 913 3813 927 3827
rect 953 3814 967 3828
rect 1213 4293 1227 4307
rect 1193 4193 1207 4207
rect 1333 4353 1347 4367
rect 1473 4473 1487 4487
rect 1453 4453 1467 4467
rect 1533 4512 1547 4526
rect 1413 4433 1427 4447
rect 1493 4373 1507 4387
rect 1573 4373 1587 4387
rect 1273 4313 1287 4327
rect 1392 4313 1406 4327
rect 1413 4313 1427 4327
rect 1233 4233 1247 4247
rect 1313 4273 1327 4287
rect 1293 4193 1307 4207
rect 1213 4133 1227 4147
rect 1253 4093 1267 4107
rect 1193 4034 1207 4048
rect 1033 3893 1047 3907
rect 1113 3893 1127 3907
rect 893 3772 907 3786
rect 933 3772 947 3786
rect 893 3713 907 3727
rect 873 3653 887 3667
rect 853 3453 867 3467
rect 1193 3933 1207 3947
rect 1173 3893 1187 3907
rect 1153 3853 1167 3867
rect 1093 3814 1107 3828
rect 1133 3814 1147 3828
rect 1053 3773 1067 3787
rect 1113 3753 1127 3767
rect 1173 3753 1187 3767
rect 1033 3713 1047 3727
rect 993 3673 1007 3687
rect 953 3593 967 3607
rect 953 3553 967 3567
rect 913 3514 927 3528
rect 1073 3593 1087 3607
rect 1013 3553 1027 3567
rect 993 3513 1007 3527
rect 893 3473 907 3487
rect 873 3433 887 3447
rect 933 3472 947 3486
rect 973 3453 987 3467
rect 913 3433 927 3447
rect 893 3413 907 3427
rect 753 3393 767 3407
rect 853 3393 867 3407
rect 753 3353 767 3367
rect 713 3333 727 3347
rect 713 3294 727 3308
rect 773 3294 787 3308
rect 813 3294 827 3308
rect 593 3213 607 3227
rect 473 3173 487 3187
rect 433 3153 447 3167
rect 393 3113 407 3127
rect 353 3013 367 3027
rect 293 2952 307 2966
rect 273 2893 287 2907
rect 213 2853 227 2867
rect 253 2853 267 2867
rect 333 2813 347 2827
rect 213 2773 227 2787
rect 293 2774 307 2788
rect 113 2713 127 2727
rect 153 2673 167 2687
rect 53 2593 67 2607
rect 13 2573 27 2587
rect 33 2513 47 2527
rect 73 2474 87 2488
rect 133 2474 147 2488
rect 53 2413 67 2427
rect 33 2373 47 2387
rect 33 2253 47 2267
rect 33 2093 47 2107
rect 33 1853 47 1867
rect 113 2433 127 2447
rect 93 2373 107 2387
rect 233 2732 247 2746
rect 213 2633 227 2647
rect 313 2713 327 2727
rect 293 2673 307 2687
rect 273 2553 287 2567
rect 253 2533 267 2547
rect 213 2513 227 2527
rect 253 2474 267 2488
rect 172 2413 186 2427
rect 193 2413 207 2427
rect 73 2333 87 2347
rect 113 2333 127 2347
rect 193 2333 207 2347
rect 113 2293 127 2307
rect 153 2254 167 2268
rect 93 2212 107 2226
rect 73 2193 87 2207
rect 73 2073 87 2087
rect 253 2373 267 2387
rect 293 2373 307 2387
rect 293 2333 307 2347
rect 253 2293 267 2307
rect 273 2273 287 2287
rect 233 2254 247 2268
rect 493 3053 507 3067
rect 593 3013 607 3027
rect 513 2994 527 3008
rect 553 2994 567 3008
rect 413 2952 427 2966
rect 453 2952 467 2966
rect 493 2953 507 2967
rect 393 2873 407 2887
rect 633 2993 647 3007
rect 573 2952 587 2966
rect 633 2933 647 2947
rect 613 2913 627 2927
rect 573 2893 587 2907
rect 513 2853 527 2867
rect 553 2833 567 2847
rect 493 2813 507 2827
rect 433 2774 447 2788
rect 553 2774 567 2788
rect 593 2774 607 2788
rect 413 2732 427 2746
rect 493 2732 507 2746
rect 353 2713 367 2727
rect 573 2732 587 2746
rect 513 2693 527 2707
rect 333 2673 347 2687
rect 513 2593 527 2607
rect 693 3252 707 3266
rect 713 3233 727 3247
rect 713 3173 727 3187
rect 893 3293 907 3307
rect 873 3252 887 3266
rect 833 3233 847 3247
rect 1153 3713 1167 3727
rect 1113 3553 1127 3567
rect 1033 3453 1047 3467
rect 1093 3433 1107 3447
rect 1173 3593 1187 3607
rect 1013 3393 1027 3407
rect 1153 3393 1167 3407
rect 993 3353 1007 3367
rect 1033 3353 1047 3367
rect 1113 3353 1127 3367
rect 1153 3353 1167 3367
rect 1113 3313 1127 3327
rect 1153 3313 1167 3327
rect 1273 4034 1287 4048
rect 1253 3953 1267 3967
rect 1233 3933 1247 3947
rect 1333 4173 1347 4187
rect 1553 4273 1567 4287
rect 1473 4233 1487 4247
rect 1373 4093 1387 4107
rect 1433 4093 1447 4107
rect 1333 4053 1347 4067
rect 1433 4053 1447 4067
rect 1413 4033 1427 4047
rect 1293 3993 1307 4007
rect 1273 3893 1287 3907
rect 1273 3853 1287 3867
rect 1313 3814 1327 3828
rect 1393 3953 1407 3967
rect 1413 3933 1427 3947
rect 1733 4653 1747 4667
rect 1713 4613 1727 4627
rect 1673 4554 1687 4568
rect 1713 4554 1727 4568
rect 1733 4493 1747 4507
rect 1693 4473 1707 4487
rect 1653 4413 1667 4427
rect 1673 4393 1687 4407
rect 1633 4293 1647 4307
rect 1592 4213 1606 4227
rect 1613 4213 1627 4227
rect 1593 4192 1607 4206
rect 1573 4173 1587 4187
rect 1533 4153 1547 4167
rect 1473 4034 1487 4048
rect 1493 3992 1507 4006
rect 1553 3993 1567 4007
rect 1453 3953 1467 3967
rect 1433 3873 1447 3887
rect 1533 3873 1547 3887
rect 1513 3853 1527 3867
rect 1493 3812 1507 3826
rect 1353 3792 1367 3806
rect 1213 3772 1227 3786
rect 1253 3772 1267 3786
rect 1293 3772 1307 3786
rect 1333 3773 1347 3787
rect 1253 3633 1267 3647
rect 1233 3593 1247 3607
rect 1353 3733 1367 3747
rect 1433 3772 1447 3786
rect 1393 3733 1407 3747
rect 1373 3573 1387 3587
rect 1193 3553 1207 3567
rect 1253 3553 1267 3567
rect 1293 3553 1307 3567
rect 1333 3553 1347 3567
rect 1253 3514 1267 3528
rect 1393 3514 1407 3528
rect 1433 3514 1447 3528
rect 1513 3772 1527 3786
rect 1673 4253 1687 4267
rect 1653 4113 1667 4127
rect 1633 4034 1647 4048
rect 1713 4293 1727 4307
rect 1693 4233 1707 4247
rect 1873 5313 1887 5327
rect 1813 5293 1827 5307
rect 1933 5293 1947 5307
rect 2073 5293 2087 5307
rect 2013 5253 2027 5267
rect 2053 5253 2067 5267
rect 1912 5233 1926 5247
rect 1933 5233 1947 5247
rect 2013 5213 2027 5227
rect 1873 5193 1887 5207
rect 1913 5193 1927 5207
rect 1812 5073 1826 5087
rect 1833 5074 1847 5088
rect 1913 5074 1927 5088
rect 1953 5074 1967 5088
rect 1893 5033 1907 5047
rect 1793 5013 1807 5027
rect 1853 5013 1867 5027
rect 1773 4973 1787 4987
rect 1813 4893 1827 4907
rect 1813 4854 1827 4868
rect 1853 4812 1867 4826
rect 1873 4773 1887 4787
rect 2153 5513 2167 5527
rect 2133 5493 2147 5507
rect 2113 5253 2127 5267
rect 2073 5213 2087 5227
rect 2333 5594 2347 5608
rect 2253 5553 2267 5567
rect 2313 5533 2327 5547
rect 2453 5594 2467 5608
rect 2533 5594 2547 5608
rect 2393 5533 2407 5547
rect 2233 5513 2247 5527
rect 2273 5513 2287 5527
rect 2313 5512 2327 5526
rect 2353 5513 2367 5527
rect 2193 5493 2207 5507
rect 2253 5493 2267 5507
rect 2213 5433 2227 5447
rect 2393 5493 2407 5507
rect 2313 5453 2327 5467
rect 2273 5413 2287 5427
rect 2433 5473 2447 5487
rect 2353 5413 2367 5427
rect 2273 5373 2287 5387
rect 2313 5374 2327 5388
rect 2533 5393 2547 5407
rect 2493 5374 2507 5388
rect 2653 5594 2667 5608
rect 2673 5553 2687 5567
rect 2613 5493 2627 5507
rect 2653 5453 2667 5467
rect 2593 5413 2607 5427
rect 2153 5293 2167 5307
rect 2293 5333 2307 5347
rect 2273 5273 2287 5287
rect 2233 5253 2247 5267
rect 2193 5233 2207 5247
rect 2153 5193 2167 5207
rect 2073 5173 2087 5187
rect 2133 5173 2147 5187
rect 1913 5013 1927 5027
rect 1953 5013 1967 5027
rect 2053 5033 2067 5047
rect 2033 4993 2047 5007
rect 1973 4973 1987 4987
rect 1913 4812 1927 4826
rect 1793 4713 1807 4727
rect 1813 4693 1827 4707
rect 1833 4554 1847 4568
rect 1973 4812 1987 4826
rect 1933 4793 1947 4807
rect 1993 4773 2007 4787
rect 1993 4733 2007 4747
rect 1933 4673 1947 4687
rect 1892 4613 1906 4627
rect 1913 4613 1927 4627
rect 1873 4553 1887 4567
rect 1953 4554 1967 4568
rect 1773 4513 1787 4527
rect 1813 4512 1827 4526
rect 1893 4513 1907 4527
rect 1893 4492 1907 4506
rect 1753 4473 1767 4487
rect 1853 4473 1867 4487
rect 1853 4413 1867 4427
rect 1813 4373 1827 4387
rect 1773 4334 1787 4348
rect 1873 4393 1887 4407
rect 1873 4333 1887 4347
rect 1733 4253 1747 4267
rect 1733 4232 1747 4246
rect 1573 3953 1587 3967
rect 1613 3953 1627 3967
rect 1593 3933 1607 3947
rect 1593 3893 1607 3907
rect 1553 3813 1567 3827
rect 1633 3893 1647 3907
rect 1633 3853 1647 3867
rect 1633 3813 1647 3827
rect 1533 3733 1547 3747
rect 1533 3673 1547 3687
rect 1573 3772 1587 3786
rect 1613 3693 1627 3707
rect 1553 3593 1567 3607
rect 1613 3593 1627 3607
rect 1553 3572 1567 3586
rect 1573 3553 1587 3567
rect 1273 3433 1287 3447
rect 1453 3473 1467 3487
rect 1413 3433 1427 3447
rect 1453 3433 1467 3447
rect 1373 3393 1387 3407
rect 1233 3353 1247 3367
rect 1173 3293 1187 3307
rect 973 3252 987 3266
rect 833 3193 847 3207
rect 913 3193 927 3207
rect 773 3153 787 3167
rect 793 3073 807 3087
rect 753 3053 767 3067
rect 713 3013 727 3027
rect 673 2993 687 3007
rect 792 2993 806 3007
rect 813 2994 827 3008
rect 673 2913 687 2927
rect 813 2933 827 2947
rect 813 2873 827 2887
rect 733 2833 747 2847
rect 773 2793 787 2807
rect 673 2773 687 2787
rect 733 2774 747 2788
rect 673 2653 687 2667
rect 653 2613 667 2627
rect 753 2732 767 2746
rect 1133 3252 1147 3266
rect 1213 3253 1227 3267
rect 1253 3333 1267 3347
rect 1293 3294 1307 3308
rect 1353 3293 1367 3307
rect 1053 3213 1067 3227
rect 1193 3213 1207 3227
rect 953 3113 967 3127
rect 1013 3113 1027 3127
rect 913 3033 927 3047
rect 873 2994 887 3008
rect 1013 3073 1027 3087
rect 953 2993 967 3007
rect 1093 3013 1107 3027
rect 1133 2994 1147 3008
rect 1173 2994 1187 3008
rect 1313 3252 1327 3266
rect 1293 3233 1307 3247
rect 1253 3193 1267 3207
rect 853 2933 867 2947
rect 933 2952 947 2966
rect 893 2873 907 2887
rect 853 2793 867 2807
rect 833 2773 847 2787
rect 1033 2952 1047 2966
rect 1093 2953 1107 2967
rect 1093 2932 1107 2946
rect 1073 2913 1087 2927
rect 1053 2833 1067 2847
rect 973 2813 987 2827
rect 953 2773 967 2787
rect 993 2774 1007 2788
rect 833 2733 847 2747
rect 733 2613 747 2627
rect 813 2613 827 2627
rect 713 2573 727 2587
rect 473 2553 487 2567
rect 633 2553 647 2567
rect 393 2513 407 2527
rect 353 2474 367 2488
rect 453 2473 467 2487
rect 413 2413 427 2427
rect 353 2333 367 2347
rect 393 2333 407 2347
rect 373 2293 387 2307
rect 313 2273 327 2287
rect 353 2273 367 2287
rect 133 2113 147 2127
rect 93 2013 107 2027
rect 113 1954 127 1968
rect 233 2212 247 2226
rect 233 2173 247 2187
rect 213 2133 227 2147
rect 313 2212 327 2226
rect 293 2193 307 2207
rect 193 2113 207 2127
rect 273 2113 287 2127
rect 173 1953 187 1967
rect 113 1893 127 1907
rect 93 1853 107 1867
rect 173 1913 187 1927
rect 133 1853 147 1867
rect 113 1833 127 1847
rect 53 1793 67 1807
rect 53 1733 67 1747
rect 113 1734 127 1748
rect 153 1734 167 1748
rect 333 2173 347 2187
rect 293 2053 307 2067
rect 293 2013 307 2027
rect 253 1954 267 1968
rect 293 1954 307 1968
rect 213 1913 227 1927
rect 193 1893 207 1907
rect 33 1172 47 1186
rect 33 1093 47 1107
rect 33 1013 47 1027
rect 313 1913 327 1927
rect 273 1833 287 1847
rect 233 1793 247 1807
rect 253 1773 267 1787
rect 213 1733 227 1747
rect 713 2552 727 2566
rect 513 2474 527 2488
rect 633 2474 647 2488
rect 673 2474 687 2488
rect 573 2453 587 2467
rect 473 2373 487 2387
rect 453 2273 467 2287
rect 393 2253 407 2267
rect 433 2254 447 2268
rect 533 2373 547 2387
rect 693 2433 707 2447
rect 673 2413 687 2427
rect 613 2373 627 2387
rect 573 2333 587 2347
rect 513 2273 527 2287
rect 673 2273 687 2287
rect 613 2254 627 2268
rect 653 2253 667 2267
rect 373 2212 387 2226
rect 413 2212 427 2226
rect 433 2193 447 2207
rect 393 1973 407 1987
rect 353 1953 367 1967
rect 513 2212 527 2226
rect 453 2153 467 2167
rect 553 2212 567 2226
rect 593 2173 607 2187
rect 593 2113 607 2127
rect 593 2053 607 2067
rect 533 2013 547 2027
rect 493 1973 507 1987
rect 433 1954 447 1968
rect 533 1954 547 1968
rect 353 1913 367 1927
rect 613 2013 627 2027
rect 333 1853 347 1867
rect 313 1753 327 1767
rect 293 1734 307 1748
rect 133 1692 147 1706
rect 193 1692 207 1706
rect 273 1692 287 1706
rect 93 1573 107 1587
rect 153 1553 167 1567
rect 333 1553 347 1567
rect 113 1513 127 1527
rect 213 1513 227 1527
rect 253 1493 267 1507
rect 313 1493 327 1507
rect 233 1392 247 1406
rect 133 1353 147 1367
rect 113 1313 127 1327
rect 93 1233 107 1247
rect 333 1392 347 1406
rect 313 1353 327 1367
rect 313 1332 327 1346
rect 193 1253 207 1267
rect 273 1253 287 1267
rect 153 1214 167 1228
rect 253 1214 267 1228
rect 53 993 67 1007
rect 93 1172 107 1186
rect 133 1172 147 1186
rect 193 1172 207 1186
rect 233 1172 247 1186
rect 413 1912 427 1926
rect 513 1912 527 1926
rect 373 1893 387 1907
rect 593 1912 607 1926
rect 553 1873 567 1887
rect 433 1833 447 1847
rect 493 1753 507 1767
rect 553 1753 567 1767
rect 373 1693 387 1707
rect 573 1734 587 1748
rect 413 1692 427 1706
rect 453 1692 467 1706
rect 493 1692 507 1706
rect 373 1633 387 1647
rect 393 1593 407 1607
rect 433 1673 447 1687
rect 413 1573 427 1587
rect 473 1553 487 1567
rect 433 1513 447 1527
rect 433 1434 447 1448
rect 353 1313 367 1327
rect 593 1693 607 1707
rect 593 1593 607 1607
rect 553 1453 567 1467
rect 513 1434 527 1448
rect 713 2413 727 2427
rect 713 2373 727 2387
rect 693 2253 707 2267
rect 1013 2732 1027 2746
rect 973 2713 987 2727
rect 913 2693 927 2707
rect 993 2673 1007 2687
rect 873 2593 887 2607
rect 833 2553 847 2567
rect 753 2513 767 2527
rect 813 2513 827 2527
rect 753 2393 767 2407
rect 733 2353 747 2367
rect 793 2353 807 2367
rect 853 2393 867 2407
rect 833 2293 847 2307
rect 753 2273 767 2287
rect 833 2272 847 2286
rect 693 2213 707 2227
rect 773 2212 787 2226
rect 693 2173 707 2187
rect 733 2173 747 2187
rect 973 2553 987 2567
rect 893 2533 907 2547
rect 933 2513 947 2527
rect 1033 2533 1047 2547
rect 1013 2474 1027 2488
rect 1193 2952 1207 2966
rect 1133 2873 1147 2887
rect 1153 2873 1167 2887
rect 1093 2773 1107 2787
rect 1173 2793 1187 2807
rect 1113 2732 1127 2746
rect 1073 2673 1087 2687
rect 1153 2673 1167 2687
rect 1113 2533 1127 2547
rect 1173 2533 1187 2547
rect 1133 2513 1147 2527
rect 893 2393 907 2407
rect 1053 2474 1067 2488
rect 1033 2433 1047 2447
rect 1013 2413 1027 2427
rect 913 2333 927 2347
rect 953 2333 967 2347
rect 873 2273 887 2287
rect 953 2312 967 2326
rect 853 2173 867 2187
rect 773 2133 787 2147
rect 693 2013 707 2027
rect 773 2013 787 2027
rect 632 1953 646 1967
rect 653 1954 667 1968
rect 793 1993 807 2007
rect 893 2212 907 2226
rect 933 2213 947 2227
rect 893 2033 907 2047
rect 773 1973 787 1987
rect 753 1953 767 1967
rect 633 1913 647 1927
rect 673 1912 687 1926
rect 713 1833 727 1847
rect 713 1793 727 1807
rect 633 1733 647 1747
rect 673 1734 687 1748
rect 813 1954 827 1968
rect 853 1954 867 1968
rect 913 1993 927 2007
rect 893 1953 907 1967
rect 793 1913 807 1927
rect 773 1873 787 1887
rect 873 1912 887 1926
rect 913 1913 927 1927
rect 853 1893 867 1907
rect 833 1873 847 1887
rect 853 1813 867 1827
rect 793 1753 807 1767
rect 873 1753 887 1767
rect 753 1734 767 1748
rect 813 1734 827 1748
rect 653 1692 667 1706
rect 733 1692 747 1706
rect 753 1673 767 1687
rect 793 1673 807 1687
rect 693 1633 707 1647
rect 713 1473 727 1487
rect 653 1453 667 1467
rect 633 1434 647 1448
rect 693 1453 707 1467
rect 473 1333 487 1347
rect 493 1293 507 1307
rect 333 1213 347 1227
rect 373 1214 387 1228
rect 413 1214 427 1228
rect 533 1273 547 1287
rect 553 1233 567 1247
rect 93 1053 107 1067
rect 153 993 167 1007
rect 73 933 87 947
rect 313 993 327 1007
rect 253 953 267 967
rect 213 933 227 947
rect 193 913 207 927
rect 53 853 67 867
rect 53 753 67 767
rect 33 713 47 727
rect 173 873 187 887
rect 133 853 147 867
rect 113 733 127 747
rect 93 713 107 727
rect 233 872 247 886
rect 313 872 327 886
rect 273 773 287 787
rect 193 733 207 747
rect 173 694 187 708
rect 53 652 67 666
rect 93 652 107 666
rect 33 613 47 627
rect 133 613 147 627
rect 113 473 127 487
rect 153 413 167 427
rect 393 1133 407 1147
rect 473 1173 487 1187
rect 433 1073 447 1087
rect 393 1053 407 1067
rect 413 1013 427 1027
rect 393 933 407 947
rect 373 914 387 928
rect 353 873 367 887
rect 513 1172 527 1186
rect 633 1253 647 1267
rect 693 1373 707 1387
rect 673 1353 687 1367
rect 713 1353 727 1367
rect 673 1332 687 1346
rect 653 1233 667 1247
rect 873 1692 887 1706
rect 833 1553 847 1567
rect 813 1473 827 1487
rect 873 1453 887 1467
rect 833 1392 847 1406
rect 873 1392 887 1406
rect 913 1793 927 1807
rect 1053 2413 1067 2427
rect 1033 2313 1047 2327
rect 1193 2493 1207 2507
rect 1233 2873 1247 2887
rect 1353 3153 1367 3167
rect 1313 2994 1327 3008
rect 1293 2913 1307 2927
rect 1373 3053 1387 3067
rect 1373 2953 1387 2967
rect 1333 2873 1347 2887
rect 1253 2833 1267 2847
rect 1333 2813 1347 2827
rect 1293 2774 1307 2788
rect 1273 2613 1287 2627
rect 1313 2593 1327 2607
rect 1573 3514 1587 3528
rect 1473 3393 1487 3407
rect 1433 3294 1447 3308
rect 1473 3294 1487 3308
rect 1553 3472 1567 3486
rect 1713 4093 1727 4107
rect 1693 3893 1707 3907
rect 1693 3853 1707 3867
rect 1673 3813 1687 3827
rect 1833 4292 1847 4306
rect 1913 4473 1927 4487
rect 1893 4233 1907 4247
rect 1793 4073 1807 4087
rect 1973 4413 1987 4427
rect 2113 5113 2127 5127
rect 2193 5173 2207 5187
rect 2153 5074 2167 5088
rect 2313 5313 2327 5327
rect 2293 5233 2307 5247
rect 2193 4993 2207 5007
rect 2293 5033 2307 5047
rect 2133 4973 2147 4987
rect 2253 4973 2267 4987
rect 2293 4953 2307 4967
rect 2073 4893 2087 4907
rect 2153 4893 2167 4907
rect 2073 4812 2087 4826
rect 2113 4773 2127 4787
rect 2133 4753 2147 4767
rect 2113 4713 2127 4727
rect 2093 4693 2107 4707
rect 2053 4554 2067 4568
rect 2413 5333 2427 5347
rect 2453 5333 2467 5347
rect 2333 5293 2347 5307
rect 2433 5293 2447 5307
rect 2333 5233 2347 5247
rect 2353 5093 2367 5107
rect 2393 5093 2407 5107
rect 2333 5053 2347 5067
rect 2473 5273 2487 5287
rect 2573 5293 2587 5307
rect 2552 5253 2566 5267
rect 2573 5253 2587 5267
rect 2513 5153 2527 5167
rect 2613 5393 2627 5407
rect 2673 5393 2687 5407
rect 2773 5852 2787 5866
rect 3033 6072 3047 6086
rect 3073 6072 3087 6086
rect 2993 6033 3007 6047
rect 2973 5913 2987 5927
rect 3213 6072 3227 6086
rect 3033 5894 3047 5908
rect 2993 5873 3007 5887
rect 2873 5852 2887 5866
rect 2733 5793 2747 5807
rect 2853 5793 2867 5807
rect 2833 5713 2847 5727
rect 2753 5633 2767 5647
rect 2733 5593 2747 5607
rect 2793 5594 2807 5608
rect 2773 5552 2787 5566
rect 2793 5533 2807 5547
rect 2713 5413 2727 5427
rect 2713 5374 2727 5388
rect 2753 5374 2767 5388
rect 2853 5693 2867 5707
rect 2913 5813 2927 5827
rect 3153 5913 3167 5927
rect 3193 5894 3207 5908
rect 3133 5852 3147 5866
rect 3173 5852 3187 5866
rect 3053 5753 3067 5767
rect 3093 5753 3107 5767
rect 2913 5693 2927 5707
rect 3013 5693 3027 5707
rect 2953 5594 2967 5608
rect 2993 5594 3007 5608
rect 2873 5533 2887 5547
rect 2953 5533 2967 5547
rect 2933 5493 2947 5507
rect 2873 5453 2887 5467
rect 2853 5433 2867 5447
rect 2633 5332 2647 5346
rect 2673 5332 2687 5346
rect 2653 5293 2667 5307
rect 2613 5253 2627 5267
rect 2613 5193 2627 5207
rect 2593 5173 2607 5187
rect 2513 5113 2527 5127
rect 2573 5113 2587 5127
rect 2553 5074 2567 5088
rect 2673 5153 2687 5167
rect 2813 5332 2827 5346
rect 2893 5374 2907 5388
rect 3093 5633 3107 5647
rect 3133 5633 3147 5647
rect 3013 5513 3027 5527
rect 3053 5513 3067 5527
rect 2993 5453 3007 5467
rect 3033 5453 3047 5467
rect 3033 5373 3047 5387
rect 2773 5313 2787 5327
rect 2773 5213 2787 5227
rect 2713 5193 2727 5207
rect 2753 5173 2767 5187
rect 2633 5113 2647 5127
rect 2693 5113 2707 5127
rect 2613 5093 2627 5107
rect 2613 5072 2627 5086
rect 2453 5032 2467 5046
rect 2353 5013 2367 5027
rect 2413 5013 2427 5027
rect 2413 4973 2427 4987
rect 2393 4913 2407 4927
rect 2353 4893 2367 4907
rect 2213 4854 2227 4868
rect 2273 4853 2287 4867
rect 2193 4812 2207 4826
rect 2233 4812 2247 4826
rect 2333 4873 2347 4887
rect 2433 4893 2447 4907
rect 2293 4812 2307 4826
rect 2253 4733 2267 4747
rect 2193 4673 2207 4687
rect 2153 4573 2167 4587
rect 2133 4554 2147 4568
rect 2113 4512 2127 4526
rect 1993 4353 2007 4367
rect 1733 4053 1747 4067
rect 1873 4053 1887 4067
rect 1913 4054 1927 4068
rect 1973 4273 1987 4287
rect 1993 4213 2007 4227
rect 1973 4193 1987 4207
rect 1813 4034 1827 4048
rect 1793 3992 1807 4006
rect 1773 3973 1787 3987
rect 1793 3953 1807 3967
rect 1833 3953 1847 3967
rect 1773 3933 1787 3947
rect 1753 3913 1767 3927
rect 1753 3873 1767 3887
rect 1733 3853 1747 3867
rect 1713 3833 1727 3847
rect 1913 4033 1927 4047
rect 1893 3992 1907 4006
rect 1973 4034 1987 4048
rect 2073 4473 2087 4487
rect 2173 4513 2187 4527
rect 2213 4573 2227 4587
rect 2193 4493 2207 4507
rect 2172 4473 2186 4487
rect 2193 4472 2207 4486
rect 2153 4453 2167 4467
rect 2133 4393 2147 4407
rect 2073 4273 2087 4287
rect 2093 4233 2107 4247
rect 2053 4113 2067 4127
rect 1853 3933 1867 3947
rect 1893 3873 1907 3887
rect 1853 3853 1867 3867
rect 1773 3813 1787 3827
rect 1913 3853 1927 3867
rect 1893 3813 1907 3827
rect 1673 3772 1687 3786
rect 1713 3772 1727 3786
rect 1773 3773 1787 3787
rect 1693 3751 1707 3765
rect 1673 3733 1687 3747
rect 1753 3732 1767 3746
rect 1653 3653 1667 3667
rect 1713 3653 1727 3667
rect 1653 3632 1667 3646
rect 1733 3613 1747 3627
rect 1833 3772 1847 3786
rect 2053 4034 2067 4048
rect 2193 4233 2207 4247
rect 2113 4113 2127 4127
rect 1973 3953 1987 3967
rect 2093 3993 2107 4007
rect 2033 3933 2047 3947
rect 2013 3853 2027 3867
rect 1933 3812 1947 3826
rect 1973 3814 1987 3828
rect 1793 3733 1807 3747
rect 1833 3733 1847 3747
rect 1773 3713 1787 3727
rect 1913 3753 1927 3767
rect 1793 3693 1807 3707
rect 1833 3693 1847 3707
rect 1813 3673 1827 3687
rect 1753 3593 1767 3607
rect 1733 3573 1747 3587
rect 1713 3533 1727 3547
rect 1673 3514 1687 3528
rect 1533 3373 1547 3387
rect 1613 3373 1627 3387
rect 1513 3293 1527 3307
rect 1413 3133 1427 3147
rect 1493 3252 1507 3266
rect 1493 3193 1507 3207
rect 1453 3113 1467 3127
rect 1453 2994 1467 3008
rect 1493 2994 1507 3008
rect 1433 2952 1447 2966
rect 1513 2953 1527 2967
rect 1393 2913 1407 2927
rect 1473 2913 1487 2927
rect 1493 2793 1507 2807
rect 1553 3333 1567 3347
rect 1613 3333 1627 3347
rect 1573 3252 1587 3266
rect 1653 3472 1667 3486
rect 1773 3514 1787 3528
rect 1873 3653 1887 3667
rect 1853 3553 1867 3567
rect 1733 3493 1747 3507
rect 1713 3453 1727 3467
rect 1773 3453 1787 3467
rect 1653 3433 1667 3447
rect 1733 3433 1747 3447
rect 1753 3333 1767 3347
rect 1653 3313 1667 3327
rect 1713 3313 1727 3327
rect 1653 3292 1667 3306
rect 1833 3472 1847 3486
rect 1793 3433 1807 3447
rect 1793 3313 1807 3327
rect 1773 3293 1787 3307
rect 1673 3253 1687 3267
rect 1653 3193 1667 3207
rect 1673 3173 1687 3187
rect 1713 3213 1727 3227
rect 1633 3133 1647 3147
rect 1693 3133 1707 3147
rect 1773 3253 1787 3267
rect 1733 3193 1747 3207
rect 1713 3113 1727 3127
rect 1673 3093 1687 3107
rect 1613 3073 1627 3087
rect 1753 3073 1767 3087
rect 1672 3053 1686 3067
rect 1693 3053 1707 3067
rect 1613 3033 1627 3047
rect 1727 3013 1741 3027
rect 1693 2993 1707 3007
rect 1793 3193 1807 3207
rect 1773 3053 1787 3067
rect 1893 3593 1907 3607
rect 1993 3772 2007 3786
rect 2033 3753 2047 3767
rect 1953 3693 1967 3707
rect 1973 3633 1987 3647
rect 1953 3613 1967 3627
rect 1913 3573 1927 3587
rect 1893 3513 1907 3527
rect 2093 3953 2107 3967
rect 2093 3753 2107 3767
rect 2133 4053 2147 4067
rect 2173 4113 2187 4127
rect 2413 4813 2427 4827
rect 2373 4793 2387 4807
rect 2393 4733 2407 4747
rect 2353 4693 2367 4707
rect 2333 4653 2347 4667
rect 2293 4613 2307 4627
rect 2293 4473 2307 4487
rect 2293 4413 2307 4427
rect 2253 4133 2267 4147
rect 2253 4112 2267 4126
rect 2213 4053 2227 4067
rect 2153 4034 2167 4048
rect 2213 4032 2227 4046
rect 2433 4713 2447 4727
rect 2413 4693 2427 4707
rect 2393 4653 2407 4667
rect 2433 4613 2447 4627
rect 2373 4593 2387 4607
rect 2353 4554 2367 4568
rect 2493 5032 2507 5046
rect 2573 5032 2587 5046
rect 2473 4913 2487 4927
rect 2512 4913 2526 4927
rect 2533 4913 2547 4927
rect 2593 4913 2607 4927
rect 2613 4893 2627 4907
rect 2593 4873 2607 4887
rect 2613 4793 2627 4807
rect 2533 4753 2547 4767
rect 2533 4593 2547 4607
rect 2613 4593 2627 4607
rect 2453 4533 2467 4547
rect 2353 4493 2367 4507
rect 2453 4453 2467 4467
rect 2473 4433 2487 4447
rect 2433 4413 2447 4427
rect 2493 4413 2507 4427
rect 2533 4413 2547 4427
rect 2413 4393 2427 4407
rect 2453 4373 2467 4387
rect 2433 4353 2447 4367
rect 2353 4333 2367 4347
rect 2413 4333 2427 4347
rect 2693 5074 2707 5088
rect 2713 5032 2727 5046
rect 2853 5332 2867 5346
rect 2873 5333 2887 5347
rect 2953 5333 2967 5347
rect 2873 5273 2887 5287
rect 2833 5093 2847 5107
rect 2813 5074 2827 5088
rect 2913 5313 2927 5327
rect 2893 5253 2907 5267
rect 2933 5253 2947 5267
rect 2913 5193 2927 5207
rect 2813 5013 2827 5027
rect 2793 4893 2807 4907
rect 2753 4853 2767 4867
rect 2673 4812 2687 4826
rect 2713 4812 2727 4826
rect 2693 4653 2707 4667
rect 2653 4593 2667 4607
rect 2753 4812 2767 4826
rect 2733 4633 2747 4647
rect 2653 4433 2667 4447
rect 2693 4433 2707 4447
rect 2633 4393 2647 4407
rect 2373 4213 2387 4227
rect 2293 4073 2307 4087
rect 2333 4073 2347 4087
rect 2333 4034 2347 4048
rect 2133 3953 2147 3967
rect 2173 3873 2187 3887
rect 2233 3913 2247 3927
rect 2213 3833 2227 3847
rect 2353 3993 2367 4007
rect 2273 3873 2287 3887
rect 2253 3833 2267 3847
rect 2193 3813 2207 3827
rect 2233 3813 2247 3827
rect 2192 3772 2206 3786
rect 2213 3772 2227 3786
rect 2153 3753 2167 3767
rect 2092 3713 2106 3727
rect 2113 3713 2127 3727
rect 2033 3513 2047 3527
rect 2213 3751 2227 3765
rect 2133 3693 2147 3707
rect 2153 3653 2167 3667
rect 1833 3433 1847 3447
rect 1873 3433 1887 3447
rect 1953 3472 1967 3486
rect 1933 3413 1947 3427
rect 1893 3373 1907 3387
rect 1873 3353 1887 3367
rect 1833 3293 1847 3307
rect 1913 3294 1927 3308
rect 2053 3453 2067 3467
rect 2033 3413 2047 3427
rect 2013 3393 2027 3407
rect 1993 3373 2007 3387
rect 2013 3353 2027 3367
rect 2013 3332 2027 3346
rect 2133 3473 2147 3487
rect 2113 3453 2127 3467
rect 2133 3433 2147 3447
rect 2073 3393 2087 3407
rect 2193 3573 2207 3587
rect 2413 4293 2427 4307
rect 2673 4393 2687 4407
rect 2733 4413 2747 4427
rect 2713 4393 2727 4407
rect 2693 4353 2707 4367
rect 2733 4373 2747 4387
rect 2913 5033 2927 5047
rect 3033 5333 3047 5347
rect 3013 5233 3027 5247
rect 3193 5813 3207 5827
rect 3173 5594 3187 5608
rect 3233 5793 3247 5807
rect 3233 5753 3247 5767
rect 3233 5673 3247 5687
rect 3373 6173 3387 6187
rect 3293 6133 3307 6147
rect 3333 6133 3347 6147
rect 3453 6114 3467 6128
rect 3493 6114 3507 6128
rect 3713 6153 3727 6167
rect 3813 6153 3827 6167
rect 3573 6114 3587 6128
rect 3613 6114 3627 6128
rect 3653 6114 3667 6128
rect 3293 6073 3307 6087
rect 3393 6033 3407 6047
rect 3453 6033 3467 6047
rect 3493 5973 3507 5987
rect 3273 5933 3287 5947
rect 3353 5933 3367 5947
rect 3333 5894 3347 5908
rect 3373 5894 3387 5908
rect 3453 5894 3467 5908
rect 3553 5993 3567 6007
rect 3513 5913 3527 5927
rect 3673 6072 3687 6086
rect 3773 6114 3787 6128
rect 3633 6033 3647 6047
rect 3713 6033 3727 6047
rect 3773 6013 3787 6027
rect 3573 5973 3587 5987
rect 3753 5973 3767 5987
rect 3613 5913 3627 5927
rect 3673 5913 3687 5927
rect 3693 5893 3707 5907
rect 3793 5993 3807 6007
rect 3673 5873 3687 5887
rect 3313 5852 3327 5866
rect 3353 5852 3367 5866
rect 3353 5831 3367 5845
rect 3273 5773 3287 5787
rect 3333 5733 3347 5747
rect 3253 5633 3267 5647
rect 3393 5813 3407 5827
rect 3413 5793 3427 5807
rect 3373 5713 3387 5727
rect 3353 5653 3367 5667
rect 3273 5593 3287 5607
rect 3333 5594 3347 5608
rect 3213 5552 3227 5566
rect 3173 5493 3187 5507
rect 3133 5473 3147 5487
rect 3073 5453 3087 5467
rect 3233 5473 3247 5487
rect 3213 5433 3227 5447
rect 3193 5413 3207 5427
rect 3133 5393 3147 5407
rect 3173 5393 3187 5407
rect 3153 5332 3167 5346
rect 3193 5333 3207 5347
rect 3093 5273 3107 5287
rect 3213 5273 3227 5287
rect 3173 5233 3187 5247
rect 3213 5233 3227 5247
rect 3053 5213 3067 5227
rect 2973 5173 2987 5187
rect 3013 5173 3027 5187
rect 2973 5152 2987 5166
rect 2973 5074 2987 5088
rect 3013 5074 3027 5088
rect 2933 4973 2947 4987
rect 2833 4953 2847 4967
rect 2833 4893 2847 4907
rect 2833 4854 2847 4868
rect 2873 4854 2887 4868
rect 2793 4813 2807 4827
rect 2853 4812 2867 4826
rect 2893 4733 2907 4747
rect 2873 4633 2887 4647
rect 2813 4554 2827 4568
rect 2833 4512 2847 4526
rect 2813 4493 2827 4507
rect 2793 4433 2807 4447
rect 2773 4393 2787 4407
rect 2793 4373 2807 4387
rect 2753 4334 2767 4348
rect 2793 4333 2807 4347
rect 2913 4693 2927 4707
rect 2993 5032 3007 5046
rect 3113 5153 3127 5167
rect 3153 5153 3167 5167
rect 3053 5013 3067 5027
rect 2953 4953 2967 4967
rect 3053 4953 3067 4967
rect 2993 4893 3007 4907
rect 3053 4893 3067 4907
rect 3033 4854 3047 4868
rect 2973 4793 2987 4807
rect 2933 4633 2947 4647
rect 2933 4593 2947 4607
rect 2953 4573 2967 4587
rect 2893 4553 2907 4567
rect 3033 4793 3047 4807
rect 3013 4713 3027 4727
rect 3033 4693 3047 4707
rect 3013 4573 3027 4587
rect 2873 4453 2887 4467
rect 2913 4512 2927 4526
rect 2953 4512 2967 4526
rect 3013 4512 3027 4526
rect 2913 4473 2927 4487
rect 3093 5032 3107 5046
rect 3173 5032 3187 5046
rect 3173 4933 3187 4947
rect 3133 4913 3147 4927
rect 3313 5552 3327 5566
rect 3333 5513 3347 5527
rect 3273 5433 3287 5447
rect 3293 5393 3307 5407
rect 3353 5473 3367 5487
rect 3393 5473 3407 5487
rect 3353 5452 3367 5466
rect 3333 5373 3347 5387
rect 3253 5333 3267 5347
rect 3313 5332 3327 5346
rect 3333 5233 3347 5247
rect 3253 5193 3267 5207
rect 3273 5133 3287 5147
rect 3293 5074 3307 5088
rect 3373 5393 3387 5407
rect 3513 5852 3527 5866
rect 3553 5853 3567 5867
rect 3553 5813 3567 5827
rect 3473 5773 3487 5787
rect 3433 5653 3447 5667
rect 3513 5653 3527 5667
rect 3473 5594 3487 5608
rect 3633 5852 3647 5866
rect 3693 5852 3707 5866
rect 3593 5773 3607 5787
rect 3593 5752 3607 5766
rect 3553 5594 3567 5608
rect 3433 5533 3447 5547
rect 3413 5393 3427 5407
rect 3472 5493 3486 5507
rect 3493 5493 3507 5507
rect 3493 5472 3507 5486
rect 3573 5553 3587 5567
rect 3553 5533 3567 5547
rect 3533 5453 3547 5467
rect 3533 5413 3547 5427
rect 3493 5393 3507 5407
rect 3533 5373 3547 5387
rect 3573 5473 3587 5487
rect 3593 5453 3607 5467
rect 3653 5773 3667 5787
rect 3793 5852 3807 5866
rect 3693 5713 3707 5727
rect 3673 5653 3687 5667
rect 3693 5594 3707 5608
rect 3633 5553 3647 5567
rect 3673 5552 3687 5566
rect 3653 5513 3667 5527
rect 3633 5492 3647 5506
rect 3633 5433 3647 5447
rect 3593 5374 3607 5388
rect 3373 5333 3387 5347
rect 3353 5213 3367 5227
rect 3273 5032 3287 5046
rect 3353 5032 3367 5046
rect 3313 5013 3327 5027
rect 3213 4953 3227 4967
rect 3193 4893 3207 4907
rect 3153 4854 3167 4868
rect 3073 4653 3087 4667
rect 3093 4593 3107 4607
rect 3093 4553 3107 4567
rect 3193 4812 3207 4826
rect 3173 4793 3187 4807
rect 3233 4853 3247 4867
rect 3153 4553 3167 4567
rect 3073 4512 3087 4526
rect 3133 4493 3147 4507
rect 2933 4433 2947 4447
rect 3033 4433 3047 4447
rect 2913 4373 2927 4387
rect 2893 4333 2907 4347
rect 2693 4293 2707 4307
rect 2653 4273 2667 4287
rect 2493 4253 2507 4267
rect 2433 4133 2447 4147
rect 2473 4093 2487 4107
rect 2473 4053 2487 4067
rect 2332 3813 2346 3827
rect 2353 3814 2367 3828
rect 2273 3773 2287 3787
rect 2312 3772 2326 3786
rect 2333 3773 2347 3787
rect 2373 3753 2387 3767
rect 2293 3733 2307 3747
rect 2333 3733 2347 3747
rect 2273 3573 2287 3587
rect 2233 3514 2247 3528
rect 2313 3713 2327 3727
rect 2293 3513 2307 3527
rect 2293 3473 2307 3487
rect 2253 3433 2267 3447
rect 2273 3413 2287 3427
rect 2213 3393 2227 3407
rect 2253 3393 2267 3407
rect 2193 3333 2207 3347
rect 2053 3313 2067 3327
rect 2153 3313 2167 3327
rect 1953 3294 1967 3308
rect 2013 3294 2027 3308
rect 2133 3294 2147 3308
rect 1833 3253 1847 3267
rect 1813 3013 1827 3027
rect 1573 2953 1587 2967
rect 1553 2933 1567 2947
rect 1553 2873 1567 2887
rect 1553 2813 1567 2827
rect 1433 2774 1447 2788
rect 1533 2773 1547 2787
rect 1493 2732 1507 2746
rect 1533 2733 1547 2747
rect 1453 2693 1467 2707
rect 1413 2673 1427 2687
rect 1393 2573 1407 2587
rect 1373 2553 1387 2567
rect 1253 2493 1267 2507
rect 1233 2473 1247 2487
rect 1313 2474 1327 2488
rect 1093 2393 1107 2407
rect 1133 2393 1147 2407
rect 1113 2373 1127 2387
rect 1153 2373 1167 2387
rect 1072 2353 1086 2367
rect 1093 2353 1107 2367
rect 1013 2254 1027 2268
rect 1053 2254 1067 2268
rect 973 2213 987 2227
rect 1073 2173 1087 2187
rect 1333 2432 1347 2446
rect 1373 2433 1387 2447
rect 1373 2393 1387 2407
rect 1233 2373 1247 2387
rect 1333 2333 1347 2347
rect 1173 2313 1187 2327
rect 1273 2313 1287 2327
rect 1153 2293 1167 2307
rect 1193 2293 1207 2307
rect 1173 2254 1187 2268
rect 1213 2254 1227 2268
rect 1333 2254 1347 2268
rect 1413 2513 1427 2527
rect 1393 2333 1407 2347
rect 1493 2493 1507 2507
rect 1413 2313 1427 2327
rect 1693 2953 1707 2967
rect 1633 2933 1647 2947
rect 1673 2893 1687 2907
rect 1633 2873 1647 2887
rect 1613 2853 1627 2867
rect 1593 2813 1607 2827
rect 1653 2833 1667 2847
rect 1573 2773 1587 2787
rect 1573 2733 1587 2747
rect 1613 2732 1627 2746
rect 1553 2573 1567 2587
rect 1573 2553 1587 2567
rect 1513 2413 1527 2427
rect 1473 2353 1487 2367
rect 1553 2353 1567 2367
rect 1453 2333 1467 2347
rect 1433 2273 1447 2287
rect 1493 2273 1507 2287
rect 1153 2173 1167 2187
rect 1233 2212 1247 2226
rect 1273 2212 1287 2226
rect 1313 2212 1327 2226
rect 1313 2173 1327 2187
rect 1113 2153 1127 2167
rect 1193 2153 1207 2167
rect 1273 2153 1287 2167
rect 1313 2113 1327 2127
rect 1033 2053 1047 2067
rect 993 1993 1007 2007
rect 953 1954 967 1968
rect 1373 2193 1387 2207
rect 1353 2033 1367 2047
rect 1153 1973 1167 1987
rect 1313 1973 1327 1987
rect 1033 1954 1047 1968
rect 973 1912 987 1926
rect 1013 1912 1027 1926
rect 953 1793 967 1807
rect 933 1733 947 1747
rect 1113 1954 1127 1968
rect 1233 1954 1247 1968
rect 1273 1954 1287 1968
rect 1173 1912 1187 1926
rect 1073 1873 1087 1887
rect 1133 1873 1147 1887
rect 1073 1813 1087 1827
rect 993 1734 1007 1748
rect 973 1692 987 1706
rect 1093 1692 1107 1706
rect 1353 1953 1367 1967
rect 1253 1813 1267 1827
rect 1153 1773 1167 1787
rect 1013 1673 1027 1687
rect 1133 1673 1147 1687
rect 993 1593 1007 1607
rect 1033 1593 1047 1607
rect 993 1553 1007 1567
rect 913 1473 927 1487
rect 953 1453 967 1467
rect 793 1353 807 1367
rect 853 1293 867 1307
rect 713 1273 727 1287
rect 753 1273 767 1287
rect 813 1253 827 1267
rect 733 1213 747 1227
rect 773 1214 787 1228
rect 853 1213 867 1227
rect 613 1172 627 1186
rect 653 1172 667 1186
rect 713 1172 727 1186
rect 553 1133 567 1147
rect 353 773 367 787
rect 473 872 487 886
rect 533 872 547 886
rect 573 872 587 886
rect 653 1133 667 1147
rect 633 933 647 947
rect 433 833 447 847
rect 613 833 627 847
rect 393 753 407 767
rect 393 694 407 708
rect 433 694 447 708
rect 493 693 507 707
rect 313 652 327 666
rect 353 652 367 666
rect 413 633 427 647
rect 353 613 367 627
rect 453 613 467 627
rect 273 573 287 587
rect 413 493 427 507
rect 253 473 267 487
rect 213 413 227 427
rect 193 393 207 407
rect 313 413 327 427
rect 133 352 147 366
rect 233 313 247 327
rect 93 273 107 287
rect 133 273 147 287
rect 13 233 27 247
rect 93 233 107 247
rect 493 433 507 447
rect 533 753 547 767
rect 573 773 587 787
rect 553 733 567 747
rect 533 693 547 707
rect 613 733 627 747
rect 633 693 647 707
rect 553 652 567 666
rect 593 633 607 647
rect 593 573 607 587
rect 553 493 567 507
rect 513 394 527 408
rect 613 433 627 447
rect 433 352 447 366
rect 313 313 327 327
rect 393 313 407 327
rect 273 233 287 247
rect 253 213 267 227
rect 573 352 587 366
rect 533 293 547 307
rect 493 273 507 287
rect 413 233 427 247
rect 393 193 407 207
rect 273 173 287 187
rect 313 173 327 187
rect 373 174 387 188
rect 413 174 427 188
rect 533 253 547 267
rect 113 132 127 146
rect 153 132 167 146
rect 233 132 247 146
rect 353 132 367 146
rect 393 132 407 146
rect 473 113 487 127
rect 633 394 647 408
rect 633 353 647 367
rect 693 914 707 928
rect 793 1172 807 1186
rect 833 1172 847 1186
rect 953 1373 967 1387
rect 933 1353 947 1367
rect 913 1214 927 1228
rect 1013 1333 1027 1347
rect 973 1253 987 1267
rect 933 1153 947 1167
rect 873 1133 887 1147
rect 853 1093 867 1107
rect 833 1073 847 1087
rect 853 1053 867 1067
rect 773 953 787 967
rect 853 933 867 947
rect 893 914 907 928
rect 773 873 787 887
rect 993 1173 1007 1187
rect 833 872 847 886
rect 933 872 947 886
rect 813 833 827 847
rect 873 833 887 847
rect 793 773 807 787
rect 713 753 727 767
rect 753 733 767 747
rect 673 693 687 707
rect 973 1033 987 1047
rect 1073 1513 1087 1527
rect 1053 1473 1067 1487
rect 1053 1373 1067 1387
rect 1213 1773 1227 1787
rect 1333 1912 1347 1926
rect 1473 2212 1487 2226
rect 1512 2212 1526 2226
rect 1533 2213 1547 2227
rect 1433 2193 1447 2207
rect 1393 2153 1407 2167
rect 1393 2073 1407 2087
rect 1413 2053 1427 2067
rect 1393 1953 1407 1967
rect 1453 2033 1467 2047
rect 1533 2133 1547 2147
rect 1713 2933 1727 2947
rect 1733 2913 1747 2927
rect 1813 2933 1827 2947
rect 1893 3252 1907 3266
rect 1853 3133 1867 3147
rect 1853 3093 1867 3107
rect 1913 3093 1927 3107
rect 1893 3033 1907 3047
rect 1953 3113 1967 3127
rect 1933 3033 1947 3047
rect 1933 2993 1947 3007
rect 1833 2893 1847 2907
rect 1913 2952 1927 2966
rect 1993 3252 2007 3266
rect 2013 3233 2027 3247
rect 2053 3233 2067 3247
rect 2073 3253 2087 3267
rect 2073 3213 2087 3227
rect 2053 3193 2067 3207
rect 2013 3153 2027 3167
rect 1993 3033 2007 3047
rect 1953 2933 1967 2947
rect 1873 2873 1887 2887
rect 1793 2793 1807 2807
rect 1773 2774 1787 2788
rect 1833 2774 1847 2788
rect 1693 2733 1707 2747
rect 1753 2732 1767 2746
rect 1793 2732 1807 2746
rect 1673 2713 1687 2727
rect 1732 2713 1746 2727
rect 1653 2693 1667 2707
rect 1633 2633 1647 2647
rect 1693 2593 1707 2607
rect 1653 2573 1667 2587
rect 1593 2533 1607 2547
rect 1613 2474 1627 2488
rect 1713 2493 1727 2507
rect 1693 2474 1707 2488
rect 1633 2413 1647 2427
rect 1693 2433 1707 2447
rect 1593 2373 1607 2387
rect 1673 2373 1687 2387
rect 1713 2413 1727 2427
rect 1853 2753 1867 2767
rect 1833 2693 1847 2707
rect 1873 2713 1887 2727
rect 1853 2653 1867 2667
rect 1813 2593 1827 2607
rect 1853 2593 1867 2607
rect 1793 2573 1807 2587
rect 1813 2553 1827 2567
rect 1753 2533 1767 2547
rect 1833 2533 1847 2547
rect 1813 2513 1827 2527
rect 1773 2493 1787 2507
rect 1753 2473 1767 2487
rect 1813 2474 1827 2488
rect 1753 2432 1767 2446
rect 1733 2393 1747 2407
rect 1733 2372 1747 2386
rect 1653 2333 1667 2347
rect 1693 2333 1707 2347
rect 1693 2312 1707 2326
rect 1653 2293 1667 2307
rect 1633 2273 1647 2287
rect 1833 2432 1847 2446
rect 1793 2413 1807 2427
rect 1893 2693 1907 2707
rect 1893 2653 1907 2667
rect 1913 2593 1927 2607
rect 2033 3033 2047 3047
rect 2013 2993 2027 3007
rect 2133 3233 2147 3247
rect 2113 3193 2127 3207
rect 2073 3053 2087 3067
rect 2173 3253 2187 3267
rect 2193 3233 2207 3247
rect 2173 3173 2187 3187
rect 2153 3153 2167 3167
rect 2333 3693 2347 3707
rect 2313 3373 2327 3387
rect 2253 3353 2267 3367
rect 2733 4253 2747 4267
rect 2653 4213 2667 4227
rect 2693 4213 2707 4227
rect 2533 4173 2547 4187
rect 2573 4153 2587 4167
rect 2633 4113 2647 4127
rect 2613 4053 2627 4067
rect 2713 4153 2727 4167
rect 2693 4093 2707 4107
rect 2673 4072 2687 4086
rect 2653 4053 2667 4067
rect 2633 4033 2647 4047
rect 2573 3992 2587 4006
rect 2533 3893 2547 3907
rect 2613 3893 2627 3907
rect 2653 3893 2667 3907
rect 2553 3853 2567 3867
rect 2473 3833 2487 3847
rect 2513 3833 2527 3847
rect 2453 3813 2467 3827
rect 2613 3852 2627 3866
rect 2593 3814 2607 3828
rect 2633 3813 2647 3827
rect 2393 3733 2407 3747
rect 2413 3673 2427 3687
rect 2352 3633 2366 3647
rect 2373 3633 2387 3647
rect 2373 3573 2387 3587
rect 2353 3513 2367 3527
rect 2493 3773 2507 3787
rect 2453 3753 2467 3767
rect 2433 3653 2447 3667
rect 2433 3593 2447 3607
rect 2413 3513 2427 3527
rect 2393 3472 2407 3486
rect 2273 3333 2287 3347
rect 2333 3333 2347 3347
rect 2233 3253 2247 3267
rect 2233 3193 2247 3207
rect 2273 3193 2287 3207
rect 2313 3193 2327 3207
rect 2253 3153 2267 3167
rect 2213 3113 2227 3127
rect 2133 3093 2147 3107
rect 2113 2993 2127 3007
rect 2072 2952 2086 2966
rect 2093 2953 2107 2967
rect 2033 2933 2047 2947
rect 2013 2873 2027 2887
rect 1973 2773 1987 2787
rect 2053 2853 2067 2867
rect 2053 2813 2067 2827
rect 1993 2732 2007 2746
rect 2013 2713 2027 2727
rect 2013 2673 2027 2687
rect 1953 2493 1967 2507
rect 1892 2473 1906 2487
rect 1913 2474 1927 2488
rect 1993 2453 2007 2467
rect 1893 2433 1907 2447
rect 1873 2393 1887 2407
rect 1853 2373 1867 2387
rect 1813 2313 1827 2327
rect 1753 2293 1767 2307
rect 1793 2293 1807 2307
rect 1713 2254 1727 2268
rect 1773 2254 1787 2268
rect 1873 2333 1887 2347
rect 1852 2273 1866 2287
rect 1913 2413 1927 2427
rect 1973 2433 1987 2447
rect 1933 2393 1947 2407
rect 1953 2373 1967 2387
rect 1913 2333 1927 2347
rect 1933 2273 1947 2287
rect 1593 2153 1607 2167
rect 1653 2212 1667 2226
rect 1893 2253 1907 2267
rect 1973 2353 1987 2367
rect 2033 2613 2047 2627
rect 2093 2833 2107 2847
rect 2133 2953 2147 2967
rect 2193 3073 2207 3087
rect 2173 3033 2187 3047
rect 2313 3172 2327 3186
rect 2313 3093 2327 3107
rect 2372 3373 2386 3387
rect 2393 3373 2407 3387
rect 2433 3373 2447 3387
rect 2473 3613 2487 3627
rect 2553 3753 2567 3767
rect 2533 3693 2547 3707
rect 2493 3593 2507 3607
rect 2573 3733 2587 3747
rect 2653 3753 2667 3767
rect 2633 3633 2647 3647
rect 2573 3533 2587 3547
rect 2553 3513 2567 3527
rect 2753 4034 2767 4048
rect 2813 4293 2827 4307
rect 2793 4273 2807 4287
rect 2693 3992 2707 4006
rect 2733 3992 2747 4006
rect 2773 3973 2787 3987
rect 2753 3873 2767 3887
rect 2693 3853 2707 3867
rect 2713 3833 2727 3847
rect 2693 3813 2707 3827
rect 2873 4173 2887 4187
rect 2833 4093 2847 4107
rect 2853 4073 2867 4087
rect 2813 4053 2827 4067
rect 2853 4034 2867 4048
rect 2893 4153 2907 4167
rect 2793 3853 2807 3867
rect 2793 3832 2807 3846
rect 2833 3992 2847 4006
rect 2873 3993 2887 4007
rect 2873 3953 2887 3967
rect 3053 4413 3067 4427
rect 2933 4333 2947 4347
rect 2973 4293 2987 4307
rect 3013 4253 3027 4267
rect 2953 4193 2967 4207
rect 3013 4153 3027 4167
rect 2933 4033 2947 4047
rect 2913 3993 2927 4007
rect 2933 3893 2947 3907
rect 2913 3873 2927 3887
rect 2893 3833 2907 3847
rect 2853 3814 2867 3828
rect 2693 3773 2707 3787
rect 2653 3593 2667 3607
rect 2573 3493 2587 3507
rect 2473 3473 2487 3487
rect 2453 3353 2467 3367
rect 2373 3292 2387 3306
rect 2433 3294 2447 3308
rect 2513 3453 2527 3467
rect 2593 3473 2607 3487
rect 2573 3433 2587 3447
rect 2513 3393 2527 3407
rect 2493 3333 2507 3347
rect 2473 3293 2487 3307
rect 2353 3173 2367 3187
rect 2393 3213 2407 3227
rect 2433 3213 2447 3227
rect 2373 3133 2387 3147
rect 2413 3093 2427 3107
rect 2273 3053 2287 3067
rect 2293 3033 2307 3047
rect 2233 2994 2247 3008
rect 2393 3053 2407 3067
rect 2313 3013 2327 3027
rect 2333 2994 2347 3008
rect 2193 2933 2207 2947
rect 2173 2913 2187 2927
rect 2153 2873 2167 2887
rect 2173 2853 2187 2867
rect 2133 2813 2147 2827
rect 2273 2953 2287 2967
rect 2233 2913 2247 2927
rect 2233 2873 2247 2887
rect 2213 2833 2227 2847
rect 2173 2793 2187 2807
rect 2093 2773 2107 2787
rect 2133 2774 2147 2788
rect 2073 2593 2087 2607
rect 2013 2433 2027 2447
rect 2013 2353 2027 2367
rect 2013 2293 2027 2307
rect 2013 2272 2027 2286
rect 1953 2253 1967 2267
rect 1753 2193 1767 2207
rect 1793 2193 1807 2207
rect 1653 2173 1667 2187
rect 1713 2173 1727 2187
rect 1613 2133 1627 2147
rect 1613 2112 1627 2126
rect 1593 2073 1607 2087
rect 1533 2053 1547 2067
rect 1573 2053 1587 2067
rect 1473 1993 1487 2007
rect 1733 2153 1747 2167
rect 1673 2133 1687 2147
rect 1653 2053 1667 2067
rect 1592 2033 1606 2047
rect 1613 2033 1627 2047
rect 1493 1953 1507 1967
rect 1533 1954 1547 1968
rect 1713 2093 1727 2107
rect 1613 1954 1627 1968
rect 1713 1993 1727 2007
rect 1693 1954 1707 1968
rect 1313 1873 1327 1887
rect 1373 1873 1387 1887
rect 1293 1733 1307 1747
rect 1193 1693 1207 1707
rect 1173 1513 1187 1527
rect 1093 1473 1107 1487
rect 1153 1473 1167 1487
rect 1093 1433 1107 1447
rect 1233 1692 1247 1706
rect 1273 1653 1287 1667
rect 1393 1793 1407 1807
rect 1333 1753 1347 1767
rect 1533 1873 1547 1887
rect 1453 1773 1467 1787
rect 1493 1773 1507 1787
rect 1433 1753 1447 1767
rect 1333 1713 1347 1727
rect 1433 1713 1447 1727
rect 1373 1653 1387 1667
rect 1413 1593 1427 1607
rect 1313 1533 1327 1547
rect 1233 1473 1247 1487
rect 1333 1473 1347 1487
rect 1373 1473 1387 1487
rect 1193 1434 1207 1448
rect 1273 1434 1287 1448
rect 1093 1393 1107 1407
rect 1033 1293 1047 1307
rect 1033 1213 1047 1227
rect 1013 1153 1027 1167
rect 993 993 1007 1007
rect 1073 1313 1087 1327
rect 1153 1373 1167 1387
rect 1253 1373 1267 1387
rect 1113 1333 1127 1347
rect 1253 1313 1267 1327
rect 1093 1273 1107 1287
rect 1133 1273 1147 1287
rect 1193 1273 1207 1287
rect 1093 1214 1107 1228
rect 1073 1173 1087 1187
rect 1053 1153 1067 1167
rect 1053 993 1067 1007
rect 1033 933 1047 947
rect 1013 914 1027 928
rect 1333 1373 1347 1387
rect 1353 1293 1367 1307
rect 1293 1253 1307 1267
rect 1333 1253 1347 1267
rect 1293 1214 1307 1228
rect 1153 1153 1167 1167
rect 1313 1173 1327 1187
rect 1273 1113 1287 1127
rect 1113 1073 1127 1087
rect 1273 1073 1287 1087
rect 1193 993 1207 1007
rect 1073 973 1087 987
rect 1233 973 1247 987
rect 1093 933 1107 947
rect 1153 933 1167 947
rect 953 853 967 867
rect 933 773 947 787
rect 832 733 846 747
rect 853 733 867 747
rect 813 693 827 707
rect 733 652 747 666
rect 673 633 687 647
rect 773 613 787 627
rect 833 573 847 587
rect 793 473 807 487
rect 693 394 707 408
rect 733 394 747 408
rect 1033 853 1047 867
rect 1293 953 1307 967
rect 1493 1734 1507 1748
rect 1553 1813 1567 1827
rect 1593 1813 1607 1827
rect 1573 1793 1587 1807
rect 1573 1733 1587 1747
rect 1553 1692 1567 1706
rect 1513 1633 1527 1647
rect 1633 1913 1647 1927
rect 1613 1752 1627 1766
rect 1653 1813 1667 1827
rect 1633 1733 1647 1747
rect 1852 2213 1866 2227
rect 1873 2213 1887 2227
rect 1833 2093 1847 2107
rect 1853 1953 1867 1967
rect 1693 1873 1707 1887
rect 1753 1893 1767 1907
rect 1713 1853 1727 1867
rect 1693 1813 1707 1827
rect 1673 1793 1687 1807
rect 1693 1753 1707 1767
rect 1772 1853 1786 1867
rect 1793 1853 1807 1867
rect 1753 1712 1767 1726
rect 1613 1653 1627 1667
rect 1593 1573 1607 1587
rect 1493 1533 1507 1547
rect 1433 1473 1447 1487
rect 1473 1473 1487 1487
rect 1673 1692 1687 1706
rect 1713 1673 1727 1687
rect 1553 1513 1567 1527
rect 1612 1513 1626 1527
rect 1633 1513 1647 1527
rect 1513 1493 1527 1507
rect 1493 1453 1507 1467
rect 1593 1493 1607 1507
rect 1433 1392 1447 1406
rect 1513 1392 1527 1406
rect 1453 1373 1467 1387
rect 1613 1392 1627 1406
rect 1553 1373 1567 1387
rect 1573 1373 1587 1387
rect 1553 1293 1567 1307
rect 1513 1253 1527 1267
rect 1433 1214 1447 1228
rect 1613 1233 1627 1247
rect 1613 1193 1627 1207
rect 1373 1172 1387 1186
rect 1413 1172 1427 1186
rect 1353 1153 1367 1167
rect 1473 1173 1487 1187
rect 1453 1153 1467 1167
rect 1473 1113 1487 1127
rect 1413 1093 1427 1107
rect 1513 1093 1527 1107
rect 1333 1033 1347 1047
rect 1613 1073 1627 1087
rect 1373 973 1387 987
rect 1333 953 1347 967
rect 1333 914 1347 928
rect 1373 914 1387 928
rect 1133 872 1147 886
rect 1093 793 1107 807
rect 1153 793 1167 807
rect 1093 733 1107 747
rect 893 694 907 708
rect 933 694 947 708
rect 993 694 1007 708
rect 1053 694 1067 708
rect 873 653 887 667
rect 913 652 927 666
rect 1133 693 1147 707
rect 913 593 927 607
rect 953 573 967 587
rect 1073 573 1087 587
rect 873 533 887 547
rect 853 453 867 467
rect 1233 872 1247 886
rect 1313 872 1327 886
rect 1173 733 1187 747
rect 1233 733 1247 747
rect 1293 733 1307 747
rect 1273 713 1287 727
rect 1193 694 1207 708
rect 1233 694 1247 708
rect 1573 973 1587 987
rect 1573 933 1587 947
rect 1533 914 1547 928
rect 1633 1013 1647 1027
rect 1633 953 1647 967
rect 1813 1813 1827 1827
rect 1833 1753 1847 1767
rect 1913 2212 1927 2226
rect 1953 2213 1967 2227
rect 1993 2213 2007 2227
rect 1893 2173 1907 2187
rect 1973 2132 1987 2146
rect 1893 2113 1907 2127
rect 2113 2733 2127 2747
rect 2153 2713 2167 2727
rect 2153 2653 2167 2667
rect 2133 2573 2147 2587
rect 2133 2533 2147 2547
rect 2093 2493 2107 2507
rect 2133 2493 2147 2507
rect 2153 2473 2167 2487
rect 2093 2432 2107 2446
rect 2053 2393 2067 2407
rect 2092 2353 2106 2367
rect 2113 2353 2127 2367
rect 2113 2313 2127 2327
rect 2213 2613 2227 2627
rect 2193 2493 2207 2507
rect 2253 2833 2267 2847
rect 2373 2953 2387 2967
rect 2353 2933 2367 2947
rect 2393 2933 2407 2947
rect 2333 2853 2347 2867
rect 2313 2833 2327 2847
rect 2293 2813 2307 2827
rect 2273 2793 2287 2807
rect 2473 3253 2487 3267
rect 2453 3133 2467 3147
rect 2553 3373 2567 3387
rect 2533 3353 2547 3367
rect 2513 3173 2527 3187
rect 2473 3093 2487 3107
rect 2473 3033 2487 3047
rect 2633 3413 2647 3427
rect 2553 3332 2567 3346
rect 2593 3333 2607 3347
rect 2553 3293 2567 3307
rect 2593 3294 2607 3308
rect 2573 3252 2587 3266
rect 2573 3231 2587 3245
rect 2613 3233 2627 3247
rect 2593 3153 2607 3167
rect 2573 3113 2587 3127
rect 2513 2952 2527 2966
rect 2453 2933 2467 2947
rect 2433 2913 2447 2927
rect 2413 2893 2427 2907
rect 2393 2853 2407 2867
rect 2353 2773 2367 2787
rect 2473 2913 2487 2927
rect 2413 2774 2427 2788
rect 2253 2693 2267 2707
rect 2333 2733 2347 2747
rect 2273 2633 2287 2647
rect 2233 2553 2247 2567
rect 2213 2473 2227 2487
rect 2313 2593 2327 2607
rect 2293 2533 2307 2547
rect 2253 2473 2267 2487
rect 2253 2433 2267 2447
rect 2213 2413 2227 2427
rect 2193 2293 2207 2307
rect 2093 2254 2107 2268
rect 2152 2253 2166 2267
rect 2033 2153 2047 2167
rect 1992 2093 2006 2107
rect 2013 2093 2027 2107
rect 1973 2073 1987 2087
rect 1933 1954 1947 1968
rect 1893 1933 1907 1947
rect 1953 1912 1967 1926
rect 1973 1873 1987 1887
rect 1933 1813 1947 1827
rect 1953 1753 1967 1767
rect 1813 1673 1827 1687
rect 1753 1633 1767 1647
rect 1733 1613 1747 1627
rect 1772 1573 1786 1587
rect 1793 1573 1807 1587
rect 1713 1434 1727 1448
rect 1673 1393 1687 1407
rect 1733 1392 1747 1406
rect 1853 1553 1867 1567
rect 1793 1513 1807 1527
rect 1853 1513 1867 1527
rect 1933 1692 1947 1706
rect 1913 1633 1927 1647
rect 1993 1813 2007 1827
rect 2033 2073 2047 2087
rect 2033 2033 2047 2047
rect 2073 2212 2087 2226
rect 2092 2073 2106 2087
rect 2113 2073 2127 2087
rect 2093 2033 2107 2047
rect 2073 2013 2087 2027
rect 2073 1973 2087 1987
rect 2113 1973 2127 1987
rect 2173 2252 2187 2266
rect 2433 2732 2447 2746
rect 2413 2713 2427 2727
rect 2373 2633 2387 2647
rect 2433 2693 2447 2707
rect 2493 2893 2507 2907
rect 2413 2593 2427 2607
rect 2413 2572 2427 2586
rect 2353 2493 2367 2507
rect 2333 2473 2347 2487
rect 2453 2673 2467 2687
rect 2433 2553 2447 2567
rect 2433 2473 2447 2487
rect 2333 2433 2347 2447
rect 2393 2432 2407 2446
rect 2433 2432 2447 2446
rect 2333 2393 2347 2407
rect 2313 2373 2327 2387
rect 2353 2333 2367 2347
rect 2253 2273 2267 2287
rect 2293 2273 2307 2287
rect 2412 2293 2426 2307
rect 2433 2293 2447 2307
rect 2373 2273 2387 2287
rect 2192 2193 2206 2207
rect 2213 2193 2227 2207
rect 2153 2073 2167 2087
rect 2153 2033 2167 2047
rect 2153 1992 2167 2006
rect 2093 1954 2107 1968
rect 2133 1954 2147 1968
rect 2053 1893 2067 1907
rect 2033 1873 2047 1887
rect 2093 1853 2107 1867
rect 2013 1754 2027 1768
rect 2273 2173 2287 2187
rect 2233 2153 2247 2167
rect 2213 2113 2227 2127
rect 2233 2053 2247 2067
rect 2213 2033 2227 2047
rect 2233 1993 2247 2007
rect 2353 2193 2367 2207
rect 2333 2173 2347 2187
rect 2293 2153 2307 2167
rect 2353 2153 2367 2167
rect 2333 2013 2347 2027
rect 2293 1993 2307 2007
rect 2233 1954 2247 1968
rect 2313 1933 2327 1947
rect 2233 1893 2247 1907
rect 2213 1853 2227 1867
rect 2113 1833 2127 1847
rect 2193 1833 2207 1847
rect 2113 1773 2127 1787
rect 2173 1773 2187 1787
rect 2013 1733 2027 1747
rect 2053 1734 2067 1748
rect 2093 1734 2107 1748
rect 1993 1692 2007 1706
rect 2073 1673 2087 1687
rect 2133 1734 2147 1748
rect 2213 1733 2227 1747
rect 2113 1693 2127 1707
rect 1953 1593 1967 1607
rect 2093 1593 2107 1607
rect 1913 1533 1927 1547
rect 1933 1513 1947 1527
rect 2153 1692 2167 1706
rect 2193 1692 2207 1706
rect 2153 1613 2167 1627
rect 2153 1533 2167 1547
rect 2132 1513 2146 1527
rect 1852 1453 1866 1467
rect 1793 1433 1807 1447
rect 1873 1452 1887 1466
rect 1893 1453 1907 1467
rect 1913 1434 1927 1448
rect 1813 1392 1827 1406
rect 2053 1493 2067 1507
rect 2013 1434 2027 1448
rect 2153 1512 2167 1526
rect 2153 1453 2167 1467
rect 2173 1434 2187 1448
rect 2333 1853 2347 1867
rect 2313 1773 2327 1787
rect 2293 1734 2307 1748
rect 2233 1633 2247 1647
rect 2313 1692 2327 1706
rect 2273 1653 2287 1667
rect 2293 1633 2307 1647
rect 2313 1593 2327 1607
rect 2293 1553 2307 1567
rect 2213 1493 2227 1507
rect 2253 1493 2267 1507
rect 2273 1434 2287 1448
rect 1933 1393 1947 1407
rect 1853 1373 1867 1387
rect 1913 1373 1927 1387
rect 1813 1353 1827 1367
rect 2033 1392 2047 1406
rect 2093 1392 2107 1406
rect 1993 1353 2007 1367
rect 1813 1313 1827 1327
rect 1973 1313 1987 1327
rect 1773 1293 1787 1307
rect 1853 1253 1867 1267
rect 1693 1233 1707 1247
rect 1733 1214 1747 1228
rect 1793 1213 1807 1227
rect 1853 1214 1867 1228
rect 1913 1213 1927 1227
rect 2053 1233 2067 1247
rect 2013 1213 2027 1227
rect 2213 1393 2227 1407
rect 2113 1353 2127 1367
rect 2153 1353 2167 1367
rect 2113 1313 2127 1327
rect 2153 1293 2167 1307
rect 2153 1253 2167 1267
rect 2113 1233 2127 1247
rect 1693 1013 1707 1027
rect 1653 933 1667 947
rect 1633 914 1647 928
rect 1713 993 1727 1007
rect 1793 1172 1807 1186
rect 1833 1172 1847 1186
rect 1753 953 1767 967
rect 1713 914 1727 928
rect 1753 914 1767 928
rect 1853 1093 1867 1107
rect 1393 833 1407 847
rect 1353 694 1367 708
rect 1393 694 1407 708
rect 1513 872 1527 886
rect 1573 872 1587 886
rect 1653 872 1667 886
rect 1693 872 1707 886
rect 1733 872 1747 886
rect 1733 813 1747 827
rect 1513 793 1527 807
rect 1473 693 1487 707
rect 1653 773 1667 787
rect 1553 694 1567 708
rect 1653 694 1667 708
rect 1253 652 1267 666
rect 1293 652 1307 666
rect 1373 652 1387 666
rect 1413 653 1427 667
rect 1213 633 1227 647
rect 1153 613 1167 627
rect 1213 533 1227 547
rect 993 513 1007 527
rect 1093 513 1107 527
rect 1133 513 1147 527
rect 953 493 967 507
rect 893 453 907 467
rect 933 453 947 467
rect 673 353 687 367
rect 653 333 667 347
rect 713 333 727 347
rect 673 313 687 327
rect 613 293 627 307
rect 653 273 667 287
rect 593 213 607 227
rect 733 253 747 267
rect 793 353 807 367
rect 833 352 847 366
rect 1033 493 1047 507
rect 813 313 827 327
rect 753 213 767 227
rect 953 353 967 367
rect 1013 352 1027 366
rect 933 313 947 327
rect 913 273 927 287
rect 833 253 847 267
rect 893 253 907 267
rect 593 132 607 146
rect 633 132 647 146
rect 513 113 527 127
rect 559 113 573 127
rect 733 73 747 87
rect 313 53 327 67
rect 813 193 827 207
rect 793 174 807 188
rect 873 213 887 227
rect 873 173 887 187
rect 813 132 827 146
rect 853 132 867 146
rect 913 153 927 167
rect 993 253 1007 267
rect 1053 253 1067 267
rect 1173 493 1187 507
rect 1173 453 1187 467
rect 1113 393 1127 407
rect 1373 493 1387 507
rect 1273 453 1287 467
rect 1213 393 1227 407
rect 1313 394 1327 408
rect 1113 353 1127 367
rect 1153 352 1167 366
rect 1193 352 1207 366
rect 1253 352 1267 366
rect 1113 313 1127 327
rect 1273 313 1287 327
rect 1233 273 1247 287
rect 1093 233 1107 247
rect 1173 233 1187 247
rect 993 174 1007 188
rect 1113 174 1127 188
rect 1153 173 1167 187
rect 933 133 947 147
rect 973 132 987 146
rect 1053 132 1067 146
rect 1833 872 1847 886
rect 1773 773 1787 787
rect 1813 773 1827 787
rect 1813 733 1827 747
rect 1913 1073 1927 1087
rect 1913 1033 1927 1047
rect 1893 973 1907 987
rect 1933 933 1947 947
rect 2033 1173 2047 1187
rect 2253 1392 2267 1406
rect 2213 1372 2227 1386
rect 2333 1553 2347 1567
rect 2373 2093 2387 2107
rect 2533 2873 2547 2887
rect 2513 2813 2527 2827
rect 2633 3113 2647 3127
rect 2633 3053 2647 3067
rect 2673 3333 2687 3347
rect 2793 3773 2807 3787
rect 2973 3992 2987 4006
rect 3213 4773 3227 4787
rect 3293 4973 3307 4987
rect 3293 4933 3307 4947
rect 3313 4893 3327 4907
rect 3313 4854 3327 4868
rect 3293 4812 3307 4826
rect 3293 4753 3307 4767
rect 3273 4693 3287 4707
rect 3273 4653 3287 4667
rect 3253 4633 3267 4647
rect 3233 4553 3247 4567
rect 3173 4493 3187 4507
rect 3413 5332 3427 5346
rect 3433 5313 3447 5327
rect 3393 5193 3407 5207
rect 3493 5332 3507 5346
rect 3573 5332 3587 5346
rect 3613 5332 3627 5346
rect 3453 5253 3467 5267
rect 3613 5293 3627 5307
rect 3493 5233 3507 5247
rect 3513 5193 3527 5207
rect 3433 5153 3447 5167
rect 3393 5073 3407 5087
rect 3473 5074 3487 5088
rect 3533 5173 3547 5187
rect 3633 5173 3647 5187
rect 3553 5133 3567 5147
rect 3593 5133 3607 5147
rect 3553 5093 3567 5107
rect 3593 5074 3607 5088
rect 3673 5493 3687 5507
rect 3393 4953 3407 4967
rect 3493 5032 3507 5046
rect 3533 5033 3547 5047
rect 3493 4993 3507 5007
rect 3473 4973 3487 4987
rect 3473 4933 3487 4947
rect 3393 4913 3407 4927
rect 3453 4913 3467 4927
rect 3433 4893 3447 4907
rect 3613 5032 3627 5046
rect 3633 5013 3647 5027
rect 3553 4973 3567 4987
rect 3593 4973 3607 4987
rect 3553 4854 3567 4868
rect 3613 4853 3627 4867
rect 3413 4773 3427 4787
rect 3453 4773 3467 4787
rect 3353 4753 3367 4767
rect 3333 4713 3347 4727
rect 3313 4553 3327 4567
rect 3493 4593 3507 4607
rect 3533 4812 3547 4826
rect 3573 4733 3587 4747
rect 3553 4673 3567 4687
rect 3552 4633 3566 4647
rect 3573 4633 3587 4647
rect 3613 4773 3627 4787
rect 3613 4693 3627 4707
rect 3613 4553 3627 4567
rect 3313 4473 3327 4487
rect 3213 4413 3227 4427
rect 3293 4413 3307 4427
rect 3293 4373 3307 4387
rect 3273 4253 3287 4267
rect 3193 4233 3207 4247
rect 3253 4193 3267 4207
rect 3253 4113 3267 4127
rect 3173 4036 3187 4050
rect 3233 4036 3247 4050
rect 3113 3893 3127 3907
rect 3413 4393 3427 4407
rect 3333 4373 3347 4387
rect 3453 4373 3467 4387
rect 3373 4334 3387 4348
rect 3413 4334 3427 4348
rect 3313 4093 3327 4107
rect 3293 4073 3307 4087
rect 3333 4073 3347 4087
rect 3353 4053 3367 4067
rect 3373 4034 3387 4048
rect 3553 4473 3567 4487
rect 3613 4473 3627 4487
rect 3573 4433 3587 4447
rect 3533 4373 3547 4387
rect 3493 4334 3507 4348
rect 3593 4393 3607 4407
rect 3573 4333 3587 4347
rect 3453 4233 3467 4247
rect 3553 4292 3567 4306
rect 3573 4273 3587 4287
rect 3573 4193 3587 4207
rect 3793 5793 3807 5807
rect 3853 5773 3867 5787
rect 3793 5753 3807 5767
rect 3853 5713 3867 5727
rect 3793 5594 3807 5608
rect 3833 5593 3847 5607
rect 3773 5473 3787 5487
rect 3733 5453 3747 5467
rect 3713 5374 3727 5388
rect 3753 5374 3767 5388
rect 4373 6233 4387 6247
rect 4433 6233 4447 6247
rect 4353 6213 4367 6227
rect 3893 6153 3907 6167
rect 4013 6153 4027 6167
rect 4293 6153 4307 6167
rect 3892 6114 3906 6128
rect 3913 6114 3927 6128
rect 3953 6114 3967 6128
rect 3993 6114 4007 6128
rect 4033 6114 4047 6128
rect 4093 6114 4107 6128
rect 3893 6073 3907 6087
rect 3933 6072 3947 6086
rect 3973 6053 3987 6067
rect 4013 6053 4027 6067
rect 3973 5933 3987 5947
rect 3913 5852 3927 5866
rect 4132 6113 4146 6127
rect 4153 6114 4167 6128
rect 4193 6114 4207 6128
rect 4233 6114 4247 6128
rect 4133 6053 4147 6067
rect 4253 6072 4267 6086
rect 4373 6193 4387 6207
rect 4393 6153 4407 6167
rect 4353 6114 4367 6128
rect 4233 6053 4247 6067
rect 4213 6033 4227 6047
rect 4153 6013 4167 6027
rect 4293 6053 4307 6067
rect 4273 6033 4287 6047
rect 4193 5993 4207 6007
rect 4233 5993 4247 6007
rect 4193 5953 4207 5967
rect 4033 5933 4047 5947
rect 4133 5933 4147 5947
rect 4333 6013 4347 6027
rect 4332 5992 4346 6006
rect 4353 5993 4367 6007
rect 4253 5913 4267 5927
rect 4293 5913 4307 5927
rect 4093 5894 4107 5908
rect 4133 5894 4147 5908
rect 4213 5894 4227 5908
rect 4073 5852 4087 5866
rect 3953 5833 3967 5847
rect 4013 5833 4027 5847
rect 3933 5753 3947 5767
rect 3893 5733 3907 5747
rect 3873 5593 3887 5607
rect 4073 5813 4087 5827
rect 4172 5853 4186 5867
rect 4193 5852 4207 5866
rect 4273 5853 4287 5867
rect 4393 6033 4407 6047
rect 4373 5913 4387 5927
rect 4933 6213 4947 6227
rect 4793 6153 4807 6167
rect 4493 6114 4507 6128
rect 4553 6113 4567 6127
rect 4833 6114 4847 6128
rect 4893 6114 4907 6128
rect 4453 6072 4467 6086
rect 4513 6072 4527 6086
rect 4553 6072 4567 6086
rect 4433 5993 4447 6007
rect 4492 6033 4506 6047
rect 4513 6033 4527 6047
rect 4473 5973 4487 5987
rect 4453 5953 4467 5967
rect 4433 5913 4447 5927
rect 4493 5933 4507 5947
rect 4533 5933 4547 5947
rect 4573 6033 4587 6047
rect 4633 5973 4647 5987
rect 4613 5933 4627 5947
rect 4613 5893 4627 5907
rect 4333 5852 4347 5866
rect 4373 5852 4387 5866
rect 4473 5852 4487 5866
rect 4513 5852 4527 5866
rect 4113 5793 4127 5807
rect 4273 5793 4287 5807
rect 4373 5793 4387 5807
rect 4053 5773 4067 5787
rect 4033 5753 4047 5767
rect 3953 5693 3967 5707
rect 3993 5693 4007 5707
rect 3933 5673 3947 5687
rect 3933 5594 3947 5608
rect 3852 5553 3866 5567
rect 3873 5553 3887 5567
rect 3853 5513 3867 5527
rect 3812 5373 3826 5387
rect 3833 5373 3847 5387
rect 3873 5493 3887 5507
rect 3953 5553 3967 5567
rect 4013 5653 4027 5667
rect 4033 5633 4047 5647
rect 4013 5593 4027 5607
rect 4233 5713 4247 5727
rect 4093 5594 4107 5608
rect 4133 5594 4147 5608
rect 4193 5594 4207 5608
rect 4373 5633 4387 5647
rect 4273 5594 4287 5608
rect 4313 5594 4327 5608
rect 4353 5594 4367 5608
rect 4013 5553 4027 5567
rect 3993 5513 4007 5527
rect 3913 5473 3927 5487
rect 3893 5453 3907 5467
rect 3933 5433 3947 5447
rect 3973 5433 3987 5447
rect 4033 5513 4047 5527
rect 4073 5513 4087 5527
rect 4173 5533 4187 5547
rect 4253 5533 4267 5547
rect 4153 5473 4167 5487
rect 4213 5473 4227 5487
rect 4073 5433 4087 5447
rect 3933 5373 3947 5387
rect 3733 5253 3747 5267
rect 3713 5233 3727 5247
rect 3912 5332 3926 5346
rect 3933 5332 3947 5346
rect 3813 5293 3827 5307
rect 3773 5213 3787 5227
rect 3713 5153 3727 5167
rect 3813 5153 3827 5167
rect 3693 5113 3707 5127
rect 3773 5113 3787 5127
rect 3673 5013 3687 5027
rect 3653 4973 3667 4987
rect 3733 5074 3747 5088
rect 3833 5113 3847 5127
rect 3713 5033 3727 5047
rect 3713 4993 3727 5007
rect 3753 4973 3767 4987
rect 3693 4873 3707 4887
rect 3653 4853 3667 4867
rect 3713 4854 3727 4868
rect 3913 5253 3927 5267
rect 3873 5233 3887 5247
rect 3933 5233 3947 5247
rect 4013 5332 4027 5346
rect 4093 5413 4107 5427
rect 3993 5293 4007 5307
rect 4073 5293 4087 5307
rect 3973 5273 3987 5287
rect 3973 5233 3987 5247
rect 3893 5133 3907 5147
rect 3873 5073 3887 5087
rect 3953 5173 3967 5187
rect 3953 5113 3967 5127
rect 3933 5073 3947 5087
rect 3853 5013 3867 5027
rect 3892 5013 3906 5027
rect 3913 5013 3927 5027
rect 3793 4993 3807 5007
rect 3813 4973 3827 4987
rect 3773 4933 3787 4947
rect 3813 4933 3827 4947
rect 3793 4913 3807 4927
rect 3753 4853 3767 4867
rect 3833 4854 3847 4868
rect 3653 4773 3667 4787
rect 3733 4812 3747 4826
rect 3813 4812 3827 4826
rect 3793 4793 3807 4807
rect 3773 4713 3787 4727
rect 3693 4693 3707 4707
rect 3653 4673 3667 4687
rect 3633 4353 3647 4367
rect 3693 4672 3707 4686
rect 3733 4554 3747 4568
rect 3773 4513 3787 4527
rect 3713 4433 3727 4447
rect 3713 4393 3727 4407
rect 3613 4253 3627 4267
rect 3693 4334 3707 4348
rect 3733 4336 3747 4350
rect 3653 4293 3667 4307
rect 3713 4293 3727 4307
rect 3672 4253 3686 4267
rect 3693 4253 3707 4267
rect 3653 4193 3667 4207
rect 3633 4173 3647 4187
rect 3593 4133 3607 4147
rect 3653 4133 3667 4147
rect 3513 4113 3527 4127
rect 3493 4093 3507 4107
rect 3293 4013 3307 4027
rect 3153 3993 3167 4007
rect 3033 3853 3047 3867
rect 3073 3853 3087 3867
rect 3133 3853 3147 3867
rect 2993 3833 3007 3847
rect 3053 3833 3067 3847
rect 2953 3813 2967 3827
rect 2833 3772 2847 3786
rect 2853 3753 2867 3767
rect 2793 3693 2807 3707
rect 2733 3633 2747 3647
rect 2933 3772 2947 3786
rect 2973 3772 2987 3786
rect 3013 3772 3027 3786
rect 2893 3753 2907 3767
rect 2993 3693 3007 3707
rect 2893 3673 2907 3687
rect 2913 3653 2927 3667
rect 2873 3613 2887 3627
rect 2853 3573 2867 3587
rect 2753 3533 2767 3547
rect 2853 3513 2867 3527
rect 2873 3533 2887 3547
rect 3033 3673 3047 3687
rect 3013 3573 3027 3587
rect 2953 3514 2967 3528
rect 2993 3514 3007 3528
rect 2833 3493 2847 3507
rect 2813 3433 2827 3447
rect 2773 3413 2787 3427
rect 2733 3373 2747 3387
rect 2713 3353 2727 3367
rect 2693 3313 2707 3327
rect 2773 3353 2787 3367
rect 2753 3313 2767 3327
rect 2733 3293 2747 3307
rect 2673 3253 2687 3267
rect 2733 3253 2747 3267
rect 2713 3213 2727 3227
rect 2693 3193 2707 3207
rect 2673 3113 2687 3127
rect 2653 3013 2667 3027
rect 2693 3033 2707 3047
rect 2613 2933 2627 2947
rect 2553 2813 2567 2827
rect 2693 2953 2707 2967
rect 2893 3472 2907 3486
rect 2973 3453 2987 3467
rect 2933 3393 2947 3407
rect 2893 3373 2907 3387
rect 2833 3353 2847 3367
rect 2813 3313 2827 3327
rect 2873 3313 2887 3327
rect 2833 3294 2847 3308
rect 2813 3252 2827 3266
rect 2853 3252 2867 3266
rect 2993 3433 3007 3447
rect 3013 3373 3027 3387
rect 3053 3633 3067 3647
rect 3093 3813 3107 3827
rect 3353 3992 3367 4006
rect 3393 3993 3407 4007
rect 3513 4033 3527 4047
rect 3553 4036 3567 4050
rect 3613 4036 3627 4050
rect 3293 3953 3307 3967
rect 3433 3990 3447 4004
rect 3493 3990 3507 4004
rect 3413 3953 3427 3967
rect 3293 3913 3307 3927
rect 3393 3913 3407 3927
rect 3193 3893 3207 3907
rect 3213 3873 3227 3887
rect 3193 3853 3207 3867
rect 3213 3813 3227 3827
rect 3173 3772 3187 3786
rect 3093 3753 3107 3767
rect 3213 3753 3227 3767
rect 3173 3733 3187 3747
rect 3193 3693 3207 3707
rect 3173 3633 3187 3647
rect 3172 3593 3186 3607
rect 3193 3593 3207 3607
rect 3493 3933 3507 3947
rect 3633 3993 3647 4007
rect 3633 3953 3647 3967
rect 3433 3913 3447 3927
rect 3513 3913 3527 3927
rect 3413 3893 3427 3907
rect 3313 3833 3327 3847
rect 3453 3893 3467 3907
rect 3613 3893 3627 3907
rect 3433 3813 3447 3827
rect 3313 3773 3327 3787
rect 3352 3770 3366 3784
rect 3373 3773 3387 3787
rect 3473 3873 3487 3887
rect 3313 3733 3327 3747
rect 3413 3770 3427 3784
rect 3453 3770 3467 3784
rect 3493 3833 3507 3847
rect 3513 3814 3527 3828
rect 3493 3773 3507 3787
rect 3473 3753 3487 3767
rect 3353 3673 3367 3687
rect 3273 3653 3287 3667
rect 3313 3653 3327 3667
rect 3253 3633 3267 3647
rect 3233 3593 3247 3607
rect 3073 3553 3087 3567
rect 3153 3553 3167 3567
rect 3213 3553 3227 3567
rect 3113 3514 3127 3528
rect 3153 3513 3167 3527
rect 3193 3514 3207 3528
rect 3253 3513 3267 3527
rect 2913 3333 2927 3347
rect 2973 3333 2987 3347
rect 3073 3333 3087 3347
rect 2773 3233 2787 3247
rect 2893 3233 2907 3247
rect 2873 3213 2887 3227
rect 2853 3193 2867 3207
rect 2773 3153 2787 3167
rect 2813 3153 2827 3167
rect 2753 3093 2767 3107
rect 2833 3113 2847 3127
rect 2833 3073 2847 3087
rect 2733 2993 2747 3007
rect 2773 2994 2787 3008
rect 2813 2993 2827 3007
rect 2713 2913 2727 2927
rect 2653 2853 2667 2867
rect 2733 2833 2747 2847
rect 2733 2793 2747 2807
rect 2613 2773 2627 2787
rect 2693 2774 2707 2788
rect 2513 2713 2527 2727
rect 2493 2673 2507 2687
rect 2533 2693 2547 2707
rect 2553 2673 2567 2687
rect 2633 2753 2647 2767
rect 2673 2732 2687 2746
rect 2713 2732 2727 2746
rect 2833 2953 2847 2967
rect 2793 2913 2807 2927
rect 2793 2892 2807 2906
rect 2893 3173 2907 3187
rect 2873 3113 2887 3127
rect 2973 3294 2987 3308
rect 2953 3252 2967 3266
rect 2933 3213 2947 3227
rect 2933 3153 2947 3167
rect 2913 3053 2927 3067
rect 2893 3033 2907 3047
rect 3013 3213 3027 3227
rect 2993 3073 3007 3087
rect 2973 3013 2987 3027
rect 2993 2993 3007 3007
rect 2873 2953 2887 2967
rect 2853 2893 2867 2907
rect 2913 2952 2927 2966
rect 3152 3473 3166 3487
rect 3173 3473 3187 3487
rect 3153 3433 3167 3447
rect 3133 3413 3147 3427
rect 3113 3393 3127 3407
rect 3093 3313 3107 3327
rect 3133 3333 3147 3347
rect 3133 3252 3147 3266
rect 3093 3213 3107 3227
rect 3033 3193 3047 3207
rect 3133 3173 3147 3187
rect 3033 3133 3047 3147
rect 3073 3133 3087 3147
rect 3053 3113 3067 3127
rect 3033 3053 3047 3067
rect 3193 3453 3207 3467
rect 3253 3473 3267 3487
rect 3213 3433 3227 3447
rect 3573 3733 3587 3747
rect 3673 4113 3687 4127
rect 3773 4193 3787 4207
rect 3713 4153 3727 4167
rect 3693 4033 3707 4047
rect 3873 4813 3887 4827
rect 3853 4773 3867 4787
rect 3813 4613 3827 4627
rect 3873 4593 3887 4607
rect 3933 4913 3947 4927
rect 3913 4893 3927 4907
rect 4033 5213 4047 5227
rect 4033 5173 4047 5187
rect 4013 5153 4027 5167
rect 4013 5113 4027 5127
rect 4052 5113 4066 5127
rect 4073 5113 4087 5127
rect 4193 5374 4207 5388
rect 4333 5552 4347 5566
rect 4373 5513 4387 5527
rect 4413 5813 4427 5827
rect 4593 5852 4607 5866
rect 4633 5852 4647 5866
rect 4593 5693 4607 5707
rect 4413 5673 4427 5687
rect 4553 5673 4567 5687
rect 4393 5433 4407 5447
rect 4513 5633 4527 5647
rect 4433 5594 4447 5608
rect 4473 5594 4487 5608
rect 4633 5594 4647 5608
rect 4673 6033 4687 6047
rect 4813 6072 4827 6086
rect 5193 6253 5207 6267
rect 5073 6233 5087 6247
rect 5113 6233 5127 6247
rect 4953 6193 4967 6207
rect 4973 6153 4987 6167
rect 5013 6133 5027 6147
rect 4933 6033 4947 6047
rect 4793 5993 4807 6007
rect 4853 5993 4867 6007
rect 4893 5993 4907 6007
rect 4733 5973 4747 5987
rect 4713 5953 4727 5967
rect 4673 5893 4687 5907
rect 4773 5953 4787 5967
rect 4753 5893 4767 5907
rect 5033 6072 5047 6086
rect 4993 5973 5007 5987
rect 4833 5933 4847 5947
rect 4913 5933 4927 5947
rect 4793 5893 4807 5907
rect 4873 5894 4887 5908
rect 4693 5852 4707 5866
rect 4733 5852 4747 5866
rect 4773 5852 4787 5866
rect 4813 5852 4827 5866
rect 4853 5852 4867 5866
rect 4813 5813 4827 5827
rect 4813 5733 4827 5747
rect 4733 5713 4747 5727
rect 4693 5633 4707 5647
rect 4433 5513 4447 5527
rect 4493 5552 4507 5566
rect 4653 5553 4667 5567
rect 4613 5533 4627 5547
rect 4593 5513 4607 5527
rect 4633 5513 4647 5527
rect 4453 5493 4467 5507
rect 4533 5493 4547 5507
rect 4533 5433 4547 5447
rect 4413 5413 4427 5427
rect 4633 5473 4647 5487
rect 4853 5693 4867 5707
rect 4813 5673 4827 5687
rect 4773 5594 4787 5608
rect 4833 5633 4847 5647
rect 4693 5493 4707 5507
rect 4673 5473 4687 5487
rect 4613 5413 4627 5427
rect 4433 5374 4447 5388
rect 4493 5373 4507 5387
rect 4553 5374 4567 5388
rect 4593 5374 4607 5388
rect 4112 5333 4126 5347
rect 4133 5332 4147 5346
rect 4173 5332 4187 5346
rect 4253 5333 4267 5347
rect 4213 5293 4227 5307
rect 4313 5332 4327 5346
rect 4373 5333 4387 5347
rect 4293 5313 4307 5327
rect 4353 5293 4367 5307
rect 4233 5253 4247 5267
rect 4153 5213 4167 5227
rect 4173 5193 4187 5207
rect 4133 5153 4147 5167
rect 4113 5133 4127 5147
rect 4153 5133 4167 5147
rect 4093 5093 4107 5107
rect 4133 5093 4147 5107
rect 4113 5074 4127 5088
rect 4013 5033 4027 5047
rect 4013 4973 4027 4987
rect 4073 5013 4087 5027
rect 3993 4913 4007 4927
rect 4053 4913 4067 4927
rect 3973 4873 3987 4887
rect 4033 4873 4047 4887
rect 3993 4854 4007 4868
rect 4133 5033 4147 5047
rect 4113 4993 4127 5007
rect 4093 4973 4107 4987
rect 4133 4933 4147 4947
rect 4113 4913 4127 4927
rect 4193 5152 4207 5166
rect 4333 5233 4347 5247
rect 4293 5193 4307 5207
rect 4333 5193 4347 5207
rect 4253 5173 4267 5187
rect 4233 5093 4247 5107
rect 4493 5332 4507 5346
rect 4533 5332 4547 5346
rect 4453 5293 4467 5307
rect 4413 5273 4427 5287
rect 4373 5213 4387 5227
rect 4473 5253 4487 5267
rect 4453 5213 4467 5227
rect 4413 5133 4427 5147
rect 4413 5093 4427 5107
rect 4233 5032 4247 5046
rect 4213 4993 4227 5007
rect 4193 4953 4207 4967
rect 4193 4913 4207 4927
rect 4173 4893 4187 4907
rect 4193 4873 4207 4887
rect 4073 4854 4087 4868
rect 4133 4854 4147 4868
rect 4193 4852 4207 4866
rect 4313 5033 4327 5047
rect 4273 4973 4287 4987
rect 4233 4953 4247 4967
rect 4313 4953 4327 4967
rect 4213 4833 4227 4847
rect 3973 4812 3987 4826
rect 4013 4812 4027 4826
rect 4073 4813 4087 4827
rect 3953 4753 3967 4767
rect 3933 4713 3947 4727
rect 3913 4673 3927 4687
rect 3813 4554 3827 4568
rect 3793 4153 3807 4167
rect 3753 4073 3767 4087
rect 3733 3992 3747 4006
rect 3833 4513 3847 4527
rect 3853 4473 3867 4487
rect 3893 4473 3907 4487
rect 3993 4693 4007 4707
rect 3993 4653 4007 4667
rect 4073 4773 4087 4787
rect 4053 4713 4067 4727
rect 4013 4554 4027 4568
rect 3933 4453 3947 4467
rect 3993 4493 4007 4507
rect 3973 4413 3987 4427
rect 3953 4393 3967 4407
rect 3953 4353 3967 4367
rect 3833 4333 3847 4347
rect 3833 4293 3847 4307
rect 3873 4293 3887 4307
rect 3813 4113 3827 4127
rect 3913 4253 3927 4267
rect 3673 3893 3687 3907
rect 3653 3833 3667 3847
rect 3733 3833 3747 3847
rect 3673 3814 3687 3828
rect 3653 3753 3667 3767
rect 3333 3613 3347 3627
rect 3373 3613 3387 3627
rect 3493 3613 3507 3627
rect 3533 3613 3547 3627
rect 3613 3613 3627 3627
rect 3693 3693 3707 3707
rect 3653 3593 3667 3607
rect 3573 3553 3587 3567
rect 3333 3514 3347 3528
rect 3373 3514 3387 3528
rect 3433 3514 3447 3528
rect 3493 3514 3507 3528
rect 3533 3514 3547 3528
rect 3293 3473 3307 3487
rect 3273 3453 3287 3467
rect 3253 3413 3267 3427
rect 3193 3393 3207 3407
rect 3313 3453 3327 3467
rect 3253 3373 3267 3387
rect 3293 3373 3307 3387
rect 3213 3333 3227 3347
rect 3193 3313 3207 3327
rect 3133 3093 3147 3107
rect 3173 3093 3187 3107
rect 3293 3294 3307 3308
rect 3213 3252 3227 3266
rect 3273 3252 3287 3266
rect 3233 3233 3247 3247
rect 3293 3233 3307 3247
rect 3273 3193 3287 3207
rect 3253 3173 3267 3187
rect 3253 3113 3267 3127
rect 3233 3053 3247 3067
rect 3172 3033 3186 3047
rect 3193 3033 3207 3047
rect 3093 2994 3107 3008
rect 3153 2994 3167 3008
rect 3033 2953 3047 2967
rect 3013 2913 3027 2927
rect 2953 2873 2967 2887
rect 2873 2853 2887 2867
rect 2893 2813 2907 2827
rect 2973 2813 2987 2827
rect 2833 2774 2847 2788
rect 2913 2773 2927 2787
rect 3013 2774 3027 2788
rect 2773 2732 2787 2746
rect 2573 2653 2587 2667
rect 2593 2633 2607 2647
rect 2553 2613 2567 2627
rect 2513 2533 2527 2547
rect 2513 2512 2527 2526
rect 2473 2473 2487 2487
rect 2533 2432 2547 2446
rect 2493 2373 2507 2387
rect 2633 2673 2647 2687
rect 2753 2693 2767 2707
rect 2693 2653 2707 2667
rect 2713 2633 2727 2647
rect 2693 2613 2707 2627
rect 2693 2573 2707 2587
rect 2673 2553 2687 2567
rect 2713 2513 2727 2527
rect 2633 2493 2647 2507
rect 2613 2474 2627 2488
rect 2673 2474 2687 2488
rect 2713 2473 2727 2487
rect 2493 2352 2507 2366
rect 2593 2353 2607 2367
rect 2653 2353 2667 2367
rect 2473 2313 2487 2327
rect 2673 2333 2687 2347
rect 2593 2313 2607 2327
rect 2433 2233 2447 2247
rect 2413 2153 2427 2167
rect 2433 2133 2447 2147
rect 2413 2113 2427 2127
rect 2473 2113 2487 2127
rect 2513 2113 2527 2127
rect 2393 1993 2407 2007
rect 2553 2193 2567 2207
rect 2553 2093 2567 2107
rect 2533 2073 2547 2087
rect 2453 2053 2467 2067
rect 2513 2053 2527 2067
rect 2433 2033 2447 2047
rect 2453 2013 2467 2027
rect 2433 1993 2447 2007
rect 2533 1993 2547 2007
rect 2713 2393 2727 2407
rect 2713 2293 2727 2307
rect 2713 2233 2727 2247
rect 2633 2212 2647 2226
rect 2633 2173 2647 2187
rect 2753 2493 2767 2507
rect 2853 2732 2867 2746
rect 2893 2733 2907 2747
rect 2813 2693 2827 2707
rect 2793 2653 2807 2667
rect 2993 2732 3007 2746
rect 2913 2693 2927 2707
rect 2953 2693 2967 2707
rect 2893 2653 2907 2667
rect 2853 2593 2867 2607
rect 2793 2573 2807 2587
rect 2853 2553 2867 2567
rect 2833 2513 2847 2527
rect 2973 2673 2987 2687
rect 2953 2653 2967 2667
rect 2933 2573 2947 2587
rect 2893 2473 2907 2487
rect 3073 2952 3087 2966
rect 3193 2994 3207 3008
rect 3233 2994 3247 3008
rect 3313 3153 3327 3167
rect 3393 3473 3407 3487
rect 3913 4073 3927 4087
rect 3833 4034 3847 4048
rect 3873 4034 3887 4048
rect 4013 4473 4027 4487
rect 4013 4433 4027 4447
rect 4053 4413 4067 4427
rect 4153 4812 4167 4826
rect 4193 4813 4207 4827
rect 4113 4793 4127 4807
rect 4173 4793 4187 4807
rect 4093 4653 4107 4667
rect 4153 4613 4167 4627
rect 4113 4554 4127 4568
rect 4193 4713 4207 4727
rect 4293 4933 4307 4947
rect 4353 5033 4367 5047
rect 4313 4812 4327 4826
rect 4333 4773 4347 4787
rect 4233 4733 4247 4747
rect 4273 4733 4287 4747
rect 4213 4693 4227 4707
rect 4193 4653 4207 4667
rect 4173 4553 4187 4567
rect 4373 4973 4387 4987
rect 4433 5013 4447 5027
rect 4393 4893 4407 4907
rect 4453 4973 4467 4987
rect 4493 5233 4507 5247
rect 4513 5193 4527 5207
rect 4553 5173 4567 5187
rect 4573 5153 4587 5167
rect 4553 5113 4567 5127
rect 4492 5073 4506 5087
rect 4513 5074 4527 5088
rect 4573 5074 4587 5088
rect 4493 5033 4507 5047
rect 4533 5033 4547 5047
rect 4473 4873 4487 4887
rect 4433 4854 4447 4868
rect 4513 4873 4527 4887
rect 4493 4853 4507 4867
rect 4413 4812 4427 4826
rect 4453 4813 4467 4827
rect 4453 4773 4467 4787
rect 4553 4953 4567 4967
rect 4713 5433 4727 5447
rect 4813 5553 4827 5567
rect 4772 5493 4786 5507
rect 4793 5493 4807 5507
rect 4773 5453 4787 5467
rect 4833 5513 4847 5527
rect 4953 5913 4967 5927
rect 4933 5893 4947 5907
rect 5033 5894 5047 5908
rect 5013 5853 5027 5867
rect 4953 5733 4967 5747
rect 4933 5673 4947 5687
rect 4853 5493 4867 5507
rect 4913 5593 4927 5607
rect 4852 5453 4866 5467
rect 4873 5453 4887 5467
rect 4753 5413 4767 5427
rect 4832 5413 4846 5427
rect 4853 5413 4867 5427
rect 4653 5332 4667 5346
rect 4713 5313 4727 5327
rect 4653 5213 4667 5227
rect 4633 5153 4647 5167
rect 4793 5374 4807 5388
rect 4873 5374 4887 5388
rect 4753 5313 4767 5327
rect 4793 5313 4807 5327
rect 4733 5213 4747 5227
rect 4773 5173 4787 5187
rect 4693 5074 4707 5088
rect 4633 5013 4647 5027
rect 4613 4933 4627 4947
rect 4633 4913 4647 4927
rect 4713 5032 4727 5046
rect 4873 5293 4887 5307
rect 4933 5552 4947 5566
rect 4913 5473 4927 5487
rect 4893 5253 4907 5267
rect 5133 6114 5147 6128
rect 5113 6072 5127 6086
rect 5093 6053 5107 6067
rect 5113 6033 5127 6047
rect 5173 6073 5187 6087
rect 5653 6233 5667 6247
rect 5333 6193 5347 6207
rect 5273 6153 5287 6167
rect 5213 6133 5227 6147
rect 5213 6073 5227 6087
rect 5293 6073 5307 6087
rect 5193 6053 5207 6067
rect 5213 6033 5227 6047
rect 5153 6013 5167 6027
rect 5213 5993 5227 6007
rect 5113 5953 5127 5967
rect 5113 5893 5127 5907
rect 5153 5894 5167 5908
rect 5253 5933 5267 5947
rect 5213 5893 5227 5907
rect 5313 5894 5327 5908
rect 5133 5852 5147 5866
rect 5093 5833 5107 5847
rect 5173 5833 5187 5847
rect 5113 5773 5127 5787
rect 5153 5773 5167 5787
rect 5093 5753 5107 5767
rect 5073 5673 5087 5687
rect 5053 5613 5067 5627
rect 5153 5733 5167 5747
rect 5133 5693 5147 5707
rect 5113 5633 5127 5647
rect 5153 5653 5167 5667
rect 5153 5593 5167 5607
rect 5073 5552 5087 5566
rect 5113 5552 5127 5566
rect 5033 5513 5047 5527
rect 5013 5493 5027 5507
rect 4953 5374 4967 5388
rect 5013 5413 5027 5427
rect 5073 5453 5087 5467
rect 4993 5373 5007 5387
rect 4993 5333 5007 5347
rect 4973 5313 4987 5327
rect 4973 5253 4987 5267
rect 4973 5213 4987 5227
rect 4913 5193 4927 5207
rect 5013 5313 5027 5327
rect 4933 5153 4947 5167
rect 4993 5153 5007 5167
rect 4833 5113 4847 5127
rect 4813 5093 4827 5107
rect 4913 5093 4927 5107
rect 4873 5074 4887 5088
rect 4733 5013 4747 5027
rect 4773 5013 4787 5027
rect 4673 4973 4687 4987
rect 4553 4893 4567 4907
rect 4653 4893 4667 4907
rect 4553 4854 4567 4868
rect 4593 4854 4607 4868
rect 4533 4813 4547 4827
rect 4553 4793 4567 4807
rect 4373 4753 4387 4767
rect 4413 4753 4427 4767
rect 4533 4753 4547 4767
rect 4353 4693 4367 4707
rect 4333 4673 4347 4687
rect 4333 4633 4347 4647
rect 4273 4613 4287 4627
rect 4253 4554 4267 4568
rect 4293 4554 4307 4568
rect 4193 4512 4207 4526
rect 4233 4512 4247 4526
rect 4132 4493 4146 4507
rect 4153 4493 4167 4507
rect 4073 4353 4087 4367
rect 4053 4334 4067 4348
rect 4093 4334 4107 4348
rect 4373 4512 4387 4526
rect 4213 4473 4227 4487
rect 4292 4473 4306 4487
rect 4313 4473 4327 4487
rect 3993 4292 4007 4306
rect 4033 4292 4047 4306
rect 3973 4253 3987 4267
rect 4013 4153 4027 4167
rect 4133 4293 4147 4307
rect 4093 4253 4107 4267
rect 4073 4113 4087 4127
rect 3973 4073 3987 4087
rect 4013 4073 4027 4087
rect 3953 4033 3967 4047
rect 3833 3993 3847 4007
rect 3853 3973 3867 3987
rect 3833 3933 3847 3947
rect 3752 3813 3766 3827
rect 3773 3813 3787 3827
rect 3813 3813 3827 3827
rect 3893 3913 3907 3927
rect 3933 3913 3947 3927
rect 3873 3853 3887 3867
rect 3853 3813 3867 3827
rect 3793 3772 3807 3786
rect 3853 3773 3867 3787
rect 3753 3733 3767 3747
rect 3693 3533 3707 3547
rect 3733 3533 3747 3547
rect 3633 3514 3647 3528
rect 3753 3514 3767 3528
rect 3793 3513 3807 3527
rect 3373 3453 3387 3467
rect 3433 3413 3447 3427
rect 3393 3333 3407 3347
rect 3433 3313 3447 3327
rect 3413 3294 3427 3308
rect 3473 3472 3487 3486
rect 3473 3393 3487 3407
rect 3493 3313 3507 3327
rect 3473 3293 3487 3307
rect 3373 3193 3387 3207
rect 3433 3252 3447 3266
rect 3493 3252 3507 3266
rect 3573 3472 3587 3486
rect 3653 3472 3667 3486
rect 3693 3472 3707 3486
rect 3773 3473 3787 3487
rect 3573 3433 3587 3447
rect 3733 3433 3747 3447
rect 3553 3313 3567 3327
rect 3613 3313 3627 3327
rect 3693 3313 3707 3327
rect 3733 3313 3747 3327
rect 3573 3252 3587 3266
rect 3613 3253 3627 3267
rect 3793 3333 3807 3347
rect 3933 3814 3947 3828
rect 4053 4053 4067 4067
rect 4073 4033 4087 4047
rect 4033 3992 4047 4006
rect 4133 4193 4147 4207
rect 4113 4073 4127 4087
rect 3993 3973 4007 3987
rect 4093 3973 4107 3987
rect 4073 3853 4087 3867
rect 4013 3816 4027 3830
rect 4193 4293 4207 4307
rect 4193 4173 4207 4187
rect 4173 4113 4187 4127
rect 4373 4433 4387 4447
rect 4233 4413 4247 4427
rect 4293 4373 4307 4387
rect 4393 4353 4407 4367
rect 4253 4233 4267 4247
rect 4233 4153 4247 4167
rect 4233 4113 4247 4127
rect 4313 4113 4327 4127
rect 4213 4053 4227 4067
rect 4133 4033 4147 4047
rect 4193 4034 4207 4048
rect 4353 4093 4367 4107
rect 4253 4034 4267 4048
rect 4133 3993 4147 4007
rect 4113 3833 4127 3847
rect 4213 3992 4227 4006
rect 4373 4073 4387 4087
rect 4213 3913 4227 3927
rect 4173 3893 4187 3907
rect 4213 3892 4227 3906
rect 4153 3816 4167 3830
rect 3993 3793 4007 3807
rect 3893 3773 3907 3787
rect 3893 3673 3907 3687
rect 3953 3772 3967 3786
rect 3893 3633 3907 3647
rect 3873 3533 3887 3547
rect 4013 3693 4027 3707
rect 3933 3513 3947 3527
rect 4013 3493 4027 3507
rect 3833 3413 3847 3427
rect 3953 3470 3967 3484
rect 4213 3773 4227 3787
rect 4213 3752 4227 3766
rect 4093 3713 4107 3727
rect 4053 3673 4067 3687
rect 4153 3653 4167 3667
rect 4073 3533 4087 3547
rect 4173 3573 4187 3587
rect 4033 3453 4047 3467
rect 4073 3453 4087 3467
rect 4053 3413 4067 3427
rect 3913 3393 3927 3407
rect 3993 3353 4007 3367
rect 3873 3333 3887 3347
rect 3673 3252 3687 3266
rect 3653 3233 3667 3247
rect 3513 3213 3527 3227
rect 3433 3193 3447 3207
rect 3393 3153 3407 3167
rect 3313 3013 3327 3027
rect 3353 3013 3367 3027
rect 3153 2933 3167 2947
rect 3073 2913 3087 2927
rect 3113 2913 3127 2927
rect 3053 2573 3067 2587
rect 3213 2952 3227 2966
rect 3253 2952 3267 2966
rect 3293 2953 3307 2967
rect 3233 2933 3247 2947
rect 3173 2893 3187 2907
rect 3173 2833 3187 2847
rect 3233 2732 3247 2746
rect 3293 2893 3307 2907
rect 3373 2994 3387 3008
rect 3353 2853 3367 2867
rect 3393 2853 3407 2867
rect 3313 2793 3327 2807
rect 3353 2774 3367 2788
rect 3413 2793 3427 2807
rect 3393 2773 3407 2787
rect 3093 2653 3107 2667
rect 3113 2593 3127 2607
rect 3073 2513 3087 2527
rect 2933 2453 2947 2467
rect 2753 2431 2767 2445
rect 2792 2431 2806 2445
rect 2813 2433 2827 2447
rect 2913 2413 2927 2427
rect 2853 2373 2867 2387
rect 2833 2353 2847 2367
rect 2833 2313 2847 2327
rect 2813 2293 2827 2307
rect 2893 2254 2907 2268
rect 2933 2254 2947 2268
rect 2753 2213 2767 2227
rect 2913 2212 2927 2226
rect 2733 2193 2747 2207
rect 2773 2193 2787 2207
rect 2613 2153 2627 2167
rect 2472 1953 2486 1967
rect 2513 1954 2527 1968
rect 2593 1973 2607 1987
rect 2573 1954 2587 1968
rect 2433 1912 2447 1926
rect 2493 1912 2507 1926
rect 2393 1893 2407 1907
rect 2453 1853 2467 1867
rect 2553 1853 2567 1867
rect 2373 1833 2387 1847
rect 2392 1813 2406 1827
rect 2413 1813 2427 1827
rect 2413 1773 2427 1787
rect 2393 1753 2407 1767
rect 2493 1793 2507 1807
rect 2373 1692 2387 1706
rect 2473 1693 2487 1707
rect 2273 1353 2287 1367
rect 2313 1353 2327 1367
rect 2212 1233 2226 1247
rect 2233 1233 2247 1247
rect 2172 1213 2186 1227
rect 2193 1214 2207 1228
rect 2313 1293 2327 1307
rect 2413 1533 2427 1547
rect 2373 1434 2387 1448
rect 2433 1513 2447 1527
rect 2433 1473 2447 1487
rect 2293 1213 2307 1227
rect 2113 1172 2127 1186
rect 2153 1172 2167 1186
rect 2213 1172 2227 1186
rect 2253 1172 2267 1186
rect 2293 1172 2307 1186
rect 2073 1153 2087 1167
rect 2033 1073 2047 1087
rect 1993 953 2007 967
rect 2093 1033 2107 1047
rect 2073 993 2087 1007
rect 2033 914 2047 928
rect 2193 993 2207 1007
rect 2153 973 2167 987
rect 2133 953 2147 967
rect 1913 872 1927 886
rect 1953 872 1967 886
rect 1993 872 2007 886
rect 1953 813 1967 827
rect 1932 773 1946 787
rect 1953 773 1967 787
rect 1913 753 1927 767
rect 1833 713 1847 727
rect 1753 693 1767 707
rect 1793 694 1807 708
rect 1573 652 1587 666
rect 1493 633 1507 647
rect 1473 613 1487 627
rect 1673 652 1687 666
rect 1733 653 1747 667
rect 1773 653 1787 667
rect 1753 633 1767 647
rect 1633 613 1647 627
rect 1493 593 1507 607
rect 1653 573 1667 587
rect 1613 553 1627 567
rect 1413 453 1427 467
rect 1573 433 1587 447
rect 1393 413 1407 427
rect 1473 394 1487 408
rect 1413 373 1427 387
rect 1393 333 1407 347
rect 1373 313 1387 327
rect 1493 293 1507 307
rect 1473 253 1487 267
rect 1293 233 1307 247
rect 1333 174 1347 188
rect 1393 174 1407 188
rect 1433 174 1447 188
rect 1213 132 1227 146
rect 1273 113 1287 127
rect 893 93 907 107
rect 1213 93 1227 107
rect 1253 92 1267 106
rect 1413 132 1427 146
rect 1473 132 1487 146
rect 1373 113 1387 127
rect 1533 273 1547 287
rect 1513 233 1527 247
rect 1853 652 1867 666
rect 1813 533 1827 547
rect 1693 493 1707 507
rect 1653 394 1667 408
rect 1913 693 1927 707
rect 1993 733 2007 747
rect 2173 953 2187 967
rect 2093 872 2107 886
rect 2153 872 2167 886
rect 2053 853 2067 867
rect 2073 793 2087 807
rect 2153 793 2167 807
rect 1933 652 1947 666
rect 1973 593 1987 607
rect 1893 573 1907 587
rect 2053 693 2067 707
rect 2113 694 2127 708
rect 2233 914 2247 928
rect 2413 1373 2427 1387
rect 2333 1233 2347 1247
rect 2393 1233 2407 1247
rect 2313 1153 2327 1167
rect 2373 1214 2387 1228
rect 2553 1734 2567 1748
rect 2673 2093 2687 2107
rect 2713 2013 2727 2027
rect 2673 1954 2687 1968
rect 2753 2073 2767 2087
rect 2753 1933 2767 1947
rect 2653 1913 2667 1927
rect 3033 2493 3047 2507
rect 2973 2473 2987 2487
rect 3013 2474 3027 2488
rect 2993 2433 3007 2447
rect 2973 2393 2987 2407
rect 2973 2353 2987 2367
rect 3073 2432 3087 2446
rect 3033 2413 3047 2427
rect 3073 2411 3087 2425
rect 2993 2313 3007 2327
rect 3033 2313 3047 2327
rect 2993 2254 3007 2268
rect 3213 2573 3227 2587
rect 3173 2474 3187 2488
rect 3133 2373 3147 2387
rect 3113 2353 3127 2367
rect 3073 2254 3087 2268
rect 3173 2254 3187 2268
rect 2993 2213 3007 2227
rect 3053 2193 3067 2207
rect 3153 2193 3167 2207
rect 3173 2173 3187 2187
rect 2973 2153 2987 2167
rect 2953 2133 2967 2147
rect 2853 1973 2867 1987
rect 2913 1954 2927 1968
rect 2953 1954 2967 1968
rect 3013 1954 3027 1968
rect 3073 1954 3087 1968
rect 2633 1793 2647 1807
rect 2633 1753 2647 1767
rect 2713 1833 2727 1847
rect 2693 1793 2707 1807
rect 2753 1813 2767 1827
rect 2713 1773 2727 1787
rect 2653 1733 2667 1747
rect 2693 1734 2707 1748
rect 2533 1692 2547 1706
rect 2493 1653 2507 1667
rect 2612 1692 2626 1706
rect 2633 1693 2647 1707
rect 2673 1692 2687 1706
rect 2733 1692 2747 1706
rect 2973 1912 2987 1926
rect 2873 1893 2887 1907
rect 2913 1893 2927 1907
rect 2972 1891 2986 1905
rect 2993 1893 3007 1907
rect 2833 1853 2847 1867
rect 2913 1833 2927 1847
rect 2793 1793 2807 1807
rect 2853 1773 2867 1787
rect 2813 1692 2827 1706
rect 2673 1653 2687 1667
rect 2573 1633 2587 1647
rect 2613 1633 2627 1647
rect 2472 1453 2486 1467
rect 2493 1453 2507 1467
rect 2573 1453 2587 1467
rect 2473 1432 2487 1446
rect 2513 1434 2527 1448
rect 2633 1453 2647 1467
rect 2673 1434 2687 1448
rect 2533 1392 2547 1406
rect 2513 1353 2527 1367
rect 2613 1353 2627 1367
rect 2473 1253 2487 1267
rect 2333 1093 2347 1107
rect 2333 1072 2347 1086
rect 2293 913 2307 927
rect 2393 1172 2407 1186
rect 2433 1172 2447 1186
rect 2513 1233 2527 1247
rect 2553 1214 2567 1228
rect 2813 1633 2827 1647
rect 2893 1692 2907 1706
rect 2873 1533 2887 1547
rect 2833 1453 2847 1467
rect 2753 1434 2767 1448
rect 2793 1434 2807 1448
rect 2753 1373 2767 1387
rect 2793 1373 2807 1387
rect 2733 1353 2747 1367
rect 2753 1333 2767 1347
rect 2673 1313 2687 1327
rect 2653 1293 2667 1307
rect 2633 1213 2647 1227
rect 2713 1233 2727 1247
rect 2873 1393 2887 1407
rect 2813 1333 2827 1347
rect 2853 1333 2867 1347
rect 2753 1293 2767 1307
rect 2793 1293 2807 1307
rect 2733 1213 2747 1227
rect 2373 1093 2387 1107
rect 2373 1053 2387 1067
rect 2353 1033 2367 1047
rect 2533 1153 2547 1167
rect 2573 1153 2587 1167
rect 2513 1053 2527 1067
rect 2453 1013 2467 1027
rect 2453 953 2467 967
rect 2393 914 2407 928
rect 2433 913 2447 927
rect 2373 872 2387 886
rect 2253 813 2267 827
rect 2193 773 2207 787
rect 2393 793 2407 807
rect 2373 753 2387 767
rect 2193 733 2207 747
rect 2253 733 2267 747
rect 2293 733 2307 747
rect 2353 733 2367 747
rect 2033 553 2047 567
rect 2013 533 2027 547
rect 2033 513 2047 527
rect 1853 473 1867 487
rect 1713 453 1727 467
rect 1813 453 1827 467
rect 1733 394 1747 408
rect 1773 394 1787 408
rect 1973 433 1987 447
rect 1853 394 1867 408
rect 1933 394 1947 408
rect 1833 352 1847 366
rect 1953 352 1967 366
rect 1733 333 1747 347
rect 2093 633 2107 647
rect 2133 593 2147 607
rect 2053 394 2067 408
rect 2213 713 2227 727
rect 2213 652 2227 666
rect 2273 652 2287 666
rect 2313 652 2327 666
rect 2193 633 2207 647
rect 2273 553 2287 567
rect 2373 693 2387 707
rect 2553 973 2567 987
rect 2533 953 2547 967
rect 2553 914 2567 928
rect 2453 873 2467 887
rect 2473 813 2487 827
rect 2433 733 2447 747
rect 2413 713 2427 727
rect 2473 693 2487 707
rect 2453 652 2467 666
rect 2533 872 2547 886
rect 2633 1053 2647 1067
rect 2673 1053 2687 1067
rect 2773 1273 2787 1287
rect 2753 1153 2767 1167
rect 2693 973 2707 987
rect 2853 1253 2867 1267
rect 3033 1853 3047 1867
rect 3013 1833 3027 1847
rect 2993 1773 3007 1787
rect 2933 1733 2947 1747
rect 2933 1633 2947 1647
rect 2913 1593 2927 1607
rect 2973 1553 2987 1567
rect 2973 1453 2987 1467
rect 3073 1793 3087 1807
rect 3153 1913 3167 1927
rect 3113 1873 3127 1887
rect 3153 1873 3167 1887
rect 3113 1773 3127 1787
rect 3093 1753 3107 1767
rect 3093 1692 3107 1706
rect 3153 1653 3167 1667
rect 3073 1613 3087 1627
rect 3073 1453 3087 1467
rect 3033 1433 3047 1447
rect 3113 1434 3127 1448
rect 3152 1434 3166 1448
rect 3273 2673 3287 2687
rect 3333 2733 3347 2747
rect 3313 2713 3327 2727
rect 3313 2633 3327 2647
rect 3293 2593 3307 2607
rect 3313 2573 3327 2587
rect 3273 2533 3287 2547
rect 3393 2733 3407 2747
rect 3373 2633 3387 2647
rect 3373 2593 3387 2607
rect 3333 2553 3347 2567
rect 3293 2493 3307 2507
rect 3353 2533 3367 2547
rect 3333 2474 3347 2488
rect 3273 2432 3287 2446
rect 3313 2413 3327 2427
rect 3593 3093 3607 3107
rect 3533 3053 3547 3067
rect 3453 3033 3467 3047
rect 3493 2994 3507 3008
rect 3773 3252 3787 3266
rect 3713 3113 3727 3127
rect 3833 3294 3847 3308
rect 3933 3313 3947 3327
rect 4033 3294 4047 3308
rect 3853 3252 3867 3266
rect 3893 3252 3907 3266
rect 3933 3252 3947 3266
rect 4013 3252 4027 3266
rect 3973 3233 3987 3247
rect 3833 3213 3847 3227
rect 3993 3213 4007 3227
rect 3833 3173 3847 3187
rect 3833 3133 3847 3147
rect 3793 3093 3807 3107
rect 3813 3073 3827 3087
rect 3693 2994 3707 3008
rect 3813 2994 3827 3008
rect 3453 2952 3467 2966
rect 3513 2952 3527 2966
rect 3453 2853 3467 2867
rect 3433 2773 3447 2787
rect 3493 2774 3507 2788
rect 3513 2732 3527 2746
rect 3473 2713 3487 2727
rect 3413 2533 3427 2547
rect 3593 2952 3607 2966
rect 3633 2952 3647 2966
rect 3573 2933 3587 2947
rect 3753 2950 3767 2964
rect 3733 2893 3747 2907
rect 4313 3992 4327 4006
rect 4353 3992 4367 4006
rect 4253 3813 4267 3827
rect 4273 3770 4287 3784
rect 4233 3713 4247 3727
rect 4353 3653 4367 3667
rect 4333 3633 4347 3647
rect 4253 3613 4267 3627
rect 4233 3513 4247 3527
rect 4492 4713 4506 4727
rect 4513 4713 4527 4727
rect 4493 4653 4507 4667
rect 4452 4593 4466 4607
rect 4473 4593 4487 4607
rect 4453 4554 4467 4568
rect 4533 4613 4547 4627
rect 4513 4573 4527 4587
rect 4493 4453 4507 4467
rect 4473 4413 4487 4427
rect 4453 4393 4467 4407
rect 4513 4433 4527 4447
rect 4512 4373 4526 4387
rect 4533 4373 4547 4387
rect 4573 4773 4587 4787
rect 4733 4973 4747 4987
rect 4713 4953 4727 4967
rect 4733 4933 4747 4947
rect 4773 4933 4787 4947
rect 4733 4873 4747 4887
rect 4713 4854 4727 4868
rect 4753 4854 4767 4868
rect 4813 5032 4827 5046
rect 4853 4993 4867 5007
rect 4833 4973 4847 4987
rect 4673 4832 4687 4846
rect 4773 4812 4787 4826
rect 4673 4773 4687 4787
rect 4653 4753 4667 4767
rect 4633 4713 4647 4727
rect 4693 4713 4707 4727
rect 4613 4673 4627 4687
rect 4613 4652 4627 4666
rect 4573 4593 4587 4607
rect 4573 4553 4587 4567
rect 4653 4633 4667 4647
rect 4633 4613 4647 4627
rect 4633 4573 4647 4587
rect 4573 4513 4587 4527
rect 4593 4493 4607 4507
rect 4573 4473 4587 4487
rect 4553 4353 4567 4367
rect 4613 4473 4627 4487
rect 4593 4433 4607 4447
rect 4712 4693 4726 4707
rect 4733 4693 4747 4707
rect 4813 4673 4827 4687
rect 4853 4873 4867 4887
rect 4993 5113 5007 5127
rect 5033 5293 5047 5307
rect 5153 5493 5167 5507
rect 5153 5433 5167 5447
rect 5133 5373 5147 5387
rect 5233 5852 5247 5866
rect 5273 5852 5287 5866
rect 5193 5813 5207 5827
rect 5293 5813 5307 5827
rect 5193 5753 5207 5767
rect 5293 5733 5307 5747
rect 5233 5713 5247 5727
rect 5193 5673 5207 5687
rect 5253 5693 5267 5707
rect 5233 5613 5247 5627
rect 5273 5653 5287 5667
rect 5313 5693 5327 5707
rect 5293 5633 5307 5647
rect 5273 5593 5287 5607
rect 5213 5552 5227 5566
rect 5193 5512 5207 5526
rect 5193 5473 5207 5487
rect 5193 5393 5207 5407
rect 5173 5373 5187 5387
rect 5093 5333 5107 5347
rect 5073 5273 5087 5287
rect 5053 5253 5067 5267
rect 5053 5213 5067 5227
rect 5033 5173 5047 5187
rect 4993 5032 5007 5046
rect 4953 4973 4967 4987
rect 4933 4893 4947 4907
rect 4933 4853 4947 4867
rect 4893 4812 4907 4826
rect 4873 4773 4887 4787
rect 4893 4753 4907 4767
rect 4873 4673 4887 4687
rect 4733 4592 4747 4606
rect 4813 4593 4827 4607
rect 4713 4573 4727 4587
rect 4653 4493 4667 4507
rect 4633 4433 4647 4447
rect 4613 4413 4627 4427
rect 4593 4353 4607 4367
rect 4693 4512 4707 4526
rect 4673 4473 4687 4487
rect 4653 4413 4667 4427
rect 4633 4393 4647 4407
rect 4693 4353 4707 4367
rect 4552 4293 4566 4307
rect 4573 4293 4587 4307
rect 4633 4334 4647 4348
rect 4673 4334 4687 4348
rect 4893 4573 4907 4587
rect 4773 4473 4787 4487
rect 4753 4453 4767 4467
rect 4733 4413 4747 4427
rect 4733 4392 4747 4406
rect 4613 4293 4627 4307
rect 4473 4233 4487 4247
rect 4513 4213 4527 4227
rect 4453 4113 4467 4127
rect 4413 4073 4427 4087
rect 4393 4033 4407 4047
rect 4393 3993 4407 4007
rect 4553 4113 4567 4127
rect 4593 4034 4607 4048
rect 4693 4292 4707 4306
rect 4633 4273 4647 4287
rect 4673 4273 4687 4287
rect 4633 4133 4647 4147
rect 4633 4112 4647 4126
rect 4413 3933 4427 3947
rect 4433 3893 4447 3907
rect 4413 3814 4427 3828
rect 4493 3814 4507 3828
rect 4393 3753 4407 3767
rect 4573 3992 4587 4006
rect 4613 3993 4627 4007
rect 4553 3952 4567 3966
rect 4593 3953 4607 3967
rect 4773 4393 4787 4407
rect 4813 4453 4827 4467
rect 4813 4373 4827 4387
rect 4993 4933 5007 4947
rect 5073 5193 5087 5207
rect 5053 5013 5067 5027
rect 5033 4913 5047 4927
rect 4993 4854 5007 4868
rect 5033 4854 5047 4868
rect 5133 5233 5147 5247
rect 5113 5153 5127 5167
rect 5233 5453 5247 5467
rect 5313 5493 5327 5507
rect 5253 5413 5267 5427
rect 5233 5393 5247 5407
rect 5213 5373 5227 5387
rect 5273 5393 5287 5407
rect 5253 5332 5267 5346
rect 5213 5273 5227 5287
rect 5173 5113 5187 5127
rect 5153 5093 5167 5107
rect 5093 5073 5107 5087
rect 5193 5093 5207 5107
rect 5093 5033 5107 5047
rect 5073 4853 5087 4867
rect 4993 4793 5007 4807
rect 4973 4593 4987 4607
rect 4953 4573 4967 4587
rect 5073 4813 5087 4827
rect 5013 4713 5027 4727
rect 5073 4633 5087 4647
rect 5173 5032 5187 5046
rect 5153 5013 5167 5027
rect 5133 4953 5147 4967
rect 5113 4913 5127 4927
rect 5613 6173 5627 6187
rect 5593 6153 5607 6167
rect 5433 6133 5447 6147
rect 5473 6133 5487 6147
rect 5513 6133 5527 6147
rect 5553 6133 5567 6147
rect 5393 6114 5407 6128
rect 5493 6114 5507 6128
rect 5593 6113 5607 6127
rect 5373 6073 5387 6087
rect 5473 6073 5487 6087
rect 5413 6033 5427 6047
rect 5513 6072 5527 6086
rect 5573 6072 5587 6086
rect 5473 6013 5487 6027
rect 5373 5993 5387 6007
rect 5413 5993 5427 6007
rect 5373 5894 5387 5908
rect 5533 5953 5547 5967
rect 5493 5933 5507 5947
rect 5473 5894 5487 5908
rect 5393 5852 5407 5866
rect 5473 5813 5487 5827
rect 5453 5773 5467 5787
rect 5473 5713 5487 5727
rect 5453 5693 5467 5707
rect 5533 5894 5547 5908
rect 5573 5894 5587 5908
rect 5553 5852 5567 5866
rect 5513 5753 5527 5767
rect 5533 5693 5547 5707
rect 5633 6153 5647 6167
rect 5853 6253 5867 6267
rect 5893 6213 5907 6227
rect 5833 6173 5847 6187
rect 5813 6133 5827 6147
rect 5733 6114 5747 6128
rect 5793 6093 5807 6107
rect 5713 6072 5727 6086
rect 5753 6053 5767 6067
rect 5653 6033 5667 6047
rect 5733 6033 5747 6047
rect 5753 5993 5767 6007
rect 5793 5993 5807 6007
rect 5733 5973 5747 5987
rect 5653 5953 5667 5967
rect 5693 5933 5707 5947
rect 5673 5852 5687 5866
rect 5713 5852 5727 5866
rect 5673 5793 5687 5807
rect 5513 5593 5527 5607
rect 5493 5552 5507 5566
rect 5433 5513 5447 5527
rect 5413 5493 5427 5507
rect 5333 5453 5347 5467
rect 5332 5413 5346 5427
rect 5353 5413 5367 5427
rect 5393 5393 5407 5407
rect 5353 5373 5367 5387
rect 5513 5533 5527 5547
rect 5493 5453 5507 5467
rect 5433 5374 5447 5388
rect 5613 5673 5627 5687
rect 5573 5594 5587 5608
rect 5613 5593 5627 5607
rect 5593 5552 5607 5566
rect 5573 5533 5587 5547
rect 5533 5413 5547 5427
rect 5593 5473 5607 5487
rect 5573 5373 5587 5387
rect 5333 5333 5347 5347
rect 5373 5332 5387 5346
rect 5413 5332 5427 5346
rect 5513 5332 5527 5346
rect 5553 5332 5567 5346
rect 5493 5293 5507 5307
rect 5413 5273 5427 5287
rect 5413 5233 5427 5247
rect 5313 5213 5327 5227
rect 5373 5213 5387 5227
rect 5253 5193 5267 5207
rect 5372 5173 5386 5187
rect 5393 5173 5407 5187
rect 5253 5074 5267 5088
rect 5293 5074 5307 5088
rect 5352 5074 5366 5088
rect 5373 5074 5387 5088
rect 5453 5153 5467 5167
rect 5213 4973 5227 4987
rect 5173 4873 5187 4887
rect 5233 4873 5247 4887
rect 5133 4853 5147 4867
rect 5193 4854 5207 4868
rect 5313 4993 5327 5007
rect 5333 4973 5347 4987
rect 5413 5074 5427 5088
rect 5473 5113 5487 5127
rect 5453 5073 5467 5087
rect 5433 5032 5447 5046
rect 5413 4993 5427 5007
rect 5373 4973 5387 4987
rect 5353 4953 5367 4967
rect 5373 4933 5387 4947
rect 5333 4893 5347 4907
rect 5273 4873 5287 4887
rect 5253 4853 5267 4867
rect 5113 4812 5127 4826
rect 5133 4773 5147 4787
rect 5173 4812 5187 4826
rect 5433 4973 5447 4987
rect 5233 4793 5247 4807
rect 5173 4733 5187 4747
rect 5213 4733 5227 4747
rect 5213 4693 5227 4707
rect 5153 4633 5167 4647
rect 5213 4633 5227 4647
rect 5093 4613 5107 4627
rect 5193 4613 5207 4627
rect 5053 4552 5067 4566
rect 5113 4554 5127 4568
rect 5153 4554 5167 4568
rect 5033 4533 5047 4547
rect 4953 4512 4967 4526
rect 4993 4493 5007 4507
rect 4913 4433 4927 4447
rect 4913 4393 4927 4407
rect 4793 4334 4807 4348
rect 4833 4334 4847 4348
rect 4893 4334 4907 4348
rect 4993 4353 5007 4367
rect 4973 4333 4987 4347
rect 4733 4153 4747 4167
rect 4673 4113 4687 4127
rect 4653 4093 4667 4107
rect 4693 4034 4707 4048
rect 4753 4033 4767 4047
rect 4633 3973 4647 3987
rect 4613 3873 4627 3887
rect 4553 3813 4567 3827
rect 4453 3753 4467 3767
rect 4493 3733 4507 3747
rect 4413 3713 4427 3727
rect 4453 3713 4467 3727
rect 4373 3573 4387 3587
rect 4373 3514 4387 3528
rect 4213 3373 4227 3387
rect 4093 3313 4107 3327
rect 4173 3313 4187 3327
rect 4073 3173 4087 3187
rect 4053 3113 4067 3127
rect 4013 3093 4027 3107
rect 3993 3053 4007 3067
rect 3873 3033 3887 3047
rect 3933 2996 3947 3010
rect 3973 2996 3987 3010
rect 3773 2873 3787 2887
rect 3813 2873 3827 2887
rect 3673 2853 3687 2867
rect 3733 2853 3747 2867
rect 3613 2774 3627 2788
rect 3653 2774 3667 2788
rect 3713 2773 3727 2787
rect 3613 2673 3627 2687
rect 3573 2593 3587 2607
rect 3493 2493 3507 2507
rect 3553 2493 3567 2507
rect 3393 2474 3407 2488
rect 3453 2474 3467 2488
rect 3473 2433 3487 2447
rect 3373 2313 3387 2327
rect 3413 2273 3427 2287
rect 3273 2253 3287 2267
rect 3353 2254 3367 2268
rect 3393 2254 3407 2268
rect 3273 2193 3287 2207
rect 3233 2173 3247 2187
rect 3253 2153 3267 2167
rect 3213 2093 3227 2107
rect 3213 2013 3227 2027
rect 3313 2113 3327 2127
rect 3393 2053 3407 2067
rect 3573 2474 3587 2488
rect 3633 2633 3647 2647
rect 3513 2453 3527 2467
rect 3513 2413 3527 2427
rect 3553 2393 3567 2407
rect 3513 2313 3527 2327
rect 3493 2273 3507 2287
rect 3473 2253 3487 2267
rect 3533 2293 3547 2307
rect 3513 2213 3527 2227
rect 3453 2073 3467 2087
rect 3352 1993 3366 2007
rect 3373 1993 3387 2007
rect 3253 1954 3267 1968
rect 3293 1954 3307 1968
rect 3353 1954 3367 1968
rect 3413 1954 3427 1968
rect 3193 1912 3207 1926
rect 3233 1912 3247 1926
rect 3293 1893 3307 1907
rect 3293 1853 3307 1867
rect 3393 1813 3407 1827
rect 3333 1793 3347 1807
rect 3253 1773 3267 1787
rect 3253 1734 3267 1748
rect 3393 1734 3407 1748
rect 3453 1733 3467 1747
rect 3293 1692 3307 1706
rect 3333 1693 3347 1707
rect 3373 1692 3387 1706
rect 3413 1693 3427 1707
rect 3693 2732 3707 2746
rect 3693 2633 3707 2647
rect 3753 2813 3767 2827
rect 3773 2773 3787 2787
rect 3813 2774 3827 2788
rect 3793 2732 3807 2746
rect 3833 2732 3847 2746
rect 3753 2673 3767 2687
rect 3753 2593 3767 2607
rect 3773 2553 3787 2567
rect 3753 2533 3767 2547
rect 3673 2433 3687 2447
rect 3613 2333 3627 2347
rect 3653 2333 3667 2347
rect 3733 2473 3747 2487
rect 3933 2813 3947 2827
rect 3873 2774 3887 2788
rect 4033 2994 4047 3008
rect 4073 2994 4087 3008
rect 4153 3294 4167 3308
rect 4193 3294 4207 3308
rect 4232 3293 4246 3307
rect 4253 3294 4267 3308
rect 4293 3294 4307 3308
rect 4393 3473 4407 3487
rect 4373 3313 4387 3327
rect 4113 3252 4127 3266
rect 4113 3213 4127 3227
rect 4113 3153 4127 3167
rect 3993 2953 4007 2967
rect 3993 2893 4007 2907
rect 3973 2793 3987 2807
rect 3873 2733 3887 2747
rect 3913 2732 3927 2746
rect 3853 2693 3867 2707
rect 3933 2693 3947 2707
rect 3853 2653 3867 2667
rect 3833 2473 3847 2487
rect 3753 2432 3767 2446
rect 3793 2432 3807 2446
rect 3553 2273 3567 2287
rect 3593 2273 3607 2287
rect 3533 2193 3547 2207
rect 3613 2254 3627 2268
rect 3653 2256 3667 2270
rect 3573 2193 3587 2207
rect 3593 2173 3607 2187
rect 3733 2333 3747 2347
rect 3833 2333 3847 2347
rect 3713 2153 3727 2167
rect 3573 2093 3587 2107
rect 3593 2073 3607 2087
rect 3553 2033 3567 2047
rect 3513 1993 3527 2007
rect 3553 1973 3567 1987
rect 3653 2033 3667 2047
rect 3633 1973 3647 1987
rect 3533 1912 3547 1926
rect 3533 1873 3547 1887
rect 3633 1912 3647 1926
rect 3573 1853 3587 1867
rect 3493 1734 3507 1748
rect 3533 1734 3547 1748
rect 3573 1733 3587 1747
rect 3333 1672 3347 1686
rect 3233 1613 3247 1627
rect 3253 1593 3267 1607
rect 3273 1513 3287 1527
rect 3253 1493 3267 1507
rect 3193 1453 3207 1467
rect 2893 1373 2907 1387
rect 2813 1214 2827 1228
rect 2953 1392 2967 1406
rect 2993 1392 3007 1406
rect 2953 1333 2967 1347
rect 2913 1214 2927 1228
rect 2793 1173 2807 1187
rect 2873 1172 2887 1186
rect 2913 1172 2927 1186
rect 2973 1172 2987 1186
rect 3053 1392 3067 1406
rect 3093 1353 3107 1367
rect 3133 1353 3147 1367
rect 3093 1293 3107 1307
rect 3033 1253 3047 1267
rect 3093 1233 3107 1247
rect 3073 1214 3087 1228
rect 3113 1214 3127 1228
rect 3173 1433 3187 1447
rect 3253 1434 3267 1448
rect 3293 1453 3307 1467
rect 3312 1434 3326 1448
rect 3473 1692 3487 1706
rect 3693 1954 3707 1968
rect 3993 2733 4007 2747
rect 3993 2653 4007 2667
rect 3953 2553 3967 2567
rect 4053 2952 4067 2966
rect 4093 2953 4107 2967
rect 4173 3252 4187 3266
rect 4153 3213 4167 3227
rect 4133 3073 4147 3087
rect 4133 3033 4147 3047
rect 4133 2973 4147 2987
rect 4213 3173 4227 3187
rect 4213 3093 4227 3107
rect 4173 3053 4187 3067
rect 4353 3293 4367 3307
rect 4253 3253 4267 3267
rect 4313 3253 4327 3267
rect 4353 3253 4367 3267
rect 4333 3233 4347 3247
rect 4413 3453 4427 3467
rect 4433 3433 4447 3447
rect 4413 3393 4427 3407
rect 4413 3333 4427 3347
rect 4493 3633 4507 3647
rect 4573 3772 4587 3786
rect 4713 3992 4727 4006
rect 4753 3992 4767 4006
rect 4673 3973 4687 3987
rect 4653 3933 4667 3947
rect 4653 3733 4667 3747
rect 4553 3713 4567 3727
rect 4633 3713 4647 3727
rect 4533 3633 4547 3647
rect 4513 3593 4527 3607
rect 4473 3553 4487 3567
rect 4533 3553 4547 3567
rect 4493 3514 4507 3528
rect 4653 3693 4667 3707
rect 4633 3593 4647 3607
rect 4553 3513 4567 3527
rect 4473 3473 4487 3487
rect 4533 3453 4547 3467
rect 4513 3393 4527 3407
rect 4473 3333 4487 3347
rect 4453 3313 4467 3327
rect 4473 3294 4487 3308
rect 4393 3233 4407 3247
rect 4433 3233 4447 3247
rect 4373 3213 4387 3227
rect 4353 3133 4367 3147
rect 4313 3073 4327 3087
rect 4413 3113 4427 3127
rect 4293 3053 4307 3067
rect 4393 3053 4407 3067
rect 4233 3033 4247 3047
rect 4273 3033 4287 3047
rect 4233 2994 4247 3008
rect 4153 2933 4167 2947
rect 4113 2893 4127 2907
rect 4093 2873 4107 2887
rect 4033 2833 4047 2847
rect 4213 2952 4227 2966
rect 4273 2953 4287 2967
rect 4253 2933 4267 2947
rect 4413 3013 4427 3027
rect 4353 2994 4367 3008
rect 4393 2994 4407 3008
rect 4513 3133 4527 3147
rect 4493 3113 4507 3127
rect 4433 2993 4447 3007
rect 4293 2913 4307 2927
rect 4273 2873 4287 2887
rect 4173 2853 4187 2867
rect 4253 2853 4267 2867
rect 4253 2813 4267 2827
rect 4113 2793 4127 2807
rect 4093 2773 4107 2787
rect 4153 2773 4167 2787
rect 4193 2774 4207 2788
rect 4233 2774 4247 2788
rect 4413 2953 4427 2967
rect 4333 2913 4347 2927
rect 4373 2913 4387 2927
rect 4333 2873 4347 2887
rect 4273 2773 4287 2787
rect 4073 2732 4087 2746
rect 4033 2693 4047 2707
rect 4073 2573 4087 2587
rect 3893 2474 3907 2488
rect 3913 2393 3927 2407
rect 4013 2533 4027 2547
rect 4033 2493 4047 2507
rect 4093 2533 4107 2547
rect 4073 2473 4087 2487
rect 4013 2432 4027 2446
rect 4073 2432 4087 2446
rect 4053 2413 4067 2427
rect 3953 2373 3967 2387
rect 4013 2373 4027 2387
rect 3873 2293 3887 2307
rect 3933 2273 3947 2287
rect 3853 2253 3867 2267
rect 3973 2254 3987 2268
rect 4053 2333 4067 2347
rect 4033 2254 4047 2268
rect 3873 2232 3887 2246
rect 3833 2210 3847 2224
rect 3893 2213 3907 2227
rect 3873 2153 3887 2167
rect 3773 2133 3787 2147
rect 3853 2133 3867 2147
rect 3953 2212 3967 2226
rect 3993 2212 4007 2226
rect 3913 2173 3927 2187
rect 3953 2173 3967 2187
rect 4013 2173 4027 2187
rect 3933 2153 3947 2167
rect 3913 2113 3927 2127
rect 3913 1973 3927 1987
rect 3713 1912 3727 1926
rect 3713 1833 3727 1847
rect 3653 1793 3667 1807
rect 3613 1773 3627 1787
rect 3413 1553 3427 1567
rect 3433 1513 3447 1527
rect 3413 1453 3427 1467
rect 3173 1393 3187 1407
rect 3212 1393 3226 1407
rect 3153 1333 3167 1347
rect 3093 1172 3107 1186
rect 3133 1173 3147 1187
rect 2833 1153 2847 1167
rect 3013 1153 3027 1167
rect 2893 1033 2907 1047
rect 2793 1013 2807 1027
rect 2833 973 2847 987
rect 3153 1033 3167 1047
rect 3133 993 3147 1007
rect 3053 973 3067 987
rect 2893 953 2907 967
rect 2993 953 3007 967
rect 2653 872 2667 886
rect 2593 853 2607 867
rect 2633 853 2647 867
rect 2553 753 2567 767
rect 2593 694 2607 708
rect 2533 652 2547 666
rect 2413 613 2427 627
rect 2493 613 2507 627
rect 2353 533 2367 547
rect 2573 533 2587 547
rect 2353 473 2367 487
rect 2373 433 2387 447
rect 2453 433 2467 447
rect 2613 433 2627 447
rect 2213 413 2227 427
rect 2233 394 2247 408
rect 2413 394 2427 408
rect 2573 394 2587 408
rect 2093 352 2107 366
rect 2133 352 2147 366
rect 2172 352 2186 366
rect 2193 352 2207 366
rect 2253 352 2267 366
rect 2293 352 2307 366
rect 2373 353 2387 367
rect 2033 333 2047 347
rect 2073 313 2087 327
rect 1733 293 1747 307
rect 1773 293 1787 307
rect 1713 273 1727 287
rect 1633 213 1647 227
rect 1693 213 1707 227
rect 1653 193 1667 207
rect 1613 173 1627 187
rect 1513 132 1527 146
rect 1553 132 1567 146
rect 1993 273 2007 287
rect 2013 253 2027 267
rect 2113 253 2127 267
rect 1793 213 1807 227
rect 1993 213 2007 227
rect 1733 174 1747 188
rect 1713 132 1727 146
rect 1593 93 1607 107
rect 1653 93 1667 107
rect 1493 73 1507 87
rect 1753 113 1767 127
rect 1953 193 1967 207
rect 1853 174 1867 188
rect 1893 174 1907 188
rect 1933 173 1947 187
rect 1833 132 1847 146
rect 1873 132 1887 146
rect 2093 213 2107 227
rect 2053 174 2067 188
rect 1953 132 1967 146
rect 1993 132 2007 146
rect 2033 132 2047 146
rect 2073 132 2087 146
rect 2473 352 2487 366
rect 2553 352 2567 366
rect 2613 353 2627 367
rect 2593 273 2607 287
rect 2553 253 2567 267
rect 2253 233 2267 247
rect 2433 233 2447 247
rect 2213 213 2227 227
rect 2173 193 2187 207
rect 2113 132 2127 146
rect 2413 213 2427 227
rect 2453 213 2467 227
rect 2433 193 2447 207
rect 2293 174 2307 188
rect 2353 174 2367 188
rect 2473 174 2487 188
rect 2533 174 2547 188
rect 1933 93 1947 107
rect 1793 73 1807 87
rect 1713 53 1727 67
rect 2153 132 2167 146
rect 2193 132 2207 146
rect 2253 132 2267 146
rect 2313 132 2327 146
rect 2413 113 2427 127
rect 2353 93 2367 107
rect 2653 793 2667 807
rect 2753 872 2767 886
rect 2693 753 2707 767
rect 2693 732 2707 746
rect 2713 713 2727 727
rect 2693 652 2707 666
rect 2733 573 2747 587
rect 2653 553 2667 567
rect 2653 513 2667 527
rect 2753 453 2767 467
rect 2953 914 2967 928
rect 3113 953 3127 967
rect 3113 914 3127 928
rect 2933 872 2947 886
rect 3053 872 3067 886
rect 3093 872 3107 886
rect 3133 833 3147 847
rect 2973 813 2987 827
rect 3133 793 3147 807
rect 3013 733 3027 747
rect 2993 713 3007 727
rect 2973 693 2987 707
rect 2813 653 2827 667
rect 2853 652 2867 666
rect 2913 613 2927 627
rect 3093 694 3107 708
rect 3193 1333 3207 1347
rect 3233 1392 3247 1406
rect 3272 1392 3286 1406
rect 3293 1393 3307 1407
rect 3333 1433 3347 1447
rect 3373 1434 3387 1448
rect 3353 1392 3367 1406
rect 3393 1392 3407 1406
rect 3433 1393 3447 1407
rect 3313 1353 3327 1367
rect 3333 1273 3347 1287
rect 3233 1253 3247 1267
rect 3213 1233 3227 1247
rect 3193 1213 3207 1227
rect 3213 1172 3227 1186
rect 3253 1172 3267 1186
rect 3193 1153 3207 1167
rect 3253 933 3267 947
rect 3413 1233 3427 1247
rect 3353 1213 3367 1227
rect 3393 1214 3407 1228
rect 3513 1692 3527 1706
rect 3593 1692 3607 1706
rect 3553 1633 3567 1647
rect 3613 1553 3627 1567
rect 3513 1493 3527 1507
rect 3473 1434 3487 1448
rect 3553 1434 3567 1448
rect 3653 1593 3667 1607
rect 3633 1473 3647 1487
rect 3733 1493 3747 1507
rect 3693 1434 3707 1448
rect 3493 1393 3507 1407
rect 3473 1353 3487 1367
rect 3453 1273 3467 1287
rect 3613 1393 3627 1407
rect 3713 1393 3727 1407
rect 3573 1353 3587 1367
rect 3633 1353 3647 1367
rect 3673 1353 3687 1367
rect 3533 1293 3547 1307
rect 3613 1293 3627 1307
rect 3573 1253 3587 1267
rect 3493 1233 3507 1247
rect 3533 1233 3547 1247
rect 3473 1213 3487 1227
rect 3333 1193 3347 1207
rect 3413 1172 3427 1186
rect 3493 1172 3507 1186
rect 3553 1172 3567 1186
rect 3593 1172 3607 1186
rect 3633 1172 3647 1186
rect 3453 1133 3467 1147
rect 3593 1033 3607 1047
rect 3553 993 3567 1007
rect 3353 933 3367 947
rect 3313 914 3327 928
rect 3393 914 3407 928
rect 3693 1172 3707 1186
rect 3733 1153 3747 1167
rect 3693 1133 3707 1147
rect 3793 1954 3807 1968
rect 3833 1954 3847 1968
rect 3893 1954 3907 1968
rect 3773 1873 3787 1887
rect 3813 1853 3827 1867
rect 3793 1793 3807 1807
rect 3893 1873 3907 1887
rect 3853 1773 3867 1787
rect 3993 2073 4007 2087
rect 3953 1954 3967 1968
rect 4033 1913 4047 1927
rect 3973 1873 3987 1887
rect 4213 2693 4227 2707
rect 4273 2733 4287 2747
rect 4253 2673 4267 2687
rect 4173 2613 4187 2627
rect 4113 2493 4127 2507
rect 4153 2493 4167 2507
rect 4213 2474 4227 2488
rect 4273 2474 4287 2488
rect 4113 2433 4127 2447
rect 4153 2413 4167 2427
rect 4193 2353 4207 2367
rect 4313 2813 4327 2827
rect 4453 2950 4467 2964
rect 4433 2873 4447 2887
rect 4713 3772 4727 3786
rect 4813 4292 4827 4306
rect 4933 4292 4947 4306
rect 4853 4253 4867 4267
rect 4893 4253 4907 4267
rect 4953 4253 4967 4267
rect 4793 4213 4807 4227
rect 4833 4213 4847 4227
rect 4793 4173 4807 4187
rect 4793 4152 4807 4166
rect 4873 4093 4887 4107
rect 4833 4034 4847 4048
rect 4933 4153 4947 4167
rect 4933 4113 4947 4127
rect 5053 4493 5067 4507
rect 5053 4373 5067 4387
rect 5033 4353 5047 4367
rect 5093 4473 5107 4487
rect 5173 4513 5187 4527
rect 5093 4433 5107 4447
rect 5133 4433 5147 4447
rect 5073 4353 5087 4367
rect 5133 4393 5147 4407
rect 5113 4373 5127 4387
rect 5093 4334 5107 4348
rect 5013 4293 5027 4307
rect 4993 4213 5007 4227
rect 5053 4253 5067 4267
rect 5033 4233 5047 4247
rect 5053 4173 5067 4187
rect 5093 4273 5107 4287
rect 5073 4133 5087 4147
rect 5013 4113 5027 4127
rect 4973 4073 4987 4087
rect 5073 4073 5087 4087
rect 4893 4033 4907 4047
rect 4833 3973 4847 3987
rect 4793 3933 4807 3947
rect 4853 3953 4867 3967
rect 4873 3933 4887 3947
rect 4773 3633 4787 3647
rect 4793 3593 4807 3607
rect 4693 3553 4707 3567
rect 4673 3513 4687 3527
rect 4753 3516 4767 3530
rect 4633 3453 4647 3467
rect 4573 3373 4587 3387
rect 4553 3313 4567 3327
rect 4613 3313 4627 3327
rect 4573 3294 4587 3308
rect 4553 3253 4567 3267
rect 4593 3252 4607 3266
rect 4553 3213 4567 3227
rect 4633 3213 4647 3227
rect 4693 3453 4707 3467
rect 4793 3433 4807 3447
rect 4813 3393 4827 3407
rect 4913 3913 4927 3927
rect 4893 3873 4907 3887
rect 5013 3913 5027 3927
rect 5153 4333 5167 4347
rect 5213 4433 5227 4447
rect 5193 4393 5207 4407
rect 5213 4334 5227 4348
rect 5273 4812 5287 4826
rect 5313 4812 5327 4826
rect 5413 4812 5427 4826
rect 5353 4773 5367 4787
rect 5253 4733 5267 4747
rect 5373 4733 5387 4747
rect 5253 4693 5267 4707
rect 5353 4653 5367 4667
rect 5353 4593 5367 4607
rect 5313 4573 5327 4587
rect 5273 4554 5287 4568
rect 5413 4593 5427 4607
rect 5373 4553 5387 4567
rect 5453 4873 5467 4887
rect 5513 5193 5527 5207
rect 5493 5073 5507 5087
rect 5713 5753 5727 5767
rect 5793 5972 5807 5986
rect 5853 5953 5867 5967
rect 5833 5894 5847 5908
rect 5873 5853 5887 5867
rect 5853 5813 5867 5827
rect 5813 5793 5827 5807
rect 5753 5693 5767 5707
rect 5853 5693 5867 5707
rect 5713 5673 5727 5687
rect 5673 5593 5687 5607
rect 5833 5633 5847 5647
rect 6073 6253 6087 6267
rect 5933 6213 5947 6227
rect 5933 6133 5947 6147
rect 5893 5833 5907 5847
rect 5873 5633 5887 5647
rect 5753 5594 5767 5608
rect 5833 5594 5847 5608
rect 5673 5553 5687 5567
rect 5793 5553 5807 5567
rect 5733 5533 5747 5547
rect 5653 5473 5667 5487
rect 5593 5153 5607 5167
rect 5633 5413 5647 5427
rect 5693 5413 5707 5427
rect 5733 5413 5747 5427
rect 5653 5374 5667 5388
rect 5853 5552 5867 5566
rect 5953 6053 5967 6067
rect 5933 5973 5947 5987
rect 5933 5933 5947 5947
rect 5973 5993 5987 6007
rect 6033 5933 6047 5947
rect 5953 5894 5967 5908
rect 5973 5852 5987 5866
rect 6033 5853 6047 5867
rect 5953 5833 5967 5847
rect 5933 5673 5947 5687
rect 5833 5513 5847 5527
rect 5873 5513 5887 5527
rect 5813 5453 5827 5467
rect 5753 5393 5767 5407
rect 5793 5393 5807 5407
rect 5673 5293 5687 5307
rect 5733 5333 5747 5347
rect 5713 5273 5727 5287
rect 5833 5373 5847 5387
rect 5813 5332 5827 5346
rect 5853 5333 5867 5347
rect 5813 5293 5827 5307
rect 5793 5273 5807 5287
rect 5753 5253 5767 5267
rect 5773 5233 5787 5247
rect 5733 5193 5747 5207
rect 5673 5173 5687 5187
rect 5613 5113 5627 5127
rect 5533 5032 5547 5046
rect 5573 5032 5587 5046
rect 5613 5032 5627 5046
rect 5513 4854 5527 4868
rect 5593 4933 5607 4947
rect 5573 4873 5587 4887
rect 5553 4853 5567 4867
rect 5433 4573 5447 4587
rect 5493 4812 5507 4826
rect 5473 4693 5487 4707
rect 5453 4554 5467 4568
rect 5553 4813 5567 4827
rect 5553 4693 5567 4707
rect 5533 4633 5547 4647
rect 5673 5133 5687 5147
rect 5713 5074 5727 5088
rect 5693 5032 5707 5046
rect 5733 4993 5747 5007
rect 5653 4973 5667 4987
rect 5713 4973 5727 4987
rect 5633 4893 5647 4907
rect 5613 4873 5627 4887
rect 5593 4853 5607 4867
rect 5693 4953 5707 4967
rect 5753 4953 5767 4967
rect 5933 5553 5947 5567
rect 5993 5633 6007 5647
rect 6113 5953 6127 5967
rect 6093 5853 6107 5867
rect 6013 5553 6027 5567
rect 5953 5513 5967 5527
rect 5993 5473 6007 5487
rect 5953 5413 5967 5427
rect 5933 5332 5947 5346
rect 5893 5293 5907 5307
rect 5873 5233 5887 5247
rect 5853 5133 5867 5147
rect 6073 5553 6087 5567
rect 6093 5473 6107 5487
rect 6033 5433 6047 5447
rect 6093 5433 6107 5447
rect 6133 5693 6147 5707
rect 6133 5393 6147 5407
rect 6113 5373 6127 5387
rect 6133 5353 6147 5367
rect 6113 5333 6127 5347
rect 6013 5273 6027 5287
rect 6053 5273 6067 5287
rect 6053 5213 6067 5227
rect 6033 5193 6047 5207
rect 5993 5113 6007 5127
rect 6093 5113 6107 5127
rect 5893 5093 5907 5107
rect 5973 5093 5987 5107
rect 5853 5074 5867 5088
rect 6033 5074 6047 5088
rect 6073 5074 6087 5088
rect 5973 5032 5987 5046
rect 5933 5013 5947 5027
rect 5833 4993 5847 5007
rect 5873 4993 5887 5007
rect 5913 4993 5927 5007
rect 5813 4953 5827 4967
rect 5793 4933 5807 4947
rect 5713 4892 5727 4906
rect 5693 4853 5707 4867
rect 5633 4812 5647 4826
rect 5693 4813 5707 4827
rect 5633 4773 5647 4787
rect 5653 4673 5667 4687
rect 5633 4653 5647 4667
rect 5513 4613 5527 4627
rect 5573 4613 5587 4627
rect 5493 4553 5507 4567
rect 5253 4513 5267 4527
rect 5253 4473 5267 4487
rect 5273 4373 5287 4387
rect 5153 4233 5167 4247
rect 5173 4213 5187 4227
rect 5133 4093 5147 4107
rect 5173 4093 5187 4107
rect 5113 4053 5127 4067
rect 5153 4053 5167 4067
rect 5353 4513 5367 4527
rect 5333 4453 5347 4467
rect 5333 4334 5347 4348
rect 5393 4493 5407 4507
rect 5473 4513 5487 4527
rect 5373 4473 5387 4487
rect 5273 4293 5287 4307
rect 5313 4292 5327 4306
rect 5253 4273 5267 4287
rect 5313 4233 5327 4247
rect 5393 4433 5407 4447
rect 5473 4473 5487 4487
rect 5413 4334 5427 4348
rect 5453 4334 5467 4348
rect 5553 4593 5567 4607
rect 5613 4554 5627 4568
rect 5653 4613 5667 4627
rect 5533 4493 5547 4507
rect 5513 4453 5527 4467
rect 5493 4333 5507 4347
rect 5373 4193 5387 4207
rect 5473 4292 5487 4306
rect 5473 4271 5487 4285
rect 5393 4133 5407 4147
rect 5433 4133 5447 4147
rect 5213 4113 5227 4127
rect 5353 4113 5367 4127
rect 5093 3992 5107 4006
rect 5133 3992 5147 4006
rect 5113 3953 5127 3967
rect 5093 3933 5107 3947
rect 5093 3893 5107 3907
rect 5073 3873 5087 3887
rect 5013 3853 5027 3867
rect 4893 3772 4907 3786
rect 4933 3772 4947 3786
rect 4933 3751 4947 3765
rect 4893 3593 4907 3607
rect 4893 3553 4907 3567
rect 4773 3353 4787 3367
rect 4733 3333 4747 3347
rect 4833 3313 4847 3327
rect 4813 3293 4827 3307
rect 4753 3252 4767 3266
rect 4693 3213 4707 3227
rect 4773 3213 4787 3227
rect 4673 3193 4687 3207
rect 4753 3193 4767 3207
rect 4653 3073 4667 3087
rect 4633 3033 4647 3047
rect 4573 2996 4587 3010
rect 4653 2993 4667 3007
rect 4553 2953 4567 2967
rect 4653 2953 4667 2967
rect 4553 2913 4567 2927
rect 4533 2893 4547 2907
rect 4593 2853 4607 2867
rect 4533 2833 4547 2847
rect 4513 2813 4527 2827
rect 4553 2813 4567 2827
rect 4453 2773 4467 2787
rect 4513 2774 4527 2788
rect 4373 2732 4387 2746
rect 4433 2733 4447 2747
rect 4413 2693 4427 2707
rect 4333 2573 4347 2587
rect 4393 2573 4407 2587
rect 4393 2552 4407 2566
rect 4313 2533 4327 2547
rect 4393 2473 4407 2487
rect 4273 2333 4287 2347
rect 4113 2313 4127 2327
rect 4153 2313 4167 2327
rect 4193 2313 4207 2327
rect 4293 2313 4307 2327
rect 4093 2273 4107 2287
rect 4133 2212 4147 2226
rect 4093 2193 4107 2207
rect 4073 2113 4087 2127
rect 4153 2013 4167 2027
rect 4093 1973 4107 1987
rect 4173 1993 4187 2007
rect 4093 1912 4107 1926
rect 3973 1852 3987 1866
rect 4053 1853 4067 1867
rect 3833 1734 3847 1748
rect 3893 1734 3907 1748
rect 3933 1734 3947 1748
rect 4053 1832 4067 1846
rect 3993 1793 4007 1807
rect 3853 1692 3867 1706
rect 3973 1733 3987 1747
rect 3913 1693 3927 1707
rect 3813 1593 3827 1607
rect 3853 1593 3867 1607
rect 3793 1513 3807 1527
rect 3773 1434 3787 1448
rect 3813 1434 3827 1448
rect 3773 1373 3787 1387
rect 3793 1353 3807 1367
rect 3853 1353 3867 1367
rect 3913 1613 3927 1627
rect 3973 1693 3987 1707
rect 3953 1453 3967 1467
rect 3933 1434 3947 1448
rect 3973 1434 3987 1448
rect 4073 1793 4087 1807
rect 4053 1753 4067 1767
rect 4033 1734 4047 1748
rect 4133 1773 4147 1787
rect 4213 2273 4227 2287
rect 4253 2254 4267 2268
rect 4333 2432 4347 2446
rect 4373 2432 4387 2446
rect 4433 2633 4447 2647
rect 4453 2613 4467 2627
rect 4533 2732 4547 2746
rect 4573 2733 4587 2747
rect 4573 2693 4587 2707
rect 4533 2573 4547 2587
rect 4493 2553 4507 2567
rect 4453 2533 4467 2547
rect 4493 2513 4507 2527
rect 4453 2474 4467 2488
rect 4693 2950 4707 2964
rect 4673 2853 4687 2867
rect 4653 2813 4667 2827
rect 4633 2774 4647 2788
rect 4753 2853 4767 2867
rect 4793 3113 4807 3127
rect 4793 2993 4807 3007
rect 5013 3733 5027 3747
rect 5093 3814 5107 3828
rect 5373 4053 5387 4067
rect 5253 4034 5267 4048
rect 5233 3993 5247 4007
rect 5213 3913 5227 3927
rect 5273 3953 5287 3967
rect 5253 3913 5267 3927
rect 5233 3853 5247 3867
rect 5053 3773 5067 3787
rect 5033 3673 5047 3687
rect 5013 3653 5027 3667
rect 5013 3613 5027 3627
rect 5133 3733 5147 3747
rect 5073 3693 5087 3707
rect 4993 3516 5007 3530
rect 5113 3553 5127 3567
rect 5033 3513 5047 3527
rect 5012 3473 5026 3487
rect 4893 3353 4907 3367
rect 4873 3313 4887 3327
rect 4913 3313 4927 3327
rect 4973 3293 4987 3307
rect 4933 3252 4947 3266
rect 4973 3233 4987 3247
rect 4873 3173 4887 3187
rect 4953 3173 4967 3187
rect 4893 3153 4907 3167
rect 4933 3153 4947 3167
rect 4853 3093 4867 3107
rect 4873 3033 4887 3047
rect 4913 3113 4927 3127
rect 4893 3013 4907 3027
rect 4873 2996 4887 3010
rect 4893 2952 4907 2966
rect 4893 2893 4907 2907
rect 4833 2853 4847 2867
rect 4733 2833 4747 2847
rect 4773 2833 4787 2847
rect 4713 2813 4727 2827
rect 4693 2773 4707 2787
rect 4653 2732 4667 2746
rect 4693 2733 4707 2747
rect 4633 2613 4647 2627
rect 4613 2593 4627 2607
rect 4613 2533 4627 2547
rect 4633 2513 4647 2527
rect 4553 2493 4567 2507
rect 4593 2494 4607 2508
rect 4533 2453 4547 2467
rect 4353 2413 4367 2427
rect 4353 2373 4367 2387
rect 4333 2353 4347 2367
rect 4313 2253 4327 2267
rect 4273 2212 4287 2226
rect 4353 2253 4367 2267
rect 4413 2432 4427 2446
rect 4473 2432 4487 2446
rect 4473 2333 4487 2347
rect 4533 2333 4547 2347
rect 4433 2254 4447 2268
rect 4373 2153 4387 2167
rect 4333 2093 4347 2107
rect 4473 2213 4487 2227
rect 4453 2113 4467 2127
rect 4213 2073 4227 2087
rect 4413 2073 4427 2087
rect 4493 2113 4507 2127
rect 4253 1993 4267 2007
rect 4313 1993 4327 2007
rect 4247 1973 4261 1987
rect 4213 1953 4227 1967
rect 4273 1954 4287 1968
rect 4473 1992 4487 2006
rect 4333 1973 4347 1987
rect 4393 1954 4407 1968
rect 4433 1954 4447 1968
rect 4333 1933 4347 1947
rect 4253 1912 4267 1926
rect 4313 1913 4327 1927
rect 4213 1873 4227 1887
rect 4293 1873 4307 1887
rect 4193 1753 4207 1767
rect 4273 1853 4287 1867
rect 4053 1692 4067 1706
rect 4133 1692 4147 1706
rect 4033 1673 4047 1687
rect 4093 1673 4107 1687
rect 3913 1392 3927 1406
rect 3873 1333 3887 1347
rect 3953 1353 3967 1367
rect 3913 1313 3927 1327
rect 4173 1692 4187 1706
rect 4233 1673 4247 1687
rect 4153 1653 4167 1667
rect 4173 1513 4187 1527
rect 4073 1434 4087 1448
rect 4133 1434 4147 1448
rect 4033 1392 4047 1406
rect 4093 1392 4107 1406
rect 4353 1913 4367 1927
rect 4333 1893 4347 1907
rect 4313 1813 4327 1827
rect 4373 1893 4387 1907
rect 4433 1893 4447 1907
rect 4413 1853 4427 1867
rect 4353 1773 4367 1787
rect 4413 1773 4427 1787
rect 4293 1753 4307 1767
rect 4353 1734 4367 1748
rect 4353 1653 4367 1667
rect 4333 1613 4347 1627
rect 4373 1593 4387 1607
rect 4353 1573 4367 1587
rect 4293 1553 4307 1567
rect 4313 1493 4327 1507
rect 4193 1473 4207 1487
rect 4273 1473 4287 1487
rect 4173 1273 4187 1287
rect 3893 1253 3907 1267
rect 3953 1253 3967 1267
rect 4013 1253 4027 1267
rect 3813 1214 3827 1228
rect 3853 1214 3867 1228
rect 3993 1214 4007 1228
rect 4113 1253 4127 1267
rect 4053 1213 4067 1227
rect 4153 1214 4167 1228
rect 3933 1172 3947 1186
rect 3973 1172 3987 1186
rect 4033 1172 4047 1186
rect 3833 1153 3847 1167
rect 3753 1033 3767 1047
rect 3673 993 3687 1007
rect 3653 933 3667 947
rect 3713 933 3727 947
rect 3753 913 3767 927
rect 3633 893 3647 907
rect 3173 872 3187 886
rect 3273 872 3287 886
rect 3333 872 3347 886
rect 3373 872 3387 886
rect 3173 773 3187 787
rect 3233 773 3247 787
rect 3453 872 3467 886
rect 3533 872 3547 886
rect 3573 872 3587 886
rect 3693 872 3707 886
rect 3213 733 3227 747
rect 3253 733 3267 747
rect 3353 733 3367 747
rect 3413 733 3427 747
rect 3393 694 3407 708
rect 3433 693 3447 707
rect 2993 652 3007 666
rect 3033 652 3047 666
rect 2973 593 2987 607
rect 2953 573 2967 587
rect 2833 433 2847 447
rect 2853 433 2867 447
rect 2753 394 2767 408
rect 3193 652 3207 666
rect 3233 652 3247 666
rect 3273 613 3287 627
rect 3333 613 3347 627
rect 3433 633 3447 647
rect 3513 833 3527 847
rect 3553 813 3567 827
rect 3593 813 3607 827
rect 3733 813 3747 827
rect 3553 733 3567 747
rect 3633 773 3647 787
rect 3613 733 3627 747
rect 3613 693 3627 707
rect 3673 713 3687 727
rect 3733 713 3747 727
rect 3533 652 3547 666
rect 3593 653 3607 667
rect 3653 652 3667 666
rect 3693 652 3707 666
rect 3753 693 3767 707
rect 3953 1133 3967 1147
rect 3953 1073 3967 1087
rect 3833 973 3847 987
rect 3873 914 3887 928
rect 4033 953 4047 967
rect 3993 914 4007 928
rect 4133 1153 4147 1167
rect 4253 1434 4267 1448
rect 4593 2473 4607 2487
rect 4713 2633 4727 2647
rect 4813 2813 4827 2827
rect 4773 2774 4787 2788
rect 5053 3470 5067 3484
rect 5073 3393 5087 3407
rect 5033 3353 5047 3367
rect 5033 3294 5047 3308
rect 5013 3253 5027 3267
rect 4993 3213 5007 3227
rect 5033 3213 5047 3227
rect 4973 3073 4987 3087
rect 4973 3033 4987 3047
rect 5013 3033 5027 3047
rect 4953 2993 4967 3007
rect 4992 2994 5006 3008
rect 5013 2993 5027 3007
rect 4913 2813 4927 2827
rect 4833 2773 4847 2787
rect 4753 2733 4767 2747
rect 4693 2573 4707 2587
rect 4653 2432 4667 2446
rect 4693 2432 4707 2446
rect 4833 2733 4847 2747
rect 4813 2713 4827 2727
rect 4793 2693 4807 2707
rect 4813 2673 4827 2687
rect 4753 2553 4767 2567
rect 4773 2474 4787 2488
rect 4913 2730 4927 2744
rect 4853 2713 4867 2727
rect 4953 2713 4967 2727
rect 5093 3153 5107 3167
rect 5153 3713 5167 3727
rect 5153 3673 5167 3687
rect 5273 3893 5287 3907
rect 5293 3873 5307 3887
rect 5273 3833 5287 3847
rect 5253 3773 5267 3787
rect 5273 3733 5287 3747
rect 5253 3653 5267 3667
rect 5213 3613 5227 3627
rect 5253 3613 5267 3627
rect 5173 3533 5187 3547
rect 5153 3513 5167 3527
rect 5193 3513 5207 3527
rect 5273 3593 5287 3607
rect 5153 3473 5167 3487
rect 5253 3473 5267 3487
rect 5133 3393 5147 3407
rect 5133 3353 5147 3367
rect 5633 4513 5647 4527
rect 5573 4453 5587 4467
rect 5593 4413 5607 4427
rect 5633 4413 5647 4427
rect 5633 4373 5647 4387
rect 5653 4353 5667 4367
rect 5753 4873 5767 4887
rect 5873 4953 5887 4967
rect 5773 4854 5787 4868
rect 5813 4854 5827 4868
rect 5753 4813 5767 4827
rect 5833 4812 5847 4826
rect 5793 4773 5807 4787
rect 5673 4333 5687 4347
rect 5533 4292 5547 4306
rect 5573 4292 5587 4306
rect 5613 4273 5627 4287
rect 5633 4273 5647 4287
rect 5553 4233 5567 4247
rect 5593 4233 5607 4247
rect 5513 4173 5527 4187
rect 5533 4133 5547 4147
rect 5473 4093 5487 4107
rect 5533 4053 5547 4067
rect 5573 4173 5587 4187
rect 5393 4012 5407 4026
rect 5373 3813 5387 3827
rect 5313 3753 5327 3767
rect 5293 3553 5307 3567
rect 5293 3532 5307 3546
rect 5293 3472 5307 3486
rect 5273 3413 5287 3427
rect 5253 3393 5267 3407
rect 5253 3372 5267 3386
rect 5213 3333 5227 3347
rect 5153 3292 5167 3306
rect 5353 3733 5367 3747
rect 5413 3853 5427 3867
rect 5473 3853 5487 3867
rect 5533 3853 5547 3867
rect 5493 3833 5507 3847
rect 5453 3814 5467 3828
rect 5513 3814 5527 3828
rect 5613 4073 5627 4087
rect 5613 4033 5627 4047
rect 5673 4293 5687 4307
rect 5673 4233 5687 4247
rect 5653 4213 5667 4227
rect 5713 4633 5727 4647
rect 5833 4633 5847 4647
rect 5713 4573 5727 4587
rect 5713 4493 5727 4507
rect 5833 4493 5847 4507
rect 5713 4433 5727 4447
rect 5813 4433 5827 4447
rect 5713 4393 5727 4407
rect 5773 4393 5787 4407
rect 5733 4353 5747 4367
rect 5773 4334 5787 4348
rect 5713 4293 5727 4307
rect 5593 3993 5607 4007
rect 5633 3873 5647 3887
rect 5593 3853 5607 3867
rect 5413 3733 5427 3747
rect 5513 3733 5527 3747
rect 5473 3713 5487 3727
rect 5433 3533 5447 3547
rect 5393 3513 5407 3527
rect 5373 3472 5387 3486
rect 5413 3433 5427 3447
rect 5393 3413 5407 3427
rect 5333 3373 5347 3387
rect 5313 3333 5327 3347
rect 5313 3294 5327 3308
rect 5133 3193 5147 3207
rect 5053 3113 5067 3127
rect 5073 3093 5087 3107
rect 5053 3053 5067 3067
rect 5033 2933 5047 2947
rect 5073 2913 5087 2927
rect 5033 2793 5047 2807
rect 5073 2773 5087 2787
rect 5053 2733 5067 2747
rect 4913 2673 4927 2687
rect 4953 2673 4967 2687
rect 4833 2493 4847 2507
rect 4873 2493 4887 2507
rect 4953 2633 4967 2647
rect 4933 2593 4947 2607
rect 4993 2553 5007 2567
rect 4973 2533 4987 2547
rect 4833 2453 4847 2467
rect 4713 2413 4727 2427
rect 4653 2373 4667 2387
rect 4713 2333 4727 2347
rect 4573 2254 4587 2268
rect 4633 2253 4647 2267
rect 4613 2210 4627 2224
rect 4593 2153 4607 2167
rect 4613 2133 4627 2147
rect 4613 2093 4627 2107
rect 4713 2093 4727 2107
rect 4593 2073 4607 2087
rect 4553 2013 4567 2027
rect 4533 1973 4547 1987
rect 4713 2033 4727 2047
rect 4613 2013 4627 2027
rect 4593 1953 4607 1967
rect 4553 1912 4567 1926
rect 4513 1873 4527 1887
rect 4473 1853 4487 1867
rect 4473 1813 4487 1827
rect 4513 1734 4527 1748
rect 4553 1873 4567 1887
rect 4413 1673 4427 1687
rect 4493 1673 4507 1687
rect 4513 1653 4527 1667
rect 4793 2432 4807 2446
rect 4753 2413 4767 2427
rect 4813 2333 4827 2347
rect 4813 2312 4827 2326
rect 4773 2254 4787 2268
rect 4873 2273 4887 2287
rect 4833 2254 4847 2268
rect 4853 2173 4867 2187
rect 4793 2153 4807 2167
rect 4833 2133 4847 2147
rect 4753 2053 4767 2067
rect 4633 1973 4647 1987
rect 4733 1973 4747 1987
rect 4653 1953 4667 1967
rect 4693 1954 4707 1968
rect 4633 1873 4647 1887
rect 4613 1853 4627 1867
rect 4633 1813 4647 1827
rect 4593 1753 4607 1767
rect 4693 1773 4707 1787
rect 4653 1753 4667 1767
rect 4592 1692 4606 1706
rect 4613 1693 4627 1707
rect 4553 1593 4567 1607
rect 4413 1493 4427 1507
rect 4333 1453 4347 1467
rect 4393 1453 4407 1467
rect 4273 1353 4287 1367
rect 4573 1453 4587 1467
rect 4533 1434 4547 1448
rect 4593 1433 4607 1447
rect 4433 1392 4447 1406
rect 4473 1393 4487 1407
rect 4553 1392 4567 1406
rect 4493 1373 4507 1387
rect 4393 1353 4407 1367
rect 4333 1273 4347 1287
rect 4233 1233 4247 1247
rect 4213 1213 4227 1227
rect 4273 1214 4287 1228
rect 4093 1133 4107 1147
rect 4193 1133 4207 1147
rect 4213 973 4227 987
rect 4333 1113 4347 1127
rect 4393 1172 4407 1186
rect 4433 1172 4447 1186
rect 4433 1133 4447 1147
rect 4293 1073 4307 1087
rect 4353 1073 4367 1087
rect 4333 1053 4347 1067
rect 4293 1013 4307 1027
rect 4253 953 4267 967
rect 4333 953 4347 967
rect 4153 933 4167 947
rect 4053 914 4067 928
rect 4113 914 4127 928
rect 3853 872 3867 886
rect 3893 872 3907 886
rect 3953 873 3967 887
rect 4193 913 4207 927
rect 4293 913 4307 927
rect 4013 872 4027 886
rect 4052 872 4066 886
rect 4093 872 4107 886
rect 4053 813 4067 827
rect 3793 773 3807 787
rect 4013 753 4027 767
rect 3853 733 3867 747
rect 3813 694 3827 708
rect 3133 593 3147 607
rect 3373 593 3387 607
rect 3453 593 3467 607
rect 3493 593 3507 607
rect 3113 553 3127 567
rect 3373 553 3387 567
rect 3373 513 3387 527
rect 3693 513 3707 527
rect 3193 453 3207 467
rect 3273 453 3287 467
rect 3013 433 3027 447
rect 3073 433 3087 447
rect 3053 413 3067 427
rect 3153 413 3167 427
rect 3213 433 3227 447
rect 3253 413 3267 427
rect 3233 394 3247 408
rect 2793 373 2807 387
rect 2973 373 2987 387
rect 2653 353 2667 367
rect 2693 352 2707 366
rect 2733 352 2747 366
rect 2853 352 2867 366
rect 2753 333 2767 347
rect 2793 333 2807 347
rect 2713 293 2727 307
rect 2673 213 2687 227
rect 2633 193 2647 207
rect 2833 313 2847 327
rect 2813 273 2827 287
rect 2613 132 2627 146
rect 2673 132 2687 146
rect 2733 132 2747 146
rect 2533 113 2547 127
rect 2573 113 2587 127
rect 2773 113 2787 127
rect 2453 93 2467 107
rect 3033 352 3047 366
rect 3073 333 3087 347
rect 3133 333 3147 347
rect 3233 353 3247 367
rect 3213 333 3227 347
rect 3173 313 3187 327
rect 3233 313 3247 327
rect 3293 413 3307 427
rect 3473 473 3487 487
rect 3693 473 3707 487
rect 3413 394 3427 408
rect 3573 453 3587 467
rect 3533 413 3547 427
rect 3633 413 3647 427
rect 3733 652 3747 666
rect 3833 652 3847 666
rect 3993 652 4007 666
rect 3873 613 3887 627
rect 3913 613 3927 627
rect 3773 453 3787 467
rect 3813 433 3827 447
rect 3973 433 3987 447
rect 3713 413 3727 427
rect 3753 394 3767 408
rect 3853 394 3867 408
rect 3933 394 3947 408
rect 3393 352 3407 366
rect 3473 352 3487 366
rect 3313 313 3327 327
rect 3353 313 3367 327
rect 3433 313 3447 327
rect 3033 293 3047 307
rect 3253 293 3267 307
rect 2893 273 2907 287
rect 2933 193 2947 207
rect 3233 273 3247 287
rect 3273 273 3287 287
rect 3213 253 3227 267
rect 3253 253 3267 267
rect 2893 174 2907 188
rect 2973 173 2987 187
rect 3033 174 3047 188
rect 3073 174 3087 188
rect 3133 173 3147 187
rect 3513 293 3527 307
rect 3413 233 3427 247
rect 3373 213 3387 227
rect 3373 173 3387 187
rect 2833 132 2847 146
rect 2873 132 2887 146
rect 2913 132 2927 146
rect 2973 132 2987 146
rect 3153 153 3167 167
rect 3013 132 3027 146
rect 3053 132 3067 146
rect 3133 132 3147 146
rect 3633 352 3647 366
rect 3673 352 3687 366
rect 3693 333 3707 347
rect 4033 393 4047 407
rect 3653 313 3667 327
rect 3753 313 3767 327
rect 3573 293 3587 307
rect 3553 273 3567 287
rect 3533 233 3547 247
rect 3193 132 3207 146
rect 3233 132 3247 146
rect 3393 133 3407 147
rect 2993 93 3007 107
rect 3153 93 3167 107
rect 3193 73 3207 87
rect 2413 53 2427 67
rect 2813 53 2827 67
rect 3513 133 3527 147
rect 3553 213 3567 227
rect 3553 173 3567 187
rect 3613 174 3627 188
rect 3833 333 3847 347
rect 3993 352 4007 366
rect 3953 333 3967 347
rect 3933 313 3947 327
rect 3793 253 3807 267
rect 3733 213 3747 227
rect 3833 213 3847 227
rect 4093 773 4107 787
rect 4073 733 4087 747
rect 4073 652 4087 666
rect 4193 873 4207 887
rect 4273 872 4287 886
rect 4333 873 4347 887
rect 4233 853 4247 867
rect 4313 773 4327 787
rect 4253 753 4267 767
rect 4133 733 4147 747
rect 4293 713 4307 727
rect 4193 695 4207 709
rect 4113 673 4127 687
rect 4093 593 4107 607
rect 4233 653 4247 667
rect 4153 573 4167 587
rect 4113 513 4127 527
rect 4153 433 4167 447
rect 4373 973 4387 987
rect 4373 913 4387 927
rect 4513 1233 4527 1247
rect 4493 1213 4507 1227
rect 4533 1172 4547 1186
rect 4452 1113 4466 1127
rect 4473 1113 4487 1127
rect 4393 872 4407 886
rect 4453 793 4467 807
rect 4493 1013 4507 1027
rect 4553 1053 4567 1067
rect 4493 913 4507 927
rect 4673 1693 4687 1707
rect 4653 1653 4667 1667
rect 4653 1573 4667 1587
rect 4633 1473 4647 1487
rect 4733 1913 4747 1927
rect 4713 1753 4727 1767
rect 4793 1954 4807 1968
rect 4953 2393 4967 2407
rect 4913 2373 4927 2387
rect 5113 3093 5127 3107
rect 5353 3252 5367 3266
rect 5233 3213 5247 3227
rect 5273 3213 5287 3227
rect 5373 3213 5387 3227
rect 5193 3173 5207 3187
rect 5153 3073 5167 3087
rect 5113 3013 5127 3027
rect 5133 2994 5147 3008
rect 5133 2933 5147 2947
rect 5113 2913 5127 2927
rect 5153 2893 5167 2907
rect 5133 2853 5147 2867
rect 5313 3173 5327 3187
rect 5193 3013 5207 3027
rect 5273 3013 5287 3027
rect 5333 3153 5347 3167
rect 5393 3173 5407 3187
rect 5313 2994 5327 3008
rect 5353 3133 5367 3147
rect 5493 3453 5507 3467
rect 5453 3413 5467 3427
rect 5433 3393 5447 3407
rect 5453 3373 5467 3387
rect 5433 3293 5447 3307
rect 5693 3993 5707 4007
rect 5653 3833 5667 3847
rect 5573 3773 5587 3787
rect 5553 3593 5567 3607
rect 5613 3772 5627 3786
rect 5753 4273 5767 4287
rect 5893 4933 5907 4947
rect 5893 4653 5907 4667
rect 6093 5013 6107 5027
rect 6073 4993 6087 5007
rect 6013 4913 6027 4927
rect 6093 4853 6107 4867
rect 6133 5273 6147 5287
rect 6133 4893 6147 4907
rect 6053 4753 6067 4767
rect 5913 4613 5927 4627
rect 6093 4653 6107 4667
rect 6133 4573 6147 4587
rect 5893 4553 5907 4567
rect 5933 4554 5947 4568
rect 5873 4493 5887 4507
rect 5913 4512 5927 4526
rect 5893 4473 5907 4487
rect 5953 4413 5967 4427
rect 5933 4373 5947 4387
rect 5913 4353 5927 4367
rect 5873 4333 5887 4347
rect 6073 4554 6087 4568
rect 6133 4552 6147 4566
rect 6053 4512 6067 4526
rect 6113 4513 6127 4527
rect 6093 4473 6107 4487
rect 5993 4453 6007 4467
rect 6093 4452 6107 4466
rect 6013 4413 6027 4427
rect 5973 4333 5987 4347
rect 6073 4373 6087 4387
rect 5893 4293 5907 4307
rect 5813 4253 5827 4267
rect 5753 4113 5767 4127
rect 5793 4113 5807 4127
rect 5793 4092 5807 4106
rect 5753 4073 5767 4087
rect 5733 4033 5747 4047
rect 5793 4034 5807 4048
rect 5733 3993 5747 4007
rect 5713 3832 5727 3846
rect 5653 3733 5667 3747
rect 5593 3653 5607 3667
rect 5573 3573 5587 3587
rect 5533 3513 5547 3527
rect 5553 3533 5567 3547
rect 5533 3473 5547 3487
rect 5513 3393 5527 3407
rect 5493 3314 5507 3328
rect 5573 3472 5587 3486
rect 5593 3453 5607 3467
rect 5553 3393 5567 3407
rect 5493 3293 5507 3307
rect 5473 3252 5487 3266
rect 5513 3252 5527 3266
rect 5433 3173 5447 3187
rect 5413 3073 5427 3087
rect 5393 3033 5407 3047
rect 5233 2952 5247 2966
rect 5193 2873 5207 2887
rect 5173 2833 5187 2847
rect 5173 2812 5187 2826
rect 5153 2793 5167 2807
rect 5233 2873 5247 2887
rect 5153 2732 5167 2746
rect 5093 2712 5107 2726
rect 5073 2593 5087 2607
rect 4993 2473 5007 2487
rect 5053 2493 5067 2507
rect 5073 2474 5087 2488
rect 4993 2433 5007 2447
rect 4973 2353 4987 2367
rect 4993 2333 5007 2347
rect 4973 2273 4987 2287
rect 4933 2093 4947 2107
rect 4873 2013 4887 2027
rect 4813 1912 4827 1926
rect 4833 1893 4847 1907
rect 4773 1833 4787 1847
rect 4753 1753 4767 1767
rect 5053 2432 5067 2446
rect 5093 2433 5107 2447
rect 5073 2393 5087 2407
rect 5053 2333 5067 2347
rect 5013 2273 5027 2287
rect 5193 2693 5207 2707
rect 5373 2993 5387 3007
rect 5313 2853 5327 2867
rect 5253 2813 5267 2827
rect 5253 2773 5267 2787
rect 5293 2774 5307 2788
rect 5353 2952 5367 2966
rect 5413 2953 5427 2967
rect 5413 2893 5427 2907
rect 5353 2873 5367 2887
rect 5393 2853 5407 2867
rect 5353 2772 5367 2786
rect 5133 2613 5147 2627
rect 5233 2613 5247 2627
rect 5313 2732 5327 2746
rect 5213 2553 5227 2567
rect 5173 2513 5187 2527
rect 5133 2473 5147 2487
rect 5113 2373 5127 2387
rect 5113 2333 5127 2347
rect 5093 2313 5107 2327
rect 5073 2273 5087 2287
rect 5033 2212 5047 2226
rect 5153 2432 5167 2446
rect 5153 2313 5167 2327
rect 5353 2693 5367 2707
rect 5333 2553 5347 2567
rect 5373 2553 5387 2567
rect 5253 2533 5267 2547
rect 5293 2474 5307 2488
rect 5333 2474 5347 2488
rect 5373 2473 5387 2487
rect 5273 2433 5287 2447
rect 5253 2413 5267 2427
rect 5253 2373 5267 2387
rect 5213 2273 5227 2287
rect 5093 2233 5107 2247
rect 5033 2173 5047 2187
rect 4893 1973 4907 1987
rect 4973 1973 4987 1987
rect 5013 1973 5027 1987
rect 4873 1813 4887 1827
rect 4933 1954 4947 1968
rect 4953 1913 4967 1927
rect 4933 1893 4947 1907
rect 4853 1753 4867 1767
rect 4833 1733 4847 1747
rect 4793 1692 4807 1706
rect 4833 1693 4847 1707
rect 4833 1553 4847 1567
rect 4753 1513 4767 1527
rect 4893 1493 4907 1507
rect 4693 1473 4707 1487
rect 4773 1433 4787 1447
rect 4633 1392 4647 1406
rect 4673 1392 4687 1406
rect 4613 1353 4627 1367
rect 4673 1333 4687 1347
rect 4713 1293 4727 1307
rect 4853 1434 4867 1448
rect 4973 1813 4987 1827
rect 5013 1813 5027 1827
rect 5133 2193 5147 2207
rect 5113 2093 5127 2107
rect 5073 2053 5087 2067
rect 5173 1993 5187 2007
rect 5093 1973 5107 1987
rect 5073 1953 5087 1967
rect 5193 1954 5207 1968
rect 5113 1912 5127 1926
rect 5053 1893 5067 1907
rect 5093 1893 5107 1907
rect 5213 1913 5227 1927
rect 5073 1833 5087 1847
rect 4973 1773 4987 1787
rect 4953 1733 4967 1747
rect 5053 1733 5067 1747
rect 4933 1673 4947 1687
rect 4913 1453 4927 1467
rect 5053 1693 5067 1707
rect 5033 1673 5047 1687
rect 4973 1633 4987 1647
rect 4953 1513 4967 1527
rect 5033 1513 5047 1527
rect 4953 1492 4967 1506
rect 4933 1433 4947 1447
rect 4793 1393 4807 1407
rect 4873 1392 4887 1406
rect 4933 1393 4947 1407
rect 4913 1353 4927 1367
rect 4793 1333 4807 1347
rect 4673 1214 4687 1228
rect 4713 1216 4727 1230
rect 4773 1216 4787 1230
rect 4813 1293 4827 1307
rect 4813 1213 4827 1227
rect 4813 1173 4827 1187
rect 4973 1453 4987 1467
rect 4953 1373 4967 1387
rect 4953 1333 4967 1347
rect 4893 1170 4907 1184
rect 4793 1133 4807 1147
rect 4672 1113 4686 1127
rect 4693 1113 4707 1127
rect 4633 1093 4647 1107
rect 4593 1033 4607 1047
rect 4613 993 4627 1007
rect 4533 872 4547 886
rect 4573 872 4587 886
rect 4693 1073 4707 1087
rect 4753 1073 4767 1087
rect 4673 953 4687 967
rect 4713 953 4727 967
rect 4633 914 4647 928
rect 4673 914 4687 928
rect 4833 993 4847 1007
rect 4773 973 4787 987
rect 4633 873 4647 887
rect 4693 872 4707 886
rect 4753 873 4767 887
rect 4873 914 4887 928
rect 4633 833 4647 847
rect 4773 833 4787 847
rect 4813 833 4827 847
rect 4613 813 4627 827
rect 4573 773 4587 787
rect 4473 733 4487 747
rect 4573 733 4587 747
rect 4353 713 4367 727
rect 4393 694 4407 708
rect 4453 693 4467 707
rect 4493 694 4507 708
rect 4313 652 4327 666
rect 4413 652 4427 666
rect 4473 653 4487 667
rect 4453 613 4467 627
rect 4513 633 4527 647
rect 4473 573 4487 587
rect 4733 793 4747 807
rect 4693 713 4707 727
rect 4653 633 4667 647
rect 4613 613 4627 627
rect 4593 593 4607 607
rect 4593 553 4607 567
rect 4573 533 4587 547
rect 4373 513 4387 527
rect 4493 493 4507 507
rect 4313 473 4327 487
rect 4113 394 4127 408
rect 4213 394 4227 408
rect 4253 394 4267 408
rect 4293 394 4307 408
rect 4053 313 4067 327
rect 4193 352 4207 366
rect 4233 352 4247 366
rect 4093 253 4107 267
rect 4033 213 4047 227
rect 3653 173 3667 187
rect 3773 174 3787 188
rect 3693 153 3707 167
rect 3633 132 3647 146
rect 3533 113 3547 127
rect 3593 113 3607 127
rect 3693 93 3707 107
rect 3793 132 3807 146
rect 4133 193 4147 207
rect 4093 174 4107 188
rect 4153 174 4167 188
rect 4213 174 4227 188
rect 4253 174 4267 188
rect 4033 132 4047 146
rect 4073 132 4087 146
rect 4193 132 4207 146
rect 4233 132 4247 146
rect 4113 93 4127 107
rect 4153 93 4167 107
rect 4213 93 4227 107
rect 4073 73 4087 87
rect 4353 453 4367 467
rect 4393 413 4407 427
rect 4433 394 4447 408
rect 4313 353 4327 367
rect 4533 394 4547 408
rect 4813 773 4827 787
rect 4773 713 4787 727
rect 4953 1153 4967 1167
rect 4953 1053 4967 1067
rect 4953 993 4967 1007
rect 4933 973 4947 987
rect 4953 953 4967 967
rect 5073 1633 5087 1647
rect 5053 1453 5067 1467
rect 5013 1373 5027 1387
rect 5073 1393 5087 1407
rect 5053 1353 5067 1367
rect 5053 1213 5067 1227
rect 5013 1172 5027 1186
rect 4993 1053 5007 1067
rect 4973 933 4987 947
rect 5173 1853 5187 1867
rect 5113 1793 5127 1807
rect 5193 1833 5207 1847
rect 5253 2333 5267 2347
rect 5353 2432 5367 2446
rect 5513 3053 5527 3067
rect 5453 3033 5467 3047
rect 5433 2813 5447 2827
rect 5473 2993 5487 3007
rect 5573 3353 5587 3367
rect 5653 3433 5667 3447
rect 5633 3353 5647 3367
rect 5613 3333 5627 3347
rect 5573 3293 5587 3307
rect 5653 3294 5667 3308
rect 5573 3253 5587 3267
rect 5553 3173 5567 3187
rect 5633 3213 5647 3227
rect 5813 3993 5827 4007
rect 5773 3953 5787 3967
rect 5793 3873 5807 3887
rect 5773 3853 5787 3867
rect 5733 3813 5747 3827
rect 5873 4273 5887 4287
rect 5853 4253 5867 4267
rect 5833 3933 5847 3947
rect 5833 3853 5847 3867
rect 5793 3772 5807 3786
rect 5773 3753 5787 3767
rect 5733 3613 5747 3627
rect 5713 3593 5727 3607
rect 5793 3573 5807 3587
rect 5693 3513 5707 3527
rect 5733 3514 5747 3528
rect 5773 3514 5787 3528
rect 5813 3513 5827 3527
rect 5693 3473 5707 3487
rect 5753 3472 5767 3486
rect 5793 3472 5807 3486
rect 5713 3413 5727 3427
rect 5773 3413 5787 3427
rect 5713 3373 5727 3387
rect 5753 3373 5767 3387
rect 5713 3333 5727 3347
rect 5753 3313 5767 3327
rect 5733 3294 5747 3308
rect 5793 3293 5807 3307
rect 5693 3233 5707 3247
rect 5593 3193 5607 3207
rect 5573 3133 5587 3147
rect 5553 3093 5567 3107
rect 5573 3073 5587 3087
rect 5553 3053 5567 3067
rect 5533 2993 5547 3007
rect 5613 2993 5627 3007
rect 5553 2952 5567 2966
rect 5593 2933 5607 2947
rect 5653 3173 5667 3187
rect 5793 3253 5807 3267
rect 5773 3233 5787 3247
rect 5753 3153 5767 3167
rect 5753 3093 5767 3107
rect 5693 2994 5707 3008
rect 5633 2953 5647 2967
rect 5533 2873 5547 2887
rect 5613 2873 5627 2887
rect 5713 2952 5727 2966
rect 5473 2833 5487 2847
rect 5553 2833 5567 2847
rect 5613 2833 5627 2847
rect 5453 2793 5467 2807
rect 5473 2774 5487 2788
rect 5553 2792 5567 2806
rect 5613 2793 5627 2807
rect 5413 2733 5427 2747
rect 5493 2732 5507 2746
rect 5453 2633 5467 2647
rect 5553 2732 5567 2746
rect 5633 2733 5647 2747
rect 5593 2713 5607 2727
rect 5593 2653 5607 2667
rect 5433 2533 5447 2547
rect 5413 2473 5427 2487
rect 5493 2493 5507 2507
rect 5533 2553 5547 2567
rect 5513 2473 5527 2487
rect 5553 2493 5567 2507
rect 5312 2413 5326 2427
rect 5333 2413 5347 2427
rect 5293 2353 5307 2367
rect 5273 2313 5287 2327
rect 5353 2333 5367 2347
rect 5333 2253 5347 2267
rect 5273 2173 5287 2187
rect 5253 2073 5267 2087
rect 5233 1773 5247 1787
rect 5153 1653 5167 1667
rect 5173 1553 5187 1567
rect 5133 1513 5147 1527
rect 5113 1473 5127 1487
rect 5213 1693 5227 1707
rect 5193 1533 5207 1547
rect 5193 1473 5207 1487
rect 5173 1434 5187 1448
rect 5113 1393 5127 1407
rect 5153 1253 5167 1267
rect 5293 2053 5307 2067
rect 5333 2213 5347 2227
rect 5452 2432 5466 2446
rect 5473 2433 5487 2447
rect 5533 2433 5547 2447
rect 5913 4273 5927 4287
rect 5893 4153 5907 4167
rect 5973 4293 5987 4307
rect 5953 4233 5967 4247
rect 5953 4113 5967 4127
rect 5913 4033 5927 4047
rect 5973 4033 5987 4047
rect 5873 3993 5887 4007
rect 5873 3953 5887 3967
rect 5933 3953 5947 3967
rect 5973 3933 5987 3947
rect 5893 3853 5907 3867
rect 5933 3853 5947 3867
rect 5853 3833 5867 3847
rect 5893 3814 5907 3828
rect 5953 3813 5967 3827
rect 5853 3733 5867 3747
rect 5913 3733 5927 3747
rect 5873 3653 5887 3667
rect 5853 3613 5867 3627
rect 5833 3413 5847 3427
rect 5933 3593 5947 3607
rect 5893 3553 5907 3567
rect 5873 3513 5887 3527
rect 5953 3513 5967 3527
rect 5873 3473 5887 3487
rect 5853 3373 5867 3387
rect 5933 3453 5947 3467
rect 5913 3433 5927 3447
rect 5833 3333 5847 3347
rect 5873 3333 5887 3347
rect 5813 3233 5827 3247
rect 5793 3173 5807 3187
rect 5793 3053 5807 3067
rect 5773 2993 5787 3007
rect 5893 3313 5907 3327
rect 5932 3313 5946 3327
rect 5953 3313 5967 3327
rect 5873 3233 5887 3247
rect 5893 3213 5907 3227
rect 5873 3173 5887 3187
rect 5853 3113 5867 3127
rect 5833 2993 5847 3007
rect 5773 2953 5787 2967
rect 5753 2893 5767 2907
rect 5713 2833 5727 2847
rect 5833 2953 5847 2967
rect 5953 3253 5967 3267
rect 5933 3233 5947 3247
rect 5913 3193 5927 3207
rect 5893 3113 5907 3127
rect 5893 3092 5907 3106
rect 5873 3033 5887 3047
rect 5933 3053 5947 3067
rect 5913 3013 5927 3027
rect 5953 2993 5967 3007
rect 5893 2933 5907 2947
rect 5853 2913 5867 2927
rect 5873 2853 5887 2867
rect 5793 2813 5807 2827
rect 5833 2813 5847 2827
rect 5773 2793 5787 2807
rect 5953 2953 5967 2967
rect 5933 2913 5947 2927
rect 5913 2853 5927 2867
rect 5853 2774 5867 2788
rect 5893 2773 5907 2787
rect 5653 2653 5667 2667
rect 5633 2493 5647 2507
rect 5693 2713 5707 2727
rect 5753 2573 5767 2587
rect 5693 2493 5707 2507
rect 5613 2432 5627 2446
rect 5553 2413 5567 2427
rect 5593 2413 5607 2427
rect 5493 2353 5507 2367
rect 5473 2333 5487 2347
rect 5673 2433 5687 2447
rect 5653 2393 5667 2407
rect 5593 2333 5607 2347
rect 5653 2333 5667 2347
rect 5433 2254 5447 2268
rect 5573 2313 5587 2327
rect 5573 2273 5587 2287
rect 5513 2254 5527 2268
rect 5553 2254 5567 2268
rect 5593 2254 5607 2268
rect 5453 2212 5467 2226
rect 5373 2173 5387 2187
rect 5373 2093 5387 2107
rect 5353 2073 5367 2087
rect 5272 1953 5286 1967
rect 5293 1954 5307 1968
rect 5333 1954 5347 1968
rect 5573 2212 5587 2226
rect 5593 2193 5607 2207
rect 5513 2173 5527 2187
rect 5433 2153 5447 2167
rect 5413 2113 5427 2127
rect 5393 2053 5407 2067
rect 5393 1993 5407 2007
rect 5353 1912 5367 1926
rect 5273 1893 5287 1907
rect 5373 1833 5387 1847
rect 5313 1793 5327 1807
rect 5573 2093 5587 2107
rect 5573 2053 5587 2067
rect 5453 2013 5467 2027
rect 5433 1953 5447 1967
rect 5533 1973 5547 1987
rect 5493 1954 5507 1968
rect 5553 1953 5567 1967
rect 5412 1913 5426 1927
rect 5593 1973 5607 1987
rect 5653 2153 5667 2167
rect 5733 2493 5747 2507
rect 5813 2733 5827 2747
rect 5773 2533 5787 2547
rect 5873 2732 5887 2746
rect 5813 2633 5827 2647
rect 5913 2613 5927 2627
rect 5873 2593 5887 2607
rect 5833 2553 5847 2567
rect 5713 2473 5727 2487
rect 5793 2493 5807 2507
rect 5693 2413 5707 2427
rect 5733 2413 5747 2427
rect 5713 2393 5727 2407
rect 5793 2432 5807 2446
rect 5853 2493 5867 2507
rect 5773 2253 5787 2267
rect 5833 2432 5847 2446
rect 5833 2393 5847 2407
rect 5913 2573 5927 2587
rect 5953 2853 5967 2867
rect 5953 2793 5967 2807
rect 6033 4233 6047 4247
rect 6033 4113 6047 4127
rect 6013 4033 6027 4047
rect 6113 4413 6127 4427
rect 6093 4073 6107 4087
rect 6073 4033 6087 4047
rect 6133 4053 6147 4067
rect 6053 3992 6067 4006
rect 6033 3973 6047 3987
rect 6013 3873 6027 3887
rect 6053 3913 6067 3927
rect 6093 3913 6107 3927
rect 5993 3813 6007 3827
rect 6033 3833 6047 3847
rect 6073 3873 6087 3887
rect 6053 3813 6067 3827
rect 6013 3673 6027 3687
rect 6053 3773 6067 3787
rect 6033 3633 6047 3647
rect 6093 3833 6107 3847
rect 6133 3953 6147 3967
rect 6133 3913 6147 3927
rect 6113 3673 6127 3687
rect 6093 3653 6107 3667
rect 6113 3633 6127 3647
rect 6093 3593 6107 3607
rect 6073 3553 6087 3567
rect 6033 3533 6047 3547
rect 5993 3513 6007 3527
rect 6113 3513 6127 3527
rect 6013 3373 6027 3387
rect 6073 3472 6087 3486
rect 6053 3333 6067 3347
rect 6113 3333 6127 3347
rect 6033 3313 6047 3327
rect 6013 3293 6027 3307
rect 6013 3253 6027 3267
rect 5993 3213 6007 3227
rect 5993 3153 6007 3167
rect 6033 3233 6047 3247
rect 6093 3233 6107 3247
rect 6073 3153 6087 3167
rect 6033 3053 6047 3067
rect 6053 3033 6067 3047
rect 6013 2993 6027 3007
rect 6113 3193 6127 3207
rect 6113 3153 6127 3167
rect 6093 3013 6107 3027
rect 6133 3053 6147 3067
rect 6133 3013 6147 3027
rect 6013 2953 6027 2967
rect 5993 2933 6007 2947
rect 6073 2952 6087 2966
rect 6133 2952 6147 2966
rect 6093 2933 6107 2947
rect 6033 2893 6047 2907
rect 6013 2813 6027 2827
rect 6053 2813 6067 2827
rect 5993 2793 6007 2807
rect 5933 2493 5947 2507
rect 6013 2732 6027 2746
rect 6013 2653 6027 2667
rect 6013 2613 6027 2627
rect 5993 2573 6007 2587
rect 6073 2653 6087 2667
rect 6053 2573 6067 2587
rect 6053 2533 6067 2547
rect 5993 2473 6007 2487
rect 6073 2473 6087 2487
rect 5873 2433 5887 2447
rect 5853 2313 5867 2327
rect 5933 2432 5947 2446
rect 5973 2433 5987 2447
rect 5993 2433 6007 2447
rect 5893 2393 5907 2407
rect 5973 2353 5987 2367
rect 5913 2313 5927 2327
rect 5953 2313 5967 2327
rect 5733 2173 5747 2187
rect 5773 2113 5787 2127
rect 5673 2053 5687 2067
rect 5773 2013 5787 2027
rect 5633 1993 5647 2007
rect 5673 1993 5687 2007
rect 5653 1954 5667 1968
rect 5733 1954 5747 1968
rect 5593 1933 5607 1947
rect 5433 1912 5447 1926
rect 5473 1912 5487 1926
rect 5513 1912 5527 1926
rect 5573 1912 5587 1926
rect 5253 1733 5267 1747
rect 5313 1753 5327 1767
rect 5393 1752 5407 1766
rect 5453 1893 5467 1907
rect 5613 1913 5627 1927
rect 5473 1873 5487 1887
rect 5592 1873 5606 1887
rect 5453 1853 5467 1867
rect 5433 1733 5447 1747
rect 5233 1593 5247 1607
rect 5293 1653 5307 1667
rect 5273 1613 5287 1627
rect 5273 1533 5287 1547
rect 5313 1533 5327 1547
rect 5232 1433 5246 1447
rect 5253 1433 5267 1447
rect 5133 1173 5147 1187
rect 5113 1073 5127 1087
rect 5093 993 5107 1007
rect 5052 932 5066 946
rect 5073 933 5087 947
rect 4993 914 5007 928
rect 5033 913 5047 927
rect 4973 872 4987 886
rect 5033 872 5047 886
rect 5033 833 5047 847
rect 4973 713 4987 727
rect 4852 693 4866 707
rect 4873 694 4887 708
rect 4933 694 4947 708
rect 4833 652 4847 666
rect 4813 633 4827 647
rect 4733 573 4747 587
rect 4713 413 4727 427
rect 4773 396 4787 410
rect 4413 333 4427 347
rect 4373 313 4387 327
rect 4353 253 4367 267
rect 4313 173 4327 187
rect 4393 174 4407 188
rect 4433 174 4447 188
rect 4373 132 4387 146
rect 4313 113 4327 127
rect 4413 113 4427 127
rect 4553 352 4567 366
rect 4593 350 4607 364
rect 5033 693 5047 707
rect 4873 633 4887 647
rect 4853 396 4867 410
rect 4813 333 4827 347
rect 4673 313 4687 327
rect 4833 213 4847 227
rect 4553 174 4567 188
rect 4633 174 4647 188
rect 4493 132 4507 146
rect 4913 253 4927 267
rect 4973 613 4987 627
rect 4993 573 5007 587
rect 5013 553 5027 567
rect 4973 473 4987 487
rect 5153 1073 5167 1087
rect 5153 973 5167 987
rect 5112 933 5126 947
rect 5133 933 5147 947
rect 5073 912 5087 926
rect 5293 1353 5307 1367
rect 5312 1214 5326 1228
rect 5373 1693 5387 1707
rect 5353 1673 5367 1687
rect 5373 1493 5387 1507
rect 5353 1433 5367 1447
rect 5433 1533 5447 1547
rect 5413 1493 5427 1507
rect 5613 1872 5627 1886
rect 5673 1912 5687 1926
rect 5713 1873 5727 1887
rect 5813 2213 5827 2227
rect 5793 1973 5807 1987
rect 5853 2093 5867 2107
rect 5853 1973 5867 1987
rect 5873 1953 5887 1967
rect 5753 1913 5767 1927
rect 5793 1893 5807 1907
rect 5733 1853 5747 1867
rect 5633 1833 5647 1847
rect 5693 1833 5707 1847
rect 5633 1793 5647 1807
rect 5493 1773 5507 1787
rect 5613 1773 5627 1787
rect 5513 1734 5527 1748
rect 5553 1734 5567 1748
rect 5593 1734 5607 1748
rect 5653 1714 5667 1728
rect 5473 1673 5487 1687
rect 5473 1613 5487 1627
rect 5453 1473 5467 1487
rect 5573 1673 5587 1687
rect 5671 1673 5685 1687
rect 5533 1633 5547 1647
rect 5393 1453 5407 1467
rect 5493 1453 5507 1467
rect 5413 1434 5427 1448
rect 5873 1893 5887 1907
rect 5853 1873 5867 1887
rect 5913 2253 5927 2267
rect 6013 2393 6027 2407
rect 6073 2433 6087 2447
rect 6053 2393 6067 2407
rect 6033 2373 6047 2387
rect 6013 2313 6027 2327
rect 5993 2273 6007 2287
rect 6013 2253 6027 2267
rect 5913 2213 5927 2227
rect 5933 2053 5947 2067
rect 5953 2013 5967 2027
rect 5913 1953 5927 1967
rect 6013 2213 6027 2227
rect 6053 2313 6067 2327
rect 6053 2273 6067 2287
rect 6033 2013 6047 2027
rect 5933 1912 5947 1926
rect 5973 1873 5987 1887
rect 5913 1833 5927 1847
rect 5953 1833 5967 1847
rect 5813 1813 5827 1827
rect 5853 1813 5867 1827
rect 5893 1813 5907 1827
rect 5973 1813 5987 1827
rect 5713 1753 5727 1767
rect 5973 1733 5987 1747
rect 5853 1712 5867 1726
rect 5953 1713 5967 1727
rect 5993 1713 6007 1727
rect 6113 2913 6127 2927
rect 6093 2393 6107 2407
rect 6093 2353 6107 2367
rect 6073 1912 6087 1926
rect 5713 1673 5727 1687
rect 5973 1653 5987 1667
rect 5693 1633 5707 1647
rect 5713 1573 5727 1587
rect 5713 1513 5727 1527
rect 5593 1453 5607 1467
rect 5953 1513 5967 1527
rect 5933 1473 5947 1487
rect 5473 1412 5487 1426
rect 5533 1412 5547 1426
rect 5573 1412 5587 1426
rect 5333 1213 5347 1227
rect 5253 1153 5267 1167
rect 5307 1153 5321 1167
rect 5273 1133 5287 1147
rect 5213 1033 5227 1047
rect 5193 953 5207 967
rect 5173 872 5187 886
rect 5393 1392 5407 1406
rect 5413 1253 5427 1267
rect 5493 1393 5507 1407
rect 5473 1353 5487 1367
rect 5473 1273 5487 1287
rect 5373 1213 5387 1227
rect 5453 1213 5467 1227
rect 5373 1173 5387 1187
rect 5433 1172 5447 1186
rect 5473 1173 5487 1187
rect 5293 1113 5307 1127
rect 5353 1113 5367 1127
rect 5533 1373 5547 1387
rect 5553 1353 5567 1367
rect 5533 1293 5547 1307
rect 5733 1414 5747 1428
rect 5853 1412 5867 1426
rect 5593 1373 5607 1387
rect 5573 1313 5587 1327
rect 5673 1313 5687 1327
rect 5713 1313 5727 1327
rect 5553 1273 5567 1287
rect 5513 1214 5527 1228
rect 5553 1214 5567 1228
rect 5693 1293 5707 1307
rect 5693 1213 5707 1227
rect 5953 1333 5967 1347
rect 6033 1673 6047 1687
rect 6073 1513 6087 1527
rect 6053 1473 6067 1487
rect 6013 1434 6027 1448
rect 6033 1392 6047 1406
rect 5973 1313 5987 1327
rect 5853 1293 5867 1307
rect 6013 1333 6027 1347
rect 5613 1194 5627 1208
rect 5673 1194 5687 1208
rect 5713 1194 5727 1208
rect 5533 1172 5547 1186
rect 5513 1153 5527 1167
rect 5993 1213 6007 1227
rect 6053 1213 6067 1227
rect 6133 2853 6147 2867
rect 6133 2593 6147 2607
rect 6133 2533 6147 2547
rect 6133 2353 6147 2367
rect 6113 2313 6127 2327
rect 6093 1273 6107 1287
rect 5873 1192 5887 1206
rect 5973 1193 5987 1207
rect 6013 1193 6027 1207
rect 5513 1113 5527 1127
rect 5453 1033 5467 1047
rect 5493 1033 5507 1047
rect 5393 993 5407 1007
rect 5433 993 5447 1007
rect 5493 993 5507 1007
rect 5293 953 5307 967
rect 5333 953 5347 967
rect 5293 914 5307 928
rect 5353 933 5367 947
rect 5333 913 5347 927
rect 5473 893 5487 907
rect 5213 872 5227 886
rect 5273 872 5287 886
rect 5093 793 5107 807
rect 5233 793 5247 807
rect 5073 733 5087 747
rect 5133 733 5147 747
rect 5093 713 5107 727
rect 5273 773 5287 787
rect 5273 733 5287 747
rect 5353 873 5367 887
rect 5413 872 5427 886
rect 5453 853 5467 867
rect 5273 694 5287 708
rect 5313 694 5327 708
rect 5393 694 5407 708
rect 5433 694 5447 708
rect 5473 694 5487 708
rect 5113 652 5127 666
rect 5053 633 5067 647
rect 5053 433 5067 447
rect 5033 413 5047 427
rect 5093 394 5107 408
rect 5253 652 5267 666
rect 5213 613 5227 627
rect 5373 633 5387 647
rect 5253 593 5267 607
rect 5453 573 5467 587
rect 5593 1093 5607 1107
rect 5553 933 5567 947
rect 5733 1153 5747 1167
rect 6093 1153 6107 1167
rect 5713 1133 5727 1147
rect 6009 1133 6023 1147
rect 6053 1113 6067 1127
rect 5853 1073 5867 1087
rect 5933 1073 5947 1087
rect 5713 993 5727 1007
rect 5813 993 5827 1007
rect 5853 993 5867 1007
rect 5713 953 5727 967
rect 5513 793 5527 807
rect 5613 853 5627 867
rect 5552 733 5566 747
rect 5573 733 5587 747
rect 5633 753 5647 767
rect 5613 733 5627 747
rect 5693 913 5707 927
rect 5733 853 5747 867
rect 5713 753 5727 767
rect 5613 693 5627 707
rect 5533 652 5547 666
rect 5573 593 5587 607
rect 5493 553 5507 567
rect 5153 493 5167 507
rect 5373 493 5387 507
rect 5413 493 5427 507
rect 5653 713 5667 727
rect 5753 713 5767 727
rect 5673 653 5687 667
rect 5653 593 5667 607
rect 5713 553 5727 567
rect 5693 533 5707 547
rect 5153 433 5167 447
rect 5033 352 5047 366
rect 5073 333 5087 347
rect 5133 333 5147 347
rect 5193 394 5207 408
rect 5593 473 5607 487
rect 5553 453 5567 467
rect 5433 413 5447 427
rect 5493 413 5507 427
rect 5613 413 5627 427
rect 5693 393 5707 407
rect 5593 373 5607 387
rect 5013 253 5027 267
rect 5153 253 5167 267
rect 5193 253 5207 267
rect 4953 213 4967 227
rect 4913 176 4927 190
rect 5013 174 5027 188
rect 5253 350 5267 364
rect 5213 213 5227 227
rect 5373 213 5387 227
rect 5293 176 5307 190
rect 5673 350 5687 364
rect 5373 174 5387 188
rect 5513 174 5527 188
rect 5593 174 5607 188
rect 5773 633 5787 647
rect 5773 533 5787 547
rect 5733 453 5747 467
rect 5773 493 5787 507
rect 5793 473 5807 487
rect 5853 953 5867 967
rect 5913 793 5927 807
rect 5873 573 5887 587
rect 6033 1033 6047 1047
rect 5993 993 6007 1007
rect 5993 914 6007 928
rect 5973 694 5987 708
rect 5993 633 6007 647
rect 5933 533 5947 547
rect 6013 493 6027 507
rect 5933 433 5947 447
rect 5813 413 5827 427
rect 5873 413 5887 427
rect 5773 352 5787 366
rect 5713 293 5727 307
rect 5773 293 5787 307
rect 5813 293 5827 307
rect 5973 394 5987 408
rect 5873 352 5887 366
rect 5913 352 5927 366
rect 5953 313 5967 327
rect 6033 352 6047 366
rect 6013 313 6027 327
rect 6073 433 6087 447
rect 5973 273 5987 287
rect 6053 273 6067 287
rect 4433 93 4447 107
rect 4013 53 4027 67
rect 4293 53 4307 67
rect 4533 53 4547 67
rect 753 33 767 47
rect 1333 33 1347 47
rect 2133 33 2147 47
rect 2773 33 2787 47
rect 2853 33 2867 47
rect 3393 33 3407 47
rect 3453 33 3467 47
rect 3753 33 3767 47
rect 4733 130 4747 144
rect 4793 130 4807 144
rect 4832 130 4846 144
rect 4853 130 4867 144
rect 5113 130 5127 144
rect 5173 130 5187 144
rect 5213 130 5227 144
rect 5853 132 5867 146
rect 5933 132 5947 146
rect 6133 1113 6147 1127
rect 6133 1073 6147 1087
rect 6113 493 6127 507
rect 6093 394 6107 408
rect 6133 293 6147 307
<< metal3 >>
rect 3347 6256 3873 6264
rect 4867 6256 5193 6264
rect 5867 6256 6073 6264
rect 3547 6236 3853 6244
rect 3867 6236 4373 6244
rect 4447 6236 4964 6244
rect 307 6216 653 6224
rect 667 6216 913 6224
rect 4367 6216 4933 6224
rect 4956 6224 4964 6236
rect 5087 6236 5113 6244
rect 5136 6236 5653 6244
rect 5136 6224 5144 6236
rect 4956 6216 5144 6224
rect 5907 6216 5933 6224
rect 767 6196 1433 6204
rect 1447 6196 1993 6204
rect 2007 6196 2073 6204
rect 2247 6196 2384 6204
rect 2376 6187 2384 6196
rect 3207 6196 3253 6204
rect 3267 6196 3533 6204
rect 4387 6196 4953 6204
rect 4967 6196 5333 6204
rect 527 6176 733 6184
rect 2047 6176 2253 6184
rect 2387 6176 2473 6184
rect 3107 6176 3373 6184
rect 5627 6176 5833 6184
rect 107 6156 253 6164
rect 267 6156 393 6164
rect 887 6156 1093 6164
rect 1207 6156 1373 6164
rect 1667 6156 1773 6164
rect 1787 6156 1873 6164
rect 2787 6156 2853 6164
rect 3727 6156 3813 6164
rect 3907 6156 4013 6164
rect 4307 6156 4393 6164
rect 4407 6156 4793 6164
rect 4807 6156 4973 6164
rect 5287 6156 5593 6164
rect 5647 6156 5824 6164
rect 5816 6147 5824 6156
rect 607 6136 753 6144
rect 807 6136 853 6144
rect 3307 6136 3333 6144
rect 5027 6136 5213 6144
rect 5447 6136 5473 6144
rect 5527 6136 5553 6144
rect 5827 6136 5933 6144
rect 187 6117 213 6125
rect 256 6116 292 6124
rect 256 6104 264 6116
rect 327 6117 353 6125
rect 527 6116 644 6124
rect 236 6096 264 6104
rect 636 6104 644 6116
rect 967 6117 1013 6125
rect 1147 6116 1233 6124
rect 1416 6116 1473 6124
rect 636 6096 684 6104
rect 236 6086 244 6096
rect 287 6076 313 6084
rect 427 6075 473 6083
rect 676 6086 684 6096
rect 607 6076 633 6084
rect 696 6084 704 6114
rect 836 6096 873 6104
rect 696 6076 773 6084
rect 836 6084 844 6096
rect 827 6076 844 6084
rect 947 6076 1113 6084
rect 1336 6084 1344 6114
rect 1236 6076 1344 6084
rect 1236 6064 1244 6076
rect 867 6056 1244 6064
rect 1267 6056 1333 6064
rect 1416 6064 1424 6116
rect 1527 6117 1573 6125
rect 1747 6117 1813 6125
rect 1927 6117 1953 6125
rect 2127 6117 2173 6125
rect 2467 6117 2573 6125
rect 2747 6117 2773 6125
rect 2967 6116 3033 6124
rect 1447 6075 1493 6083
rect 1687 6075 1713 6083
rect 1727 6076 1793 6084
rect 1927 6075 2093 6083
rect 2187 6076 2253 6084
rect 2276 6084 2284 6113
rect 2276 6076 2353 6084
rect 2367 6076 2513 6084
rect 2816 6084 2824 6114
rect 3467 6117 3493 6125
rect 3587 6117 3613 6125
rect 3667 6116 3773 6124
rect 3787 6117 3892 6125
rect 3927 6117 3953 6125
rect 4007 6117 4033 6125
rect 4107 6116 4132 6124
rect 4167 6117 4193 6125
rect 4247 6116 4353 6124
rect 3676 6096 3964 6104
rect 2727 6076 2824 6084
rect 3047 6075 3073 6083
rect 3227 6076 3293 6084
rect 3676 6086 3684 6096
rect 3907 6076 3933 6084
rect 3956 6084 3964 6096
rect 3956 6076 4253 6084
rect 1347 6056 1424 6064
rect 1987 6056 2033 6064
rect 3987 6056 4013 6064
rect 4147 6056 4233 6064
rect 4336 6064 4344 6116
rect 4507 6116 4553 6124
rect 4847 6117 4893 6125
rect 5036 6116 5133 6124
rect 5036 6086 5044 6116
rect 5536 6116 5593 6124
rect 5396 6087 5404 6114
rect 5496 6087 5504 6114
rect 5536 6104 5544 6116
rect 4467 6075 4513 6083
rect 4567 6075 4813 6083
rect 5127 6076 5173 6084
rect 5227 6076 5293 6084
rect 5387 6076 5404 6087
rect 5387 6073 5400 6076
rect 5487 6076 5504 6087
rect 5516 6096 5544 6104
rect 5736 6104 5744 6114
rect 5736 6096 5793 6104
rect 5516 6086 5524 6096
rect 5487 6073 5500 6076
rect 5587 6076 5713 6084
rect 4307 6056 4344 6064
rect 5107 6056 5193 6064
rect 5767 6056 5953 6064
rect 547 6036 633 6044
rect 787 6036 1493 6044
rect 1507 6036 1833 6044
rect 1847 6036 2713 6044
rect 2727 6036 2753 6044
rect 3007 6036 3393 6044
rect 3407 6036 3453 6044
rect 3647 6036 3713 6044
rect 4227 6036 4273 6044
rect 4407 6036 4492 6044
rect 4527 6036 4573 6044
rect 4587 6036 4673 6044
rect 4947 6036 5113 6044
rect 5227 6036 5413 6044
rect 5667 6036 5733 6044
rect 807 6016 973 6024
rect 987 6016 1393 6024
rect 1747 6016 1953 6024
rect 3787 6016 4153 6024
rect 4167 6016 4333 6024
rect 4347 6016 5153 6024
rect 5167 6016 5473 6024
rect 607 5996 853 6004
rect 1367 5996 1573 6004
rect 2067 5996 3553 6004
rect 3807 5996 4193 6004
rect 4247 5996 4332 6004
rect 4367 5996 4433 6004
rect 4807 5996 4853 6004
rect 4907 5996 5213 6004
rect 5387 5996 5413 6004
rect 5767 5996 5793 6004
rect 5807 5996 5973 6004
rect 667 5976 793 5984
rect 1027 5976 1193 5984
rect 1207 5976 1413 5984
rect 3507 5976 3573 5984
rect 3587 5976 3753 5984
rect 3767 5976 4473 5984
rect 4647 5976 4733 5984
rect 4747 5976 4993 5984
rect 5747 5976 5793 5984
rect 5807 5976 5933 5984
rect 387 5956 633 5964
rect 1787 5956 1873 5964
rect 2147 5956 2433 5964
rect 4207 5956 4453 5964
rect 4727 5956 4773 5964
rect 4816 5956 5113 5964
rect 1007 5936 1073 5944
rect 1407 5936 1633 5944
rect 1907 5936 2113 5944
rect 2567 5936 2633 5944
rect 2647 5936 2833 5944
rect 3287 5936 3353 5944
rect 3987 5936 4033 5944
rect 4047 5936 4133 5944
rect 4147 5936 4444 5944
rect 127 5916 393 5924
rect 4436 5927 4444 5936
rect 4507 5936 4533 5944
rect 4816 5944 4824 5956
rect 5547 5956 5653 5964
rect 5867 5956 6113 5964
rect 4627 5936 4824 5944
rect 4847 5936 4913 5944
rect 4927 5936 5253 5944
rect 5507 5936 5693 5944
rect 5947 5936 6033 5944
rect 407 5916 553 5924
rect 1136 5916 1233 5924
rect 1136 5908 1144 5916
rect 2987 5916 3153 5924
rect 3167 5916 3364 5924
rect 156 5864 164 5894
rect 227 5896 273 5904
rect 347 5897 393 5905
rect 447 5896 493 5904
rect 747 5896 813 5904
rect 827 5896 893 5904
rect 1067 5897 1133 5905
rect 1307 5897 1393 5905
rect 1567 5897 1613 5905
rect 1887 5897 1993 5905
rect 2267 5896 2353 5904
rect 2367 5896 2453 5904
rect 936 5884 944 5894
rect 1676 5884 1684 5894
rect 1816 5884 1824 5894
rect 2467 5896 2524 5904
rect 936 5876 1004 5884
rect 1676 5876 1824 5884
rect 156 5856 293 5864
rect 427 5856 533 5864
rect 547 5856 564 5864
rect 347 5836 393 5844
rect 556 5844 564 5856
rect 587 5855 613 5863
rect 996 5864 1004 5876
rect 1816 5867 1824 5876
rect 996 5856 1213 5864
rect 1227 5856 1313 5864
rect 1427 5856 1473 5864
rect 1607 5856 1693 5864
rect 1807 5856 1824 5867
rect 1807 5853 1820 5856
rect 1847 5856 1973 5864
rect 2027 5856 2113 5864
rect 2387 5856 2473 5864
rect 2516 5864 2524 5896
rect 2547 5897 2573 5905
rect 2687 5896 2713 5904
rect 3047 5896 3164 5904
rect 2516 5856 2613 5864
rect 2667 5856 2773 5864
rect 2993 5863 3007 5873
rect 2887 5855 3133 5863
rect 3156 5864 3164 5896
rect 3207 5896 3324 5904
rect 3316 5866 3324 5896
rect 3356 5904 3364 5916
rect 3527 5916 3564 5924
rect 3356 5896 3373 5904
rect 3556 5904 3564 5916
rect 3627 5916 3673 5924
rect 4267 5916 4293 5924
rect 4387 5916 4424 5924
rect 3556 5896 3693 5904
rect 3156 5856 3173 5864
rect 556 5836 713 5844
rect 927 5836 1033 5844
rect 1387 5836 2053 5844
rect 3336 5845 3344 5894
rect 3456 5864 3464 5894
rect 4147 5896 4204 5904
rect 3516 5876 3673 5884
rect 3516 5866 3524 5876
rect 4096 5884 4104 5894
rect 4096 5880 4183 5884
rect 4096 5876 4187 5880
rect 4173 5867 4187 5876
rect 3367 5856 3464 5864
rect 3567 5856 3633 5864
rect 3707 5855 3793 5863
rect 3927 5856 4073 5864
rect 4186 5860 4187 5867
rect 4196 5866 4204 5896
rect 4416 5904 4424 5916
rect 4447 5916 4953 5924
rect 4416 5896 4613 5904
rect 4216 5864 4224 5894
rect 4687 5904 4700 5907
rect 4740 5904 4753 5907
rect 4687 5893 4704 5904
rect 4216 5856 4273 5864
rect 4696 5866 4704 5893
rect 4736 5893 4753 5904
rect 4807 5896 4864 5904
rect 4736 5866 4744 5893
rect 4856 5866 4864 5896
rect 4887 5896 4933 5904
rect 5036 5867 5044 5894
rect 5127 5904 5140 5907
rect 5127 5893 5144 5904
rect 5167 5896 5204 5904
rect 4347 5855 4373 5863
rect 4487 5855 4513 5863
rect 4607 5855 4633 5863
rect 4787 5855 4813 5863
rect 5027 5856 5044 5867
rect 5136 5866 5144 5893
rect 5027 5853 5040 5856
rect 5196 5864 5204 5896
rect 5227 5896 5284 5904
rect 5276 5866 5284 5896
rect 5327 5897 5373 5905
rect 5487 5897 5533 5905
rect 5716 5896 5833 5904
rect 5196 5856 5233 5864
rect 5407 5856 5553 5864
rect 5576 5864 5584 5894
rect 5716 5866 5724 5896
rect 5956 5884 5964 5894
rect 5876 5880 5964 5884
rect 5873 5876 5964 5880
rect 5873 5867 5887 5876
rect 5576 5856 5673 5864
rect 5987 5856 6033 5864
rect 6047 5856 6093 5864
rect 3336 5833 3353 5845
rect 3967 5836 4013 5844
rect 5107 5836 5173 5844
rect 5907 5836 5953 5844
rect 107 5816 193 5824
rect 207 5816 373 5824
rect 487 5816 553 5824
rect 567 5816 613 5824
rect 1267 5816 1353 5824
rect 1567 5816 1873 5824
rect 1887 5816 2273 5824
rect 2527 5816 2913 5824
rect 3207 5816 3393 5824
rect 3407 5816 3553 5824
rect 4087 5816 4413 5824
rect 4427 5816 4813 5824
rect 5207 5816 5293 5824
rect 5487 5816 5853 5824
rect 727 5796 773 5804
rect 2747 5796 2853 5804
rect 3247 5796 3413 5804
rect 3807 5796 4113 5804
rect 4127 5796 4273 5804
rect 4387 5796 4924 5804
rect 187 5776 253 5784
rect 716 5784 724 5793
rect 267 5776 724 5784
rect 1287 5776 1533 5784
rect 1547 5776 1913 5784
rect 3287 5776 3473 5784
rect 3607 5776 3653 5784
rect 3667 5776 3853 5784
rect 3867 5776 4053 5784
rect 4916 5784 4924 5796
rect 5687 5796 5813 5804
rect 4916 5776 5113 5784
rect 5167 5776 5453 5784
rect 3067 5756 3093 5764
rect 3107 5756 3233 5764
rect 3607 5756 3793 5764
rect 3947 5756 4033 5764
rect 5107 5756 5193 5764
rect 5527 5756 5713 5764
rect 1747 5736 1793 5744
rect 1807 5736 2233 5744
rect 3347 5736 3893 5744
rect 4827 5736 4953 5744
rect 4967 5736 5153 5744
rect 5307 5736 5564 5744
rect 167 5716 473 5724
rect 487 5716 613 5724
rect 1767 5716 1913 5724
rect 2427 5716 2833 5724
rect 3387 5716 3693 5724
rect 3867 5716 4233 5724
rect 4247 5716 4733 5724
rect 5247 5716 5473 5724
rect 5556 5724 5564 5736
rect 5556 5716 6124 5724
rect 6116 5707 6124 5716
rect 307 5696 813 5704
rect 1947 5696 2853 5704
rect 2867 5696 2913 5704
rect 3027 5696 3953 5704
rect 4007 5696 4593 5704
rect 4867 5696 5133 5704
rect 5267 5696 5313 5704
rect 5467 5696 5533 5704
rect 5547 5696 5753 5704
rect 5767 5696 5853 5704
rect 6116 5696 6133 5707
rect 6120 5693 6133 5696
rect 1107 5676 1153 5684
rect 1787 5676 1993 5684
rect 3247 5676 3933 5684
rect 4427 5676 4553 5684
rect 4827 5676 4933 5684
rect 5087 5676 5193 5684
rect 5627 5676 5713 5684
rect 5727 5676 5933 5684
rect 227 5656 273 5664
rect 867 5656 1253 5664
rect 2447 5656 2693 5664
rect 3367 5656 3433 5664
rect 3527 5656 3673 5664
rect 5076 5664 5084 5673
rect 4027 5656 5084 5664
rect 5167 5656 5273 5664
rect 587 5636 633 5644
rect 807 5636 1033 5644
rect 2496 5636 2593 5644
rect 2496 5627 2504 5636
rect 2636 5636 2753 5644
rect 107 5616 204 5624
rect 87 5596 173 5604
rect 196 5564 204 5616
rect 1147 5616 1233 5624
rect 1627 5616 1793 5624
rect 1856 5616 1953 5624
rect 247 5597 293 5605
rect 336 5584 344 5594
rect 407 5604 420 5607
rect 407 5593 424 5604
rect 447 5597 533 5605
rect 547 5596 673 5604
rect 827 5596 913 5604
rect 1167 5597 1193 5605
rect 1487 5596 1573 5604
rect 1587 5596 1653 5604
rect 336 5576 384 5584
rect 376 5567 384 5576
rect 196 5556 213 5564
rect 307 5556 353 5564
rect 376 5556 393 5567
rect 380 5553 393 5556
rect 416 5564 424 5593
rect 796 5576 853 5584
rect 416 5556 613 5564
rect 796 5566 804 5576
rect 727 5556 753 5564
rect 1087 5556 1133 5564
rect 1256 5564 1264 5593
rect 1227 5556 1264 5564
rect 1316 5564 1324 5594
rect 1856 5604 1864 5616
rect 2133 5616 2233 5624
rect 2133 5608 2147 5616
rect 2247 5616 2284 5624
rect 1847 5596 1864 5604
rect 1887 5597 1933 5605
rect 2067 5596 2133 5604
rect 2187 5597 2213 5605
rect 2276 5604 2284 5616
rect 2407 5616 2493 5624
rect 2636 5624 2644 5636
rect 3107 5636 3133 5644
rect 3147 5636 3253 5644
rect 4047 5636 4373 5644
rect 4527 5636 4693 5644
rect 4847 5636 5024 5644
rect 2567 5616 2644 5624
rect 5016 5624 5024 5636
rect 5127 5636 5293 5644
rect 5847 5636 5873 5644
rect 5887 5636 5993 5644
rect 5016 5616 5053 5624
rect 5067 5616 5233 5624
rect 2276 5596 2333 5604
rect 2467 5597 2533 5605
rect 2667 5596 2684 5604
rect 1936 5584 1944 5594
rect 1396 5576 1944 5584
rect 1396 5564 1404 5576
rect 2676 5567 2684 5596
rect 2967 5597 2993 5605
rect 3187 5597 3273 5605
rect 2733 5584 2747 5593
rect 2733 5580 2784 5584
rect 2736 5576 2784 5580
rect 1316 5556 1404 5564
rect 1547 5556 1593 5564
rect 1667 5555 1713 5563
rect 1867 5556 1913 5564
rect 2167 5556 2253 5564
rect 2776 5566 2784 5576
rect 2796 5547 2804 5594
rect 3287 5597 3333 5605
rect 3807 5596 3833 5604
rect 3227 5556 3304 5564
rect 487 5536 533 5544
rect 1967 5536 2113 5544
rect 2327 5536 2393 5544
rect 2887 5536 2953 5544
rect 3296 5544 3304 5556
rect 3476 5564 3484 5594
rect 3556 5584 3564 5594
rect 3696 5584 3704 5594
rect 3556 5580 3584 5584
rect 3636 5580 3704 5584
rect 3556 5576 3587 5580
rect 3327 5556 3484 5564
rect 3573 5567 3587 5576
rect 3633 5576 3704 5580
rect 3633 5567 3647 5576
rect 3876 5567 3884 5593
rect 3936 5567 3944 5594
rect 4107 5597 4133 5605
rect 4287 5597 4313 5605
rect 4447 5597 4473 5605
rect 4756 5596 4773 5604
rect 4016 5567 4024 5593
rect 3687 5556 3852 5564
rect 3936 5556 3953 5567
rect 3940 5553 3953 5556
rect 4196 5564 4204 5594
rect 4196 5556 4333 5564
rect 4356 5564 4364 5594
rect 4636 5567 4644 5594
rect 4356 5556 4493 5564
rect 4636 5556 4653 5567
rect 4640 5553 4653 5556
rect 3296 5536 3433 5544
rect 3476 5536 3553 5544
rect 47 5516 133 5524
rect 887 5516 933 5524
rect 947 5516 1333 5524
rect 1347 5516 1393 5524
rect 1507 5516 1693 5524
rect 2167 5516 2233 5524
rect 2287 5516 2313 5524
rect 2327 5516 2353 5524
rect 3027 5516 3053 5524
rect 3476 5524 3484 5536
rect 4187 5536 4253 5544
rect 4756 5544 4764 5596
rect 5036 5596 5153 5604
rect 4916 5584 4924 5593
rect 5036 5584 5044 5596
rect 5287 5596 5404 5604
rect 4816 5580 5044 5584
rect 4813 5576 5044 5580
rect 5396 5584 5404 5596
rect 5527 5596 5573 5604
rect 5600 5604 5613 5607
rect 5596 5593 5613 5604
rect 5816 5596 5833 5604
rect 5396 5576 5424 5584
rect 4813 5567 4827 5576
rect 4947 5556 5073 5564
rect 5127 5555 5213 5563
rect 5416 5564 5424 5576
rect 5596 5566 5604 5593
rect 5676 5567 5684 5593
rect 5416 5556 5493 5564
rect 5756 5564 5764 5594
rect 5756 5556 5793 5564
rect 4627 5536 4764 5544
rect 5527 5536 5573 5544
rect 5816 5544 5824 5596
rect 5867 5556 5933 5564
rect 6027 5556 6073 5564
rect 5747 5536 5824 5544
rect 3347 5516 3484 5524
rect 3667 5516 3853 5524
rect 4007 5516 4033 5524
rect 4087 5516 4373 5524
rect 4387 5516 4433 5524
rect 4447 5516 4593 5524
rect 4647 5516 4833 5524
rect 5047 5516 5193 5524
rect 5447 5516 5833 5524
rect 5887 5516 5953 5524
rect 1467 5496 1633 5504
rect 1727 5496 1893 5504
rect 1947 5496 2133 5504
rect 2207 5496 2253 5504
rect 2267 5496 2393 5504
rect 2627 5496 2933 5504
rect 3187 5496 3472 5504
rect 3507 5496 3633 5504
rect 3687 5496 3873 5504
rect 4467 5496 4533 5504
rect 4707 5496 4772 5504
rect 4807 5496 4853 5504
rect 5027 5496 5153 5504
rect 5327 5496 5413 5504
rect 107 5476 133 5484
rect 367 5476 393 5484
rect 407 5476 453 5484
rect 467 5476 653 5484
rect 1707 5476 2433 5484
rect 3147 5476 3233 5484
rect 3367 5476 3393 5484
rect 207 5456 293 5464
rect 1367 5456 1452 5464
rect 1487 5456 1952 5464
rect 1987 5456 2313 5464
rect 2667 5456 2804 5464
rect 67 5436 253 5444
rect 1007 5436 1113 5444
rect 2027 5436 2213 5444
rect 2796 5444 2804 5456
rect 2887 5456 2993 5464
rect 3007 5456 3033 5464
rect 3087 5456 3353 5464
rect 3396 5464 3404 5473
rect 3507 5476 3573 5484
rect 3587 5476 3773 5484
rect 3927 5476 4153 5484
rect 4227 5476 4633 5484
rect 4687 5476 4913 5484
rect 5207 5476 5504 5484
rect 5496 5467 5504 5476
rect 5607 5476 5653 5484
rect 6007 5476 6093 5484
rect 3396 5456 3533 5464
rect 3547 5456 3593 5464
rect 3747 5456 3893 5464
rect 4787 5456 4852 5464
rect 4887 5456 5073 5464
rect 5247 5456 5333 5464
rect 5507 5456 5813 5464
rect 2796 5436 2853 5444
rect 3227 5436 3273 5444
rect 3647 5436 3933 5444
rect 3987 5436 4073 5444
rect 4216 5436 4393 5444
rect 307 5416 413 5424
rect 567 5416 753 5424
rect 767 5416 833 5424
rect 927 5416 1173 5424
rect 1767 5416 1793 5424
rect 2287 5416 2353 5424
rect 2607 5416 2713 5424
rect 3207 5416 3533 5424
rect 4216 5424 4224 5436
rect 4547 5436 4713 5444
rect 5167 5436 6033 5444
rect 6047 5436 6093 5444
rect 6107 5436 6184 5444
rect 4107 5416 4224 5424
rect 4427 5416 4613 5424
rect 4767 5416 4832 5424
rect 4867 5416 5013 5424
rect 5267 5416 5332 5424
rect 5367 5416 5533 5424
rect 5647 5416 5693 5424
rect 5747 5416 5953 5424
rect 227 5396 273 5404
rect 587 5396 613 5404
rect 627 5396 673 5404
rect 2547 5396 2613 5404
rect 3147 5396 3173 5404
rect 3307 5396 3373 5404
rect 3427 5404 3440 5407
rect 3427 5393 3444 5404
rect 5207 5396 5233 5404
rect 5287 5396 5393 5404
rect 5767 5396 5793 5404
rect 6147 5396 6204 5404
rect 27 5377 133 5385
rect 416 5376 513 5384
rect 227 5335 273 5343
rect 416 5327 424 5376
rect 727 5376 773 5384
rect 887 5376 924 5384
rect 916 5364 924 5376
rect 947 5377 973 5385
rect 1027 5376 1073 5384
rect 1196 5376 1273 5384
rect 916 5356 964 5364
rect 587 5335 613 5343
rect 667 5335 753 5343
rect 956 5344 964 5356
rect 1196 5346 1204 5376
rect 1327 5376 1393 5384
rect 1567 5376 1633 5384
rect 1647 5376 1753 5384
rect 1847 5376 1873 5384
rect 1887 5377 1913 5385
rect 2027 5377 2053 5385
rect 2507 5376 2544 5384
rect 956 5336 993 5344
rect 167 5316 193 5324
rect 616 5324 624 5332
rect 616 5316 813 5324
rect 1807 5316 1873 5324
rect 2276 5324 2284 5373
rect 2316 5364 2324 5374
rect 2296 5360 2324 5364
rect 2293 5356 2324 5360
rect 2293 5347 2307 5356
rect 2427 5336 2453 5344
rect 2536 5344 2544 5376
rect 2676 5346 2684 5393
rect 2727 5377 2753 5385
rect 2896 5347 2904 5374
rect 3047 5376 3184 5384
rect 3176 5364 3184 5376
rect 3436 5384 3444 5393
rect 3436 5376 3464 5384
rect 3176 5360 3264 5364
rect 3176 5356 3267 5360
rect 3253 5347 3267 5356
rect 2536 5336 2633 5344
rect 2827 5335 2853 5343
rect 2887 5336 2904 5347
rect 2887 5333 2900 5336
rect 2967 5336 3033 5344
rect 3167 5336 3193 5344
rect 3336 5344 3344 5373
rect 3327 5336 3344 5344
rect 3387 5335 3413 5343
rect 3456 5327 3464 5376
rect 3496 5346 3504 5393
rect 3547 5376 3584 5384
rect 3576 5346 3584 5376
rect 3607 5376 3713 5384
rect 3767 5376 3812 5384
rect 3847 5376 3924 5384
rect 3916 5364 3924 5376
rect 3947 5376 4144 5384
rect 3916 5360 4123 5364
rect 3916 5356 4127 5360
rect 4113 5347 4127 5356
rect 3627 5336 3912 5344
rect 3947 5335 4013 5343
rect 4126 5340 4127 5347
rect 4136 5346 4144 5376
rect 4207 5376 4433 5384
rect 4447 5376 4493 5384
rect 4567 5376 4584 5384
rect 4576 5364 4584 5376
rect 4607 5377 4793 5385
rect 4887 5377 4953 5385
rect 5036 5376 5133 5384
rect 4576 5356 4664 5364
rect 4187 5336 4253 5344
rect 4327 5336 4373 5344
rect 4656 5346 4664 5356
rect 4996 5347 5004 5373
rect 4507 5335 4533 5343
rect 5036 5327 5044 5376
rect 5367 5376 5404 5384
rect 5176 5344 5184 5373
rect 5107 5336 5184 5344
rect 5216 5344 5224 5373
rect 5396 5364 5404 5376
rect 5560 5384 5573 5387
rect 5447 5376 5524 5384
rect 5396 5356 5424 5364
rect 5216 5336 5253 5344
rect 5416 5346 5424 5356
rect 5516 5346 5524 5376
rect 5556 5373 5573 5384
rect 5556 5346 5564 5373
rect 5347 5336 5373 5344
rect 5656 5344 5664 5374
rect 6100 5384 6113 5387
rect 6096 5373 6113 5384
rect 5656 5336 5733 5344
rect 5836 5344 5844 5373
rect 6096 5347 6104 5373
rect 6176 5364 6184 5384
rect 6147 5356 6184 5364
rect 5827 5336 5844 5344
rect 5867 5336 5933 5344
rect 6096 5336 6113 5347
rect 6100 5333 6113 5336
rect 6196 5344 6204 5396
rect 6176 5336 6204 5344
rect 2276 5316 2313 5324
rect 2787 5316 2913 5324
rect 3447 5316 3464 5327
rect 3447 5313 3460 5316
rect 4307 5316 4713 5324
rect 4727 5316 4753 5324
rect 4807 5316 4973 5324
rect 5027 5316 5044 5327
rect 5027 5313 5040 5316
rect 196 5304 204 5313
rect 196 5296 393 5304
rect 707 5296 853 5304
rect 987 5296 1033 5304
rect 1087 5296 1293 5304
rect 1827 5296 1933 5304
rect 2087 5296 2153 5304
rect 2167 5296 2333 5304
rect 2447 5296 2573 5304
rect 2776 5304 2784 5313
rect 2667 5296 2784 5304
rect 3436 5304 3444 5313
rect 3436 5296 3613 5304
rect 3827 5296 3993 5304
rect 4087 5296 4213 5304
rect 4367 5296 4453 5304
rect 4756 5296 4873 5304
rect 107 5276 312 5284
rect 347 5276 533 5284
rect 1167 5276 1253 5284
rect 2287 5276 2473 5284
rect 2887 5276 3093 5284
rect 3107 5276 3213 5284
rect 3227 5276 3973 5284
rect 4756 5284 4764 5296
rect 4887 5296 5033 5304
rect 5507 5296 5673 5304
rect 5827 5296 5893 5304
rect 4427 5276 4764 5284
rect 5087 5276 5213 5284
rect 5427 5276 5713 5284
rect 5807 5276 6013 5284
rect 6067 5276 6133 5284
rect 447 5256 1473 5264
rect 1587 5256 1773 5264
rect 1787 5256 2013 5264
rect 2067 5256 2113 5264
rect 2247 5256 2552 5264
rect 2587 5256 2613 5264
rect 2627 5256 2804 5264
rect 436 5244 444 5253
rect 27 5236 444 5244
rect 567 5236 933 5244
rect 1147 5236 1233 5244
rect 1507 5236 1653 5244
rect 1667 5236 1912 5244
rect 1947 5236 2193 5244
rect 2307 5236 2333 5244
rect 2796 5244 2804 5256
rect 2907 5256 2933 5264
rect 3467 5256 3733 5264
rect 3927 5256 4233 5264
rect 4487 5256 4893 5264
rect 4987 5256 5053 5264
rect 5116 5256 5753 5264
rect 2796 5236 3013 5244
rect 3187 5236 3213 5244
rect 3347 5236 3493 5244
rect 3507 5236 3713 5244
rect 3887 5236 3933 5244
rect 3987 5236 4333 5244
rect 5116 5244 5124 5256
rect 4507 5236 5124 5244
rect 5147 5236 5413 5244
rect 5787 5236 5873 5244
rect 207 5216 353 5224
rect 2027 5216 2073 5224
rect 2787 5216 3053 5224
rect 3367 5216 3773 5224
rect 4047 5216 4153 5224
rect 4387 5216 4453 5224
rect 4667 5216 4733 5224
rect 4747 5216 4973 5224
rect 5067 5216 5313 5224
rect 5387 5216 6053 5224
rect 527 5196 693 5204
rect 1107 5196 1173 5204
rect 1547 5196 1873 5204
rect 1927 5196 2153 5204
rect 2627 5196 2713 5204
rect 2927 5196 3253 5204
rect 3407 5196 3513 5204
rect 4187 5196 4293 5204
rect 4347 5196 4513 5204
rect 4927 5196 5073 5204
rect 5267 5196 5513 5204
rect 5527 5196 5733 5204
rect 5747 5196 6033 5204
rect 1407 5176 2073 5184
rect 2147 5176 2193 5184
rect 2607 5176 2753 5184
rect 2987 5176 3013 5184
rect 3547 5176 3633 5184
rect 3967 5176 4033 5184
rect 4267 5176 4553 5184
rect 4787 5176 5004 5184
rect 4996 5167 5004 5176
rect 5047 5176 5372 5184
rect 5407 5176 5673 5184
rect 787 5156 973 5164
rect 1107 5156 1373 5164
rect 1467 5156 1613 5164
rect 2527 5156 2673 5164
rect 2987 5156 3113 5164
rect 3167 5156 3433 5164
rect 3727 5156 3813 5164
rect 4027 5156 4133 5164
rect 4207 5156 4573 5164
rect 4647 5156 4933 5164
rect 5007 5156 5113 5164
rect 5467 5156 5593 5164
rect 107 5136 333 5144
rect 467 5136 553 5144
rect 3287 5136 3553 5144
rect 3607 5136 3893 5144
rect 4127 5136 4153 5144
rect 4167 5136 4413 5144
rect 5687 5136 5853 5144
rect 1167 5116 1353 5124
rect 1767 5116 2113 5124
rect 2127 5116 2204 5124
rect 367 5096 673 5104
rect 1307 5096 1333 5104
rect 1487 5096 1533 5104
rect 2196 5104 2204 5116
rect 2527 5116 2573 5124
rect 2647 5116 2693 5124
rect 3707 5116 3773 5124
rect 3847 5116 3953 5124
rect 4000 5124 4013 5127
rect 3996 5113 4013 5124
rect 4066 5113 4067 5120
rect 4087 5116 4224 5124
rect 2196 5096 2353 5104
rect 2407 5096 2613 5104
rect 67 5077 133 5085
rect 147 5076 253 5084
rect 307 5077 513 5085
rect 727 5077 753 5085
rect 827 5076 873 5084
rect 896 5076 1093 5084
rect 896 5064 904 5076
rect 1427 5077 1453 5085
rect 1627 5077 1653 5085
rect 1667 5076 1753 5084
rect 1826 5073 1827 5080
rect 1927 5077 1953 5085
rect 2167 5076 2304 5084
rect 1813 5064 1827 5073
rect 836 5056 904 5064
rect 1756 5060 1827 5064
rect 1756 5056 1823 5060
rect 836 5046 844 5056
rect 47 5035 153 5043
rect 167 5036 233 5044
rect 1367 5036 1593 5044
rect 1756 5044 1764 5056
rect 1747 5036 1764 5044
rect 1836 5044 1844 5074
rect 2296 5047 2304 5076
rect 2556 5064 2564 5074
rect 2347 5056 2564 5064
rect 1787 5036 1844 5044
rect 1907 5036 2053 5044
rect 2576 5046 2584 5096
rect 2796 5096 2833 5104
rect 2627 5076 2693 5084
rect 2796 5064 2804 5096
rect 3996 5104 4004 5113
rect 3567 5096 4004 5104
rect 4053 5104 4067 5113
rect 4053 5100 4093 5104
rect 4055 5096 4093 5100
rect 4147 5096 4204 5104
rect 2827 5076 2973 5084
rect 3307 5076 3393 5084
rect 3016 5064 3024 5074
rect 3487 5076 3593 5084
rect 3796 5076 3873 5084
rect 3736 5064 3744 5074
rect 2796 5056 2824 5064
rect 3016 5056 3084 5064
rect 2467 5035 2493 5043
rect 2587 5036 2713 5044
rect 2816 5027 2824 5056
rect 2927 5036 2993 5044
rect 3076 5044 3084 5056
rect 3696 5056 3744 5064
rect 3076 5036 3093 5044
rect 3187 5035 3273 5043
rect 3367 5035 3493 5043
rect 3507 5036 3533 5044
rect 3696 5044 3704 5056
rect 3627 5036 3704 5044
rect 3796 5044 3804 5076
rect 3947 5084 3960 5087
rect 3947 5073 3964 5084
rect 3727 5036 3804 5044
rect 3956 5044 3964 5073
rect 4116 5047 4124 5074
rect 3956 5036 4013 5044
rect 4116 5036 4133 5047
rect 4120 5033 4133 5036
rect 4196 5044 4204 5096
rect 4216 5084 4224 5116
rect 4567 5116 4833 5124
rect 5007 5116 5173 5124
rect 5487 5116 5613 5124
rect 5627 5116 5993 5124
rect 6007 5116 6093 5124
rect 4247 5096 4344 5104
rect 4336 5084 4344 5096
rect 4427 5096 4587 5104
rect 4573 5088 4587 5096
rect 4827 5096 4913 5104
rect 5167 5096 5193 5104
rect 5836 5096 5893 5104
rect 4216 5076 4244 5084
rect 4336 5076 4492 5084
rect 4236 5064 4244 5076
rect 4356 5064 4364 5076
rect 4527 5076 4544 5084
rect 4236 5056 4344 5064
rect 4356 5056 4384 5064
rect 4336 5047 4344 5056
rect 4196 5036 4233 5044
rect 4247 5036 4313 5044
rect 4336 5036 4353 5047
rect 4340 5033 4353 5036
rect 4376 5044 4384 5056
rect 4536 5047 4544 5076
rect 4587 5076 4693 5084
rect 4376 5036 4493 5044
rect 4727 5036 4813 5044
rect 4876 5044 4884 5074
rect 5176 5076 5253 5084
rect 5096 5047 5104 5073
rect 4876 5036 4993 5044
rect 5176 5046 5184 5076
rect 5307 5077 5352 5085
rect 5387 5077 5413 5085
rect 5440 5084 5453 5087
rect 5436 5073 5453 5084
rect 5596 5076 5713 5084
rect 5436 5046 5444 5073
rect 5496 5044 5504 5073
rect 5596 5064 5604 5076
rect 5836 5084 5844 5096
rect 5907 5096 5973 5104
rect 5727 5076 5844 5084
rect 5867 5076 5984 5084
rect 5576 5056 5604 5064
rect 5576 5046 5584 5056
rect 5976 5046 5984 5076
rect 6047 5077 6073 5085
rect 5496 5036 5533 5044
rect 5627 5035 5693 5043
rect 127 5016 353 5024
rect 707 5016 773 5024
rect 887 5016 993 5024
rect 1227 5016 1253 5024
rect 1307 5016 1333 5024
rect 1347 5016 1473 5024
rect 1807 5016 1853 5024
rect 1927 5016 1953 5024
rect 2367 5016 2413 5024
rect 3067 5016 3313 5024
rect 3647 5016 3673 5024
rect 3867 5016 3892 5024
rect 3927 5016 4073 5024
rect 4447 5016 4633 5024
rect 4747 5016 4773 5024
rect 5067 5016 5153 5024
rect 5947 5016 6093 5024
rect 507 4996 633 5004
rect 1587 4996 1673 5004
rect 1687 4996 1753 5004
rect 2047 4996 2193 5004
rect 3507 4996 3713 5004
rect 3916 5004 3924 5013
rect 3807 4996 3924 5004
rect 4127 4996 4213 5004
rect 4867 4996 5304 5004
rect 287 4976 433 4984
rect 927 4976 1064 4984
rect 427 4956 513 4964
rect 587 4956 753 4964
rect 767 4956 792 4964
rect 827 4956 953 4964
rect 1056 4964 1064 4976
rect 1087 4976 1173 4984
rect 1607 4976 1773 4984
rect 1987 4976 2133 4984
rect 2147 4976 2253 4984
rect 2427 4976 2933 4984
rect 3307 4976 3473 4984
rect 3567 4976 3593 4984
rect 3667 4976 3753 4984
rect 3827 4976 4013 4984
rect 4027 4976 4093 4984
rect 4107 4976 4273 4984
rect 4387 4976 4453 4984
rect 4467 4976 4673 4984
rect 4747 4976 4833 4984
rect 4967 4976 5213 4984
rect 5296 4984 5304 4996
rect 5327 4996 5413 5004
rect 5747 4996 5833 5004
rect 5887 4996 5913 5004
rect 5927 4996 6073 5004
rect 5296 4976 5333 4984
rect 5387 4976 5433 4984
rect 5667 4976 5713 4984
rect 1056 4956 1733 4964
rect 2307 4956 2833 4964
rect 2847 4956 2953 4964
rect 2967 4956 3053 4964
rect 3227 4956 3393 4964
rect 4207 4956 4233 4964
rect 4327 4956 4553 4964
rect 4676 4964 4684 4973
rect 4676 4956 4713 4964
rect 5147 4956 5353 4964
rect 5707 4956 5753 4964
rect 5827 4956 5873 4964
rect 1027 4936 1273 4944
rect 1467 4936 1713 4944
rect 3187 4936 3293 4944
rect 3487 4936 3773 4944
rect 3787 4936 3813 4944
rect 4147 4936 4293 4944
rect 4627 4936 4733 4944
rect 4787 4936 4993 4944
rect 5387 4936 5593 4944
rect 5807 4936 5893 4944
rect 1327 4916 1653 4924
rect 2407 4916 2473 4924
rect 2487 4916 2512 4924
rect 2547 4916 2593 4924
rect 3147 4916 3393 4924
rect 3467 4916 3793 4924
rect 3947 4916 3993 4924
rect 4067 4916 4113 4924
rect 4207 4916 4633 4924
rect 5047 4916 5113 4924
rect 6027 4916 6124 4924
rect 6116 4907 6124 4916
rect 407 4896 493 4904
rect 1567 4896 1693 4904
rect 1707 4896 1813 4904
rect 2087 4896 2153 4904
rect 2367 4896 2433 4904
rect 2627 4896 2793 4904
rect 2847 4896 2993 4904
rect 3007 4896 3053 4904
rect 3207 4896 3313 4904
rect 3447 4896 3913 4904
rect 4187 4896 4393 4904
rect 4567 4896 4653 4904
rect 4947 4896 5333 4904
rect 5647 4896 5713 4904
rect 6116 4896 6133 4907
rect 6120 4893 6133 4896
rect 187 4876 233 4884
rect 247 4876 553 4884
rect 567 4876 693 4884
rect 976 4876 1013 4884
rect 127 4856 164 4864
rect 156 4827 164 4856
rect 287 4856 313 4864
rect 387 4857 473 4865
rect 576 4856 593 4864
rect 576 4844 584 4856
rect 747 4856 853 4864
rect 976 4844 984 4876
rect 2607 4876 2684 4884
rect 1107 4857 1113 4865
rect 1127 4857 1133 4865
rect 1207 4856 1313 4864
rect 1367 4857 1413 4865
rect 1607 4856 1653 4864
rect 2227 4856 2273 4864
rect 516 4836 584 4844
rect 876 4836 984 4844
rect 1816 4844 1824 4854
rect 1816 4836 1964 4844
rect 327 4815 393 4823
rect 516 4824 524 4836
rect 447 4820 564 4824
rect 447 4816 567 4820
rect 553 4807 567 4816
rect 667 4816 813 4824
rect 876 4826 884 4836
rect 976 4826 984 4836
rect 1027 4816 1153 4824
rect 1547 4816 1713 4824
rect 1727 4816 1853 4824
rect 1867 4815 1913 4823
rect 1956 4824 1964 4836
rect 1956 4816 1973 4824
rect 2087 4816 2193 4824
rect 2247 4815 2293 4823
rect 2336 4824 2344 4873
rect 2336 4816 2413 4824
rect 2676 4826 2684 4876
rect 3707 4876 3824 4884
rect 2767 4856 2833 4864
rect 3047 4856 3124 4864
rect 2876 4844 2884 4854
rect 2876 4836 3004 4844
rect 2727 4815 2753 4823
rect 2807 4815 2853 4823
rect 2996 4824 3004 4836
rect 2996 4816 3024 4824
rect 147 4796 173 4804
rect 1347 4796 1453 4804
rect 1467 4796 1933 4804
rect 2387 4796 2613 4804
rect 2853 4804 2867 4812
rect 3016 4807 3024 4816
rect 2853 4796 2973 4804
rect 3016 4796 3033 4807
rect 3020 4793 3033 4796
rect 3116 4804 3124 4856
rect 3167 4856 3233 4864
rect 3327 4856 3524 4864
rect 3516 4844 3524 4856
rect 3567 4856 3613 4864
rect 3667 4856 3713 4864
rect 3516 4836 3544 4844
rect 3536 4826 3544 4836
rect 3207 4815 3293 4823
rect 3547 4816 3733 4824
rect 3116 4796 3173 4804
rect 3756 4804 3764 4853
rect 3816 4826 3824 4876
rect 4047 4876 4193 4884
rect 3847 4856 3884 4864
rect 3876 4827 3884 4856
rect 3976 4826 3984 4873
rect 4007 4856 4064 4864
rect 4056 4844 4064 4856
rect 4087 4857 4133 4865
rect 4056 4836 4164 4844
rect 4027 4816 4073 4824
rect 4156 4826 4164 4836
rect 4176 4807 4184 4876
rect 4487 4876 4513 4884
rect 4747 4876 4853 4884
rect 5187 4876 5233 4884
rect 5247 4876 5273 4884
rect 5587 4876 5613 4884
rect 5767 4876 5804 4884
rect 4196 4827 4204 4852
rect 4436 4844 4444 4854
rect 4607 4856 4713 4864
rect 4736 4856 4753 4864
rect 4227 4836 4444 4844
rect 4327 4816 4413 4824
rect 4427 4816 4453 4824
rect 3756 4796 3793 4804
rect 4127 4796 4173 4804
rect 4496 4804 4504 4853
rect 4556 4844 4564 4854
rect 4536 4840 4564 4844
rect 4533 4836 4564 4840
rect 4533 4827 4547 4836
rect 4736 4844 4744 4856
rect 4947 4856 4993 4864
rect 5016 4856 5033 4864
rect 5016 4844 5024 4856
rect 5147 4856 5193 4864
rect 5453 4864 5467 4873
rect 5453 4860 5513 4864
rect 5456 4856 5513 4860
rect 4687 4836 4744 4844
rect 4996 4836 5024 4844
rect 4787 4816 4893 4824
rect 4996 4807 5004 4836
rect 5076 4827 5084 4853
rect 5127 4815 5173 4823
rect 5256 4824 5264 4853
rect 5556 4827 5564 4853
rect 5593 4844 5607 4853
rect 5593 4840 5644 4844
rect 5596 4836 5644 4840
rect 5236 4820 5264 4824
rect 5233 4816 5264 4820
rect 5233 4807 5247 4816
rect 5287 4815 5313 4823
rect 5427 4815 5493 4823
rect 5636 4826 5644 4836
rect 5696 4827 5704 4853
rect 5776 4844 5784 4854
rect 5756 4840 5784 4844
rect 5753 4836 5784 4840
rect 5796 4844 5804 4876
rect 5827 4856 6093 4864
rect 5796 4836 5844 4844
rect 5753 4827 5767 4836
rect 5836 4826 5844 4836
rect 4496 4796 4553 4804
rect 267 4776 333 4784
rect 727 4776 873 4784
rect 1267 4776 1393 4784
rect 1647 4776 1873 4784
rect 2007 4776 2113 4784
rect 3227 4776 3413 4784
rect 3467 4776 3613 4784
rect 3667 4776 3853 4784
rect 4087 4776 4333 4784
rect 4467 4776 4573 4784
rect 4687 4776 4873 4784
rect 5147 4776 5353 4784
rect 5647 4776 5793 4784
rect 1107 4756 1553 4764
rect 1567 4756 1593 4764
rect 2147 4756 2533 4764
rect 3307 4756 3353 4764
rect 3967 4756 4373 4764
rect 4387 4756 4413 4764
rect 4520 4764 4533 4767
rect 4516 4753 4533 4764
rect 4667 4756 4844 4764
rect 107 4736 193 4744
rect 207 4736 213 4744
rect 227 4736 533 4744
rect 547 4736 733 4744
rect 1367 4736 1993 4744
rect 2007 4736 2253 4744
rect 2276 4736 2393 4744
rect 347 4716 573 4724
rect 767 4716 1053 4724
rect 1256 4716 1353 4724
rect 787 4696 1193 4704
rect 1256 4704 1264 4716
rect 1407 4716 1793 4724
rect 2276 4724 2284 4736
rect 2907 4736 3573 4744
rect 3916 4736 4233 4744
rect 2127 4716 2284 4724
rect 2447 4716 3013 4724
rect 3027 4716 3333 4724
rect 3916 4724 3924 4736
rect 4516 4744 4524 4753
rect 4287 4736 4524 4744
rect 4836 4744 4844 4756
rect 4907 4756 6053 4764
rect 4836 4736 5173 4744
rect 5227 4736 5253 4744
rect 5267 4736 5373 4744
rect 3787 4716 3924 4724
rect 3947 4716 4053 4724
rect 4207 4716 4492 4724
rect 4527 4716 4633 4724
rect 4707 4716 5013 4724
rect 1207 4696 1264 4704
rect 1307 4696 1813 4704
rect 1827 4696 2093 4704
rect 2176 4696 2353 4704
rect 487 4676 613 4684
rect 1507 4676 1613 4684
rect 1627 4676 1673 4684
rect 2176 4684 2184 4696
rect 2427 4696 2913 4704
rect 3047 4696 3273 4704
rect 3627 4696 3693 4704
rect 4007 4696 4213 4704
rect 4367 4696 4712 4704
rect 4747 4696 5213 4704
rect 5267 4696 5473 4704
rect 5487 4696 5553 4704
rect 1947 4676 2184 4684
rect 2207 4676 2944 4684
rect 27 4656 773 4664
rect 1227 4656 1293 4664
rect 1747 4656 2333 4664
rect 2407 4656 2693 4664
rect 2936 4664 2944 4676
rect 3567 4676 3653 4684
rect 3667 4676 3693 4684
rect 3927 4676 4333 4684
rect 4627 4676 4813 4684
rect 4887 4676 5653 4684
rect 2936 4656 3073 4664
rect 3287 4656 3993 4664
rect 4107 4656 4193 4664
rect 4507 4656 4613 4664
rect 5367 4656 5633 4664
rect 5907 4656 6093 4664
rect 887 4636 1153 4644
rect 1407 4636 1593 4644
rect 1607 4636 2733 4644
rect 2887 4636 2933 4644
rect 3267 4636 3552 4644
rect 3587 4636 4184 4644
rect 507 4616 973 4624
rect 1727 4616 1892 4624
rect 1927 4616 2184 4624
rect 87 4596 233 4604
rect 1047 4596 1073 4604
rect 2176 4604 2184 4616
rect 2307 4616 2433 4624
rect 3827 4616 4153 4624
rect 4176 4624 4184 4636
rect 4347 4636 4653 4644
rect 5087 4636 5153 4644
rect 5227 4636 5533 4644
rect 5727 4636 5833 4644
rect 4176 4616 4273 4624
rect 4547 4616 4633 4624
rect 5107 4616 5193 4624
rect 5527 4616 5573 4624
rect 5667 4616 5913 4624
rect 2176 4596 2373 4604
rect 2547 4596 2613 4604
rect 2667 4596 2933 4604
rect 3107 4596 3493 4604
rect 3887 4596 4452 4604
rect 4487 4596 4573 4604
rect 4747 4596 4813 4604
rect 4987 4596 5353 4604
rect 5427 4596 5553 4604
rect 747 4576 1084 4584
rect 47 4557 73 4565
rect 127 4557 152 4565
rect 307 4556 393 4564
rect 447 4556 513 4564
rect 567 4556 673 4564
rect 176 4524 184 4553
rect 516 4544 524 4554
rect 716 4544 724 4554
rect 787 4556 813 4564
rect 1047 4564 1060 4567
rect 1076 4564 1084 4576
rect 1147 4576 1213 4584
rect 2167 4576 2213 4584
rect 2967 4576 3013 4584
rect 4396 4576 4513 4584
rect 1047 4553 1064 4564
rect 1076 4556 1224 4564
rect 516 4536 724 4544
rect 1056 4544 1064 4553
rect 1056 4536 1204 4544
rect 176 4516 213 4524
rect 327 4516 373 4524
rect 547 4516 693 4524
rect 607 4496 633 4504
rect 716 4504 724 4536
rect 807 4516 1033 4524
rect 1196 4526 1204 4536
rect 1107 4515 1172 4523
rect 1216 4524 1224 4556
rect 1267 4557 1313 4565
rect 1567 4556 1673 4564
rect 1696 4556 1713 4564
rect 1516 4544 1524 4554
rect 1696 4544 1704 4556
rect 1476 4540 1524 4544
rect 1473 4536 1524 4540
rect 1536 4536 1704 4544
rect 1473 4527 1487 4536
rect 1216 4516 1233 4524
rect 1327 4516 1373 4524
rect 1536 4526 1544 4536
rect 1787 4516 1813 4524
rect 716 4496 893 4504
rect 1836 4504 1844 4554
rect 1887 4556 1953 4564
rect 1967 4557 2053 4565
rect 2367 4557 2813 4565
rect 2827 4556 2893 4564
rect 1907 4516 2113 4524
rect 2136 4524 2144 4554
rect 3056 4556 3093 4564
rect 3056 4544 3064 4556
rect 3167 4556 3233 4564
rect 3327 4556 3613 4564
rect 3747 4557 3813 4565
rect 4027 4556 4113 4564
rect 4160 4564 4173 4567
rect 4156 4553 4173 4564
rect 4267 4557 4293 4565
rect 2467 4536 2704 4544
rect 2136 4516 2173 4524
rect 2696 4524 2704 4536
rect 2996 4536 3064 4544
rect 2696 4516 2833 4524
rect 2847 4516 2913 4524
rect 2996 4524 3004 4536
rect 2967 4516 3004 4524
rect 3027 4515 3073 4523
rect 3787 4516 3833 4524
rect 4156 4507 4164 4553
rect 4396 4544 4404 4576
rect 4647 4576 4713 4584
rect 4907 4576 4953 4584
rect 5113 4576 5313 4584
rect 5113 4568 5127 4576
rect 6147 4584 6160 4587
rect 6147 4573 6164 4584
rect 4467 4556 4564 4564
rect 4376 4536 4404 4544
rect 4556 4544 4564 4556
rect 4587 4556 5024 4564
rect 5016 4547 5024 4556
rect 5067 4557 5113 4565
rect 5360 4564 5373 4567
rect 4556 4540 4584 4544
rect 4556 4536 4587 4540
rect 5016 4536 5033 4547
rect 4376 4526 4384 4536
rect 4573 4527 4587 4536
rect 5020 4533 5033 4536
rect 4207 4515 4233 4523
rect 5156 4527 5164 4554
rect 5276 4527 5284 4554
rect 5356 4553 5373 4564
rect 5356 4527 5364 4553
rect 4707 4515 4953 4523
rect 5156 4516 5173 4527
rect 5160 4513 5173 4516
rect 5267 4516 5284 4527
rect 5267 4513 5280 4516
rect 5436 4524 5444 4573
rect 5467 4556 5493 4564
rect 5627 4556 5644 4564
rect 5636 4527 5644 4556
rect 5436 4516 5473 4524
rect 5716 4507 5724 4573
rect 5947 4556 6064 4564
rect 5893 4544 5907 4553
rect 5893 4540 5924 4544
rect 5896 4536 5924 4540
rect 5916 4526 5924 4536
rect 6056 4526 6064 4556
rect 6087 4557 6133 4565
rect 6156 4544 6164 4573
rect 6116 4540 6164 4544
rect 6113 4536 6164 4540
rect 6113 4527 6127 4536
rect 1747 4496 1844 4504
rect 1907 4496 2193 4504
rect 2367 4496 2813 4504
rect 3147 4496 3173 4504
rect 4007 4496 4132 4504
rect 4607 4496 4653 4504
rect 5007 4496 5053 4504
rect 5407 4496 5533 4504
rect 5847 4496 5873 4504
rect 187 4476 293 4484
rect 827 4476 853 4484
rect 1067 4476 1233 4484
rect 1487 4476 1693 4484
rect 1767 4476 1853 4484
rect 1867 4476 1913 4484
rect 2087 4476 2172 4484
rect 2207 4476 2293 4484
rect 2927 4476 3313 4484
rect 3327 4476 3553 4484
rect 3627 4476 3853 4484
rect 3907 4476 4013 4484
rect 4227 4476 4292 4484
rect 4327 4476 4573 4484
rect 4627 4476 4673 4484
rect 4787 4476 5093 4484
rect 5107 4476 5253 4484
rect 5387 4476 5473 4484
rect 5907 4476 6093 4484
rect 107 4456 413 4464
rect 427 4456 533 4464
rect 587 4456 773 4464
rect 1167 4456 1453 4464
rect 2167 4456 2453 4464
rect 2887 4456 3933 4464
rect 4507 4456 4753 4464
rect 4827 4456 5333 4464
rect 5347 4456 5513 4464
rect 5527 4456 5573 4464
rect 6007 4456 6093 4464
rect 1187 4436 1312 4444
rect 1347 4436 1413 4444
rect 2487 4436 2653 4444
rect 2707 4436 2793 4444
rect 2947 4436 3033 4444
rect 3587 4436 3713 4444
rect 4027 4436 4373 4444
rect 4527 4436 4593 4444
rect 4647 4436 4913 4444
rect 5107 4436 5133 4444
rect 5227 4436 5393 4444
rect 5727 4436 5813 4444
rect 987 4416 1112 4424
rect 1147 4416 1653 4424
rect 1867 4416 1973 4424
rect 2307 4416 2433 4424
rect 2507 4416 2533 4424
rect 2747 4416 3053 4424
rect 3067 4416 3213 4424
rect 3307 4416 3973 4424
rect 4067 4416 4233 4424
rect 4487 4416 4613 4424
rect 4667 4416 4733 4424
rect 5607 4416 5633 4424
rect 5967 4416 6013 4424
rect 6027 4416 6113 4424
rect 627 4396 653 4404
rect 667 4396 873 4404
rect 967 4396 993 4404
rect 1007 4396 1673 4404
rect 1887 4396 2133 4404
rect 2427 4396 2633 4404
rect 2687 4396 2713 4404
rect 2727 4396 2773 4404
rect 3427 4396 3593 4404
rect 3727 4396 3953 4404
rect 4467 4396 4633 4404
rect 4747 4396 4773 4404
rect 4927 4396 5133 4404
rect 5147 4396 5193 4404
rect 5727 4396 5773 4404
rect 247 4376 373 4384
rect 867 4376 1493 4384
rect 1587 4376 1813 4384
rect 2467 4376 2733 4384
rect 2807 4376 2913 4384
rect 3307 4376 3333 4384
rect 3467 4376 3533 4384
rect 4307 4376 4512 4384
rect 4547 4376 4813 4384
rect 5067 4376 5113 4384
rect 5287 4376 5633 4384
rect 5947 4376 6073 4384
rect 307 4356 453 4364
rect 747 4356 793 4364
rect 1107 4356 1153 4364
rect 1207 4356 1333 4364
rect 2007 4364 2020 4367
rect 2007 4353 2024 4364
rect 2447 4356 2693 4364
rect 3967 4356 4073 4364
rect 4407 4356 4553 4364
rect 4607 4356 4693 4364
rect 5007 4356 5033 4364
rect 5667 4356 5724 4364
rect 67 4337 93 4345
rect 167 4336 224 4344
rect 127 4296 173 4304
rect 216 4306 224 4336
rect 256 4324 264 4353
rect 287 4337 312 4345
rect 333 4324 347 4333
rect 476 4336 533 4344
rect 256 4316 324 4324
rect 333 4320 384 4324
rect 336 4316 384 4320
rect 316 4304 324 4316
rect 316 4296 353 4304
rect 376 4304 384 4316
rect 476 4307 484 4336
rect 1187 4336 1204 4344
rect 676 4307 684 4334
rect 1196 4307 1204 4336
rect 1836 4336 1873 4344
rect 1287 4316 1392 4324
rect 376 4296 433 4304
rect 676 4296 693 4307
rect 680 4293 693 4296
rect 827 4295 1013 4303
rect 1067 4295 1093 4303
rect 1196 4296 1213 4307
rect 1200 4293 1213 4296
rect 1413 4304 1427 4313
rect 1413 4300 1633 4304
rect 1416 4296 1633 4300
rect 1776 4304 1784 4334
rect 1836 4306 1844 4336
rect 2016 4344 2024 4353
rect 2016 4336 2353 4344
rect 2696 4336 2753 4344
rect 2416 4307 2424 4333
rect 2696 4307 2704 4336
rect 2807 4344 2820 4347
rect 2807 4333 2824 4344
rect 2907 4336 2933 4344
rect 2976 4336 3373 4344
rect 2816 4307 2824 4333
rect 2976 4307 2984 4336
rect 3427 4336 3493 4344
rect 3560 4344 3573 4347
rect 3556 4333 3573 4344
rect 1727 4296 1784 4304
rect 3556 4306 3564 4333
rect 3636 4307 3644 4353
rect 3696 4307 3704 4334
rect 3636 4296 3653 4307
rect 3640 4293 3653 4296
rect 3696 4296 3713 4307
rect 3700 4293 3713 4296
rect 407 4276 553 4284
rect 567 4276 613 4284
rect 787 4276 933 4284
rect 947 4276 1004 4284
rect 467 4256 513 4264
rect 996 4264 1004 4276
rect 1327 4276 1553 4284
rect 1987 4276 2073 4284
rect 2667 4276 2793 4284
rect 3736 4284 3744 4336
rect 4696 4336 4793 4344
rect 3836 4307 3844 4333
rect 4056 4324 4064 4334
rect 3976 4316 4064 4324
rect 3976 4304 3984 4316
rect 3887 4296 3984 4304
rect 4007 4295 4033 4303
rect 4096 4304 4104 4334
rect 4096 4296 4133 4304
rect 4207 4296 4552 4304
rect 4587 4296 4613 4304
rect 4636 4287 4644 4334
rect 4676 4287 4684 4334
rect 4696 4306 4704 4336
rect 4847 4337 4893 4345
rect 4907 4336 4973 4344
rect 5076 4324 5084 4353
rect 5016 4320 5084 4324
rect 5013 4316 5084 4320
rect 5013 4307 5027 4316
rect 4827 4296 4933 4304
rect 5096 4287 5104 4334
rect 5167 4336 5213 4344
rect 5347 4336 5413 4344
rect 5287 4296 5313 4304
rect 3587 4276 3744 4284
rect 5136 4276 5253 4284
rect 996 4256 1153 4264
rect 1687 4256 1733 4264
rect 2507 4256 2733 4264
rect 3027 4256 3273 4264
rect 3627 4256 3672 4264
rect 3707 4256 3913 4264
rect 3987 4256 4093 4264
rect 4867 4256 4893 4264
rect 4907 4256 4953 4264
rect 5136 4264 5144 4276
rect 5456 4285 5464 4334
rect 5496 4304 5504 4333
rect 5676 4307 5684 4333
rect 5716 4307 5724 4356
rect 5747 4356 5913 4364
rect 5787 4336 5873 4344
rect 5896 4307 5904 4356
rect 5976 4307 5984 4333
rect 5487 4296 5504 4304
rect 5547 4295 5573 4303
rect 5456 4276 5473 4285
rect 5460 4273 5473 4276
rect 5627 4276 5633 4284
rect 5647 4276 5753 4284
rect 5887 4276 5913 4284
rect 5067 4256 5144 4264
rect 5827 4256 5853 4264
rect 607 4236 713 4244
rect 767 4236 1073 4244
rect 1247 4236 1473 4244
rect 1707 4236 1733 4244
rect 1747 4236 1893 4244
rect 2107 4236 2193 4244
rect 3207 4236 3453 4244
rect 4267 4236 4473 4244
rect 5047 4236 5153 4244
rect 5327 4236 5553 4244
rect 5607 4236 5673 4244
rect 5967 4236 6033 4244
rect 1147 4216 1592 4224
rect 1627 4216 1993 4224
rect 2387 4216 2653 4224
rect 2707 4216 2784 4224
rect 667 4196 773 4204
rect 1207 4196 1293 4204
rect 1607 4196 1973 4204
rect 2776 4204 2784 4216
rect 4527 4216 4793 4224
rect 4847 4216 4993 4224
rect 5187 4216 5653 4224
rect 2776 4196 2953 4204
rect 3267 4196 3573 4204
rect 3667 4196 3773 4204
rect 4147 4196 5373 4204
rect 807 4176 913 4184
rect 1127 4176 1333 4184
rect 1587 4176 2533 4184
rect 2716 4176 2873 4184
rect 2716 4167 2724 4176
rect 3647 4176 4193 4184
rect 4807 4176 5053 4184
rect 5527 4176 5573 4184
rect 1547 4156 2264 4164
rect 2256 4147 2264 4156
rect 2587 4156 2713 4164
rect 2907 4156 3013 4164
rect 3116 4156 3713 4164
rect 707 4136 893 4144
rect 907 4136 1093 4144
rect 1107 4136 1213 4144
rect 2267 4136 2433 4144
rect 3116 4144 3124 4156
rect 3807 4156 4013 4164
rect 4247 4156 4733 4164
rect 4807 4156 4933 4164
rect 5696 4156 5893 4164
rect 2447 4136 3124 4144
rect 3607 4136 3653 4144
rect 4647 4136 5073 4144
rect 5407 4136 5433 4144
rect 5696 4144 5704 4156
rect 5547 4136 5704 4144
rect 1667 4116 2053 4124
rect 2067 4116 2113 4124
rect 2187 4116 2253 4124
rect 2267 4116 2364 4124
rect 1087 4096 1253 4104
rect 1267 4096 1373 4104
rect 1447 4096 1713 4104
rect 2356 4104 2364 4116
rect 2647 4116 3253 4124
rect 3527 4116 3673 4124
rect 3687 4116 3813 4124
rect 3827 4116 4073 4124
rect 4187 4116 4233 4124
rect 4327 4116 4453 4124
rect 4467 4116 4553 4124
rect 4647 4116 4673 4124
rect 4947 4116 5013 4124
rect 5227 4116 5353 4124
rect 5767 4116 5793 4124
rect 5807 4116 5953 4124
rect 5967 4116 6033 4124
rect 2356 4096 2473 4104
rect 2707 4096 2833 4104
rect 3327 4096 3493 4104
rect 4367 4096 4653 4104
rect 4887 4096 5133 4104
rect 5147 4096 5173 4104
rect 5487 4096 5793 4104
rect 127 4076 313 4084
rect 327 4076 393 4084
rect 507 4076 753 4084
rect 1807 4076 2293 4084
rect 216 4056 253 4064
rect 167 4037 193 4045
rect 216 4007 224 4056
rect 1347 4056 1433 4064
rect 1616 4056 1733 4064
rect 247 4036 333 4044
rect 347 4036 493 4044
rect 507 4037 533 4045
rect 587 4036 673 4044
rect 1207 4037 1273 4045
rect 1427 4036 1473 4044
rect 787 4016 953 4024
rect 67 3996 93 4004
rect 516 4000 553 4004
rect 513 3996 553 4000
rect 513 3987 527 3996
rect 1307 3996 1493 4004
rect 1616 4004 1624 4056
rect 1887 4056 1913 4064
rect 1647 4036 1813 4044
rect 1836 4036 1913 4044
rect 1836 4024 1844 4036
rect 1936 4024 1944 4076
rect 2347 4076 2673 4084
rect 2867 4076 3293 4084
rect 3307 4076 3333 4084
rect 3767 4076 3913 4084
rect 3927 4076 3973 4084
rect 4027 4076 4113 4084
rect 4387 4076 4413 4084
rect 4987 4076 5073 4084
rect 5627 4076 5753 4084
rect 5796 4084 5804 4092
rect 5796 4076 6093 4084
rect 2147 4056 2213 4064
rect 2487 4056 2613 4064
rect 2627 4056 2653 4064
rect 2736 4056 2813 4064
rect 1987 4037 2053 4045
rect 2167 4036 2213 4044
rect 2227 4036 2333 4044
rect 2633 4024 2647 4033
rect 1796 4016 1844 4024
rect 1896 4016 1944 4024
rect 2536 4020 2647 4024
rect 2736 4024 2744 4056
rect 4067 4056 4207 4064
rect 2767 4036 2853 4044
rect 2867 4036 2933 4044
rect 2536 4016 2644 4020
rect 2736 4016 2844 4024
rect 1796 4006 1804 4016
rect 1896 4006 1904 4016
rect 1567 3996 1624 4004
rect 2107 3996 2353 4004
rect 2536 4004 2544 4016
rect 2836 4006 2844 4016
rect 3176 4007 3184 4036
rect 3236 4024 3244 4036
rect 3236 4016 3293 4024
rect 2367 3996 2544 4004
rect 2587 3995 2693 4003
rect 2747 4000 2784 4004
rect 2747 3996 2787 4000
rect 2773 3987 2787 3996
rect 2887 3996 2913 4004
rect 2927 3996 2973 4004
rect 3167 3996 3184 4007
rect 3356 4006 3364 4053
rect 3376 4007 3384 4034
rect 3527 4036 3553 4044
rect 4193 4048 4207 4056
rect 4227 4056 4284 4064
rect 3627 4036 3693 4044
rect 3616 4007 3624 4036
rect 3847 4037 3873 4045
rect 4207 4037 4253 4045
rect 3167 3993 3180 3996
rect 3376 3996 3393 4007
rect 3380 3993 3393 3996
rect 3447 3993 3493 4001
rect 3616 3996 3633 4007
rect 3620 3993 3633 3996
rect 3747 3996 3833 4004
rect 147 3976 253 3984
rect 727 3976 1013 3984
rect 1716 3976 1773 3984
rect 487 3956 673 3964
rect 1267 3956 1393 3964
rect 1467 3956 1573 3964
rect 1716 3964 1724 3976
rect 3956 3984 3964 4033
rect 4076 4004 4084 4033
rect 4136 4007 4144 4033
rect 4047 3996 4084 4004
rect 4276 4004 4284 4056
rect 5127 4056 5153 4064
rect 5387 4056 5533 4064
rect 5956 4056 6084 4064
rect 4607 4036 4693 4044
rect 4767 4036 4833 4044
rect 4856 4036 4893 4044
rect 4396 4007 4404 4033
rect 4856 4024 4864 4036
rect 5236 4036 5253 4044
rect 4836 4016 4864 4024
rect 4227 3996 4284 4004
rect 4327 3995 4353 4003
rect 4587 3996 4613 4004
rect 4727 3995 4753 4003
rect 4836 3987 4844 4016
rect 5236 4007 5244 4036
rect 5396 4040 5613 4044
rect 5393 4036 5613 4040
rect 5393 4026 5407 4036
rect 5807 4036 5824 4044
rect 5736 4007 5744 4033
rect 5816 4007 5824 4036
rect 5956 4044 5964 4056
rect 6076 4047 6084 4056
rect 5927 4036 5964 4044
rect 5987 4044 6000 4047
rect 5987 4033 6004 4044
rect 5107 3995 5133 4003
rect 5607 3996 5693 4004
rect 5916 4004 5924 4033
rect 5887 3996 5924 4004
rect 5996 4004 6004 4033
rect 6013 4024 6027 4033
rect 6013 4020 6064 4024
rect 6016 4016 6064 4020
rect 6056 4006 6064 4016
rect 5996 4000 6044 4004
rect 5996 3996 6047 4000
rect 6033 3987 6047 3996
rect 6136 4004 6144 4053
rect 6136 3996 6164 4004
rect 3867 3976 3964 3984
rect 4007 3976 4093 3984
rect 4647 3976 4673 3984
rect 1627 3956 1724 3964
rect 1807 3956 1833 3964
rect 1987 3956 2093 3964
rect 2147 3956 2873 3964
rect 3307 3956 3413 3964
rect 3427 3956 3633 3964
rect 3647 3956 4553 3964
rect 4607 3956 4853 3964
rect 5127 3956 5273 3964
rect 5787 3956 5873 3964
rect 5947 3956 6133 3964
rect 27 3936 413 3944
rect 507 3936 693 3944
rect 827 3936 873 3944
rect 1007 3936 1193 3944
rect 1247 3936 1413 3944
rect 1607 3936 1773 3944
rect 1867 3936 2033 3944
rect 3436 3940 3493 3944
rect 3433 3936 3493 3940
rect 3433 3927 3447 3936
rect 3847 3936 4413 3944
rect 4667 3936 4793 3944
rect 4887 3936 5093 3944
rect 5847 3936 5973 3944
rect 6156 3927 6164 3996
rect 127 3916 333 3924
rect 687 3916 853 3924
rect 896 3916 1753 3924
rect 167 3896 273 3904
rect 287 3896 753 3904
rect 896 3904 904 3916
rect 2247 3916 2664 3924
rect 2656 3907 2664 3916
rect 3307 3916 3393 3924
rect 3527 3916 3893 3924
rect 3947 3916 4213 3924
rect 4927 3916 5013 3924
rect 5227 3916 5253 3924
rect 6067 3916 6093 3924
rect 6147 3916 6164 3927
rect 6147 3913 6160 3916
rect 767 3896 904 3904
rect 1047 3896 1113 3904
rect 1187 3896 1273 3904
rect 1607 3896 1633 3904
rect 1647 3896 1693 3904
rect 2547 3896 2613 3904
rect 2667 3896 2933 3904
rect 3127 3896 3193 3904
rect 3427 3896 3453 3904
rect 3627 3896 3673 3904
rect 4187 3896 4213 3904
rect 4916 3904 4924 3913
rect 4447 3896 4924 3904
rect 5107 3896 5273 3904
rect 387 3876 513 3884
rect 527 3876 833 3884
rect 1447 3876 1533 3884
rect 1767 3876 1893 3884
rect 2187 3876 2273 3884
rect 2767 3876 2913 3884
rect 3227 3876 3473 3884
rect 4627 3876 4893 3884
rect 5087 3876 5293 3884
rect 5647 3876 5793 3884
rect 6027 3876 6073 3884
rect 907 3856 1153 3864
rect 1287 3856 1513 3864
rect 1647 3856 1693 3864
rect 1747 3856 1853 3864
rect 1927 3856 2013 3864
rect 2567 3856 2613 3864
rect 2707 3856 2793 3864
rect 2807 3856 3033 3864
rect 3087 3856 3133 3864
rect 3207 3856 3544 3864
rect 67 3836 253 3844
rect 267 3836 413 3844
rect 607 3836 633 3844
rect 647 3836 813 3844
rect 2227 3836 2253 3844
rect 2487 3836 2513 3844
rect 2727 3836 2793 3844
rect 307 3816 353 3824
rect 587 3816 604 3824
rect 67 3775 93 3783
rect 196 3784 204 3813
rect 596 3787 604 3816
rect 720 3824 733 3827
rect 716 3813 733 3824
rect 856 3816 913 3824
rect 196 3776 253 3784
rect 407 3776 513 3784
rect 527 3775 553 3783
rect 596 3776 613 3787
rect 600 3773 613 3776
rect 656 3784 664 3813
rect 716 3786 724 3813
rect 856 3787 864 3816
rect 967 3816 1093 3824
rect 1147 3816 1304 3824
rect 656 3776 673 3784
rect 767 3775 793 3783
rect 907 3775 933 3783
rect 947 3776 1053 3784
rect 1296 3786 1304 3816
rect 1316 3787 1324 3814
rect 1507 3816 1553 3824
rect 1576 3816 1633 3824
rect 1576 3804 1584 3816
rect 1687 3824 1700 3827
rect 1687 3813 1704 3824
rect 1367 3796 1584 3804
rect 1227 3775 1253 3783
rect 1316 3776 1333 3787
rect 1320 3773 1333 3776
rect 1447 3775 1513 3783
rect 1587 3775 1673 3783
rect 713 3764 727 3772
rect 387 3756 727 3764
rect 1127 3756 1173 3764
rect 1696 3765 1704 3813
rect 1716 3804 1724 3833
rect 2807 3836 2893 3844
rect 3007 3836 3053 3844
rect 3327 3836 3493 3844
rect 1773 3804 1787 3813
rect 1716 3796 1744 3804
rect 1773 3800 1804 3804
rect 1776 3796 1804 3800
rect 1736 3784 1744 3796
rect 1736 3776 1773 3784
rect 1796 3784 1804 3796
rect 1796 3776 1833 3784
rect 1896 3784 1904 3813
rect 1947 3817 1973 3825
rect 1987 3816 2193 3824
rect 2367 3816 2444 3824
rect 2233 3804 2247 3813
rect 2216 3800 2247 3804
rect 2216 3796 2244 3800
rect 2216 3786 2224 3796
rect 2335 3787 2343 3813
rect 1896 3776 1993 3784
rect 2007 3775 2192 3783
rect 2287 3776 2312 3784
rect 1716 3764 1724 3772
rect 2436 3767 2444 3816
rect 2607 3816 2633 3824
rect 2456 3784 2464 3813
rect 2696 3787 2704 3813
rect 2456 3776 2493 3784
rect 2807 3775 2833 3783
rect 2856 3767 2864 3814
rect 2967 3816 3093 3824
rect 3213 3804 3227 3813
rect 2916 3800 3227 3804
rect 3376 3816 3433 3824
rect 2916 3796 3224 3800
rect 2916 3767 2924 3796
rect 3376 3787 3384 3816
rect 3536 3824 3544 3856
rect 3887 3856 4073 3864
rect 5027 3856 5233 3864
rect 5427 3856 5473 3864
rect 5547 3856 5593 3864
rect 5787 3856 5833 3864
rect 5907 3856 5933 3864
rect 3667 3836 3733 3844
rect 5287 3836 5493 3844
rect 5616 3836 5653 3844
rect 3527 3816 3544 3824
rect 3687 3816 3752 3824
rect 3896 3816 3933 3824
rect 2947 3775 2973 3783
rect 3027 3776 3173 3784
rect 3327 3776 3352 3784
rect 3427 3773 3453 3781
rect 3776 3784 3784 3813
rect 3507 3776 3784 3784
rect 3816 3784 3824 3813
rect 3856 3787 3864 3813
rect 3896 3787 3904 3816
rect 4113 3827 4127 3833
rect 4027 3819 4153 3827
rect 4116 3816 4124 3819
rect 4427 3817 4493 3825
rect 4253 3804 4267 3813
rect 3807 3776 3824 3784
rect 3993 3784 4007 3793
rect 3967 3780 4007 3784
rect 4196 3800 4267 3804
rect 4196 3796 4264 3800
rect 3967 3776 4004 3780
rect 4196 3767 4204 3796
rect 4556 3784 4564 3813
rect 5096 3804 5104 3814
rect 5387 3816 5444 3824
rect 5036 3796 5104 3804
rect 5436 3804 5444 3816
rect 5467 3817 5513 3825
rect 5436 3800 5584 3804
rect 5436 3796 5587 3800
rect 4227 3773 4273 3781
rect 4556 3776 4573 3784
rect 4727 3775 4893 3783
rect 5036 3784 5044 3796
rect 5573 3787 5587 3796
rect 4947 3776 5044 3784
rect 5067 3776 5253 3784
rect 5616 3786 5624 3836
rect 5727 3836 5853 3844
rect 6047 3836 6093 3844
rect 5747 3816 5784 3824
rect 5776 3767 5784 3816
rect 5796 3816 5893 3824
rect 5796 3786 5804 3816
rect 5967 3816 5993 3824
rect 6056 3787 6064 3813
rect 1716 3756 1913 3764
rect 2047 3756 2093 3764
rect 2107 3756 2153 3764
rect 2227 3756 2373 3764
rect 2436 3756 2453 3767
rect 2440 3753 2453 3756
rect 2567 3756 2653 3764
rect 2907 3756 2924 3767
rect 2907 3753 2920 3756
rect 3107 3756 3213 3764
rect 3487 3756 3653 3764
rect 4196 3766 4220 3767
rect 4196 3756 4213 3766
rect 4200 3753 4213 3756
rect 4407 3756 4453 3764
rect 4947 3756 5313 3764
rect 187 3736 313 3744
rect 327 3736 833 3744
rect 847 3736 1353 3744
rect 1407 3736 1533 3744
rect 1687 3736 1753 3744
rect 1807 3736 1833 3744
rect 2307 3736 2333 3744
rect 2407 3736 2573 3744
rect 3187 3736 3313 3744
rect 3587 3736 3753 3744
rect 4507 3736 4653 3744
rect 5027 3736 5133 3744
rect 5287 3736 5353 3744
rect 5427 3736 5513 3744
rect 5527 3736 5653 3744
rect 5867 3736 5913 3744
rect 607 3716 673 3724
rect 687 3716 893 3724
rect 1047 3716 1153 3724
rect 1787 3716 2092 3724
rect 2127 3716 2313 3724
rect 4107 3716 4233 3724
rect 4427 3716 4453 3724
rect 4567 3716 4633 3724
rect 5167 3716 5473 3724
rect 1627 3696 1793 3704
rect 1847 3696 1953 3704
rect 1967 3696 2024 3704
rect 1007 3676 1533 3684
rect 1547 3676 1813 3684
rect 2016 3684 2024 3696
rect 2147 3696 2333 3704
rect 2547 3696 2793 3704
rect 3007 3696 3193 3704
rect 3707 3696 4013 3704
rect 4667 3696 5073 3704
rect 2016 3676 2413 3684
rect 2427 3676 2893 3684
rect 3047 3676 3353 3684
rect 3907 3676 4053 3684
rect 5047 3676 5153 3684
rect 6027 3676 6113 3684
rect 707 3656 873 3664
rect 1667 3656 1713 3664
rect 1887 3656 2144 3664
rect 1267 3636 1644 3644
rect 27 3616 333 3624
rect 347 3616 433 3624
rect 1636 3624 1644 3636
rect 1667 3636 1973 3644
rect 2136 3644 2144 3656
rect 2167 3656 2433 3664
rect 2927 3656 3273 3664
rect 3327 3656 3564 3664
rect 2136 3636 2352 3644
rect 2387 3636 2633 3644
rect 2747 3636 3053 3644
rect 3187 3636 3253 3644
rect 3556 3644 3564 3656
rect 4167 3656 4353 3664
rect 4367 3656 5013 3664
rect 5267 3656 5593 3664
rect 5887 3656 6093 3664
rect 3556 3636 3893 3644
rect 4347 3636 4493 3644
rect 4547 3636 4773 3644
rect 6047 3636 6113 3644
rect 1636 3616 1733 3624
rect 1967 3616 2473 3624
rect 2887 3616 3333 3624
rect 3387 3616 3493 3624
rect 3547 3616 3613 3624
rect 3627 3616 4253 3624
rect 5027 3616 5213 3624
rect 5227 3616 5253 3624
rect 5747 3616 5853 3624
rect 207 3596 753 3604
rect 967 3596 1073 3604
rect 1187 3596 1233 3604
rect 1567 3596 1613 3604
rect 1767 3596 1893 3604
rect 2447 3596 2493 3604
rect 2667 3596 3172 3604
rect 3207 3596 3233 3604
rect 3667 3596 4513 3604
rect 4647 3596 4793 3604
rect 4907 3596 5273 3604
rect 5567 3596 5713 3604
rect 5947 3596 6093 3604
rect 287 3576 353 3584
rect 1387 3576 1553 3584
rect 1747 3576 1913 3584
rect 2207 3576 2273 3584
rect 2287 3576 2373 3584
rect 2867 3576 3013 3584
rect 4187 3576 4373 3584
rect 5587 3576 5793 3584
rect 616 3556 673 3564
rect 616 3547 624 3556
rect 787 3556 953 3564
rect 1027 3556 1113 3564
rect 1207 3556 1253 3564
rect 1307 3556 1333 3564
rect 1347 3556 1573 3564
rect 1756 3556 1853 3564
rect 547 3536 613 3544
rect 1756 3544 1764 3556
rect 3087 3556 3153 3564
rect 3227 3556 3573 3564
rect 4487 3556 4533 3564
rect 4707 3556 4893 3564
rect 5127 3556 5293 3564
rect 5907 3556 6073 3564
rect 1727 3536 1764 3544
rect 2587 3536 2753 3544
rect 2767 3536 2873 3544
rect 3707 3536 3733 3544
rect 3887 3536 4073 3544
rect 5187 3536 5293 3544
rect 5307 3536 5433 3544
rect 5447 3536 5553 3544
rect 6020 3544 6033 3547
rect 6016 3533 6033 3544
rect 147 3516 233 3524
rect 447 3517 493 3525
rect 536 3516 633 3524
rect 536 3504 544 3516
rect 847 3517 913 3525
rect 516 3496 544 3504
rect 67 3474 73 3482
rect 87 3474 93 3482
rect 367 3476 433 3484
rect 516 3486 524 3496
rect 676 3487 684 3513
rect 736 3504 744 3514
rect 1267 3516 1393 3524
rect 1587 3516 1673 3524
rect 736 3496 884 3504
rect 876 3487 884 3496
rect 807 3476 833 3484
rect 876 3476 893 3487
rect 880 3473 893 3476
rect 996 3484 1004 3513
rect 947 3476 1004 3484
rect 1436 3487 1444 3514
rect 1556 3496 1733 3504
rect 1436 3476 1453 3487
rect 1440 3473 1453 3476
rect 1556 3486 1564 3496
rect 1776 3484 1784 3514
rect 2047 3516 2233 3524
rect 2367 3516 2404 3524
rect 1893 3504 1907 3513
rect 1893 3500 1984 3504
rect 1896 3496 1984 3500
rect 1667 3476 1784 3484
rect 1847 3476 1953 3484
rect 1976 3484 1984 3496
rect 2296 3487 2304 3513
rect 1976 3476 2133 3484
rect 2396 3486 2404 3516
rect 2967 3517 2993 3525
rect 2413 3504 2427 3513
rect 2413 3500 2484 3504
rect 2416 3496 2487 3500
rect 2473 3487 2487 3496
rect 2556 3484 2564 3513
rect 2587 3496 2833 3504
rect 2853 3504 2867 3513
rect 2853 3500 2904 3504
rect 2856 3496 2904 3500
rect 2556 3476 2593 3484
rect 2896 3486 2904 3496
rect 3116 3484 3124 3514
rect 3153 3504 3167 3513
rect 3153 3500 3184 3504
rect 3156 3496 3187 3500
rect 3173 3487 3187 3496
rect 3116 3476 3152 3484
rect 3196 3467 3204 3514
rect 3447 3517 3493 3525
rect 3547 3516 3633 3524
rect 3767 3516 3793 3524
rect 3256 3487 3264 3513
rect 3336 3504 3344 3514
rect 3296 3500 3344 3504
rect 3293 3496 3344 3500
rect 3293 3487 3307 3496
rect 3376 3467 3384 3514
rect 4247 3516 4373 3524
rect 4387 3516 4493 3524
rect 4767 3516 4993 3524
rect 5207 3516 5264 3524
rect 3933 3504 3947 3513
rect 3456 3496 3964 3504
rect 3456 3484 3464 3496
rect 3407 3476 3464 3484
rect 3487 3475 3573 3483
rect 3667 3475 3693 3483
rect 3707 3476 3773 3484
rect 3956 3484 3964 3496
rect 4027 3496 4364 3504
rect 4356 3484 4364 3496
rect 4356 3476 4393 3484
rect 4556 3484 4564 3513
rect 4487 3476 4564 3484
rect 4676 3484 4684 3513
rect 5033 3504 5047 3513
rect 5033 3500 5064 3504
rect 5036 3496 5064 3500
rect 4676 3476 5012 3484
rect 5056 3484 5064 3496
rect 5156 3487 5164 3513
rect 5256 3487 5264 3516
rect 5547 3516 5584 3524
rect 5393 3504 5407 3513
rect 5393 3500 5544 3504
rect 5396 3496 5547 3500
rect 5533 3487 5547 3496
rect 5307 3475 5373 3483
rect 5576 3486 5584 3516
rect 5787 3516 5813 3524
rect 5696 3487 5704 3513
rect 167 3456 233 3464
rect 247 3456 653 3464
rect 867 3456 973 3464
rect 987 3456 1033 3464
rect 1727 3456 1773 3464
rect 2067 3456 2113 3464
rect 2527 3456 2973 3464
rect 3287 3456 3313 3464
rect 4047 3456 4073 3464
rect 4427 3456 4533 3464
rect 4647 3456 4693 3464
rect 5507 3456 5593 3464
rect 47 3436 593 3444
rect 887 3436 913 3444
rect 1107 3436 1273 3444
rect 1287 3436 1413 3444
rect 1467 3436 1653 3444
rect 1747 3436 1793 3444
rect 1847 3436 1873 3444
rect 2147 3436 2253 3444
rect 2267 3436 2573 3444
rect 2827 3436 2993 3444
rect 3167 3436 3213 3444
rect 3587 3436 3733 3444
rect 4447 3436 4793 3444
rect 5427 3436 5653 3444
rect 5736 3444 5744 3514
rect 5967 3516 5993 3524
rect 5876 3487 5884 3513
rect 6016 3504 6024 3533
rect 5976 3496 6024 3504
rect 6076 3516 6113 3524
rect 5767 3475 5793 3483
rect 5976 3484 5984 3496
rect 6076 3486 6084 3516
rect 5936 3480 5984 3484
rect 5933 3476 5984 3480
rect 5933 3467 5947 3476
rect 5736 3436 5913 3444
rect 647 3416 692 3424
rect 727 3416 893 3424
rect 1947 3416 2033 3424
rect 2287 3416 2633 3424
rect 2787 3416 3133 3424
rect 3267 3416 3433 3424
rect 3847 3416 4053 3424
rect 5287 3416 5393 3424
rect 5467 3416 5713 3424
rect 5787 3416 5833 3424
rect 127 3396 753 3404
rect 867 3396 1013 3404
rect 1167 3396 1373 3404
rect 1487 3396 2013 3404
rect 2087 3396 2213 3404
rect 2267 3396 2513 3404
rect 2947 3396 3113 3404
rect 3127 3396 3193 3404
rect 3207 3396 3473 3404
rect 3927 3396 4413 3404
rect 4527 3396 4813 3404
rect 5087 3396 5133 3404
rect 5267 3396 5433 3404
rect 5527 3396 5553 3404
rect 1547 3376 1613 3384
rect 1907 3376 1993 3384
rect 2327 3376 2372 3384
rect 2407 3376 2433 3384
rect 2567 3376 2733 3384
rect 2907 3376 3013 3384
rect 3267 3376 3293 3384
rect 4227 3376 4573 3384
rect 5267 3376 5333 3384
rect 5347 3376 5453 3384
rect 5727 3376 5753 3384
rect 5867 3376 6013 3384
rect 387 3356 533 3364
rect 767 3356 993 3364
rect 1047 3356 1113 3364
rect 1167 3356 1233 3364
rect 1247 3356 1873 3364
rect 2027 3356 2253 3364
rect 2467 3356 2533 3364
rect 2727 3356 2773 3364
rect 2847 3356 3284 3364
rect 427 3336 473 3344
rect 627 3336 713 3344
rect 1267 3336 1553 3344
rect 1627 3336 1753 3344
rect 2027 3336 2193 3344
rect 2207 3336 2273 3344
rect 2347 3336 2493 3344
rect 2567 3336 2593 3344
rect 2607 3336 2673 3344
rect 2927 3336 2973 3344
rect 2987 3336 3073 3344
rect 3147 3336 3213 3344
rect 3276 3344 3284 3356
rect 3876 3356 3993 3364
rect 3876 3347 3884 3356
rect 4787 3356 4893 3364
rect 5047 3356 5133 3364
rect 5587 3356 5633 3364
rect 3276 3336 3393 3344
rect 3807 3336 3873 3344
rect 4427 3336 4473 3344
rect 4487 3336 4733 3344
rect 5227 3336 5313 3344
rect 5627 3336 5713 3344
rect 5847 3336 5873 3344
rect 6067 3336 6113 3344
rect 207 3316 233 3324
rect 1127 3316 1153 3324
rect 1667 3316 1713 3324
rect 1807 3316 1904 3324
rect 47 3296 73 3304
rect 96 3296 153 3304
rect 96 3266 104 3296
rect 287 3296 373 3304
rect 587 3296 713 3304
rect 727 3296 764 3304
rect 356 3276 453 3284
rect 356 3266 364 3276
rect 756 3284 764 3296
rect 787 3297 813 3305
rect 907 3296 1024 3304
rect 756 3276 784 3284
rect 307 3256 353 3264
rect 407 3256 553 3264
rect 627 3255 693 3263
rect 776 3264 784 3276
rect 776 3256 873 3264
rect 887 3256 973 3264
rect 1016 3264 1024 3296
rect 1307 3296 1353 3304
rect 1376 3296 1433 3304
rect 1173 3284 1187 3293
rect 1376 3284 1384 3296
rect 1173 3280 1224 3284
rect 1176 3276 1227 3280
rect 1213 3267 1227 3276
rect 1016 3256 1133 3264
rect 1316 3276 1384 3284
rect 1476 3284 1484 3294
rect 1527 3296 1653 3304
rect 1896 3304 1904 3316
rect 2067 3324 2080 3327
rect 2067 3313 2084 3324
rect 2167 3316 2244 3324
rect 1896 3296 1913 3304
rect 1967 3297 2013 3305
rect 1476 3276 1604 3284
rect 1316 3266 1324 3276
rect 1507 3256 1573 3264
rect 1596 3264 1604 3276
rect 1776 3267 1784 3293
rect 1836 3267 1844 3293
rect 2076 3267 2084 3313
rect 2147 3296 2184 3304
rect 2176 3267 2184 3296
rect 2236 3267 2244 3316
rect 2767 3316 2813 3324
rect 3107 3316 3193 3324
rect 3447 3316 3493 3324
rect 3507 3316 3553 3324
rect 3627 3316 3693 3324
rect 3747 3316 3933 3324
rect 4107 3316 4173 3324
rect 4387 3316 4453 3324
rect 4467 3316 4553 3324
rect 4627 3316 4833 3324
rect 4887 3316 4913 3324
rect 5507 3324 5520 3327
rect 5507 3314 5524 3324
rect 5500 3313 5524 3314
rect 5767 3316 5893 3324
rect 6047 3324 6060 3327
rect 6047 3313 6064 3324
rect 2387 3296 2433 3304
rect 2607 3296 2684 3304
rect 2476 3267 2484 3293
rect 2553 3284 2567 3293
rect 2553 3280 2584 3284
rect 2556 3276 2584 3280
rect 1596 3256 1673 3264
rect 1907 3256 1993 3264
rect 2576 3266 2584 3276
rect 2676 3267 2684 3296
rect 2696 3264 2704 3313
rect 2747 3296 2804 3304
rect 2796 3284 2804 3296
rect 2873 3304 2887 3313
rect 2847 3300 2887 3304
rect 2847 3296 2884 3300
rect 2987 3296 3144 3304
rect 2796 3276 2824 3284
rect 2696 3256 2733 3264
rect 2816 3266 2824 3276
rect 3136 3266 3144 3296
rect 3307 3296 3413 3304
rect 2867 3256 2953 3264
rect 3227 3255 3273 3263
rect 1313 3247 1327 3252
rect 727 3236 833 3244
rect 1307 3233 1327 3247
rect 2027 3236 2053 3244
rect 2147 3236 2193 3244
rect 2587 3236 2613 3244
rect 2853 3244 2867 3252
rect 3296 3247 3304 3294
rect 3487 3296 3684 3304
rect 3447 3255 3493 3263
rect 3587 3256 3613 3264
rect 3676 3266 3684 3296
rect 3736 3296 3833 3304
rect 2787 3236 2867 3244
rect 2907 3236 3233 3244
rect 3736 3244 3744 3296
rect 4047 3296 4153 3304
rect 4207 3296 4232 3304
rect 4267 3297 4293 3305
rect 4487 3296 4504 3304
rect 4356 3267 4364 3293
rect 3787 3255 3853 3263
rect 3907 3255 3933 3263
rect 3947 3256 4013 3264
rect 4127 3255 4173 3263
rect 4267 3256 4313 3264
rect 4496 3264 4504 3296
rect 4496 3256 4553 3264
rect 3667 3236 3744 3244
rect 3853 3244 3867 3252
rect 3853 3236 3973 3244
rect 4347 3236 4393 3244
rect 4576 3244 4584 3294
rect 4827 3296 4973 3304
rect 5047 3296 5153 3304
rect 5176 3296 5313 3304
rect 5176 3284 5184 3296
rect 5447 3296 5493 3304
rect 4976 3276 5184 3284
rect 4607 3256 4753 3264
rect 4767 3256 4933 3264
rect 4976 3247 4984 3276
rect 5516 3266 5524 3313
rect 5667 3297 5733 3305
rect 5576 3267 5584 3293
rect 5796 3267 5804 3293
rect 5027 3256 5353 3264
rect 5367 3256 5473 3264
rect 5936 3247 5944 3313
rect 5956 3267 5964 3313
rect 6016 3267 6024 3293
rect 6056 3247 6064 3313
rect 4447 3236 4584 3244
rect 5707 3236 5773 3244
rect 5827 3236 5873 3244
rect 6047 3244 6064 3247
rect 6047 3236 6093 3244
rect 6047 3233 6060 3236
rect 147 3216 193 3224
rect 207 3216 253 3224
rect 607 3216 944 3224
rect 847 3196 913 3204
rect 936 3204 944 3216
rect 1067 3216 1193 3224
rect 1727 3216 2073 3224
rect 2407 3216 2433 3224
rect 2727 3216 2873 3224
rect 2947 3216 3013 3224
rect 3027 3216 3093 3224
rect 3527 3216 3833 3224
rect 4007 3216 4113 3224
rect 4167 3216 4373 3224
rect 4567 3216 4633 3224
rect 4707 3216 4773 3224
rect 5007 3216 5033 3224
rect 5247 3216 5273 3224
rect 5387 3216 5633 3224
rect 5907 3216 5993 3224
rect 936 3196 1253 3204
rect 1507 3196 1653 3204
rect 1747 3196 1793 3204
rect 1807 3196 2053 3204
rect 2127 3196 2233 3204
rect 2287 3196 2313 3204
rect 2707 3196 2853 3204
rect 3047 3196 3273 3204
rect 3387 3196 3433 3204
rect 4687 3196 4753 3204
rect 5147 3196 5593 3204
rect 5927 3196 6113 3204
rect 487 3176 713 3184
rect 1687 3176 2173 3184
rect 2327 3176 2353 3184
rect 2527 3176 2893 3184
rect 3147 3176 3253 3184
rect 3847 3176 4073 3184
rect 4227 3176 4873 3184
rect 4967 3176 5193 3184
rect 5327 3176 5393 3184
rect 5447 3176 5553 3184
rect 5667 3176 5793 3184
rect 5807 3176 5873 3184
rect 327 3156 433 3164
rect 447 3156 773 3164
rect 787 3156 1353 3164
rect 2027 3156 2153 3164
rect 2167 3156 2253 3164
rect 2607 3156 2773 3164
rect 2787 3156 2813 3164
rect 2947 3156 3313 3164
rect 3327 3156 3393 3164
rect 4127 3156 4893 3164
rect 4947 3156 5093 3164
rect 5347 3156 5753 3164
rect 6007 3156 6073 3164
rect 6087 3156 6113 3164
rect 1427 3136 1633 3144
rect 1707 3136 1853 3144
rect 1867 3136 2373 3144
rect 2467 3136 3033 3144
rect 3087 3136 3833 3144
rect 4367 3136 4513 3144
rect 5367 3136 5573 3144
rect 187 3116 393 3124
rect 967 3116 1013 3124
rect 1467 3116 1713 3124
rect 1967 3116 2213 3124
rect 2587 3116 2633 3124
rect 2687 3116 2833 3124
rect 2887 3116 3053 3124
rect 3267 3116 3713 3124
rect 4067 3116 4413 3124
rect 4507 3116 4793 3124
rect 4927 3116 5053 3124
rect 5867 3116 5893 3124
rect 1687 3096 1844 3104
rect 807 3076 1013 3084
rect 1627 3076 1753 3084
rect 1836 3084 1844 3096
rect 1867 3096 1913 3104
rect 2147 3096 2313 3104
rect 2427 3096 2473 3104
rect 2767 3096 3133 3104
rect 3187 3096 3593 3104
rect 3807 3096 4013 3104
rect 4027 3096 4213 3104
rect 4867 3096 5073 3104
rect 5127 3096 5553 3104
rect 5767 3096 5893 3104
rect 1836 3076 2193 3084
rect 2847 3076 2993 3084
rect 3827 3076 4133 3084
rect 4327 3076 4653 3084
rect 4667 3076 4973 3084
rect 5167 3076 5413 3084
rect 5427 3076 5573 3084
rect 507 3056 753 3064
rect 1387 3056 1672 3064
rect 1707 3056 1773 3064
rect 2087 3056 2273 3064
rect 2407 3056 2633 3064
rect 2927 3056 3033 3064
rect 3247 3056 3533 3064
rect 4007 3056 4173 3064
rect 4307 3056 4393 3064
rect 5067 3056 5513 3064
rect 5567 3056 5793 3064
rect 5947 3056 6033 3064
rect 6147 3064 6160 3067
rect 6147 3053 6164 3064
rect 756 3044 764 3053
rect 756 3036 913 3044
rect 1336 3036 1613 3044
rect 367 3016 593 3024
rect 607 3016 713 3024
rect 1336 3024 1344 3036
rect 1907 3036 1933 3044
rect 1947 3036 1993 3044
rect 2047 3036 2173 3044
rect 2187 3036 2293 3044
rect 2487 3036 2693 3044
rect 2907 3036 3172 3044
rect 3207 3036 3453 3044
rect 3887 3036 4133 3044
rect 4247 3036 4273 3044
rect 4647 3036 4873 3044
rect 4987 3036 5013 3044
rect 5407 3036 5453 3044
rect 5887 3036 6053 3044
rect 1107 3016 1344 3024
rect 1741 3016 1813 3024
rect 2300 3024 2313 3027
rect 2296 3013 2313 3024
rect 2987 3016 3107 3024
rect 147 2997 173 3005
rect 227 2997 273 3005
rect 527 2997 553 3005
rect 620 3004 633 3007
rect 616 2993 633 3004
rect 687 2996 792 3004
rect 827 2997 873 3005
rect 940 3004 953 3007
rect 936 2993 953 3004
rect 1187 2996 1313 3004
rect 1416 2996 1453 3004
rect 616 2984 624 2993
rect 576 2976 624 2984
rect 47 2955 73 2963
rect 127 2956 293 2964
rect 307 2956 413 2964
rect 467 2956 493 2964
rect 576 2966 584 2976
rect 936 2966 944 2993
rect 1047 2956 1093 2964
rect 647 2936 813 2944
rect 933 2944 947 2952
rect 867 2936 947 2944
rect 1136 2944 1144 2994
rect 1416 2984 1424 2996
rect 1507 2996 1524 3004
rect 1356 2976 1424 2984
rect 1356 2964 1364 2976
rect 1516 2967 1524 2996
rect 1693 2984 1707 2993
rect 1676 2980 1707 2984
rect 1896 2996 1933 3004
rect 1676 2976 1704 2980
rect 1207 2956 1364 2964
rect 1387 2956 1433 2964
rect 1676 2964 1684 2976
rect 1587 2956 1684 2964
rect 1896 2964 1904 2996
rect 2100 3004 2113 3007
rect 2096 2993 2113 3004
rect 2296 3004 2304 3013
rect 2256 2996 2304 3004
rect 1707 2956 1904 2964
rect 2016 2964 2024 2993
rect 2096 2967 2104 2993
rect 2236 2984 2244 2994
rect 2136 2980 2244 2984
rect 2133 2976 2244 2980
rect 2133 2967 2147 2976
rect 1927 2956 2072 2964
rect 2256 2964 2264 2996
rect 2653 3004 2667 3013
rect 3093 3008 3107 3016
rect 3327 3016 3353 3024
rect 4427 3016 4464 3024
rect 2576 3000 2667 3004
rect 2576 2996 2664 3000
rect 2336 2984 2344 2994
rect 2576 2984 2584 2996
rect 2733 2984 2747 2993
rect 2316 2976 2344 2984
rect 2376 2980 2584 2984
rect 2373 2976 2584 2980
rect 2616 2980 2747 2984
rect 2616 2976 2744 2980
rect 2216 2956 2264 2964
rect 2216 2947 2224 2956
rect 2316 2964 2324 2976
rect 2287 2956 2324 2964
rect 2373 2967 2387 2976
rect 2616 2964 2624 2976
rect 2527 2956 2624 2964
rect 2636 2956 2693 2964
rect 2636 2947 2644 2956
rect 2776 2964 2784 2994
rect 2827 2996 2864 3004
rect 2856 2984 2864 2996
rect 2916 2996 2993 3004
rect 2856 2980 2884 2984
rect 2856 2976 2887 2980
rect 2873 2967 2887 2976
rect 2776 2956 2833 2964
rect 2916 2966 2924 2996
rect 3107 2996 3144 3004
rect 3136 2984 3144 2996
rect 3167 2997 3193 3005
rect 3247 2996 3373 3004
rect 3507 2996 3693 3004
rect 3707 2997 3813 3005
rect 3947 2999 3973 3007
rect 4247 2996 4353 3004
rect 4036 2984 4044 2994
rect 3136 2976 3224 2984
rect 3216 2966 3224 2976
rect 3976 2976 4044 2984
rect 3047 2955 3073 2963
rect 3267 2956 3293 2964
rect 3467 2955 3513 2963
rect 3607 2955 3633 2963
rect 3976 2964 3984 2976
rect 4076 2967 4084 2994
rect 4147 2976 4184 2984
rect 3767 2956 3984 2964
rect 4007 2956 4053 2964
rect 4076 2956 4093 2967
rect 4080 2953 4093 2956
rect 4176 2964 4184 2976
rect 4176 2956 4213 2964
rect 4236 2964 4244 2994
rect 4396 2967 4404 2994
rect 4236 2956 4273 2964
rect 4396 2956 4413 2967
rect 4400 2953 4413 2956
rect 1107 2936 1144 2944
rect 1567 2936 1633 2944
rect 1727 2936 1813 2944
rect 1967 2936 2033 2944
rect 2207 2936 2224 2947
rect 2207 2933 2220 2936
rect 2367 2936 2393 2944
rect 2407 2936 2453 2944
rect 2627 2936 2644 2947
rect 2627 2933 2640 2936
rect 3167 2936 3233 2944
rect 3587 2936 4153 2944
rect 4436 2944 4444 2993
rect 4456 2964 4464 3016
rect 4907 3016 5113 3024
rect 5207 3016 5273 3024
rect 5900 3024 5913 3027
rect 5896 3013 5913 3024
rect 6107 3016 6133 3024
rect 4576 2967 4584 2996
rect 4887 2996 4953 3004
rect 4967 2996 4992 3004
rect 5027 2996 5124 3004
rect 4656 2967 4664 2993
rect 4567 2956 4584 2967
rect 4567 2953 4580 2956
rect 4796 2964 4804 2993
rect 5116 2984 5124 2996
rect 5147 2997 5313 3005
rect 5487 2996 5533 3004
rect 5627 2996 5693 3004
rect 5373 2984 5387 2993
rect 5116 2976 5364 2984
rect 5373 2980 5424 2984
rect 5376 2976 5427 2980
rect 5356 2966 5364 2976
rect 5413 2967 5427 2976
rect 5776 2967 5784 2993
rect 5836 2967 5844 2993
rect 4707 2956 4804 2964
rect 4907 2955 5233 2963
rect 5567 2960 5604 2964
rect 5567 2956 5607 2960
rect 5593 2947 5607 2956
rect 5647 2956 5713 2964
rect 5896 2947 5904 3013
rect 5956 2967 5964 2993
rect 6016 2967 6024 2993
rect 6087 2955 6133 2963
rect 4267 2936 4444 2944
rect 5047 2936 5133 2944
rect 6007 2936 6093 2944
rect 627 2916 673 2924
rect 1087 2916 1293 2924
rect 1407 2916 1473 2924
rect 1636 2924 1644 2933
rect 1636 2916 1733 2924
rect 2187 2916 2233 2924
rect 2447 2916 2473 2924
rect 2727 2916 2793 2924
rect 3027 2916 3073 2924
rect 3087 2916 3113 2924
rect 4307 2916 4333 2924
rect 4387 2916 4553 2924
rect 5087 2916 5113 2924
rect 5867 2916 5933 2924
rect 6156 2924 6164 3053
rect 6127 2916 6164 2924
rect 147 2896 273 2904
rect 287 2896 573 2904
rect 1687 2896 1833 2904
rect 2427 2896 2493 2904
rect 2807 2896 2853 2904
rect 3187 2896 3293 2904
rect 3307 2896 3733 2904
rect 4007 2896 4113 2904
rect 4547 2896 4893 2904
rect 5167 2896 5413 2904
rect 5767 2896 6033 2904
rect 407 2876 813 2884
rect 907 2876 1133 2884
rect 1147 2876 1153 2884
rect 1247 2876 1333 2884
rect 1567 2876 1633 2884
rect 1887 2876 2013 2884
rect 2167 2876 2233 2884
rect 2547 2876 2953 2884
rect 3787 2876 3813 2884
rect 4107 2876 4273 2884
rect 4347 2876 4433 2884
rect 5207 2876 5233 2884
rect 5247 2876 5353 2884
rect 5547 2876 5613 2884
rect 227 2856 253 2864
rect 267 2856 513 2864
rect 1876 2864 1884 2873
rect 1627 2856 1884 2864
rect 2067 2856 2173 2864
rect 2347 2856 2393 2864
rect 2667 2856 2873 2864
rect 3036 2856 3353 2864
rect 567 2836 733 2844
rect 1067 2836 1253 2844
rect 1667 2836 2093 2844
rect 2227 2836 2253 2844
rect 2276 2836 2313 2844
rect 187 2816 333 2824
rect 507 2816 973 2824
rect 1347 2816 1553 2824
rect 1607 2816 2053 2824
rect 2116 2816 2133 2824
rect 787 2796 853 2804
rect 1187 2796 1307 2804
rect 1293 2788 1307 2796
rect 1507 2800 1544 2804
rect 1507 2796 1547 2800
rect 67 2776 93 2784
rect 227 2784 240 2787
rect 227 2773 244 2784
rect 307 2776 424 2784
rect 236 2746 244 2773
rect 416 2746 424 2776
rect 447 2776 553 2784
rect 607 2776 624 2784
rect 167 2736 233 2744
rect 507 2735 573 2743
rect 616 2744 624 2776
rect 687 2776 733 2784
rect 967 2776 993 2784
rect 1007 2776 1093 2784
rect 836 2747 844 2773
rect 1036 2764 1044 2776
rect 1307 2776 1433 2784
rect 1533 2787 1547 2796
rect 2116 2804 2124 2816
rect 2276 2824 2284 2836
rect 3036 2844 3044 2856
rect 3407 2856 3453 2864
rect 3687 2856 3733 2864
rect 4187 2856 4253 2864
rect 4536 2856 4593 2864
rect 4536 2847 4544 2856
rect 4687 2856 4753 2864
rect 4847 2856 5133 2864
rect 5327 2856 5393 2864
rect 5887 2856 5913 2864
rect 5967 2856 6133 2864
rect 2747 2836 3044 2844
rect 3187 2836 4033 2844
rect 4236 2836 4533 2844
rect 2147 2816 2284 2824
rect 2307 2816 2504 2824
rect 1807 2796 2124 2804
rect 2187 2796 2273 2804
rect 2496 2804 2504 2816
rect 2527 2816 2553 2824
rect 2907 2816 2973 2824
rect 3767 2816 3933 2824
rect 4236 2824 4244 2836
rect 4747 2836 4773 2844
rect 4796 2836 5173 2844
rect 4176 2816 4244 2824
rect 2496 2796 2733 2804
rect 3327 2796 3413 2804
rect 4176 2804 4184 2816
rect 4267 2816 4313 2824
rect 4527 2816 4553 2824
rect 4667 2816 4713 2824
rect 4796 2824 4804 2836
rect 5487 2836 5553 2844
rect 5627 2836 5713 2844
rect 4736 2816 4804 2824
rect 4736 2804 4744 2816
rect 4827 2816 4913 2824
rect 5016 2816 5173 2824
rect 5016 2804 5024 2816
rect 5267 2816 5433 2824
rect 5807 2816 5833 2824
rect 6027 2816 6053 2824
rect 4127 2796 4184 2804
rect 4656 2796 4744 2804
rect 4936 2796 5024 2804
rect 1787 2777 1833 2785
rect 2107 2777 2133 2785
rect 2427 2776 2604 2784
rect 1036 2756 1064 2764
rect 616 2736 753 2744
rect 976 2740 1013 2744
rect 973 2736 1013 2740
rect 973 2727 987 2736
rect 1056 2744 1064 2756
rect 1576 2747 1584 2773
rect 1656 2756 1804 2764
rect 1056 2736 1113 2744
rect 1507 2735 1533 2743
rect 1656 2744 1664 2756
rect 1627 2736 1664 2744
rect 1796 2746 1804 2756
rect 1973 2764 1987 2773
rect 2353 2764 2367 2773
rect 1867 2760 1987 2764
rect 2316 2760 2367 2764
rect 2596 2764 2604 2776
rect 2627 2776 2693 2784
rect 2716 2776 2833 2784
rect 1867 2756 1984 2760
rect 2316 2756 2364 2760
rect 2596 2756 2624 2764
rect 1707 2736 1753 2744
rect 2007 2740 2024 2744
rect 2007 2736 2027 2740
rect 127 2716 313 2724
rect 327 2716 353 2724
rect 1687 2716 1732 2724
rect 1753 2724 1767 2732
rect 2013 2727 2027 2736
rect 2316 2744 2324 2756
rect 2127 2736 2324 2744
rect 2347 2736 2433 2744
rect 2616 2744 2624 2756
rect 2716 2764 2724 2776
rect 2927 2776 3013 2784
rect 3367 2776 3393 2784
rect 2647 2756 2724 2764
rect 3356 2747 3364 2774
rect 3507 2776 3613 2784
rect 3667 2776 3713 2784
rect 3827 2777 3873 2785
rect 2616 2736 2673 2744
rect 1753 2716 1873 2724
rect 2167 2716 2413 2724
rect 2616 2724 2624 2736
rect 2727 2735 2773 2743
rect 2867 2736 2893 2744
rect 3007 2735 3233 2743
rect 3347 2736 3364 2747
rect 3347 2733 3360 2736
rect 3436 2744 3444 2773
rect 3407 2736 3513 2744
rect 3527 2735 3693 2743
rect 3776 2744 3784 2773
rect 3976 2747 3984 2793
rect 4167 2776 4193 2784
rect 4247 2776 4264 2784
rect 3776 2736 3793 2744
rect 3847 2735 3873 2743
rect 3887 2735 3913 2743
rect 3976 2736 3993 2747
rect 3980 2733 3993 2736
rect 4096 2744 4104 2773
rect 4087 2736 4104 2744
rect 4256 2747 4264 2776
rect 4287 2776 4384 2784
rect 4256 2736 4273 2747
rect 4260 2733 4273 2736
rect 4376 2746 4384 2776
rect 4467 2776 4513 2784
rect 4536 2776 4633 2784
rect 4536 2746 4544 2776
rect 4656 2784 4664 2796
rect 4647 2776 4664 2784
rect 4756 2776 4773 2784
rect 4696 2747 4704 2773
rect 4756 2747 4764 2776
rect 4836 2747 4844 2773
rect 4447 2736 4533 2744
rect 4587 2736 4653 2744
rect 4936 2744 4944 2796
rect 5076 2800 5153 2804
rect 5033 2784 5047 2793
rect 5073 2796 5153 2800
rect 5073 2787 5087 2796
rect 5467 2796 5553 2804
rect 5567 2796 5613 2804
rect 5967 2796 5993 2804
rect 5033 2780 5064 2784
rect 5036 2776 5064 2780
rect 5056 2747 5064 2776
rect 5096 2776 5253 2784
rect 4927 2736 4944 2744
rect 2527 2716 2624 2724
rect 3327 2716 3473 2724
rect 4827 2716 4853 2724
rect 4867 2716 4953 2724
rect 5096 2726 5104 2776
rect 5307 2776 5353 2784
rect 5416 2776 5473 2784
rect 5416 2747 5424 2776
rect 5773 2784 5787 2793
rect 5773 2780 5853 2784
rect 5776 2776 5853 2780
rect 5776 2764 5784 2776
rect 5636 2760 5784 2764
rect 5633 2756 5784 2760
rect 5633 2747 5647 2756
rect 5167 2736 5313 2744
rect 5507 2735 5553 2743
rect 5827 2736 5873 2744
rect 5896 2744 5904 2773
rect 5896 2736 6013 2744
rect 5316 2724 5324 2732
rect 5493 2724 5507 2732
rect 5316 2716 5507 2724
rect 5607 2716 5693 2724
rect 527 2696 913 2704
rect 1467 2696 1653 2704
rect 1847 2696 1893 2704
rect 2267 2696 2433 2704
rect 2547 2696 2753 2704
rect 2827 2696 2913 2704
rect 2927 2696 2953 2704
rect 3867 2696 3933 2704
rect 4047 2696 4213 2704
rect 4427 2696 4573 2704
rect 4596 2696 4793 2704
rect 27 2676 153 2684
rect 307 2676 333 2684
rect 1007 2676 1073 2684
rect 1087 2676 1153 2684
rect 1167 2676 1413 2684
rect 2027 2676 2453 2684
rect 2467 2676 2493 2684
rect 2567 2676 2633 2684
rect 2987 2676 3273 2684
rect 3627 2676 3753 2684
rect 4596 2684 4604 2696
rect 5207 2696 5353 2704
rect 4267 2676 4604 2684
rect 4696 2676 4813 2684
rect 687 2656 1784 2664
rect 227 2636 1633 2644
rect 1776 2644 1784 2656
rect 1867 2656 1893 2664
rect 2167 2656 2573 2664
rect 2596 2660 2693 2664
rect 2593 2656 2693 2660
rect 2593 2647 2607 2656
rect 2807 2656 2893 2664
rect 2967 2656 3093 2664
rect 3867 2656 3993 2664
rect 4696 2664 4704 2676
rect 4927 2676 4953 2684
rect 4007 2656 4704 2664
rect 5607 2656 5653 2664
rect 5667 2656 6013 2664
rect 6027 2656 6073 2664
rect 1776 2636 2273 2644
rect 2287 2636 2373 2644
rect 2727 2636 3313 2644
rect 3387 2636 3633 2644
rect 3707 2636 4433 2644
rect 4727 2636 4953 2644
rect 5467 2636 5813 2644
rect 667 2616 733 2624
rect 827 2616 1273 2624
rect 2047 2616 2213 2624
rect 2567 2616 2693 2624
rect 4187 2616 4453 2624
rect 4647 2616 5133 2624
rect 5147 2616 5233 2624
rect 5927 2616 6013 2624
rect 67 2596 513 2604
rect 887 2596 1313 2604
rect 1707 2596 1813 2604
rect 1867 2596 1913 2604
rect 2087 2596 2313 2604
rect 2427 2596 2853 2604
rect 3127 2596 3293 2604
rect 3387 2596 3573 2604
rect 3767 2596 4613 2604
rect 4947 2596 5073 2604
rect 5887 2596 6133 2604
rect 27 2576 713 2584
rect 1407 2576 1553 2584
rect 1667 2576 1793 2584
rect 2147 2576 2413 2584
rect 2707 2576 2793 2584
rect 2947 2576 3053 2584
rect 3227 2576 3313 2584
rect 4087 2576 4333 2584
rect 4347 2576 4393 2584
rect 4547 2576 4693 2584
rect 5767 2576 5913 2584
rect 6007 2576 6053 2584
rect 287 2556 473 2564
rect 487 2556 633 2564
rect 727 2556 833 2564
rect 987 2556 1373 2564
rect 1387 2556 1573 2564
rect 1827 2556 2233 2564
rect 2447 2556 2673 2564
rect 2867 2556 3333 2564
rect 3787 2556 3953 2564
rect 3967 2556 4393 2564
rect 4407 2556 4493 2564
rect 4507 2556 4753 2564
rect 4767 2556 4993 2564
rect 5227 2556 5333 2564
rect 5387 2556 5533 2564
rect 5776 2556 5833 2564
rect 5776 2547 5784 2556
rect 267 2536 893 2544
rect 1047 2536 1113 2544
rect 1187 2536 1424 2544
rect 1416 2527 1424 2536
rect 1607 2536 1753 2544
rect 1847 2536 2133 2544
rect 2307 2536 2513 2544
rect 3287 2536 3353 2544
rect 3427 2536 3753 2544
rect 4027 2536 4093 2544
rect 4327 2536 4453 2544
rect 4627 2536 4973 2544
rect 5267 2536 5433 2544
rect 5636 2536 5773 2544
rect 47 2516 213 2524
rect 407 2516 753 2524
rect 767 2516 813 2524
rect 947 2516 1133 2524
rect 1427 2516 1813 2524
rect 2527 2516 2713 2524
rect 2847 2516 3073 2524
rect 4507 2516 4633 2524
rect 5636 2524 5644 2536
rect 6067 2536 6133 2544
rect 5187 2516 5644 2524
rect 1207 2496 1253 2504
rect 1507 2496 1713 2504
rect 1787 2496 1953 2504
rect 2036 2496 2093 2504
rect 87 2476 124 2484
rect 116 2447 124 2476
rect 147 2476 253 2484
rect 367 2476 453 2484
rect 467 2476 513 2484
rect 1027 2477 1053 2485
rect 636 2464 644 2474
rect 587 2456 644 2464
rect 676 2447 684 2474
rect 1247 2477 1313 2485
rect 1627 2477 1693 2485
rect 1827 2476 1892 2484
rect 676 2436 693 2447
rect 680 2433 693 2436
rect 1047 2436 1333 2444
rect 1387 2436 1693 2444
rect 1756 2446 1764 2473
rect 1816 2464 1824 2474
rect 1816 2456 1884 2464
rect 1767 2435 1833 2443
rect 67 2416 172 2424
rect 207 2416 413 2424
rect 687 2416 713 2424
rect 1027 2416 1053 2424
rect 1527 2416 1633 2424
rect 1727 2416 1793 2424
rect 1876 2424 1884 2456
rect 1916 2447 1924 2474
rect 2036 2464 2044 2496
rect 2147 2496 2193 2504
rect 2207 2496 2353 2504
rect 2536 2496 2633 2504
rect 2267 2484 2280 2487
rect 2267 2473 2284 2484
rect 2447 2476 2473 2484
rect 2153 2464 2167 2473
rect 2007 2456 2044 2464
rect 2096 2460 2167 2464
rect 2096 2456 2164 2460
rect 1907 2436 1924 2447
rect 1907 2433 1920 2436
rect 1987 2436 2013 2444
rect 2096 2446 2104 2456
rect 2216 2444 2224 2473
rect 2216 2436 2253 2444
rect 1876 2416 1913 2424
rect 2276 2424 2284 2473
rect 2336 2447 2344 2473
rect 2536 2446 2544 2496
rect 2767 2496 3033 2504
rect 3156 2496 3293 2504
rect 2627 2477 2673 2485
rect 2907 2476 2973 2484
rect 2713 2464 2727 2473
rect 2713 2460 2933 2464
rect 2716 2456 2933 2460
rect 3016 2447 3024 2474
rect 2407 2435 2433 2443
rect 2767 2434 2792 2442
rect 2827 2440 2924 2444
rect 2827 2436 2927 2440
rect 2227 2416 2284 2424
rect 2913 2427 2927 2436
rect 3007 2436 3024 2447
rect 3007 2433 3020 2436
rect 3156 2444 3164 2496
rect 3507 2496 3553 2504
rect 4047 2496 4113 2504
rect 4127 2496 4153 2504
rect 4567 2496 4593 2504
rect 4756 2496 4833 2504
rect 3187 2476 3284 2484
rect 3276 2446 3284 2476
rect 3347 2477 3393 2485
rect 3467 2476 3484 2484
rect 3476 2447 3484 2476
rect 3576 2464 3584 2474
rect 3747 2476 3833 2484
rect 3856 2476 3893 2484
rect 3856 2464 3864 2476
rect 4227 2477 4273 2485
rect 4336 2476 4393 2484
rect 3527 2456 3584 2464
rect 3796 2456 3864 2464
rect 3087 2436 3164 2444
rect 3796 2446 3804 2456
rect 4076 2446 4084 2473
rect 3687 2436 3753 2444
rect 4027 2435 4073 2443
rect 4336 2446 4344 2476
rect 4467 2476 4524 2484
rect 4516 2467 4524 2476
rect 4756 2484 4764 2496
rect 4847 2496 4873 2504
rect 5507 2496 5553 2504
rect 5647 2496 5693 2504
rect 5707 2496 5733 2504
rect 5807 2504 5820 2507
rect 5807 2493 5824 2504
rect 5867 2496 5933 2504
rect 4676 2476 4764 2484
rect 4516 2456 4533 2467
rect 4520 2453 4533 2456
rect 4127 2436 4284 2444
rect 3047 2416 3073 2424
rect 767 2396 853 2404
rect 907 2396 1093 2404
rect 1147 2396 1373 2404
rect 1676 2396 1733 2404
rect 1676 2387 1684 2396
rect 1887 2396 1933 2404
rect 2216 2404 2224 2413
rect 3327 2416 3513 2424
rect 4067 2416 4153 2424
rect 4276 2424 4284 2436
rect 4387 2435 4413 2443
rect 4596 2444 4604 2473
rect 4487 2436 4604 2444
rect 4676 2444 4684 2476
rect 4787 2476 4824 2484
rect 4816 2467 4824 2476
rect 4816 2456 4833 2467
rect 4820 2453 4833 2456
rect 4996 2447 5004 2473
rect 4667 2436 4684 2444
rect 4707 2435 4793 2443
rect 5056 2446 5064 2493
rect 5076 2447 5084 2474
rect 5147 2484 5160 2487
rect 5147 2473 5164 2484
rect 5076 2436 5093 2447
rect 5080 2433 5093 2436
rect 5156 2446 5164 2473
rect 5276 2476 5293 2484
rect 5276 2447 5284 2476
rect 5336 2427 5344 2474
rect 5427 2476 5464 2484
rect 5373 2464 5387 2473
rect 5356 2460 5387 2464
rect 5356 2456 5384 2460
rect 5356 2446 5364 2456
rect 5456 2446 5464 2476
rect 5513 2464 5527 2473
rect 5476 2460 5527 2464
rect 5473 2456 5524 2460
rect 5473 2447 5487 2456
rect 5547 2436 5613 2444
rect 5716 2444 5724 2473
rect 5816 2464 5824 2493
rect 5816 2460 5884 2464
rect 5816 2456 5887 2460
rect 5873 2447 5887 2456
rect 5996 2447 6004 2473
rect 6076 2447 6084 2473
rect 5687 2436 5724 2444
rect 5807 2435 5833 2443
rect 5947 2436 5973 2444
rect 4276 2416 4353 2424
rect 4727 2416 4753 2424
rect 5267 2416 5312 2424
rect 5567 2416 5593 2424
rect 5707 2416 5733 2424
rect 2067 2396 2224 2404
rect 2347 2396 2713 2404
rect 2987 2396 3553 2404
rect 3927 2396 4953 2404
rect 4967 2396 5073 2404
rect 5667 2396 5713 2404
rect 5727 2396 5833 2404
rect 5907 2396 6013 2404
rect 6067 2396 6093 2404
rect 47 2376 93 2384
rect 267 2376 293 2384
rect 487 2376 533 2384
rect 547 2376 613 2384
rect 627 2376 713 2384
rect 727 2376 1113 2384
rect 1167 2376 1233 2384
rect 1607 2376 1673 2384
rect 1747 2376 1853 2384
rect 1967 2376 2313 2384
rect 2507 2376 2853 2384
rect 2867 2376 3133 2384
rect 3967 2376 4013 2384
rect 4367 2376 4653 2384
rect 4927 2376 5113 2384
rect 5267 2376 6033 2384
rect 747 2356 793 2364
rect 807 2356 1072 2364
rect 1107 2356 1473 2364
rect 1567 2356 1973 2364
rect 2027 2356 2092 2364
rect 2127 2356 2493 2364
rect 2507 2356 2593 2364
rect 2667 2356 2833 2364
rect 2987 2356 3113 2364
rect 4207 2356 4333 2364
rect 4987 2356 5293 2364
rect 5507 2356 5973 2364
rect 6107 2356 6133 2364
rect 87 2336 113 2344
rect 207 2336 293 2344
rect 307 2336 353 2344
rect 407 2336 573 2344
rect 587 2336 913 2344
rect 927 2336 953 2344
rect 1347 2336 1393 2344
rect 1467 2336 1653 2344
rect 1707 2336 1824 2344
rect 1816 2327 1824 2336
rect 1887 2336 1913 2344
rect 1927 2336 2353 2344
rect 2687 2336 3613 2344
rect 3667 2336 3733 2344
rect 4067 2336 4273 2344
rect 4487 2336 4533 2344
rect 4727 2336 4813 2344
rect 5007 2336 5053 2344
rect 5127 2336 5253 2344
rect 5367 2336 5473 2344
rect 5607 2336 5653 2344
rect 967 2316 1033 2324
rect 1187 2316 1273 2324
rect 1287 2316 1413 2324
rect 1427 2316 1693 2324
rect 1827 2316 2113 2324
rect 2487 2316 2593 2324
rect 2847 2316 2993 2324
rect 3007 2316 3033 2324
rect 3056 2316 3373 2324
rect 127 2296 253 2304
rect 387 2296 464 2304
rect 456 2287 464 2296
rect 847 2296 1153 2304
rect 1207 2296 1444 2304
rect 1436 2287 1444 2296
rect 1667 2296 1753 2304
rect 1807 2296 2013 2304
rect 2207 2296 2412 2304
rect 2447 2296 2713 2304
rect 3056 2304 3064 2316
rect 3387 2316 3513 2324
rect 3833 2324 3847 2333
rect 3833 2320 4113 2324
rect 3836 2316 4113 2320
rect 4167 2316 4193 2324
rect 4207 2316 4293 2324
rect 4827 2316 5093 2324
rect 5107 2316 5153 2324
rect 5167 2316 5273 2324
rect 5287 2316 5573 2324
rect 5867 2316 5913 2324
rect 5967 2316 6013 2324
rect 6067 2316 6113 2324
rect 2827 2296 3064 2304
rect 3547 2296 3873 2304
rect 327 2276 353 2284
rect 467 2276 513 2284
rect 687 2276 753 2284
rect -24 2256 33 2264
rect 167 2257 233 2265
rect -24 2204 -16 2224
rect 107 2215 233 2223
rect 276 2207 284 2273
rect 847 2276 873 2284
rect 1447 2276 1493 2284
rect 1507 2276 1633 2284
rect 1947 2276 2013 2284
rect 407 2264 420 2267
rect 407 2253 424 2264
rect 447 2256 464 2264
rect 416 2226 424 2253
rect 327 2215 373 2223
rect 456 2207 464 2256
rect 627 2256 653 2264
rect 707 2256 1013 2264
rect 1067 2256 1173 2264
rect 1227 2256 1333 2264
rect 1347 2256 1504 2264
rect 696 2227 704 2253
rect 527 2215 553 2223
rect 787 2216 893 2224
rect 947 2216 973 2224
rect 1247 2215 1273 2223
rect 1327 2216 1473 2224
rect 1496 2224 1504 2256
rect 1727 2257 1773 2265
rect 1855 2227 1863 2273
rect 2307 2276 2373 2284
rect 3427 2276 3493 2284
rect 3567 2276 3593 2284
rect 3947 2276 4064 2284
rect 2107 2256 2152 2264
rect 1893 2244 1907 2253
rect 1876 2240 1907 2244
rect 1876 2236 1904 2240
rect 1876 2227 1884 2236
rect 1956 2227 1964 2253
rect 2253 2264 2267 2273
rect 2187 2260 2267 2264
rect 2187 2256 2264 2260
rect 2907 2257 2933 2265
rect 3007 2257 3073 2265
rect 3187 2256 3273 2264
rect 3367 2257 3393 2265
rect 3627 2256 3653 2264
rect 3840 2264 3853 2267
rect 1996 2240 2433 2244
rect 1993 2236 2433 2240
rect 1993 2227 2007 2236
rect 3473 2244 3487 2253
rect 3836 2253 3853 2264
rect 3987 2257 4033 2265
rect 3473 2240 3524 2244
rect 3476 2236 3527 2240
rect 1496 2216 1512 2224
rect 1547 2216 1653 2224
rect 1887 2216 1913 2224
rect 2087 2220 2203 2224
rect 2216 2220 2633 2224
rect 2087 2216 2207 2220
rect 2193 2207 2207 2216
rect -24 2196 73 2204
rect 276 2196 293 2207
rect 280 2193 293 2196
rect 447 2196 464 2207
rect 447 2193 460 2196
rect 1387 2196 1433 2204
rect 1767 2196 1793 2204
rect 2206 2200 2207 2207
rect 2213 2216 2633 2220
rect 2213 2207 2227 2216
rect 2713 2224 2727 2233
rect 3513 2227 3527 2236
rect 2713 2220 2753 2224
rect 2716 2216 2753 2220
rect 2927 2216 2993 2224
rect 3836 2224 3844 2253
rect 4056 2244 4064 2276
rect 4107 2276 4213 2284
rect 4253 2276 4873 2284
rect 4253 2268 4267 2276
rect 4987 2276 5013 2284
rect 5087 2276 5213 2284
rect 6007 2276 6053 2284
rect 4256 2244 4264 2254
rect 4367 2256 4424 2264
rect 4313 2244 4327 2253
rect 3887 2236 4004 2244
rect 4056 2236 4264 2244
rect 4276 2240 4327 2244
rect 4416 2244 4424 2256
rect 4447 2257 4573 2265
rect 4620 2264 4633 2267
rect 4616 2253 4633 2264
rect 4787 2257 4833 2265
rect 5447 2256 5513 2264
rect 5527 2257 5553 2265
rect 4416 2240 4484 2244
rect 4276 2236 4324 2240
rect 4416 2236 4487 2240
rect 3996 2226 4004 2236
rect 3907 2216 3953 2224
rect 4236 2224 4244 2236
rect 4276 2226 4284 2236
rect 4473 2227 4487 2236
rect 4147 2216 4244 2224
rect 4616 2224 4624 2253
rect 5036 2236 5093 2244
rect 5036 2226 5044 2236
rect 5336 2227 5344 2253
rect 5216 2216 5304 2224
rect 2367 2196 2553 2204
rect 2747 2196 2773 2204
rect 3067 2196 3153 2204
rect 3287 2196 3533 2204
rect 3587 2196 4093 2204
rect 5216 2204 5224 2216
rect 5147 2196 5224 2204
rect 5296 2204 5304 2216
rect 5576 2226 5584 2273
rect 5607 2256 5624 2264
rect 5356 2216 5453 2224
rect 5356 2204 5364 2216
rect 5616 2207 5624 2256
rect 5787 2256 5824 2264
rect 5816 2227 5824 2256
rect 5916 2227 5924 2253
rect 6016 2227 6024 2253
rect 5296 2196 5364 2204
rect 5607 2196 5624 2207
rect 5607 2193 5620 2196
rect 247 2176 333 2184
rect 607 2176 693 2184
rect 747 2176 853 2184
rect 1087 2176 1153 2184
rect 1167 2176 1313 2184
rect 1667 2176 1713 2184
rect 1907 2176 2273 2184
rect 2347 2176 2633 2184
rect 3187 2176 3233 2184
rect 3607 2176 3913 2184
rect 3967 2176 4013 2184
rect 4867 2176 5033 2184
rect 5287 2176 5373 2184
rect 5527 2176 5733 2184
rect 736 2164 744 2173
rect 467 2156 744 2164
rect 1127 2156 1193 2164
rect 1287 2156 1393 2164
rect 1607 2156 1733 2164
rect 2047 2156 2233 2164
rect 2307 2156 2353 2164
rect 2427 2156 2613 2164
rect 2987 2156 3253 2164
rect 3727 2156 3873 2164
rect 3947 2156 4373 2164
rect 4607 2156 4793 2164
rect 5447 2156 5653 2164
rect 227 2136 773 2144
rect 1416 2136 1533 2144
rect 147 2116 193 2124
rect 287 2116 593 2124
rect 1416 2124 1424 2136
rect 1627 2136 1673 2144
rect 1987 2136 2324 2144
rect 1327 2116 1424 2124
rect 1436 2116 1613 2124
rect 1436 2104 1444 2116
rect 1907 2116 2213 2124
rect 2316 2124 2324 2136
rect 2447 2136 2953 2144
rect 3787 2136 3853 2144
rect 4627 2136 4833 2144
rect 2316 2116 2413 2124
rect 2427 2116 2473 2124
rect 2527 2116 3313 2124
rect 3927 2116 4073 2124
rect 4467 2116 4493 2124
rect 5427 2116 5773 2124
rect 47 2096 1444 2104
rect 1636 2096 1704 2104
rect 87 2076 1393 2084
rect 1636 2084 1644 2096
rect 1607 2076 1644 2084
rect 1696 2084 1704 2096
rect 1727 2096 1833 2104
rect 1847 2096 1992 2104
rect 2027 2096 2373 2104
rect 2567 2096 2673 2104
rect 3227 2096 3573 2104
rect 4347 2096 4613 2104
rect 4727 2096 4933 2104
rect 5127 2096 5373 2104
rect 5587 2096 5853 2104
rect 1696 2076 1973 2084
rect 2047 2076 2092 2084
rect 2127 2076 2153 2084
rect 2547 2076 2753 2084
rect 2767 2076 3453 2084
rect 3607 2076 3993 2084
rect 4007 2076 4213 2084
rect 4427 2076 4593 2084
rect 5267 2076 5353 2084
rect 307 2056 593 2064
rect 1047 2056 1413 2064
rect 1547 2056 1573 2064
rect 1667 2056 2233 2064
rect 2467 2056 2513 2064
rect 3407 2056 4753 2064
rect 5087 2056 5293 2064
rect 5407 2056 5573 2064
rect 5687 2056 5933 2064
rect 907 2036 1353 2044
rect 1467 2036 1592 2044
rect 1627 2036 2033 2044
rect 2107 2036 2153 2044
rect 2227 2036 2433 2044
rect 3567 2036 3653 2044
rect 4536 2036 4713 2044
rect 107 2016 293 2024
rect 547 2016 613 2024
rect 707 2016 773 2024
rect 2087 2016 2333 2024
rect 807 1996 913 2004
rect 1007 1996 1164 2004
rect 1156 1987 1164 1996
rect 1487 1996 1713 2004
rect 2153 2006 2167 2016
rect 2467 2016 2713 2024
rect 2727 2016 3213 2024
rect 3227 2016 3384 2024
rect 3376 2007 3384 2016
rect 4536 2024 4544 2036
rect 4167 2016 4384 2024
rect 2247 1996 2284 2004
rect 407 1976 493 1984
rect 507 1976 773 1984
rect 1167 1976 1313 1984
rect 2087 1976 2113 1984
rect 2276 1984 2284 1996
rect 2307 1996 2393 2004
rect 2547 1996 3352 2004
rect 3387 1996 3513 2004
rect 4267 1996 4313 2004
rect 4376 2004 4384 2016
rect 4516 2016 4544 2024
rect 4376 1996 4473 2004
rect 2433 1984 2447 1993
rect 2276 1980 2447 1984
rect 2276 1976 2444 1980
rect 2607 1976 2853 1984
rect 3567 1976 3633 1984
rect 3676 1976 3913 1984
rect 116 1907 124 1954
rect 307 1956 324 1964
rect 176 1927 184 1953
rect 256 1924 264 1954
rect 316 1927 324 1956
rect 447 1956 533 1964
rect 646 1953 647 1960
rect 667 1956 753 1964
rect 356 1927 364 1953
rect 633 1944 647 1953
rect 816 1944 824 1954
rect 633 1940 664 1944
rect 796 1940 824 1944
rect 636 1936 664 1940
rect 656 1927 664 1936
rect 227 1916 264 1924
rect 427 1916 513 1924
rect 527 1915 593 1923
rect 647 1924 664 1927
rect 793 1936 824 1940
rect 793 1927 807 1936
rect 647 1916 673 1924
rect 647 1913 660 1916
rect 856 1907 864 1954
rect 967 1957 1033 1965
rect 1247 1957 1273 1965
rect 1340 1964 1353 1967
rect 893 1944 907 1953
rect 876 1940 907 1944
rect 876 1936 904 1940
rect 876 1926 884 1936
rect 927 1916 973 1924
rect 1116 1924 1124 1954
rect 1336 1953 1353 1964
rect 1507 1956 1533 1964
rect 1627 1957 1693 1965
rect 1867 1956 1924 1964
rect 1336 1926 1344 1953
rect 1393 1944 1407 1953
rect 1393 1940 1893 1944
rect 1396 1936 1893 1940
rect 1916 1944 1924 1956
rect 1947 1956 2093 1964
rect 2147 1957 2233 1965
rect 2247 1956 2472 1964
rect 2527 1957 2573 1965
rect 2927 1957 2953 1965
rect 3027 1957 3073 1965
rect 3267 1957 3293 1965
rect 3367 1957 3413 1965
rect 3676 1964 3684 1976
rect 4173 1984 4187 1993
rect 4516 1987 4524 2016
rect 4567 2016 4613 2024
rect 4887 2016 5453 2024
rect 5787 2016 5953 2024
rect 5967 2016 6033 2024
rect 5187 1996 5393 2004
rect 5647 1996 5673 2004
rect 4107 1980 4187 1984
rect 4107 1976 4184 1980
rect 4261 1976 4333 1984
rect 4516 1976 4533 1987
rect 4520 1973 4533 1976
rect 4647 1976 4733 1984
rect 4907 1976 4973 1984
rect 5027 1976 5093 1984
rect 5547 1976 5593 1984
rect 5807 1976 5853 1984
rect 3427 1956 3684 1964
rect 3707 1956 3793 1964
rect 3847 1957 3893 1965
rect 1916 1936 2313 1944
rect 2676 1927 2684 1954
rect 3956 1944 3964 1954
rect 2767 1936 2984 1944
rect 1027 1916 1124 1924
rect 1187 1916 1333 1924
rect 1647 1916 1953 1924
rect 2447 1915 2493 1923
rect 2667 1916 2684 1927
rect 2976 1926 2984 1936
rect 3616 1936 3964 1944
rect 2667 1913 2680 1916
rect 3167 1916 3193 1924
rect 3207 1915 3233 1923
rect 3616 1924 3624 1936
rect 3547 1916 3624 1924
rect 3647 1915 3713 1923
rect 4047 1916 4093 1924
rect 4216 1924 4224 1953
rect 4276 1944 4284 1954
rect 4276 1936 4304 1944
rect 4296 1927 4304 1936
rect 4347 1944 4360 1947
rect 4347 1940 4364 1944
rect 4347 1933 4367 1940
rect 4353 1927 4367 1933
rect 4216 1916 4253 1924
rect 4296 1916 4313 1927
rect 4300 1913 4313 1916
rect 207 1896 373 1904
rect 1767 1896 2053 1904
rect 2247 1896 2393 1904
rect 2887 1896 2913 1904
rect 2927 1896 2972 1904
rect 3007 1896 3293 1904
rect 4347 1896 4373 1904
rect 4396 1904 4404 1954
rect 4436 1924 4444 1954
rect 4607 1956 4653 1964
rect 4807 1956 4884 1964
rect 4436 1916 4553 1924
rect 4696 1924 4704 1954
rect 4876 1944 4884 1956
rect 4936 1944 4944 1954
rect 5073 1944 5087 1953
rect 4876 1936 4944 1944
rect 4696 1916 4733 1924
rect 4827 1920 4844 1924
rect 4827 1916 4847 1920
rect 4833 1907 4847 1916
rect 4936 1907 4944 1936
rect 5036 1940 5087 1944
rect 5156 1956 5193 1964
rect 5036 1936 5084 1940
rect 5036 1924 5044 1936
rect 4967 1916 5044 1924
rect 5156 1924 5164 1956
rect 5127 1916 5164 1924
rect 5275 1924 5283 1953
rect 5227 1916 5283 1924
rect 5296 1907 5304 1954
rect 4396 1896 4433 1904
rect 5067 1896 5093 1904
rect 5287 1896 5304 1907
rect 5336 1904 5344 1954
rect 5507 1956 5553 1964
rect 5667 1957 5733 1965
rect 5887 1956 5913 1964
rect 5433 1944 5447 1953
rect 5433 1940 5593 1944
rect 5436 1936 5593 1940
rect 5367 1916 5412 1924
rect 5447 1915 5473 1923
rect 5527 1915 5573 1923
rect 5627 1916 5673 1924
rect 5767 1916 5933 1924
rect 5947 1915 6073 1923
rect 5336 1896 5453 1904
rect 5287 1893 5300 1896
rect 5807 1896 5873 1904
rect 396 1876 553 1884
rect 47 1856 93 1864
rect 147 1856 333 1864
rect 396 1864 404 1876
rect 787 1876 833 1884
rect 1087 1876 1133 1884
rect 1327 1876 1373 1884
rect 1547 1876 1693 1884
rect 1987 1876 2033 1884
rect 2556 1876 3113 1884
rect 2556 1867 2564 1876
rect 3167 1876 3533 1884
rect 3547 1876 3773 1884
rect 3907 1876 3973 1884
rect 3987 1876 4213 1884
rect 4227 1876 4293 1884
rect 4307 1876 4513 1884
rect 4567 1876 4633 1884
rect 5487 1876 5592 1884
rect 5627 1876 5713 1884
rect 5867 1876 5973 1884
rect 347 1856 404 1864
rect 1727 1856 1772 1864
rect 1807 1856 2093 1864
rect 2227 1856 2333 1864
rect 2467 1856 2553 1864
rect 2847 1856 3033 1864
rect 3307 1856 3573 1864
rect 3827 1856 3973 1864
rect 4067 1856 4273 1864
rect 4427 1856 4473 1864
rect 4627 1856 5173 1864
rect 5467 1856 5733 1864
rect 127 1836 273 1844
rect 287 1836 433 1844
rect 447 1836 713 1844
rect 2127 1836 2193 1844
rect 2207 1836 2373 1844
rect 2387 1836 2713 1844
rect 2927 1836 3013 1844
rect 3727 1836 4053 1844
rect 4787 1836 5073 1844
rect 5207 1836 5373 1844
rect 5647 1836 5693 1844
rect 5927 1836 5953 1844
rect 867 1816 1073 1824
rect 1087 1816 1253 1824
rect 1267 1816 1553 1824
rect 1607 1816 1653 1824
rect 1707 1816 1813 1824
rect 1947 1816 1993 1824
rect 2007 1816 2392 1824
rect 2427 1816 2753 1824
rect 3407 1816 4313 1824
rect 4327 1816 4473 1824
rect 4487 1816 4633 1824
rect 4887 1816 4973 1824
rect 5027 1816 5104 1824
rect 5096 1807 5104 1816
rect 5907 1816 5973 1824
rect 67 1796 233 1804
rect 727 1796 913 1804
rect 927 1796 953 1804
rect 1407 1796 1573 1804
rect 1587 1796 1673 1804
rect 2507 1796 2633 1804
rect 2707 1796 2793 1804
rect 2807 1796 3073 1804
rect 3087 1796 3333 1804
rect 3667 1796 3793 1804
rect 4007 1796 4073 1804
rect 5096 1796 5113 1807
rect 5100 1793 5113 1796
rect 5327 1796 5633 1804
rect 267 1776 404 1784
rect 396 1764 404 1776
rect 1167 1776 1213 1784
rect 1467 1776 1493 1784
rect 2127 1776 2173 1784
rect 2327 1776 2413 1784
rect 2727 1776 2853 1784
rect 2867 1776 2993 1784
rect 3127 1776 3253 1784
rect 3627 1776 3853 1784
rect 3867 1776 4133 1784
rect 4367 1776 4413 1784
rect 4707 1776 4973 1784
rect 5220 1784 5233 1787
rect 5216 1773 5233 1784
rect 5507 1776 5613 1784
rect 327 1756 384 1764
rect 396 1756 444 1764
rect 67 1736 113 1744
rect 167 1736 213 1744
rect 227 1736 293 1744
rect 376 1744 384 1756
rect 376 1736 424 1744
rect 147 1695 193 1703
rect 207 1696 273 1704
rect 296 1704 304 1734
rect 296 1696 373 1704
rect 416 1706 424 1736
rect 436 1687 444 1756
rect 507 1756 553 1764
rect 807 1756 873 1764
rect 887 1756 1333 1764
rect 1347 1756 1433 1764
rect 1627 1756 1693 1764
rect 1707 1756 1833 1764
rect 1967 1756 2013 1764
rect 2407 1756 2633 1764
rect 3107 1756 3164 1764
rect 576 1707 584 1734
rect 647 1744 660 1747
rect 647 1733 664 1744
rect 687 1737 753 1745
rect 827 1736 933 1744
rect 1196 1736 1293 1744
rect 467 1695 493 1703
rect 576 1696 593 1707
rect 580 1693 593 1696
rect 656 1706 664 1733
rect 747 1696 873 1704
rect 887 1695 973 1703
rect 996 1704 1004 1734
rect 1196 1707 1204 1736
rect 1456 1736 1493 1744
rect 1456 1727 1464 1736
rect 1560 1744 1573 1747
rect 1236 1716 1333 1724
rect 996 1696 1093 1704
rect 1236 1706 1244 1716
rect 1447 1716 1464 1727
rect 1556 1733 1573 1744
rect 1647 1736 1684 1744
rect 1756 1740 2013 1744
rect 1447 1713 1460 1716
rect 1556 1706 1564 1733
rect 1676 1706 1684 1736
rect 1753 1736 2013 1740
rect 1753 1726 1767 1736
rect 2107 1737 2133 1745
rect 2176 1736 2213 1744
rect 1947 1695 1993 1703
rect 2056 1704 2064 1734
rect 2176 1724 2184 1736
rect 2236 1736 2293 1744
rect 2236 1724 2244 1736
rect 2556 1724 2564 1734
rect 2667 1736 2693 1744
rect 2707 1736 2933 1744
rect 2156 1716 2184 1724
rect 2196 1716 2244 1724
rect 2496 1716 2564 1724
rect 2056 1696 2113 1704
rect 2156 1706 2164 1716
rect 2196 1706 2204 1716
rect 2496 1707 2504 1716
rect 2327 1695 2373 1703
rect 2487 1696 2504 1707
rect 2487 1693 2500 1696
rect 2547 1695 2612 1703
rect 2647 1696 2673 1704
rect 2747 1696 2813 1704
rect 2907 1695 3093 1703
rect 3156 1704 3164 1756
rect 4207 1756 4293 1764
rect 4607 1764 4620 1767
rect 4607 1753 4624 1764
rect 4667 1764 4680 1767
rect 4667 1753 4684 1764
rect 4727 1756 4753 1764
rect 4767 1756 4853 1764
rect 3267 1736 3393 1744
rect 3440 1744 3453 1747
rect 3436 1733 3453 1744
rect 3507 1737 3533 1745
rect 3547 1736 3573 1744
rect 3847 1737 3893 1745
rect 3436 1724 3444 1733
rect 3936 1724 3944 1734
rect 3416 1720 3444 1724
rect 3916 1720 3944 1724
rect 3413 1716 3444 1720
rect 3913 1716 3944 1720
rect 3413 1707 3427 1716
rect 3156 1696 3284 1704
rect 767 1676 793 1684
rect 1027 1676 1133 1684
rect 1727 1676 1813 1684
rect 1827 1676 2073 1684
rect 3276 1684 3284 1696
rect 3307 1696 3333 1704
rect 3347 1695 3373 1703
rect 3913 1707 3927 1716
rect 3976 1707 3984 1733
rect 3487 1695 3513 1703
rect 3607 1695 3853 1703
rect 4036 1687 4044 1734
rect 4056 1706 4064 1753
rect 4076 1736 4353 1744
rect 3276 1676 3333 1684
rect 1136 1664 1144 1673
rect 4076 1684 4084 1736
rect 4147 1695 4173 1703
rect 4516 1704 4524 1734
rect 4616 1707 4624 1753
rect 4676 1707 4684 1753
rect 4796 1736 4833 1744
rect 4516 1696 4592 1704
rect 4796 1706 4804 1736
rect 4953 1724 4967 1733
rect 4916 1720 4967 1724
rect 4916 1716 4964 1720
rect 4916 1704 4924 1716
rect 5056 1707 5064 1733
rect 5216 1707 5224 1773
rect 5327 1756 5393 1764
rect 5407 1756 5567 1764
rect 5553 1748 5567 1756
rect 5816 1764 5824 1813
rect 5727 1756 5824 1764
rect 5496 1736 5513 1744
rect 5253 1724 5267 1733
rect 5253 1720 5384 1724
rect 5256 1716 5387 1720
rect 5373 1707 5387 1716
rect 4847 1696 4924 1704
rect 4047 1676 4084 1684
rect 4107 1676 4233 1684
rect 4427 1676 4493 1684
rect 4947 1676 5033 1684
rect 5436 1684 5444 1733
rect 5496 1687 5504 1736
rect 5567 1737 5593 1745
rect 5856 1726 5864 1813
rect 5656 1704 5664 1714
rect 5876 1716 5953 1724
rect 5876 1704 5884 1716
rect 5616 1696 5664 1704
rect 5676 1700 5884 1704
rect 5673 1696 5884 1700
rect 5367 1676 5444 1684
rect 5487 1676 5504 1687
rect 5487 1673 5500 1676
rect 5616 1684 5624 1696
rect 5673 1687 5687 1696
rect 5587 1676 5624 1684
rect 5685 1680 5687 1687
rect 1136 1656 1273 1664
rect 1387 1656 1613 1664
rect 2287 1656 2493 1664
rect 2576 1656 2673 1664
rect 2576 1647 2584 1656
rect 2687 1656 3153 1664
rect 4167 1656 4353 1664
rect 4527 1656 4653 1664
rect 5167 1656 5293 1664
rect 387 1636 693 1644
rect 1527 1636 1753 1644
rect 1927 1636 2233 1644
rect 2307 1636 2573 1644
rect 2627 1636 2813 1644
rect 2947 1636 3553 1644
rect 4987 1636 5073 1644
rect 5547 1636 5693 1644
rect 1076 1616 1733 1624
rect 407 1596 593 1604
rect 607 1596 993 1604
rect 1076 1604 1084 1616
rect 2167 1616 2524 1624
rect 1047 1596 1084 1604
rect 1427 1596 1953 1604
rect 2107 1596 2313 1604
rect 2516 1604 2524 1616
rect 3087 1616 3233 1624
rect 3927 1616 4333 1624
rect 5287 1616 5473 1624
rect 2516 1596 2913 1604
rect 3267 1596 3653 1604
rect 3667 1596 3813 1604
rect 3827 1596 3853 1604
rect 3867 1596 4373 1604
rect 4387 1596 4553 1604
rect 5156 1596 5233 1604
rect 107 1576 413 1584
rect 1607 1576 1772 1584
rect 1807 1576 2084 1584
rect 167 1556 333 1564
rect 487 1556 833 1564
rect 1007 1556 1853 1564
rect 2076 1564 2084 1576
rect 4367 1576 4653 1584
rect 5156 1584 5164 1596
rect 5716 1587 5724 1673
rect 5976 1667 5984 1733
rect 6007 1716 6044 1724
rect 6036 1687 6044 1716
rect 4667 1576 5164 1584
rect 2076 1556 2293 1564
rect 2347 1556 2973 1564
rect 3427 1556 3613 1564
rect 4307 1556 4833 1564
rect 4847 1556 5173 1564
rect 1327 1536 1493 1544
rect 1616 1536 1913 1544
rect 1616 1527 1624 1536
rect 2336 1544 2344 1553
rect 2167 1536 2344 1544
rect 2427 1536 2873 1544
rect 5207 1536 5273 1544
rect 5327 1536 5433 1544
rect 127 1516 213 1524
rect 227 1516 433 1524
rect 1087 1516 1173 1524
rect 1567 1516 1612 1524
rect 1647 1516 1793 1524
rect 1867 1516 1933 1524
rect 1947 1516 2132 1524
rect 2416 1524 2424 1533
rect 2167 1516 2424 1524
rect 2447 1516 2864 1524
rect 267 1496 313 1504
rect 1527 1496 1593 1504
rect 2067 1496 2213 1504
rect 2227 1496 2253 1504
rect 2856 1504 2864 1516
rect 3287 1516 3433 1524
rect 3807 1516 4173 1524
rect 4767 1516 4953 1524
rect 4967 1516 5033 1524
rect 5047 1516 5133 1524
rect 5967 1516 6073 1524
rect 2856 1496 3253 1504
rect 3527 1496 3733 1504
rect 4327 1496 4413 1504
rect 4907 1496 4953 1504
rect 4967 1496 5373 1504
rect 5387 1496 5413 1504
rect 727 1476 813 1484
rect 927 1476 1053 1484
rect 1107 1476 1153 1484
rect 1247 1476 1333 1484
rect 1387 1476 1433 1484
rect 1487 1476 2433 1484
rect 3296 1476 3633 1484
rect 3296 1467 3304 1476
rect 4207 1476 4273 1484
rect 4647 1476 4693 1484
rect 5127 1476 5193 1484
rect 5467 1476 5624 1484
rect 567 1456 653 1464
rect 707 1456 873 1464
rect 887 1456 953 1464
rect 967 1456 1364 1464
rect 447 1436 513 1444
rect 527 1437 633 1445
rect 1207 1437 1273 1445
rect 1356 1444 1364 1456
rect 1507 1456 1852 1464
rect 1887 1456 1893 1464
rect 1907 1456 2153 1464
rect 2256 1456 2472 1464
rect 1356 1436 1713 1444
rect 1927 1437 2013 1445
rect 2256 1444 2264 1456
rect 2507 1456 2573 1464
rect 2587 1456 2633 1464
rect 2847 1456 2973 1464
rect 2987 1456 3073 1464
rect 3207 1456 3293 1464
rect 4347 1456 4393 1464
rect 4407 1456 4573 1464
rect 4927 1456 4973 1464
rect 5067 1464 5080 1467
rect 5067 1453 5084 1464
rect 5507 1456 5593 1464
rect 2187 1436 2264 1444
rect 2287 1436 2364 1444
rect 1096 1407 1104 1433
rect 1793 1424 1807 1433
rect 1776 1420 1807 1424
rect 1776 1416 1804 1420
rect 247 1395 333 1403
rect 847 1395 873 1403
rect 1447 1395 1513 1403
rect 1627 1396 1673 1404
rect 1776 1404 1784 1416
rect 1747 1396 1784 1404
rect 1827 1396 1933 1404
rect 2047 1395 2093 1403
rect 707 1376 953 1384
rect 1067 1376 1153 1384
rect 1167 1376 1253 1384
rect 1347 1376 1453 1384
rect 1567 1373 1573 1387
rect 1867 1376 1913 1384
rect 2176 1384 2184 1434
rect 2356 1424 2364 1436
rect 2387 1436 2473 1444
rect 2487 1436 2513 1444
rect 2556 1436 2673 1444
rect 2356 1416 2424 1424
rect 2227 1396 2253 1404
rect 2416 1387 2424 1416
rect 2556 1404 2564 1436
rect 2767 1437 2793 1445
rect 2956 1436 3033 1444
rect 2956 1424 2964 1436
rect 3127 1437 3152 1445
rect 3267 1437 3312 1445
rect 3347 1444 3360 1447
rect 3347 1433 3364 1444
rect 3413 1444 3427 1453
rect 3387 1440 3427 1444
rect 3387 1436 3424 1440
rect 3487 1437 3553 1445
rect 3707 1437 3773 1445
rect 3827 1436 3933 1444
rect 3173 1424 3187 1433
rect 3356 1424 3364 1433
rect 2936 1416 2964 1424
rect 2976 1416 3164 1424
rect 3173 1420 3204 1424
rect 3176 1416 3204 1420
rect 3356 1420 3504 1424
rect 3356 1416 3507 1420
rect 2547 1396 2564 1404
rect 2936 1404 2944 1416
rect 2887 1396 2944 1404
rect 2976 1404 2984 1416
rect 3156 1407 3164 1416
rect 3196 1407 3204 1416
rect 3493 1407 3507 1416
rect 2967 1396 2984 1404
rect 3007 1396 3053 1404
rect 3156 1396 3173 1407
rect 3160 1393 3173 1396
rect 3196 1396 3212 1407
rect 3200 1393 3212 1396
rect 3247 1395 3272 1403
rect 3307 1396 3353 1404
rect 3407 1396 3433 1404
rect 3627 1396 3713 1404
rect 2176 1376 2213 1384
rect 2767 1376 2793 1384
rect 2993 1384 3007 1392
rect 2907 1376 3007 1384
rect 3496 1384 3504 1393
rect 3956 1404 3964 1453
rect 3987 1436 4073 1444
rect 4147 1436 4253 1444
rect 3927 1396 3964 1404
rect 4047 1395 4093 1403
rect 4447 1396 4473 1404
rect 3496 1376 3773 1384
rect 4536 1384 4544 1434
rect 4787 1436 4853 1444
rect 4596 1404 4604 1433
rect 4936 1407 4944 1433
rect 5076 1407 5084 1453
rect 5187 1436 5232 1444
rect 4567 1396 4604 1404
rect 4647 1395 4673 1403
rect 4807 1396 4873 1404
rect 5256 1404 5264 1433
rect 5127 1396 5264 1404
rect 5356 1404 5364 1433
rect 5396 1424 5404 1453
rect 5427 1436 5464 1444
rect 5456 1424 5464 1436
rect 5396 1416 5444 1424
rect 5456 1416 5473 1424
rect 5356 1396 5393 1404
rect 5436 1404 5444 1416
rect 5547 1415 5573 1423
rect 5436 1396 5493 1404
rect 4507 1376 4544 1384
rect 4967 1376 5013 1384
rect 5547 1376 5593 1384
rect 147 1356 313 1364
rect 327 1356 673 1364
rect 727 1356 793 1364
rect 807 1356 933 1364
rect 947 1356 1813 1364
rect 2007 1356 2113 1364
rect 2167 1356 2273 1364
rect 2327 1356 2513 1364
rect 2627 1356 2733 1364
rect 3107 1356 3133 1364
rect 3327 1356 3473 1364
rect 3587 1356 3633 1364
rect 3647 1356 3673 1364
rect 3807 1356 3853 1364
rect 3967 1356 4273 1364
rect 4287 1356 4393 1364
rect 4627 1356 4904 1364
rect 327 1336 473 1344
rect 487 1336 673 1344
rect 1027 1336 1113 1344
rect 2767 1336 2813 1344
rect 2867 1336 2953 1344
rect 2967 1336 3153 1344
rect 3167 1336 3193 1344
rect 3207 1336 3873 1344
rect 4687 1336 4793 1344
rect 4896 1344 4904 1356
rect 4927 1356 5053 1364
rect 5067 1356 5293 1364
rect 5307 1356 5473 1364
rect 5616 1364 5624 1476
rect 5716 1424 5724 1513
rect 5947 1476 6053 1484
rect 5916 1436 6013 1444
rect 5716 1416 5733 1424
rect 5916 1424 5924 1436
rect 5867 1416 5924 1424
rect 6176 1404 6184 1444
rect 6047 1396 6184 1404
rect 5567 1356 5624 1364
rect 4896 1336 4953 1344
rect 5967 1336 6013 1344
rect 127 1316 353 1324
rect 1087 1316 1253 1324
rect 1827 1316 1973 1324
rect 2127 1316 2673 1324
rect 2687 1316 3913 1324
rect 5587 1316 5673 1324
rect 5727 1316 5973 1324
rect 507 1296 853 1304
rect 867 1296 1033 1304
rect 1367 1296 1553 1304
rect 1567 1296 1773 1304
rect 2167 1296 2313 1304
rect 2667 1296 2753 1304
rect 2807 1296 3093 1304
rect 3107 1296 3344 1304
rect 3336 1287 3344 1296
rect 3547 1296 3613 1304
rect 4727 1296 4813 1304
rect 5547 1296 5693 1304
rect 5867 1296 5964 1304
rect 547 1276 713 1284
rect 727 1276 753 1284
rect 1107 1276 1133 1284
rect 1147 1276 1193 1284
rect 2476 1276 2773 1284
rect 2476 1267 2484 1276
rect 3347 1276 3453 1284
rect 4187 1276 4333 1284
rect 5487 1276 5553 1284
rect 5956 1284 5964 1296
rect 5956 1276 6093 1284
rect 207 1256 273 1264
rect 647 1256 813 1264
rect 827 1256 973 1264
rect 1307 1256 1333 1264
rect 1527 1256 1853 1264
rect 2167 1256 2473 1264
rect 2867 1256 3033 1264
rect 3047 1256 3233 1264
rect 3587 1256 3893 1264
rect 3907 1256 3953 1264
rect 4027 1256 4113 1264
rect 5167 1256 5413 1264
rect 567 1236 653 1244
rect 1627 1236 1693 1244
rect 2067 1236 2113 1244
rect 2226 1233 2227 1240
rect 2247 1236 2333 1244
rect 2527 1236 2713 1244
rect 3156 1236 3213 1244
rect 96 1186 104 1233
rect 167 1216 253 1224
rect 267 1216 333 1224
rect 356 1216 373 1224
rect 356 1204 364 1216
rect 236 1196 364 1204
rect 236 1186 244 1196
rect -24 1176 33 1184
rect 147 1175 193 1183
rect 416 1184 424 1214
rect 747 1216 773 1224
rect 840 1224 853 1227
rect 836 1213 853 1224
rect 416 1176 473 1184
rect 836 1186 844 1213
rect 916 1204 924 1214
rect 1047 1216 1093 1224
rect 1136 1216 1293 1224
rect 1136 1204 1144 1216
rect 1316 1216 1433 1224
rect 916 1196 964 1204
rect 1076 1200 1144 1204
rect 527 1176 613 1184
rect 667 1175 713 1183
rect 727 1176 793 1184
rect 956 1184 964 1196
rect 1073 1196 1144 1200
rect 1073 1187 1087 1196
rect 1316 1187 1324 1216
rect 1747 1216 1793 1224
rect 1867 1216 1913 1224
rect 2027 1224 2040 1227
rect 2027 1213 2044 1224
rect 2186 1213 2187 1220
rect 2213 1224 2227 1233
rect 2207 1220 2227 1224
rect 2207 1216 2223 1220
rect 2307 1216 2373 1224
rect 1476 1200 1613 1204
rect 1473 1196 1613 1200
rect 1473 1187 1487 1196
rect 2036 1187 2044 1213
rect 2173 1204 2187 1213
rect 2173 1200 2224 1204
rect 2176 1196 2224 1200
rect 956 1176 993 1184
rect 1387 1175 1413 1183
rect 1807 1175 1833 1183
rect 2216 1186 2224 1196
rect 2396 1186 2404 1233
rect 2436 1216 2553 1224
rect 2436 1186 2444 1216
rect 2647 1216 2733 1224
rect 2927 1217 3073 1225
rect 2816 1187 2824 1214
rect 2127 1175 2153 1183
rect 2267 1175 2293 1183
rect 2807 1176 2824 1187
rect 3096 1186 3104 1233
rect 3127 1216 3144 1224
rect 3136 1187 3144 1216
rect 3156 1204 3164 1236
rect 3427 1236 3493 1244
rect 3507 1236 3533 1244
rect 4247 1236 4513 1244
rect 3367 1216 3393 1224
rect 3156 1196 3184 1204
rect 2807 1173 2820 1176
rect 2887 1175 2913 1183
rect 2927 1176 2973 1184
rect 3176 1167 3184 1196
rect 3196 1184 3204 1213
rect 3256 1196 3333 1204
rect 3256 1186 3264 1196
rect 3473 1204 3487 1213
rect 3736 1216 3813 1224
rect 3473 1200 3524 1204
rect 3476 1196 3524 1200
rect 3196 1176 3213 1184
rect 3427 1175 3493 1183
rect 3516 1184 3524 1196
rect 3516 1176 3553 1184
rect 3607 1175 3633 1183
rect 3736 1184 3744 1216
rect 3867 1216 3944 1224
rect 3936 1186 3944 1216
rect 4007 1216 4053 1224
rect 4167 1216 4213 1224
rect 4287 1216 4404 1224
rect 4396 1186 4404 1216
rect 4436 1186 4444 1236
rect 4687 1216 4713 1224
rect 4727 1219 4773 1227
rect 5067 1216 5312 1224
rect 5347 1216 5373 1224
rect 5527 1217 5553 1225
rect 5707 1216 5744 1224
rect 3707 1176 3744 1184
rect 3987 1175 4033 1183
rect 4496 1184 4504 1213
rect 4816 1187 4824 1213
rect 5453 1204 5467 1213
rect 5453 1200 5613 1204
rect 5456 1196 5613 1200
rect 5687 1197 5713 1205
rect 5736 1204 5744 1216
rect 5936 1216 5993 1224
rect 5736 1196 5873 1204
rect 4496 1176 4533 1184
rect 947 1156 1013 1164
rect 1067 1156 1153 1164
rect 1367 1156 1453 1164
rect 2087 1156 2313 1164
rect 2327 1156 2533 1164
rect 2587 1156 2753 1164
rect 2847 1156 3013 1164
rect 3176 1156 3193 1167
rect 3180 1153 3193 1156
rect 3747 1156 3833 1164
rect 3933 1164 3947 1172
rect 4907 1176 5013 1184
rect 5147 1176 5373 1184
rect 5447 1176 5473 1184
rect 5616 1184 5624 1194
rect 5547 1176 5624 1184
rect 3933 1156 4133 1164
rect 4967 1156 5253 1164
rect 5321 1156 5513 1164
rect 5720 1164 5733 1167
rect 5716 1160 5733 1164
rect 5713 1153 5733 1160
rect 5713 1147 5727 1153
rect 407 1136 553 1144
rect 667 1136 873 1144
rect 3467 1136 3693 1144
rect 3967 1136 4093 1144
rect 4207 1136 4433 1144
rect 4807 1136 5273 1144
rect 1287 1116 1473 1124
rect 4347 1116 4452 1124
rect 4487 1116 4672 1124
rect 4707 1116 5293 1124
rect 5367 1116 5513 1124
rect 47 1096 853 1104
rect 1427 1096 1513 1104
rect 1867 1096 2333 1104
rect 2387 1096 4633 1104
rect 5096 1096 5593 1104
rect 447 1076 833 1084
rect 1127 1076 1273 1084
rect 1627 1076 1913 1084
rect 2047 1076 2333 1084
rect 3967 1076 4293 1084
rect 4367 1076 4693 1084
rect 5096 1084 5104 1096
rect 5936 1087 5944 1216
rect 6067 1216 6124 1224
rect 6027 1196 6104 1204
rect 5976 1144 5984 1193
rect 6096 1167 6104 1196
rect 5976 1136 6009 1144
rect 6116 1144 6124 1216
rect 6023 1136 6024 1144
rect 6116 1136 6164 1144
rect 6067 1116 6133 1124
rect 6156 1087 6164 1136
rect 4767 1076 5104 1084
rect 5127 1076 5153 1084
rect 5167 1076 5853 1084
rect 6147 1076 6164 1087
rect 6147 1073 6160 1076
rect 107 1056 393 1064
rect 867 1056 2373 1064
rect 2527 1056 2633 1064
rect 2647 1056 2673 1064
rect 4347 1056 4553 1064
rect 4967 1056 4993 1064
rect 987 1036 1333 1044
rect 1927 1036 2093 1044
rect 2367 1036 2893 1044
rect 3167 1036 3593 1044
rect 3607 1036 3753 1044
rect 4607 1036 5213 1044
rect 5227 1036 5453 1044
rect 5507 1036 6033 1044
rect 47 1016 413 1024
rect 1647 1016 1693 1024
rect 2176 1016 2453 1024
rect 67 996 153 1004
rect 167 996 313 1004
rect 1007 996 1053 1004
rect 1067 996 1193 1004
rect 1727 996 2073 1004
rect 2176 1004 2184 1016
rect 2536 1016 2793 1024
rect 2087 996 2184 1004
rect 2536 1004 2544 1016
rect 4307 1016 4493 1024
rect 2207 996 2544 1004
rect 3147 996 3553 1004
rect 3567 996 3673 1004
rect 4627 996 4833 1004
rect 4967 996 5084 1004
rect 1087 976 1233 984
rect 1387 976 1573 984
rect 1756 976 1893 984
rect 1756 967 1764 976
rect 2167 976 2553 984
rect 2707 976 2833 984
rect 2847 976 3053 984
rect 3067 976 3833 984
rect 4227 976 4373 984
rect 4787 976 4933 984
rect 5076 984 5084 996
rect 5107 996 5393 1004
rect 5447 996 5493 1004
rect 5727 996 5813 1004
rect 5867 996 5993 1004
rect 5076 976 5153 984
rect 267 956 773 964
rect 1307 956 1333 964
rect 1647 956 1753 964
rect 2007 956 2133 964
rect 2187 956 2453 964
rect 2467 956 2533 964
rect 2907 956 2993 964
rect 3127 956 4033 964
rect 4267 956 4333 964
rect 4687 956 4713 964
rect 4967 956 5193 964
rect 5307 956 5333 964
rect 5727 956 5853 964
rect 87 936 213 944
rect 407 936 633 944
rect 867 936 1033 944
rect 1047 936 1093 944
rect 1107 936 1153 944
rect 1587 936 1653 944
rect 1667 936 1933 944
rect 3267 936 3353 944
rect 3667 936 3713 944
rect 3856 936 4153 944
rect 180 924 193 927
rect 176 913 193 924
rect 907 916 1013 924
rect 1347 917 1373 925
rect 1547 916 1633 924
rect 1727 917 1753 925
rect 2047 917 2233 925
rect 176 887 184 913
rect 376 887 384 914
rect 247 875 313 883
rect 367 876 384 887
rect 367 873 380 876
rect 487 875 533 883
rect 696 884 704 914
rect 2407 916 2433 924
rect 2567 916 2664 924
rect 587 876 704 884
rect 787 876 833 884
rect 947 875 1133 883
rect 1247 875 1313 883
rect 1527 875 1573 883
rect 1667 876 1693 884
rect 1707 875 1733 883
rect 1847 875 1913 883
rect 1967 875 1993 883
rect 2107 875 2153 883
rect 2296 884 2304 913
rect 2296 876 2373 884
rect 2656 886 2664 916
rect 2967 916 3113 924
rect 3327 917 3393 925
rect 3696 916 3753 924
rect 3576 896 3633 904
rect 3576 886 3584 896
rect 3696 886 3704 916
rect 3856 886 3864 936
rect 4987 936 5052 944
rect 5087 936 5112 944
rect 5367 936 5553 944
rect 3887 916 3993 924
rect 4067 917 4113 925
rect 4207 916 4293 924
rect 4387 924 4400 927
rect 4387 913 4404 924
rect 4507 916 4544 924
rect 2467 876 2533 884
rect 2767 875 2933 883
rect 3067 875 3093 883
rect 3187 875 3273 883
rect 3347 875 3373 883
rect 3467 875 3533 883
rect 3907 876 3953 884
rect 4027 875 4052 883
rect 4107 876 4193 884
rect 4287 876 4333 884
rect 4396 886 4404 913
rect 4536 886 4544 916
rect 4647 917 4673 925
rect 5007 916 5033 924
rect 4587 876 4633 884
rect 4707 876 4753 884
rect 4876 884 4884 914
rect 5133 924 5147 933
rect 5087 920 5147 924
rect 5087 916 5144 920
rect 5296 904 5304 914
rect 5347 916 5693 924
rect 6007 916 6184 924
rect 5296 896 5473 904
rect 4876 876 4973 884
rect 5047 875 5173 883
rect 5227 875 5273 883
rect 5367 876 5413 884
rect 67 856 133 864
rect 967 856 1033 864
rect 1733 864 1747 872
rect 1733 856 2053 864
rect 2607 856 2633 864
rect 4056 864 4064 872
rect 4056 856 4233 864
rect 5173 864 5187 872
rect 5173 856 5453 864
rect 5467 856 5613 864
rect 5627 856 5733 864
rect 447 836 613 844
rect 827 836 873 844
rect 887 836 1393 844
rect 3147 836 3513 844
rect 4647 836 4773 844
rect 4827 836 5033 844
rect 1747 816 1953 824
rect 2267 816 2473 824
rect 2987 816 3553 824
rect 3607 816 3733 824
rect 4067 816 4613 824
rect 1107 796 1153 804
rect 1527 796 2073 804
rect 2087 796 2153 804
rect 2167 796 2393 804
rect 2667 796 3133 804
rect 4467 796 4733 804
rect 5107 796 5233 804
rect 5527 796 5913 804
rect 287 776 353 784
rect 367 776 573 784
rect 807 776 933 784
rect 1667 776 1773 784
rect 1827 776 1932 784
rect 1967 776 2193 784
rect 3187 776 3233 784
rect 3247 776 3633 784
rect 3807 776 4093 784
rect 4327 776 4573 784
rect 4827 776 5273 784
rect 67 756 393 764
rect 407 756 533 764
rect 547 756 713 764
rect 1927 756 2373 764
rect 2387 756 2553 764
rect 2567 756 2693 764
rect 4027 756 4253 764
rect 5647 756 5713 764
rect 127 736 193 744
rect 567 736 613 744
rect 767 736 832 744
rect 867 736 1093 744
rect 1187 736 1233 744
rect 1307 736 1813 744
rect 2007 736 2193 744
rect 2207 736 2253 744
rect 2307 736 2353 744
rect 2447 736 2693 744
rect 3027 736 3213 744
rect 3267 736 3353 744
rect 3367 736 3413 744
rect 3567 736 3613 744
rect 3867 736 4073 744
rect 4087 736 4133 744
rect 4487 736 4573 744
rect 5087 736 5133 744
rect 5287 736 5552 744
rect 5587 736 5613 744
rect 47 716 93 724
rect 1847 716 2213 724
rect 2227 716 2413 724
rect 2427 716 2464 724
rect 187 697 393 705
rect 447 696 493 704
rect 547 704 560 707
rect 547 693 564 704
rect 647 696 673 704
rect 736 696 813 704
rect 556 666 564 693
rect 736 666 744 696
rect 876 696 893 704
rect 876 667 884 696
rect 947 697 993 705
rect 67 655 93 663
rect 327 655 353 663
rect 1056 664 1064 694
rect 1147 696 1193 704
rect 1273 704 1287 713
rect 1247 700 1287 704
rect 1247 696 1284 700
rect 1296 696 1353 704
rect 1296 684 1304 696
rect 1407 696 1424 704
rect 1256 676 1304 684
rect 1256 666 1264 676
rect 1416 667 1424 696
rect 1487 696 1553 704
rect 927 656 1064 664
rect 1307 655 1373 663
rect 1656 664 1664 694
rect 1767 696 1793 704
rect 1927 704 1940 707
rect 1927 693 1944 704
rect 2067 696 2113 704
rect 1587 656 1664 664
rect 1687 656 1733 664
rect 1936 666 1944 693
rect 1787 656 1853 664
rect 2227 655 2273 663
rect 2376 664 2384 693
rect 2456 666 2464 716
rect 2727 716 2993 724
rect 3687 716 3733 724
rect 4307 716 4353 724
rect 4707 716 4773 724
rect 4987 716 5093 724
rect 5476 716 5653 724
rect 2607 696 2973 704
rect 2473 684 2487 693
rect 2473 680 2544 684
rect 2476 676 2544 680
rect 2536 666 2544 676
rect 2696 666 2704 696
rect 3407 696 3433 704
rect 3096 684 3104 694
rect 3396 684 3404 694
rect 3627 696 3684 704
rect 3096 676 3264 684
rect 2327 656 2384 664
rect 2827 656 2853 664
rect 3007 655 3033 663
rect 3207 655 3233 663
rect 3256 664 3264 676
rect 3376 676 3404 684
rect 3676 684 3684 696
rect 3767 696 3813 704
rect 5476 708 5484 716
rect 5667 716 5753 724
rect 3676 676 3704 684
rect 3376 664 3384 676
rect 3256 656 3384 664
rect 3547 656 3593 664
rect 3696 666 3704 676
rect 4196 684 4204 695
rect 4407 696 4453 704
rect 4840 704 4852 707
rect 4127 676 4204 684
rect 4236 680 4324 684
rect 4233 676 4324 680
rect 4233 667 4247 676
rect 3607 656 3653 664
rect 3747 655 3833 663
rect 4007 655 4073 663
rect 4316 666 4324 676
rect 4496 667 4504 694
rect 4327 655 4413 663
rect 4487 656 4504 667
rect 4836 693 4852 704
rect 4887 697 4933 705
rect 5047 696 5273 704
rect 5327 697 5393 705
rect 5447 697 5473 705
rect 5536 696 5613 704
rect 4836 666 4844 693
rect 5536 666 5544 696
rect 5676 696 5973 704
rect 5676 667 5684 696
rect 4487 653 4500 656
rect 5127 656 5253 664
rect 336 636 413 644
rect 47 616 133 624
rect 336 624 344 636
rect 607 636 673 644
rect 1296 644 1304 652
rect 1227 636 1304 644
rect 1507 636 1753 644
rect 2107 636 2193 644
rect 3447 636 3484 644
rect 147 616 344 624
rect 367 616 453 624
rect 787 616 1153 624
rect 1487 616 1633 624
rect 2427 616 2493 624
rect 2927 616 3273 624
rect 3287 616 3333 624
rect 3476 624 3484 636
rect 4527 636 4653 644
rect 4827 636 4873 644
rect 5067 636 5373 644
rect 5787 636 5993 644
rect 3476 616 3873 624
rect 3887 616 3913 624
rect 4467 616 4613 624
rect 4987 616 5213 624
rect 927 596 1493 604
rect 1987 596 2133 604
rect 2416 604 2424 613
rect 2147 596 2424 604
rect 2987 596 3133 604
rect 3387 596 3453 604
rect 3467 596 3493 604
rect 4107 596 4593 604
rect 5267 596 5573 604
rect 5587 596 5653 604
rect 287 576 593 584
rect 847 576 953 584
rect 967 576 1073 584
rect 1667 576 1893 584
rect 2747 576 2953 584
rect 4167 576 4473 584
rect 4747 576 4993 584
rect 5467 576 5873 584
rect 1627 556 2033 564
rect 2287 556 2653 564
rect 3127 556 3373 564
rect 4607 556 5013 564
rect 5507 556 5713 564
rect 887 536 1213 544
rect 1827 536 2013 544
rect 2367 536 2573 544
rect 4587 536 5693 544
rect 5787 536 5933 544
rect 1007 516 1093 524
rect 1107 516 1133 524
rect 2047 516 2653 524
rect 2667 516 3373 524
rect 3707 516 4113 524
rect 4127 516 4373 524
rect 427 496 553 504
rect 567 496 953 504
rect 1047 496 1173 504
rect 1387 496 1693 504
rect 4507 496 5153 504
rect 5387 496 5413 504
rect 5787 496 6013 504
rect 6027 496 6113 504
rect 127 476 253 484
rect 267 476 793 484
rect 1867 476 2353 484
rect 3487 476 3693 484
rect 4327 476 4973 484
rect 5607 476 5793 484
rect 867 456 893 464
rect 907 456 933 464
rect 1187 456 1273 464
rect 1287 456 1413 464
rect 1727 456 1813 464
rect 2767 456 3193 464
rect 3287 456 3573 464
rect 3787 456 4353 464
rect 5567 456 5733 464
rect 507 436 613 444
rect 1587 436 1973 444
rect 2387 436 2453 444
rect 2627 436 2833 444
rect 2847 436 2853 444
rect 2867 436 3013 444
rect 3087 436 3213 444
rect 3827 436 3973 444
rect 3987 436 4153 444
rect 5067 436 5153 444
rect 5947 436 6073 444
rect 167 416 213 424
rect 227 416 313 424
rect 1176 416 1393 424
rect 156 396 193 404
rect 156 364 164 396
rect 436 396 513 404
rect 436 366 444 396
rect 647 397 693 405
rect 147 356 164 364
rect 587 356 633 364
rect 736 364 744 394
rect 1116 367 1124 393
rect 1176 384 1184 416
rect 2456 424 2464 433
rect 2456 416 3053 424
rect 3067 416 3153 424
rect 3267 416 3293 424
rect 3547 416 3633 424
rect 3647 416 3713 424
rect 4407 416 4713 424
rect 5447 416 5493 424
rect 5507 416 5613 424
rect 5827 416 5873 424
rect 1200 404 1213 407
rect 1156 376 1184 384
rect 1196 393 1213 404
rect 1327 397 1473 405
rect 1556 396 1653 404
rect 687 356 744 364
rect 807 356 833 364
rect 967 356 1013 364
rect 1156 366 1164 376
rect 1196 366 1204 393
rect 1556 384 1564 396
rect 1747 397 1773 405
rect 1867 396 1933 404
rect 2213 405 2227 413
rect 2067 397 2233 405
rect 2216 396 2224 397
rect 2587 396 2753 404
rect 3247 397 3413 405
rect 3767 397 3853 405
rect 3867 396 3933 404
rect 1427 376 1564 384
rect 1936 384 1944 394
rect 2416 384 2424 394
rect 4047 396 4113 404
rect 4127 396 4213 404
rect 4267 397 4293 405
rect 4447 396 4533 404
rect 4787 399 4853 407
rect 1936 376 2744 384
rect 1207 356 1253 364
rect 1847 356 1953 364
rect 1976 364 1984 376
rect 1976 356 2093 364
rect 2147 355 2172 363
rect 2207 355 2253 363
rect 2307 356 2373 364
rect 2487 356 2553 364
rect 2567 356 2613 364
rect 2736 366 2744 376
rect 2807 376 2973 384
rect 2667 356 2693 364
rect 2747 356 2853 364
rect 3047 356 3233 364
rect 3407 355 3473 363
rect 3647 355 3673 363
rect 4007 356 4193 364
rect 4247 356 4313 364
rect 5036 366 5044 413
rect 5107 396 5193 404
rect 5680 404 5693 407
rect 5676 393 5693 404
rect 5987 397 6093 405
rect 5256 376 5593 384
rect 4567 356 4593 364
rect 667 336 713 344
rect 1407 336 1733 344
rect 1953 344 1967 352
rect 5256 364 5264 376
rect 5676 364 5684 393
rect 5787 355 5873 363
rect 5927 355 6033 363
rect 1953 336 2033 344
rect 2767 336 2793 344
rect 3087 336 3133 344
rect 3147 336 3213 344
rect 3707 336 3833 344
rect 3847 336 3953 344
rect 4427 336 4813 344
rect 4827 336 5073 344
rect 5087 336 5133 344
rect 247 316 313 324
rect 407 316 673 324
rect 687 316 813 324
rect 947 316 1113 324
rect 1287 316 1373 324
rect 2087 316 2833 324
rect 3187 316 3233 324
rect 3327 316 3353 324
rect 3367 316 3433 324
rect 3447 316 3653 324
rect 3667 316 3753 324
rect 3947 316 4053 324
rect 4387 316 4673 324
rect 5967 316 6013 324
rect 547 296 613 304
rect 1507 296 1733 304
rect 1787 296 2713 304
rect 3047 296 3253 304
rect 3527 296 3573 304
rect 5727 296 5773 304
rect 5827 296 6133 304
rect 107 276 133 284
rect 147 276 493 284
rect 507 276 653 284
rect 927 276 1233 284
rect 1547 276 1713 284
rect 1727 276 1993 284
rect 2607 276 2813 284
rect 2907 276 3233 284
rect 3287 276 3553 284
rect 5987 276 6053 284
rect 547 256 733 264
rect 847 256 893 264
rect 1007 256 1053 264
rect 1067 256 1473 264
rect 1516 256 2013 264
rect 1516 247 1524 256
rect 2027 256 2113 264
rect 2567 256 3213 264
rect 3267 256 3793 264
rect 3807 256 4093 264
rect 4107 256 4353 264
rect 4927 256 5013 264
rect 5167 256 5193 264
rect 27 236 93 244
rect 287 236 413 244
rect 1107 236 1173 244
rect 1307 236 1513 244
rect 2267 236 2433 244
rect 2616 236 3413 244
rect 267 216 593 224
rect 607 216 753 224
rect 767 216 873 224
rect 887 216 1633 224
rect 1707 216 1793 224
rect 2007 216 2093 224
rect 2227 216 2413 224
rect 2616 224 2624 236
rect 3427 236 3533 244
rect 2467 216 2624 224
rect 2687 216 3373 224
rect 3567 216 3733 224
rect 3747 216 3833 224
rect 4047 216 4244 224
rect 1667 196 1953 204
rect 1967 196 2173 204
rect 2447 196 2633 204
rect 2920 204 2933 207
rect 2916 196 2933 204
rect 2920 193 2933 196
rect 2947 196 3064 204
rect 116 176 273 184
rect 116 146 124 176
rect 327 176 373 184
rect 396 146 404 193
rect 427 176 793 184
rect 816 146 824 193
rect 860 184 873 187
rect 856 173 873 184
rect 1007 176 1084 184
rect 856 146 864 173
rect 1076 164 1084 176
rect 1127 176 1153 184
rect 1347 177 1393 185
rect 1447 176 1613 184
rect 1747 176 1853 184
rect 1907 176 1933 184
rect 1956 176 2053 184
rect 1956 164 1964 176
rect 2307 177 2353 185
rect 2487 177 2533 185
rect 2756 176 2893 184
rect 2756 164 2764 176
rect 2987 176 3033 184
rect 927 156 1064 164
rect 1076 156 1104 164
rect 167 136 233 144
rect 247 136 353 144
rect 607 135 633 143
rect 1056 146 1064 156
rect 947 136 973 144
rect 1096 144 1104 156
rect 1876 156 3024 164
rect 1876 146 1884 156
rect 3016 146 3024 156
rect 3056 146 3064 196
rect 3087 176 3133 184
rect 3387 176 3553 184
rect 3640 184 3653 187
rect 3167 156 3244 164
rect 3236 146 3244 156
rect 1096 136 1213 144
rect 1427 135 1473 143
rect 1527 135 1553 143
rect 1727 136 1833 144
rect 1967 135 1993 143
rect 2047 135 2073 143
rect 2127 135 2153 143
rect 2207 135 2253 143
rect 2327 136 2613 144
rect 2687 135 2733 143
rect 2847 135 2873 143
rect 2927 135 2973 143
rect 3147 135 3193 143
rect 3407 136 3513 144
rect 353 124 367 132
rect 353 116 473 124
rect 527 116 559 124
rect 1287 116 1373 124
rect 1873 124 1887 132
rect 1767 116 1887 124
rect 2427 116 2533 124
rect 2547 116 2573 124
rect 2613 124 2627 132
rect 2613 116 2773 124
rect 3547 116 3593 124
rect 3616 124 3624 174
rect 3636 173 3653 184
rect 4133 184 4147 193
rect 4107 180 4147 184
rect 4107 176 4144 180
rect 4167 177 4213 185
rect 3636 146 3644 173
rect 3776 164 3784 174
rect 3707 156 3784 164
rect 4236 146 4244 216
rect 4847 216 4953 224
rect 5227 216 5373 224
rect 4267 176 4313 184
rect 4407 177 4433 185
rect 4567 177 4633 185
rect 4927 176 5013 184
rect 5307 176 5373 184
rect 5527 177 5593 185
rect 4736 156 4864 164
rect 3807 135 4033 143
rect 4087 136 4193 144
rect 4387 136 4493 144
rect 4736 144 4744 156
rect 4856 144 4864 156
rect 4807 133 4832 141
rect 4867 133 5113 141
rect 5187 133 5213 141
rect 5867 135 5933 143
rect 3616 116 3684 124
rect 907 96 1213 104
rect 1267 96 1593 104
rect 1607 96 1653 104
rect 1947 96 2353 104
rect 2367 96 2453 104
rect 3007 96 3153 104
rect 3676 104 3684 116
rect 4327 116 4413 124
rect 3676 96 3693 104
rect 3707 96 4113 104
rect 4127 96 4153 104
rect 4227 96 4433 104
rect 747 76 1493 84
rect 1807 76 2344 84
rect 327 56 1713 64
rect 2336 64 2344 76
rect 3207 76 4073 84
rect 2336 56 2413 64
rect 2827 56 4013 64
rect 4307 56 4533 64
rect 767 36 1333 44
rect 2147 36 2773 44
rect 2867 36 3393 44
rect 3467 36 3753 44
use INVX1  _889_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 5390 0 -1 1830
box -12 -8 72 272
use NOR2X1  _890_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 5070 0 1 1310
box -12 -8 92 272
use NAND2X1  _891_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 5190 0 1 1310
box -12 -8 92 272
use INVX1  _892_
timestamp 1727136778
transform 1 0 5410 0 -1 1310
box -12 -8 72 272
use INVX1  _893_
timestamp 1727136778
transform -1 0 5310 0 1 1310
box -12 -8 72 272
use INVX2  _894_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 5530 0 -1 1310
box -12 -8 72 272
use NOR2X1  _895_
timestamp 1727136778
transform -1 0 5330 0 -1 1830
box -12 -8 92 272
use NAND2X1  _896_
timestamp 1727136778
transform -1 0 5210 0 -1 1830
box -12 -8 92 272
use INVX1  _897_
timestamp 1727136778
transform 1 0 5150 0 1 2350
box -12 -8 72 272
use NOR2X1  _898_
timestamp 1727136778
transform -1 0 5570 0 -1 1830
box -12 -8 92 272
use AOI21X1  _899_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 5290 0 1 1830
box -12 -8 112 272
use NOR2X1  _900_
timestamp 1727136778
transform -1 0 5950 0 1 2350
box -12 -8 92 272
use OAI21X1  _901_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 5810 0 1 2350
box -12 -8 112 272
use INVX1  _902_
timestamp 1727136778
transform 1 0 5830 0 -1 2350
box -12 -8 72 272
use INVX4  _903_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 4930 0 1 1830
box -12 -8 92 272
use OAI21X1  _904_
timestamp 1727136778
transform -1 0 5450 0 1 1310
box -12 -8 112 272
use INVX1  _905_
timestamp 1727136778
transform -1 0 5770 0 -1 2350
box -12 -8 72 272
use NOR2X1  _906_
timestamp 1727136778
transform -1 0 4310 0 -1 2350
box -12 -8 92 272
use INVX1  _907_
timestamp 1727136778
transform 1 0 5010 0 -1 2350
box -12 -8 72 272
use INVX1  _908_
timestamp 1727136778
transform 1 0 5990 0 -1 2870
box -12 -8 72 272
use OAI21X1  _909_
timestamp 1727136778
transform 1 0 5630 0 1 1830
box -12 -8 112 272
use OAI21X1  _910_
timestamp 1727136778
transform 1 0 5550 0 -1 2350
box -12 -8 112 272
use AOI22X1  _911_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 5450 0 1 1830
box -14 -8 132 272
use NAND2X1  _912_
timestamp 1727136778
transform 1 0 5790 0 1 1830
box -12 -8 92 272
use OAI21X1  _913_
timestamp 1727136778
transform -1 0 5670 0 1 2350
box -12 -8 112 272
use OAI21X1  _914_
timestamp 1727136778
transform -1 0 5370 0 1 2350
box -12 -8 112 272
use NAND2X1  _915_
timestamp 1727136778
transform 1 0 5270 0 -1 2350
box -12 -8 92 272
use NOR2X1  _916_
timestamp 1727136778
transform -1 0 5730 0 1 2870
box -12 -8 92 272
use NOR2X1  _917_
timestamp 1727136778
transform 1 0 5850 0 -1 2870
box -12 -8 92 272
use OAI22X1  _918_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 5530 0 -1 2870
box -12 -8 132 272
use OR2X2  _919_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 5430 0 1 2350
box -12 -8 112 272
use INVX1  _920_
timestamp 1727136778
transform -1 0 5630 0 -1 2870
box -12 -8 72 272
use AOI22X1  _921_
timestamp 1727136778
transform 1 0 5690 0 -1 2870
box -14 -8 132 272
use NAND3X1  _922_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 5410 0 -1 2350
box -12 -8 112 272
use AND2X2  _923_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 5930 0 -1 2350
box -12 -8 112 273
use OAI21X1  _924_
timestamp 1727136778
transform 1 0 5930 0 1 1830
box -12 -8 112 272
use INVX1  _925_
timestamp 1727136778
transform -1 0 6050 0 1 1310
box -12 -8 72 272
use INVX1  _926_
timestamp 1727136778
transform -1 0 4390 0 1 4430
box -12 -8 72 272
use NAND2X1  _927_
timestamp 1727136778
transform 1 0 4890 0 -1 3390
box -12 -8 92 272
use OAI21X1  _928_
timestamp 1727136778
transform 1 0 4730 0 -1 3390
box -12 -8 112 272
use INVX1  _929_
timestamp 1727136778
transform 1 0 4230 0 1 4430
box -12 -8 72 272
use NAND2X1  _930_
timestamp 1727136778
transform 1 0 3710 0 1 3910
box -12 -8 92 272
use OAI21X1  _931_
timestamp 1727136778
transform -1 0 3950 0 1 3910
box -12 -8 112 272
use INVX1  _932_
timestamp 1727136778
transform 1 0 4150 0 -1 4430
box -12 -8 72 272
use NAND2X1  _933_
timestamp 1727136778
transform -1 0 4510 0 -1 3390
box -12 -8 92 272
use OAI21X1  _934_
timestamp 1727136778
transform 1 0 4570 0 -1 3390
box -12 -8 112 272
use INVX1  _935_
timestamp 1727136778
transform -1 0 5450 0 1 4950
box -12 -8 72 272
use NAND2X1  _936_
timestamp 1727136778
transform 1 0 4110 0 1 4430
box -12 -8 92 272
use OAI21X1  _937_
timestamp 1727136778
transform -1 0 4110 0 -1 4430
box -12 -8 112 272
use INVX1  _938_
timestamp 1727136778
transform -1 0 4050 0 -1 5470
box -12 -8 72 272
use NAND2X1  _939_
timestamp 1727136778
transform 1 0 3690 0 1 4430
box -12 -8 92 272
use OAI21X1  _940_
timestamp 1727136778
transform 1 0 3490 0 -1 4430
box -12 -8 112 272
use INVX1  _941_
timestamp 1727136778
transform -1 0 3330 0 -1 4950
box -12 -8 72 272
use NAND2X1  _942_
timestamp 1727136778
transform 1 0 3650 0 -1 3910
box -12 -8 92 272
use OAI21X1  _943_
timestamp 1727136778
transform 1 0 3510 0 -1 3910
box -12 -8 112 272
use INVX1  _944_
timestamp 1727136778
transform -1 0 5390 0 1 3390
box -12 -8 72 272
use NAND2X1  _945_
timestamp 1727136778
transform 1 0 5590 0 -1 3390
box -12 -8 92 272
use OAI21X1  _946_
timestamp 1727136778
transform 1 0 5450 0 -1 3390
box -12 -8 112 272
use INVX4  _947_
timestamp 1727136778
transform 1 0 5690 0 1 790
box -12 -8 92 272
use NAND2X1  _948_
timestamp 1727136778
transform 1 0 5270 0 -1 2870
box -12 -8 92 272
use OAI21X1  _949_
timestamp 1727136778
transform 1 0 5130 0 -1 2870
box -12 -8 112 272
use INVX1  _950_
timestamp 1727136778
transform -1 0 4730 0 1 1830
box -12 -8 72 272
use INVX1  _951_
timestamp 1727136778
transform 1 0 3930 0 -1 1830
box -12 -8 72 272
use INVX2  _952_
timestamp 1727136778
transform 1 0 2370 0 1 3390
box -12 -8 72 272
use NOR2X1  _953_
timestamp 1727136778
transform 1 0 2670 0 -1 1310
box -12 -8 92 272
use AND2X2  _954_
timestamp 1727136778
transform -1 0 2590 0 1 1310
box -12 -8 112 273
use NAND2X1  _955_
timestamp 1727136778
transform 1 0 2790 0 1 790
box -12 -8 92 272
use NAND2X1  _956_
timestamp 1727136778
transform 1 0 3210 0 1 1830
box -12 -8 92 272
use NAND2X1  _957_
timestamp 1727136778
transform 1 0 3510 0 -1 1830
box -12 -8 92 272
use OR2X2  _958_
timestamp 1727136778
transform 1 0 3650 0 -1 1830
box -12 -8 112 272
use NAND2X1  _959_
timestamp 1727136778
transform 1 0 3650 0 1 1310
box -12 -8 92 272
use AND2X2  _960_
timestamp 1727136778
transform 1 0 3190 0 1 1310
box -12 -8 112 273
use OAI21X1  _961_
timestamp 1727136778
transform -1 0 3590 0 1 1310
box -12 -8 112 272
use NAND2X1  _962_
timestamp 1727136778
transform 1 0 3810 0 -1 1830
box -12 -8 92 272
use INVX1  _963_
timestamp 1727136778
transform 1 0 2950 0 -1 1310
box -12 -8 72 272
use NAND2X1  _964_
timestamp 1727136778
transform -1 0 2730 0 1 1830
box -12 -8 92 272
use NAND2X1  _965_
timestamp 1727136778
transform 1 0 2530 0 1 1830
box -12 -8 92 272
use OR2X2  _966_
timestamp 1727136778
transform 1 0 3370 0 -1 1830
box -12 -8 112 272
use INVX1  _967_
timestamp 1727136778
transform -1 0 2990 0 1 1830
box -12 -8 72 272
use INVX1  _968_
timestamp 1727136778
transform 1 0 2610 0 1 3390
box -12 -8 72 272
use OAI21X1  _969_
timestamp 1727136778
transform -1 0 2890 0 1 1830
box -12 -8 112 272
use NAND3X1  _970_
timestamp 1727136778
transform 1 0 3050 0 -1 1310
box -12 -8 112 272
use NOR2X1  _971_
timestamp 1727136778
transform 1 0 3070 0 -1 1830
box -12 -8 92 272
use AND2X2  _972_
timestamp 1727136778
transform -1 0 3310 0 -1 1830
box -12 -8 112 273
use OAI21X1  _973_
timestamp 1727136778
transform 1 0 3050 0 1 1310
box -12 -8 112 272
use NAND3X1  _974_
timestamp 1727136778
transform -1 0 3610 0 1 790
box -12 -8 112 272
use INVX1  _975_
timestamp 1727136778
transform 1 0 3090 0 1 790
box -12 -8 72 272
use NAND2X1  _976_
timestamp 1727136778
transform 1 0 2630 0 1 1310
box -12 -8 92 272
use INVX2  _977_
timestamp 1727136778
transform 1 0 2150 0 1 3910
box -12 -8 72 272
use NAND2X1  _978_
timestamp 1727136778
transform 1 0 2530 0 -1 1830
box -12 -8 92 272
use OAI21X1  _979_
timestamp 1727136778
transform 1 0 2110 0 1 1310
box -12 -8 112 272
use OAI21X1  _980_
timestamp 1727136778
transform 1 0 2930 0 1 790
box -12 -8 112 272
use AOI21X1  _981_
timestamp 1727136778
transform 1 0 3670 0 1 790
box -12 -8 112 272
use OAI21X1  _982_
timestamp 1727136778
transform -1 0 3570 0 -1 790
box -12 -8 112 272
use OAI21X1  _983_
timestamp 1727136778
transform -1 0 2870 0 1 1310
box -12 -8 112 272
use AND2X2  _984_
timestamp 1727136778
transform -1 0 2550 0 -1 2350
box -12 -8 112 273
use NAND3X1  _985_
timestamp 1727136778
transform -1 0 2470 0 1 1830
box -12 -8 112 272
use AOI22X1  _986_
timestamp 1727136778
transform -1 0 1850 0 -1 2350
box -14 -8 132 272
use INVX1  _987_
timestamp 1727136778
transform -1 0 1670 0 1 790
box -12 -8 72 272
use NAND2X1  _988_
timestamp 1727136778
transform -1 0 1470 0 1 1310
box -12 -8 92 272
use INVX1  _989_
timestamp 1727136778
transform -1 0 1870 0 -1 1310
box -12 -8 72 272
use NAND3X1  _990_
timestamp 1727136778
transform 1 0 1890 0 1 790
box -12 -8 112 272
use NAND2X1  _991_
timestamp 1727136778
transform 1 0 2430 0 1 3910
box -12 -8 92 272
use NOR2X1  _992_
timestamp 1727136778
transform -1 0 2470 0 -1 1830
box -12 -8 92 272
use OAI21X1  _993_
timestamp 1727136778
transform 1 0 2050 0 1 790
box -12 -8 112 272
use NAND3X1  _994_
timestamp 1727136778
transform 1 0 2630 0 1 790
box -12 -8 112 272
use AOI21X1  _995_
timestamp 1727136778
transform -1 0 2890 0 -1 1310
box -12 -8 112 272
use OAI21X1  _996_
timestamp 1727136778
transform 1 0 1730 0 1 790
box -12 -8 112 272
use NAND3X1  _997_
timestamp 1727136778
transform -1 0 1550 0 1 790
box -12 -8 112 272
use NAND3X1  _998_
timestamp 1727136778
transform 1 0 1630 0 -1 790
box -12 -8 112 272
use NAND2X1  _999_
timestamp 1727136778
transform 1 0 2230 0 1 1830
box -12 -8 92 272
use INVX1  _1000_
timestamp 1727136778
transform 1 0 2250 0 1 1310
box -12 -8 72 272
use AND2X2  _1001_
timestamp 1727136778
transform 1 0 2810 0 -1 1830
box -12 -8 112 273
use NAND2X1  _1002_
timestamp 1727136778
transform 1 0 2370 0 1 1310
box -12 -8 92 272
use INVX1  _1003_
timestamp 1727136778
transform -1 0 3010 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1004_
timestamp 1727136778
transform 1 0 2510 0 -1 1310
box -12 -8 112 272
use NAND3X1  _1005_
timestamp 1727136778
transform -1 0 2450 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1006_
timestamp 1727136778
transform 1 0 2050 0 -1 1310
box -12 -8 112 272
use INVX1  _1007_
timestamp 1727136778
transform -1 0 1750 0 1 1310
box -12 -8 72 272
use OAI21X1  _1008_
timestamp 1727136778
transform 1 0 1810 0 1 1310
box -12 -8 112 272
use NAND3X1  _1009_
timestamp 1727136778
transform -1 0 2070 0 1 1310
box -12 -8 112 272
use AND2X2  _1010_
timestamp 1727136778
transform 1 0 2330 0 1 790
box -12 -8 112 273
use NAND3X1  _1011_
timestamp 1727136778
transform -1 0 2330 0 -1 790
box -12 -8 112 272
use AOI21X1  _1012_
timestamp 1727136778
transform -1 0 1590 0 -1 790
box -12 -8 112 272
use AOI21X1  _1013_
timestamp 1727136778
transform -1 0 2570 0 1 790
box -12 -8 112 272
use NAND2X1  _1014_
timestamp 1727136778
transform -1 0 2290 0 1 790
box -12 -8 92 272
use OAI21X1  _1015_
timestamp 1727136778
transform -1 0 2170 0 -1 790
box -12 -8 112 272
use NAND3X1  _1016_
timestamp 1727136778
transform -1 0 2170 0 1 270
box -12 -8 112 272
use AOI21X1  _1017_
timestamp 1727136778
transform 1 0 2230 0 1 270
box -12 -8 112 272
use OAI21X1  _1018_
timestamp 1727136778
transform -1 0 2490 0 1 270
box -12 -8 112 272
use AOI21X1  _1019_
timestamp 1727136778
transform -1 0 1870 0 -1 790
box -12 -8 112 272
use OAI21X1  _1020_
timestamp 1727136778
transform -1 0 1630 0 1 1310
box -12 -8 112 272
use AND2X2  _1021_
timestamp 1727136778
transform -1 0 1550 0 1 3910
box -12 -8 112 273
use NAND2X1  _1022_
timestamp 1727136778
transform -1 0 1470 0 1 1830
box -12 -8 92 272
use INVX1  _1023_
timestamp 1727136778
transform 1 0 1170 0 1 2350
box -12 -8 72 272
use INVX2  _1024_
timestamp 1727136778
transform 1 0 1530 0 -1 4950
box -12 -8 72 272
use NAND2X1  _1025_
timestamp 1727136778
transform 1 0 1470 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1026_
timestamp 1727136778
transform 1 0 1290 0 1 2350
box -12 -8 112 272
use NAND2X1  _1027_
timestamp 1727136778
transform 1 0 1530 0 1 1830
box -12 -8 92 272
use INVX1  _1028_
timestamp 1727136778
transform 1 0 1070 0 -1 1830
box -12 -8 72 272
use NAND3X1  _1029_
timestamp 1727136778
transform -1 0 1030 0 -1 1830
box -12 -8 112 272
use NOR2X1  _1030_
timestamp 1727136778
transform -1 0 1690 0 -1 2350
box -12 -8 92 272
use AOI22X1  _1031_
timestamp 1727136778
transform 1 0 1310 0 -1 2350
box -14 -8 132 272
use OAI21X1  _1032_
timestamp 1727136778
transform -1 0 1350 0 1 1830
box -12 -8 112 272
use AOI21X1  _1033_
timestamp 1727136778
transform -1 0 1190 0 1 1310
box -12 -8 112 272
use AOI21X1  _1034_
timestamp 1727136778
transform -1 0 1770 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1035_
timestamp 1727136778
transform -1 0 1190 0 1 1830
box -12 -8 112 272
use NAND3X1  _1036_
timestamp 1727136778
transform -1 0 1290 0 -1 1830
box -12 -8 112 272
use AOI21X1  _1037_
timestamp 1727136778
transform -1 0 1170 0 -1 1310
box -12 -8 112 272
use NAND2X1  _1038_
timestamp 1727136778
transform 1 0 1650 0 1 1830
box -12 -8 92 272
use INVX1  _1039_
timestamp 1727136778
transform -1 0 1410 0 -1 1830
box -12 -8 72 272
use AND2X2  _1040_
timestamp 1727136778
transform -1 0 2170 0 1 1830
box -12 -8 112 273
use AND2X2  _1041_
timestamp 1727136778
transform -1 0 2750 0 -1 1830
box -12 -8 112 273
use NAND2X1  _1042_
timestamp 1727136778
transform 1 0 1930 0 1 1830
box -12 -8 92 272
use INVX2  _1043_
timestamp 1727136778
transform 1 0 2330 0 -1 2350
box -12 -8 72 272
use NAND2X1  _1044_
timestamp 1727136778
transform 1 0 2270 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1045_
timestamp 1727136778
transform 1 0 2130 0 -1 1830
box -12 -8 112 272
use NAND3X1  _1046_
timestamp 1727136778
transform -1 0 1730 0 -1 1830
box -12 -8 112 272
use OAI21X1  _1047_
timestamp 1727136778
transform 1 0 1770 0 1 1830
box -12 -8 112 272
use OAI21X1  _1048_
timestamp 1727136778
transform -1 0 2070 0 -1 1830
box -12 -8 112 272
use NAND3X1  _1049_
timestamp 1727136778
transform -1 0 1570 0 -1 1830
box -12 -8 112 272
use AND2X2  _1050_
timestamp 1727136778
transform 1 0 1510 0 -1 1310
box -12 -8 112 273
use OAI21X1  _1051_
timestamp 1727136778
transform -1 0 810 0 -1 790
box -12 -8 112 272
use NAND3X1  _1052_
timestamp 1727136778
transform 1 0 1230 0 -1 1310
box -12 -8 112 272
use NAND3X1  _1053_
timestamp 1727136778
transform 1 0 1230 0 1 1310
box -12 -8 112 272
use NAND2X1  _1054_
timestamp 1727136778
transform -1 0 1470 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1055_
timestamp 1727136778
transform -1 0 1070 0 1 790
box -12 -8 112 272
use NAND3X1  _1056_
timestamp 1727136778
transform 1 0 1030 0 -1 790
box -12 -8 112 272
use OAI21X1  _1057_
timestamp 1727136778
transform -1 0 2010 0 -1 790
box -12 -8 112 272
use NAND3X1  _1058_
timestamp 1727136778
transform 1 0 1290 0 1 790
box -12 -8 112 272
use OAI21X1  _1059_
timestamp 1727136778
transform 1 0 1130 0 1 790
box -12 -8 112 272
use NAND3X1  _1060_
timestamp 1727136778
transform -1 0 1270 0 -1 790
box -12 -8 112 272
use INVX4  _1061_
timestamp 1727136778
transform -1 0 3030 0 1 3910
box -12 -8 92 272
use NOR2X1  _1062_
timestamp 1727136778
transform -1 0 2010 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1063_
timestamp 1727136778
transform 1 0 2190 0 -1 1310
box -12 -8 112 272
use XNOR2X1  _1064_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727153789
transform 1 0 1410 0 1 270
box -12 -8 152 272
use INVX1  _1065_
timestamp 1727136778
transform -1 0 1010 0 -1 270
box -12 -8 72 272
use NAND3X1  _1066_
timestamp 1727136778
transform 1 0 1050 0 -1 270
box -12 -8 112 272
use AOI21X1  _1067_
timestamp 1727136778
transform 1 0 1330 0 -1 790
box -12 -8 112 272
use AOI21X1  _1068_
timestamp 1727136778
transform -1 0 970 0 -1 790
box -12 -8 112 272
use OAI21X1  _1069_
timestamp 1727136778
transform 1 0 1250 0 1 270
box -12 -8 112 272
use NAND3X1  _1070_
timestamp 1727136778
transform 1 0 1990 0 -1 270
box -12 -8 112 272
use NAND2X1  _1071_
timestamp 1727136778
transform 1 0 1610 0 1 270
box -12 -8 92 272
use INVX1  _1072_
timestamp 1727136778
transform -1 0 270 0 -1 270
box -12 -8 72 272
use OAI21X1  _1073_
timestamp 1727136778
transform -1 0 1070 0 1 270
box -12 -8 112 272
use AOI21X1  _1074_
timestamp 1727136778
transform -1 0 910 0 1 790
box -12 -8 112 272
use OAI21X1  _1075_
timestamp 1727136778
transform -1 0 890 0 1 1830
box -12 -8 112 272
use NAND3X1  _1076_
timestamp 1727136778
transform -1 0 1090 0 -1 2350
box -12 -8 112 272
use AOI22X1  _1077_
timestamp 1727136778
transform 1 0 1150 0 -1 2350
box -14 -8 132 272
use INVX1  _1078_
timestamp 1727136778
transform -1 0 550 0 1 2350
box -12 -8 72 272
use NAND2X1  _1079_
timestamp 1727136778
transform -1 0 990 0 1 2350
box -12 -8 92 272
use INVX1  _1080_
timestamp 1727136778
transform -1 0 930 0 -1 2350
box -12 -8 72 272
use NAND3X1  _1081_
timestamp 1727136778
transform -1 0 330 0 -1 2350
box -12 -8 112 272
use NAND2X1  _1082_
timestamp 1727136778
transform -1 0 1110 0 1 2350
box -12 -8 92 272
use NOR2X1  _1083_
timestamp 1727136778
transform -1 0 850 0 1 2350
box -12 -8 92 272
use OAI21X1  _1084_
timestamp 1727136778
transform -1 0 490 0 -1 2350
box -12 -8 112 272
use AOI21X1  _1085_
timestamp 1727136778
transform -1 0 450 0 1 1830
box -12 -8 112 272
use OAI21X1  _1086_
timestamp 1727136778
transform 1 0 710 0 -1 2350
box -12 -8 112 272
use NAND3X1  _1087_
timestamp 1727136778
transform 1 0 550 0 -1 2350
box -12 -8 112 272
use AOI22X1  _1088_
timestamp 1727136778
transform -1 0 750 0 -1 1830
box -14 -8 132 272
use NAND2X1  _1089_
timestamp 1727136778
transform 1 0 1990 0 -1 2870
box -12 -8 92 272
use INVX1  _1090_
timestamp 1727136778
transform 1 0 1590 0 -1 2870
box -12 -8 72 272
use AND2X2  _1091_
timestamp 1727136778
transform -1 0 1990 0 -1 2350
box -12 -8 112 273
use AND2X2  _1092_
timestamp 1727136778
transform -1 0 2150 0 1 2350
box -12 -8 112 273
use NAND2X1  _1093_
timestamp 1727136778
transform 1 0 1910 0 1 2350
box -12 -8 92 272
use AOI22X1  _1094_
timestamp 1727136778
transform 1 0 2190 0 1 3390
box -14 -8 132 272
use INVX1  _1095_
timestamp 1727136778
transform -1 0 1930 0 -1 2870
box -12 -8 72 272
use NAND3X1  _1096_
timestamp 1727136778
transform -1 0 1810 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1097_
timestamp 1727136778
transform -1 0 1690 0 1 2350
box -12 -8 112 272
use OAI21X1  _1098_
timestamp 1727136778
transform -1 0 1850 0 1 2350
box -12 -8 112 272
use NAND3X1  _1099_
timestamp 1727136778
transform -1 0 1550 0 1 2350
box -12 -8 112 272
use AND2X2  _1100_
timestamp 1727136778
transform -1 0 150 0 1 2350
box -12 -8 112 273
use OAI21X1  _1101_
timestamp 1727136778
transform -1 0 170 0 -1 1830
box -12 -8 112 272
use AOI21X1  _1102_
timestamp 1727136778
transform -1 0 1050 0 1 1830
box -12 -8 112 272
use NAND3X1  _1103_
timestamp 1727136778
transform 1 0 650 0 1 1830
box -12 -8 112 272
use NAND3X1  _1104_
timestamp 1727136778
transform 1 0 490 0 1 1830
box -12 -8 112 272
use NAND2X1  _1105_
timestamp 1727136778
transform 1 0 210 0 1 2350
box -12 -8 92 272
use NAND3X1  _1106_
timestamp 1727136778
transform -1 0 170 0 1 1830
box -12 -8 112 272
use NAND3X1  _1107_
timestamp 1727136778
transform 1 0 210 0 1 790
box -12 -8 112 272
use OAI21X1  _1108_
timestamp 1727136778
transform 1 0 910 0 -1 1310
box -12 -8 112 272
use NAND3X1  _1109_
timestamp 1727136778
transform -1 0 470 0 -1 1830
box -12 -8 112 272
use OAI21X1  _1110_
timestamp 1727136778
transform -1 0 310 0 -1 1830
box -12 -8 112 272
use NAND3X1  _1111_
timestamp 1727136778
transform -1 0 170 0 1 1310
box -12 -8 112 272
use NAND2X1  _1112_
timestamp 1727136778
transform -1 0 2130 0 -1 2350
box -12 -8 92 272
use INVX1  _1113_
timestamp 1727136778
transform 1 0 490 0 -1 1310
box -12 -8 72 272
use AOI22X1  _1114_
timestamp 1727136778
transform -1 0 1910 0 -1 1830
box -14 -8 132 272
use INVX1  _1115_
timestamp 1727136778
transform -1 0 590 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1116_
timestamp 1727136778
transform -1 0 730 0 1 1310
box -12 -8 112 272
use NOR2X1  _1117_
timestamp 1727136778
transform 1 0 790 0 1 1310
box -12 -8 92 272
use NAND2X1  _1118_
timestamp 1727136778
transform -1 0 450 0 1 1310
box -12 -8 92 272
use NAND3X1  _1119_
timestamp 1727136778
transform 1 0 510 0 1 790
box -12 -8 112 272
use NAND2X1  _1120_
timestamp 1727136778
transform 1 0 510 0 1 1310
box -12 -8 92 272
use OAI21X1  _1121_
timestamp 1727136778
transform 1 0 930 0 1 1310
box -12 -8 112 272
use NAND3X1  _1122_
timestamp 1727136778
transform -1 0 850 0 -1 1310
box -12 -8 112 272
use NAND2X1  _1123_
timestamp 1727136778
transform -1 0 750 0 1 790
box -12 -8 92 272
use NAND3X1  _1124_
timestamp 1727136778
transform 1 0 550 0 -1 790
box -12 -8 112 272
use AOI21X1  _1125_
timestamp 1727136778
transform 1 0 210 0 1 1310
box -12 -8 112 272
use AOI21X1  _1126_
timestamp 1727136778
transform -1 0 170 0 1 790
box -12 -8 112 272
use NAND3X1  _1127_
timestamp 1727136778
transform 1 0 610 0 -1 1310
box -12 -8 112 272
use NAND3X1  _1128_
timestamp 1727136778
transform -1 0 450 0 -1 1310
box -12 -8 112 272
use NAND2X1  _1129_
timestamp 1727136778
transform -1 0 290 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1130_
timestamp 1727136778
transform 1 0 390 0 -1 790
box -12 -8 112 272
use AOI21X1  _1131_
timestamp 1727136778
transform -1 0 470 0 1 270
box -12 -8 112 272
use AOI21X1  _1132_
timestamp 1727136778
transform -1 0 910 0 1 270
box -12 -8 112 272
use OAI21X1  _1133_
timestamp 1727136778
transform -1 0 170 0 -1 790
box -12 -8 112 272
use NAND3X1  _1134_
timestamp 1727136778
transform -1 0 330 0 -1 790
box -12 -8 112 272
use AOI21X1  _1135_
timestamp 1727136778
transform 1 0 210 0 1 270
box -12 -8 112 272
use OAI21X1  _1136_
timestamp 1727136778
transform -1 0 430 0 -1 270
box -12 -8 112 272
use NAND3X1  _1137_
timestamp 1727136778
transform -1 0 170 0 1 270
box -12 -8 112 272
use NAND3X1  _1138_
timestamp 1727136778
transform 1 0 510 0 1 270
box -12 -8 112 272
use NAND3X1  _1139_
timestamp 1727136778
transform 1 0 630 0 -1 270
box -12 -8 112 272
use AOI21X1  _1140_
timestamp 1727136778
transform 1 0 1830 0 -1 270
box -12 -8 112 272
use INVX1  _1141_
timestamp 1727136778
transform 1 0 2290 0 -1 270
box -12 -8 72 272
use INVX1  _1142_
timestamp 1727136778
transform 1 0 2550 0 1 270
box -12 -8 72 272
use NOR2X1  _1143_
timestamp 1727136778
transform 1 0 3350 0 1 1310
box -12 -8 92 272
use INVX1  _1144_
timestamp 1727136778
transform 1 0 3670 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1145_
timestamp 1727136778
transform 1 0 3050 0 1 1830
box -12 -8 112 272
use AOI21X1  _1146_
timestamp 1727136778
transform -1 0 3470 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1147_
timestamp 1727136778
transform -1 0 3010 0 1 1310
box -12 -8 112 272
use NAND3X1  _1148_
timestamp 1727136778
transform 1 0 3210 0 -1 1310
box -12 -8 112 272
use AOI21X1  _1149_
timestamp 1727136778
transform -1 0 3310 0 1 790
box -12 -8 112 272
use AND2X2  _1150_
timestamp 1727136778
transform 1 0 2850 0 -1 790
box -12 -8 112 273
use NAND3X1  _1151_
timestamp 1727136778
transform 1 0 3350 0 1 790
box -12 -8 112 272
use AOI21X1  _1152_
timestamp 1727136778
transform -1 0 3290 0 -1 790
box -12 -8 112 272
use OAI21X1  _1153_
timestamp 1727136778
transform 1 0 2390 0 -1 790
box -12 -8 112 272
use NAND3X1  _1154_
timestamp 1727136778
transform 1 0 2530 0 -1 790
box -12 -8 112 272
use NAND3X1  _1155_
timestamp 1727136778
transform 1 0 2690 0 -1 790
box -12 -8 112 272
use NAND3X1  _1156_
timestamp 1727136778
transform -1 0 2770 0 1 270
box -12 -8 112 272
use OAI21X1  _1157_
timestamp 1727136778
transform -1 0 1210 0 1 270
box -12 -8 112 272
use NAND3X1  _1158_
timestamp 1727136778
transform 1 0 1210 0 -1 270
box -12 -8 112 272
use AOI22X1  _1159_
timestamp 1727136778
transform -1 0 1870 0 1 270
box -14 -8 132 272
use NAND3X1  _1160_
timestamp 1727136778
transform 1 0 470 0 -1 270
box -12 -8 112 272
use OAI21X1  _1161_
timestamp 1727136778
transform 1 0 790 0 -1 270
box -12 -8 112 272
use AOI21X1  _1162_
timestamp 1727136778
transform 1 0 1370 0 -1 270
box -12 -8 112 272
use NAND3X1  _1163_
timestamp 1727136778
transform 1 0 3330 0 -1 790
box -12 -8 112 272
use NAND3X1  _1164_
timestamp 1727136778
transform 1 0 3790 0 -1 1310
box -12 -8 112 272
use NAND2X1  _1165_
timestamp 1727136778
transform -1 0 4010 0 1 1830
box -12 -8 92 272
use OR2X2  _1166_
timestamp 1727136778
transform 1 0 4170 0 -1 1830
box -12 -8 112 272
use NAND2X1  _1167_
timestamp 1727136778
transform 1 0 4330 0 -1 1830
box -12 -8 92 272
use AOI22X1  _1168_
timestamp 1727136778
transform -1 0 3610 0 1 1830
box -14 -8 132 272
use OAI21X1  _1169_
timestamp 1727136778
transform 1 0 4030 0 -1 1830
box -12 -8 112 272
use OAI21X1  _1170_
timestamp 1727136778
transform 1 0 3530 0 -1 1310
box -12 -8 112 272
use NAND3X1  _1171_
timestamp 1727136778
transform 1 0 4090 0 -1 1310
box -12 -8 112 272
use AOI21X1  _1172_
timestamp 1727136778
transform 1 0 3930 0 -1 1310
box -12 -8 112 272
use OAI21X1  _1173_
timestamp 1727136778
transform 1 0 4090 0 1 790
box -12 -8 112 272
use OAI21X1  _1174_
timestamp 1727136778
transform 1 0 3630 0 -1 790
box -12 -8 112 272
use NAND3X1  _1175_
timestamp 1727136778
transform -1 0 3890 0 -1 790
box -12 -8 112 272
use INVX1  _1176_
timestamp 1727136778
transform 1 0 3670 0 1 270
box -12 -8 72 272
use AOI22X1  _1177_
timestamp 1727136778
transform -1 0 3130 0 -1 790
box -14 -8 132 272
use OAI21X1  _1178_
timestamp 1727136778
transform -1 0 3090 0 1 270
box -12 -8 112 272
use NAND3X1  _1179_
timestamp 1727136778
transform 1 0 3370 0 1 270
box -12 -8 112 272
use AOI21X1  _1180_
timestamp 1727136778
transform 1 0 2150 0 -1 270
box -12 -8 112 272
use NOR3X1  _1181_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 3330 0 -1 270
box -12 -8 192 273
use INVX1  _1182_
timestamp 1727136778
transform -1 0 4030 0 1 790
box -12 -8 72 272
use NAND3X1  _1183_
timestamp 1727136778
transform 1 0 3830 0 1 790
box -12 -8 112 272
use INVX1  _1184_
timestamp 1727136778
transform -1 0 3730 0 1 1830
box -12 -8 72 272
use OAI21X1  _1185_
timestamp 1727136778
transform -1 0 3870 0 1 1830
box -12 -8 112 272
use OR2X2  _1186_
timestamp 1727136778
transform 1 0 4070 0 1 1310
box -12 -8 112 272
use NAND2X1  _1187_
timestamp 1727136778
transform -1 0 3430 0 1 1830
box -12 -8 92 272
use NOR2X1  _1188_
timestamp 1727136778
transform -1 0 4530 0 -1 1830
box -12 -8 92 272
use INVX1  _1189_
timestamp 1727136778
transform 1 0 3790 0 1 1310
box -12 -8 72 272
use OAI21X1  _1190_
timestamp 1727136778
transform 1 0 3910 0 1 1310
box -12 -8 112 272
use NAND3X1  _1191_
timestamp 1727136778
transform -1 0 4310 0 1 1310
box -12 -8 112 272
use INVX1  _1192_
timestamp 1727136778
transform 1 0 4510 0 -1 1310
box -12 -8 72 272
use INVX1  _1193_
timestamp 1727136778
transform 1 0 4390 0 1 790
box -12 -8 72 272
use OAI21X1  _1194_
timestamp 1727136778
transform 1 0 4230 0 1 790
box -12 -8 112 272
use NAND3X1  _1195_
timestamp 1727136778
transform 1 0 4510 0 1 790
box -12 -8 112 272
use AOI21X1  _1196_
timestamp 1727136778
transform 1 0 3950 0 -1 790
box -12 -8 112 272
use NOR3X1  _1197_
timestamp 1727136778
transform -1 0 4290 0 -1 790
box -12 -8 192 273
use OAI21X1  _1198_
timestamp 1727136778
transform 1 0 3130 0 1 270
box -12 -8 112 272
use NAND3X1  _1199_
timestamp 1727136778
transform 1 0 2830 0 1 270
box -12 -8 112 272
use NAND3X1  _1200_
timestamp 1727136778
transform 1 0 3530 0 1 270
box -12 -8 112 272
use NAND3X1  _1201_
timestamp 1727136778
transform -1 0 3870 0 1 270
box -12 -8 112 272
use INVX1  _1202_
timestamp 1727136778
transform 1 0 4090 0 1 270
box -12 -8 72 272
use OAI21X1  _1203_
timestamp 1727136778
transform 1 0 3570 0 -1 270
box -12 -8 112 272
use AOI21X1  _1204_
timestamp 1727136778
transform -1 0 3810 0 -1 270
box -12 -8 112 272
use OAI21X1  _1205_
timestamp 1727136778
transform 1 0 2710 0 -1 270
box -12 -8 112 272
use AOI21X1  _1206_
timestamp 1727136778
transform -1 0 170 0 -1 270
box -12 -8 112 272
use NAND2X1  _1207_
timestamp 1727136778
transform 1 0 790 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1208_
timestamp 1727136778
transform -1 0 170 0 -1 1310
box -12 -8 112 272
use NAND2X1  _1209_
timestamp 1727136778
transform 1 0 2410 0 -1 3390
box -12 -8 92 272
use INVX1  _1210_
timestamp 1727136778
transform -1 0 1610 0 -1 3390
box -12 -8 72 272
use NOR2X1  _1211_
timestamp 1727136778
transform -1 0 2270 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1212_
timestamp 1727136778
transform 1 0 1870 0 1 2870
box -12 -8 112 272
use NAND2X1  _1213_
timestamp 1727136778
transform 1 0 2110 0 -1 3390
box -12 -8 92 272
use OR2X2  _1214_
timestamp 1727136778
transform 1 0 2250 0 -1 3390
box -12 -8 112 272
use NAND3X1  _1215_
timestamp 1727136778
transform -1 0 1510 0 -1 3390
box -12 -8 112 272
use AND2X2  _1216_
timestamp 1727136778
transform -1 0 2070 0 -1 3390
box -12 -8 112 273
use NOR2X1  _1217_
timestamp 1727136778
transform 1 0 2030 0 1 2870
box -12 -8 92 272
use OAI21X1  _1218_
timestamp 1727136778
transform -1 0 1930 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1219_
timestamp 1727136778
transform 1 0 1270 0 -1 3390
box -12 -8 92 272
use AOI21X1  _1220_
timestamp 1727136778
transform -1 0 310 0 1 1830
box -12 -8 112 272
use NAND2X1  _1221_
timestamp 1727136778
transform -1 0 1630 0 -1 3910
box -12 -8 92 272
use AND2X2  _1222_
timestamp 1727136778
transform -1 0 2030 0 -1 4430
box -12 -8 112 273
use OAI21X1  _1223_
timestamp 1727136778
transform 1 0 1810 0 -1 3910
box -12 -8 112 272
use AND2X2  _1224_
timestamp 1727136778
transform -1 0 2230 0 -1 3910
box -12 -8 112 273
use OAI21X1  _1225_
timestamp 1727136778
transform 1 0 1970 0 -1 3910
box -12 -8 112 272
use NAND3X1  _1226_
timestamp 1727136778
transform -1 0 1770 0 -1 3910
box -12 -8 112 272
use INVX1  _1227_
timestamp 1727136778
transform 1 0 1610 0 1 3910
box -12 -8 72 272
use NAND2X1  _1228_
timestamp 1727136778
transform 1 0 2010 0 1 3910
box -12 -8 92 272
use AOI22X1  _1229_
timestamp 1727136778
transform 1 0 2250 0 1 3910
box -14 -8 132 272
use INVX1  _1230_
timestamp 1727136778
transform 1 0 1890 0 1 3910
box -12 -8 72 272
use NAND3X1  _1231_
timestamp 1727136778
transform -1 0 1830 0 1 3910
box -12 -8 112 272
use NAND2X1  _1232_
timestamp 1727136778
transform 1 0 790 0 -1 3910
box -12 -8 92 272
use AOI21X1  _1233_
timestamp 1727136778
transform 1 0 350 0 1 2350
box -12 -8 112 272
use NAND2X1  _1234_
timestamp 1727136778
transform 1 0 1150 0 -1 4430
box -12 -8 92 272
use XOR2X1  _1235_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727152697
transform 1 0 950 0 1 3910
box -12 -8 151 272
use NAND2X1  _1236_
timestamp 1727136778
transform -1 0 390 0 1 3390
box -12 -8 92 272
use OAI21X1  _1237_
timestamp 1727136778
transform 1 0 610 0 1 2350
box -12 -8 112 272
use XNOR2X1  _1238_
timestamp 1727153789
transform 1 0 770 0 1 3910
box -12 -8 152 272
use NAND2X1  _1239_
timestamp 1727136778
transform -1 0 610 0 -1 3910
box -12 -8 92 272
use NAND3X1  _1240_
timestamp 1727136778
transform -1 0 550 0 1 3390
box -12 -8 112 272
use AND2X2  _1241_
timestamp 1727136778
transform -1 0 330 0 -1 3910
box -12 -8 112 273
use NAND2X1  _1242_
timestamp 1727136778
transform 1 0 670 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1243_
timestamp 1727136778
transform 1 0 390 0 -1 3910
box -12 -8 92 272
use NAND3X1  _1244_
timestamp 1727136778
transform 1 0 230 0 1 3910
box -12 -8 112 272
use NAND3X1  _1245_
timestamp 1727136778
transform -1 0 310 0 -1 3390
box -12 -8 112 272
use OAI21X1  _1246_
timestamp 1727136778
transform -1 0 170 0 -1 2350
box -12 -8 112 272
use AOI22X1  _1247_
timestamp 1727136778
transform -1 0 190 0 -1 3910
box -14 -8 132 272
use AOI21X1  _1248_
timestamp 1727136778
transform 1 0 590 0 1 3390
box -12 -8 112 272
use OAI21X1  _1249_
timestamp 1727136778
transform 1 0 70 0 1 2870
box -12 -8 112 272
use NAND3X1  _1250_
timestamp 1727136778
transform -1 0 330 0 1 2870
box -12 -8 112 272
use AND2X2  _1251_
timestamp 1727136778
transform -1 0 1210 0 -1 3390
box -12 -8 112 273
use NAND3X1  _1252_
timestamp 1727136778
transform 1 0 510 0 -1 3390
box -12 -8 112 272
use OAI21X1  _1253_
timestamp 1727136778
transform 1 0 70 0 -1 3390
box -12 -8 112 272
use NAND3X1  _1254_
timestamp 1727136778
transform -1 0 750 0 -1 3390
box -12 -8 112 272
use NAND3X1  _1255_
timestamp 1727136778
transform -1 0 170 0 -1 2870
box -12 -8 112 272
use AOI21X1  _1256_
timestamp 1727136778
transform 1 0 370 0 1 790
box -12 -8 112 272
use AOI22X1  _1257_
timestamp 1727136778
transform -1 0 1070 0 -1 3390
box -14 -8 132 272
use AOI21X1  _1258_
timestamp 1727136778
transform 1 0 390 0 1 2870
box -12 -8 112 272
use OAI21X1  _1259_
timestamp 1727136778
transform -1 0 950 0 1 2870
box -12 -8 112 272
use AOI21X1  _1260_
timestamp 1727136778
transform -1 0 930 0 -1 2870
box -12 -8 112 272
use INVX1  _1261_
timestamp 1727136778
transform 1 0 990 0 -1 2870
box -12 -8 72 272
use NAND3X1  _1262_
timestamp 1727136778
transform 1 0 230 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1263_
timestamp 1727136778
transform -1 0 790 0 1 2870
box -12 -8 112 272
use AOI21X1  _1264_
timestamp 1727136778
transform 1 0 530 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1265_
timestamp 1727136778
transform -1 0 790 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1266_
timestamp 1727136778
transform -1 0 770 0 1 270
box -12 -8 112 272
use NAND3X1  _1267_
timestamp 1727136778
transform -1 0 470 0 -1 2870
box -12 -8 112 272
use NAND3X1  _1268_
timestamp 1727136778
transform 1 0 1110 0 -1 2870
box -12 -8 112 272
use NAND3X1  _1269_
timestamp 1727136778
transform 1 0 1270 0 -1 2870
box -12 -8 112 272
use AND2X2  _1270_
timestamp 1727136778
transform 1 0 2370 0 -1 2870
box -12 -8 112 273
use XOR2X1  _1271_
timestamp 1727152697
transform -1 0 3250 0 -1 2870
box -12 -8 151 272
use NOR2X1  _1272_
timestamp 1727136778
transform 1 0 5030 0 -1 3390
box -12 -8 92 272
use NOR2X1  _1273_
timestamp 1727136778
transform -1 0 4830 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1274_
timestamp 1727136778
transform 1 0 4190 0 -1 2870
box -12 -8 112 272
use AOI21X1  _1275_
timestamp 1727136778
transform 1 0 3990 0 1 2350
box -12 -8 112 272
use OAI21X1  _1276_
timestamp 1727136778
transform -1 0 4570 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1277_
timestamp 1727136778
transform 1 0 4150 0 1 2350
box -12 -8 112 272
use NAND2X1  _1278_
timestamp 1727136778
transform 1 0 4790 0 1 1830
box -12 -8 92 272
use OAI21X1  _1279_
timestamp 1727136778
transform 1 0 4730 0 -1 1830
box -12 -8 112 272
use INVX1  _1280_
timestamp 1727136778
transform -1 0 3630 0 -1 2350
box -12 -8 72 272
use INVX1  _1281_
timestamp 1727136778
transform -1 0 3930 0 1 2350
box -12 -8 72 272
use OAI21X1  _1282_
timestamp 1727136778
transform -1 0 4170 0 -1 2350
box -12 -8 112 272
use OAI21X1  _1283_
timestamp 1727136778
transform -1 0 3810 0 1 2350
box -12 -8 112 272
use NAND3X1  _1284_
timestamp 1727136778
transform -1 0 1770 0 -1 270
box -12 -8 112 272
use INVX1  _1285_
timestamp 1727136778
transform -1 0 3330 0 1 270
box -12 -8 72 272
use NAND2X1  _1286_
timestamp 1727136778
transform -1 0 1610 0 -1 270
box -12 -8 92 272
use NAND3X1  _1287_
timestamp 1727136778
transform 1 0 1930 0 1 270
box -12 -8 112 272
use NAND3X1  _1288_
timestamp 1727136778
transform 1 0 3010 0 -1 270
box -12 -8 112 272
use AOI21X1  _1289_
timestamp 1727136778
transform 1 0 2870 0 -1 270
box -12 -8 112 272
use OAI21X1  _1290_
timestamp 1727136778
transform -1 0 3270 0 -1 270
box -12 -8 112 272
use AOI21X1  _1291_
timestamp 1727136778
transform -1 0 2510 0 -1 270
box -12 -8 112 272
use NAND2X1  _1292_
timestamp 1727136778
transform -1 0 2330 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1293_
timestamp 1727136778
transform -1 0 2750 0 -1 2870
box -12 -8 112 272
use INVX1  _1294_
timestamp 1727136778
transform 1 0 1290 0 1 2870
box -12 -8 72 272
use AOI21X1  _1295_
timestamp 1727136778
transform 1 0 1130 0 1 2870
box -12 -8 112 272
use OAI21X1  _1296_
timestamp 1727136778
transform -1 0 1770 0 -1 3390
box -12 -8 112 272
use INVX1  _1297_
timestamp 1727136778
transform 1 0 1650 0 1 3390
box -12 -8 72 272
use AOI21X1  _1298_
timestamp 1727136778
transform 1 0 350 0 -1 3390
box -12 -8 112 272
use OAI21X1  _1299_
timestamp 1727136778
transform 1 0 810 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1300_
timestamp 1727136778
transform -1 0 1710 0 -1 4430
box -12 -8 92 272
use NOR2X1  _1301_
timestamp 1727136778
transform 1 0 2070 0 1 3390
box -12 -8 92 272
use NAND2X1  _1302_
timestamp 1727136778
transform -1 0 2010 0 1 4430
box -12 -8 92 272
use NAND2X1  _1303_
timestamp 1727136778
transform -1 0 2170 0 -1 4430
box -12 -8 92 272
use OAI22X1  _1304_
timestamp 1727136778
transform -1 0 1870 0 -1 4430
box -12 -8 132 272
use XNOR2X1  _1305_
timestamp 1727153789
transform -1 0 1570 0 -1 4430
box -12 -8 152 272
use XNOR2X1  _1306_
timestamp 1727153789
transform 1 0 810 0 -1 4430
box -12 -8 152 272
use NOR2X1  _1307_
timestamp 1727136778
transform 1 0 370 0 1 3910
box -12 -8 92 272
use AOI21X1  _1308_
timestamp 1727136778
transform -1 0 170 0 1 3910
box -12 -8 112 272
use NAND2X1  _1309_
timestamp 1727136778
transform 1 0 1350 0 1 4430
box -12 -8 92 272
use NAND2X1  _1310_
timestamp 1727136778
transform 1 0 1630 0 -1 4950
box -12 -8 92 272
use INVX1  _1311_
timestamp 1727136778
transform 1 0 1130 0 -1 4950
box -12 -8 72 272
use AND2X2  _1312_
timestamp 1727136778
transform -1 0 1870 0 -1 4950
box -12 -8 112 273
use AND2X2  _1313_
timestamp 1727136778
transform -1 0 1470 0 -1 4950
box -12 -8 112 273
use NAND2X1  _1314_
timestamp 1727136778
transform -1 0 1310 0 -1 4950
box -12 -8 92 272
use AOI22X1  _1315_
timestamp 1727136778
transform 1 0 1330 0 1 4950
box -14 -8 132 272
use INVX1  _1316_
timestamp 1727136778
transform -1 0 850 0 1 4950
box -12 -8 72 272
use AOI21X1  _1317_
timestamp 1727136778
transform 1 0 970 0 -1 4950
box -12 -8 112 272
use INVX2  _1318_
timestamp 1727136778
transform 1 0 2810 0 1 4430
box -12 -8 72 272
use OAI21X1  _1319_
timestamp 1727136778
transform -1 0 2170 0 1 4430
box -12 -8 112 272
use OAI21X1  _1320_
timestamp 1727136778
transform -1 0 1870 0 1 4430
box -12 -8 112 272
use AOI21X1  _1321_
timestamp 1727136778
transform -1 0 1730 0 1 4430
box -12 -8 112 272
use OAI22X1  _1322_
timestamp 1727136778
transform -1 0 1290 0 1 4430
box -12 -8 132 272
use NAND3X1  _1323_
timestamp 1727136778
transform -1 0 1570 0 1 4430
box -12 -8 112 272
use NAND3X1  _1324_
timestamp 1727136778
transform -1 0 930 0 -1 4950
box -12 -8 112 272
use NOR2X1  _1325_
timestamp 1727136778
transform -1 0 1110 0 1 4430
box -12 -8 92 272
use NAND3X1  _1326_
timestamp 1727136778
transform -1 0 770 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1327_
timestamp 1727136778
transform -1 0 150 0 -1 4950
box -12 -8 92 272
use NOR2X1  _1328_
timestamp 1727136778
transform -1 0 150 0 -1 4430
box -12 -8 92 272
use NOR2X1  _1329_
timestamp 1727136778
transform 1 0 650 0 1 3910
box -12 -8 92 272
use OAI21X1  _1330_
timestamp 1727136778
transform -1 0 610 0 1 3910
box -12 -8 112 272
use AOI21X1  _1331_
timestamp 1727136778
transform 1 0 210 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1332_
timestamp 1727136778
transform 1 0 490 0 -1 4430
box -12 -8 112 272
use XOR2X1  _1333_
timestamp 1727152697
transform 1 0 830 0 1 4430
box -12 -8 151 272
use NAND3X1  _1334_
timestamp 1727136778
transform 1 0 530 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1335_
timestamp 1727136778
transform -1 0 130 0 1 4430
box -12 -8 92 272
use NAND3X1  _1336_
timestamp 1727136778
transform 1 0 510 0 1 4430
box -12 -8 112 272
use NAND3X1  _1337_
timestamp 1727136778
transform 1 0 1150 0 1 3910
box -12 -8 112 272
use NOR3X1  _1338_
timestamp 1727136778
transform 1 0 70 0 1 3390
box -12 -8 192 273
use AOI21X1  _1339_
timestamp 1727136778
transform 1 0 730 0 1 3390
box -12 -8 112 272
use AOI21X1  _1340_
timestamp 1727136778
transform 1 0 670 0 1 4430
box -12 -8 112 272
use NAND3X1  _1341_
timestamp 1727136778
transform 1 0 190 0 1 4430
box -12 -8 112 272
use OAI21X1  _1342_
timestamp 1727136778
transform -1 0 290 0 -1 4430
box -12 -8 112 272
use AOI21X1  _1343_
timestamp 1727136778
transform 1 0 350 0 -1 4430
box -12 -8 112 272
use OAI21X1  _1344_
timestamp 1727136778
transform -1 0 990 0 1 3390
box -12 -8 112 272
use NAND3X1  _1345_
timestamp 1727136778
transform -1 0 1590 0 1 3390
box -12 -8 112 272
use NAND3X1  _1346_
timestamp 1727136778
transform 1 0 930 0 -1 3910
box -12 -8 112 272
use OAI21X1  _1347_
timestamp 1727136778
transform 1 0 1050 0 1 3390
box -12 -8 112 272
use NAND3X1  _1348_
timestamp 1727136778
transform -1 0 1450 0 1 3390
box -12 -8 112 272
use NAND3X1  _1349_
timestamp 1727136778
transform -1 0 1510 0 1 2870
box -12 -8 112 272
use AOI21X1  _1350_
timestamp 1727136778
transform 1 0 550 0 1 2870
box -12 -8 112 272
use OAI21X1  _1351_
timestamp 1727136778
transform 1 0 990 0 1 2870
box -12 -8 112 272
use NAND3X1  _1352_
timestamp 1727136778
transform 1 0 1770 0 1 3390
box -12 -8 112 272
use NAND3X1  _1353_
timestamp 1727136778
transform -1 0 1310 0 1 3390
box -12 -8 112 272
use NAND3X1  _1354_
timestamp 1727136778
transform 1 0 1710 0 1 2870
box -12 -8 112 272
use NAND2X1  _1355_
timestamp 1727136778
transform -1 0 2250 0 1 2870
box -12 -8 92 272
use AND2X2  _1356_
timestamp 1727136778
transform 1 0 3310 0 -1 2870
box -12 -8 112 273
use OAI21X1  _1357_
timestamp 1727136778
transform 1 0 3450 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1358_
timestamp 1727136778
transform 1 0 3610 0 -1 2870
box -12 -8 112 272
use AND2X2  _1359_
timestamp 1727136778
transform 1 0 4590 0 -1 1830
box -12 -8 112 273
use NAND2X1  _1360_
timestamp 1727136778
transform 1 0 4530 0 1 1830
box -12 -8 92 272
use OAI21X1  _1361_
timestamp 1727136778
transform -1 0 4310 0 1 1830
box -12 -8 112 272
use OAI21X1  _1362_
timestamp 1727136778
transform 1 0 4370 0 1 1830
box -12 -8 112 272
use AOI21X1  _1363_
timestamp 1727136778
transform -1 0 4170 0 1 1830
box -12 -8 112 272
use AOI22X1  _1364_
timestamp 1727136778
transform 1 0 3910 0 -1 2350
box -14 -8 132 272
use OAI21X1  _1365_
timestamp 1727136778
transform -1 0 4930 0 1 1310
box -12 -8 112 272
use AOI21X1  _1366_
timestamp 1727136778
transform -1 0 1670 0 1 2870
box -12 -8 112 272
use AOI22X1  _1367_
timestamp 1727136778
transform 1 0 1410 0 -1 2870
box -14 -8 132 272
use NOR2X1  _1368_
timestamp 1727136778
transform 1 0 2130 0 -1 2870
box -12 -8 92 272
use NAND3X1  _1369_
timestamp 1727136778
transform 1 0 2950 0 -1 2870
box -12 -8 112 272
use AOI21X1  _1370_
timestamp 1727136778
transform 1 0 2290 0 1 2870
box -12 -8 112 272
use INVX1  _1371_
timestamp 1727136778
transform 1 0 2530 0 -1 2870
box -12 -8 72 272
use NAND2X1  _1372_
timestamp 1727136778
transform -1 0 1370 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1373_
timestamp 1727136778
transform 1 0 990 0 -1 4430
box -12 -8 112 272
use INVX1  _1374_
timestamp 1727136778
transform -1 0 590 0 1 4950
box -12 -8 72 272
use AOI21X1  _1375_
timestamp 1727136778
transform -1 0 450 0 1 4430
box -12 -8 112 272
use NAND2X1  _1376_
timestamp 1727136778
transform -1 0 1370 0 1 5470
box -12 -8 92 272
use INVX1  _1377_
timestamp 1727136778
transform -1 0 950 0 1 5470
box -12 -8 72 272
use NOR2X1  _1378_
timestamp 1727136778
transform -1 0 1270 0 1 4950
box -12 -8 92 272
use OAI21X1  _1379_
timestamp 1727136778
transform -1 0 1130 0 1 4950
box -12 -8 112 272
use NAND2X1  _1380_
timestamp 1727136778
transform -1 0 1250 0 1 5470
box -12 -8 92 272
use OR2X2  _1381_
timestamp 1727136778
transform -1 0 1110 0 1 5470
box -12 -8 112 272
use NAND3X1  _1382_
timestamp 1727136778
transform -1 0 830 0 1 5470
box -12 -8 112 272
use AND2X2  _1383_
timestamp 1727136778
transform -1 0 1110 0 -1 5990
box -12 -8 112 273
use NOR2X1  _1384_
timestamp 1727136778
transform -1 0 1250 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1385_
timestamp 1727136778
transform -1 0 950 0 -1 5990
box -12 -8 112 272
use NAND2X1  _1386_
timestamp 1727136778
transform -1 0 310 0 -1 5990
box -12 -8 92 272
use OR2X2  _1387_
timestamp 1727136778
transform 1 0 650 0 -1 4430
box -12 -8 112 272
use NAND2X1  _1388_
timestamp 1727136778
transform 1 0 1610 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1389_
timestamp 1727136778
transform -1 0 1890 0 1 4950
box -12 -8 92 272
use NAND2X1  _1390_
timestamp 1727136778
transform -1 0 1770 0 1 4950
box -12 -8 92 272
use AOI22X1  _1391_
timestamp 1727136778
transform -1 0 1630 0 1 4950
box -14 -8 132 272
use INVX1  _1392_
timestamp 1727136778
transform 1 0 2050 0 -1 5470
box -12 -8 72 272
use OAI21X1  _1393_
timestamp 1727136778
transform 1 0 1910 0 -1 5470
box -12 -8 112 272
use XNOR2X1  _1394_
timestamp 1727153789
transform 1 0 1410 0 -1 5470
box -12 -8 152 272
use AOI21X1  _1395_
timestamp 1727136778
transform 1 0 430 0 1 5470
box -12 -8 112 272
use NAND3X1  _1396_
timestamp 1727136778
transform -1 0 690 0 1 5470
box -12 -8 112 272
use INVX1  _1397_
timestamp 1727136778
transform -1 0 130 0 1 5990
box -12 -8 72 272
use OAI21X1  _1398_
timestamp 1727136778
transform -1 0 430 0 1 5990
box -12 -8 112 272
use AND2X2  _1399_
timestamp 1727136778
transform -1 0 790 0 -1 5990
box -12 -8 112 273
use NAND2X1  _1400_
timestamp 1727136778
transform -1 0 390 0 1 5470
box -12 -8 92 272
use INVX1  _1401_
timestamp 1727136778
transform -1 0 110 0 1 5470
box -12 -8 72 272
use NAND2X1  _1402_
timestamp 1727136778
transform -1 0 250 0 1 5470
box -12 -8 92 272
use NAND3X1  _1403_
timestamp 1727136778
transform 1 0 370 0 -1 5990
box -12 -8 112 272
use NAND3X1  _1404_
timestamp 1727136778
transform -1 0 590 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1405_
timestamp 1727136778
transform 1 0 370 0 -1 4950
box -12 -8 112 272
use AOI22X1  _1406_
timestamp 1727136778
transform -1 0 190 0 -1 5990
box -14 -8 132 272
use OR2X2  _1407_
timestamp 1727136778
transform -1 0 170 0 -1 5470
box -12 -8 112 272
use NAND2X1  _1408_
timestamp 1727136778
transform -1 0 450 0 -1 5470
box -12 -8 92 272
use AOI21X1  _1409_
timestamp 1727136778
transform -1 0 330 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1410_
timestamp 1727136778
transform 1 0 230 0 1 4950
box -12 -8 112 272
use NAND3X1  _1411_
timestamp 1727136778
transform -1 0 470 0 1 4950
box -12 -8 112 272
use NAND3X1  _1412_
timestamp 1727136778
transform 1 0 650 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1413_
timestamp 1727136778
transform -1 0 170 0 1 4950
box -12 -8 112 272
use NAND3X1  _1414_
timestamp 1727136778
transform -1 0 730 0 1 4950
box -12 -8 112 272
use NAND2X1  _1415_
timestamp 1727136778
transform -1 0 1390 0 1 3910
box -12 -8 92 272
use NAND3X1  _1416_
timestamp 1727136778
transform 1 0 1930 0 1 3390
box -12 -8 112 272
use AOI21X1  _1417_
timestamp 1727136778
transform 1 0 1070 0 -1 3910
box -12 -8 112 272
use OAI21X1  _1418_
timestamp 1727136778
transform -1 0 1330 0 -1 3910
box -12 -8 112 272
use NAND3X1  _1419_
timestamp 1727136778
transform 1 0 1390 0 -1 3910
box -12 -8 112 272
use NAND2X1  _1420_
timestamp 1727136778
transform -1 0 2550 0 1 3390
box -12 -8 92 272
use AOI21X1  _1421_
timestamp 1727136778
transform -1 0 2570 0 1 2350
box -12 -8 112 272
use NAND2X1  _1422_
timestamp 1727136778
transform 1 0 2810 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1423_
timestamp 1727136778
transform -1 0 2710 0 1 2350
box -12 -8 112 272
use INVX1  _1424_
timestamp 1727136778
transform 1 0 2890 0 -1 2350
box -12 -8 72 272
use NOR2X1  _1425_
timestamp 1727136778
transform -1 0 3090 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1426_
timestamp 1727136778
transform 1 0 3130 0 -1 2350
box -12 -8 112 272
use NOR2X1  _1427_
timestamp 1727136778
transform 1 0 4630 0 -1 2870
box -12 -8 92 272
use NOR2X1  _1428_
timestamp 1727136778
transform -1 0 4390 0 1 2350
box -12 -8 92 272
use AOI21X1  _1429_
timestamp 1727136778
transform 1 0 4370 0 1 1310
box -12 -8 112 272
use OAI21X1  _1430_
timestamp 1727136778
transform 1 0 4510 0 1 1310
box -12 -8 112 272
use NOR2X1  _1431_
timestamp 1727136778
transform -1 0 4810 0 1 2350
box -12 -8 92 272
use NOR2X1  _1432_
timestamp 1727136778
transform 1 0 4770 0 -1 2350
box -12 -8 92 272
use AOI22X1  _1433_
timestamp 1727136778
transform -1 0 4470 0 -1 2350
box -14 -8 132 272
use OAI21X1  _1434_
timestamp 1727136778
transform 1 0 4670 0 1 1310
box -12 -8 112 272
use INVX1  _1435_
timestamp 1727136778
transform 1 0 5970 0 -1 790
box -12 -8 72 272
use INVX1  _1436_
timestamp 1727136778
transform -1 0 5830 0 1 2870
box -12 -8 72 272
use OAI21X1  _1437_
timestamp 1727136778
transform -1 0 3990 0 -1 2870
box -12 -8 112 272
use INVX1  _1438_
timestamp 1727136778
transform 1 0 2690 0 -1 3390
box -12 -8 72 272
use OAI21X1  _1439_
timestamp 1727136778
transform 1 0 1290 0 -1 5990
box -12 -8 112 272
use INVX1  _1440_
timestamp 1727136778
transform -1 0 1270 0 1 5990
box -12 -8 72 272
use AOI21X1  _1441_
timestamp 1727136778
transform 1 0 530 0 -1 5990
box -12 -8 112 272
use NAND2X1  _1442_
timestamp 1727136778
transform 1 0 1830 0 1 5470
box -12 -8 92 272
use INVX1  _1443_
timestamp 1727136778
transform -1 0 2150 0 -1 5990
box -12 -8 72 272
use NOR2X1  _1444_
timestamp 1727136778
transform -1 0 1510 0 1 5470
box -12 -8 92 272
use OAI22X1  _1445_
timestamp 1727136778
transform -1 0 1850 0 -1 5470
box -12 -8 132 272
use NAND2X1  _1446_
timestamp 1727136778
transform 1 0 1570 0 1 5470
box -12 -8 92 272
use NOR2X1  _1447_
timestamp 1727136778
transform 1 0 1710 0 1 5470
box -12 -8 92 272
use INVX1  _1448_
timestamp 1727136778
transform 1 0 1810 0 -1 5990
box -12 -8 72 272
use NAND3X1  _1449_
timestamp 1727136778
transform -1 0 2030 0 -1 5990
box -12 -8 112 272
use INVX1  _1450_
timestamp 1727136778
transform -1 0 1630 0 -1 5990
box -12 -8 72 272
use OAI21X1  _1451_
timestamp 1727136778
transform 1 0 1670 0 -1 5990
box -12 -8 112 272
use NAND2X1  _1452_
timestamp 1727136778
transform 1 0 1930 0 -1 4950
box -12 -8 92 272
use NAND2X1  _1453_
timestamp 1727136778
transform 1 0 2110 0 1 4950
box -12 -8 92 272
use OR2X2  _1454_
timestamp 1727136778
transform 1 0 1950 0 1 4950
box -12 -8 112 272
use INVX1  _1455_
timestamp 1727136778
transform 1 0 2890 0 -1 5470
box -12 -8 72 272
use OAI21X1  _1456_
timestamp 1727136778
transform -1 0 2270 0 -1 5470
box -12 -8 112 272
use AND2X2  _1457_
timestamp 1727136778
transform -1 0 2070 0 1 5470
box -12 -8 112 273
use AOI21X1  _1458_
timestamp 1727136778
transform -1 0 1710 0 1 5990
box -12 -8 112 272
use INVX1  _1459_
timestamp 1727136778
transform -1 0 550 0 1 5990
box -12 -8 72 272
use NAND3X1  _1460_
timestamp 1727136778
transform 1 0 1770 0 1 5990
box -12 -8 112 272
use NAND3X1  _1461_
timestamp 1727136778
transform 1 0 750 0 1 5990
box -12 -8 112 272
use OAI21X1  _1462_
timestamp 1727136778
transform -1 0 290 0 1 5990
box -12 -8 112 272
use INVX1  _1463_
timestamp 1727136778
transform -1 0 1510 0 -1 5990
box -12 -8 72 272
use OAI21X1  _1464_
timestamp 1727136778
transform -1 0 990 0 1 5990
box -12 -8 112 272
use NAND3X1  _1465_
timestamp 1727136778
transform -1 0 1150 0 1 5990
box -12 -8 112 272
use NAND3X1  _1466_
timestamp 1727136778
transform -1 0 710 0 1 5990
box -12 -8 112 272
use OAI21X1  _1467_
timestamp 1727136778
transform -1 0 1410 0 1 5990
box -12 -8 112 272
use NAND3X1  _1468_
timestamp 1727136778
transform 1 0 1470 0 1 5990
box -12 -8 112 272
use NAND2X1  _1469_
timestamp 1727136778
transform -1 0 1210 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1470_
timestamp 1727136778
transform -1 0 990 0 1 4950
box -12 -8 112 272
use AOI21X1  _1471_
timestamp 1727136778
transform 1 0 810 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1472_
timestamp 1727136778
transform 1 0 970 0 -1 5470
box -12 -8 112 272
use NAND3X1  _1473_
timestamp 1727136778
transform 1 0 1250 0 -1 5470
box -12 -8 112 272
use NAND2X1  _1474_
timestamp 1727136778
transform 1 0 2810 0 -1 3390
box -12 -8 92 272
use NOR3X1  _1475_
timestamp 1727136778
transform 1 0 2770 0 1 2350
box -12 -8 192 273
use AOI21X1  _1476_
timestamp 1727136778
transform 1 0 3010 0 1 2350
box -12 -8 112 272
use INVX1  _1477_
timestamp 1727136778
transform 1 0 3150 0 1 2350
box -12 -8 72 272
use OAI21X1  _1478_
timestamp 1727136778
transform 1 0 3270 0 1 2350
box -12 -8 112 272
use OAI21X1  _1479_
timestamp 1727136778
transform 1 0 3550 0 1 2350
box -12 -8 112 272
use NAND2X1  _1480_
timestamp 1727136778
transform -1 0 4310 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1481_
timestamp 1727136778
transform -1 0 4450 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1482_
timestamp 1727136778
transform 1 0 4670 0 1 790
box -12 -8 92 272
use NAND2X1  _1483_
timestamp 1727136778
transform 1 0 5390 0 1 790
box -12 -8 92 272
use OAI21X1  _1484_
timestamp 1727136778
transform -1 0 5630 0 1 790
box -12 -8 112 272
use AOI21X1  _1485_
timestamp 1727136778
transform 1 0 5530 0 -1 790
box -12 -8 112 272
use AOI22X1  _1486_
timestamp 1727136778
transform -1 0 5790 0 -1 790
box -14 -8 132 272
use INVX1  _1487_
timestamp 1727136778
transform 1 0 5850 0 -1 790
box -12 -8 72 272
use OAI21X1  _1488_
timestamp 1727136778
transform 1 0 2210 0 -1 5990
box -12 -8 112 272
use INVX1  _1489_
timestamp 1727136778
transform 1 0 2350 0 -1 5990
box -12 -8 72 272
use INVX1  _1490_
timestamp 1727136778
transform -1 0 2430 0 1 4950
box -12 -8 72 272
use NAND2X1  _1491_
timestamp 1727136778
transform -1 0 2970 0 1 5470
box -12 -8 92 272
use OAI21X1  _1492_
timestamp 1727136778
transform -1 0 2210 0 1 5470
box -12 -8 112 272
use OAI21X1  _1493_
timestamp 1727136778
transform -1 0 2370 0 1 5470
box -12 -8 112 272
use OR2X2  _1494_
timestamp 1727136778
transform 1 0 2590 0 1 5470
box -12 -8 112 272
use INVX1  _1495_
timestamp 1727136778
transform 1 0 2990 0 -1 5470
box -12 -8 72 272
use OAI21X1  _1496_
timestamp 1727136778
transform 1 0 2430 0 1 5470
box -12 -8 112 272
use NAND2X1  _1497_
timestamp 1727136778
transform 1 0 2630 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1498_
timestamp 1727136778
transform 1 0 2750 0 -1 5470
box -12 -8 112 272
use INVX1  _1499_
timestamp 1727136778
transform 1 0 2250 0 1 4950
box -12 -8 72 272
use NAND3X1  _1500_
timestamp 1727136778
transform 1 0 2470 0 -1 5470
box -12 -8 112 272
use NAND2X1  _1501_
timestamp 1727136778
transform 1 0 2750 0 1 5470
box -12 -8 92 272
use NOR2X1  _1502_
timestamp 1727136778
transform 1 0 2750 0 -1 5990
box -12 -8 92 272
use NAND2X1  _1503_
timestamp 1727136778
transform 1 0 2810 0 1 5990
box -12 -8 92 272
use INVX1  _1504_
timestamp 1727136778
transform 1 0 2890 0 -1 5990
box -12 -8 72 272
use OAI21X1  _1505_
timestamp 1727136778
transform -1 0 2550 0 -1 5990
box -12 -8 112 272
use OR2X2  _1506_
timestamp 1727136778
transform -1 0 2750 0 1 5990
box -12 -8 112 272
use NAND3X1  _1507_
timestamp 1727136778
transform -1 0 2590 0 1 5990
box -12 -8 112 272
use NAND2X1  _1508_
timestamp 1727136778
transform -1 0 2290 0 1 5990
box -12 -8 92 272
use NAND3X1  _1509_
timestamp 1727136778
transform 1 0 2070 0 1 5990
box -12 -8 112 272
use NAND2X1  _1510_
timestamp 1727136778
transform -1 0 2010 0 1 5990
box -12 -8 92 272
use NAND3X1  _1511_
timestamp 1727136778
transform 1 0 2330 0 1 5990
box -12 -8 112 272
use NAND2X1  _1512_
timestamp 1727136778
transform -1 0 2810 0 1 3390
box -12 -8 92 272
use NOR2X1  _1513_
timestamp 1727136778
transform 1 0 3350 0 1 2870
box -12 -8 92 272
use NOR2X1  _1514_
timestamp 1727136778
transform -1 0 3130 0 1 2870
box -12 -8 92 272
use NAND3X1  _1515_
timestamp 1727136778
transform 1 0 3190 0 1 2870
box -12 -8 112 272
use NAND2X1  _1516_
timestamp 1727136778
transform -1 0 2630 0 -1 3390
box -12 -8 92 272
use AOI22X1  _1517_
timestamp 1727136778
transform 1 0 2890 0 1 2870
box -14 -8 132 272
use AOI21X1  _1518_
timestamp 1727136778
transform -1 0 3330 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1519_
timestamp 1727136778
transform 1 0 2950 0 -1 3390
box -12 -8 92 272
use OAI21X1  _1520_
timestamp 1727136778
transform 1 0 3070 0 -1 3390
box -12 -8 112 272
use AOI21X1  _1521_
timestamp 1727136778
transform 1 0 2590 0 1 2870
box -12 -8 112 272
use OAI21X1  _1522_
timestamp 1727136778
transform 1 0 2750 0 1 2870
box -12 -8 112 272
use AOI22X1  _1523_
timestamp 1727136778
transform 1 0 2870 0 1 3390
box -14 -8 132 272
use OAI21X1  _1524_
timestamp 1727136778
transform 1 0 3310 0 1 3390
box -12 -8 112 272
use OR2X2  _1525_
timestamp 1727136778
transform -1 0 5590 0 1 2870
box -12 -8 112 272
use NAND3X1  _1526_
timestamp 1727136778
transform -1 0 5090 0 1 2350
box -12 -8 112 272
use INVX1  _1527_
timestamp 1727136778
transform 1 0 4490 0 -1 790
box -12 -8 72 272
use OAI21X1  _1528_
timestamp 1727136778
transform 1 0 4350 0 -1 790
box -12 -8 112 272
use NAND2X1  _1529_
timestamp 1727136778
transform 1 0 4610 0 -1 790
box -12 -8 92 272
use NAND2X1  _1530_
timestamp 1727136778
transform -1 0 4930 0 1 2350
box -12 -8 92 272
use OAI21X1  _1531_
timestamp 1727136778
transform -1 0 5190 0 1 790
box -12 -8 112 272
use AOI21X1  _1532_
timestamp 1727136778
transform 1 0 5250 0 1 790
box -12 -8 112 272
use AOI22X1  _1533_
timestamp 1727136778
transform -1 0 5470 0 -1 790
box -14 -8 132 272
use INVX1  _1534_
timestamp 1727136778
transform -1 0 5230 0 1 270
box -12 -8 72 272
use INVX1  _1535_
timestamp 1727136778
transform -1 0 3830 0 -1 2870
box -12 -8 72 272
use NAND2X1  _1536_
timestamp 1727136778
transform 1 0 3190 0 1 3390
box -12 -8 92 272
use INVX1  _1537_
timestamp 1727136778
transform 1 0 2830 0 1 3910
box -12 -8 72 272
use AOI21X1  _1538_
timestamp 1727136778
transform 1 0 2610 0 -1 5990
box -12 -8 112 272
use OAI21X1  _1539_
timestamp 1727136778
transform 1 0 2310 0 -1 5470
box -12 -8 112 272
use NOR2X1  _1540_
timestamp 1727136778
transform -1 0 2730 0 1 4950
box -12 -8 92 272
use NAND3X1  _1541_
timestamp 1727136778
transform -1 0 2910 0 -1 4950
box -12 -8 112 272
use OAI22X1  _1542_
timestamp 1727136778
transform -1 0 2590 0 1 4950
box -12 -8 132 272
use NAND2X1  _1543_
timestamp 1727136778
transform 1 0 2670 0 -1 4950
box -12 -8 92 272
use XNOR2X1  _1544_
timestamp 1727153789
transform 1 0 2470 0 -1 4950
box -12 -8 152 272
use XOR2X1  _1545_
timestamp 1727152697
transform -1 0 2610 0 1 4430
box -12 -8 151 272
use XOR2X1  _1546_
timestamp 1727152697
transform -1 0 2650 0 -1 4430
box -12 -8 151 272
use NOR2X1  _1547_
timestamp 1727136778
transform -1 0 2770 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1548_
timestamp 1727136778
transform -1 0 3150 0 1 3390
box -12 -8 112 272
use OAI21X1  _1549_
timestamp 1727136778
transform -1 0 2910 0 -1 3910
box -12 -8 112 272
use NAND3X1  _1550_
timestamp 1727136778
transform 1 0 3490 0 1 2870
box -12 -8 112 272
use AOI21X1  _1551_
timestamp 1727136778
transform 1 0 3930 0 1 270
box -12 -8 112 272
use OAI21X1  _1552_
timestamp 1727136778
transform 1 0 4190 0 1 270
box -12 -8 112 272
use INVX1  _1553_
timestamp 1727136778
transform -1 0 5130 0 1 1830
box -12 -8 72 272
use AOI21X1  _1554_
timestamp 1727136778
transform 1 0 5250 0 -1 1310
box -12 -8 112 272
use AOI21X1  _1555_
timestamp 1727136778
transform 1 0 5210 0 -1 790
box -12 -8 112 272
use AOI22X1  _1556_
timestamp 1727136778
transform -1 0 5110 0 1 270
box -14 -8 132 272
use INVX1  _1557_
timestamp 1727136778
transform -1 0 4930 0 1 270
box -12 -8 72 272
use NAND3X1  _1558_
timestamp 1727136778
transform 1 0 2530 0 -1 3910
box -12 -8 112 272
use INVX1  _1559_
timestamp 1727136778
transform 1 0 3550 0 -1 3390
box -12 -8 72 272
use NAND3X1  _1560_
timestamp 1727136778
transform 1 0 3670 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1561_
timestamp 1727136778
transform -1 0 2770 0 1 3910
box -12 -8 92 272
use OAI21X1  _1562_
timestamp 1727136778
transform 1 0 2710 0 -1 4430
box -12 -8 112 272
use INVX1  _1563_
timestamp 1727136778
transform 1 0 3730 0 1 3390
box -12 -8 72 272
use INVX1  _1564_
timestamp 1727136778
transform -1 0 2110 0 -1 4950
box -12 -8 72 272
use NAND2X1  _1565_
timestamp 1727136778
transform -1 0 2250 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1566_
timestamp 1727136778
transform -1 0 2410 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1567_
timestamp 1727136778
transform 1 0 2910 0 1 4430
box -12 -8 112 272
use XOR2X1  _1568_
timestamp 1727152697
transform 1 0 3350 0 1 4430
box -12 -8 151 272
use NAND3X1  _1569_
timestamp 1727136778
transform 1 0 3970 0 -1 3390
box -12 -8 112 272
use AOI21X1  _1570_
timestamp 1727136778
transform 1 0 3390 0 -1 3390
box -12 -8 112 272
use INVX1  _1571_
timestamp 1727136778
transform -1 0 3670 0 1 3390
box -12 -8 72 272
use OAI21X1  _1572_
timestamp 1727136778
transform 1 0 3470 0 1 3390
box -12 -8 112 272
use NAND3X1  _1573_
timestamp 1727136778
transform 1 0 4130 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1574_
timestamp 1727136778
transform -1 0 4130 0 -1 270
box -12 -8 92 272
use NOR2X1  _1575_
timestamp 1727136778
transform 1 0 4350 0 -1 270
box -12 -8 92 272
use AOI21X1  _1576_
timestamp 1727136778
transform 1 0 4190 0 -1 270
box -12 -8 112 272
use OAI21X1  _1577_
timestamp 1727136778
transform 1 0 4470 0 -1 270
box -12 -8 112 272
use NOR2X1  _1578_
timestamp 1727136778
transform 1 0 5730 0 -1 3390
box -12 -8 92 272
use NOR2X1  _1579_
timestamp 1727136778
transform -1 0 5210 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1580_
timestamp 1727136778
transform -1 0 5170 0 -1 790
box -12 -8 112 272
use AOI22X1  _1581_
timestamp 1727136778
transform 1 0 4910 0 -1 790
box -14 -8 132 272
use INVX1  _1582_
timestamp 1727136778
transform -1 0 4570 0 1 270
box -12 -8 72 272
use AOI21X1  _1583_
timestamp 1727136778
transform -1 0 3910 0 -1 3390
box -12 -8 112 272
use NAND3X1  _1584_
timestamp 1727136778
transform 1 0 2970 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1585_
timestamp 1727136778
transform 1 0 3130 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1586_
timestamp 1727136778
transform 1 0 3630 0 1 2870
box -12 -8 112 272
use NAND2X1  _1587_
timestamp 1727136778
transform 1 0 2570 0 -1 270
box -12 -8 92 272
use XNOR2X1  _1588_
timestamp 1727153789
transform -1 0 4010 0 -1 270
box -12 -8 152 272
use NAND2X1  _1589_
timestamp 1727136778
transform 1 0 4950 0 1 790
box -12 -8 92 272
use OAI21X1  _1590_
timestamp 1727136778
transform 1 0 4810 0 1 790
box -12 -8 112 272
use AOI21X1  _1591_
timestamp 1727136778
transform -1 0 4850 0 -1 790
box -12 -8 112 272
use AOI22X1  _1592_
timestamp 1727136778
transform -1 0 4450 0 1 270
box -14 -8 132 272
use NAND2X1  _1593_
timestamp 1727136778
transform -1 0 4430 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1594_
timestamp 1727136778
transform 1 0 4330 0 1 2870
box -12 -8 112 272
use NAND2X1  _1595_
timestamp 1727136778
transform 1 0 4010 0 1 3910
box -12 -8 92 272
use OAI21X1  _1596_
timestamp 1727136778
transform -1 0 4230 0 1 3910
box -12 -8 112 272
use NAND2X1  _1597_
timestamp 1727136778
transform 1 0 4030 0 1 2870
box -12 -8 92 272
use OAI21X1  _1598_
timestamp 1727136778
transform -1 0 4270 0 1 2870
box -12 -8 112 272
use NAND2X1  _1599_
timestamp 1727136778
transform -1 0 3970 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1600_
timestamp 1727136778
transform -1 0 4130 0 -1 3910
box -12 -8 112 272
use NAND2X1  _1601_
timestamp 1727136778
transform 1 0 3330 0 1 3910
box -12 -8 92 272
use OAI21X1  _1602_
timestamp 1727136778
transform -1 0 3430 0 -1 4430
box -12 -8 112 272
use NAND2X1  _1603_
timestamp 1727136778
transform 1 0 2970 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1604_
timestamp 1727136778
transform -1 0 3210 0 -1 3910
box -12 -8 112 272
use NAND2X1  _1605_
timestamp 1727136778
transform -1 0 4550 0 1 3390
box -12 -8 92 272
use OAI21X1  _1606_
timestamp 1727136778
transform -1 0 5270 0 -1 3390
box -12 -8 112 272
use NAND2X1  _1607_
timestamp 1727136778
transform 1 0 4450 0 1 2350
box -12 -8 92 272
use OAI21X1  _1608_
timestamp 1727136778
transform -1 0 4670 0 1 2350
box -12 -8 112 272
use DFFPOSX1  _1609_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1726828622
transform -1 0 4790 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1610_
timestamp 1726828622
transform -1 0 3650 0 1 3910
box -13 -8 253 272
use DFFPOSX1  _1611_
timestamp 1726828622
transform -1 0 4910 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1612_
timestamp 1726828622
transform -1 0 3950 0 -1 4430
box -13 -8 253 272
use DFFPOSX1  _1613_
timestamp 1726828622
transform -1 0 3290 0 -1 4430
box -13 -8 253 272
use DFFPOSX1  _1614_
timestamp 1726828622
transform -1 0 3450 0 -1 3910
box -13 -8 253 272
use DFFPOSX1  _1615_
timestamp 1726828622
transform -1 0 5270 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1616_
timestamp 1726828622
transform 1 0 4830 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1617_
timestamp 1726828622
transform -1 0 5070 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1618_
timestamp 1726828622
transform -1 0 3870 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1619_
timestamp 1726828622
transform -1 0 4930 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1620_
timestamp 1726828622
transform 1 0 5470 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1621_
timestamp 1726828622
transform -1 0 5470 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1622_
timestamp 1726828622
transform 1 0 5090 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1623_
timestamp 1726828622
transform 1 0 4710 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1624_
timestamp 1726828622
transform -1 0 4810 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1625_
timestamp 1726828622
transform -1 0 4670 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1626_
timestamp 1726828622
transform -1 0 4370 0 -1 3910
box -13 -8 253 272
use DFFPOSX1  _1627_
timestamp 1726828622
transform -1 0 3970 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1628_
timestamp 1726828622
transform -1 0 4170 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1629_
timestamp 1726828622
transform -1 0 3050 0 -1 4430
box -13 -8 253 272
use DFFPOSX1  _1630_
timestamp 1726828622
transform -1 0 3270 0 1 3910
box -13 -8 253 272
use DFFPOSX1  _1631_
timestamp 1726828622
transform -1 0 5030 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1632_
timestamp 1726828622
transform -1 0 4710 0 -1 2350
box -13 -8 253 272
use DFFSR  _1633_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727133863
transform -1 0 5930 0 1 1310
box -12 -8 492 273
use DFFSR  _1634_
timestamp 1727133863
transform -1 0 6070 0 -1 1310
box -12 -8 492 273
use DFFSR  _1635_
timestamp 1727133863
transform -1 0 6050 0 -1 1830
box -12 -8 492 273
use INVX1  _1636_
timestamp 1727136778
transform -1 0 5970 0 -1 5470
box -12 -8 72 272
use INVX4  _1637_
timestamp 1727136778
transform 1 0 5930 0 1 5990
box -12 -8 92 272
use OAI21X1  _1638_
timestamp 1727136778
transform -1 0 5450 0 -1 5470
box -12 -8 112 272
use NOR2X1  _1639_
timestamp 1727136778
transform 1 0 5230 0 -1 5470
box -12 -8 92 272
use INVX1  _1640_
timestamp 1727136778
transform 1 0 5230 0 1 5470
box -12 -8 72 272
use INVX2  _1641_
timestamp 1727136778
transform -1 0 3810 0 1 5470
box -12 -8 72 272
use NAND2X1  _1642_
timestamp 1727136778
transform -1 0 3250 0 1 5470
box -12 -8 92 272
use INVX2  _1643_
timestamp 1727136778
transform -1 0 3070 0 -1 5990
box -12 -8 72 272
use NAND2X1  _1644_
timestamp 1727136778
transform -1 0 3950 0 1 5470
box -12 -8 92 272
use NAND2X1  _1645_
timestamp 1727136778
transform -1 0 4470 0 -1 5470
box -12 -8 92 272
use AOI22X1  _1646_
timestamp 1727136778
transform -1 0 4230 0 -1 5470
box -14 -8 132 272
use INVX2  _1647_
timestamp 1727136778
transform 1 0 3190 0 1 5990
box -12 -8 72 272
use INVX1  _1648_
timestamp 1727136778
transform 1 0 5790 0 -1 5470
box -12 -8 72 272
use INVX1  _1649_
timestamp 1727136778
transform -1 0 4350 0 -1 5470
box -12 -8 72 272
use OAI21X1  _1650_
timestamp 1727136778
transform -1 0 4550 0 1 5470
box -12 -8 112 272
use NAND2X1  _1651_
timestamp 1727136778
transform 1 0 4310 0 1 5470
box -12 -8 92 272
use NAND2X1  _1652_
timestamp 1727136778
transform -1 0 3710 0 1 5470
box -12 -8 92 272
use OAI21X1  _1653_
timestamp 1727136778
transform 1 0 4170 0 1 5470
box -12 -8 112 272
use OAI21X1  _1654_
timestamp 1727136778
transform 1 0 5810 0 1 5470
box -12 -8 112 272
use AOI21X1  _1655_
timestamp 1727136778
transform -1 0 5770 0 1 5470
box -12 -8 112 272
use NOR2X1  _1656_
timestamp 1727136778
transform 1 0 5950 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1657_
timestamp 1727136778
transform 1 0 5790 0 -1 5990
box -12 -8 112 272
use OAI21X1  _1658_
timestamp 1727136778
transform 1 0 5650 0 -1 5990
box -12 -8 112 272
use XOR2X1  _1659_
timestamp 1727152697
transform -1 0 5490 0 1 5470
box -12 -8 151 272
use NOR2X1  _1660_
timestamp 1727136778
transform -1 0 5590 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1661_
timestamp 1727136778
transform 1 0 5370 0 -1 5990
box -12 -8 112 272
use NAND2X1  _1662_
timestamp 1727136778
transform -1 0 3550 0 1 5990
box -12 -8 92 272
use NAND3X1  _1663_
timestamp 1727136778
transform -1 0 3390 0 1 5470
box -12 -8 112 272
use AOI22X1  _1664_
timestamp 1727136778
transform -1 0 3570 0 1 5470
box -14 -8 132 272
use INVX1  _1665_
timestamp 1727136778
transform -1 0 3710 0 -1 4430
box -12 -8 72 272
use NOR2X1  _1666_
timestamp 1727136778
transform -1 0 3910 0 1 4430
box -12 -8 92 272
use OAI21X1  _1667_
timestamp 1727136778
transform 1 0 3850 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1668_
timestamp 1727136778
transform 1 0 3730 0 -1 5990
box -12 -8 112 272
use OAI21X1  _1669_
timestamp 1727136778
transform -1 0 4150 0 -1 5990
box -12 -8 112 272
use AOI21X1  _1670_
timestamp 1727136778
transform 1 0 4190 0 -1 5990
box -12 -8 112 272
use INVX1  _1671_
timestamp 1727136778
transform 1 0 5250 0 1 5990
box -12 -8 72 272
use OAI21X1  _1672_
timestamp 1727136778
transform -1 0 5770 0 1 5990
box -12 -8 112 272
use MUX2X1  _1673_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform 1 0 5490 0 1 5990
box -12 -8 131 272
use NAND2X1  _1674_
timestamp 1727136778
transform -1 0 5450 0 1 5990
box -12 -8 92 272
use INVX1  _1675_
timestamp 1727136778
transform -1 0 5610 0 1 5470
box -12 -8 72 272
use OAI21X1  _1676_
timestamp 1727136778
transform 1 0 5490 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1677_
timestamp 1727136778
transform -1 0 4990 0 1 5470
box -12 -8 112 272
use MUX2X1  _1678_
timestamp 1727136778
transform -1 0 5050 0 -1 5470
box -12 -8 131 272
use NAND2X1  _1679_
timestamp 1727136778
transform -1 0 4590 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1680_
timestamp 1727136778
transform 1 0 4650 0 -1 5470
box -12 -8 92 272
use AOI21X1  _1681_
timestamp 1727136778
transform -1 0 4110 0 1 5470
box -12 -8 112 272
use NAND2X1  _1682_
timestamp 1727136778
transform 1 0 4590 0 1 5470
box -12 -8 92 272
use NAND3X1  _1683_
timestamp 1727136778
transform 1 0 4730 0 1 5470
box -12 -8 112 272
use AOI22X1  _1684_
timestamp 1727136778
transform 1 0 5050 0 1 5470
box -14 -8 132 272
use OAI21X1  _1685_
timestamp 1727136778
transform -1 0 4270 0 1 5990
box -12 -8 112 272
use OAI21X1  _1686_
timestamp 1727136778
transform 1 0 4330 0 1 5990
box -12 -8 112 272
use NAND2X1  _1687_
timestamp 1727136778
transform -1 0 5190 0 -1 5990
box -12 -8 92 272
use NAND2X1  _1688_
timestamp 1727136778
transform 1 0 5230 0 -1 5990
box -12 -8 92 272
use INVX1  _1689_
timestamp 1727136778
transform 1 0 4910 0 -1 2350
box -12 -8 72 272
use NOR2X1  _1690_
timestamp 1727136778
transform 1 0 5110 0 1 5990
box -12 -8 92 272
use OAI21X1  _1691_
timestamp 1727136778
transform -1 0 5050 0 1 5990
box -12 -8 112 272
use NAND2X1  _1692_
timestamp 1727136778
transform 1 0 3590 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1693_
timestamp 1727136778
transform 1 0 3130 0 -1 5990
box -12 -8 112 272
use AOI22X1  _1694_
timestamp 1727136778
transform -1 0 3410 0 -1 5990
box -14 -8 132 272
use INVX1  _1695_
timestamp 1727136778
transform -1 0 2990 0 1 5990
box -12 -8 72 272
use NOR2X1  _1696_
timestamp 1727136778
transform -1 0 3130 0 1 5990
box -12 -8 92 272
use OAI21X1  _1697_
timestamp 1727136778
transform -1 0 3410 0 1 5990
box -12 -8 112 272
use OAI21X1  _1698_
timestamp 1727136778
transform 1 0 3450 0 -1 5990
box -12 -8 112 272
use OAI21X1  _1699_
timestamp 1727136778
transform -1 0 3990 0 -1 5990
box -12 -8 112 272
use AOI21X1  _1700_
timestamp 1727136778
transform -1 0 4010 0 1 5990
box -12 -8 112 272
use OAI21X1  _1701_
timestamp 1727136778
transform -1 0 3690 0 1 5990
box -12 -8 112 272
use OAI21X1  _1702_
timestamp 1727136778
transform 1 0 3750 0 1 5990
box -12 -8 112 272
use XOR2X1  _1703_
timestamp 1727152697
transform -1 0 4730 0 1 5990
box -12 -8 151 272
use INVX1  _1704_
timestamp 1727136778
transform -1 0 4850 0 -1 3910
box -12 -8 72 272
use INVX1  _1705_
timestamp 1727136778
transform 1 0 4070 0 1 5990
box -12 -8 72 272
use OAI21X1  _1706_
timestamp 1727136778
transform -1 0 4450 0 -1 5990
box -12 -8 112 272
use INVX1  _1707_
timestamp 1727136778
transform -1 0 4530 0 1 5990
box -12 -8 72 272
use AOI22X1  _1708_
timestamp 1727136778
transform 1 0 4510 0 -1 5990
box -14 -8 132 272
use NAND2X1  _1709_
timestamp 1727136778
transform -1 0 3750 0 -1 4950
box -12 -8 92 272
use AND2X2  _1710_
timestamp 1727136778
transform -1 0 3970 0 1 4950
box -12 -8 112 273
use NAND2X1  _1711_
timestamp 1727136778
transform -1 0 3650 0 1 4950
box -12 -8 92 272
use AOI22X1  _1712_
timestamp 1727136778
transform -1 0 3830 0 1 4950
box -14 -8 132 272
use OAI21X1  _1713_
timestamp 1727136778
transform -1 0 3510 0 1 4950
box -12 -8 112 272
use OAI21X1  _1714_
timestamp 1727136778
transform 1 0 3790 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1715_
timestamp 1727136778
transform -1 0 4050 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1716_
timestamp 1727136778
transform 1 0 4110 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1717_
timestamp 1727136778
transform -1 0 4530 0 1 4430
box -12 -8 112 272
use OAI21X1  _1718_
timestamp 1727136778
transform 1 0 4590 0 1 4430
box -12 -8 112 272
use XOR2X1  _1719_
timestamp 1727152697
transform 1 0 4750 0 1 4430
box -12 -8 151 272
use XNOR2X1  _1720_
timestamp 1727153789
transform 1 0 4250 0 -1 4430
box -12 -8 152 272
use NAND2X1  _1721_
timestamp 1727136778
transform 1 0 4690 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1722_
timestamp 1727136778
transform 1 0 4790 0 1 5990
box -12 -8 112 272
use NAND3X1  _1723_
timestamp 1727136778
transform 1 0 4810 0 -1 5990
box -12 -8 112 272
use NAND2X1  _1724_
timestamp 1727136778
transform -1 0 4890 0 1 3910
box -12 -8 92 272
use OAI21X1  _1725_
timestamp 1727136778
transform 1 0 4450 0 -1 4430
box -12 -8 112 272
use INVX1  _1726_
timestamp 1727136778
transform -1 0 4330 0 1 3910
box -12 -8 72 272
use OAI21X1  _1727_
timestamp 1727136778
transform -1 0 4490 0 1 3910
box -12 -8 112 272
use NAND2X1  _1728_
timestamp 1727136778
transform -1 0 3110 0 1 5470
box -12 -8 92 272
use AND2X2  _1729_
timestamp 1727136778
transform 1 0 3090 0 -1 5470
box -12 -8 112 273
use NAND2X1  _1730_
timestamp 1727136778
transform -1 0 3330 0 -1 5470
box -12 -8 92 272
use AOI22X1  _1731_
timestamp 1727136778
transform -1 0 3510 0 -1 5470
box -14 -8 132 272
use OAI21X1  _1732_
timestamp 1727136778
transform 1 0 3550 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1733_
timestamp 1727136778
transform 1 0 3710 0 -1 5470
box -12 -8 112 272
use OAI21X1  _1734_
timestamp 1727136778
transform 1 0 4990 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1735_
timestamp 1727136778
transform 1 0 4930 0 1 4430
box -12 -8 112 272
use OAI21X1  _1736_
timestamp 1727136778
transform -1 0 5350 0 1 4430
box -12 -8 112 272
use OAI21X1  _1737_
timestamp 1727136778
transform 1 0 5090 0 1 4430
box -12 -8 112 272
use INVX1  _1738_
timestamp 1727136778
transform 1 0 5130 0 1 3910
box -12 -8 72 272
use XOR2X1  _1739_
timestamp 1727152697
transform 1 0 4930 0 1 3910
box -12 -8 151 272
use INVX1  _1740_
timestamp 1727136778
transform -1 0 5230 0 -1 4430
box -12 -8 72 272
use AOI21X1  _1741_
timestamp 1727136778
transform 1 0 5250 0 1 3910
box -12 -8 112 272
use NAND2X1  _1742_
timestamp 1727136778
transform 1 0 3530 0 -1 4950
box -12 -8 92 272
use AND2X2  _1743_
timestamp 1727136778
transform -1 0 2890 0 1 4950
box -12 -8 112 273
use NAND2X1  _1744_
timestamp 1727136778
transform -1 0 3030 0 1 4950
box -12 -8 92 272
use AOI22X1  _1745_
timestamp 1727136778
transform -1 0 3350 0 1 4950
box -14 -8 132 272
use OAI21X1  _1746_
timestamp 1727136778
transform 1 0 3090 0 1 4950
box -12 -8 112 272
use OAI21X1  _1747_
timestamp 1727136778
transform 1 0 3390 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1748_
timestamp 1727136778
transform -1 0 5190 0 1 4950
box -12 -8 112 272
use AOI21X1  _1749_
timestamp 1727136778
transform 1 0 5250 0 1 4950
box -12 -8 112 272
use OAI21X1  _1750_
timestamp 1727136778
transform 1 0 5470 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1751_
timestamp 1727136778
transform 1 0 5390 0 1 4430
box -12 -8 112 272
use INVX1  _1752_
timestamp 1727136778
transform -1 0 5350 0 -1 4430
box -12 -8 72 272
use XOR2X1  _1753_
timestamp 1727152697
transform 1 0 5410 0 1 3910
box -12 -8 151 272
use INVX1  _1754_
timestamp 1727136778
transform 1 0 5170 0 1 1830
box -12 -8 72 272
use OAI21X1  _1755_
timestamp 1727136778
transform 1 0 5410 0 -1 4430
box -12 -8 112 272
use INVX1  _1756_
timestamp 1727136778
transform 1 0 4870 0 -1 4950
box -12 -8 72 272
use AND2X2  _1757_
timestamp 1727136778
transform -1 0 4490 0 -1 4950
box -12 -8 112 273
use NAND2X1  _1758_
timestamp 1727136778
transform 1 0 4270 0 -1 4950
box -12 -8 92 272
use AOI22X1  _1759_
timestamp 1727136778
transform 1 0 4030 0 1 4950
box -14 -8 132 272
use OAI21X1  _1760_
timestamp 1727136778
transform 1 0 4550 0 -1 4950
box -12 -8 112 272
use OAI22X1  _1761_
timestamp 1727136778
transform -1 0 4810 0 -1 4950
box -12 -8 132 272
use OAI21X1  _1762_
timestamp 1727136778
transform -1 0 5250 0 -1 4950
box -12 -8 112 272
use AOI21X1  _1763_
timestamp 1727136778
transform 1 0 5310 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1764_
timestamp 1727136778
transform 1 0 5610 0 -1 4950
box -12 -8 112 272
use OAI21X1  _1765_
timestamp 1727136778
transform 1 0 5770 0 -1 4950
box -12 -8 112 272
use NAND2X1  _1766_
timestamp 1727136778
transform 1 0 5870 0 -1 3910
box -12 -8 92 272
use INVX1  _1767_
timestamp 1727136778
transform 1 0 4910 0 -1 4430
box -12 -8 72 272
use AOI21X1  _1768_
timestamp 1727136778
transform -1 0 4870 0 -1 4430
box -12 -8 112 272
use AOI21X1  _1769_
timestamp 1727136778
transform -1 0 4710 0 -1 4430
box -12 -8 112 272
use OAI21X1  _1770_
timestamp 1727136778
transform -1 0 5110 0 -1 4430
box -12 -8 112 272
use OR2X2  _1771_
timestamp 1727136778
transform 1 0 5550 0 1 4430
box -12 -8 112 272
use AOI22X1  _1772_
timestamp 1727136778
transform 1 0 5570 0 -1 4430
box -14 -8 132 272
use INVX1  _1773_
timestamp 1727136778
transform -1 0 5870 0 1 5990
box -12 -8 72 272
use NAND2X1  _1774_
timestamp 1727136778
transform -1 0 5690 0 1 3910
box -12 -8 92 272
use NAND2X1  _1775_
timestamp 1727136778
transform -1 0 5810 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1776_
timestamp 1727136778
transform 1 0 5730 0 -1 4430
box -12 -8 112 272
use NAND2X1  _1777_
timestamp 1727136778
transform 1 0 4970 0 1 4950
box -12 -8 92 272
use AND2X2  _1778_
timestamp 1727136778
transform 1 0 4510 0 1 4950
box -12 -8 112 273
use NAND2X1  _1779_
timestamp 1727136778
transform 1 0 4370 0 1 4950
box -12 -8 92 272
use AOI22X1  _1780_
timestamp 1727136778
transform 1 0 4210 0 1 4950
box -14 -8 132 272
use OAI21X1  _1781_
timestamp 1727136778
transform 1 0 4670 0 1 4950
box -12 -8 112 272
use OAI21X1  _1782_
timestamp 1727136778
transform 1 0 4810 0 1 4950
box -12 -8 112 272
use OAI21X1  _1783_
timestamp 1727136778
transform 1 0 5650 0 -1 5470
box -12 -8 112 272
use AOI21X1  _1784_
timestamp 1727136778
transform 1 0 5510 0 1 4950
box -12 -8 112 272
use OAI21X1  _1785_
timestamp 1727136778
transform -1 0 5930 0 1 4950
box -12 -8 112 272
use OAI21X1  _1786_
timestamp 1727136778
transform 1 0 5970 0 1 4950
box -12 -8 112 272
use NAND2X1  _1787_
timestamp 1727136778
transform -1 0 5990 0 -1 270
box -12 -8 92 272
use NAND2X1  _1788_
timestamp 1727136778
transform 1 0 5750 0 1 3910
box -12 -8 92 272
use INVX1  _1789_
timestamp 1727136778
transform 1 0 6010 0 -1 4430
box -12 -8 72 272
use NAND3X1  _1790_
timestamp 1727136778
transform 1 0 6030 0 1 3910
box -12 -8 112 272
use NAND2X1  _1791_
timestamp 1727136778
transform 1 0 6010 0 1 2350
box -12 -8 92 272
use NOR2X1  _1792_
timestamp 1727136778
transform 1 0 4670 0 1 3910
box -12 -8 92 272
use NAND2X1  _1793_
timestamp 1727136778
transform 1 0 4550 0 1 3910
box -12 -8 92 272
use NOR2X1  _1794_
timestamp 1727136778
transform 1 0 4910 0 -1 3910
box -12 -8 92 272
use NAND3X1  _1795_
timestamp 1727136778
transform -1 0 5670 0 -1 3910
box -12 -8 112 272
use NOR2X1  _1796_
timestamp 1727136778
transform 1 0 5450 0 -1 3910
box -12 -8 92 272
use AND2X2  _1797_
timestamp 1727136778
transform -1 0 5150 0 -1 3910
box -12 -8 112 273
use NAND3X1  _1798_
timestamp 1727136778
transform -1 0 5970 0 1 3910
box -12 -8 112 272
use NAND2X1  _1799_
timestamp 1727136778
transform -1 0 5970 0 -1 4430
box -12 -8 92 272
use NAND2X1  _1800_
timestamp 1727136778
transform -1 0 5950 0 1 3390
box -12 -8 92 272
use NAND2X1  _1801_
timestamp 1727136778
transform 1 0 5430 0 1 3390
box -12 -8 92 272
use NOR2X1  _1802_
timestamp 1727136778
transform 1 0 4790 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1803_
timestamp 1727136778
transform 1 0 5910 0 1 270
box -12 -8 112 272
use NOR2X1  _1804_
timestamp 1727136778
transform -1 0 5970 0 1 4430
box -12 -8 92 272
use AOI21X1  _1805_
timestamp 1727136778
transform 1 0 6030 0 1 4430
box -12 -8 112 272
use XOR2X1  _1806_
timestamp 1727152697
transform -1 0 5850 0 1 4430
box -12 -8 151 272
use OAI21X1  _1807_
timestamp 1727136778
transform 1 0 5710 0 1 3390
box -12 -8 112 272
use NAND3X1  _1808_
timestamp 1727136778
transform 1 0 5550 0 1 3390
box -12 -8 112 272
use AOI21X1  _1809_
timestamp 1727136778
transform 1 0 5670 0 1 4950
box -12 -8 112 272
use XOR2X1  _1810_
timestamp 1727152697
transform 1 0 5930 0 -1 4950
box -12 -8 151 272
use NAND3X1  _1811_
timestamp 1727136778
transform 1 0 5750 0 1 270
box -12 -8 112 272
use INVX1  _1812_
timestamp 1727136778
transform 1 0 6010 0 -1 3910
box -12 -8 72 272
use NAND3X1  _1813_
timestamp 1727136778
transform -1 0 6110 0 1 3390
box -12 -8 112 272
use NAND2X1  _1814_
timestamp 1727136778
transform -1 0 6090 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1815_
timestamp 1727136778
transform 1 0 5870 0 -1 3390
box -12 -8 112 272
use NAND3X1  _1816_
timestamp 1727136778
transform -1 0 6110 0 1 2870
box -12 -8 112 272
use NAND2X1  _1817_
timestamp 1727136778
transform -1 0 5950 0 1 2870
box -12 -8 92 272
use BUFX2  _1818_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 3370 0 -1 2350
box -12 -8 92 272
use BUFX2  _1819_
timestamp 1727136778
transform -1 0 2690 0 -1 2350
box -12 -8 92 272
use BUFX2  _1820_
timestamp 1727136778
transform -1 0 4690 0 -1 1310
box -12 -8 92 272
use BUFX2  _1821_
timestamp 1727136778
transform -1 0 5730 0 -1 270
box -12 -8 92 272
use BUFX2  _1822_
timestamp 1727136778
transform 1 0 5510 0 -1 270
box -12 -8 92 272
use BUFX2  _1823_
timestamp 1727136778
transform 1 0 5370 0 -1 270
box -12 -8 92 272
use BUFX2  _1824_
timestamp 1727136778
transform 1 0 5010 0 -1 270
box -12 -8 92 272
use BUFX2  _1825_
timestamp 1727136778
transform 1 0 4630 0 -1 270
box -12 -8 92 272
use BUFX2  _1826_
timestamp 1727136778
transform 1 0 5770 0 -1 270
box -12 -8 92 272
use BUFX2  BUFX2_insert0
timestamp 1727136778
transform 1 0 3970 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert1
timestamp 1727136778
transform -1 0 2310 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert2
timestamp 1727136778
transform -1 0 2410 0 1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert3
timestamp 1727136778
transform -1 0 2370 0 -1 3910
box -12 -8 92 272
use BUFX2  BUFX2_insert4
timestamp 1727136778
transform -1 0 4510 0 -1 3910
box -12 -8 92 272
use BUFX2  BUFX2_insert5
timestamp 1727136778
transform -1 0 3850 0 -1 3910
box -12 -8 92 272
use BUFX2  BUFX2_insert6
timestamp 1727136778
transform -1 0 2830 0 -1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert7
timestamp 1727136778
transform -1 0 3510 0 -1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert13
timestamp 1727136778
transform 1 0 5230 0 1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert14
timestamp 1727136778
transform -1 0 3930 0 1 3390
box -12 -8 92 272
use BUFX2  BUFX2_insert15
timestamp 1727136778
transform -1 0 4430 0 1 3390
box -12 -8 92 272
use BUFX2  BUFX2_insert16
timestamp 1727136778
transform -1 0 4130 0 -1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert17
timestamp 1727136778
transform 1 0 2570 0 1 3910
box -12 -8 92 272
use BUFX2  BUFX2_insert18
timestamp 1727136778
transform -1 0 2430 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert19
timestamp 1727136778
transform 1 0 3070 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert20
timestamp 1727136778
transform -1 0 2530 0 1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert21
timestamp 1727136778
transform 1 0 5350 0 1 2870
box -12 -8 92 272
use BUFX2  BUFX2_insert22
timestamp 1727136778
transform -1 0 4310 0 1 3390
box -12 -8 92 272
use BUFX2  BUFX2_insert23
timestamp 1727136778
transform 1 0 4290 0 -1 3390
box -12 -8 92 272
use BUFX2  BUFX2_insert24
timestamp 1727136778
transform 1 0 5310 0 -1 3390
box -12 -8 92 272
use BUFX2  BUFX2_insert25
timestamp 1727136778
transform -1 0 2450 0 -1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert26
timestamp 1727136778
transform -1 0 2750 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert27
timestamp 1727136778
transform -1 0 2490 0 -1 3910
box -12 -8 92 272
use BUFX2  BUFX2_insert28
timestamp 1727136778
transform 1 0 3210 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert29
timestamp 1727136778
transform -1 0 2290 0 1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert30
timestamp 1727136778
transform 1 0 3410 0 1 2350
box -12 -8 92 272
use BUFX2  BUFX2_insert31
timestamp 1727136778
transform -1 0 2310 0 -1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert32
timestamp 1727136778
transform 1 0 3550 0 1 4430
box -12 -8 92 272
use BUFX2  BUFX2_insert33
timestamp 1727136778
transform -1 0 5170 0 -1 5470
box -12 -8 92 272
use BUFX2  BUFX2_insert34
timestamp 1727136778
transform -1 0 6110 0 -1 5470
box -12 -8 92 272
use BUFX2  BUFX2_insert35
timestamp 1727136778
transform -1 0 5050 0 -1 5990
box -12 -8 92 272
use BUFX2  BUFX2_insert36
timestamp 1727136778
transform -1 0 6050 0 1 5470
box -12 -8 92 272
use CLKBUF1  CLKBUF1_insert8 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1727136778
transform -1 0 4750 0 -1 3910
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert9
timestamp 1727136778
transform -1 0 5170 0 1 2870
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert10
timestamp 1727136778
transform -1 0 6030 0 1 790
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert11
timestamp 1727136778
transform -1 0 5390 0 -1 3910
box -12 -8 212 272
use CLKBUF1  CLKBUF1_insert12
timestamp 1727136778
transform -1 0 5190 0 -1 1310
box -12 -8 212 272
use FILL  FILL89850x150 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1700315010
transform -1 0 6010 0 -1 270
box -12 -8 32 272
use FILL  FILL90150x150
timestamp 1700315010
transform -1 0 6030 0 -1 270
box -12 -8 32 272
use FILL  FILL90150x4050
timestamp 1700315010
transform 1 0 6010 0 1 270
box -12 -8 32 272
use FILL  FILL90150x89850
timestamp 1700315010
transform 1 0 6010 0 1 5990
box -12 -8 32 272
use FILL  FILL90450x150
timestamp 1700315010
transform -1 0 6050 0 -1 270
box -12 -8 32 272
use FILL  FILL90450x4050
timestamp 1700315010
transform 1 0 6030 0 1 270
box -12 -8 32 272
use FILL  FILL90450x7950
timestamp 1700315010
transform -1 0 6050 0 -1 790
box -12 -8 32 272
use FILL  FILL90450x11850
timestamp 1700315010
transform 1 0 6030 0 1 790
box -12 -8 32 272
use FILL  FILL90450x27450
timestamp 1700315010
transform 1 0 6030 0 1 1830
box -12 -8 32 272
use FILL  FILL90450x31350
timestamp 1700315010
transform -1 0 6050 0 -1 2350
box -12 -8 32 272
use FILL  FILL90450x85950
timestamp 1700315010
transform -1 0 6050 0 -1 5990
box -12 -8 32 272
use FILL  FILL90450x89850
timestamp 1700315010
transform 1 0 6030 0 1 5990
box -12 -8 32 272
use FILL  FILL90750x150
timestamp 1700315010
transform -1 0 6070 0 -1 270
box -12 -8 32 272
use FILL  FILL90750x4050
timestamp 1700315010
transform 1 0 6050 0 1 270
box -12 -8 32 272
use FILL  FILL90750x7950
timestamp 1700315010
transform -1 0 6070 0 -1 790
box -12 -8 32 272
use FILL  FILL90750x11850
timestamp 1700315010
transform 1 0 6050 0 1 790
box -12 -8 32 272
use FILL  FILL90750x19650
timestamp 1700315010
transform 1 0 6050 0 1 1310
box -12 -8 32 272
use FILL  FILL90750x23550
timestamp 1700315010
transform -1 0 6070 0 -1 1830
box -12 -8 32 272
use FILL  FILL90750x27450
timestamp 1700315010
transform 1 0 6050 0 1 1830
box -12 -8 32 272
use FILL  FILL90750x31350
timestamp 1700315010
transform -1 0 6070 0 -1 2350
box -12 -8 32 272
use FILL  FILL90750x39150
timestamp 1700315010
transform -1 0 6070 0 -1 2870
box -12 -8 32 272
use FILL  FILL90750x82050
timestamp 1700315010
transform 1 0 6050 0 1 5470
box -12 -8 32 272
use FILL  FILL90750x85950
timestamp 1700315010
transform -1 0 6070 0 -1 5990
box -12 -8 32 272
use FILL  FILL90750x89850
timestamp 1700315010
transform 1 0 6050 0 1 5990
box -12 -8 32 272
use FILL  FILL91050x150
timestamp 1700315010
transform -1 0 6090 0 -1 270
box -12 -8 32 272
use FILL  FILL91050x4050
timestamp 1700315010
transform 1 0 6070 0 1 270
box -12 -8 32 272
use FILL  FILL91050x7950
timestamp 1700315010
transform -1 0 6090 0 -1 790
box -12 -8 32 272
use FILL  FILL91050x11850
timestamp 1700315010
transform 1 0 6070 0 1 790
box -12 -8 32 272
use FILL  FILL91050x15750
timestamp 1700315010
transform -1 0 6090 0 -1 1310
box -12 -8 32 272
use FILL  FILL91050x19650
timestamp 1700315010
transform 1 0 6070 0 1 1310
box -12 -8 32 272
use FILL  FILL91050x23550
timestamp 1700315010
transform -1 0 6090 0 -1 1830
box -12 -8 32 272
use FILL  FILL91050x27450
timestamp 1700315010
transform 1 0 6070 0 1 1830
box -12 -8 32 272
use FILL  FILL91050x31350
timestamp 1700315010
transform -1 0 6090 0 -1 2350
box -12 -8 32 272
use FILL  FILL91050x39150
timestamp 1700315010
transform -1 0 6090 0 -1 2870
box -12 -8 32 272
use FILL  FILL91050x54750
timestamp 1700315010
transform -1 0 6090 0 -1 3910
box -12 -8 32 272
use FILL  FILL91050x62550
timestamp 1700315010
transform -1 0 6090 0 -1 4430
box -12 -8 32 272
use FILL  FILL91050x70350
timestamp 1700315010
transform -1 0 6090 0 -1 4950
box -12 -8 32 272
use FILL  FILL91050x74250
timestamp 1700315010
transform 1 0 6070 0 1 4950
box -12 -8 32 272
use FILL  FILL91050x82050
timestamp 1700315010
transform 1 0 6070 0 1 5470
box -12 -8 32 272
use FILL  FILL91050x85950
timestamp 1700315010
transform -1 0 6090 0 -1 5990
box -12 -8 32 272
use FILL  FILL91050x89850
timestamp 1700315010
transform 1 0 6070 0 1 5990
box -12 -8 32 272
use FILL  FILL91350x150
timestamp 1700315010
transform -1 0 6110 0 -1 270
box -12 -8 32 272
use FILL  FILL91350x4050
timestamp 1700315010
transform 1 0 6090 0 1 270
box -12 -8 32 272
use FILL  FILL91350x7950
timestamp 1700315010
transform -1 0 6110 0 -1 790
box -12 -8 32 272
use FILL  FILL91350x11850
timestamp 1700315010
transform 1 0 6090 0 1 790
box -12 -8 32 272
use FILL  FILL91350x15750
timestamp 1700315010
transform -1 0 6110 0 -1 1310
box -12 -8 32 272
use FILL  FILL91350x19650
timestamp 1700315010
transform 1 0 6090 0 1 1310
box -12 -8 32 272
use FILL  FILL91350x23550
timestamp 1700315010
transform -1 0 6110 0 -1 1830
box -12 -8 32 272
use FILL  FILL91350x27450
timestamp 1700315010
transform 1 0 6090 0 1 1830
box -12 -8 32 272
use FILL  FILL91350x31350
timestamp 1700315010
transform -1 0 6110 0 -1 2350
box -12 -8 32 272
use FILL  FILL91350x35250
timestamp 1700315010
transform 1 0 6090 0 1 2350
box -12 -8 32 272
use FILL  FILL91350x39150
timestamp 1700315010
transform -1 0 6110 0 -1 2870
box -12 -8 32 272
use FILL  FILL91350x46950
timestamp 1700315010
transform -1 0 6110 0 -1 3390
box -12 -8 32 272
use FILL  FILL91350x54750
timestamp 1700315010
transform -1 0 6110 0 -1 3910
box -12 -8 32 272
use FILL  FILL91350x62550
timestamp 1700315010
transform -1 0 6110 0 -1 4430
box -12 -8 32 272
use FILL  FILL91350x70350
timestamp 1700315010
transform -1 0 6110 0 -1 4950
box -12 -8 32 272
use FILL  FILL91350x74250
timestamp 1700315010
transform 1 0 6090 0 1 4950
box -12 -8 32 272
use FILL  FILL91350x82050
timestamp 1700315010
transform 1 0 6090 0 1 5470
box -12 -8 32 272
use FILL  FILL91350x85950
timestamp 1700315010
transform -1 0 6110 0 -1 5990
box -12 -8 32 272
use FILL  FILL91350x89850
timestamp 1700315010
transform 1 0 6090 0 1 5990
box -12 -8 32 272
use FILL  FILL91650x150
timestamp 1700315010
transform -1 0 6130 0 -1 270
box -12 -8 32 272
use FILL  FILL91650x4050
timestamp 1700315010
transform 1 0 6110 0 1 270
box -12 -8 32 272
use FILL  FILL91650x7950
timestamp 1700315010
transform -1 0 6130 0 -1 790
box -12 -8 32 272
use FILL  FILL91650x11850
timestamp 1700315010
transform 1 0 6110 0 1 790
box -12 -8 32 272
use FILL  FILL91650x15750
timestamp 1700315010
transform -1 0 6130 0 -1 1310
box -12 -8 32 272
use FILL  FILL91650x19650
timestamp 1700315010
transform 1 0 6110 0 1 1310
box -12 -8 32 272
use FILL  FILL91650x23550
timestamp 1700315010
transform -1 0 6130 0 -1 1830
box -12 -8 32 272
use FILL  FILL91650x27450
timestamp 1700315010
transform 1 0 6110 0 1 1830
box -12 -8 32 272
use FILL  FILL91650x31350
timestamp 1700315010
transform -1 0 6130 0 -1 2350
box -12 -8 32 272
use FILL  FILL91650x35250
timestamp 1700315010
transform 1 0 6110 0 1 2350
box -12 -8 32 272
use FILL  FILL91650x39150
timestamp 1700315010
transform -1 0 6130 0 -1 2870
box -12 -8 32 272
use FILL  FILL91650x43050
timestamp 1700315010
transform 1 0 6110 0 1 2870
box -12 -8 32 272
use FILL  FILL91650x46950
timestamp 1700315010
transform -1 0 6130 0 -1 3390
box -12 -8 32 272
use FILL  FILL91650x50850
timestamp 1700315010
transform 1 0 6110 0 1 3390
box -12 -8 32 272
use FILL  FILL91650x54750
timestamp 1700315010
transform -1 0 6130 0 -1 3910
box -12 -8 32 272
use FILL  FILL91650x62550
timestamp 1700315010
transform -1 0 6130 0 -1 4430
box -12 -8 32 272
use FILL  FILL91650x70350
timestamp 1700315010
transform -1 0 6130 0 -1 4950
box -12 -8 32 272
use FILL  FILL91650x74250
timestamp 1700315010
transform 1 0 6110 0 1 4950
box -12 -8 32 272
use FILL  FILL91650x78150
timestamp 1700315010
transform -1 0 6130 0 -1 5470
box -12 -8 32 272
use FILL  FILL91650x82050
timestamp 1700315010
transform 1 0 6110 0 1 5470
box -12 -8 32 272
use FILL  FILL91650x85950
timestamp 1700315010
transform -1 0 6130 0 -1 5990
box -12 -8 32 272
use FILL  FILL91650x89850
timestamp 1700315010
transform 1 0 6110 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__889_
timestamp 1700315010
transform 1 0 5330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__890_
timestamp 1700315010
transform -1 0 4950 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__891_
timestamp 1700315010
transform -1 0 5090 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__892_
timestamp 1700315010
transform 1 0 5350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__893_
timestamp 1700315010
transform -1 0 5210 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__894_
timestamp 1700315010
transform 1 0 5470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__895_
timestamp 1700315010
transform -1 0 5230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__896_
timestamp 1700315010
transform -1 0 5090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__897_
timestamp 1700315010
transform 1 0 5090 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__898_
timestamp 1700315010
transform -1 0 5470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__899_
timestamp 1700315010
transform 1 0 5230 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__900_
timestamp 1700315010
transform -1 0 5830 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__901_
timestamp 1700315010
transform -1 0 5690 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__902_
timestamp 1700315010
transform 1 0 5770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__903_
timestamp 1700315010
transform 1 0 4870 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__904_
timestamp 1700315010
transform -1 0 5330 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__905_
timestamp 1700315010
transform -1 0 5670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__906_
timestamp 1700315010
transform -1 0 4190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__907_
timestamp 1700315010
transform 1 0 4970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__908_
timestamp 1700315010
transform 1 0 5930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__909_
timestamp 1700315010
transform 1 0 5570 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__910_
timestamp 1700315010
transform 1 0 5510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__911_
timestamp 1700315010
transform 1 0 5390 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__912_
timestamp 1700315010
transform 1 0 5730 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__913_
timestamp 1700315010
transform -1 0 5550 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__914_
timestamp 1700315010
transform -1 0 5230 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__915_
timestamp 1700315010
transform 1 0 5210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__916_
timestamp 1700315010
transform -1 0 5610 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__917_
timestamp 1700315010
transform 1 0 5810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__918_
timestamp 1700315010
transform -1 0 5370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__919_
timestamp 1700315010
transform 1 0 5370 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__920_
timestamp 1700315010
transform -1 0 5550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__921_
timestamp 1700315010
transform 1 0 5630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__922_
timestamp 1700315010
transform 1 0 5350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__923_
timestamp 1700315010
transform 1 0 5890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__924_
timestamp 1700315010
transform 1 0 5870 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__925_
timestamp 1700315010
transform -1 0 5950 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__926_
timestamp 1700315010
transform -1 0 4310 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__927_
timestamp 1700315010
transform 1 0 4830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__928_
timestamp 1700315010
transform 1 0 4670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__929_
timestamp 1700315010
transform 1 0 4190 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__930_
timestamp 1700315010
transform 1 0 3650 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__931_
timestamp 1700315010
transform -1 0 3810 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__932_
timestamp 1700315010
transform 1 0 4110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__933_
timestamp 1700315010
transform -1 0 4390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__934_
timestamp 1700315010
transform 1 0 4510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__935_
timestamp 1700315010
transform -1 0 5370 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__936_
timestamp 1700315010
transform 1 0 4050 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__937_
timestamp 1700315010
transform -1 0 3970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__938_
timestamp 1700315010
transform -1 0 3970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__939_
timestamp 1700315010
transform 1 0 3630 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__940_
timestamp 1700315010
transform 1 0 3430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__941_
timestamp 1700315010
transform -1 0 3230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__942_
timestamp 1700315010
transform 1 0 3610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__943_
timestamp 1700315010
transform 1 0 3450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__944_
timestamp 1700315010
transform -1 0 5290 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__945_
timestamp 1700315010
transform 1 0 5550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__946_
timestamp 1700315010
transform 1 0 5390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__947_
timestamp 1700315010
transform 1 0 5630 0 1 790
box -12 -8 32 272
use FILL  FILL_0__948_
timestamp 1700315010
transform 1 0 5230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__949_
timestamp 1700315010
transform 1 0 5070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__950_
timestamp 1700315010
transform -1 0 4630 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__951_
timestamp 1700315010
transform 1 0 3890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__952_
timestamp 1700315010
transform 1 0 2310 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__953_
timestamp 1700315010
transform 1 0 2610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__954_
timestamp 1700315010
transform -1 0 2470 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__955_
timestamp 1700315010
transform 1 0 2730 0 1 790
box -12 -8 32 272
use FILL  FILL_0__956_
timestamp 1700315010
transform 1 0 3150 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__957_
timestamp 1700315010
transform 1 0 3470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__958_
timestamp 1700315010
transform 1 0 3590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__959_
timestamp 1700315010
transform 1 0 3590 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__960_
timestamp 1700315010
transform 1 0 3150 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__961_
timestamp 1700315010
transform -1 0 3450 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__962_
timestamp 1700315010
transform 1 0 3750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__963_
timestamp 1700315010
transform 1 0 2890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__964_
timestamp 1700315010
transform -1 0 2630 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__965_
timestamp 1700315010
transform 1 0 2470 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__966_
timestamp 1700315010
transform 1 0 3310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__967_
timestamp 1700315010
transform -1 0 2910 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__968_
timestamp 1700315010
transform 1 0 2550 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__969_
timestamp 1700315010
transform -1 0 2750 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__970_
timestamp 1700315010
transform 1 0 3010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__971_
timestamp 1700315010
transform 1 0 3010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__972_
timestamp 1700315010
transform -1 0 3170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__973_
timestamp 1700315010
transform 1 0 3010 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__974_
timestamp 1700315010
transform -1 0 3470 0 1 790
box -12 -8 32 272
use FILL  FILL_0__975_
timestamp 1700315010
transform 1 0 3030 0 1 790
box -12 -8 32 272
use FILL  FILL_0__976_
timestamp 1700315010
transform 1 0 2590 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__977_
timestamp 1700315010
transform 1 0 2090 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__978_
timestamp 1700315010
transform 1 0 2470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__979_
timestamp 1700315010
transform 1 0 2070 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__980_
timestamp 1700315010
transform 1 0 2870 0 1 790
box -12 -8 32 272
use FILL  FILL_0__981_
timestamp 1700315010
transform 1 0 3610 0 1 790
box -12 -8 32 272
use FILL  FILL_0__982_
timestamp 1700315010
transform -1 0 3450 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__983_
timestamp 1700315010
transform -1 0 2730 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__984_
timestamp 1700315010
transform -1 0 2410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__985_
timestamp 1700315010
transform -1 0 2330 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__986_
timestamp 1700315010
transform -1 0 1710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__987_
timestamp 1700315010
transform -1 0 1570 0 1 790
box -12 -8 32 272
use FILL  FILL_0__988_
timestamp 1700315010
transform -1 0 1350 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__989_
timestamp 1700315010
transform -1 0 1790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__990_
timestamp 1700315010
transform 1 0 1830 0 1 790
box -12 -8 32 272
use FILL  FILL_0__991_
timestamp 1700315010
transform 1 0 2370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__992_
timestamp 1700315010
transform -1 0 2370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__993_
timestamp 1700315010
transform 1 0 1990 0 1 790
box -12 -8 32 272
use FILL  FILL_0__994_
timestamp 1700315010
transform 1 0 2570 0 1 790
box -12 -8 32 272
use FILL  FILL_0__995_
timestamp 1700315010
transform -1 0 2770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__996_
timestamp 1700315010
transform 1 0 1670 0 1 790
box -12 -8 32 272
use FILL  FILL_0__997_
timestamp 1700315010
transform -1 0 1410 0 1 790
box -12 -8 32 272
use FILL  FILL_0__998_
timestamp 1700315010
transform 1 0 1590 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__999_
timestamp 1700315010
transform 1 0 2170 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1000_
timestamp 1700315010
transform 1 0 2210 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1001_
timestamp 1700315010
transform 1 0 2750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1002_
timestamp 1700315010
transform 1 0 2310 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1003_
timestamp 1700315010
transform -1 0 2930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1004_
timestamp 1700315010
transform 1 0 2450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1005_
timestamp 1700315010
transform -1 0 2310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1006_
timestamp 1700315010
transform 1 0 2010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1007_
timestamp 1700315010
transform -1 0 1650 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1008_
timestamp 1700315010
transform 1 0 1750 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1009_
timestamp 1700315010
transform -1 0 1930 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1010_
timestamp 1700315010
transform 1 0 2290 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1011_
timestamp 1700315010
transform -1 0 2190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1012_
timestamp 1700315010
transform -1 0 1450 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1013_
timestamp 1700315010
transform -1 0 2450 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1014_
timestamp 1700315010
transform -1 0 2170 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1015_
timestamp 1700315010
transform -1 0 2030 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1016_
timestamp 1700315010
transform -1 0 2050 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1017_
timestamp 1700315010
transform 1 0 2170 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1018_
timestamp 1700315010
transform -1 0 2350 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1019_
timestamp 1700315010
transform -1 0 1750 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1020_
timestamp 1700315010
transform -1 0 1490 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1021_
timestamp 1700315010
transform -1 0 1410 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1022_
timestamp 1700315010
transform -1 0 1370 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1023_
timestamp 1700315010
transform 1 0 1110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1024_
timestamp 1700315010
transform 1 0 1470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1025_
timestamp 1700315010
transform 1 0 1430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1026_
timestamp 1700315010
transform 1 0 1230 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1027_
timestamp 1700315010
transform 1 0 1470 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1028_
timestamp 1700315010
transform 1 0 1030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1029_
timestamp 1700315010
transform -1 0 890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1030_
timestamp 1700315010
transform -1 0 1570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1031_
timestamp 1700315010
transform 1 0 1270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1032_
timestamp 1700315010
transform -1 0 1210 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1033_
timestamp 1700315010
transform -1 0 1050 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1034_
timestamp 1700315010
transform -1 0 1630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1035_
timestamp 1700315010
transform -1 0 1070 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1036_
timestamp 1700315010
transform -1 0 1150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1037_
timestamp 1700315010
transform -1 0 1030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1038_
timestamp 1700315010
transform 1 0 1610 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1039_
timestamp 1700315010
transform -1 0 1310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1040_
timestamp 1700315010
transform -1 0 2030 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1041_
timestamp 1700315010
transform -1 0 2630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1042_
timestamp 1700315010
transform 1 0 1870 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1043_
timestamp 1700315010
transform 1 0 2270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1044_
timestamp 1700315010
transform 1 0 2230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1045_
timestamp 1700315010
transform 1 0 2070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1046_
timestamp 1700315010
transform -1 0 1590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1047_
timestamp 1700315010
transform 1 0 1730 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1048_
timestamp 1700315010
transform -1 0 1930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1049_
timestamp 1700315010
transform -1 0 1430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1050_
timestamp 1700315010
transform 1 0 1470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1051_
timestamp 1700315010
transform -1 0 670 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1052_
timestamp 1700315010
transform 1 0 1170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1053_
timestamp 1700315010
transform 1 0 1190 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1054_
timestamp 1700315010
transform -1 0 1350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1055_
timestamp 1700315010
transform -1 0 930 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1056_
timestamp 1700315010
transform 1 0 970 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1057_
timestamp 1700315010
transform -1 0 1890 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1058_
timestamp 1700315010
transform 1 0 1230 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1059_
timestamp 1700315010
transform 1 0 1070 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1060_
timestamp 1700315010
transform -1 0 1150 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1061_
timestamp 1700315010
transform -1 0 2910 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1062_
timestamp 1700315010
transform -1 0 1890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1063_
timestamp 1700315010
transform 1 0 2150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1064_
timestamp 1700315010
transform 1 0 1350 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1065_
timestamp 1700315010
transform -1 0 910 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1066_
timestamp 1700315010
transform 1 0 1010 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1067_
timestamp 1700315010
transform 1 0 1270 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1068_
timestamp 1700315010
transform -1 0 830 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1069_
timestamp 1700315010
transform 1 0 1210 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1070_
timestamp 1700315010
transform 1 0 1930 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1071_
timestamp 1700315010
transform 1 0 1550 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1072_
timestamp 1700315010
transform -1 0 190 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1073_
timestamp 1700315010
transform -1 0 930 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1074_
timestamp 1700315010
transform -1 0 770 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1075_
timestamp 1700315010
transform -1 0 770 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1076_
timestamp 1700315010
transform -1 0 950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1077_
timestamp 1700315010
transform 1 0 1090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1078_
timestamp 1700315010
transform -1 0 470 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1079_
timestamp 1700315010
transform -1 0 870 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1080_
timestamp 1700315010
transform -1 0 830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1081_
timestamp 1700315010
transform -1 0 190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1082_
timestamp 1700315010
transform -1 0 1010 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1083_
timestamp 1700315010
transform -1 0 730 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1084_
timestamp 1700315010
transform -1 0 350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1085_
timestamp 1700315010
transform -1 0 330 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1086_
timestamp 1700315010
transform 1 0 650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1087_
timestamp 1700315010
transform 1 0 490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1088_
timestamp 1700315010
transform -1 0 610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1089_
timestamp 1700315010
transform 1 0 1930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1090_
timestamp 1700315010
transform 1 0 1530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1091_
timestamp 1700315010
transform -1 0 1870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1092_
timestamp 1700315010
transform -1 0 2010 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1093_
timestamp 1700315010
transform 1 0 1850 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1094_
timestamp 1700315010
transform 1 0 2150 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1095_
timestamp 1700315010
transform -1 0 1830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1096_
timestamp 1700315010
transform -1 0 1670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1097_
timestamp 1700315010
transform -1 0 1570 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1098_
timestamp 1700315010
transform -1 0 1710 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1099_
timestamp 1700315010
transform -1 0 1410 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1100_
timestamp 1700315010
transform -1 0 30 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1101_
timestamp 1700315010
transform -1 0 30 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1102_
timestamp 1700315010
transform -1 0 910 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1103_
timestamp 1700315010
transform 1 0 590 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1104_
timestamp 1700315010
transform 1 0 450 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1105_
timestamp 1700315010
transform 1 0 150 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1106_
timestamp 1700315010
transform -1 0 30 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1107_
timestamp 1700315010
transform 1 0 170 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1108_
timestamp 1700315010
transform 1 0 850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1109_
timestamp 1700315010
transform -1 0 330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1110_
timestamp 1700315010
transform -1 0 190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1111_
timestamp 1700315010
transform -1 0 30 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1112_
timestamp 1700315010
transform -1 0 2010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1113_
timestamp 1700315010
transform 1 0 450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1114_
timestamp 1700315010
transform -1 0 1750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1115_
timestamp 1700315010
transform -1 0 490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1116_
timestamp 1700315010
transform -1 0 610 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1117_
timestamp 1700315010
transform 1 0 730 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1118_
timestamp 1700315010
transform -1 0 330 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1119_
timestamp 1700315010
transform 1 0 470 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1120_
timestamp 1700315010
transform 1 0 450 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1121_
timestamp 1700315010
transform 1 0 870 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1122_
timestamp 1700315010
transform -1 0 730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1123_
timestamp 1700315010
transform -1 0 630 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1124_
timestamp 1700315010
transform 1 0 490 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1125_
timestamp 1700315010
transform 1 0 170 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1126_
timestamp 1700315010
transform -1 0 30 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1127_
timestamp 1700315010
transform 1 0 550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1128_
timestamp 1700315010
transform -1 0 310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1129_
timestamp 1700315010
transform -1 0 190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1130_
timestamp 1700315010
transform 1 0 330 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1131_
timestamp 1700315010
transform -1 0 330 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1132_
timestamp 1700315010
transform -1 0 790 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1133_
timestamp 1700315010
transform -1 0 30 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1134_
timestamp 1700315010
transform -1 0 190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1135_
timestamp 1700315010
transform 1 0 170 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1136_
timestamp 1700315010
transform -1 0 290 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1137_
timestamp 1700315010
transform -1 0 30 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1138_
timestamp 1700315010
transform 1 0 470 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1139_
timestamp 1700315010
transform 1 0 570 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1140_
timestamp 1700315010
transform 1 0 1770 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1141_
timestamp 1700315010
transform 1 0 2250 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1142_
timestamp 1700315010
transform 1 0 2490 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1143_
timestamp 1700315010
transform 1 0 3290 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1144_
timestamp 1700315010
transform 1 0 3630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1145_
timestamp 1700315010
transform 1 0 2990 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1146_
timestamp 1700315010
transform -1 0 3330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1147_
timestamp 1700315010
transform -1 0 2890 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1148_
timestamp 1700315010
transform 1 0 3150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1149_
timestamp 1700315010
transform -1 0 3170 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1150_
timestamp 1700315010
transform 1 0 2790 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1151_
timestamp 1700315010
transform 1 0 3310 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1152_
timestamp 1700315010
transform -1 0 3150 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1153_
timestamp 1700315010
transform 1 0 2330 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1154_
timestamp 1700315010
transform 1 0 2490 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1155_
timestamp 1700315010
transform 1 0 2630 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1156_
timestamp 1700315010
transform -1 0 2630 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1157_
timestamp 1700315010
transform -1 0 1090 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1158_
timestamp 1700315010
transform 1 0 1150 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1159_
timestamp 1700315010
transform -1 0 1710 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1160_
timestamp 1700315010
transform 1 0 430 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1161_
timestamp 1700315010
transform 1 0 730 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1162_
timestamp 1700315010
transform 1 0 1310 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1163_
timestamp 1700315010
transform 1 0 3290 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1164_
timestamp 1700315010
transform 1 0 3730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1165_
timestamp 1700315010
transform -1 0 3890 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1166_
timestamp 1700315010
transform 1 0 4130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1167_
timestamp 1700315010
transform 1 0 4270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1168_
timestamp 1700315010
transform -1 0 3450 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1169_
timestamp 1700315010
transform 1 0 3990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1170_
timestamp 1700315010
transform 1 0 3470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1171_
timestamp 1700315010
transform 1 0 4030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1172_
timestamp 1700315010
transform 1 0 3890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1173_
timestamp 1700315010
transform 1 0 4030 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1174_
timestamp 1700315010
transform 1 0 3570 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1175_
timestamp 1700315010
transform -1 0 3750 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1176_
timestamp 1700315010
transform 1 0 3630 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1177_
timestamp 1700315010
transform -1 0 2970 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1178_
timestamp 1700315010
transform -1 0 2950 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1179_
timestamp 1700315010
transform 1 0 3330 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1180_
timestamp 1700315010
transform 1 0 2090 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1181_
timestamp 1700315010
transform 1 0 3270 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1182_
timestamp 1700315010
transform -1 0 3950 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1183_
timestamp 1700315010
transform 1 0 3770 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1184_
timestamp 1700315010
transform -1 0 3630 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1185_
timestamp 1700315010
transform -1 0 3750 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1186_
timestamp 1700315010
transform 1 0 4010 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1187_
timestamp 1700315010
transform -1 0 3310 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1188_
timestamp 1700315010
transform -1 0 4430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1189_
timestamp 1700315010
transform 1 0 3730 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1190_
timestamp 1700315010
transform 1 0 3850 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1191_
timestamp 1700315010
transform -1 0 4190 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1192_
timestamp 1700315010
transform 1 0 4450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1193_
timestamp 1700315010
transform 1 0 4330 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1194_
timestamp 1700315010
transform 1 0 4190 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1195_
timestamp 1700315010
transform 1 0 4450 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1196_
timestamp 1700315010
transform 1 0 3890 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1197_
timestamp 1700315010
transform -1 0 4070 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1198_
timestamp 1700315010
transform 1 0 3090 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1199_
timestamp 1700315010
transform 1 0 2770 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1200_
timestamp 1700315010
transform 1 0 3470 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1201_
timestamp 1700315010
transform -1 0 3750 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1202_
timestamp 1700315010
transform 1 0 4030 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1203_
timestamp 1700315010
transform 1 0 3510 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1204_
timestamp 1700315010
transform -1 0 3690 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1205_
timestamp 1700315010
transform 1 0 2650 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1206_
timestamp 1700315010
transform -1 0 30 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1207_
timestamp 1700315010
transform 1 0 750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1208_
timestamp 1700315010
transform -1 0 30 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1209_
timestamp 1700315010
transform 1 0 2350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1210_
timestamp 1700315010
transform -1 0 1530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1211_
timestamp 1700315010
transform -1 0 2150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1212_
timestamp 1700315010
transform 1 0 1810 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1213_
timestamp 1700315010
transform 1 0 2070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1214_
timestamp 1700315010
transform 1 0 2190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1215_
timestamp 1700315010
transform -1 0 1370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1216_
timestamp 1700315010
transform -1 0 1950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1217_
timestamp 1700315010
transform 1 0 1970 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1218_
timestamp 1700315010
transform -1 0 1790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1219_
timestamp 1700315010
transform 1 0 1210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1220_
timestamp 1700315010
transform -1 0 190 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1221_
timestamp 1700315010
transform -1 0 1510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1222_
timestamp 1700315010
transform -1 0 1890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1223_
timestamp 1700315010
transform 1 0 1770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1224_
timestamp 1700315010
transform -1 0 2090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1225_
timestamp 1700315010
transform 1 0 1910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1226_
timestamp 1700315010
transform -1 0 1650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1227_
timestamp 1700315010
transform 1 0 1550 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1228_
timestamp 1700315010
transform 1 0 1950 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1229_
timestamp 1700315010
transform 1 0 2210 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1230_
timestamp 1700315010
transform 1 0 1830 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1231_
timestamp 1700315010
transform -1 0 1690 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1232_
timestamp 1700315010
transform 1 0 750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1233_
timestamp 1700315010
transform 1 0 290 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1234_
timestamp 1700315010
transform 1 0 1090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1235_
timestamp 1700315010
transform 1 0 910 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1236_
timestamp 1700315010
transform -1 0 270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1237_
timestamp 1700315010
transform 1 0 550 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1238_
timestamp 1700315010
transform 1 0 730 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1239_
timestamp 1700315010
transform -1 0 490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1240_
timestamp 1700315010
transform -1 0 410 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1241_
timestamp 1700315010
transform -1 0 210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1242_
timestamp 1700315010
transform 1 0 610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1243_
timestamp 1700315010
transform 1 0 330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1244_
timestamp 1700315010
transform 1 0 170 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1245_
timestamp 1700315010
transform -1 0 190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1246_
timestamp 1700315010
transform -1 0 30 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1247_
timestamp 1700315010
transform -1 0 30 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1248_
timestamp 1700315010
transform 1 0 550 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1249_
timestamp 1700315010
transform 1 0 10 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1250_
timestamp 1700315010
transform -1 0 190 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1251_
timestamp 1700315010
transform -1 0 1090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1252_
timestamp 1700315010
transform 1 0 450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1253_
timestamp 1700315010
transform 1 0 10 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1254_
timestamp 1700315010
transform -1 0 630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1255_
timestamp 1700315010
transform -1 0 30 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1256_
timestamp 1700315010
transform 1 0 310 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1257_
timestamp 1700315010
transform -1 0 930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1258_
timestamp 1700315010
transform 1 0 330 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1259_
timestamp 1700315010
transform -1 0 810 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1260_
timestamp 1700315010
transform -1 0 810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1261_
timestamp 1700315010
transform 1 0 930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1262_
timestamp 1700315010
transform 1 0 170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1263_
timestamp 1700315010
transform -1 0 670 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1264_
timestamp 1700315010
transform 1 0 470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1265_
timestamp 1700315010
transform -1 0 650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1266_
timestamp 1700315010
transform -1 0 630 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1267_
timestamp 1700315010
transform -1 0 350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1268_
timestamp 1700315010
transform 1 0 1050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1269_
timestamp 1700315010
transform 1 0 1210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1270_
timestamp 1700315010
transform 1 0 2330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1271_
timestamp 1700315010
transform -1 0 3070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1272_
timestamp 1700315010
transform 1 0 4970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1273_
timestamp 1700315010
transform -1 0 4730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1274_
timestamp 1700315010
transform 1 0 4130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1275_
timestamp 1700315010
transform 1 0 3930 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1276_
timestamp 1700315010
transform -1 0 4450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1277_
timestamp 1700315010
transform 1 0 4090 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1278_
timestamp 1700315010
transform 1 0 4730 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1279_
timestamp 1700315010
transform 1 0 4690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1280_
timestamp 1700315010
transform -1 0 3530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1281_
timestamp 1700315010
transform -1 0 3830 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1282_
timestamp 1700315010
transform -1 0 4050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1283_
timestamp 1700315010
transform -1 0 3670 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1284_
timestamp 1700315010
transform -1 0 1630 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1285_
timestamp 1700315010
transform -1 0 3250 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1286_
timestamp 1700315010
transform -1 0 1490 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1287_
timestamp 1700315010
transform 1 0 1870 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1288_
timestamp 1700315010
transform 1 0 2970 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1289_
timestamp 1700315010
transform 1 0 2810 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1290_
timestamp 1700315010
transform -1 0 3130 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1291_
timestamp 1700315010
transform -1 0 2370 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1292_
timestamp 1700315010
transform -1 0 2230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1293_
timestamp 1700315010
transform -1 0 2610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1294_
timestamp 1700315010
transform 1 0 1230 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1295_
timestamp 1700315010
transform 1 0 1090 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1296_
timestamp 1700315010
transform -1 0 1630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1297_
timestamp 1700315010
transform 1 0 1590 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1298_
timestamp 1700315010
transform 1 0 310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1299_
timestamp 1700315010
transform 1 0 750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1300_
timestamp 1700315010
transform -1 0 1590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1301_
timestamp 1700315010
transform 1 0 2030 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1302_
timestamp 1700315010
transform -1 0 1890 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1303_
timestamp 1700315010
transform -1 0 2050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1304_
timestamp 1700315010
transform -1 0 1730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1305_
timestamp 1700315010
transform -1 0 1390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1306_
timestamp 1700315010
transform 1 0 750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1307_
timestamp 1700315010
transform 1 0 330 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1308_
timestamp 1700315010
transform -1 0 30 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1309_
timestamp 1700315010
transform 1 0 1290 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1310_
timestamp 1700315010
transform 1 0 1590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1311_
timestamp 1700315010
transform 1 0 1070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1312_
timestamp 1700315010
transform -1 0 1730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1313_
timestamp 1700315010
transform -1 0 1330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1314_
timestamp 1700315010
transform -1 0 1210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1315_
timestamp 1700315010
transform 1 0 1270 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1316_
timestamp 1700315010
transform -1 0 750 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1317_
timestamp 1700315010
transform 1 0 930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1318_
timestamp 1700315010
transform 1 0 2750 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1319_
timestamp 1700315010
transform -1 0 2030 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1320_
timestamp 1700315010
transform -1 0 1750 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1321_
timestamp 1700315010
transform -1 0 1590 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1322_
timestamp 1700315010
transform -1 0 1130 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1323_
timestamp 1700315010
transform -1 0 1450 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1324_
timestamp 1700315010
transform -1 0 790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1325_
timestamp 1700315010
transform -1 0 990 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1326_
timestamp 1700315010
transform -1 0 650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1327_
timestamp 1700315010
transform -1 0 30 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1328_
timestamp 1700315010
transform -1 0 30 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1329_
timestamp 1700315010
transform 1 0 610 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1330_
timestamp 1700315010
transform -1 0 470 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1331_
timestamp 1700315010
transform 1 0 150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1332_
timestamp 1700315010
transform 1 0 450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1333_
timestamp 1700315010
transform 1 0 770 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1334_
timestamp 1700315010
transform 1 0 470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1335_
timestamp 1700315010
transform -1 0 30 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1336_
timestamp 1700315010
transform 1 0 450 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1337_
timestamp 1700315010
transform 1 0 1090 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1338_
timestamp 1700315010
transform 1 0 10 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1339_
timestamp 1700315010
transform 1 0 690 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1340_
timestamp 1700315010
transform 1 0 610 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1341_
timestamp 1700315010
transform 1 0 130 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1342_
timestamp 1700315010
transform -1 0 170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1343_
timestamp 1700315010
transform 1 0 290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1344_
timestamp 1700315010
transform -1 0 850 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1345_
timestamp 1700315010
transform -1 0 1470 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1346_
timestamp 1700315010
transform 1 0 870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1347_
timestamp 1700315010
transform 1 0 990 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1348_
timestamp 1700315010
transform -1 0 1330 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1349_
timestamp 1700315010
transform -1 0 1370 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1350_
timestamp 1700315010
transform 1 0 490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1351_
timestamp 1700315010
transform 1 0 950 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1352_
timestamp 1700315010
transform 1 0 1710 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1353_
timestamp 1700315010
transform -1 0 1170 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1354_
timestamp 1700315010
transform 1 0 1670 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1355_
timestamp 1700315010
transform -1 0 2130 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1356_
timestamp 1700315010
transform 1 0 3250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1357_
timestamp 1700315010
transform 1 0 3410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1358_
timestamp 1700315010
transform 1 0 3550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1359_
timestamp 1700315010
transform 1 0 4530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1360_
timestamp 1700315010
transform 1 0 4470 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1361_
timestamp 1700315010
transform -1 0 4190 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1362_
timestamp 1700315010
transform 1 0 4310 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1363_
timestamp 1700315010
transform -1 0 4030 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1364_
timestamp 1700315010
transform 1 0 3870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1365_
timestamp 1700315010
transform -1 0 4790 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1366_
timestamp 1700315010
transform -1 0 1530 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1367_
timestamp 1700315010
transform 1 0 1370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1368_
timestamp 1700315010
transform 1 0 2070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1369_
timestamp 1700315010
transform 1 0 2890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1370_
timestamp 1700315010
transform 1 0 2250 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1371_
timestamp 1700315010
transform 1 0 2470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1372_
timestamp 1700315010
transform -1 0 1250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1373_
timestamp 1700315010
transform 1 0 950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1374_
timestamp 1700315010
transform -1 0 490 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1375_
timestamp 1700315010
transform -1 0 310 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1376_
timestamp 1700315010
transform -1 0 1270 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1377_
timestamp 1700315010
transform -1 0 850 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1378_
timestamp 1700315010
transform -1 0 1150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1379_
timestamp 1700315010
transform -1 0 1010 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1380_
timestamp 1700315010
transform -1 0 1130 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1381_
timestamp 1700315010
transform -1 0 970 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1382_
timestamp 1700315010
transform -1 0 710 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1383_
timestamp 1700315010
transform -1 0 970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1384_
timestamp 1700315010
transform -1 0 1130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1385_
timestamp 1700315010
transform -1 0 810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1386_
timestamp 1700315010
transform -1 0 210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1387_
timestamp 1700315010
transform 1 0 590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1388_
timestamp 1700315010
transform 1 0 1550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1389_
timestamp 1700315010
transform -1 0 1790 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1390_
timestamp 1700315010
transform -1 0 1650 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1391_
timestamp 1700315010
transform -1 0 1470 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1392_
timestamp 1700315010
transform 1 0 2010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1393_
timestamp 1700315010
transform 1 0 1850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1394_
timestamp 1700315010
transform 1 0 1350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1395_
timestamp 1700315010
transform 1 0 390 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1396_
timestamp 1700315010
transform -1 0 550 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1397_
timestamp 1700315010
transform -1 0 30 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1398_
timestamp 1700315010
transform -1 0 310 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1399_
timestamp 1700315010
transform -1 0 650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1400_
timestamp 1700315010
transform -1 0 270 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1401_
timestamp 1700315010
transform -1 0 30 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1402_
timestamp 1700315010
transform -1 0 130 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1403_
timestamp 1700315010
transform 1 0 310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1404_
timestamp 1700315010
transform -1 0 470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1405_
timestamp 1700315010
transform 1 0 310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1406_
timestamp 1700315010
transform -1 0 30 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1407_
timestamp 1700315010
transform -1 0 30 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1408_
timestamp 1700315010
transform -1 0 350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1409_
timestamp 1700315010
transform -1 0 190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1410_
timestamp 1700315010
transform 1 0 170 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1411_
timestamp 1700315010
transform -1 0 350 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1412_
timestamp 1700315010
transform 1 0 590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1413_
timestamp 1700315010
transform -1 0 30 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1414_
timestamp 1700315010
transform -1 0 610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1415_
timestamp 1700315010
transform -1 0 1270 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1416_
timestamp 1700315010
transform 1 0 1870 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1417_
timestamp 1700315010
transform 1 0 1030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1418_
timestamp 1700315010
transform -1 0 1190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1419_
timestamp 1700315010
transform 1 0 1330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1420_
timestamp 1700315010
transform -1 0 2450 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1421_
timestamp 1700315010
transform -1 0 2430 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1422_
timestamp 1700315010
transform 1 0 2750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1423_
timestamp 1700315010
transform -1 0 2590 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1424_
timestamp 1700315010
transform 1 0 2830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1425_
timestamp 1700315010
transform -1 0 2970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1426_
timestamp 1700315010
transform 1 0 3090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1427_
timestamp 1700315010
transform 1 0 4570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1428_
timestamp 1700315010
transform -1 0 4270 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1429_
timestamp 1700315010
transform 1 0 4310 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1430_
timestamp 1700315010
transform 1 0 4470 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1431_
timestamp 1700315010
transform -1 0 4690 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1432_
timestamp 1700315010
transform 1 0 4710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1433_
timestamp 1700315010
transform -1 0 4330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1434_
timestamp 1700315010
transform 1 0 4610 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1435_
timestamp 1700315010
transform 1 0 5910 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1436_
timestamp 1700315010
transform -1 0 5750 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1437_
timestamp 1700315010
transform -1 0 3850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1438_
timestamp 1700315010
transform 1 0 2630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1439_
timestamp 1700315010
transform 1 0 1250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1440_
timestamp 1700315010
transform -1 0 1170 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1441_
timestamp 1700315010
transform 1 0 470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1442_
timestamp 1700315010
transform 1 0 1790 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1443_
timestamp 1700315010
transform -1 0 2050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1444_
timestamp 1700315010
transform -1 0 1390 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1445_
timestamp 1700315010
transform -1 0 1710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1446_
timestamp 1700315010
transform 1 0 1510 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1447_
timestamp 1700315010
transform 1 0 1650 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1448_
timestamp 1700315010
transform 1 0 1770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1449_
timestamp 1700315010
transform -1 0 1890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1450_
timestamp 1700315010
transform -1 0 1530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1451_
timestamp 1700315010
transform 1 0 1630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1452_
timestamp 1700315010
transform 1 0 1870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1453_
timestamp 1700315010
transform 1 0 2050 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1454_
timestamp 1700315010
transform 1 0 1890 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1455_
timestamp 1700315010
transform 1 0 2850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1456_
timestamp 1700315010
transform -1 0 2130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1457_
timestamp 1700315010
transform -1 0 1930 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1458_
timestamp 1700315010
transform -1 0 1590 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1459_
timestamp 1700315010
transform -1 0 450 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1460_
timestamp 1700315010
transform 1 0 1710 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1461_
timestamp 1700315010
transform 1 0 710 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1462_
timestamp 1700315010
transform -1 0 150 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1463_
timestamp 1700315010
transform -1 0 1410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1464_
timestamp 1700315010
transform -1 0 870 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1465_
timestamp 1700315010
transform -1 0 1010 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1466_
timestamp 1700315010
transform -1 0 570 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1467_
timestamp 1700315010
transform -1 0 1290 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1468_
timestamp 1700315010
transform 1 0 1410 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1469_
timestamp 1700315010
transform -1 0 1090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1470_
timestamp 1700315010
transform -1 0 870 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1471_
timestamp 1700315010
transform 1 0 750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1472_
timestamp 1700315010
transform 1 0 910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1473_
timestamp 1700315010
transform 1 0 1210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1474_
timestamp 1700315010
transform 1 0 2750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1475_
timestamp 1700315010
transform 1 0 2710 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1476_
timestamp 1700315010
transform 1 0 2950 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1477_
timestamp 1700315010
transform 1 0 3110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1478_
timestamp 1700315010
transform 1 0 3210 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1479_
timestamp 1700315010
transform 1 0 3490 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1480_
timestamp 1700315010
transform -1 0 4210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1481_
timestamp 1700315010
transform -1 0 4330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1482_
timestamp 1700315010
transform 1 0 4610 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1483_
timestamp 1700315010
transform 1 0 5350 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1484_
timestamp 1700315010
transform -1 0 5490 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1485_
timestamp 1700315010
transform 1 0 5470 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1486_
timestamp 1700315010
transform -1 0 5650 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1487_
timestamp 1700315010
transform 1 0 5790 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1488_
timestamp 1700315010
transform 1 0 2150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1489_
timestamp 1700315010
transform 1 0 2310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1490_
timestamp 1700315010
transform -1 0 2330 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1491_
timestamp 1700315010
transform -1 0 2850 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1492_
timestamp 1700315010
transform -1 0 2090 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1493_
timestamp 1700315010
transform -1 0 2230 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1494_
timestamp 1700315010
transform 1 0 2530 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1495_
timestamp 1700315010
transform 1 0 2950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1496_
timestamp 1700315010
transform 1 0 2370 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1497_
timestamp 1700315010
transform 1 0 2570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1498_
timestamp 1700315010
transform 1 0 2710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1499_
timestamp 1700315010
transform 1 0 2190 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1500_
timestamp 1700315010
transform 1 0 2410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1501_
timestamp 1700315010
transform 1 0 2690 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1502_
timestamp 1700315010
transform 1 0 2710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1503_
timestamp 1700315010
transform 1 0 2750 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1504_
timestamp 1700315010
transform 1 0 2830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1505_
timestamp 1700315010
transform -1 0 2430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1506_
timestamp 1700315010
transform -1 0 2610 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1507_
timestamp 1700315010
transform -1 0 2450 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1508_
timestamp 1700315010
transform -1 0 2190 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1509_
timestamp 1700315010
transform 1 0 2010 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1510_
timestamp 1700315010
transform -1 0 1890 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1511_
timestamp 1700315010
transform 1 0 2290 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1512_
timestamp 1700315010
transform -1 0 2690 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1513_
timestamp 1700315010
transform 1 0 3290 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1514_
timestamp 1700315010
transform -1 0 3030 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1515_
timestamp 1700315010
transform 1 0 3130 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1516_
timestamp 1700315010
transform -1 0 2510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1517_
timestamp 1700315010
transform 1 0 2850 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1518_
timestamp 1700315010
transform -1 0 3190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1519_
timestamp 1700315010
transform 1 0 2890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1520_
timestamp 1700315010
transform 1 0 3030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1521_
timestamp 1700315010
transform 1 0 2530 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1522_
timestamp 1700315010
transform 1 0 2690 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1523_
timestamp 1700315010
transform 1 0 2810 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1524_
timestamp 1700315010
transform 1 0 3270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1525_
timestamp 1700315010
transform -1 0 5450 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1526_
timestamp 1700315010
transform -1 0 4950 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1527_
timestamp 1700315010
transform 1 0 4450 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1528_
timestamp 1700315010
transform 1 0 4290 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1529_
timestamp 1700315010
transform 1 0 4550 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1530_
timestamp 1700315010
transform -1 0 4830 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1531_
timestamp 1700315010
transform -1 0 5050 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1532_
timestamp 1700315010
transform 1 0 5190 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1533_
timestamp 1700315010
transform -1 0 5330 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1534_
timestamp 1700315010
transform -1 0 5130 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1535_
timestamp 1700315010
transform -1 0 3730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1536_
timestamp 1700315010
transform 1 0 3150 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1537_
timestamp 1700315010
transform 1 0 2770 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1538_
timestamp 1700315010
transform 1 0 2550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1539_
timestamp 1700315010
transform 1 0 2270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1540_
timestamp 1700315010
transform -1 0 2610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1541_
timestamp 1700315010
transform -1 0 2770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1542_
timestamp 1700315010
transform -1 0 2450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1543_
timestamp 1700315010
transform 1 0 2610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1544_
timestamp 1700315010
transform 1 0 2410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1545_
timestamp 1700315010
transform -1 0 2450 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1546_
timestamp 1700315010
transform -1 0 2470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1547_
timestamp 1700315010
transform -1 0 2650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1548_
timestamp 1700315010
transform -1 0 3010 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1549_
timestamp 1700315010
transform -1 0 2790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1550_
timestamp 1700315010
transform 1 0 3430 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1551_
timestamp 1700315010
transform 1 0 3870 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1552_
timestamp 1700315010
transform 1 0 4150 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1553_
timestamp 1700315010
transform -1 0 5030 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1554_
timestamp 1700315010
transform 1 0 5190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1555_
timestamp 1700315010
transform 1 0 5170 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1556_
timestamp 1700315010
transform -1 0 4950 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1557_
timestamp 1700315010
transform -1 0 4830 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1558_
timestamp 1700315010
transform 1 0 2490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1559_
timestamp 1700315010
transform 1 0 3490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1560_
timestamp 1700315010
transform 1 0 3610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1561_
timestamp 1700315010
transform -1 0 2670 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1562_
timestamp 1700315010
transform 1 0 2650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1563_
timestamp 1700315010
transform 1 0 3670 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1564_
timestamp 1700315010
transform -1 0 2030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1565_
timestamp 1700315010
transform -1 0 2130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1566_
timestamp 1700315010
transform -1 0 2270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1567_
timestamp 1700315010
transform 1 0 2870 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1568_
timestamp 1700315010
transform 1 0 3290 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1569_
timestamp 1700315010
transform 1 0 3910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1570_
timestamp 1700315010
transform 1 0 3330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1571_
timestamp 1700315010
transform -1 0 3590 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1572_
timestamp 1700315010
transform 1 0 3410 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1573_
timestamp 1700315010
transform 1 0 4070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1574_
timestamp 1700315010
transform -1 0 4030 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1575_
timestamp 1700315010
transform 1 0 4290 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1576_
timestamp 1700315010
transform 1 0 4130 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1577_
timestamp 1700315010
transform 1 0 4430 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1578_
timestamp 1700315010
transform 1 0 5670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1579_
timestamp 1700315010
transform -1 0 5090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1580_
timestamp 1700315010
transform -1 0 5050 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1581_
timestamp 1700315010
transform 1 0 4850 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1582_
timestamp 1700315010
transform -1 0 4470 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1583_
timestamp 1700315010
transform -1 0 3790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1584_
timestamp 1700315010
transform 1 0 2910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1585_
timestamp 1700315010
transform 1 0 3070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1586_
timestamp 1700315010
transform 1 0 3590 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1587_
timestamp 1700315010
transform 1 0 2510 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1588_
timestamp 1700315010
transform -1 0 3830 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1589_
timestamp 1700315010
transform 1 0 4910 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1590_
timestamp 1700315010
transform 1 0 4750 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1591_
timestamp 1700315010
transform -1 0 4710 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1592_
timestamp 1700315010
transform -1 0 4310 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1593_
timestamp 1700315010
transform -1 0 4310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1594_
timestamp 1700315010
transform 1 0 4270 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1595_
timestamp 1700315010
transform 1 0 3950 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1596_
timestamp 1700315010
transform -1 0 4110 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1597_
timestamp 1700315010
transform 1 0 3970 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1598_
timestamp 1700315010
transform -1 0 4130 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1599_
timestamp 1700315010
transform -1 0 3870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1600_
timestamp 1700315010
transform -1 0 3990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1601_
timestamp 1700315010
transform 1 0 3270 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1602_
timestamp 1700315010
transform -1 0 3310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1603_
timestamp 1700315010
transform 1 0 2910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1604_
timestamp 1700315010
transform -1 0 3070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1605_
timestamp 1700315010
transform -1 0 4450 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1606_
timestamp 1700315010
transform -1 0 5130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1607_
timestamp 1700315010
transform 1 0 4390 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1608_
timestamp 1700315010
transform -1 0 4550 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1636_
timestamp 1700315010
transform -1 0 5870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1637_
timestamp 1700315010
transform 1 0 5870 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1638_
timestamp 1700315010
transform -1 0 5330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1639_
timestamp 1700315010
transform 1 0 5170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1640_
timestamp 1700315010
transform 1 0 5170 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1641_
timestamp 1700315010
transform -1 0 3730 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1642_
timestamp 1700315010
transform -1 0 3130 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1643_
timestamp 1700315010
transform -1 0 2970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1644_
timestamp 1700315010
transform -1 0 3830 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1645_
timestamp 1700315010
transform -1 0 4370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1646_
timestamp 1700315010
transform -1 0 4070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1647_
timestamp 1700315010
transform 1 0 3130 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1648_
timestamp 1700315010
transform 1 0 5750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1649_
timestamp 1700315010
transform -1 0 4250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1650_
timestamp 1700315010
transform -1 0 4410 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1651_
timestamp 1700315010
transform 1 0 4270 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1652_
timestamp 1700315010
transform -1 0 3590 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1653_
timestamp 1700315010
transform 1 0 4110 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1654_
timestamp 1700315010
transform 1 0 5770 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1655_
timestamp 1700315010
transform -1 0 5630 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1656_
timestamp 1700315010
transform 1 0 5890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1657_
timestamp 1700315010
transform 1 0 5750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1658_
timestamp 1700315010
transform 1 0 5590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1659_
timestamp 1700315010
transform -1 0 5310 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1660_
timestamp 1700315010
transform -1 0 5490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1661_
timestamp 1700315010
transform 1 0 5310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1662_
timestamp 1700315010
transform -1 0 3430 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1663_
timestamp 1700315010
transform -1 0 3270 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1664_
timestamp 1700315010
transform -1 0 3410 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1665_
timestamp 1700315010
transform -1 0 3610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1666_
timestamp 1700315010
transform -1 0 3790 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1667_
timestamp 1700315010
transform 1 0 3810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1668_
timestamp 1700315010
transform 1 0 3670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1669_
timestamp 1700315010
transform -1 0 4010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1670_
timestamp 1700315010
transform 1 0 4150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1671_
timestamp 1700315010
transform 1 0 5190 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1672_
timestamp 1700315010
transform -1 0 5630 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1673_
timestamp 1700315010
transform 1 0 5450 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1674_
timestamp 1700315010
transform -1 0 5330 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1675_
timestamp 1700315010
transform -1 0 5510 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1676_
timestamp 1700315010
transform 1 0 5450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1677_
timestamp 1700315010
transform -1 0 4850 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1678_
timestamp 1700315010
transform -1 0 4890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1679_
timestamp 1700315010
transform -1 0 4490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1680_
timestamp 1700315010
transform 1 0 4590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1681_
timestamp 1700315010
transform -1 0 3970 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1682_
timestamp 1700315010
transform 1 0 4550 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1683_
timestamp 1700315010
transform 1 0 4670 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1684_
timestamp 1700315010
transform 1 0 4990 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1685_
timestamp 1700315010
transform -1 0 4150 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1686_
timestamp 1700315010
transform 1 0 4270 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1687_
timestamp 1700315010
transform -1 0 5070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1688_
timestamp 1700315010
transform 1 0 5190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1689_
timestamp 1700315010
transform 1 0 4850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1690_
timestamp 1700315010
transform 1 0 5050 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1691_
timestamp 1700315010
transform -1 0 4910 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1692_
timestamp 1700315010
transform 1 0 3550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1693_
timestamp 1700315010
transform 1 0 3070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1694_
timestamp 1700315010
transform -1 0 3250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1695_
timestamp 1700315010
transform -1 0 2910 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1696_
timestamp 1700315010
transform -1 0 3010 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1697_
timestamp 1700315010
transform -1 0 3270 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1698_
timestamp 1700315010
transform 1 0 3410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1699_
timestamp 1700315010
transform -1 0 3850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1700_
timestamp 1700315010
transform -1 0 3870 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1701_
timestamp 1700315010
transform -1 0 3570 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1702_
timestamp 1700315010
transform 1 0 3690 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1703_
timestamp 1700315010
transform -1 0 4550 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1704_
timestamp 1700315010
transform -1 0 4770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1705_
timestamp 1700315010
transform 1 0 4010 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1706_
timestamp 1700315010
transform -1 0 4310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1707_
timestamp 1700315010
transform -1 0 4450 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1708_
timestamp 1700315010
transform 1 0 4450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1709_
timestamp 1700315010
transform -1 0 3630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1710_
timestamp 1700315010
transform -1 0 3850 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1711_
timestamp 1700315010
transform -1 0 3530 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1712_
timestamp 1700315010
transform -1 0 3670 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1713_
timestamp 1700315010
transform -1 0 3370 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1714_
timestamp 1700315010
transform 1 0 3750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1715_
timestamp 1700315010
transform -1 0 3910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1716_
timestamp 1700315010
transform 1 0 4050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1717_
timestamp 1700315010
transform -1 0 4410 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1718_
timestamp 1700315010
transform 1 0 4530 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1719_
timestamp 1700315010
transform 1 0 4690 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1720_
timestamp 1700315010
transform 1 0 4210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1721_
timestamp 1700315010
transform 1 0 4630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1722_
timestamp 1700315010
transform 1 0 4730 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1723_
timestamp 1700315010
transform 1 0 4770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1724_
timestamp 1700315010
transform -1 0 4770 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1725_
timestamp 1700315010
transform 1 0 4390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1726_
timestamp 1700315010
transform -1 0 4250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1727_
timestamp 1700315010
transform -1 0 4350 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1728_
timestamp 1700315010
transform -1 0 2990 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1729_
timestamp 1700315010
transform 1 0 3050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1730_
timestamp 1700315010
transform -1 0 3210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1731_
timestamp 1700315010
transform -1 0 3350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1732_
timestamp 1700315010
transform 1 0 3510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1733_
timestamp 1700315010
transform 1 0 3650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1734_
timestamp 1700315010
transform 1 0 4930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1735_
timestamp 1700315010
transform 1 0 4890 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1736_
timestamp 1700315010
transform -1 0 5210 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1737_
timestamp 1700315010
transform 1 0 5030 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1738_
timestamp 1700315010
transform 1 0 5070 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1739_
timestamp 1700315010
transform 1 0 4890 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1740_
timestamp 1700315010
transform -1 0 5130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1741_
timestamp 1700315010
transform 1 0 5190 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1742_
timestamp 1700315010
transform 1 0 3490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1743_
timestamp 1700315010
transform -1 0 2750 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1744_
timestamp 1700315010
transform -1 0 2910 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1745_
timestamp 1700315010
transform -1 0 3210 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1746_
timestamp 1700315010
transform 1 0 3030 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1747_
timestamp 1700315010
transform 1 0 3330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1748_
timestamp 1700315010
transform -1 0 5070 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1749_
timestamp 1700315010
transform 1 0 5190 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1750_
timestamp 1700315010
transform 1 0 5410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1751_
timestamp 1700315010
transform 1 0 5350 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1752_
timestamp 1700315010
transform -1 0 5250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1753_
timestamp 1700315010
transform 1 0 5350 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1754_
timestamp 1700315010
transform 1 0 5130 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1755_
timestamp 1700315010
transform 1 0 5350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1756_
timestamp 1700315010
transform 1 0 4810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1757_
timestamp 1700315010
transform -1 0 4370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1758_
timestamp 1700315010
transform 1 0 4210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1759_
timestamp 1700315010
transform 1 0 3970 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1760_
timestamp 1700315010
transform 1 0 4490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1761_
timestamp 1700315010
transform -1 0 4670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1762_
timestamp 1700315010
transform -1 0 5110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1763_
timestamp 1700315010
transform 1 0 5250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1764_
timestamp 1700315010
transform 1 0 5570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1765_
timestamp 1700315010
transform 1 0 5710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1766_
timestamp 1700315010
transform 1 0 5810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1767_
timestamp 1700315010
transform 1 0 4870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1768_
timestamp 1700315010
transform -1 0 4730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1769_
timestamp 1700315010
transform -1 0 4570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1770_
timestamp 1700315010
transform -1 0 4990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1771_
timestamp 1700315010
transform 1 0 5490 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1772_
timestamp 1700315010
transform 1 0 5510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1773_
timestamp 1700315010
transform -1 0 5790 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1774_
timestamp 1700315010
transform -1 0 5570 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1775_
timestamp 1700315010
transform -1 0 5690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1776_
timestamp 1700315010
transform 1 0 5690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1777_
timestamp 1700315010
transform 1 0 4910 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1778_
timestamp 1700315010
transform 1 0 4450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1779_
timestamp 1700315010
transform 1 0 4330 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1780_
timestamp 1700315010
transform 1 0 4150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1781_
timestamp 1700315010
transform 1 0 4610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1782_
timestamp 1700315010
transform 1 0 4770 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1783_
timestamp 1700315010
transform 1 0 5590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1784_
timestamp 1700315010
transform 1 0 5450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1785_
timestamp 1700315010
transform -1 0 5790 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1786_
timestamp 1700315010
transform 1 0 5930 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1787_
timestamp 1700315010
transform -1 0 5870 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1788_
timestamp 1700315010
transform 1 0 5690 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1789_
timestamp 1700315010
transform 1 0 5970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1790_
timestamp 1700315010
transform 1 0 5970 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1791_
timestamp 1700315010
transform 1 0 5950 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1792_
timestamp 1700315010
transform 1 0 4630 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1793_
timestamp 1700315010
transform 1 0 4490 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1794_
timestamp 1700315010
transform 1 0 4850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1795_
timestamp 1700315010
transform -1 0 5550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1796_
timestamp 1700315010
transform 1 0 5390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1797_
timestamp 1700315010
transform -1 0 5010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1798_
timestamp 1700315010
transform -1 0 5850 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1799_
timestamp 1700315010
transform -1 0 5850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1800_
timestamp 1700315010
transform -1 0 5830 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1801_
timestamp 1700315010
transform 1 0 5390 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1802_
timestamp 1700315010
transform 1 0 4730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1803_
timestamp 1700315010
transform 1 0 5850 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1804_
timestamp 1700315010
transform -1 0 5870 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1805_
timestamp 1700315010
transform 1 0 5970 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1806_
timestamp 1700315010
transform -1 0 5670 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1807_
timestamp 1700315010
transform 1 0 5650 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1808_
timestamp 1700315010
transform 1 0 5510 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1809_
timestamp 1700315010
transform 1 0 5610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1810_
timestamp 1700315010
transform 1 0 5870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1811_
timestamp 1700315010
transform 1 0 5710 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1812_
timestamp 1700315010
transform 1 0 5950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1813_
timestamp 1700315010
transform -1 0 5970 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1814_
timestamp 1700315010
transform -1 0 5990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1815_
timestamp 1700315010
transform 1 0 5810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1816_
timestamp 1700315010
transform -1 0 5970 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1817_
timestamp 1700315010
transform -1 0 5850 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1818_
timestamp 1700315010
transform -1 0 3250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1819_
timestamp 1700315010
transform -1 0 2570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1820_
timestamp 1700315010
transform -1 0 4590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1821_
timestamp 1700315010
transform -1 0 5610 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1822_
timestamp 1700315010
transform 1 0 5450 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1823_
timestamp 1700315010
transform 1 0 5330 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1824_
timestamp 1700315010
transform 1 0 4950 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1825_
timestamp 1700315010
transform 1 0 4570 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1826_
timestamp 1700315010
transform 1 0 5730 0 -1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert0
timestamp 1700315010
transform 1 0 3910 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert1
timestamp 1700315010
transform -1 0 2190 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert2
timestamp 1700315010
transform -1 0 2310 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert3
timestamp 1700315010
transform -1 0 2250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert4
timestamp 1700315010
transform -1 0 4390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert5
timestamp 1700315010
transform -1 0 3750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert6
timestamp 1700315010
transform -1 0 2710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert7
timestamp 1700315010
transform -1 0 3390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert13
timestamp 1700315010
transform 1 0 5170 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert14
timestamp 1700315010
transform -1 0 3810 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert15
timestamp 1700315010
transform -1 0 4330 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert16
timestamp 1700315010
transform -1 0 4010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert17
timestamp 1700315010
transform 1 0 2510 0 1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert18
timestamp 1700315010
transform -1 0 2330 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert19
timestamp 1700315010
transform 1 0 3010 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert20
timestamp 1700315010
transform -1 0 2410 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert21
timestamp 1700315010
transform 1 0 5310 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert22
timestamp 1700315010
transform -1 0 4190 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert23
timestamp 1700315010
transform 1 0 4230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert24
timestamp 1700315010
transform 1 0 5270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert25
timestamp 1700315010
transform -1 0 2330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert26
timestamp 1700315010
transform -1 0 2630 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert27
timestamp 1700315010
transform -1 0 2390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert28
timestamp 1700315010
transform 1 0 3150 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert29
timestamp 1700315010
transform -1 0 2170 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert30
timestamp 1700315010
transform 1 0 3370 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert31
timestamp 1700315010
transform -1 0 2190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert32
timestamp 1700315010
transform 1 0 3490 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert33
timestamp 1700315010
transform -1 0 5070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert34
timestamp 1700315010
transform -1 0 5990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert35
timestamp 1700315010
transform -1 0 4930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert36
timestamp 1700315010
transform -1 0 5930 0 1 5470
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1700315010
transform -1 0 4530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1700315010
transform -1 0 4930 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 5790 0 1 790
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert11
timestamp 1700315010
transform -1 0 5170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 4950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__889_
timestamp 1700315010
transform 1 0 5350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__890_
timestamp 1700315010
transform -1 0 4970 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__891_
timestamp 1700315010
transform -1 0 5110 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__892_
timestamp 1700315010
transform 1 0 5370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__893_
timestamp 1700315010
transform -1 0 5230 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__894_
timestamp 1700315010
transform 1 0 5490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__895_
timestamp 1700315010
transform -1 0 5250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__896_
timestamp 1700315010
transform -1 0 5110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__897_
timestamp 1700315010
transform 1 0 5110 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__898_
timestamp 1700315010
transform -1 0 5490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__899_
timestamp 1700315010
transform 1 0 5250 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__900_
timestamp 1700315010
transform -1 0 5850 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__901_
timestamp 1700315010
transform -1 0 5710 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__902_
timestamp 1700315010
transform 1 0 5790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__903_
timestamp 1700315010
transform 1 0 4890 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__904_
timestamp 1700315010
transform -1 0 5350 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__905_
timestamp 1700315010
transform -1 0 5690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__906_
timestamp 1700315010
transform -1 0 4210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__907_
timestamp 1700315010
transform 1 0 4990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__908_
timestamp 1700315010
transform 1 0 5950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__909_
timestamp 1700315010
transform 1 0 5590 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__910_
timestamp 1700315010
transform 1 0 5530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__911_
timestamp 1700315010
transform 1 0 5410 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__912_
timestamp 1700315010
transform 1 0 5750 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__913_
timestamp 1700315010
transform -1 0 5570 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__914_
timestamp 1700315010
transform -1 0 5250 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__915_
timestamp 1700315010
transform 1 0 5230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__916_
timestamp 1700315010
transform -1 0 5630 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__917_
timestamp 1700315010
transform 1 0 5830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__918_
timestamp 1700315010
transform -1 0 5390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__919_
timestamp 1700315010
transform 1 0 5390 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__920_
timestamp 1700315010
transform -1 0 5570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__921_
timestamp 1700315010
transform 1 0 5650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__922_
timestamp 1700315010
transform 1 0 5370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__923_
timestamp 1700315010
transform 1 0 5910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__924_
timestamp 1700315010
transform 1 0 5890 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__925_
timestamp 1700315010
transform -1 0 5970 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__926_
timestamp 1700315010
transform -1 0 4330 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__927_
timestamp 1700315010
transform 1 0 4850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__928_
timestamp 1700315010
transform 1 0 4690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__929_
timestamp 1700315010
transform 1 0 4210 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__930_
timestamp 1700315010
transform 1 0 3670 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__931_
timestamp 1700315010
transform -1 0 3830 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__932_
timestamp 1700315010
transform 1 0 4130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__933_
timestamp 1700315010
transform -1 0 4410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__934_
timestamp 1700315010
transform 1 0 4530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__935_
timestamp 1700315010
transform -1 0 5390 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__936_
timestamp 1700315010
transform 1 0 4070 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__937_
timestamp 1700315010
transform -1 0 3990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__938_
timestamp 1700315010
transform -1 0 3990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__939_
timestamp 1700315010
transform 1 0 3650 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__940_
timestamp 1700315010
transform 1 0 3450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__941_
timestamp 1700315010
transform -1 0 3250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__942_
timestamp 1700315010
transform 1 0 3630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__943_
timestamp 1700315010
transform 1 0 3470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__944_
timestamp 1700315010
transform -1 0 5310 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__945_
timestamp 1700315010
transform 1 0 5570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__946_
timestamp 1700315010
transform 1 0 5410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__947_
timestamp 1700315010
transform 1 0 5650 0 1 790
box -12 -8 32 272
use FILL  FILL_1__948_
timestamp 1700315010
transform 1 0 5250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__949_
timestamp 1700315010
transform 1 0 5090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__950_
timestamp 1700315010
transform -1 0 4650 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__951_
timestamp 1700315010
transform 1 0 3910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__952_
timestamp 1700315010
transform 1 0 2330 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__953_
timestamp 1700315010
transform 1 0 2630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__954_
timestamp 1700315010
transform -1 0 2490 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__955_
timestamp 1700315010
transform 1 0 2750 0 1 790
box -12 -8 32 272
use FILL  FILL_1__956_
timestamp 1700315010
transform 1 0 3170 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__957_
timestamp 1700315010
transform 1 0 3490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__958_
timestamp 1700315010
transform 1 0 3610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__959_
timestamp 1700315010
transform 1 0 3610 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__960_
timestamp 1700315010
transform 1 0 3170 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__961_
timestamp 1700315010
transform -1 0 3470 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__962_
timestamp 1700315010
transform 1 0 3770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__963_
timestamp 1700315010
transform 1 0 2910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__964_
timestamp 1700315010
transform -1 0 2650 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__965_
timestamp 1700315010
transform 1 0 2490 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__966_
timestamp 1700315010
transform 1 0 3330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__967_
timestamp 1700315010
transform -1 0 2930 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__968_
timestamp 1700315010
transform 1 0 2570 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__969_
timestamp 1700315010
transform -1 0 2770 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__970_
timestamp 1700315010
transform 1 0 3030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__971_
timestamp 1700315010
transform 1 0 3030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__972_
timestamp 1700315010
transform -1 0 3190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__973_
timestamp 1700315010
transform 1 0 3030 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__974_
timestamp 1700315010
transform -1 0 3490 0 1 790
box -12 -8 32 272
use FILL  FILL_1__975_
timestamp 1700315010
transform 1 0 3050 0 1 790
box -12 -8 32 272
use FILL  FILL_1__976_
timestamp 1700315010
transform 1 0 2610 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__977_
timestamp 1700315010
transform 1 0 2110 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__978_
timestamp 1700315010
transform 1 0 2490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__979_
timestamp 1700315010
transform 1 0 2090 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__980_
timestamp 1700315010
transform 1 0 2890 0 1 790
box -12 -8 32 272
use FILL  FILL_1__981_
timestamp 1700315010
transform 1 0 3630 0 1 790
box -12 -8 32 272
use FILL  FILL_1__982_
timestamp 1700315010
transform -1 0 3470 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__983_
timestamp 1700315010
transform -1 0 2750 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__984_
timestamp 1700315010
transform -1 0 2430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__985_
timestamp 1700315010
transform -1 0 2350 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__986_
timestamp 1700315010
transform -1 0 1730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__987_
timestamp 1700315010
transform -1 0 1590 0 1 790
box -12 -8 32 272
use FILL  FILL_1__988_
timestamp 1700315010
transform -1 0 1370 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__989_
timestamp 1700315010
transform -1 0 1810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__990_
timestamp 1700315010
transform 1 0 1850 0 1 790
box -12 -8 32 272
use FILL  FILL_1__991_
timestamp 1700315010
transform 1 0 2390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__992_
timestamp 1700315010
transform -1 0 2390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__993_
timestamp 1700315010
transform 1 0 2010 0 1 790
box -12 -8 32 272
use FILL  FILL_1__994_
timestamp 1700315010
transform 1 0 2590 0 1 790
box -12 -8 32 272
use FILL  FILL_1__995_
timestamp 1700315010
transform -1 0 2790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__996_
timestamp 1700315010
transform 1 0 1690 0 1 790
box -12 -8 32 272
use FILL  FILL_1__997_
timestamp 1700315010
transform -1 0 1430 0 1 790
box -12 -8 32 272
use FILL  FILL_1__998_
timestamp 1700315010
transform 1 0 1610 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__999_
timestamp 1700315010
transform 1 0 2190 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1000_
timestamp 1700315010
transform 1 0 2230 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1001_
timestamp 1700315010
transform 1 0 2770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1002_
timestamp 1700315010
transform 1 0 2330 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1003_
timestamp 1700315010
transform -1 0 2950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1004_
timestamp 1700315010
transform 1 0 2470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1005_
timestamp 1700315010
transform -1 0 2330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1006_
timestamp 1700315010
transform 1 0 2030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1007_
timestamp 1700315010
transform -1 0 1670 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1008_
timestamp 1700315010
transform 1 0 1770 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1009_
timestamp 1700315010
transform -1 0 1950 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1010_
timestamp 1700315010
transform 1 0 2310 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1011_
timestamp 1700315010
transform -1 0 2210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1012_
timestamp 1700315010
transform -1 0 1470 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1013_
timestamp 1700315010
transform -1 0 2470 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1014_
timestamp 1700315010
transform -1 0 2190 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1015_
timestamp 1700315010
transform -1 0 2050 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1016_
timestamp 1700315010
transform -1 0 2070 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1017_
timestamp 1700315010
transform 1 0 2190 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1018_
timestamp 1700315010
transform -1 0 2370 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1019_
timestamp 1700315010
transform -1 0 1770 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1020_
timestamp 1700315010
transform -1 0 1510 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1021_
timestamp 1700315010
transform -1 0 1430 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1022_
timestamp 1700315010
transform -1 0 1390 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1023_
timestamp 1700315010
transform 1 0 1130 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1024_
timestamp 1700315010
transform 1 0 1490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1025_
timestamp 1700315010
transform 1 0 1450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1026_
timestamp 1700315010
transform 1 0 1250 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1027_
timestamp 1700315010
transform 1 0 1490 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1028_
timestamp 1700315010
transform 1 0 1050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1029_
timestamp 1700315010
transform -1 0 910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1030_
timestamp 1700315010
transform -1 0 1590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1031_
timestamp 1700315010
transform 1 0 1290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1032_
timestamp 1700315010
transform -1 0 1230 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1033_
timestamp 1700315010
transform -1 0 1070 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1034_
timestamp 1700315010
transform -1 0 1650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1035_
timestamp 1700315010
transform -1 0 1090 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1036_
timestamp 1700315010
transform -1 0 1170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1037_
timestamp 1700315010
transform -1 0 1050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1038_
timestamp 1700315010
transform 1 0 1630 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1039_
timestamp 1700315010
transform -1 0 1330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1040_
timestamp 1700315010
transform -1 0 2050 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1041_
timestamp 1700315010
transform -1 0 2650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1042_
timestamp 1700315010
transform 1 0 1890 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1043_
timestamp 1700315010
transform 1 0 2290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1044_
timestamp 1700315010
transform 1 0 2250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1045_
timestamp 1700315010
transform 1 0 2090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1046_
timestamp 1700315010
transform -1 0 1610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1047_
timestamp 1700315010
transform 1 0 1750 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1048_
timestamp 1700315010
transform -1 0 1950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1049_
timestamp 1700315010
transform -1 0 1450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1050_
timestamp 1700315010
transform 1 0 1490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1051_
timestamp 1700315010
transform -1 0 690 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1052_
timestamp 1700315010
transform 1 0 1190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1053_
timestamp 1700315010
transform 1 0 1210 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1054_
timestamp 1700315010
transform -1 0 1370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1055_
timestamp 1700315010
transform -1 0 950 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1056_
timestamp 1700315010
transform 1 0 990 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1057_
timestamp 1700315010
transform -1 0 1910 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1058_
timestamp 1700315010
transform 1 0 1250 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1059_
timestamp 1700315010
transform 1 0 1090 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1060_
timestamp 1700315010
transform -1 0 1170 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1061_
timestamp 1700315010
transform -1 0 2930 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1062_
timestamp 1700315010
transform -1 0 1910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1063_
timestamp 1700315010
transform 1 0 2170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1064_
timestamp 1700315010
transform 1 0 1370 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1065_
timestamp 1700315010
transform -1 0 930 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1066_
timestamp 1700315010
transform 1 0 1030 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1067_
timestamp 1700315010
transform 1 0 1290 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1068_
timestamp 1700315010
transform -1 0 850 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1069_
timestamp 1700315010
transform 1 0 1230 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1070_
timestamp 1700315010
transform 1 0 1950 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1071_
timestamp 1700315010
transform 1 0 1570 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1072_
timestamp 1700315010
transform -1 0 210 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1073_
timestamp 1700315010
transform -1 0 950 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1074_
timestamp 1700315010
transform -1 0 790 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1075_
timestamp 1700315010
transform -1 0 790 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1076_
timestamp 1700315010
transform -1 0 970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1077_
timestamp 1700315010
transform 1 0 1110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1078_
timestamp 1700315010
transform -1 0 490 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1079_
timestamp 1700315010
transform -1 0 890 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1080_
timestamp 1700315010
transform -1 0 850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1081_
timestamp 1700315010
transform -1 0 210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1082_
timestamp 1700315010
transform -1 0 1030 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1083_
timestamp 1700315010
transform -1 0 750 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1084_
timestamp 1700315010
transform -1 0 370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1085_
timestamp 1700315010
transform -1 0 350 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1086_
timestamp 1700315010
transform 1 0 670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1087_
timestamp 1700315010
transform 1 0 510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1088_
timestamp 1700315010
transform -1 0 630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1089_
timestamp 1700315010
transform 1 0 1950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1090_
timestamp 1700315010
transform 1 0 1550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1091_
timestamp 1700315010
transform -1 0 1890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1092_
timestamp 1700315010
transform -1 0 2030 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1093_
timestamp 1700315010
transform 1 0 1870 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1094_
timestamp 1700315010
transform 1 0 2170 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1095_
timestamp 1700315010
transform -1 0 1850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1096_
timestamp 1700315010
transform -1 0 1690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1097_
timestamp 1700315010
transform -1 0 1590 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1098_
timestamp 1700315010
transform -1 0 1730 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1099_
timestamp 1700315010
transform -1 0 1430 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1100_
timestamp 1700315010
transform -1 0 50 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1101_
timestamp 1700315010
transform -1 0 50 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1102_
timestamp 1700315010
transform -1 0 930 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1103_
timestamp 1700315010
transform 1 0 610 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1104_
timestamp 1700315010
transform 1 0 470 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1105_
timestamp 1700315010
transform 1 0 170 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1106_
timestamp 1700315010
transform -1 0 50 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1107_
timestamp 1700315010
transform 1 0 190 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1108_
timestamp 1700315010
transform 1 0 870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1109_
timestamp 1700315010
transform -1 0 350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1110_
timestamp 1700315010
transform -1 0 210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1111_
timestamp 1700315010
transform -1 0 50 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1112_
timestamp 1700315010
transform -1 0 2030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1113_
timestamp 1700315010
transform 1 0 470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1114_
timestamp 1700315010
transform -1 0 1770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1115_
timestamp 1700315010
transform -1 0 510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1116_
timestamp 1700315010
transform -1 0 630 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1117_
timestamp 1700315010
transform 1 0 750 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1118_
timestamp 1700315010
transform -1 0 350 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1119_
timestamp 1700315010
transform 1 0 490 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1120_
timestamp 1700315010
transform 1 0 470 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1121_
timestamp 1700315010
transform 1 0 890 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1122_
timestamp 1700315010
transform -1 0 750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1123_
timestamp 1700315010
transform -1 0 650 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1124_
timestamp 1700315010
transform 1 0 510 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1125_
timestamp 1700315010
transform 1 0 190 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1126_
timestamp 1700315010
transform -1 0 50 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1127_
timestamp 1700315010
transform 1 0 570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1128_
timestamp 1700315010
transform -1 0 330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1129_
timestamp 1700315010
transform -1 0 210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1130_
timestamp 1700315010
transform 1 0 350 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1131_
timestamp 1700315010
transform -1 0 350 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1132_
timestamp 1700315010
transform -1 0 810 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1133_
timestamp 1700315010
transform -1 0 50 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1134_
timestamp 1700315010
transform -1 0 210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1135_
timestamp 1700315010
transform 1 0 190 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1136_
timestamp 1700315010
transform -1 0 310 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1137_
timestamp 1700315010
transform -1 0 50 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1138_
timestamp 1700315010
transform 1 0 490 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1139_
timestamp 1700315010
transform 1 0 590 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1140_
timestamp 1700315010
transform 1 0 1790 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1141_
timestamp 1700315010
transform 1 0 2270 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1142_
timestamp 1700315010
transform 1 0 2510 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1143_
timestamp 1700315010
transform 1 0 3310 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1144_
timestamp 1700315010
transform 1 0 3650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1145_
timestamp 1700315010
transform 1 0 3010 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1146_
timestamp 1700315010
transform -1 0 3350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1147_
timestamp 1700315010
transform -1 0 2910 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1148_
timestamp 1700315010
transform 1 0 3170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1149_
timestamp 1700315010
transform -1 0 3190 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1150_
timestamp 1700315010
transform 1 0 2810 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1151_
timestamp 1700315010
transform 1 0 3330 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1152_
timestamp 1700315010
transform -1 0 3170 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1153_
timestamp 1700315010
transform 1 0 2350 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1154_
timestamp 1700315010
transform 1 0 2510 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1155_
timestamp 1700315010
transform 1 0 2650 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1156_
timestamp 1700315010
transform -1 0 2650 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1157_
timestamp 1700315010
transform -1 0 1110 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1158_
timestamp 1700315010
transform 1 0 1170 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1159_
timestamp 1700315010
transform -1 0 1730 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1160_
timestamp 1700315010
transform 1 0 450 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1161_
timestamp 1700315010
transform 1 0 750 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1162_
timestamp 1700315010
transform 1 0 1330 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1163_
timestamp 1700315010
transform 1 0 3310 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1164_
timestamp 1700315010
transform 1 0 3750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1165_
timestamp 1700315010
transform -1 0 3910 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1166_
timestamp 1700315010
transform 1 0 4150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1167_
timestamp 1700315010
transform 1 0 4290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1168_
timestamp 1700315010
transform -1 0 3470 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1169_
timestamp 1700315010
transform 1 0 4010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1170_
timestamp 1700315010
transform 1 0 3490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1171_
timestamp 1700315010
transform 1 0 4050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1172_
timestamp 1700315010
transform 1 0 3910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1173_
timestamp 1700315010
transform 1 0 4050 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1174_
timestamp 1700315010
transform 1 0 3590 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1175_
timestamp 1700315010
transform -1 0 3770 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1176_
timestamp 1700315010
transform 1 0 3650 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1177_
timestamp 1700315010
transform -1 0 2990 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1178_
timestamp 1700315010
transform -1 0 2970 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1179_
timestamp 1700315010
transform 1 0 3350 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1180_
timestamp 1700315010
transform 1 0 2110 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1181_
timestamp 1700315010
transform 1 0 3290 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1182_
timestamp 1700315010
transform -1 0 3970 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1183_
timestamp 1700315010
transform 1 0 3790 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1184_
timestamp 1700315010
transform -1 0 3650 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1185_
timestamp 1700315010
transform -1 0 3770 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1186_
timestamp 1700315010
transform 1 0 4030 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1187_
timestamp 1700315010
transform -1 0 3330 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1188_
timestamp 1700315010
transform -1 0 4450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1189_
timestamp 1700315010
transform 1 0 3750 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1190_
timestamp 1700315010
transform 1 0 3870 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1191_
timestamp 1700315010
transform -1 0 4210 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1192_
timestamp 1700315010
transform 1 0 4470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1193_
timestamp 1700315010
transform 1 0 4350 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1194_
timestamp 1700315010
transform 1 0 4210 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1195_
timestamp 1700315010
transform 1 0 4470 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1196_
timestamp 1700315010
transform 1 0 3910 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1197_
timestamp 1700315010
transform -1 0 4090 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1198_
timestamp 1700315010
transform 1 0 3110 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1199_
timestamp 1700315010
transform 1 0 2790 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1200_
timestamp 1700315010
transform 1 0 3490 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1201_
timestamp 1700315010
transform -1 0 3770 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1202_
timestamp 1700315010
transform 1 0 4050 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1203_
timestamp 1700315010
transform 1 0 3530 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1204_
timestamp 1700315010
transform -1 0 3710 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1205_
timestamp 1700315010
transform 1 0 2670 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1206_
timestamp 1700315010
transform -1 0 50 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1207_
timestamp 1700315010
transform 1 0 770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1208_
timestamp 1700315010
transform -1 0 50 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1209_
timestamp 1700315010
transform 1 0 2370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1210_
timestamp 1700315010
transform -1 0 1550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1211_
timestamp 1700315010
transform -1 0 2170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1212_
timestamp 1700315010
transform 1 0 1830 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1213_
timestamp 1700315010
transform 1 0 2090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1214_
timestamp 1700315010
transform 1 0 2210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1215_
timestamp 1700315010
transform -1 0 1390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1216_
timestamp 1700315010
transform -1 0 1970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1217_
timestamp 1700315010
transform 1 0 1990 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1218_
timestamp 1700315010
transform -1 0 1810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1219_
timestamp 1700315010
transform 1 0 1230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1220_
timestamp 1700315010
transform -1 0 210 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1221_
timestamp 1700315010
transform -1 0 1530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1222_
timestamp 1700315010
transform -1 0 1910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1223_
timestamp 1700315010
transform 1 0 1790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1224_
timestamp 1700315010
transform -1 0 2110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1225_
timestamp 1700315010
transform 1 0 1930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1226_
timestamp 1700315010
transform -1 0 1670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1227_
timestamp 1700315010
transform 1 0 1570 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1228_
timestamp 1700315010
transform 1 0 1970 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1229_
timestamp 1700315010
transform 1 0 2230 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1230_
timestamp 1700315010
transform 1 0 1850 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1231_
timestamp 1700315010
transform -1 0 1710 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1232_
timestamp 1700315010
transform 1 0 770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1233_
timestamp 1700315010
transform 1 0 310 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1234_
timestamp 1700315010
transform 1 0 1110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1235_
timestamp 1700315010
transform 1 0 930 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1236_
timestamp 1700315010
transform -1 0 290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1237_
timestamp 1700315010
transform 1 0 570 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1238_
timestamp 1700315010
transform 1 0 750 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1239_
timestamp 1700315010
transform -1 0 510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1240_
timestamp 1700315010
transform -1 0 430 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1241_
timestamp 1700315010
transform -1 0 230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1242_
timestamp 1700315010
transform 1 0 630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1243_
timestamp 1700315010
transform 1 0 350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1244_
timestamp 1700315010
transform 1 0 190 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1245_
timestamp 1700315010
transform -1 0 210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1246_
timestamp 1700315010
transform -1 0 50 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1247_
timestamp 1700315010
transform -1 0 50 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1248_
timestamp 1700315010
transform 1 0 570 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1249_
timestamp 1700315010
transform 1 0 30 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1250_
timestamp 1700315010
transform -1 0 210 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1251_
timestamp 1700315010
transform -1 0 1110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1252_
timestamp 1700315010
transform 1 0 470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1253_
timestamp 1700315010
transform 1 0 30 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1254_
timestamp 1700315010
transform -1 0 650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1255_
timestamp 1700315010
transform -1 0 50 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1256_
timestamp 1700315010
transform 1 0 330 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1257_
timestamp 1700315010
transform -1 0 950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1258_
timestamp 1700315010
transform 1 0 350 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1259_
timestamp 1700315010
transform -1 0 830 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1260_
timestamp 1700315010
transform -1 0 830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1261_
timestamp 1700315010
transform 1 0 950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1262_
timestamp 1700315010
transform 1 0 190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1263_
timestamp 1700315010
transform -1 0 690 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1264_
timestamp 1700315010
transform 1 0 490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1265_
timestamp 1700315010
transform -1 0 670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1266_
timestamp 1700315010
transform -1 0 650 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1267_
timestamp 1700315010
transform -1 0 370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1268_
timestamp 1700315010
transform 1 0 1070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1269_
timestamp 1700315010
transform 1 0 1230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1270_
timestamp 1700315010
transform 1 0 2350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1271_
timestamp 1700315010
transform -1 0 3090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1272_
timestamp 1700315010
transform 1 0 4990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1273_
timestamp 1700315010
transform -1 0 4750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1274_
timestamp 1700315010
transform 1 0 4150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1275_
timestamp 1700315010
transform 1 0 3950 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1276_
timestamp 1700315010
transform -1 0 4470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1277_
timestamp 1700315010
transform 1 0 4110 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1278_
timestamp 1700315010
transform 1 0 4750 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1279_
timestamp 1700315010
transform 1 0 4710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1280_
timestamp 1700315010
transform -1 0 3550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1281_
timestamp 1700315010
transform -1 0 3850 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1282_
timestamp 1700315010
transform -1 0 4070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1283_
timestamp 1700315010
transform -1 0 3690 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1284_
timestamp 1700315010
transform -1 0 1650 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1285_
timestamp 1700315010
transform -1 0 3270 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1286_
timestamp 1700315010
transform -1 0 1510 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1287_
timestamp 1700315010
transform 1 0 1890 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1288_
timestamp 1700315010
transform 1 0 2990 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1289_
timestamp 1700315010
transform 1 0 2830 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1290_
timestamp 1700315010
transform -1 0 3150 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1291_
timestamp 1700315010
transform -1 0 2390 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1292_
timestamp 1700315010
transform -1 0 2250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1293_
timestamp 1700315010
transform -1 0 2630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1294_
timestamp 1700315010
transform 1 0 1250 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1295_
timestamp 1700315010
transform 1 0 1110 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1296_
timestamp 1700315010
transform -1 0 1650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1297_
timestamp 1700315010
transform 1 0 1610 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1298_
timestamp 1700315010
transform 1 0 330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1299_
timestamp 1700315010
transform 1 0 770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1300_
timestamp 1700315010
transform -1 0 1610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1301_
timestamp 1700315010
transform 1 0 2050 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1302_
timestamp 1700315010
transform -1 0 1910 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1303_
timestamp 1700315010
transform -1 0 2070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1304_
timestamp 1700315010
transform -1 0 1750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1305_
timestamp 1700315010
transform -1 0 1410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1306_
timestamp 1700315010
transform 1 0 770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1307_
timestamp 1700315010
transform 1 0 350 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1308_
timestamp 1700315010
transform -1 0 50 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1309_
timestamp 1700315010
transform 1 0 1310 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1310_
timestamp 1700315010
transform 1 0 1610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1311_
timestamp 1700315010
transform 1 0 1090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1312_
timestamp 1700315010
transform -1 0 1750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1313_
timestamp 1700315010
transform -1 0 1350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1314_
timestamp 1700315010
transform -1 0 1230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1315_
timestamp 1700315010
transform 1 0 1290 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1316_
timestamp 1700315010
transform -1 0 770 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1317_
timestamp 1700315010
transform 1 0 950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1318_
timestamp 1700315010
transform 1 0 2770 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1319_
timestamp 1700315010
transform -1 0 2050 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1320_
timestamp 1700315010
transform -1 0 1770 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1321_
timestamp 1700315010
transform -1 0 1610 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1322_
timestamp 1700315010
transform -1 0 1150 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1323_
timestamp 1700315010
transform -1 0 1470 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1324_
timestamp 1700315010
transform -1 0 810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1325_
timestamp 1700315010
transform -1 0 1010 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1326_
timestamp 1700315010
transform -1 0 670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1327_
timestamp 1700315010
transform -1 0 50 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1328_
timestamp 1700315010
transform -1 0 50 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1329_
timestamp 1700315010
transform 1 0 630 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1330_
timestamp 1700315010
transform -1 0 490 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1331_
timestamp 1700315010
transform 1 0 170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1332_
timestamp 1700315010
transform 1 0 470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1333_
timestamp 1700315010
transform 1 0 790 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1334_
timestamp 1700315010
transform 1 0 490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1335_
timestamp 1700315010
transform -1 0 50 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1336_
timestamp 1700315010
transform 1 0 470 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1337_
timestamp 1700315010
transform 1 0 1110 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1338_
timestamp 1700315010
transform 1 0 30 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1339_
timestamp 1700315010
transform 1 0 710 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1340_
timestamp 1700315010
transform 1 0 630 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1341_
timestamp 1700315010
transform 1 0 150 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1342_
timestamp 1700315010
transform -1 0 190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1343_
timestamp 1700315010
transform 1 0 310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1344_
timestamp 1700315010
transform -1 0 870 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1345_
timestamp 1700315010
transform -1 0 1490 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1346_
timestamp 1700315010
transform 1 0 890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1347_
timestamp 1700315010
transform 1 0 1010 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1348_
timestamp 1700315010
transform -1 0 1350 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1349_
timestamp 1700315010
transform -1 0 1390 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1350_
timestamp 1700315010
transform 1 0 510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1351_
timestamp 1700315010
transform 1 0 970 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1352_
timestamp 1700315010
transform 1 0 1730 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1353_
timestamp 1700315010
transform -1 0 1190 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1354_
timestamp 1700315010
transform 1 0 1690 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1355_
timestamp 1700315010
transform -1 0 2150 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1356_
timestamp 1700315010
transform 1 0 3270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1357_
timestamp 1700315010
transform 1 0 3430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1358_
timestamp 1700315010
transform 1 0 3570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1359_
timestamp 1700315010
transform 1 0 4550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1360_
timestamp 1700315010
transform 1 0 4490 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1361_
timestamp 1700315010
transform -1 0 4210 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1362_
timestamp 1700315010
transform 1 0 4330 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1363_
timestamp 1700315010
transform -1 0 4050 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1364_
timestamp 1700315010
transform 1 0 3890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1365_
timestamp 1700315010
transform -1 0 4810 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1366_
timestamp 1700315010
transform -1 0 1550 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1367_
timestamp 1700315010
transform 1 0 1390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1368_
timestamp 1700315010
transform 1 0 2090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1369_
timestamp 1700315010
transform 1 0 2910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1370_
timestamp 1700315010
transform 1 0 2270 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1371_
timestamp 1700315010
transform 1 0 2490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1372_
timestamp 1700315010
transform -1 0 1270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1373_
timestamp 1700315010
transform 1 0 970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1374_
timestamp 1700315010
transform -1 0 510 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1375_
timestamp 1700315010
transform -1 0 330 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1376_
timestamp 1700315010
transform -1 0 1290 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1377_
timestamp 1700315010
transform -1 0 870 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1378_
timestamp 1700315010
transform -1 0 1170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1379_
timestamp 1700315010
transform -1 0 1030 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1380_
timestamp 1700315010
transform -1 0 1150 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1381_
timestamp 1700315010
transform -1 0 990 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1382_
timestamp 1700315010
transform -1 0 730 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1383_
timestamp 1700315010
transform -1 0 990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1384_
timestamp 1700315010
transform -1 0 1150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1385_
timestamp 1700315010
transform -1 0 830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1386_
timestamp 1700315010
transform -1 0 230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1387_
timestamp 1700315010
transform 1 0 610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1388_
timestamp 1700315010
transform 1 0 1570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1389_
timestamp 1700315010
transform -1 0 1810 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1390_
timestamp 1700315010
transform -1 0 1670 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1391_
timestamp 1700315010
transform -1 0 1490 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1392_
timestamp 1700315010
transform 1 0 2030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1393_
timestamp 1700315010
transform 1 0 1870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1394_
timestamp 1700315010
transform 1 0 1370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1395_
timestamp 1700315010
transform 1 0 410 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1396_
timestamp 1700315010
transform -1 0 570 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1397_
timestamp 1700315010
transform -1 0 50 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1398_
timestamp 1700315010
transform -1 0 330 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1399_
timestamp 1700315010
transform -1 0 670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1400_
timestamp 1700315010
transform -1 0 290 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1401_
timestamp 1700315010
transform -1 0 50 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1402_
timestamp 1700315010
transform -1 0 150 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1403_
timestamp 1700315010
transform 1 0 330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1404_
timestamp 1700315010
transform -1 0 490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1405_
timestamp 1700315010
transform 1 0 330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1406_
timestamp 1700315010
transform -1 0 50 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1407_
timestamp 1700315010
transform -1 0 50 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1408_
timestamp 1700315010
transform -1 0 370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1409_
timestamp 1700315010
transform -1 0 210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1410_
timestamp 1700315010
transform 1 0 190 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1411_
timestamp 1700315010
transform -1 0 370 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1412_
timestamp 1700315010
transform 1 0 610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1413_
timestamp 1700315010
transform -1 0 50 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1414_
timestamp 1700315010
transform -1 0 630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1415_
timestamp 1700315010
transform -1 0 1290 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1416_
timestamp 1700315010
transform 1 0 1890 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1417_
timestamp 1700315010
transform 1 0 1050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1418_
timestamp 1700315010
transform -1 0 1210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1419_
timestamp 1700315010
transform 1 0 1350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1420_
timestamp 1700315010
transform -1 0 2470 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1421_
timestamp 1700315010
transform -1 0 2450 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1422_
timestamp 1700315010
transform 1 0 2770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1423_
timestamp 1700315010
transform -1 0 2610 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1424_
timestamp 1700315010
transform 1 0 2850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1425_
timestamp 1700315010
transform -1 0 2990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1426_
timestamp 1700315010
transform 1 0 3110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1427_
timestamp 1700315010
transform 1 0 4590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1428_
timestamp 1700315010
transform -1 0 4290 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1429_
timestamp 1700315010
transform 1 0 4330 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1430_
timestamp 1700315010
transform 1 0 4490 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1431_
timestamp 1700315010
transform -1 0 4710 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1432_
timestamp 1700315010
transform 1 0 4730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1433_
timestamp 1700315010
transform -1 0 4350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1434_
timestamp 1700315010
transform 1 0 4630 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1435_
timestamp 1700315010
transform 1 0 5930 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1436_
timestamp 1700315010
transform -1 0 5770 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1437_
timestamp 1700315010
transform -1 0 3870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1438_
timestamp 1700315010
transform 1 0 2650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1439_
timestamp 1700315010
transform 1 0 1270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1440_
timestamp 1700315010
transform -1 0 1190 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1441_
timestamp 1700315010
transform 1 0 490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1442_
timestamp 1700315010
transform 1 0 1810 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1443_
timestamp 1700315010
transform -1 0 2070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1444_
timestamp 1700315010
transform -1 0 1410 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1445_
timestamp 1700315010
transform -1 0 1730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1446_
timestamp 1700315010
transform 1 0 1530 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1447_
timestamp 1700315010
transform 1 0 1670 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1448_
timestamp 1700315010
transform 1 0 1790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1449_
timestamp 1700315010
transform -1 0 1910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1450_
timestamp 1700315010
transform -1 0 1550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1451_
timestamp 1700315010
transform 1 0 1650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1452_
timestamp 1700315010
transform 1 0 1890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1453_
timestamp 1700315010
transform 1 0 2070 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1454_
timestamp 1700315010
transform 1 0 1910 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1455_
timestamp 1700315010
transform 1 0 2870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1456_
timestamp 1700315010
transform -1 0 2150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1457_
timestamp 1700315010
transform -1 0 1950 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1458_
timestamp 1700315010
transform -1 0 1610 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1459_
timestamp 1700315010
transform -1 0 470 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1460_
timestamp 1700315010
transform 1 0 1730 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1461_
timestamp 1700315010
transform 1 0 730 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1462_
timestamp 1700315010
transform -1 0 170 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1463_
timestamp 1700315010
transform -1 0 1430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1464_
timestamp 1700315010
transform -1 0 890 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1465_
timestamp 1700315010
transform -1 0 1030 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1466_
timestamp 1700315010
transform -1 0 590 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1467_
timestamp 1700315010
transform -1 0 1310 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1468_
timestamp 1700315010
transform 1 0 1430 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1469_
timestamp 1700315010
transform -1 0 1110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1470_
timestamp 1700315010
transform -1 0 890 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1471_
timestamp 1700315010
transform 1 0 770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1472_
timestamp 1700315010
transform 1 0 930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1473_
timestamp 1700315010
transform 1 0 1230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1474_
timestamp 1700315010
transform 1 0 2770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1475_
timestamp 1700315010
transform 1 0 2730 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1476_
timestamp 1700315010
transform 1 0 2970 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1477_
timestamp 1700315010
transform 1 0 3130 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1478_
timestamp 1700315010
transform 1 0 3230 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1479_
timestamp 1700315010
transform 1 0 3510 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1480_
timestamp 1700315010
transform -1 0 4230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1481_
timestamp 1700315010
transform -1 0 4350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1482_
timestamp 1700315010
transform 1 0 4630 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1483_
timestamp 1700315010
transform 1 0 5370 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1484_
timestamp 1700315010
transform -1 0 5510 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1485_
timestamp 1700315010
transform 1 0 5490 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1486_
timestamp 1700315010
transform -1 0 5670 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1487_
timestamp 1700315010
transform 1 0 5810 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1488_
timestamp 1700315010
transform 1 0 2170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1489_
timestamp 1700315010
transform 1 0 2330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1490_
timestamp 1700315010
transform -1 0 2350 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1491_
timestamp 1700315010
transform -1 0 2870 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1492_
timestamp 1700315010
transform -1 0 2110 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1493_
timestamp 1700315010
transform -1 0 2250 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1494_
timestamp 1700315010
transform 1 0 2550 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1495_
timestamp 1700315010
transform 1 0 2970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1496_
timestamp 1700315010
transform 1 0 2390 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1497_
timestamp 1700315010
transform 1 0 2590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1498_
timestamp 1700315010
transform 1 0 2730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1499_
timestamp 1700315010
transform 1 0 2210 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1500_
timestamp 1700315010
transform 1 0 2430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1501_
timestamp 1700315010
transform 1 0 2710 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1502_
timestamp 1700315010
transform 1 0 2730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1503_
timestamp 1700315010
transform 1 0 2770 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1504_
timestamp 1700315010
transform 1 0 2850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1505_
timestamp 1700315010
transform -1 0 2450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1506_
timestamp 1700315010
transform -1 0 2630 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1507_
timestamp 1700315010
transform -1 0 2470 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1508_
timestamp 1700315010
transform -1 0 2210 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1509_
timestamp 1700315010
transform 1 0 2030 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1510_
timestamp 1700315010
transform -1 0 1910 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1511_
timestamp 1700315010
transform 1 0 2310 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1512_
timestamp 1700315010
transform -1 0 2710 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1513_
timestamp 1700315010
transform 1 0 3310 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1514_
timestamp 1700315010
transform -1 0 3050 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1515_
timestamp 1700315010
transform 1 0 3150 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1516_
timestamp 1700315010
transform -1 0 2530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1517_
timestamp 1700315010
transform 1 0 2870 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1518_
timestamp 1700315010
transform -1 0 3210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1519_
timestamp 1700315010
transform 1 0 2910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1520_
timestamp 1700315010
transform 1 0 3050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1521_
timestamp 1700315010
transform 1 0 2550 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1522_
timestamp 1700315010
transform 1 0 2710 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1523_
timestamp 1700315010
transform 1 0 2830 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1524_
timestamp 1700315010
transform 1 0 3290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1525_
timestamp 1700315010
transform -1 0 5470 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1526_
timestamp 1700315010
transform -1 0 4970 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1527_
timestamp 1700315010
transform 1 0 4470 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1528_
timestamp 1700315010
transform 1 0 4310 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1529_
timestamp 1700315010
transform 1 0 4570 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1530_
timestamp 1700315010
transform -1 0 4850 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1531_
timestamp 1700315010
transform -1 0 5070 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1532_
timestamp 1700315010
transform 1 0 5210 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1533_
timestamp 1700315010
transform -1 0 5350 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1534_
timestamp 1700315010
transform -1 0 5150 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1535_
timestamp 1700315010
transform -1 0 3750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1536_
timestamp 1700315010
transform 1 0 3170 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1537_
timestamp 1700315010
transform 1 0 2790 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1538_
timestamp 1700315010
transform 1 0 2570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1539_
timestamp 1700315010
transform 1 0 2290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1540_
timestamp 1700315010
transform -1 0 2630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1541_
timestamp 1700315010
transform -1 0 2790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1542_
timestamp 1700315010
transform -1 0 2470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1543_
timestamp 1700315010
transform 1 0 2630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1544_
timestamp 1700315010
transform 1 0 2430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1545_
timestamp 1700315010
transform -1 0 2470 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1546_
timestamp 1700315010
transform -1 0 2490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1547_
timestamp 1700315010
transform -1 0 2670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1548_
timestamp 1700315010
transform -1 0 3030 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1549_
timestamp 1700315010
transform -1 0 2810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1550_
timestamp 1700315010
transform 1 0 3450 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1551_
timestamp 1700315010
transform 1 0 3890 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1552_
timestamp 1700315010
transform 1 0 4170 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1553_
timestamp 1700315010
transform -1 0 5050 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1554_
timestamp 1700315010
transform 1 0 5210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1555_
timestamp 1700315010
transform 1 0 5190 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1556_
timestamp 1700315010
transform -1 0 4970 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1557_
timestamp 1700315010
transform -1 0 4850 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1558_
timestamp 1700315010
transform 1 0 2510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1559_
timestamp 1700315010
transform 1 0 3510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1560_
timestamp 1700315010
transform 1 0 3630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1561_
timestamp 1700315010
transform -1 0 2690 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1562_
timestamp 1700315010
transform 1 0 2670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1563_
timestamp 1700315010
transform 1 0 3690 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1564_
timestamp 1700315010
transform -1 0 2050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1565_
timestamp 1700315010
transform -1 0 2150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1566_
timestamp 1700315010
transform -1 0 2290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1567_
timestamp 1700315010
transform 1 0 2890 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1568_
timestamp 1700315010
transform 1 0 3310 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1569_
timestamp 1700315010
transform 1 0 3930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1570_
timestamp 1700315010
transform 1 0 3350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1571_
timestamp 1700315010
transform -1 0 3610 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1572_
timestamp 1700315010
transform 1 0 3430 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1573_
timestamp 1700315010
transform 1 0 4090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1574_
timestamp 1700315010
transform -1 0 4050 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1575_
timestamp 1700315010
transform 1 0 4310 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1576_
timestamp 1700315010
transform 1 0 4150 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1577_
timestamp 1700315010
transform 1 0 4450 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1578_
timestamp 1700315010
transform 1 0 5690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1579_
timestamp 1700315010
transform -1 0 5110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1580_
timestamp 1700315010
transform -1 0 5070 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1581_
timestamp 1700315010
transform 1 0 4870 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1582_
timestamp 1700315010
transform -1 0 4490 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1583_
timestamp 1700315010
transform -1 0 3810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1584_
timestamp 1700315010
transform 1 0 2930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1585_
timestamp 1700315010
transform 1 0 3090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1586_
timestamp 1700315010
transform 1 0 3610 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1587_
timestamp 1700315010
transform 1 0 2530 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1588_
timestamp 1700315010
transform -1 0 3850 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1589_
timestamp 1700315010
transform 1 0 4930 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1590_
timestamp 1700315010
transform 1 0 4770 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1591_
timestamp 1700315010
transform -1 0 4730 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1592_
timestamp 1700315010
transform -1 0 4330 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1593_
timestamp 1700315010
transform -1 0 4330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1594_
timestamp 1700315010
transform 1 0 4290 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1595_
timestamp 1700315010
transform 1 0 3970 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1596_
timestamp 1700315010
transform -1 0 4130 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1597_
timestamp 1700315010
transform 1 0 3990 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1598_
timestamp 1700315010
transform -1 0 4150 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1599_
timestamp 1700315010
transform -1 0 3890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1600_
timestamp 1700315010
transform -1 0 4010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1601_
timestamp 1700315010
transform 1 0 3290 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1602_
timestamp 1700315010
transform -1 0 3330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1603_
timestamp 1700315010
transform 1 0 2930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1604_
timestamp 1700315010
transform -1 0 3090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1605_
timestamp 1700315010
transform -1 0 4470 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1606_
timestamp 1700315010
transform -1 0 5150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1607_
timestamp 1700315010
transform 1 0 4410 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1608_
timestamp 1700315010
transform -1 0 4570 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1636_
timestamp 1700315010
transform -1 0 5890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1637_
timestamp 1700315010
transform 1 0 5890 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1638_
timestamp 1700315010
transform -1 0 5350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1639_
timestamp 1700315010
transform 1 0 5190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1640_
timestamp 1700315010
transform 1 0 5190 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1641_
timestamp 1700315010
transform -1 0 3750 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1642_
timestamp 1700315010
transform -1 0 3150 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1643_
timestamp 1700315010
transform -1 0 2990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1644_
timestamp 1700315010
transform -1 0 3850 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1645_
timestamp 1700315010
transform -1 0 4390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1646_
timestamp 1700315010
transform -1 0 4090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1647_
timestamp 1700315010
transform 1 0 3150 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1648_
timestamp 1700315010
transform 1 0 5770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1649_
timestamp 1700315010
transform -1 0 4270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1650_
timestamp 1700315010
transform -1 0 4430 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1651_
timestamp 1700315010
transform 1 0 4290 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1652_
timestamp 1700315010
transform -1 0 3610 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1653_
timestamp 1700315010
transform 1 0 4130 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1654_
timestamp 1700315010
transform 1 0 5790 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1655_
timestamp 1700315010
transform -1 0 5650 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1656_
timestamp 1700315010
transform 1 0 5910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1657_
timestamp 1700315010
transform 1 0 5770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1658_
timestamp 1700315010
transform 1 0 5610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1659_
timestamp 1700315010
transform -1 0 5330 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1660_
timestamp 1700315010
transform -1 0 5510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1661_
timestamp 1700315010
transform 1 0 5330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1662_
timestamp 1700315010
transform -1 0 3450 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1663_
timestamp 1700315010
transform -1 0 3290 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1664_
timestamp 1700315010
transform -1 0 3430 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1665_
timestamp 1700315010
transform -1 0 3630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1666_
timestamp 1700315010
transform -1 0 3810 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1667_
timestamp 1700315010
transform 1 0 3830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1668_
timestamp 1700315010
transform 1 0 3690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1669_
timestamp 1700315010
transform -1 0 4030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1670_
timestamp 1700315010
transform 1 0 4170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1671_
timestamp 1700315010
transform 1 0 5210 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1672_
timestamp 1700315010
transform -1 0 5650 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1673_
timestamp 1700315010
transform 1 0 5470 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1674_
timestamp 1700315010
transform -1 0 5350 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1675_
timestamp 1700315010
transform -1 0 5530 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1676_
timestamp 1700315010
transform 1 0 5470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1677_
timestamp 1700315010
transform -1 0 4870 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1678_
timestamp 1700315010
transform -1 0 4910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1679_
timestamp 1700315010
transform -1 0 4510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1680_
timestamp 1700315010
transform 1 0 4610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1681_
timestamp 1700315010
transform -1 0 3990 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1682_
timestamp 1700315010
transform 1 0 4570 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1683_
timestamp 1700315010
transform 1 0 4690 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1684_
timestamp 1700315010
transform 1 0 5010 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1685_
timestamp 1700315010
transform -1 0 4170 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1686_
timestamp 1700315010
transform 1 0 4290 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1687_
timestamp 1700315010
transform -1 0 5090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1688_
timestamp 1700315010
transform 1 0 5210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1689_
timestamp 1700315010
transform 1 0 4870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1690_
timestamp 1700315010
transform 1 0 5070 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1691_
timestamp 1700315010
transform -1 0 4930 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1692_
timestamp 1700315010
transform 1 0 3570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1693_
timestamp 1700315010
transform 1 0 3090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1694_
timestamp 1700315010
transform -1 0 3270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1695_
timestamp 1700315010
transform -1 0 2930 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1696_
timestamp 1700315010
transform -1 0 3030 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1697_
timestamp 1700315010
transform -1 0 3290 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1698_
timestamp 1700315010
transform 1 0 3430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1699_
timestamp 1700315010
transform -1 0 3870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1700_
timestamp 1700315010
transform -1 0 3890 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1701_
timestamp 1700315010
transform -1 0 3590 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1702_
timestamp 1700315010
transform 1 0 3710 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1703_
timestamp 1700315010
transform -1 0 4570 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1704_
timestamp 1700315010
transform -1 0 4790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1705_
timestamp 1700315010
transform 1 0 4030 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1706_
timestamp 1700315010
transform -1 0 4330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1707_
timestamp 1700315010
transform -1 0 4470 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1708_
timestamp 1700315010
transform 1 0 4470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1709_
timestamp 1700315010
transform -1 0 3650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1710_
timestamp 1700315010
transform -1 0 3870 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1711_
timestamp 1700315010
transform -1 0 3550 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1712_
timestamp 1700315010
transform -1 0 3690 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1713_
timestamp 1700315010
transform -1 0 3390 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1714_
timestamp 1700315010
transform 1 0 3770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1715_
timestamp 1700315010
transform -1 0 3930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1716_
timestamp 1700315010
transform 1 0 4070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1717_
timestamp 1700315010
transform -1 0 4430 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1718_
timestamp 1700315010
transform 1 0 4550 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1719_
timestamp 1700315010
transform 1 0 4710 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1720_
timestamp 1700315010
transform 1 0 4230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1721_
timestamp 1700315010
transform 1 0 4650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1722_
timestamp 1700315010
transform 1 0 4750 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1723_
timestamp 1700315010
transform 1 0 4790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1724_
timestamp 1700315010
transform -1 0 4790 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1725_
timestamp 1700315010
transform 1 0 4410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1726_
timestamp 1700315010
transform -1 0 4270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1727_
timestamp 1700315010
transform -1 0 4370 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1728_
timestamp 1700315010
transform -1 0 3010 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1729_
timestamp 1700315010
transform 1 0 3070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1730_
timestamp 1700315010
transform -1 0 3230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1731_
timestamp 1700315010
transform -1 0 3370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1732_
timestamp 1700315010
transform 1 0 3530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1733_
timestamp 1700315010
transform 1 0 3670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1734_
timestamp 1700315010
transform 1 0 4950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1735_
timestamp 1700315010
transform 1 0 4910 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1736_
timestamp 1700315010
transform -1 0 5230 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1737_
timestamp 1700315010
transform 1 0 5050 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1738_
timestamp 1700315010
transform 1 0 5090 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1739_
timestamp 1700315010
transform 1 0 4910 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1740_
timestamp 1700315010
transform -1 0 5150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1741_
timestamp 1700315010
transform 1 0 5210 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1742_
timestamp 1700315010
transform 1 0 3510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1743_
timestamp 1700315010
transform -1 0 2770 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1744_
timestamp 1700315010
transform -1 0 2930 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1745_
timestamp 1700315010
transform -1 0 3230 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1746_
timestamp 1700315010
transform 1 0 3050 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1747_
timestamp 1700315010
transform 1 0 3350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1748_
timestamp 1700315010
transform -1 0 5090 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1749_
timestamp 1700315010
transform 1 0 5210 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1750_
timestamp 1700315010
transform 1 0 5430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1751_
timestamp 1700315010
transform 1 0 5370 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1752_
timestamp 1700315010
transform -1 0 5270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1753_
timestamp 1700315010
transform 1 0 5370 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1754_
timestamp 1700315010
transform 1 0 5150 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1755_
timestamp 1700315010
transform 1 0 5370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1756_
timestamp 1700315010
transform 1 0 4830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1757_
timestamp 1700315010
transform -1 0 4390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1758_
timestamp 1700315010
transform 1 0 4230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1759_
timestamp 1700315010
transform 1 0 3990 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1760_
timestamp 1700315010
transform 1 0 4510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1761_
timestamp 1700315010
transform -1 0 4690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1762_
timestamp 1700315010
transform -1 0 5130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1763_
timestamp 1700315010
transform 1 0 5270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1764_
timestamp 1700315010
transform 1 0 5590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1765_
timestamp 1700315010
transform 1 0 5730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1766_
timestamp 1700315010
transform 1 0 5830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1767_
timestamp 1700315010
transform 1 0 4890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1768_
timestamp 1700315010
transform -1 0 4750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1769_
timestamp 1700315010
transform -1 0 4590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1770_
timestamp 1700315010
transform -1 0 5010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1771_
timestamp 1700315010
transform 1 0 5510 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1772_
timestamp 1700315010
transform 1 0 5530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1773_
timestamp 1700315010
transform -1 0 5810 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1774_
timestamp 1700315010
transform -1 0 5590 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1775_
timestamp 1700315010
transform -1 0 5710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1776_
timestamp 1700315010
transform 1 0 5710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1777_
timestamp 1700315010
transform 1 0 4930 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1778_
timestamp 1700315010
transform 1 0 4470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1779_
timestamp 1700315010
transform 1 0 4350 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1780_
timestamp 1700315010
transform 1 0 4170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1781_
timestamp 1700315010
transform 1 0 4630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1782_
timestamp 1700315010
transform 1 0 4790 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1783_
timestamp 1700315010
transform 1 0 5610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1784_
timestamp 1700315010
transform 1 0 5470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1785_
timestamp 1700315010
transform -1 0 5810 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1786_
timestamp 1700315010
transform 1 0 5950 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1787_
timestamp 1700315010
transform -1 0 5890 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1788_
timestamp 1700315010
transform 1 0 5710 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1789_
timestamp 1700315010
transform 1 0 5990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1790_
timestamp 1700315010
transform 1 0 5990 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1791_
timestamp 1700315010
transform 1 0 5970 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1792_
timestamp 1700315010
transform 1 0 4650 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1793_
timestamp 1700315010
transform 1 0 4510 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1794_
timestamp 1700315010
transform 1 0 4870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1795_
timestamp 1700315010
transform -1 0 5570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1796_
timestamp 1700315010
transform 1 0 5410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1797_
timestamp 1700315010
transform -1 0 5030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1798_
timestamp 1700315010
transform -1 0 5870 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1799_
timestamp 1700315010
transform -1 0 5870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1800_
timestamp 1700315010
transform -1 0 5850 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1801_
timestamp 1700315010
transform 1 0 5410 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1802_
timestamp 1700315010
transform 1 0 4750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1803_
timestamp 1700315010
transform 1 0 5870 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1804_
timestamp 1700315010
transform -1 0 5890 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1805_
timestamp 1700315010
transform 1 0 5990 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1806_
timestamp 1700315010
transform -1 0 5690 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1807_
timestamp 1700315010
transform 1 0 5670 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1808_
timestamp 1700315010
transform 1 0 5530 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1809_
timestamp 1700315010
transform 1 0 5630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1810_
timestamp 1700315010
transform 1 0 5890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1811_
timestamp 1700315010
transform 1 0 5730 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1812_
timestamp 1700315010
transform 1 0 5970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1813_
timestamp 1700315010
transform -1 0 5990 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1814_
timestamp 1700315010
transform -1 0 6010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1815_
timestamp 1700315010
transform 1 0 5830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1816_
timestamp 1700315010
transform -1 0 5990 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1817_
timestamp 1700315010
transform -1 0 5870 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1818_
timestamp 1700315010
transform -1 0 3270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1819_
timestamp 1700315010
transform -1 0 2590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1820_
timestamp 1700315010
transform -1 0 4610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1821_
timestamp 1700315010
transform -1 0 5630 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1822_
timestamp 1700315010
transform 1 0 5470 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1823_
timestamp 1700315010
transform 1 0 5350 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1824_
timestamp 1700315010
transform 1 0 4970 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1825_
timestamp 1700315010
transform 1 0 4590 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1826_
timestamp 1700315010
transform 1 0 5750 0 -1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert0
timestamp 1700315010
transform 1 0 3930 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert1
timestamp 1700315010
transform -1 0 2210 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert2
timestamp 1700315010
transform -1 0 2330 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert3
timestamp 1700315010
transform -1 0 2270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert4
timestamp 1700315010
transform -1 0 4410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert5
timestamp 1700315010
transform -1 0 3770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert6
timestamp 1700315010
transform -1 0 2730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert7
timestamp 1700315010
transform -1 0 3410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert13
timestamp 1700315010
transform 1 0 5190 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert14
timestamp 1700315010
transform -1 0 3830 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert15
timestamp 1700315010
transform -1 0 4350 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert16
timestamp 1700315010
transform -1 0 4030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert17
timestamp 1700315010
transform 1 0 2530 0 1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert18
timestamp 1700315010
transform -1 0 2350 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert19
timestamp 1700315010
transform 1 0 3030 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert20
timestamp 1700315010
transform -1 0 2430 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert21
timestamp 1700315010
transform 1 0 5330 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert22
timestamp 1700315010
transform -1 0 4210 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert23
timestamp 1700315010
transform 1 0 4250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert24
timestamp 1700315010
transform 1 0 5290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert25
timestamp 1700315010
transform -1 0 2350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert26
timestamp 1700315010
transform -1 0 2650 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert27
timestamp 1700315010
transform -1 0 2410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert28
timestamp 1700315010
transform 1 0 3170 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert29
timestamp 1700315010
transform -1 0 2190 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert30
timestamp 1700315010
transform 1 0 3390 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert31
timestamp 1700315010
transform -1 0 2210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert32
timestamp 1700315010
transform 1 0 3510 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert33
timestamp 1700315010
transform -1 0 5090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert34
timestamp 1700315010
transform -1 0 6010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert35
timestamp 1700315010
transform -1 0 4950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert36
timestamp 1700315010
transform -1 0 5950 0 1 5470
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert8
timestamp 1700315010
transform -1 0 4550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1700315010
transform -1 0 4950 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 5810 0 1 790
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert11
timestamp 1700315010
transform -1 0 5190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 4970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__889_
timestamp 1700315010
transform 1 0 5370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__890_
timestamp 1700315010
transform -1 0 4990 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__892_
timestamp 1700315010
transform 1 0 5390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__893_
timestamp 1700315010
transform -1 0 5250 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__894_
timestamp 1700315010
transform 1 0 5510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__896_
timestamp 1700315010
transform -1 0 5130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__897_
timestamp 1700315010
transform 1 0 5130 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__899_
timestamp 1700315010
transform 1 0 5270 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__900_
timestamp 1700315010
transform -1 0 5870 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__902_
timestamp 1700315010
transform 1 0 5810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__903_
timestamp 1700315010
transform 1 0 4910 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__905_
timestamp 1700315010
transform -1 0 5710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__906_
timestamp 1700315010
transform -1 0 4230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__908_
timestamp 1700315010
transform 1 0 5970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__909_
timestamp 1700315010
transform 1 0 5610 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__911_
timestamp 1700315010
transform 1 0 5430 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__912_
timestamp 1700315010
transform 1 0 5770 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__914_
timestamp 1700315010
transform -1 0 5270 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__915_
timestamp 1700315010
transform 1 0 5250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__916_
timestamp 1700315010
transform -1 0 5650 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__918_
timestamp 1700315010
transform -1 0 5410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__919_
timestamp 1700315010
transform 1 0 5410 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__921_
timestamp 1700315010
transform 1 0 5670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__922_
timestamp 1700315010
transform 1 0 5390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__924_
timestamp 1700315010
transform 1 0 5910 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__925_
timestamp 1700315010
transform -1 0 5990 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__927_
timestamp 1700315010
transform 1 0 4870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__928_
timestamp 1700315010
transform 1 0 4710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__930_
timestamp 1700315010
transform 1 0 3690 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__931_
timestamp 1700315010
transform -1 0 3850 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__933_
timestamp 1700315010
transform -1 0 4430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__934_
timestamp 1700315010
transform 1 0 4550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__936_
timestamp 1700315010
transform 1 0 4090 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__937_
timestamp 1700315010
transform -1 0 4010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__939_
timestamp 1700315010
transform 1 0 3670 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__940_
timestamp 1700315010
transform 1 0 3470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__941_
timestamp 1700315010
transform -1 0 3270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__943_
timestamp 1700315010
transform 1 0 3490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__944_
timestamp 1700315010
transform -1 0 5330 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__946_
timestamp 1700315010
transform 1 0 5430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__947_
timestamp 1700315010
transform 1 0 5670 0 1 790
box -12 -8 32 272
use FILL  FILL_2__949_
timestamp 1700315010
transform 1 0 5110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__950_
timestamp 1700315010
transform -1 0 4670 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__952_
timestamp 1700315010
transform 1 0 2350 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__953_
timestamp 1700315010
transform 1 0 2650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__955_
timestamp 1700315010
transform 1 0 2770 0 1 790
box -12 -8 32 272
use FILL  FILL_2__956_
timestamp 1700315010
transform 1 0 3190 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__958_
timestamp 1700315010
transform 1 0 3630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__959_
timestamp 1700315010
transform 1 0 3630 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__961_
timestamp 1700315010
transform -1 0 3490 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__962_
timestamp 1700315010
transform 1 0 3790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__963_
timestamp 1700315010
transform 1 0 2930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__965_
timestamp 1700315010
transform 1 0 2510 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__966_
timestamp 1700315010
transform 1 0 3350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__968_
timestamp 1700315010
transform 1 0 2590 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__969_
timestamp 1700315010
transform -1 0 2790 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__971_
timestamp 1700315010
transform 1 0 3050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__972_
timestamp 1700315010
transform -1 0 3210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__974_
timestamp 1700315010
transform -1 0 3510 0 1 790
box -12 -8 32 272
use FILL  FILL_2__975_
timestamp 1700315010
transform 1 0 3070 0 1 790
box -12 -8 32 272
use FILL  FILL_2__977_
timestamp 1700315010
transform 1 0 2130 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__978_
timestamp 1700315010
transform 1 0 2510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__980_
timestamp 1700315010
transform 1 0 2910 0 1 790
box -12 -8 32 272
use FILL  FILL_2__981_
timestamp 1700315010
transform 1 0 3650 0 1 790
box -12 -8 32 272
use FILL  FILL_2__983_
timestamp 1700315010
transform -1 0 2770 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__984_
timestamp 1700315010
transform -1 0 2450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__985_
timestamp 1700315010
transform -1 0 2370 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__987_
timestamp 1700315010
transform -1 0 1610 0 1 790
box -12 -8 32 272
use FILL  FILL_2__988_
timestamp 1700315010
transform -1 0 1390 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__990_
timestamp 1700315010
transform 1 0 1870 0 1 790
box -12 -8 32 272
use FILL  FILL_2__991_
timestamp 1700315010
transform 1 0 2410 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__993_
timestamp 1700315010
transform 1 0 2030 0 1 790
box -12 -8 32 272
use FILL  FILL_2__994_
timestamp 1700315010
transform 1 0 2610 0 1 790
box -12 -8 32 272
use FILL  FILL_2__996_
timestamp 1700315010
transform 1 0 1710 0 1 790
box -12 -8 32 272
use FILL  FILL_2__997_
timestamp 1700315010
transform -1 0 1450 0 1 790
box -12 -8 32 272
use FILL  FILL_2__999_
timestamp 1700315010
transform 1 0 2210 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1001_
timestamp 1700315010
transform 1 0 2790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1002_
timestamp 1700315010
transform 1 0 2350 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1004_
timestamp 1700315010
transform 1 0 2490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1005_
timestamp 1700315010
transform -1 0 2350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1007_
timestamp 1700315010
transform -1 0 1690 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1008_
timestamp 1700315010
transform 1 0 1790 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1009_
timestamp 1700315010
transform -1 0 1970 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1011_
timestamp 1700315010
transform -1 0 2230 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1012_
timestamp 1700315010
transform -1 0 1490 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1014_
timestamp 1700315010
transform -1 0 2210 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1015_
timestamp 1700315010
transform -1 0 2070 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1017_
timestamp 1700315010
transform 1 0 2210 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1018_
timestamp 1700315010
transform -1 0 2390 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1020_
timestamp 1700315010
transform -1 0 1530 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1021_
timestamp 1700315010
transform -1 0 1450 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1023_
timestamp 1700315010
transform 1 0 1150 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1024_
timestamp 1700315010
transform 1 0 1510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1026_
timestamp 1700315010
transform 1 0 1270 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1027_
timestamp 1700315010
transform 1 0 1510 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1029_
timestamp 1700315010
transform -1 0 930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1030_
timestamp 1700315010
transform -1 0 1610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1032_
timestamp 1700315010
transform -1 0 1250 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1033_
timestamp 1700315010
transform -1 0 1090 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1034_
timestamp 1700315010
transform -1 0 1670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1036_
timestamp 1700315010
transform -1 0 1190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1037_
timestamp 1700315010
transform -1 0 1070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1039_
timestamp 1700315010
transform -1 0 1350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1040_
timestamp 1700315010
transform -1 0 2070 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1042_
timestamp 1700315010
transform 1 0 1910 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1043_
timestamp 1700315010
transform 1 0 2310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1045_
timestamp 1700315010
transform 1 0 2110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1046_
timestamp 1700315010
transform -1 0 1630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1048_
timestamp 1700315010
transform -1 0 1970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1049_
timestamp 1700315010
transform -1 0 1470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1051_
timestamp 1700315010
transform -1 0 710 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1052_
timestamp 1700315010
transform 1 0 1210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1054_
timestamp 1700315010
transform -1 0 1390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1055_
timestamp 1700315010
transform -1 0 970 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1056_
timestamp 1700315010
transform 1 0 1010 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1058_
timestamp 1700315010
transform 1 0 1270 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1059_
timestamp 1700315010
transform 1 0 1110 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1061_
timestamp 1700315010
transform -1 0 2950 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1062_
timestamp 1700315010
transform -1 0 1930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1064_
timestamp 1700315010
transform 1 0 1390 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1065_
timestamp 1700315010
transform -1 0 950 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1067_
timestamp 1700315010
transform 1 0 1310 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1068_
timestamp 1700315010
transform -1 0 870 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1070_
timestamp 1700315010
transform 1 0 1970 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1071_
timestamp 1700315010
transform 1 0 1590 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1073_
timestamp 1700315010
transform -1 0 970 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1074_
timestamp 1700315010
transform -1 0 810 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1076_
timestamp 1700315010
transform -1 0 990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1077_
timestamp 1700315010
transform 1 0 1130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1079_
timestamp 1700315010
transform -1 0 910 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1080_
timestamp 1700315010
transform -1 0 870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1081_
timestamp 1700315010
transform -1 0 230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1083_
timestamp 1700315010
transform -1 0 770 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1084_
timestamp 1700315010
transform -1 0 390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1086_
timestamp 1700315010
transform 1 0 690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1087_
timestamp 1700315010
transform 1 0 530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1089_
timestamp 1700315010
transform 1 0 1970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1090_
timestamp 1700315010
transform 1 0 1570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1092_
timestamp 1700315010
transform -1 0 2050 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1093_
timestamp 1700315010
transform 1 0 1890 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1095_
timestamp 1700315010
transform -1 0 1870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1096_
timestamp 1700315010
transform -1 0 1710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1098_
timestamp 1700315010
transform -1 0 1750 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1099_
timestamp 1700315010
transform -1 0 1450 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1101_
timestamp 1700315010
transform -1 0 70 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1102_
timestamp 1700315010
transform -1 0 950 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1103_
timestamp 1700315010
transform 1 0 630 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1105_
timestamp 1700315010
transform 1 0 190 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1106_
timestamp 1700315010
transform -1 0 70 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1108_
timestamp 1700315010
transform 1 0 890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1109_
timestamp 1700315010
transform -1 0 370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1111_
timestamp 1700315010
transform -1 0 70 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1112_
timestamp 1700315010
transform -1 0 2050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1114_
timestamp 1700315010
transform -1 0 1790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1115_
timestamp 1700315010
transform -1 0 530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1117_
timestamp 1700315010
transform 1 0 770 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1118_
timestamp 1700315010
transform -1 0 370 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1120_
timestamp 1700315010
transform 1 0 490 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1121_
timestamp 1700315010
transform 1 0 910 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1123_
timestamp 1700315010
transform -1 0 670 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1124_
timestamp 1700315010
transform 1 0 530 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1126_
timestamp 1700315010
transform -1 0 70 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1127_
timestamp 1700315010
transform 1 0 590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1128_
timestamp 1700315010
transform -1 0 350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1130_
timestamp 1700315010
transform 1 0 370 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1131_
timestamp 1700315010
transform -1 0 370 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1133_
timestamp 1700315010
transform -1 0 70 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1134_
timestamp 1700315010
transform -1 0 230 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1136_
timestamp 1700315010
transform -1 0 330 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1137_
timestamp 1700315010
transform -1 0 70 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1139_
timestamp 1700315010
transform 1 0 610 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1140_
timestamp 1700315010
transform 1 0 1810 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1142_
timestamp 1700315010
transform 1 0 2530 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1143_
timestamp 1700315010
transform 1 0 3330 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1145_
timestamp 1700315010
transform 1 0 3030 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1146_
timestamp 1700315010
transform -1 0 3370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1148_
timestamp 1700315010
transform 1 0 3190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1149_
timestamp 1700315010
transform -1 0 3210 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1150_
timestamp 1700315010
transform 1 0 2830 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1152_
timestamp 1700315010
transform -1 0 3190 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1153_
timestamp 1700315010
transform 1 0 2370 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1155_
timestamp 1700315010
transform 1 0 2670 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1156_
timestamp 1700315010
transform -1 0 2670 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1158_
timestamp 1700315010
transform 1 0 1190 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1159_
timestamp 1700315010
transform -1 0 1750 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1161_
timestamp 1700315010
transform 1 0 770 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1162_
timestamp 1700315010
transform 1 0 1350 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1164_
timestamp 1700315010
transform 1 0 3770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1165_
timestamp 1700315010
transform -1 0 3930 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1167_
timestamp 1700315010
transform 1 0 4310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1168_
timestamp 1700315010
transform -1 0 3490 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1170_
timestamp 1700315010
transform 1 0 3510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1171_
timestamp 1700315010
transform 1 0 4070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1173_
timestamp 1700315010
transform 1 0 4070 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1174_
timestamp 1700315010
transform 1 0 3610 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1175_
timestamp 1700315010
transform -1 0 3790 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1177_
timestamp 1700315010
transform -1 0 3010 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1178_
timestamp 1700315010
transform -1 0 2990 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1180_
timestamp 1700315010
transform 1 0 2130 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1181_
timestamp 1700315010
transform 1 0 3310 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1183_
timestamp 1700315010
transform 1 0 3810 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1184_
timestamp 1700315010
transform -1 0 3670 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1186_
timestamp 1700315010
transform 1 0 4050 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1187_
timestamp 1700315010
transform -1 0 3350 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1189_
timestamp 1700315010
transform 1 0 3770 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1190_
timestamp 1700315010
transform 1 0 3890 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1192_
timestamp 1700315010
transform 1 0 4490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1193_
timestamp 1700315010
transform 1 0 4370 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1195_
timestamp 1700315010
transform 1 0 4490 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1196_
timestamp 1700315010
transform 1 0 3930 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1197_
timestamp 1700315010
transform -1 0 4110 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1199_
timestamp 1700315010
transform 1 0 2810 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1200_
timestamp 1700315010
transform 1 0 3510 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1202_
timestamp 1700315010
transform 1 0 4070 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1203_
timestamp 1700315010
transform 1 0 3550 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1205_
timestamp 1700315010
transform 1 0 2690 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1206_
timestamp 1700315010
transform -1 0 70 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1208_
timestamp 1700315010
transform -1 0 70 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1209_
timestamp 1700315010
transform 1 0 2390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1211_
timestamp 1700315010
transform -1 0 2190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1212_
timestamp 1700315010
transform 1 0 1850 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1214_
timestamp 1700315010
transform 1 0 2230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1215_
timestamp 1700315010
transform -1 0 1410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1217_
timestamp 1700315010
transform 1 0 2010 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1218_
timestamp 1700315010
transform -1 0 1830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1219_
timestamp 1700315010
transform 1 0 1250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1221_
timestamp 1700315010
transform -1 0 1550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1222_
timestamp 1700315010
transform -1 0 1930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1224_
timestamp 1700315010
transform -1 0 2130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1225_
timestamp 1700315010
transform 1 0 1950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1227_
timestamp 1700315010
transform 1 0 1590 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1228_
timestamp 1700315010
transform 1 0 1990 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1230_
timestamp 1700315010
transform 1 0 1870 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1231_
timestamp 1700315010
transform -1 0 1730 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1233_
timestamp 1700315010
transform 1 0 330 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1234_
timestamp 1700315010
transform 1 0 1130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1236_
timestamp 1700315010
transform -1 0 310 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1237_
timestamp 1700315010
transform 1 0 590 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1239_
timestamp 1700315010
transform -1 0 530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1240_
timestamp 1700315010
transform -1 0 450 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1242_
timestamp 1700315010
transform 1 0 650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1243_
timestamp 1700315010
transform 1 0 370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1244_
timestamp 1700315010
transform 1 0 210 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1246_
timestamp 1700315010
transform -1 0 70 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1247_
timestamp 1700315010
transform -1 0 70 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1249_
timestamp 1700315010
transform 1 0 50 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1250_
timestamp 1700315010
transform -1 0 230 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1252_
timestamp 1700315010
transform 1 0 490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1253_
timestamp 1700315010
transform 1 0 50 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1255_
timestamp 1700315010
transform -1 0 70 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1256_
timestamp 1700315010
transform 1 0 350 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1258_
timestamp 1700315010
transform 1 0 370 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1259_
timestamp 1700315010
transform -1 0 850 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1261_
timestamp 1700315010
transform 1 0 970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1262_
timestamp 1700315010
transform 1 0 210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1264_
timestamp 1700315010
transform 1 0 510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1265_
timestamp 1700315010
transform -1 0 690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1266_
timestamp 1700315010
transform -1 0 670 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1268_
timestamp 1700315010
transform 1 0 1090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1269_
timestamp 1700315010
transform 1 0 1250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1271_
timestamp 1700315010
transform -1 0 3110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1272_
timestamp 1700315010
transform 1 0 5010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1274_
timestamp 1700315010
transform 1 0 4170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1275_
timestamp 1700315010
transform 1 0 3970 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1277_
timestamp 1700315010
transform 1 0 4130 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1278_
timestamp 1700315010
transform 1 0 4770 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1280_
timestamp 1700315010
transform -1 0 3570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1281_
timestamp 1700315010
transform -1 0 3870 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1283_
timestamp 1700315010
transform -1 0 3710 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1284_
timestamp 1700315010
transform -1 0 1670 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1286_
timestamp 1700315010
transform -1 0 1530 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1287_
timestamp 1700315010
transform 1 0 1910 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1289_
timestamp 1700315010
transform 1 0 2850 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1290_
timestamp 1700315010
transform -1 0 3170 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1291_
timestamp 1700315010
transform -1 0 2410 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1293_
timestamp 1700315010
transform -1 0 2650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1294_
timestamp 1700315010
transform 1 0 1270 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1296_
timestamp 1700315010
transform -1 0 1670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1297_
timestamp 1700315010
transform 1 0 1630 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1299_
timestamp 1700315010
transform 1 0 790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1300_
timestamp 1700315010
transform -1 0 1630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1302_
timestamp 1700315010
transform -1 0 1930 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1303_
timestamp 1700315010
transform -1 0 2090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1305_
timestamp 1700315010
transform -1 0 1430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1306_
timestamp 1700315010
transform 1 0 790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1308_
timestamp 1700315010
transform -1 0 70 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1309_
timestamp 1700315010
transform 1 0 1330 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1311_
timestamp 1700315010
transform 1 0 1110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1312_
timestamp 1700315010
transform -1 0 1770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1313_
timestamp 1700315010
transform -1 0 1370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1315_
timestamp 1700315010
transform 1 0 1310 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1316_
timestamp 1700315010
transform -1 0 790 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1318_
timestamp 1700315010
transform 1 0 2790 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1319_
timestamp 1700315010
transform -1 0 2070 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1321_
timestamp 1700315010
transform -1 0 1630 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1322_
timestamp 1700315010
transform -1 0 1170 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1324_
timestamp 1700315010
transform -1 0 830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1325_
timestamp 1700315010
transform -1 0 1030 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1327_
timestamp 1700315010
transform -1 0 70 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1328_
timestamp 1700315010
transform -1 0 70 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1330_
timestamp 1700315010
transform -1 0 510 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1331_
timestamp 1700315010
transform 1 0 190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1333_
timestamp 1700315010
transform 1 0 810 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1334_
timestamp 1700315010
transform 1 0 510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1336_
timestamp 1700315010
transform 1 0 490 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1337_
timestamp 1700315010
transform 1 0 1130 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1338_
timestamp 1700315010
transform 1 0 50 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1340_
timestamp 1700315010
transform 1 0 650 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1341_
timestamp 1700315010
transform 1 0 170 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1343_
timestamp 1700315010
transform 1 0 330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1344_
timestamp 1700315010
transform -1 0 890 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1346_
timestamp 1700315010
transform 1 0 910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1347_
timestamp 1700315010
transform 1 0 1030 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1349_
timestamp 1700315010
transform -1 0 1410 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1350_
timestamp 1700315010
transform 1 0 530 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1352_
timestamp 1700315010
transform 1 0 1750 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1353_
timestamp 1700315010
transform -1 0 1210 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1355_
timestamp 1700315010
transform -1 0 2170 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1356_
timestamp 1700315010
transform 1 0 3290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1358_
timestamp 1700315010
transform 1 0 3590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1359_
timestamp 1700315010
transform 1 0 4570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1360_
timestamp 1700315010
transform 1 0 4510 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1362_
timestamp 1700315010
transform 1 0 4350 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1363_
timestamp 1700315010
transform -1 0 4070 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1365_
timestamp 1700315010
transform -1 0 4830 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1366_
timestamp 1700315010
transform -1 0 1570 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1368_
timestamp 1700315010
transform 1 0 2110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1369_
timestamp 1700315010
transform 1 0 2930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1371_
timestamp 1700315010
transform 1 0 2510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1372_
timestamp 1700315010
transform -1 0 1290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1374_
timestamp 1700315010
transform -1 0 530 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1375_
timestamp 1700315010
transform -1 0 350 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1377_
timestamp 1700315010
transform -1 0 890 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1378_
timestamp 1700315010
transform -1 0 1190 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1380_
timestamp 1700315010
transform -1 0 1170 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1381_
timestamp 1700315010
transform -1 0 1010 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1383_
timestamp 1700315010
transform -1 0 1010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1384_
timestamp 1700315010
transform -1 0 1170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1385_
timestamp 1700315010
transform -1 0 850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1387_
timestamp 1700315010
transform 1 0 630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1388_
timestamp 1700315010
transform 1 0 1590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1390_
timestamp 1700315010
transform -1 0 1690 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1391_
timestamp 1700315010
transform -1 0 1510 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1393_
timestamp 1700315010
transform 1 0 1890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1394_
timestamp 1700315010
transform 1 0 1390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1396_
timestamp 1700315010
transform -1 0 590 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1397_
timestamp 1700315010
transform -1 0 70 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1399_
timestamp 1700315010
transform -1 0 690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1400_
timestamp 1700315010
transform -1 0 310 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1402_
timestamp 1700315010
transform -1 0 170 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1403_
timestamp 1700315010
transform 1 0 350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1405_
timestamp 1700315010
transform 1 0 350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1406_
timestamp 1700315010
transform -1 0 70 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1407_
timestamp 1700315010
transform -1 0 70 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1409_
timestamp 1700315010
transform -1 0 230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1410_
timestamp 1700315010
transform 1 0 210 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1412_
timestamp 1700315010
transform 1 0 630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1413_
timestamp 1700315010
transform -1 0 70 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1415_
timestamp 1700315010
transform -1 0 1310 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1416_
timestamp 1700315010
transform 1 0 1910 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1418_
timestamp 1700315010
transform -1 0 1230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1419_
timestamp 1700315010
transform 1 0 1370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1421_
timestamp 1700315010
transform -1 0 2470 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1422_
timestamp 1700315010
transform 1 0 2790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1424_
timestamp 1700315010
transform 1 0 2870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1425_
timestamp 1700315010
transform -1 0 3010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1427_
timestamp 1700315010
transform 1 0 4610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1428_
timestamp 1700315010
transform -1 0 4310 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1429_
timestamp 1700315010
transform 1 0 4350 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1431_
timestamp 1700315010
transform -1 0 4730 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1432_
timestamp 1700315010
transform 1 0 4750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1434_
timestamp 1700315010
transform 1 0 4650 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1435_
timestamp 1700315010
transform 1 0 5950 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1437_
timestamp 1700315010
transform -1 0 3890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1438_
timestamp 1700315010
transform 1 0 2670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1440_
timestamp 1700315010
transform -1 0 1210 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1441_
timestamp 1700315010
transform 1 0 510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1443_
timestamp 1700315010
transform -1 0 2090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1444_
timestamp 1700315010
transform -1 0 1430 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1446_
timestamp 1700315010
transform 1 0 1550 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1447_
timestamp 1700315010
transform 1 0 1690 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1449_
timestamp 1700315010
transform -1 0 1930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1450_
timestamp 1700315010
transform -1 0 1570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1452_
timestamp 1700315010
transform 1 0 1910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1453_
timestamp 1700315010
transform 1 0 2090 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1454_
timestamp 1700315010
transform 1 0 1930 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1456_
timestamp 1700315010
transform -1 0 2170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1457_
timestamp 1700315010
transform -1 0 1970 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1459_
timestamp 1700315010
transform -1 0 490 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1460_
timestamp 1700315010
transform 1 0 1750 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1462_
timestamp 1700315010
transform -1 0 190 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1463_
timestamp 1700315010
transform -1 0 1450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1465_
timestamp 1700315010
transform -1 0 1050 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1466_
timestamp 1700315010
transform -1 0 610 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1468_
timestamp 1700315010
transform 1 0 1450 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1469_
timestamp 1700315010
transform -1 0 1130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1471_
timestamp 1700315010
transform 1 0 790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1472_
timestamp 1700315010
transform 1 0 950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1474_
timestamp 1700315010
transform 1 0 2790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1475_
timestamp 1700315010
transform 1 0 2750 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1476_
timestamp 1700315010
transform 1 0 2990 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1478_
timestamp 1700315010
transform 1 0 3250 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1479_
timestamp 1700315010
transform 1 0 3530 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1481_
timestamp 1700315010
transform -1 0 4370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1482_
timestamp 1700315010
transform 1 0 4650 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1484_
timestamp 1700315010
transform -1 0 5530 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1485_
timestamp 1700315010
transform 1 0 5510 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1487_
timestamp 1700315010
transform 1 0 5830 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1488_
timestamp 1700315010
transform 1 0 2190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1490_
timestamp 1700315010
transform -1 0 2370 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1491_
timestamp 1700315010
transform -1 0 2890 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1493_
timestamp 1700315010
transform -1 0 2270 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1494_
timestamp 1700315010
transform 1 0 2570 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1496_
timestamp 1700315010
transform 1 0 2410 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1497_
timestamp 1700315010
transform 1 0 2610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1499_
timestamp 1700315010
transform 1 0 2230 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1500_
timestamp 1700315010
transform 1 0 2450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1501_
timestamp 1700315010
transform 1 0 2730 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1503_
timestamp 1700315010
transform 1 0 2790 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1504_
timestamp 1700315010
transform 1 0 2870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1506_
timestamp 1700315010
transform -1 0 2650 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1507_
timestamp 1700315010
transform -1 0 2490 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1509_
timestamp 1700315010
transform 1 0 2050 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1510_
timestamp 1700315010
transform -1 0 1930 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1512_
timestamp 1700315010
transform -1 0 2730 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1513_
timestamp 1700315010
transform 1 0 3330 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1515_
timestamp 1700315010
transform 1 0 3170 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1516_
timestamp 1700315010
transform -1 0 2550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1518_
timestamp 1700315010
transform -1 0 3230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1519_
timestamp 1700315010
transform 1 0 2930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1521_
timestamp 1700315010
transform 1 0 2570 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1522_
timestamp 1700315010
transform 1 0 2730 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1523_
timestamp 1700315010
transform 1 0 2850 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1525_
timestamp 1700315010
transform -1 0 5490 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1526_
timestamp 1700315010
transform -1 0 4990 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1528_
timestamp 1700315010
transform 1 0 4330 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1529_
timestamp 1700315010
transform 1 0 4590 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1531_
timestamp 1700315010
transform -1 0 5090 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1532_
timestamp 1700315010
transform 1 0 5230 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1534_
timestamp 1700315010
transform -1 0 5170 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1535_
timestamp 1700315010
transform -1 0 3770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1537_
timestamp 1700315010
transform 1 0 2810 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1538_
timestamp 1700315010
transform 1 0 2590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1540_
timestamp 1700315010
transform -1 0 2650 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1541_
timestamp 1700315010
transform -1 0 2810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1543_
timestamp 1700315010
transform 1 0 2650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1544_
timestamp 1700315010
transform 1 0 2450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1546_
timestamp 1700315010
transform -1 0 2510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1547_
timestamp 1700315010
transform -1 0 2690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1548_
timestamp 1700315010
transform -1 0 3050 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1550_
timestamp 1700315010
transform 1 0 3470 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1551_
timestamp 1700315010
transform 1 0 3910 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1553_
timestamp 1700315010
transform -1 0 5070 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1554_
timestamp 1700315010
transform 1 0 5230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1556_
timestamp 1700315010
transform -1 0 4990 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1557_
timestamp 1700315010
transform -1 0 4870 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1559_
timestamp 1700315010
transform 1 0 3530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1560_
timestamp 1700315010
transform 1 0 3650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1562_
timestamp 1700315010
transform 1 0 2690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1563_
timestamp 1700315010
transform 1 0 3710 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1565_
timestamp 1700315010
transform -1 0 2170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1566_
timestamp 1700315010
transform -1 0 2310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1568_
timestamp 1700315010
transform 1 0 3330 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1569_
timestamp 1700315010
transform 1 0 3950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1570_
timestamp 1700315010
transform 1 0 3370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1572_
timestamp 1700315010
transform 1 0 3450 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1573_
timestamp 1700315010
transform 1 0 4110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1575_
timestamp 1700315010
transform 1 0 4330 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1576_
timestamp 1700315010
transform 1 0 4170 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1578_
timestamp 1700315010
transform 1 0 5710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1579_
timestamp 1700315010
transform -1 0 5130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1581_
timestamp 1700315010
transform 1 0 4890 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1582_
timestamp 1700315010
transform -1 0 4510 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1584_
timestamp 1700315010
transform 1 0 2950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1585_
timestamp 1700315010
transform 1 0 3110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1587_
timestamp 1700315010
transform 1 0 2550 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1588_
timestamp 1700315010
transform -1 0 3870 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1590_
timestamp 1700315010
transform 1 0 4790 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1591_
timestamp 1700315010
transform -1 0 4750 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1593_
timestamp 1700315010
transform -1 0 4350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1594_
timestamp 1700315010
transform 1 0 4310 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1595_
timestamp 1700315010
transform 1 0 3990 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1597_
timestamp 1700315010
transform 1 0 4010 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1598_
timestamp 1700315010
transform -1 0 4170 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1600_
timestamp 1700315010
transform -1 0 4030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1601_
timestamp 1700315010
transform 1 0 3310 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1603_
timestamp 1700315010
transform 1 0 2950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1604_
timestamp 1700315010
transform -1 0 3110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1606_
timestamp 1700315010
transform -1 0 5170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1607_
timestamp 1700315010
transform 1 0 4430 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1636_
timestamp 1700315010
transform -1 0 5910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1637_
timestamp 1700315010
transform 1 0 5910 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1639_
timestamp 1700315010
transform 1 0 5210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1640_
timestamp 1700315010
transform 1 0 5210 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1642_
timestamp 1700315010
transform -1 0 3170 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1643_
timestamp 1700315010
transform -1 0 3010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1644_
timestamp 1700315010
transform -1 0 3870 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1646_
timestamp 1700315010
transform -1 0 4110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1647_
timestamp 1700315010
transform 1 0 3170 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1649_
timestamp 1700315010
transform -1 0 4290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1650_
timestamp 1700315010
transform -1 0 4450 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1652_
timestamp 1700315010
transform -1 0 3630 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1653_
timestamp 1700315010
transform 1 0 4150 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1655_
timestamp 1700315010
transform -1 0 5670 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1656_
timestamp 1700315010
transform 1 0 5930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1658_
timestamp 1700315010
transform 1 0 5630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1659_
timestamp 1700315010
transform -1 0 5350 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1661_
timestamp 1700315010
transform 1 0 5350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1662_
timestamp 1700315010
transform -1 0 3470 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1664_
timestamp 1700315010
transform -1 0 3450 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1665_
timestamp 1700315010
transform -1 0 3650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1666_
timestamp 1700315010
transform -1 0 3830 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1668_
timestamp 1700315010
transform 1 0 3710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1669_
timestamp 1700315010
transform -1 0 4050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1671_
timestamp 1700315010
transform 1 0 5230 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1672_
timestamp 1700315010
transform -1 0 5670 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1674_
timestamp 1700315010
transform -1 0 5370 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1675_
timestamp 1700315010
transform -1 0 5550 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1677_
timestamp 1700315010
transform -1 0 4890 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1678_
timestamp 1700315010
transform -1 0 4930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1680_
timestamp 1700315010
transform 1 0 4630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1681_
timestamp 1700315010
transform -1 0 4010 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1683_
timestamp 1700315010
transform 1 0 4710 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1684_
timestamp 1700315010
transform 1 0 5030 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1686_
timestamp 1700315010
transform 1 0 4310 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1687_
timestamp 1700315010
transform -1 0 5110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1689_
timestamp 1700315010
transform 1 0 4890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1690_
timestamp 1700315010
transform 1 0 5090 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1691_
timestamp 1700315010
transform -1 0 4950 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1693_
timestamp 1700315010
transform 1 0 3110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1694_
timestamp 1700315010
transform -1 0 3290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1696_
timestamp 1700315010
transform -1 0 3050 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1697_
timestamp 1700315010
transform -1 0 3310 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1699_
timestamp 1700315010
transform -1 0 3890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1700_
timestamp 1700315010
transform -1 0 3910 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1702_
timestamp 1700315010
transform 1 0 3730 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1703_
timestamp 1700315010
transform -1 0 4590 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1705_
timestamp 1700315010
transform 1 0 4050 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1706_
timestamp 1700315010
transform -1 0 4350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1708_
timestamp 1700315010
transform 1 0 4490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1709_
timestamp 1700315010
transform -1 0 3670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1711_
timestamp 1700315010
transform -1 0 3570 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1712_
timestamp 1700315010
transform -1 0 3710 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1713_
timestamp 1700315010
transform -1 0 3410 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1715_
timestamp 1700315010
transform -1 0 3950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1716_
timestamp 1700315010
transform 1 0 4090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1718_
timestamp 1700315010
transform 1 0 4570 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1719_
timestamp 1700315010
transform 1 0 4730 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1721_
timestamp 1700315010
transform 1 0 4670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1722_
timestamp 1700315010
transform 1 0 4770 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1724_
timestamp 1700315010
transform -1 0 4810 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1725_
timestamp 1700315010
transform 1 0 4430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1727_
timestamp 1700315010
transform -1 0 4390 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1728_
timestamp 1700315010
transform -1 0 3030 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1730_
timestamp 1700315010
transform -1 0 3250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1731_
timestamp 1700315010
transform -1 0 3390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1733_
timestamp 1700315010
transform 1 0 3690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1734_
timestamp 1700315010
transform 1 0 4970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1736_
timestamp 1700315010
transform -1 0 5250 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1737_
timestamp 1700315010
transform 1 0 5070 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1738_
timestamp 1700315010
transform 1 0 5110 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1740_
timestamp 1700315010
transform -1 0 5170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1741_
timestamp 1700315010
transform 1 0 5230 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1743_
timestamp 1700315010
transform -1 0 2790 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1744_
timestamp 1700315010
transform -1 0 2950 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1746_
timestamp 1700315010
transform 1 0 3070 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1747_
timestamp 1700315010
transform 1 0 3370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1749_
timestamp 1700315010
transform 1 0 5230 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1750_
timestamp 1700315010
transform 1 0 5450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1752_
timestamp 1700315010
transform -1 0 5290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1753_
timestamp 1700315010
transform 1 0 5390 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1755_
timestamp 1700315010
transform 1 0 5390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1756_
timestamp 1700315010
transform 1 0 4850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1758_
timestamp 1700315010
transform 1 0 4250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1759_
timestamp 1700315010
transform 1 0 4010 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1760_
timestamp 1700315010
transform 1 0 4530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1762_
timestamp 1700315010
transform -1 0 5150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1763_
timestamp 1700315010
transform 1 0 5290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1765_
timestamp 1700315010
transform 1 0 5750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1766_
timestamp 1700315010
transform 1 0 5850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1768_
timestamp 1700315010
transform -1 0 4770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1769_
timestamp 1700315010
transform -1 0 4610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1771_
timestamp 1700315010
transform 1 0 5530 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1772_
timestamp 1700315010
transform 1 0 5550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1774_
timestamp 1700315010
transform -1 0 5610 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1775_
timestamp 1700315010
transform -1 0 5730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1777_
timestamp 1700315010
transform 1 0 4950 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1778_
timestamp 1700315010
transform 1 0 4490 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1780_
timestamp 1700315010
transform 1 0 4190 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1781_
timestamp 1700315010
transform 1 0 4650 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1783_
timestamp 1700315010
transform 1 0 5630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1784_
timestamp 1700315010
transform 1 0 5490 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1785_
timestamp 1700315010
transform -1 0 5830 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1787_
timestamp 1700315010
transform -1 0 5910 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1788_
timestamp 1700315010
transform 1 0 5730 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1790_
timestamp 1700315010
transform 1 0 6010 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1791_
timestamp 1700315010
transform 1 0 5990 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1793_
timestamp 1700315010
transform 1 0 4530 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1794_
timestamp 1700315010
transform 1 0 4890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1796_
timestamp 1700315010
transform 1 0 5430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1797_
timestamp 1700315010
transform -1 0 5050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1799_
timestamp 1700315010
transform -1 0 5890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1800_
timestamp 1700315010
transform -1 0 5870 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1802_
timestamp 1700315010
transform 1 0 4770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1803_
timestamp 1700315010
transform 1 0 5890 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1805_
timestamp 1700315010
transform 1 0 6010 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1806_
timestamp 1700315010
transform -1 0 5710 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1807_
timestamp 1700315010
transform 1 0 5690 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1809_
timestamp 1700315010
transform 1 0 5650 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1810_
timestamp 1700315010
transform 1 0 5910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1812_
timestamp 1700315010
transform 1 0 5990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1813_
timestamp 1700315010
transform -1 0 6010 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1815_
timestamp 1700315010
transform 1 0 5850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1816_
timestamp 1700315010
transform -1 0 6010 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1818_
timestamp 1700315010
transform -1 0 3290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1819_
timestamp 1700315010
transform -1 0 2610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1821_
timestamp 1700315010
transform -1 0 5650 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1822_
timestamp 1700315010
transform 1 0 5490 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1824_
timestamp 1700315010
transform 1 0 4990 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1825_
timestamp 1700315010
transform 1 0 4610 0 -1 270
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert0
timestamp 1700315010
transform 1 0 3950 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert1
timestamp 1700315010
transform -1 0 2230 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert3
timestamp 1700315010
transform -1 0 2290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert4
timestamp 1700315010
transform -1 0 4430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert6
timestamp 1700315010
transform -1 0 2750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert7
timestamp 1700315010
transform -1 0 3430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert13
timestamp 1700315010
transform 1 0 5210 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert14
timestamp 1700315010
transform -1 0 3850 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert16
timestamp 1700315010
transform -1 0 4050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert17
timestamp 1700315010
transform 1 0 2550 0 1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert19
timestamp 1700315010
transform 1 0 3050 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert20
timestamp 1700315010
transform -1 0 2450 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert22
timestamp 1700315010
transform -1 0 4230 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert23
timestamp 1700315010
transform 1 0 4270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert25
timestamp 1700315010
transform -1 0 2370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert26
timestamp 1700315010
transform -1 0 2670 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert28
timestamp 1700315010
transform 1 0 3190 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert29
timestamp 1700315010
transform -1 0 2210 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert31
timestamp 1700315010
transform -1 0 2230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert32
timestamp 1700315010
transform 1 0 3530 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert34
timestamp 1700315010
transform -1 0 6030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert35
timestamp 1700315010
transform -1 0 4970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert36
timestamp 1700315010
transform -1 0 5970 0 1 5470
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert9
timestamp 1700315010
transform -1 0 4970 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert10
timestamp 1700315010
transform -1 0 5830 0 1 790
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert12
timestamp 1700315010
transform -1 0 4990 0 -1 1310
box -12 -8 32 272
<< labels >>
flabel metal1 s 6143 2 6203 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 3336 6296 3344 6304 3 FreeSans 16 90 0 0 ABCmd_i[7]
port 2 nsew
flabel metal2 s 4856 6296 4864 6304 3 FreeSans 16 90 0 0 ABCmd_i[6]
port 3 nsew
flabel metal2 s 4956 6296 4964 6304 3 FreeSans 16 90 0 0 ABCmd_i[5]
port 4 nsew
flabel metal2 s 5116 6296 5124 6304 3 FreeSans 16 90 0 0 ABCmd_i[4]
port 5 nsew
flabel metal2 s 5816 6296 5824 6304 3 FreeSans 16 90 0 0 ABCmd_i[3]
port 6 nsew
flabel metal3 s 6176 5436 6184 5444 3 FreeSans 16 0 0 0 ABCmd_i[2]
port 7 nsew
flabel metal3 s 6176 5376 6184 5384 3 FreeSans 16 0 0 0 ABCmd_i[1]
port 8 nsew
flabel metal3 s 6176 5336 6184 5344 3 FreeSans 16 0 0 0 ABCmd_i[0]
port 9 nsew
flabel metal2 s 4656 -24 4664 -16 7 FreeSans 16 270 0 0 ACC_o[7]
port 10 nsew
flabel metal2 s 5036 -24 5044 -16 7 FreeSans 16 270 0 0 ACC_o[6]
port 11 nsew
flabel metal2 s 5396 -24 5404 -16 7 FreeSans 16 270 0 0 ACC_o[5]
port 12 nsew
flabel metal2 s 5536 -24 5544 -16 7 FreeSans 16 270 0 0 ACC_o[4]
port 13 nsew
flabel metal2 s 5676 -24 5684 -16 7 FreeSans 16 270 0 0 ACC_o[3]
port 14 nsew
flabel metal3 s -24 1176 -16 1184 7 FreeSans 16 0 0 0 ACC_o[2]
port 15 nsew
flabel metal3 s -24 2216 -16 2224 7 FreeSans 16 0 0 0 ACC_o[1]
port 16 nsew
flabel metal3 s -24 2256 -16 2264 7 FreeSans 16 0 0 0 ACC_o[0]
port 17 nsew
flabel metal2 s 5796 -24 5804 -16 7 FreeSans 16 270 0 0 Done_o
port 18 nsew
flabel metal2 s 5936 6296 5944 6304 3 FreeSans 16 90 0 0 LoadA_i
port 19 nsew
flabel metal2 s 5896 6296 5904 6304 3 FreeSans 16 90 0 0 LoadB_i
port 20 nsew
flabel metal2 s 5856 6296 5864 6304 3 FreeSans 16 90 0 0 LoadCmd_i
port 21 nsew
flabel metal3 s 6176 916 6184 924 3 FreeSans 16 0 0 0 clk
port 22 nsew
flabel metal3 s 6176 1436 6184 1444 3 FreeSans 16 0 0 0 reset
port 23 nsew
<< properties >>
string FIXED_BBOX -40 -40 6180 6300
<< end >>
