magic
tech scmos
magscale 1 2
timestamp 1726561449
<< nwell >>
rect -12 154 152 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 48 14 52 54
rect 68 14 72 54
rect 78 14 82 54
rect 100 14 104 54
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 50 166 54 246
rect 70 166 74 246
rect 78 166 82 246
rect 100 166 104 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 48 40 54
rect 24 14 26 48
rect 38 14 40 48
rect 44 14 48 54
rect 52 50 68 54
rect 52 14 54 50
rect 66 14 68 50
rect 72 14 78 54
rect 82 48 100 54
rect 82 14 84 48
rect 96 14 100 48
rect 104 14 106 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 180 26 246
rect 38 180 40 246
rect 24 166 40 180
rect 44 166 50 246
rect 54 166 56 246
rect 68 166 70 246
rect 74 166 78 246
rect 82 180 84 246
rect 98 180 100 246
rect 82 166 100 180
rect 104 166 106 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 48
rect 54 14 66 50
rect 84 14 96 48
rect 106 14 118 54
<< pdcontact >>
rect 6 166 18 246
rect 26 180 38 246
rect 56 166 68 246
rect 84 180 98 246
rect 106 166 118 246
<< psubstratepcontact >>
rect -6 -6 146 6
<< nsubstratencontact >>
rect -6 254 146 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 50 246 54 250
rect 70 246 74 250
rect 78 246 82 250
rect 100 246 104 250
rect 20 102 24 166
rect 40 162 44 166
rect 34 158 44 162
rect 34 130 39 158
rect 50 150 54 166
rect 59 138 62 150
rect 34 118 38 130
rect 34 104 40 118
rect 17 90 24 102
rect 20 54 24 90
rect 29 100 40 104
rect 29 62 33 100
rect 58 96 62 138
rect 70 116 74 166
rect 78 160 82 166
rect 100 160 104 166
rect 78 156 104 160
rect 70 104 72 116
rect 58 92 72 96
rect 29 58 44 62
rect 40 54 44 58
rect 48 54 52 72
rect 68 54 72 92
rect 100 62 104 156
rect 78 58 104 62
rect 78 54 82 58
rect 100 54 104 58
rect 20 10 24 14
rect 40 10 44 14
rect 48 10 52 14
rect 68 10 72 14
rect 78 10 82 14
rect 100 10 104 14
<< polycontact >>
rect 47 138 59 150
rect 38 118 50 130
rect 5 90 17 102
rect 72 104 84 116
rect 41 72 53 84
rect 104 116 116 128
<< metal1 >>
rect -6 266 146 268
rect -6 252 146 254
rect 26 246 38 252
rect 84 246 98 252
rect 18 166 24 172
rect 6 164 24 166
rect 68 166 78 172
rect 24 152 59 158
rect 47 150 59 152
rect 70 136 78 166
rect 98 166 106 174
rect 17 90 38 98
rect 6 60 21 70
rect 6 54 16 60
rect 59 50 65 132
rect 88 60 102 62
rect 88 54 118 60
rect 26 8 38 14
rect 84 8 96 14
rect -6 6 146 8
rect -6 -8 146 -6
<< m2contact >>
rect 24 158 38 172
rect 84 160 98 174
rect 3 102 17 116
rect 38 104 52 118
rect 38 84 52 98
rect 21 60 35 74
rect 65 122 79 136
rect 71 90 85 104
rect 103 102 117 116
rect 65 64 79 78
rect 88 62 102 76
<< metal2 >>
rect 6 116 14 134
rect 26 74 32 158
rect 66 136 74 154
rect 91 116 97 160
rect 52 110 97 116
rect 52 90 71 98
rect 91 76 97 110
rect 106 86 114 102
rect 66 46 74 64
<< m1p >>
rect -6 252 146 268
rect -6 -8 146 8
<< m2p >>
rect 66 138 74 154
rect 6 118 14 134
rect 106 86 114 100
rect 66 46 74 62
<< labels >>
rlabel metal1 -6 252 126 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 126 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal2 10 130 10 130 1 A
port 1 n signal input
rlabel metal2 70 150 70 150 1 Y
port 3 n signal output
rlabel metal2 70 50 70 50 1 Y
port 3 n signal output
rlabel metal2 110 90 110 90 5 B
port 2 n signal input
<< properties >>
string FIXED_BBOX 0 0 140 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
