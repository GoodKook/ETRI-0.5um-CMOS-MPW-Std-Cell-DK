** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/NAND2X1_TB.sch
**.subckt NAND2X1_TB
Vdd VDD GND 5
VAin A GND pwl(0 0 5n 0 6n 5 15n 5 16n 0 20n 0 21n 5 25n 5 26n 0 30n 0 31n 5 40n 5 41n 0)
R1 VDD Y 1Mega m=1
x1 B A Y VDD GND NAND2X1
VBin B GND pwl(0 0 5n 0 6n 5 15n 5 16n 0 20n 0 21n 5 35n 5 36n 0)
**** begin user architecture code



.include ~/ETRI050_DesignKit/tech/05cmos_model_240201.lib
.tran 0.01 50n
*.dc VAin 0 5 0.01
.save all



**** end user architecture code
**.ends

* expanding   symbol:  /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/NAND2X1.sym # of pins=5
** sym_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/NAND2X1.sym
** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-4_StdCell_DFFSR/Sch/NAND2X1.sch
.subckt NAND2X1 B A Y vdd gnd
*.ipin A
*.ipin B
*.opin Y
*.iopin vdd
*.iopin gnd
M1 Y A net1 GND nfet w=6u l=0.6u m=1
M2 Y A vdd VDD pfet w=6u l=0.6u m=1
M3 net1 B gnd GND nfet w=6u l=0.6u m=1
M4 Y B vdd VDD pfet w=6u l=0.6u m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
