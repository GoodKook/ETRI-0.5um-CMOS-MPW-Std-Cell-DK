magic
tech scmos
magscale 1 2
timestamp 1727572430
<< nwell >>
rect -12 194 492 273
<< ntransistor >>
rect 24 14 28 54
rect 36 14 40 54
rect 60 14 64 54
rect 72 14 76 54
rect 122 14 126 34
rect 142 14 146 34
rect 162 14 166 34
rect 212 14 216 34
rect 232 14 236 34
rect 276 14 280 34
rect 296 14 300 34
rect 350 14 354 54
rect 362 14 366 54
rect 384 14 388 54
rect 396 14 400 54
rect 444 14 448 34
<< ptransistor >>
rect 22 206 26 246
rect 42 206 46 246
rect 62 206 66 246
rect 82 206 86 246
rect 126 226 130 246
rect 146 226 150 246
rect 166 206 170 246
rect 212 206 216 246
rect 232 206 236 246
rect 276 226 280 246
rect 296 226 300 246
rect 340 206 344 246
rect 360 206 364 246
rect 380 206 384 246
rect 400 206 404 246
rect 444 206 448 246
<< ndiffusion >>
rect 20 14 24 54
rect 28 14 36 54
rect 40 14 44 54
rect 56 14 60 54
rect 64 14 72 54
rect 76 14 80 54
rect 120 14 122 34
rect 126 14 128 34
rect 140 14 142 34
rect 146 14 148 34
rect 160 14 162 34
rect 166 14 168 34
rect 210 14 212 34
rect 216 14 218 34
rect 230 14 232 34
rect 236 14 238 34
rect 274 14 276 34
rect 280 14 282 34
rect 294 14 296 34
rect 300 14 302 34
rect 346 14 350 54
rect 354 14 362 54
rect 366 14 368 54
rect 380 14 384 54
rect 388 14 396 54
rect 400 14 404 54
rect 442 14 444 34
rect 448 14 450 34
<< pdiffusion >>
rect 20 206 22 246
rect 26 206 28 246
rect 40 206 42 246
rect 46 206 48 246
rect 60 206 62 246
rect 66 206 68 246
rect 80 206 82 246
rect 86 214 88 246
rect 124 226 126 246
rect 130 226 132 246
rect 144 226 146 246
rect 150 226 152 246
rect 164 226 166 246
rect 86 206 96 214
rect 154 206 166 226
rect 170 206 172 246
rect 210 206 212 246
rect 216 206 218 246
rect 230 206 232 246
rect 236 206 238 246
rect 274 226 276 246
rect 280 226 282 246
rect 294 226 296 246
rect 300 226 302 246
rect 338 206 340 246
rect 344 206 346 246
rect 358 206 360 246
rect 364 206 366 246
rect 378 206 380 246
rect 384 206 386 246
rect 398 206 400 246
rect 404 206 406 246
rect 442 206 444 246
rect 448 206 450 246
<< ndcontact >>
rect 8 14 20 54
rect 44 14 56 54
rect 80 14 92 54
rect 108 14 120 34
rect 128 14 140 34
rect 148 14 160 34
rect 168 14 180 34
rect 198 14 210 34
rect 218 14 230 34
rect 238 14 250 34
rect 262 14 274 34
rect 282 14 294 34
rect 302 14 314 34
rect 334 14 346 54
rect 368 14 380 54
rect 404 14 416 54
rect 430 14 442 34
rect 450 14 462 34
<< pdcontact >>
rect 8 206 20 246
rect 28 206 40 246
rect 48 206 60 246
rect 68 206 80 246
rect 88 214 100 246
rect 112 226 124 246
rect 132 226 144 246
rect 152 226 164 246
rect 172 206 184 246
rect 198 206 210 246
rect 218 206 230 246
rect 238 206 250 246
rect 262 226 274 246
rect 282 226 294 246
rect 302 226 314 246
rect 326 206 338 246
rect 346 206 358 246
rect 366 206 378 246
rect 386 206 398 246
rect 406 206 418 246
rect 430 206 442 246
rect 450 206 462 246
<< psubstratepcontact >>
rect -6 -6 486 6
<< nsubstratencontact >>
rect -6 254 486 266
<< polysilicon >>
rect 22 246 26 250
rect 42 246 46 250
rect 62 246 66 250
rect 82 246 86 250
rect 126 246 130 250
rect 146 246 150 250
rect 166 246 170 250
rect 212 246 216 250
rect 232 246 236 250
rect 276 246 280 250
rect 296 246 300 250
rect 340 246 344 250
rect 360 246 364 250
rect 380 246 384 250
rect 400 246 404 250
rect 444 246 448 250
rect 22 117 26 206
rect 42 188 46 206
rect 22 105 24 117
rect 24 54 28 105
rect 44 72 48 176
rect 62 172 66 206
rect 36 54 40 60
rect 60 54 64 160
rect 82 137 86 206
rect 82 84 86 125
rect 126 116 130 226
rect 127 104 130 116
rect 146 132 150 226
rect 146 96 150 120
rect 72 80 86 84
rect 122 90 150 96
rect 166 91 170 206
rect 212 142 216 206
rect 232 166 236 206
rect 276 191 280 226
rect 256 179 280 191
rect 232 160 264 166
rect 212 132 231 142
rect 72 54 76 80
rect 122 34 126 90
rect 142 34 146 70
rect 162 34 166 79
rect 212 54 216 132
rect 260 116 264 160
rect 232 112 264 116
rect 232 80 236 112
rect 276 110 280 179
rect 296 144 300 226
rect 340 188 344 206
rect 300 132 314 138
rect 276 104 300 110
rect 192 46 216 54
rect 212 34 216 46
rect 232 34 236 68
rect 276 34 280 66
rect 296 34 300 104
rect 308 78 314 132
rect 328 84 334 188
rect 360 166 364 206
rect 380 200 384 206
rect 344 160 364 166
rect 344 134 350 160
rect 380 150 384 188
rect 400 160 404 206
rect 370 144 384 150
rect 328 78 338 84
rect 332 62 338 78
rect 344 70 350 122
rect 370 90 374 144
rect 400 102 404 148
rect 372 78 374 90
rect 344 66 366 70
rect 332 58 354 62
rect 350 54 354 58
rect 362 54 366 66
rect 370 62 374 78
rect 380 98 404 102
rect 380 70 384 98
rect 444 88 448 206
rect 404 78 448 88
rect 380 66 400 70
rect 370 58 388 62
rect 384 54 388 58
rect 396 54 400 66
rect 444 34 448 78
rect 24 10 28 14
rect 36 10 40 14
rect 60 10 64 14
rect 72 10 76 14
rect 122 10 126 14
rect 142 10 146 14
rect 162 10 166 14
rect 212 10 216 14
rect 232 10 236 14
rect 276 10 280 14
rect 296 10 300 14
rect 350 10 354 14
rect 362 10 366 14
rect 384 10 388 14
rect 396 10 400 14
rect 444 10 448 14
<< polycontact >>
rect 38 176 50 188
rect 24 105 36 117
rect 36 60 48 72
rect 60 160 72 172
rect 77 125 89 137
rect 115 104 127 116
rect 146 120 158 132
rect 244 179 256 191
rect 231 132 243 144
rect 142 70 154 82
rect 162 79 174 91
rect 288 132 300 144
rect 328 188 340 200
rect 224 68 236 80
rect 180 42 192 54
rect 276 66 288 78
rect 372 188 384 200
rect 392 148 404 160
rect 344 122 356 134
rect 308 66 320 78
rect 360 78 372 90
rect 392 78 404 90
<< metal1 >>
rect -6 266 486 268
rect -6 252 486 254
rect 8 246 20 252
rect 48 246 60 252
rect 88 246 100 252
rect 172 246 184 252
rect 218 246 230 252
rect 326 246 338 252
rect 366 246 378 252
rect 406 246 418 252
rect 450 246 462 252
rect 109 226 112 246
rect 130 226 132 246
rect 151 226 152 246
rect 109 208 115 226
rect 130 208 137 226
rect 151 208 159 226
rect 28 200 35 206
rect 8 194 35 200
rect 8 86 16 194
rect 68 186 80 206
rect 198 196 210 206
rect 50 178 166 186
rect 198 182 203 196
rect 289 200 296 212
rect 346 200 358 206
rect 289 192 328 200
rect 236 191 250 192
rect 236 179 244 191
rect 346 192 372 200
rect 158 173 166 178
rect 72 160 123 168
rect 158 166 263 173
rect 390 172 398 206
rect 317 166 416 172
rect 158 152 392 160
rect 77 148 89 149
rect 158 148 166 152
rect 77 142 166 148
rect 77 137 89 142
rect 24 117 36 123
rect 95 122 140 129
rect 95 113 103 122
rect 36 105 103 113
rect 133 112 140 122
rect 158 124 217 132
rect 294 124 300 132
rect 203 118 300 124
rect 322 122 344 134
rect 374 123 383 137
rect 322 112 328 122
rect 133 104 328 112
rect 374 104 382 123
rect 8 78 110 86
rect 8 54 16 78
rect 48 60 92 68
rect 82 54 92 60
rect 103 54 110 78
rect 120 70 127 104
rect 174 83 183 91
rect 336 96 382 104
rect 336 94 346 96
rect 224 84 346 94
rect 224 80 236 84
rect 120 62 186 70
rect 352 78 360 88
rect 372 78 392 88
rect 288 66 308 78
rect 180 54 186 62
rect 352 54 362 78
rect 410 54 416 166
rect 115 40 117 54
rect 108 34 117 40
rect 128 34 137 40
rect 148 34 159 40
rect 203 34 210 40
rect 239 34 250 40
rect 262 34 274 40
rect 283 34 294 40
rect 305 34 314 40
rect 346 46 362 54
rect 430 137 440 206
rect 430 123 443 137
rect 430 34 440 123
rect 44 8 56 14
rect 168 8 180 14
rect 218 8 230 14
rect 368 8 380 14
rect 450 8 462 14
rect -6 6 486 8
rect -6 -8 486 -6
<< m2contact >>
rect 101 194 115 208
rect 123 194 137 208
rect 145 194 159 208
rect 260 212 274 226
rect 282 212 296 226
rect 305 212 319 226
rect 203 182 217 196
rect 236 192 250 206
rect 123 158 137 172
rect 263 166 277 180
rect 303 166 317 180
rect 23 123 37 137
rect 63 123 77 137
rect 203 132 217 146
rect 243 132 257 146
rect 383 123 397 137
rect 183 83 197 97
rect 101 40 115 54
rect 123 40 137 54
rect 145 40 159 54
rect 203 40 217 54
rect 239 40 253 54
rect 261 40 275 54
rect 283 40 297 54
rect 305 40 319 54
rect 443 123 457 137
<< metal2 >>
rect 23 137 37 157
rect 63 103 77 123
rect 106 54 114 194
rect 126 172 134 194
rect 129 54 137 158
rect 149 54 157 194
rect 250 192 251 206
rect 203 146 211 182
rect 243 146 251 192
rect 266 180 274 212
rect 289 192 296 212
rect 183 97 197 117
rect 207 54 215 132
rect 243 54 251 132
rect 265 54 275 166
rect 289 54 297 192
rect 305 180 313 212
rect 305 54 313 166
rect 383 103 397 123
rect 443 103 457 123
<< m2p >>
rect 23 143 37 157
rect 63 103 77 117
rect 183 103 197 117
rect 383 103 397 117
rect 443 103 457 117
<< labels >>
rlabel metal2 23 143 37 157 0 R
port 0 nsew signal input
rlabel metal2 63 103 77 117 0 S
port 1 nsew signal input
rlabel metal2 183 103 197 117 0 D
port 2 nsew signal input
rlabel metal2 383 103 397 117 0 CLK
port 3 nsew clock input
rlabel metal2 443 103 457 117 0 Q
port 4 nsew signal output
rlabel metal1 -6 252 486 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 486 8 0 gnd
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 480 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
