magic
tech scmos
magscale 1 30
timestamp 1741148510
<< checkpaint >>
rect -1337 -644 15289 26875
rect -1200 -705 13595 -644
rect -1200 -9750 12700 -705
rect -1200 -12610 11490 -9750
<< metal3 >>
rect 0 23400 12000 25060
rect 0 21100 12000 22760
rect 0 11300 12000 19100
rect 0 0 12000 7800
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 6500 0 1 0
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1569139307
transform 1 0 500 0 1 0
box -35 0 5035 25060
use pad80_CDNS_704676826050  pad80_CDNS_704676826050_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 1750 0 1 -9150
box 0 0 8500 8500
<< end >>
