magic
tech scmos
magscale 1 2
timestamp 1726483455
<< nwell >>
rect -12 154 292 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
rect 100 14 104 54
rect 120 14 124 54
rect 140 14 144 54
rect 160 14 164 54
rect 180 14 184 54
rect 200 14 204 54
rect 220 14 224 54
rect 240 14 244 54
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 60 166 64 246
rect 80 166 84 246
rect 100 166 104 246
rect 120 166 124 246
rect 140 166 144 246
rect 160 166 164 246
rect 180 166 184 246
rect 200 166 204 246
rect 220 166 224 246
rect 240 166 244 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 26 54
rect 38 14 40 54
rect 44 14 46 54
rect 58 14 60 54
rect 64 14 66 54
rect 78 14 80 54
rect 84 14 86 54
rect 98 14 100 54
rect 104 14 106 54
rect 118 14 120 54
rect 124 14 126 54
rect 138 14 140 54
rect 144 14 146 54
rect 158 14 160 54
rect 164 14 166 54
rect 178 14 180 54
rect 184 14 186 54
rect 198 14 200 54
rect 204 14 206 54
rect 218 14 220 54
rect 224 14 226 54
rect 238 14 240 54
rect 244 14 246 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 26 246
rect 38 166 40 246
rect 44 166 46 246
rect 58 166 60 246
rect 64 166 66 246
rect 78 166 80 246
rect 84 166 86 246
rect 98 166 100 246
rect 104 166 106 246
rect 118 166 120 246
rect 124 166 126 246
rect 138 166 140 246
rect 144 166 146 246
rect 158 166 160 246
rect 164 166 166 246
rect 178 166 180 246
rect 184 166 186 246
rect 198 166 200 246
rect 204 166 206 246
rect 218 166 220 246
rect 224 166 226 246
rect 238 166 240 246
rect 244 166 246 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 54
rect 46 14 58 54
rect 66 14 78 54
rect 86 14 98 54
rect 106 14 118 54
rect 126 14 138 54
rect 146 14 158 54
rect 166 14 178 54
rect 186 14 198 54
rect 206 14 218 54
rect 226 14 238 54
rect 246 14 258 54
<< pdcontact >>
rect 6 166 18 246
rect 26 166 38 246
rect 46 166 58 246
rect 66 166 78 246
rect 86 166 98 246
rect 106 166 118 246
rect 126 166 138 246
rect 146 166 158 246
rect 166 166 178 246
rect 186 166 198 246
rect 206 166 218 246
rect 226 166 238 246
rect 246 166 258 246
<< psubstratepcontact >>
rect -6 -6 286 6
<< nsubstratencontact >>
rect -6 254 286 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 80 246 84 250
rect 100 246 104 250
rect 120 246 124 250
rect 140 246 144 250
rect 160 246 164 250
rect 180 246 184 250
rect 200 246 204 250
rect 220 246 224 250
rect 240 246 244 250
rect 20 54 24 166
rect 40 103 44 166
rect 36 91 44 103
rect 40 54 44 91
rect 60 86 64 166
rect 80 82 84 166
rect 72 74 84 82
rect 60 54 64 74
rect 80 54 84 74
rect 100 86 104 166
rect 120 82 124 166
rect 112 74 124 82
rect 100 54 104 74
rect 120 54 124 74
rect 140 86 144 166
rect 160 82 164 166
rect 152 74 164 82
rect 140 54 144 74
rect 160 54 164 74
rect 180 86 184 166
rect 200 82 204 166
rect 192 74 204 82
rect 180 54 184 74
rect 200 54 204 74
rect 220 86 224 166
rect 240 82 244 166
rect 232 74 244 82
rect 220 54 224 74
rect 240 54 244 74
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
rect 100 10 104 14
rect 120 10 124 14
rect 140 10 144 14
rect 160 10 164 14
rect 180 10 184 14
rect 200 10 204 14
rect 220 10 224 14
rect 240 10 244 14
<< polycontact >>
rect 24 91 36 103
rect 60 74 72 86
rect 100 74 112 86
rect 140 74 152 86
rect 180 74 192 86
rect 220 74 232 86
<< metal1 >>
rect -6 266 286 268
rect -6 252 286 254
rect 6 246 18 252
rect 46 246 58 252
rect 86 246 98 252
rect 126 246 138 252
rect 166 246 178 252
rect 206 246 218 252
rect 246 246 258 252
rect 26 160 38 166
rect 66 160 78 166
rect 106 160 118 166
rect 146 160 158 166
rect 186 160 198 166
rect 226 160 238 166
rect 26 152 53 160
rect 66 152 92 160
rect 106 152 132 160
rect 146 152 174 160
rect 186 152 208 160
rect 226 152 248 160
rect 45 82 53 152
rect 45 74 60 82
rect 84 82 92 152
rect 84 74 100 82
rect 124 82 132 152
rect 124 74 140 82
rect 166 82 174 152
rect 166 74 180 82
rect 200 82 208 152
rect 240 117 248 152
rect 240 103 243 117
rect 200 74 220 82
rect 45 68 53 74
rect 84 68 92 74
rect 124 68 132 74
rect 166 68 174 74
rect 200 68 208 74
rect 240 68 248 103
rect 26 60 53 68
rect 66 60 92 68
rect 106 60 132 68
rect 146 60 174 68
rect 186 60 208 68
rect 226 60 248 68
rect 26 54 38 60
rect 66 54 78 60
rect 106 54 118 60
rect 146 54 158 60
rect 186 54 198 60
rect 226 54 238 60
rect 6 8 18 14
rect 46 8 58 14
rect 86 8 98 14
rect 126 8 138 14
rect 166 8 178 14
rect 206 8 218 14
rect 246 8 258 14
rect -6 6 286 8
rect -6 -8 286 -6
<< m2contact >>
rect 23 103 37 117
rect 243 103 257 117
<< metal2 >>
rect 26 117 34 134
rect 246 117 254 134
<< m1p >>
rect -6 252 286 268
rect -6 -8 286 8
<< m2p >>
rect 26 119 34 134
rect 246 119 254 134
<< labels >>
rlabel metal1 -6 252 266 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 266 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal2 30 131 30 131 3 A
port 1 n signal input
rlabel metal2 250 131 250 131 7 Y
port 2 n signal output
<< properties >>
string FIXED_BBOX 0 0 280 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
