magic
tech scmos
magscale 1 6
timestamp 1537935238
<< checkpaint >>
rect -120 -208 1608 960
<< nwell >>
rect 647 -20 1488 648
<< psubstratepdiff >>
rect 0 756 512 792
rect 0 198 40 756
rect 472 198 512 756
rect 0 162 512 198
<< nsubstratendiff >>
rect 667 592 1469 628
rect 667 36 707 592
rect 1429 36 1469 592
rect 667 0 1469 36
<< metal1 >>
rect 0 756 512 792
rect 0 198 40 756
rect 116 698 392 738
rect 142 254 186 274
rect 262 254 306 274
rect 382 254 424 274
rect 142 214 424 254
rect 472 198 512 756
rect 0 162 512 198
rect 667 592 1469 628
rect 667 36 707 592
rect 777 536 1353 576
rect 745 92 787 112
rect 863 92 907 112
rect 983 92 1027 112
rect 1103 92 1147 112
rect 1223 92 1267 112
rect 1343 92 1385 112
rect 745 52 1385 92
rect 1429 36 1469 592
rect 667 0 1469 36
<< metal2 >>
rect 0 162 40 792
rect 226 738 290 840
rect 116 698 1140 738
rect 84 274 126 678
rect 202 274 246 678
rect 322 274 366 678
rect 172 -20 356 254
rect 472 162 512 678
rect 667 0 707 628
rect 1044 576 1140 698
rect 777 536 1353 576
rect 805 112 847 516
rect 923 112 967 516
rect 1043 112 1085 516
rect 1161 112 1205 516
rect 1283 112 1325 516
rect 745 -20 1385 92
rect 1429 0 1469 628
rect 172 -88 1385 -20
<< metal3 >>
rect 0 460 40 792
rect 84 460 126 678
rect 202 460 246 678
rect 322 460 366 678
rect 472 460 512 792
rect 667 0 707 332
rect 805 112 847 332
rect 923 112 967 332
rect 1043 111 1085 331
rect 1161 112 1205 332
rect 1283 112 1325 332
rect 1429 0 1469 332
use CONT  CONT_0
array 0 17 24 0 0 0
timestamp 1537935238
transform 1 0 47 0 1 774
box -6 -6 6 6
use CONT  CONT_1
array 0 0 0 0 10 56
timestamp 1537935238
transform 1 0 492 0 1 210
box -6 -6 6 6
use CONT  CONT_2
array 0 0 0 0 10 56
timestamp 1537935238
transform 1 0 687 0 1 24
box -6 -6 6 6
use CONT  CONT_3
array 0 0 0 0 10 56
timestamp 1537935238
transform 1 0 20 0 1 206
box -6 -6 6 6
use CONT  CONT_4
array 0 0 0 0 10 56
timestamp 1537935238
transform 1 0 1449 0 1 24
box -6 -6 6 6
use CONT  CONT_5
array 0 17 24 0 0 0
timestamp 1537935238
transform 1 0 47 0 1 180
box -6 -6 6 6
use CONT  CONT_6
array 0 12 56 0 0 0
timestamp 1537935238
transform 1 0 723 0 1 610
box -6 -6 6 6
use CONT  CONT_7
array 0 12 56 0 0 0
timestamp 1537935238
transform 1 0 723 0 1 18
box -6 -6 6 6
use NCELL1  NCELL1_0
array 0 4 60 0 0 0
timestamp 1537935238
transform -1 0 422 0 -1 676
box -2 -58 98 410
use PCELL1  PCELL1_0
array 0 9 60 0 0 0
timestamp 1537935238
transform -1 0 1383 0 -1 514
box -2 -58 98 410
use VIA1  VIA1_0
array 0 0 0 0 9 56
timestamp 1537935238
transform 1 0 1449 0 1 52
box -8 -8 8 8
use VIA1  VIA1_1
array 0 13 44 0 0 0
timestamp 1537935238
transform 1 0 766 0 1 72
box -8 -8 8 8
use VIA1  VIA1_2
array 0 4 36 0 0 0
timestamp 1537935238
transform 1 0 192 0 1 234
box -8 -8 8 8
use VIA1  VIA1_3
array 0 0 0 0 7 56
timestamp 1537935238
transform 1 0 492 0 1 238
box -8 -8 8 8
use VIA1  VIA1_4
array 0 2 120 0 5 56
timestamp 1537935238
transform 1 0 104 0 1 348
box -8 -8 8 8
use VIA1  VIA1_5
array 0 8 60 0 0 0
timestamp 1537935238
transform 1 0 825 0 1 556
box -8 -8 8 8
use VIA1  VIA1_6
array 0 3 60 0 0 0
timestamp 1537935238
transform 1 0 164 0 1 718
box -8 -8 8 8
use VIA1  VIA1_7
array 0 4 120 0 5 56
timestamp 1537935238
transform 1 0 825 0 1 186
box -8 -8 8 8
use VIA1  VIA1_8
array 0 0 0 0 9 56
timestamp 1537935238
transform 1 0 20 0 1 234
box -8 -8 8 8
use VIA1  VIA1_9
array 0 0 0 0 9 56
timestamp 1537935238
transform 1 0 687 0 1 52
box -8 -8 8 8
use VIA2  VIA2_0
array 0 0 0 0 5 56
timestamp 1537935238
transform 1 0 1449 0 1 24
box -8 -8 8 8
use VIA2  VIA2_1
array 0 0 0 0 4 56
timestamp 1537935238
transform 1 0 687 0 1 24
box -8 -8 8 8
use VIA2  VIA2_2
array 0 2 120 0 3 56
timestamp 1537935238
transform 1 0 104 0 1 488
box -8 -8 8 8
use VIA2  VIA2_3
array 0 4 120 0 2 56
timestamp 1537935238
transform 1 0 825 0 1 158
box -8 -8 8 8
use VIA2  VIA2_4
array 0 0 0 0 3 56
timestamp 1537935238
transform 1 0 492 0 1 490
box -8 -8 8 8
use VIA2  VIA2_5
array 0 0 0 0 5 56
timestamp 1537935238
transform 1 0 20 0 1 486
box -8 -8 8 8
<< end >>
