magic
tech scmos
timestamp 1702508443
<< nwell >>
rect -6 77 46 136
<< ntransistor >>
rect 9 7 11 37
rect 14 7 16 37
rect 21 7 23 37
<< ptransistor >>
rect 9 103 11 123
rect 19 103 21 123
rect 29 103 31 123
<< ndiffusion >>
rect 8 7 9 37
rect 11 7 14 37
rect 16 7 21 37
rect 23 36 30 37
rect 23 7 24 36
<< pdiffusion >>
rect 8 103 9 123
rect 11 103 12 123
rect 18 103 19 123
rect 21 105 22 123
rect 28 105 29 123
rect 21 103 29 105
rect 31 103 32 123
<< ndcontact >>
rect 2 7 8 37
rect 24 7 30 36
<< pdcontact >>
rect 2 103 8 123
rect 12 103 18 123
rect 22 105 28 123
rect 32 103 38 123
<< psubstratepcontact >>
rect -3 -3 43 3
<< nsubstratencontact >>
rect -3 127 43 133
<< polysilicon >>
rect 9 123 11 125
rect 19 123 21 125
rect 29 123 31 125
rect 9 97 11 103
rect 19 102 21 103
rect 5 95 11 97
rect 14 100 21 102
rect 5 51 8 95
rect 14 64 16 100
rect 5 40 8 45
rect 5 38 11 40
rect 9 37 11 38
rect 14 37 16 58
rect 29 51 31 103
rect 28 45 31 51
rect 26 40 28 45
rect 21 38 28 40
rect 21 37 23 38
rect 9 5 11 7
rect 14 5 16 7
rect 21 5 23 7
<< polycontact >>
rect 12 58 18 64
rect 2 45 8 51
rect 22 45 28 51
<< metal1 >>
rect -3 133 43 134
rect -3 126 43 127
rect 2 123 8 126
rect 22 123 28 126
rect 13 102 18 103
rect 32 102 35 103
rect 13 99 35 102
rect 32 58 35 99
rect 32 39 35 51
rect 24 36 35 39
rect 30 35 35 36
rect 2 4 8 7
rect -3 3 43 4
rect -3 -4 43 -3
<< m2contact >>
rect 1 51 8 58
rect 11 51 18 58
rect 21 51 28 58
rect 31 51 38 58
<< metal2 >>
rect 3 58 7 67
rect 23 58 27 67
rect 13 43 17 51
rect 33 43 37 51
<< m1p >>
rect -3 126 43 134
rect -3 -4 43 4
<< m2p >>
rect 3 59 7 67
rect 23 59 27 67
rect 13 43 17 50
rect 33 43 37 50
<< labels >>
rlabel metal2 5 65 5 65 1 A
port 1 n signal input
rlabel metal2 15 45 15 45 5 B
port 2 n signal input
rlabel metal2 25 65 25 65 1 C
port 3 n signal input
rlabel metal2 35 44 35 44 5 Y
port 4 n signal output
rlabel metal1 -3 126 43 134 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -3 -4 43 4 0 gnd
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 40 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
