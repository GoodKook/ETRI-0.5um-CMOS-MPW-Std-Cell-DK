VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ALU_wrapper
  CLASS BLOCK ;
  FOREIGN ALU_wrapper ;
  ORIGIN 6.000 6.000 ;
  SIZE 870.000 BY 879.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 19.500 830.700 21.300 840.600 ;
        RECT 29.700 830.700 31.500 840.600 ;
        RECT 51.000 830.700 52.800 837.600 ;
        RECT 58.500 830.700 60.300 834.600 ;
        RECT 74.400 830.700 76.200 835.800 ;
        RECT 100.800 830.700 102.600 835.800 ;
        RECT 118.800 830.700 120.600 834.600 ;
        RECT 139.500 830.700 141.300 840.600 ;
        RECT 152.400 830.700 154.200 835.800 ;
        RECT 171.000 830.700 172.800 837.600 ;
        RECT 178.500 830.700 180.300 834.600 ;
        RECT 196.800 830.700 198.600 834.600 ;
        RECT 206.700 830.700 208.500 840.600 ;
        RECT 238.500 830.700 240.300 840.600 ;
        RECT 256.800 830.700 258.600 835.800 ;
        RECT 274.800 830.700 276.600 834.600 ;
        RECT 292.800 830.700 294.600 835.800 ;
        RECT 305.400 830.700 307.200 834.600 ;
        RECT 325.800 830.700 327.600 834.600 ;
        RECT 331.800 831.600 333.600 834.600 ;
        RECT 332.400 830.700 333.600 831.600 ;
        RECT 343.800 830.700 345.600 834.600 ;
        RECT 349.800 830.700 351.600 834.600 ;
        RECT 367.800 830.700 369.600 835.800 ;
        RECT 385.800 830.700 387.600 834.600 ;
        RECT 398.400 830.700 400.200 835.800 ;
        RECT 419.700 830.700 421.500 834.600 ;
        RECT 427.200 830.700 429.000 837.600 ;
        RECT 437.700 830.700 439.500 837.600 ;
        RECT 455.400 831.600 457.200 834.600 ;
        RECT 455.400 830.700 456.600 831.600 ;
        RECT 461.400 830.700 463.200 834.600 ;
        RECT 487.500 830.700 489.300 840.600 ;
        RECT 502.800 830.700 504.600 834.600 ;
        RECT 520.500 830.700 522.300 837.600 ;
        RECT 530.400 830.700 532.200 837.600 ;
        RECT 536.400 830.700 538.200 837.600 ;
        RECT 542.400 830.700 544.200 837.600 ;
        RECT 548.400 830.700 550.200 837.600 ;
        RECT 554.400 830.700 556.200 837.600 ;
        RECT 562.200 830.700 564.000 834.600 ;
        RECT 574.500 830.700 576.300 837.600 ;
        RECT 597.000 830.700 598.800 834.600 ;
        RECT 604.500 830.700 606.300 834.600 ;
        RECT 623.100 830.700 624.900 837.600 ;
        RECT 646.500 830.700 648.300 837.600 ;
        RECT 652.200 830.700 654.000 834.600 ;
        RECT 664.500 830.700 666.300 837.600 ;
        RECT 687.000 830.700 688.800 834.600 ;
        RECT 694.500 830.700 696.300 834.600 ;
        RECT 713.100 830.700 714.900 837.600 ;
        RECT 736.800 830.700 738.600 835.800 ;
        RECT 751.800 830.700 753.600 834.600 ;
        RECT 757.800 830.700 759.600 834.600 ;
        RECT 767.400 830.700 769.200 834.600 ;
        RECT 787.800 830.700 789.600 834.600 ;
        RECT 794.850 830.700 796.650 834.600 ;
        RECT 803.850 830.700 805.650 834.600 ;
        RECT 810.750 830.700 812.550 834.600 ;
        RECT 820.050 830.700 821.850 834.600 ;
        RECT 833.400 830.700 835.200 837.600 ;
        RECT 858.450 830.700 867.450 866.700 ;
        RECT 0.600 828.300 867.450 830.700 ;
        RECT 11.700 824.400 13.500 828.300 ;
        RECT 19.200 821.400 21.000 828.300 ;
        RECT 40.500 818.400 42.300 828.300 ;
        RECT 58.800 823.200 60.600 828.300 ;
        RECT 79.800 823.200 81.600 828.300 ;
        RECT 97.800 824.400 99.600 828.300 ;
        RECT 107.700 818.400 109.500 828.300 ;
        RECT 131.700 824.400 133.500 828.300 ;
        RECT 139.200 821.400 141.000 828.300 ;
        RECT 154.800 824.400 156.600 828.300 ;
        RECT 161.400 827.400 162.600 828.300 ;
        RECT 160.800 824.400 162.600 827.400 ;
        RECT 170.700 821.400 172.500 828.300 ;
        RECT 193.800 821.400 195.600 828.300 ;
        RECT 202.200 821.400 204.000 828.300 ;
        RECT 212.700 821.400 214.500 828.300 ;
        RECT 230.700 818.400 232.500 828.300 ;
        RECT 251.700 818.400 253.500 828.300 ;
        RECT 280.500 821.400 282.300 828.300 ;
        RECT 301.500 818.400 303.300 828.300 ;
        RECT 311.700 818.400 313.500 828.300 ;
        RECT 332.700 821.400 334.500 828.300 ;
        RECT 355.800 824.400 357.600 828.300 ;
        RECT 365.700 818.400 367.500 828.300 ;
        RECT 386.400 824.400 388.200 828.300 ;
        RECT 412.500 818.400 414.300 828.300 ;
        RECT 433.500 818.400 435.300 828.300 ;
        RECT 451.500 821.400 453.300 828.300 ;
        RECT 466.800 824.400 468.600 828.300 ;
        RECT 473.400 827.400 474.600 828.300 ;
        RECT 472.800 824.400 474.600 827.400 ;
        RECT 482.700 821.400 484.500 828.300 ;
        RECT 508.800 823.200 510.600 828.300 ;
        RECT 529.500 821.400 531.300 828.300 ;
        RECT 547.800 823.200 549.600 828.300 ;
        RECT 568.500 821.400 570.300 828.300 ;
        RECT 581.700 824.400 583.500 828.300 ;
        RECT 589.200 821.400 591.000 828.300 ;
        RECT 604.800 824.400 606.600 828.300 ;
        RECT 619.800 824.400 621.600 828.300 ;
        RECT 629.700 818.400 631.500 828.300 ;
        RECT 655.800 824.400 657.600 828.300 ;
        RECT 668.400 823.200 670.200 828.300 ;
        RECT 689.400 823.200 691.200 828.300 ;
        RECT 710.400 823.200 712.200 828.300 ;
        RECT 735.300 821.400 737.100 828.300 ;
        RECT 749.400 824.400 751.200 828.300 ;
        RECT 755.400 824.400 757.200 828.300 ;
        RECT 767.400 824.400 769.200 828.300 ;
        RECT 773.400 824.400 775.200 828.300 ;
        RECT 785.400 827.400 786.600 828.300 ;
        RECT 785.400 824.400 787.200 827.400 ;
        RECT 791.400 824.400 793.200 828.300 ;
        RECT 809.400 822.900 811.200 828.300 ;
        RECT 835.800 821.400 837.600 828.300 ;
        RECT 844.200 821.400 846.000 828.300 ;
        RECT 10.800 758.700 12.600 762.600 ;
        RECT 16.800 758.700 18.600 762.600 ;
        RECT 34.500 758.700 36.300 765.600 ;
        RECT 47.700 758.700 49.500 762.600 ;
        RECT 55.200 758.700 57.000 765.600 ;
        RECT 65.700 758.700 67.500 768.600 ;
        RECT 93.300 758.700 95.100 765.600 ;
        RECT 115.800 758.700 117.600 763.800 ;
        RECT 131.400 758.700 133.200 763.800 ;
        RECT 156.300 758.700 158.100 765.600 ;
        RECT 170.400 758.700 172.200 762.600 ;
        RECT 176.400 758.700 178.200 762.600 ;
        RECT 191.700 758.700 193.500 762.600 ;
        RECT 199.200 758.700 201.000 765.600 ;
        RECT 220.500 758.700 222.300 768.600 ;
        RECT 230.700 758.700 232.500 765.600 ;
        RECT 255.300 758.700 257.100 765.600 ;
        RECT 280.500 758.700 282.300 768.600 ;
        RECT 290.700 758.700 292.500 765.600 ;
        RECT 316.800 758.700 318.600 763.800 ;
        RECT 337.800 758.700 339.600 763.800 ;
        RECT 350.400 758.700 352.200 762.600 ;
        RECT 356.400 758.700 358.200 762.600 ;
        RECT 372.900 758.700 374.700 765.600 ;
        RECT 400.500 758.700 402.300 768.600 ;
        RECT 410.400 758.700 412.200 762.600 ;
        RECT 425.700 758.700 427.500 765.600 ;
        RECT 443.700 758.700 445.500 765.600 ;
        RECT 461.700 758.700 463.500 768.600 ;
        RECT 493.500 758.700 495.300 768.600 ;
        RECT 504.000 758.700 505.800 765.600 ;
        RECT 511.500 758.700 513.300 762.600 ;
        RECT 532.800 758.700 534.600 763.800 ;
        RECT 553.800 758.700 555.600 763.800 ;
        RECT 573.300 758.700 575.100 765.600 ;
        RECT 592.800 758.700 594.600 762.600 ;
        RECT 602.400 758.700 604.200 762.600 ;
        RECT 608.400 758.700 610.200 762.600 ;
        RECT 623.400 758.700 625.200 764.100 ;
        RECT 647.700 758.700 649.500 762.600 ;
        RECT 655.200 758.700 657.000 765.600 ;
        RECT 665.400 758.700 667.200 762.600 ;
        RECT 681.000 758.700 682.800 765.600 ;
        RECT 689.400 758.700 691.200 765.600 ;
        RECT 707.400 758.700 709.200 763.800 ;
        RECT 726.000 758.700 727.800 765.600 ;
        RECT 733.500 758.700 735.300 762.600 ;
        RECT 749.400 758.700 751.200 763.800 ;
        RECT 767.100 758.700 768.900 765.600 ;
        RECT 785.700 758.700 787.500 762.600 ;
        RECT 793.200 758.700 795.000 762.600 ;
        RECT 815.700 758.700 817.500 765.600 ;
        RECT 828.000 758.700 829.800 762.600 ;
        RECT 839.400 758.700 841.200 762.600 ;
        RECT 858.450 758.700 867.450 828.300 ;
        RECT 0.600 756.300 867.450 758.700 ;
        RECT 16.500 749.400 18.300 756.300 ;
        RECT 34.800 751.200 36.600 756.300 ;
        RECT 50.400 751.200 52.200 756.300 ;
        RECT 71.700 752.400 73.500 756.300 ;
        RECT 79.200 749.400 81.000 756.300 ;
        RECT 100.500 746.400 102.300 756.300 ;
        RECT 110.700 749.400 112.500 756.300 ;
        RECT 128.400 752.400 130.200 756.300 ;
        RECT 143.700 746.400 145.500 756.300 ;
        RECT 164.700 749.400 166.500 756.300 ;
        RECT 182.400 755.400 183.600 756.300 ;
        RECT 182.400 752.400 184.200 755.400 ;
        RECT 188.400 752.400 190.200 756.300 ;
        RECT 211.500 749.400 213.300 756.300 ;
        RECT 223.800 752.400 225.600 756.300 ;
        RECT 229.800 752.400 231.600 756.300 ;
        RECT 247.500 749.400 249.300 756.300 ;
        RECT 257.400 752.400 259.200 756.300 ;
        RECT 283.500 746.400 285.300 756.300 ;
        RECT 298.800 752.400 300.600 756.300 ;
        RECT 305.400 755.400 306.600 756.300 ;
        RECT 304.800 752.400 306.600 755.400 ;
        RECT 314.700 749.400 316.500 756.300 ;
        RECT 332.400 752.400 334.200 756.300 ;
        RECT 338.400 752.400 340.200 756.300 ;
        RECT 358.800 751.200 360.600 756.300 ;
        RECT 371.400 752.400 373.200 756.300 ;
        RECT 391.800 752.400 393.600 756.300 ;
        RECT 401.400 752.400 403.200 756.300 ;
        RECT 407.400 752.400 409.200 756.300 ;
        RECT 419.700 749.400 421.500 756.300 ;
        RECT 445.800 751.200 447.600 756.300 ;
        RECT 458.700 749.400 460.500 756.300 ;
        RECT 484.800 751.200 486.600 756.300 ;
        RECT 502.800 752.400 504.600 756.300 ;
        RECT 523.800 750.900 525.600 756.300 ;
        RECT 536.700 749.400 538.500 756.300 ;
        RECT 556.800 749.400 558.600 756.300 ;
        RECT 562.800 749.400 564.600 756.300 ;
        RECT 572.400 752.400 574.200 756.300 ;
        RECT 578.400 752.400 580.200 756.300 ;
        RECT 590.400 752.400 592.200 756.300 ;
        RECT 596.400 752.400 598.200 756.300 ;
        RECT 616.800 751.200 618.600 756.300 ;
        RECT 629.400 752.400 631.200 756.300 ;
        RECT 649.800 752.400 651.600 756.300 ;
        RECT 659.400 752.400 661.200 756.300 ;
        RECT 665.400 752.400 667.200 756.300 ;
        RECT 677.400 752.400 679.200 756.300 ;
        RECT 683.400 752.400 685.200 756.300 ;
        RECT 703.500 749.400 705.300 756.300 ;
        RECT 710.850 752.400 712.650 756.300 ;
        RECT 719.850 752.400 721.650 756.300 ;
        RECT 726.750 752.400 728.550 756.300 ;
        RECT 736.050 752.400 737.850 756.300 ;
        RECT 749.700 749.400 751.500 756.300 ;
        RECT 775.800 751.200 777.600 756.300 ;
        RECT 793.800 752.400 795.600 756.300 ;
        RECT 806.700 749.400 808.500 756.300 ;
        RECT 824.400 751.200 826.200 756.300 ;
        RECT 842.700 749.400 844.500 756.300 ;
        RECT 19.500 686.700 21.300 696.600 ;
        RECT 30.000 686.700 31.800 693.600 ;
        RECT 37.500 686.700 39.300 690.600 ;
        RECT 53.400 686.700 55.200 691.800 ;
        RECT 74.400 686.700 76.200 691.800 ;
        RECT 92.700 686.700 94.500 696.600 ;
        RECT 113.700 686.700 115.500 696.600 ;
        RECT 135.000 686.700 136.800 693.600 ;
        RECT 142.500 686.700 144.300 690.600 ;
        RECT 158.400 686.700 160.200 691.800 ;
        RECT 184.500 686.700 186.300 693.600 ;
        RECT 194.700 686.700 196.500 696.600 ;
        RECT 217.800 686.700 219.600 690.600 ;
        RECT 223.800 686.700 225.600 690.600 ;
        RECT 244.500 686.700 246.300 696.600 ;
        RECT 257.400 686.700 259.200 692.100 ;
        RECT 289.500 686.700 291.300 696.600 ;
        RECT 302.700 686.700 304.500 690.600 ;
        RECT 310.200 686.700 312.000 693.600 ;
        RECT 320.400 686.700 322.200 690.600 ;
        RECT 335.400 686.700 337.200 690.600 ;
        RECT 353.400 686.700 355.200 691.800 ;
        RECT 376.800 686.700 378.600 693.600 ;
        RECT 386.700 686.700 388.500 693.600 ;
        RECT 415.800 686.700 417.600 692.100 ;
        RECT 436.500 686.700 438.300 693.600 ;
        RECT 446.400 687.600 448.200 690.600 ;
        RECT 446.400 686.700 447.600 687.600 ;
        RECT 452.400 686.700 454.200 690.600 ;
        RECT 472.800 686.700 474.600 690.600 ;
        RECT 482.700 686.700 484.500 696.600 ;
        RECT 503.700 686.700 505.500 693.600 ;
        RECT 526.800 686.700 528.600 693.600 ;
        RECT 536.400 686.700 538.200 690.600 ;
        RECT 551.400 686.700 553.200 690.600 ;
        RECT 557.400 686.700 559.200 690.600 ;
        RECT 577.500 686.700 579.300 693.600 ;
        RECT 587.400 686.700 589.200 690.600 ;
        RECT 593.400 686.700 595.200 690.600 ;
        RECT 605.400 686.700 607.200 690.600 ;
        RECT 611.400 686.700 613.200 690.600 ;
        RECT 623.700 686.700 625.500 693.600 ;
        RECT 639.150 686.700 640.950 690.600 ;
        RECT 648.450 686.700 650.250 690.600 ;
        RECT 655.350 686.700 657.150 690.600 ;
        RECT 664.350 686.700 666.150 690.600 ;
        RECT 677.700 686.700 679.500 693.600 ;
        RECT 695.400 686.700 697.200 690.600 ;
        RECT 707.850 686.700 709.650 690.600 ;
        RECT 716.850 686.700 718.650 690.600 ;
        RECT 723.750 686.700 725.550 690.600 ;
        RECT 733.050 686.700 734.850 690.600 ;
        RECT 746.700 686.700 748.500 693.600 ;
        RECT 772.800 686.700 774.600 691.800 ;
        RECT 790.500 686.700 792.300 693.600 ;
        RECT 808.800 686.700 810.600 690.600 ;
        RECT 816.150 686.700 817.950 690.600 ;
        RECT 825.450 686.700 827.250 690.600 ;
        RECT 832.350 686.700 834.150 690.600 ;
        RECT 841.350 686.700 843.150 690.600 ;
        RECT 858.450 686.700 867.450 756.300 ;
        RECT 0.600 684.300 867.450 686.700 ;
        RECT 16.800 679.200 18.600 684.300 ;
        RECT 32.700 680.400 34.500 684.300 ;
        RECT 40.200 677.400 42.000 684.300 ;
        RECT 52.800 680.400 54.600 684.300 ;
        RECT 58.800 680.400 60.600 684.300 ;
        RECT 76.500 677.400 78.300 684.300 ;
        RECT 97.500 674.400 99.300 684.300 ;
        RECT 107.700 674.400 109.500 684.300 ;
        RECT 128.400 680.400 130.200 684.300 ;
        RECT 143.700 674.400 145.500 684.300 ;
        RECT 164.700 674.400 166.500 684.300 ;
        RECT 185.700 674.400 187.500 684.300 ;
        RECT 206.700 677.400 208.500 684.300 ;
        RECT 224.400 680.400 226.200 684.300 ;
        RECT 247.500 677.400 249.300 684.300 ;
        RECT 257.400 677.400 259.200 684.300 ;
        RECT 275.700 680.400 277.500 684.300 ;
        RECT 283.200 677.400 285.000 684.300 ;
        RECT 304.500 674.400 306.300 684.300 ;
        RECT 314.700 677.400 316.500 684.300 ;
        RECT 340.800 679.200 342.600 684.300 ;
        RECT 361.500 677.400 363.300 684.300 ;
        RECT 378.300 677.400 380.100 684.300 ;
        RECT 397.800 677.400 399.600 684.300 ;
        RECT 406.200 677.400 408.000 684.300 ;
        RECT 416.700 677.400 418.500 684.300 ;
        RECT 437.400 680.400 439.200 684.300 ;
        RECT 443.400 680.400 445.200 684.300 ;
        RECT 458.700 677.400 460.500 684.300 ;
        RECT 473.700 677.400 475.500 684.300 ;
        RECT 491.400 677.400 493.200 684.300 ;
        RECT 509.400 679.200 511.200 684.300 ;
        RECT 527.400 683.400 528.600 684.300 ;
        RECT 527.400 680.400 529.200 683.400 ;
        RECT 533.400 680.400 535.200 684.300 ;
        RECT 551.400 679.200 553.200 684.300 ;
        RECT 577.500 677.400 579.300 684.300 ;
        RECT 592.500 677.400 594.300 684.300 ;
        RECT 608.700 677.400 610.500 684.300 ;
        RECT 631.500 677.400 633.300 684.300 ;
        RECT 649.800 679.200 651.600 684.300 ;
        RECT 662.400 677.400 664.200 684.300 ;
        RECT 668.400 677.400 670.200 684.300 ;
        RECT 674.400 677.400 676.200 684.300 ;
        RECT 680.400 677.400 682.200 684.300 ;
        RECT 686.400 677.400 688.200 684.300 ;
        RECT 695.850 680.400 697.650 684.300 ;
        RECT 704.850 680.400 706.650 684.300 ;
        RECT 711.750 680.400 713.550 684.300 ;
        RECT 721.050 680.400 722.850 684.300 ;
        RECT 742.800 679.200 744.600 684.300 ;
        RECT 755.700 677.400 757.500 684.300 ;
        RECT 776.700 677.400 778.500 684.300 ;
        RECT 788.850 680.400 790.650 684.300 ;
        RECT 797.850 680.400 799.650 684.300 ;
        RECT 804.750 680.400 806.550 684.300 ;
        RECT 814.050 680.400 815.850 684.300 ;
        RECT 830.400 679.200 832.200 684.300 ;
        RECT 11.700 614.700 13.500 618.600 ;
        RECT 19.200 614.700 21.000 621.600 ;
        RECT 40.500 614.700 42.300 624.600 ;
        RECT 58.500 614.700 60.300 621.600 ;
        RECT 79.500 614.700 81.300 624.600 ;
        RECT 97.800 614.700 99.600 619.800 ;
        RECT 115.800 614.700 117.600 621.600 ;
        RECT 124.200 614.700 126.000 621.600 ;
        RECT 134.700 614.700 136.500 621.600 ;
        RECT 156.900 614.700 158.700 621.600 ;
        RECT 184.500 614.700 186.300 624.600 ;
        RECT 199.800 614.700 201.600 618.600 ;
        RECT 214.800 614.700 216.600 618.600 ;
        RECT 232.800 614.700 234.600 619.800 ;
        RECT 256.500 614.700 258.300 624.600 ;
        RECT 266.700 614.700 268.500 621.600 ;
        RECT 292.800 614.700 294.600 619.800 ;
        RECT 305.700 614.700 307.500 621.600 ;
        RECT 331.800 614.700 333.600 619.800 ;
        RECT 347.400 614.700 349.200 619.800 ;
        RECT 372.300 614.700 374.100 621.600 ;
        RECT 387.000 614.700 388.800 621.600 ;
        RECT 395.400 614.700 397.200 621.600 ;
        RECT 411.000 614.700 412.800 621.600 ;
        RECT 419.400 614.700 421.200 621.600 ;
        RECT 434.400 614.700 436.200 618.600 ;
        RECT 457.500 614.700 459.300 621.600 ;
        RECT 474.300 614.700 476.100 621.600 ;
        RECT 496.800 614.700 498.600 619.800 ;
        RECT 512.400 614.700 514.200 619.800 ;
        RECT 535.800 614.700 537.600 618.600 ;
        RECT 553.500 614.700 555.300 621.600 ;
        RECT 563.700 614.700 565.500 621.600 ;
        RECT 589.500 614.700 591.300 621.600 ;
        RECT 599.400 614.700 601.200 618.600 ;
        RECT 617.700 614.700 619.500 621.600 ;
        RECT 632.700 614.700 634.500 621.600 ;
        RECT 658.800 614.700 660.600 619.800 ;
        RECT 668.850 614.700 670.650 618.600 ;
        RECT 677.850 614.700 679.650 618.600 ;
        RECT 684.750 614.700 686.550 618.600 ;
        RECT 694.050 614.700 695.850 618.600 ;
        RECT 712.500 614.700 714.300 621.600 ;
        RECT 723.150 614.700 724.950 618.600 ;
        RECT 732.450 614.700 734.250 618.600 ;
        RECT 739.350 614.700 741.150 618.600 ;
        RECT 748.350 614.700 750.150 618.600 ;
        RECT 764.700 614.700 766.500 621.600 ;
        RECT 782.400 614.700 784.200 619.800 ;
        RECT 800.700 614.700 802.500 621.600 ;
        RECT 826.500 614.700 828.300 621.600 ;
        RECT 839.400 614.700 841.200 619.800 ;
        RECT 858.450 614.700 867.450 684.300 ;
        RECT 0.600 612.300 867.450 614.700 ;
        RECT 19.500 602.400 21.300 612.300 ;
        RECT 30.000 605.400 31.800 612.300 ;
        RECT 37.500 608.400 39.300 612.300 ;
        RECT 50.700 602.400 52.500 612.300 ;
        RECT 74.400 607.200 76.200 612.300 ;
        RECT 92.700 605.400 94.500 612.300 ;
        RECT 110.400 608.400 112.200 612.300 ;
        RECT 116.400 608.400 118.200 612.300 ;
        RECT 128.700 605.400 130.500 612.300 ;
        RECT 154.500 605.400 156.300 612.300 ;
        RECT 175.500 602.400 177.300 612.300 ;
        RECT 186.000 605.400 187.800 612.300 ;
        RECT 193.500 608.400 195.300 612.300 ;
        RECT 209.700 608.400 211.500 612.300 ;
        RECT 217.200 605.400 219.000 612.300 ;
        RECT 230.400 607.200 232.200 612.300 ;
        RECT 248.400 608.400 250.200 612.300 ;
        RECT 263.700 605.400 265.500 612.300 ;
        RECT 288.300 605.400 290.100 612.300 ;
        RECT 302.400 605.400 304.200 612.300 ;
        RECT 322.800 605.400 324.600 612.300 ;
        RECT 331.200 605.400 333.000 612.300 ;
        RECT 346.500 605.400 348.300 612.300 ;
        RECT 362.700 605.400 364.500 612.300 ;
        RECT 382.500 605.400 384.300 612.300 ;
        RECT 403.500 605.400 405.300 612.300 ;
        RECT 418.800 608.400 420.600 612.300 ;
        RECT 425.400 611.400 426.600 612.300 ;
        RECT 424.800 608.400 426.600 611.400 ;
        RECT 439.800 608.400 441.600 612.300 ;
        RECT 446.400 611.400 447.600 612.300 ;
        RECT 445.800 608.400 447.600 611.400 ;
        RECT 458.700 608.400 460.500 612.300 ;
        RECT 466.200 605.400 468.000 612.300 ;
        RECT 487.500 602.400 489.300 612.300 ;
        RECT 502.800 608.400 504.600 612.300 ;
        RECT 523.500 602.400 525.300 612.300 ;
        RECT 534.000 605.400 535.800 612.300 ;
        RECT 541.500 608.400 543.300 612.300 ;
        RECT 557.400 607.200 559.200 612.300 ;
        RECT 575.400 608.400 577.200 612.300 ;
        RECT 581.400 608.400 583.200 612.300 ;
        RECT 596.400 607.200 598.200 612.300 ;
        RECT 614.400 605.400 616.200 612.300 ;
        RECT 620.400 605.400 622.200 612.300 ;
        RECT 626.400 605.400 628.200 612.300 ;
        RECT 632.400 605.400 634.200 612.300 ;
        RECT 638.400 605.400 640.200 612.300 ;
        RECT 658.500 605.400 660.300 612.300 ;
        RECT 676.800 607.200 678.600 612.300 ;
        RECT 689.700 605.400 691.500 612.300 ;
        RECT 715.800 607.200 717.600 612.300 ;
        RECT 731.400 607.200 733.200 612.300 ;
        RECT 749.700 605.400 751.500 612.300 ;
        RECT 770.400 607.200 772.200 612.300 ;
        RECT 788.700 605.400 790.500 612.300 ;
        RECT 811.800 608.400 813.600 612.300 ;
        RECT 821.400 605.400 823.200 612.300 ;
        RECT 827.400 605.400 829.200 612.300 ;
        RECT 842.700 605.400 844.500 612.300 ;
        RECT 13.500 542.700 15.300 549.600 ;
        RECT 34.800 542.700 36.600 547.800 ;
        RECT 55.800 542.700 57.600 547.800 ;
        RECT 71.100 542.700 73.200 546.600 ;
        RECT 77.400 542.700 79.200 546.600 ;
        RECT 104.700 542.700 106.500 546.600 ;
        RECT 112.200 542.700 114.000 549.600 ;
        RECT 133.500 542.700 135.300 552.600 ;
        RECT 148.800 542.700 150.600 549.600 ;
        RECT 157.200 542.700 159.000 549.600 ;
        RECT 174.300 542.700 176.100 549.600 ;
        RECT 199.500 542.700 201.300 552.600 ;
        RECT 214.800 542.700 216.600 546.600 ;
        RECT 232.800 542.700 234.600 547.800 ;
        RECT 253.800 542.700 255.600 547.800 ;
        RECT 271.800 542.700 273.600 546.600 ;
        RECT 277.800 543.600 279.600 546.600 ;
        RECT 278.400 542.700 279.600 543.600 ;
        RECT 287.400 542.700 289.200 546.600 ;
        RECT 293.400 542.700 295.200 546.600 ;
        RECT 305.700 542.700 307.500 549.600 ;
        RECT 327.900 542.700 329.700 549.600 ;
        RECT 346.800 542.700 348.600 546.600 ;
        RECT 352.800 542.700 354.600 546.600 ;
        RECT 362.700 542.700 364.500 549.600 ;
        RECT 380.400 542.700 382.200 546.600 ;
        RECT 403.500 542.700 405.300 549.600 ;
        RECT 416.700 542.700 418.500 546.600 ;
        RECT 424.200 542.700 426.000 549.600 ;
        RECT 442.500 542.700 444.300 549.600 ;
        RECT 453.000 542.700 454.800 549.600 ;
        RECT 461.400 542.700 463.200 549.600 ;
        RECT 476.400 542.700 478.200 546.600 ;
        RECT 482.400 542.700 484.200 546.600 ;
        RECT 497.400 542.700 499.200 547.800 ;
        RECT 517.800 542.700 519.600 546.600 ;
        RECT 523.800 542.700 525.600 546.600 ;
        RECT 533.700 542.700 535.500 552.600 ;
        RECT 554.700 542.700 556.500 552.600 ;
        RECT 575.700 542.700 577.500 552.600 ;
        RECT 600.900 542.700 602.700 549.600 ;
        RECT 620.400 542.700 622.200 547.800 ;
        RECT 635.850 542.700 637.650 546.600 ;
        RECT 644.850 542.700 646.650 546.600 ;
        RECT 651.750 542.700 653.550 546.600 ;
        RECT 661.050 542.700 662.850 546.600 ;
        RECT 671.850 542.700 673.650 546.600 ;
        RECT 680.850 542.700 682.650 546.600 ;
        RECT 687.750 542.700 689.550 546.600 ;
        RECT 697.050 542.700 698.850 546.600 ;
        RECT 707.850 542.700 709.650 546.600 ;
        RECT 716.850 542.700 718.650 546.600 ;
        RECT 723.750 542.700 725.550 546.600 ;
        RECT 733.050 542.700 734.850 546.600 ;
        RECT 749.400 542.700 751.200 547.800 ;
        RECT 767.700 542.700 769.500 549.600 ;
        RECT 785.400 542.700 787.200 546.600 ;
        RECT 797.850 542.700 799.650 546.600 ;
        RECT 806.850 542.700 808.650 546.600 ;
        RECT 813.750 542.700 815.550 546.600 ;
        RECT 823.050 542.700 824.850 546.600 ;
        RECT 836.400 542.700 838.200 546.600 ;
        RECT 858.450 542.700 867.450 612.300 ;
        RECT 0.600 540.300 867.450 542.700 ;
        RECT 11.700 536.400 13.500 540.300 ;
        RECT 19.200 533.400 21.000 540.300 ;
        RECT 29.700 530.400 31.500 540.300 ;
        RECT 50.700 530.400 52.500 540.300 ;
        RECT 72.000 533.400 73.800 540.300 ;
        RECT 79.500 536.400 81.300 540.300 ;
        RECT 95.400 535.200 97.200 540.300 ;
        RECT 113.700 530.400 115.500 540.300 ;
        RECT 135.000 533.400 136.800 540.300 ;
        RECT 142.500 536.400 144.300 540.300 ;
        RECT 160.800 536.400 162.600 540.300 ;
        RECT 171.000 533.400 172.800 540.300 ;
        RECT 179.400 533.400 181.200 540.300 ;
        RECT 194.700 530.400 196.500 540.300 ;
        RECT 223.500 533.400 225.300 540.300 ;
        RECT 240.300 533.400 242.100 540.300 ;
        RECT 255.000 533.400 256.800 540.300 ;
        RECT 263.400 533.400 265.200 540.300 ;
        RECT 286.500 533.400 288.300 540.300 ;
        RECT 296.400 536.400 298.200 540.300 ;
        RECT 302.400 536.400 304.200 540.300 ;
        RECT 322.800 535.200 324.600 540.300 ;
        RECT 335.400 536.400 337.200 540.300 ;
        RECT 350.700 533.400 352.500 540.300 ;
        RECT 369.000 533.400 370.800 540.300 ;
        RECT 376.500 536.400 378.300 540.300 ;
        RECT 389.400 536.400 391.200 540.300 ;
        RECT 404.400 536.400 406.200 540.300 ;
        RECT 410.400 536.400 412.200 540.300 ;
        RECT 425.400 535.200 427.200 540.300 ;
        RECT 443.400 536.400 445.200 540.300 ;
        RECT 458.700 530.400 460.500 540.300 ;
        RECT 480.000 533.400 481.800 540.300 ;
        RECT 487.500 536.400 489.300 540.300 ;
        RECT 500.400 536.400 502.200 540.300 ;
        RECT 516.000 533.400 517.800 540.300 ;
        RECT 523.500 536.400 525.300 540.300 ;
        RECT 536.700 530.400 538.500 540.300 ;
        RECT 560.400 535.200 562.200 540.300 ;
        RECT 580.800 533.400 582.600 540.300 ;
        RECT 586.800 533.400 588.600 540.300 ;
        RECT 592.800 533.400 594.600 540.300 ;
        RECT 598.800 533.400 600.600 540.300 ;
        RECT 604.800 533.400 606.600 540.300 ;
        RECT 616.800 533.400 618.600 540.300 ;
        RECT 622.800 533.400 624.600 540.300 ;
        RECT 628.800 533.400 630.600 540.300 ;
        RECT 634.800 533.400 636.600 540.300 ;
        RECT 640.800 533.400 642.600 540.300 ;
        RECT 653.400 535.200 655.200 540.300 ;
        RECT 671.700 533.400 673.500 540.300 ;
        RECT 692.400 535.200 694.200 540.300 ;
        RECT 710.700 533.400 712.500 540.300 ;
        RECT 725.850 536.400 727.650 540.300 ;
        RECT 734.850 536.400 736.650 540.300 ;
        RECT 741.750 536.400 743.550 540.300 ;
        RECT 751.050 536.400 752.850 540.300 ;
        RECT 765.000 533.400 766.800 540.300 ;
        RECT 772.500 536.400 774.300 540.300 ;
        RECT 788.400 535.200 790.200 540.300 ;
        RECT 806.400 536.400 808.200 540.300 ;
        RECT 824.400 535.200 826.200 540.300 ;
        RECT 842.700 533.400 844.500 540.300 ;
        RECT 16.800 470.700 18.600 475.800 ;
        RECT 32.400 470.700 34.200 475.800 ;
        RECT 50.700 470.700 52.500 480.600 ;
        RECT 82.500 470.700 84.300 480.600 ;
        RECT 93.000 470.700 94.800 477.600 ;
        RECT 100.500 470.700 102.300 474.600 ;
        RECT 118.800 470.700 120.600 474.600 ;
        RECT 129.000 470.700 130.800 477.600 ;
        RECT 136.500 470.700 138.300 474.600 ;
        RECT 152.400 470.700 154.200 475.800 ;
        RECT 170.700 470.700 172.500 480.600 ;
        RECT 199.800 470.700 201.600 475.800 ;
        RECT 217.800 470.700 219.600 474.600 ;
        RECT 232.500 470.700 234.300 477.600 ;
        RECT 256.500 470.700 258.300 480.600 ;
        RECT 271.800 470.700 273.600 474.600 ;
        RECT 285.900 470.700 287.700 477.600 ;
        RECT 302.700 470.700 304.500 477.600 ;
        RECT 328.500 470.700 330.300 477.600 ;
        RECT 346.500 470.700 348.300 477.600 ;
        RECT 356.700 470.700 358.500 480.600 ;
        RECT 378.000 470.700 379.800 477.600 ;
        RECT 385.500 470.700 387.300 474.600 ;
        RECT 406.800 470.700 408.600 475.800 ;
        RECT 421.800 470.700 423.600 474.600 ;
        RECT 427.800 470.700 429.600 474.600 ;
        RECT 442.800 470.700 444.600 474.600 ;
        RECT 453.000 470.700 454.800 477.600 ;
        RECT 460.500 470.700 462.300 474.600 ;
        RECT 476.100 470.700 478.200 474.600 ;
        RECT 482.400 470.700 484.200 474.600 ;
        RECT 511.800 470.700 513.600 474.600 ;
        RECT 524.400 470.700 526.200 475.800 ;
        RECT 539.850 470.700 541.650 474.600 ;
        RECT 548.850 470.700 550.650 474.600 ;
        RECT 555.750 470.700 557.550 474.600 ;
        RECT 565.050 470.700 566.850 474.600 ;
        RECT 575.850 470.700 577.650 474.600 ;
        RECT 584.850 470.700 586.650 474.600 ;
        RECT 591.750 470.700 593.550 474.600 ;
        RECT 601.050 470.700 602.850 474.600 ;
        RECT 622.500 470.700 624.300 477.600 ;
        RECT 640.800 470.700 642.600 475.800 ;
        RECT 653.400 470.700 655.200 474.600 ;
        RECT 673.800 470.700 675.600 474.600 ;
        RECT 691.500 470.700 693.300 477.600 ;
        RECT 709.500 470.700 711.300 477.600 ;
        RECT 720.000 470.700 721.800 477.600 ;
        RECT 728.400 470.700 730.200 477.600 ;
        RECT 751.800 470.700 753.600 475.800 ;
        RECT 769.800 470.700 771.600 474.600 ;
        RECT 781.800 470.700 783.600 474.600 ;
        RECT 787.800 470.700 789.600 474.600 ;
        RECT 800.400 470.700 802.200 475.800 ;
        RECT 826.800 470.700 828.600 475.800 ;
        RECT 841.800 470.700 843.600 474.600 ;
        RECT 847.800 470.700 849.600 474.600 ;
        RECT 858.450 470.700 867.450 540.300 ;
        RECT 0.600 468.300 867.450 470.700 ;
        RECT 15.300 461.400 17.100 468.300 ;
        RECT 29.700 461.400 31.500 468.300 ;
        RECT 58.500 458.400 60.300 468.300 ;
        RECT 71.700 464.400 73.500 468.300 ;
        RECT 79.200 461.400 81.000 468.300 ;
        RECT 100.500 458.400 102.300 468.300 ;
        RECT 110.400 464.400 112.200 468.300 ;
        RECT 133.800 463.200 135.600 468.300 ;
        RECT 148.800 464.400 150.600 468.300 ;
        RECT 154.800 464.400 156.600 468.300 ;
        RECT 164.700 461.400 166.500 468.300 ;
        RECT 193.500 458.400 195.300 468.300 ;
        RECT 203.700 461.400 205.500 468.300 ;
        RECT 222.000 461.400 223.800 468.300 ;
        RECT 230.400 461.400 232.200 468.300 ;
        RECT 250.500 461.400 252.300 468.300 ;
        RECT 274.500 458.400 276.300 468.300 ;
        RECT 287.400 463.200 289.200 468.300 ;
        RECT 313.800 463.200 315.600 468.300 ;
        RECT 330.900 461.400 332.700 468.300 ;
        RECT 351.900 461.400 353.700 468.300 ;
        RECT 376.500 461.400 378.300 468.300 ;
        RECT 394.800 463.200 396.600 468.300 ;
        RECT 410.400 463.200 412.200 468.300 ;
        RECT 431.400 463.200 433.200 468.300 ;
        RECT 454.800 464.400 456.600 468.300 ;
        RECT 467.400 463.200 469.200 468.300 ;
        RECT 488.400 463.200 490.200 468.300 ;
        RECT 509.400 463.200 511.200 468.300 ;
        RECT 532.500 461.400 534.300 468.300 ;
        RECT 547.800 461.400 549.600 468.300 ;
        RECT 553.800 461.400 555.600 468.300 ;
        RECT 566.700 461.400 568.500 468.300 ;
        RECT 581.400 464.400 583.200 468.300 ;
        RECT 598.800 464.400 600.600 468.300 ;
        RECT 604.800 464.400 606.600 468.300 ;
        RECT 614.400 464.400 616.200 468.300 ;
        RECT 631.800 464.400 633.600 468.300 ;
        RECT 637.800 464.400 639.600 468.300 ;
        RECT 650.400 463.200 652.200 468.300 ;
        RECT 676.500 461.400 678.300 468.300 ;
        RECT 687.000 461.400 688.800 468.300 ;
        RECT 695.400 461.400 697.200 468.300 ;
        RECT 713.400 463.200 715.200 468.300 ;
        RECT 731.700 461.400 733.500 468.300 ;
        RECT 749.700 458.400 751.500 468.300 ;
        RECT 770.700 458.400 772.500 468.300 ;
        RECT 799.800 463.200 801.600 468.300 ;
        RECT 820.800 463.200 822.600 468.300 ;
        RECT 833.400 467.400 834.600 468.300 ;
        RECT 833.400 464.400 835.200 467.400 ;
        RECT 839.400 464.400 841.200 468.300 ;
        RECT 16.800 398.700 18.600 403.800 ;
        RECT 40.500 398.700 42.300 408.600 ;
        RECT 53.700 398.700 55.500 402.600 ;
        RECT 61.200 398.700 63.000 405.600 ;
        RECT 79.800 398.700 81.600 403.800 ;
        RECT 97.800 398.700 99.600 402.600 ;
        RECT 115.800 398.700 117.600 403.800 ;
        RECT 131.400 398.700 133.200 403.800 ;
        RECT 157.500 398.700 159.300 405.600 ;
        RECT 167.700 398.700 169.500 405.600 ;
        RECT 185.700 398.700 187.500 405.600 ;
        RECT 210.300 398.700 212.100 405.600 ;
        RECT 225.000 398.700 226.800 405.600 ;
        RECT 233.400 398.700 235.200 405.600 ;
        RECT 251.700 398.700 253.500 405.600 ;
        RECT 269.700 398.700 271.500 405.600 ;
        RECT 292.500 398.700 294.300 405.600 ;
        RECT 310.800 398.700 312.600 403.800 ;
        RECT 323.700 398.700 325.500 405.600 ;
        RECT 348.300 398.700 350.100 405.600 ;
        RECT 362.700 398.700 364.500 405.600 ;
        RECT 381.000 398.700 382.800 405.600 ;
        RECT 388.500 398.700 390.300 402.600 ;
        RECT 406.500 398.700 408.300 405.600 ;
        RECT 422.400 398.700 424.200 403.800 ;
        RECT 443.400 398.700 445.200 403.800 ;
        RECT 466.800 398.700 468.600 402.600 ;
        RECT 473.850 398.700 475.650 402.600 ;
        RECT 482.850 398.700 484.650 402.600 ;
        RECT 489.750 398.700 491.550 402.600 ;
        RECT 499.050 398.700 500.850 402.600 ;
        RECT 515.400 398.700 517.200 403.800 ;
        RECT 533.700 398.700 535.500 405.600 ;
        RECT 553.800 398.700 555.600 402.600 ;
        RECT 559.800 398.700 561.600 402.600 ;
        RECT 574.500 398.700 576.300 405.600 ;
        RECT 595.500 398.700 597.300 405.600 ;
        RECT 608.400 398.700 610.200 403.800 ;
        RECT 631.800 398.700 633.600 405.600 ;
        RECT 640.200 398.700 642.000 405.600 ;
        RECT 653.400 398.700 655.200 403.800 ;
        RECT 679.500 398.700 681.300 405.600 ;
        RECT 692.400 398.700 694.200 403.800 ;
        RECT 718.800 398.700 720.600 403.800 ;
        RECT 734.400 398.700 736.200 403.800 ;
        RECT 743.400 398.700 745.200 406.800 ;
        RECT 755.700 398.700 757.500 405.600 ;
        RECT 778.800 398.700 780.600 405.600 ;
        RECT 793.800 398.700 795.600 405.600 ;
        RECT 811.500 398.700 813.300 405.600 ;
        RECT 821.700 398.700 823.500 405.600 ;
        RECT 843.900 398.700 845.700 405.600 ;
        RECT 858.450 398.700 867.450 468.300 ;
        RECT 0.600 396.300 867.450 398.700 ;
        RECT 19.500 386.400 21.300 396.300 ;
        RECT 30.000 389.400 31.800 396.300 ;
        RECT 37.500 392.400 39.300 396.300 ;
        RECT 61.500 386.400 63.300 396.300 ;
        RECT 76.800 389.400 78.600 396.300 ;
        RECT 85.200 389.400 87.000 396.300 ;
        RECT 98.700 392.400 100.500 396.300 ;
        RECT 106.200 389.400 108.000 396.300 ;
        RECT 121.800 392.400 123.600 396.300 ;
        RECT 139.500 389.400 141.300 396.300 ;
        RECT 160.500 386.400 162.300 396.300 ;
        RECT 170.400 392.400 172.200 396.300 ;
        RECT 176.400 392.400 178.200 396.300 ;
        RECT 196.500 389.400 198.300 396.300 ;
        RECT 211.800 392.400 213.600 396.300 ;
        RECT 226.800 392.400 228.600 396.300 ;
        RECT 247.500 386.400 249.300 396.300 ;
        RECT 262.800 389.400 264.600 396.300 ;
        RECT 271.200 389.400 273.000 396.300 ;
        RECT 286.800 392.400 288.600 396.300 ;
        RECT 307.500 386.400 309.300 396.300 ;
        RECT 320.400 391.200 322.200 396.300 ;
        RECT 345.300 389.400 347.100 396.300 ;
        RECT 364.500 389.400 366.300 396.300 ;
        RECT 381.900 389.400 383.700 396.300 ;
        RECT 403.500 389.400 405.300 396.300 ;
        RECT 416.400 392.400 418.200 396.300 ;
        RECT 432.000 389.400 433.800 396.300 ;
        RECT 440.400 389.400 442.200 396.300 ;
        RECT 452.850 392.400 454.650 396.300 ;
        RECT 461.850 392.400 463.650 396.300 ;
        RECT 468.750 392.400 470.550 396.300 ;
        RECT 478.050 392.400 479.850 396.300 ;
        RECT 494.400 391.200 496.200 396.300 ;
        RECT 513.000 389.400 514.800 396.300 ;
        RECT 520.500 392.400 522.300 396.300 ;
        RECT 541.800 391.200 543.600 396.300 ;
        RECT 562.800 391.200 564.600 396.300 ;
        RECT 577.800 388.200 579.600 396.300 ;
        RECT 586.800 391.200 588.600 396.300 ;
        RECT 599.700 389.400 601.500 396.300 ;
        RECT 620.400 391.200 622.200 396.300 ;
        RECT 639.000 389.400 640.800 396.300 ;
        RECT 647.400 389.400 649.200 396.300 ;
        RECT 673.500 386.400 675.300 396.300 ;
        RECT 686.700 389.400 688.500 396.300 ;
        RECT 709.500 389.400 711.300 396.300 ;
        RECT 719.400 392.400 721.200 396.300 ;
        RECT 739.800 392.400 741.600 396.300 ;
        RECT 755.700 389.400 757.500 396.300 ;
        RECT 770.700 389.400 772.500 396.300 ;
        RECT 796.800 391.200 798.600 396.300 ;
        RECT 810.000 389.400 811.800 396.300 ;
        RECT 818.400 389.400 820.200 396.300 ;
        RECT 833.700 389.400 835.500 396.300 ;
        RECT 19.500 326.700 21.300 336.600 ;
        RECT 37.800 326.700 39.600 331.800 ;
        RECT 53.400 326.700 55.200 331.800 ;
        RECT 82.500 326.700 84.300 336.600 ;
        RECT 100.800 326.700 102.600 331.800 ;
        RECT 113.700 326.700 115.500 336.600 ;
        RECT 137.400 326.700 139.200 331.800 ;
        RECT 166.500 326.700 168.300 336.600 ;
        RECT 187.500 326.700 189.300 336.600 ;
        RECT 197.700 326.700 199.500 333.600 ;
        RECT 223.800 326.700 225.600 331.800 ;
        RECT 236.400 326.700 238.200 330.600 ;
        RECT 242.400 326.700 244.200 330.600 ;
        RECT 262.800 326.700 264.600 331.800 ;
        RECT 283.800 326.700 285.600 331.800 ;
        RECT 299.400 326.700 301.200 331.800 ;
        RECT 325.500 326.700 327.300 333.600 ;
        RECT 342.300 326.700 344.100 333.600 ;
        RECT 364.500 326.700 366.300 333.600 ;
        RECT 374.400 326.700 376.200 333.600 ;
        RECT 389.700 326.700 391.500 333.600 ;
        RECT 410.700 326.700 412.500 333.600 ;
        RECT 430.800 326.700 432.600 330.600 ;
        RECT 442.800 326.700 444.600 330.600 ;
        RECT 448.800 326.700 450.600 330.600 ;
        RECT 463.800 326.700 465.600 333.600 ;
        RECT 472.200 326.700 474.000 333.600 ;
        RECT 484.800 326.700 486.600 330.600 ;
        RECT 490.800 326.700 492.600 330.600 ;
        RECT 502.800 326.700 504.600 330.600 ;
        RECT 508.800 326.700 510.600 330.600 ;
        RECT 521.700 326.700 523.500 330.600 ;
        RECT 529.200 326.700 531.000 333.600 ;
        RECT 544.800 326.700 546.600 330.600 ;
        RECT 557.400 326.700 559.200 331.800 ;
        RECT 583.500 326.700 585.300 333.600 ;
        RECT 596.400 326.700 598.200 331.800 ;
        RECT 622.800 326.700 624.600 331.800 ;
        RECT 635.400 326.700 637.200 330.600 ;
        RECT 641.400 326.700 643.200 330.600 ;
        RECT 661.500 326.700 663.300 333.600 ;
        RECT 676.800 326.700 678.600 333.600 ;
        RECT 685.200 326.700 687.000 333.600 ;
        RECT 696.000 326.700 697.800 333.600 ;
        RECT 704.400 326.700 706.200 333.600 ;
        RECT 727.500 326.700 729.300 333.600 ;
        RECT 744.300 326.700 746.100 333.600 ;
        RECT 759.000 326.700 760.800 333.600 ;
        RECT 767.400 326.700 769.200 333.600 ;
        RECT 783.000 326.700 784.800 333.600 ;
        RECT 791.400 326.700 793.200 333.600 ;
        RECT 814.800 326.700 816.600 331.800 ;
        RECT 830.400 326.700 832.200 331.800 ;
        RECT 858.450 326.700 867.450 396.300 ;
        RECT 0.600 324.300 867.450 326.700 ;
        RECT 11.700 320.400 13.500 324.300 ;
        RECT 19.200 317.400 21.000 324.300 ;
        RECT 29.700 314.400 31.500 324.300 ;
        RECT 53.700 320.400 55.500 324.300 ;
        RECT 61.200 317.400 63.000 324.300 ;
        RECT 79.800 319.200 81.600 324.300 ;
        RECT 99.300 317.400 101.100 324.300 ;
        RECT 113.700 317.400 115.500 324.300 ;
        RECT 131.700 317.400 133.500 324.300 ;
        RECT 157.500 317.400 159.300 324.300 ;
        RECT 178.500 314.400 180.300 324.300 ;
        RECT 199.500 314.400 201.300 324.300 ;
        RECT 214.800 320.400 216.600 324.300 ;
        RECT 229.800 317.400 231.600 324.300 ;
        RECT 238.200 317.400 240.000 324.300 ;
        RECT 256.500 317.400 258.300 324.300 ;
        RECT 271.800 317.400 273.600 324.300 ;
        RECT 280.200 317.400 282.000 324.300 ;
        RECT 301.500 314.400 303.300 324.300 ;
        RECT 314.400 319.200 316.200 324.300 ;
        RECT 340.500 317.400 342.300 324.300 ;
        RECT 361.500 314.400 363.300 324.300 ;
        RECT 374.400 319.200 376.200 324.300 ;
        RECT 396.900 317.400 398.700 324.300 ;
        RECT 413.400 320.400 415.200 324.300 ;
        RECT 428.700 317.400 430.500 324.300 ;
        RECT 446.700 317.400 448.500 324.300 ;
        RECT 467.400 319.200 469.200 324.300 ;
        RECT 485.700 317.400 487.500 324.300 ;
        RECT 504.000 317.400 505.800 324.300 ;
        RECT 511.500 320.400 513.300 324.300 ;
        RECT 527.400 319.200 529.200 324.300 ;
        RECT 545.400 320.400 547.200 324.300 ;
        RECT 551.400 320.400 553.200 324.300 ;
        RECT 574.500 314.400 576.300 324.300 ;
        RECT 584.700 317.400 586.500 324.300 ;
        RECT 613.500 314.400 615.300 324.300 ;
        RECT 631.800 319.200 633.600 324.300 ;
        RECT 652.800 319.200 654.600 324.300 ;
        RECT 672.300 317.400 674.100 324.300 ;
        RECT 689.400 319.200 691.200 324.300 ;
        RECT 707.700 317.400 709.500 324.300 ;
        RECT 733.500 317.400 735.300 324.300 ;
        RECT 751.800 319.200 753.600 324.300 ;
        RECT 767.400 319.200 769.200 324.300 ;
        RECT 788.400 319.200 790.200 324.300 ;
        RECT 813.300 317.400 815.100 324.300 ;
        RECT 831.900 317.400 833.700 324.300 ;
        RECT 11.700 254.700 13.500 258.600 ;
        RECT 19.200 254.700 21.000 261.600 ;
        RECT 29.700 254.700 31.500 264.600 ;
        RECT 53.400 254.700 55.200 259.800 ;
        RECT 74.400 254.700 76.200 259.800 ;
        RECT 92.700 254.700 94.500 264.600 ;
        RECT 113.700 254.700 115.500 264.600 ;
        RECT 134.700 254.700 136.500 264.600 ;
        RECT 156.000 254.700 157.800 261.600 ;
        RECT 163.500 254.700 165.300 258.600 ;
        RECT 179.400 254.700 181.200 259.800 ;
        RECT 200.700 254.700 202.500 258.600 ;
        RECT 208.200 254.700 210.000 261.600 ;
        RECT 223.800 254.700 225.600 258.600 ;
        RECT 240.300 254.700 242.100 261.600 ;
        RECT 254.700 254.700 256.500 261.600 ;
        RECT 277.800 254.700 279.600 258.600 ;
        RECT 283.800 255.600 285.600 258.600 ;
        RECT 284.400 254.700 285.600 255.600 ;
        RECT 293.700 254.700 295.500 261.600 ;
        RECT 319.800 254.700 321.600 259.800 ;
        RECT 334.800 254.700 336.600 258.600 ;
        RECT 340.800 254.700 342.600 258.600 ;
        RECT 353.400 254.700 355.200 259.800 ;
        RECT 371.400 254.700 373.200 258.600 ;
        RECT 377.400 254.700 379.200 258.600 ;
        RECT 389.700 254.700 391.500 261.600 ;
        RECT 412.800 254.700 414.600 258.600 ;
        RECT 430.500 254.700 432.300 261.600 ;
        RECT 443.700 254.700 445.500 258.600 ;
        RECT 451.200 254.700 453.000 261.600 ;
        RECT 466.800 254.700 468.600 261.600 ;
        RECT 475.200 254.700 477.000 261.600 ;
        RECT 485.700 254.700 487.500 261.600 ;
        RECT 503.400 254.700 505.200 258.600 ;
        RECT 509.400 254.700 511.200 258.600 ;
        RECT 521.400 254.700 523.200 258.600 ;
        RECT 527.400 254.700 529.200 258.600 ;
        RECT 547.800 254.700 549.600 259.800 ;
        RECT 565.800 254.700 567.600 261.600 ;
        RECT 574.200 254.700 576.000 261.600 ;
        RECT 585.000 254.700 586.800 261.600 ;
        RECT 592.500 254.700 594.300 258.600 ;
        RECT 613.800 254.700 615.600 259.800 ;
        RECT 634.800 254.700 636.600 259.800 ;
        RECT 647.400 254.700 649.200 258.600 ;
        RECT 662.400 254.700 664.200 258.600 ;
        RECT 685.800 254.700 687.600 259.800 ;
        RECT 699.000 254.700 700.800 261.600 ;
        RECT 706.500 254.700 708.300 258.600 ;
        RECT 722.700 254.700 724.500 261.600 ;
        RECT 740.400 254.700 742.200 259.800 ;
        RECT 759.000 254.700 760.800 261.600 ;
        RECT 766.500 254.700 768.300 258.600 ;
        RECT 782.700 254.700 784.500 261.600 ;
        RECT 799.800 254.700 801.600 258.600 ;
        RECT 805.800 254.700 807.600 258.600 ;
        RECT 820.500 254.700 822.300 261.600 ;
        RECT 841.800 254.700 843.600 259.800 ;
        RECT 858.450 254.700 867.450 324.300 ;
        RECT 0.600 252.300 867.450 254.700 ;
        RECT 16.800 247.200 18.600 252.300 ;
        RECT 32.700 248.400 34.500 252.300 ;
        RECT 40.200 245.400 42.000 252.300 ;
        RECT 53.700 248.400 55.500 252.300 ;
        RECT 61.200 245.400 63.000 252.300 ;
        RECT 71.700 242.400 73.500 252.300 ;
        RECT 103.500 242.400 105.300 252.300 ;
        RECT 116.700 248.400 118.500 252.300 ;
        RECT 124.200 245.400 126.000 252.300 ;
        RECT 137.400 247.200 139.200 252.300 ;
        RECT 156.000 245.400 157.800 252.300 ;
        RECT 163.500 248.400 165.300 252.300 ;
        RECT 176.700 242.400 178.500 252.300 ;
        RECT 200.400 247.200 202.200 252.300 ;
        RECT 221.400 247.200 223.200 252.300 ;
        RECT 239.700 242.400 241.500 252.300 ;
        RECT 261.000 245.400 262.800 252.300 ;
        RECT 268.500 248.400 270.300 252.300 ;
        RECT 281.700 242.400 283.500 252.300 ;
        RECT 303.000 245.400 304.800 252.300 ;
        RECT 310.500 248.400 312.300 252.300 ;
        RECT 323.700 242.400 325.500 252.300 ;
        RECT 347.700 248.400 349.500 252.300 ;
        RECT 355.200 245.400 357.000 252.300 ;
        RECT 365.700 242.400 367.500 252.300 ;
        RECT 391.800 248.400 393.600 252.300 ;
        RECT 409.800 247.200 411.600 252.300 ;
        RECT 425.400 247.200 427.200 252.300 ;
        RECT 443.700 245.400 445.500 252.300 ;
        RECT 469.500 245.400 471.300 252.300 ;
        RECT 483.900 245.400 485.700 252.300 ;
        RECT 503.400 247.200 505.200 252.300 ;
        RECT 524.400 247.200 526.200 252.300 ;
        RECT 542.700 245.400 544.500 252.300 ;
        RECT 565.800 248.400 567.600 252.300 ;
        RECT 580.800 248.400 582.600 252.300 ;
        RECT 587.850 248.400 589.650 252.300 ;
        RECT 596.850 248.400 598.650 252.300 ;
        RECT 603.750 248.400 605.550 252.300 ;
        RECT 613.050 248.400 614.850 252.300 ;
        RECT 626.400 248.400 628.200 252.300 ;
        RECT 641.700 245.400 643.500 252.300 ;
        RECT 667.500 245.400 669.300 252.300 ;
        RECT 680.400 247.200 682.200 252.300 ;
        RECT 689.400 244.200 691.200 252.300 ;
        RECT 709.800 247.200 711.600 252.300 ;
        RECT 725.400 247.200 727.200 252.300 ;
        RECT 746.400 247.200 748.200 252.300 ;
        RECT 767.400 247.200 769.200 252.300 ;
        RECT 786.000 245.400 787.800 252.300 ;
        RECT 793.500 248.400 795.300 252.300 ;
        RECT 809.700 248.400 811.500 252.300 ;
        RECT 817.200 245.400 819.000 252.300 ;
        RECT 830.400 247.200 832.200 252.300 ;
        RECT 16.800 182.700 18.600 187.800 ;
        RECT 29.700 182.700 31.500 192.600 ;
        RECT 50.700 182.700 52.500 192.600 ;
        RECT 74.700 182.700 76.500 186.600 ;
        RECT 82.200 182.700 84.000 189.600 ;
        RECT 100.800 182.700 102.600 187.800 ;
        RECT 121.800 182.700 123.600 187.800 ;
        RECT 134.700 182.700 136.500 192.600 ;
        RECT 162.300 182.700 164.100 189.600 ;
        RECT 176.700 182.700 178.500 189.600 ;
        RECT 202.500 182.700 204.300 189.600 ;
        RECT 212.700 182.700 214.500 189.600 ;
        RECT 238.500 182.700 240.300 189.600 ;
        RECT 251.100 182.700 253.200 186.600 ;
        RECT 257.400 182.700 259.200 186.600 ;
        RECT 281.400 182.700 283.200 186.600 ;
        RECT 299.400 182.700 301.200 187.800 ;
        RECT 322.800 182.700 324.600 186.600 ;
        RECT 333.000 182.700 334.800 189.600 ;
        RECT 340.500 182.700 342.300 186.600 ;
        RECT 361.500 182.700 363.300 189.600 ;
        RECT 379.500 182.700 381.300 189.600 ;
        RECT 391.800 182.700 393.600 186.600 ;
        RECT 397.800 182.700 399.600 186.600 ;
        RECT 410.400 182.700 412.200 188.100 ;
        RECT 436.800 182.700 438.600 189.600 ;
        RECT 446.400 182.700 448.200 186.600 ;
        RECT 452.400 182.700 454.200 186.600 ;
        RECT 469.800 182.700 471.600 189.600 ;
        RECT 478.200 182.700 480.000 189.600 ;
        RECT 493.800 182.700 495.600 186.600 ;
        RECT 500.850 182.700 502.650 186.600 ;
        RECT 509.850 182.700 511.650 186.600 ;
        RECT 516.750 182.700 518.550 186.600 ;
        RECT 526.050 182.700 527.850 186.600 ;
        RECT 544.800 182.700 546.600 186.600 ;
        RECT 557.700 182.700 559.500 186.600 ;
        RECT 565.200 182.700 567.000 189.600 ;
        RECT 583.800 182.700 585.600 187.800 ;
        RECT 598.800 182.700 600.600 186.600 ;
        RECT 604.800 182.700 606.600 186.600 ;
        RECT 621.300 182.700 623.100 189.600 ;
        RECT 646.500 182.700 648.300 192.600 ;
        RECT 656.700 182.700 658.500 189.600 ;
        RECT 674.400 182.700 676.200 186.600 ;
        RECT 680.400 182.700 682.200 186.600 ;
        RECT 695.400 182.700 697.200 187.800 ;
        RECT 716.400 182.700 718.200 187.800 ;
        RECT 734.400 182.700 736.200 186.600 ;
        RECT 752.400 182.700 754.200 188.100 ;
        RECT 775.800 182.700 777.600 186.600 ;
        RECT 781.800 182.700 783.600 186.600 ;
        RECT 799.500 182.700 801.300 189.600 ;
        RECT 812.700 182.700 814.500 186.600 ;
        RECT 820.200 182.700 822.000 189.600 ;
        RECT 830.700 182.700 832.500 189.600 ;
        RECT 853.800 182.700 855.600 186.600 ;
        RECT 858.450 182.700 867.450 252.300 ;
        RECT 0.600 180.300 867.450 182.700 ;
        RECT 16.800 175.200 18.600 180.300 ;
        RECT 40.500 170.400 42.300 180.300 ;
        RECT 51.000 173.400 52.800 180.300 ;
        RECT 58.500 176.400 60.300 180.300 ;
        RECT 72.000 173.400 73.800 180.300 ;
        RECT 79.500 176.400 81.300 180.300 ;
        RECT 92.700 170.400 94.500 180.300 ;
        RECT 116.400 175.200 118.200 180.300 ;
        RECT 134.700 170.400 136.500 180.300 ;
        RECT 160.800 173.400 162.600 180.300 ;
        RECT 169.200 173.400 171.000 180.300 ;
        RECT 179.700 170.400 181.500 180.300 ;
        RECT 201.000 173.400 202.800 180.300 ;
        RECT 208.500 176.400 210.300 180.300 ;
        RECT 221.700 173.400 223.500 180.300 ;
        RECT 239.700 170.400 241.500 180.300 ;
        RECT 263.400 175.200 265.200 180.300 ;
        RECT 281.400 176.400 283.200 180.300 ;
        RECT 296.700 170.400 298.500 180.300 ;
        RECT 318.000 173.400 319.800 180.300 ;
        RECT 325.500 176.400 327.300 180.300 ;
        RECT 341.400 175.200 343.200 180.300 ;
        RECT 362.400 175.200 364.200 180.300 ;
        RECT 380.700 170.400 382.500 180.300 ;
        RECT 401.700 173.400 403.500 180.300 ;
        RECT 419.400 176.400 421.200 180.300 ;
        RECT 425.400 176.400 427.200 180.300 ;
        RECT 437.400 176.400 439.200 180.300 ;
        RECT 460.800 175.200 462.600 180.300 ;
        RECT 474.000 173.400 475.800 180.300 ;
        RECT 481.500 176.400 483.300 180.300 ;
        RECT 497.400 175.200 499.200 180.300 ;
        RECT 520.800 173.400 522.600 180.300 ;
        RECT 529.200 173.400 531.000 180.300 ;
        RECT 544.800 176.400 546.600 180.300 ;
        RECT 551.850 176.400 553.650 180.300 ;
        RECT 560.850 176.400 562.650 180.300 ;
        RECT 567.750 176.400 569.550 180.300 ;
        RECT 577.050 176.400 578.850 180.300 ;
        RECT 592.800 176.400 594.600 180.300 ;
        RECT 598.800 176.400 600.600 180.300 ;
        RECT 608.400 179.400 609.600 180.300 ;
        RECT 608.400 176.400 610.200 179.400 ;
        RECT 614.400 176.400 616.200 180.300 ;
        RECT 640.500 170.400 642.300 180.300 ;
        RECT 650.700 173.400 652.500 180.300 ;
        RECT 668.400 176.400 670.200 180.300 ;
        RECT 686.400 175.200 688.200 180.300 ;
        RECT 709.800 176.400 711.600 180.300 ;
        RECT 719.400 176.400 721.200 180.300 ;
        RECT 735.000 173.400 736.800 180.300 ;
        RECT 742.500 176.400 744.300 180.300 ;
        RECT 755.400 176.400 757.200 180.300 ;
        RECT 773.400 175.200 775.200 180.300 ;
        RECT 794.400 175.200 796.200 180.300 ;
        RECT 812.400 176.400 814.200 180.300 ;
        RECT 818.400 176.400 820.200 180.300 ;
        RECT 833.400 175.200 835.200 180.300 ;
        RECT 13.800 110.700 15.600 114.600 ;
        RECT 24.000 110.700 25.800 117.600 ;
        RECT 31.500 110.700 33.300 114.600 ;
        RECT 44.700 110.700 46.500 120.600 ;
        RECT 65.700 110.700 67.500 120.600 ;
        RECT 94.800 110.700 96.600 115.800 ;
        RECT 107.700 110.700 109.500 120.600 ;
        RECT 129.000 110.700 130.800 117.600 ;
        RECT 136.500 110.700 138.300 114.600 ;
        RECT 157.800 110.700 159.600 115.800 ;
        RECT 172.800 110.700 174.600 114.600 ;
        RECT 178.800 110.700 180.600 114.600 ;
        RECT 196.800 110.700 198.600 115.800 ;
        RECT 214.800 110.700 216.600 114.600 ;
        RECT 229.800 110.700 231.600 114.600 ;
        RECT 235.800 111.600 237.600 114.600 ;
        RECT 236.400 110.700 237.600 111.600 ;
        RECT 245.400 110.700 247.200 114.600 ;
        RECT 251.400 110.700 253.200 114.600 ;
        RECT 265.800 110.700 267.600 114.600 ;
        RECT 271.800 110.700 273.600 114.600 ;
        RECT 281.400 111.600 283.200 114.600 ;
        RECT 281.400 110.700 282.600 111.600 ;
        RECT 287.400 110.700 289.200 114.600 ;
        RECT 305.700 110.700 307.500 114.600 ;
        RECT 313.200 110.700 315.000 117.600 ;
        RECT 323.700 110.700 325.500 120.600 ;
        RECT 348.900 110.700 350.700 117.600 ;
        RECT 370.800 110.700 372.600 114.600 ;
        RECT 383.400 110.700 385.200 115.800 ;
        RECT 404.400 110.700 406.200 115.800 ;
        RECT 430.500 110.700 432.300 117.600 ;
        RECT 441.000 110.700 442.800 117.600 ;
        RECT 448.500 110.700 450.300 114.600 ;
        RECT 461.700 110.700 463.500 120.600 ;
        RECT 484.800 110.700 486.600 117.600 ;
        RECT 490.800 110.700 492.600 117.600 ;
        RECT 501.000 110.700 502.800 117.600 ;
        RECT 508.500 110.700 510.300 114.600 ;
        RECT 524.700 110.700 526.500 114.600 ;
        RECT 532.200 110.700 534.000 117.600 ;
        RECT 547.800 110.700 549.600 114.600 ;
        RECT 557.700 110.700 559.500 117.600 ;
        RECT 578.400 110.700 580.200 115.800 ;
        RECT 604.500 110.700 606.300 117.600 ;
        RECT 622.500 110.700 624.300 117.600 ;
        RECT 633.000 110.700 634.800 117.600 ;
        RECT 640.500 110.700 642.300 114.600 ;
        RECT 658.800 110.700 660.600 114.600 ;
        RECT 676.800 110.700 678.600 115.800 ;
        RECT 696.300 110.700 698.100 117.600 ;
        RECT 721.500 110.700 723.300 120.600 ;
        RECT 736.800 110.700 738.600 114.600 ;
        RECT 751.800 110.700 753.600 114.600 ;
        RECT 769.800 110.700 771.600 115.800 ;
        RECT 790.500 110.700 792.300 117.600 ;
        RECT 808.800 110.700 810.600 115.800 ;
        RECT 829.800 110.700 831.600 115.800 ;
        RECT 845.400 110.700 847.200 115.800 ;
        RECT 858.450 110.700 867.450 180.300 ;
        RECT 0.600 108.300 867.450 110.700 ;
        RECT 13.800 104.400 15.600 108.300 ;
        RECT 31.800 103.200 33.600 108.300 ;
        RECT 55.500 98.400 57.300 108.300 ;
        RECT 66.000 101.400 67.800 108.300 ;
        RECT 73.500 104.400 75.300 108.300 ;
        RECT 89.700 104.400 91.500 108.300 ;
        RECT 97.200 101.400 99.000 108.300 ;
        RECT 118.500 98.400 120.300 108.300 ;
        RECT 139.500 98.400 141.300 108.300 ;
        RECT 157.800 103.200 159.600 108.300 ;
        RECT 173.400 103.200 175.200 108.300 ;
        RECT 199.800 103.200 201.600 108.300 ;
        RECT 223.500 98.400 225.300 108.300 ;
        RECT 236.700 104.400 238.500 108.300 ;
        RECT 244.200 101.400 246.000 108.300 ;
        RECT 262.800 103.200 264.600 108.300 ;
        RECT 275.400 104.400 277.200 108.300 ;
        RECT 290.700 98.400 292.500 108.300 ;
        RECT 322.500 98.400 324.300 108.300 ;
        RECT 333.000 101.400 334.800 108.300 ;
        RECT 340.500 104.400 342.300 108.300 ;
        RECT 361.800 103.200 363.600 108.300 ;
        RECT 374.400 104.400 376.200 108.300 ;
        RECT 397.800 103.200 399.600 108.300 ;
        RECT 413.400 103.200 415.200 108.300 ;
        RECT 442.500 98.400 444.300 108.300 ;
        RECT 453.000 101.400 454.800 108.300 ;
        RECT 460.500 104.400 462.300 108.300 ;
        RECT 481.500 101.400 483.300 108.300 ;
        RECT 491.400 104.400 493.200 108.300 ;
        RECT 514.500 101.400 516.300 108.300 ;
        RECT 527.700 104.400 529.500 108.300 ;
        RECT 535.200 101.400 537.000 108.300 ;
        RECT 548.400 103.200 550.200 108.300 ;
        RECT 574.500 101.400 576.300 108.300 ;
        RECT 591.300 101.400 593.100 108.300 ;
        RECT 605.400 104.400 607.200 108.300 ;
        RECT 611.400 104.400 613.200 108.300 ;
        RECT 625.800 104.400 627.600 108.300 ;
        RECT 631.800 104.400 633.600 108.300 ;
        RECT 641.400 104.400 643.200 108.300 ;
        RECT 647.400 104.400 649.200 108.300 ;
        RECT 659.400 104.400 661.200 108.300 ;
        RECT 665.400 104.400 667.200 108.300 ;
        RECT 678.000 101.400 679.800 108.300 ;
        RECT 685.500 104.400 687.300 108.300 ;
        RECT 701.400 103.200 703.200 108.300 ;
        RECT 719.700 101.400 721.500 108.300 ;
        RECT 742.800 104.400 744.600 108.300 ;
        RECT 755.400 103.200 757.200 108.300 ;
        RECT 784.500 98.400 786.300 108.300 ;
        RECT 795.000 101.400 796.800 108.300 ;
        RECT 802.500 104.400 804.300 108.300 ;
        RECT 815.400 104.400 817.200 108.300 ;
        RECT 830.700 101.400 832.500 108.300 ;
        RECT 853.800 104.400 855.600 108.300 ;
        RECT 19.500 38.700 21.300 48.600 ;
        RECT 30.000 38.700 31.800 45.600 ;
        RECT 37.500 38.700 39.300 42.600 ;
        RECT 53.400 38.700 55.200 43.800 ;
        RECT 82.500 38.700 84.300 48.600 ;
        RECT 97.800 38.700 99.600 45.600 ;
        RECT 106.200 38.700 108.000 45.600 ;
        RECT 124.800 38.700 126.600 43.800 ;
        RECT 148.500 38.700 150.300 48.600 ;
        RECT 159.000 38.700 160.800 45.600 ;
        RECT 166.500 38.700 168.300 42.600 ;
        RECT 187.800 38.700 189.600 43.800 ;
        RECT 211.500 38.700 213.300 48.600 ;
        RECT 224.700 38.700 226.500 42.600 ;
        RECT 232.200 38.700 234.000 45.600 ;
        RECT 249.300 38.700 251.100 45.600 ;
        RECT 263.700 38.700 265.500 45.600 ;
        RECT 282.000 38.700 283.800 45.600 ;
        RECT 289.500 38.700 291.300 42.600 ;
        RECT 302.700 38.700 304.500 48.600 ;
        RECT 323.700 38.700 325.500 45.600 ;
        RECT 346.800 38.700 348.600 42.600 ;
        RECT 356.700 38.700 358.500 48.600 ;
        RECT 388.500 38.700 390.300 48.600 ;
        RECT 398.700 38.700 400.500 45.600 ;
        RECT 417.000 38.700 418.800 45.600 ;
        RECT 424.500 38.700 426.300 42.600 ;
        RECT 438.000 38.700 439.800 45.600 ;
        RECT 446.400 38.700 448.200 45.600 ;
        RECT 458.850 38.700 460.650 42.600 ;
        RECT 467.850 38.700 469.650 42.600 ;
        RECT 474.750 38.700 476.550 42.600 ;
        RECT 484.050 38.700 485.850 42.600 ;
        RECT 497.400 38.700 499.200 42.600 ;
        RECT 513.000 38.700 514.800 45.600 ;
        RECT 521.400 38.700 523.200 45.600 ;
        RECT 539.700 38.700 541.500 45.600 ;
        RECT 559.500 38.700 561.300 45.600 ;
        RECT 583.500 38.700 585.300 48.600 ;
        RECT 601.800 38.700 603.600 43.800 ;
        RECT 614.400 38.700 616.200 42.600 ;
        RECT 640.500 38.700 642.300 48.600 ;
        RECT 650.700 38.700 652.500 45.600 ;
        RECT 676.500 38.700 678.300 45.600 ;
        RECT 694.500 38.700 696.300 45.600 ;
        RECT 715.500 38.700 717.300 48.600 ;
        RECT 726.000 38.700 727.800 45.600 ;
        RECT 733.500 38.700 735.300 42.600 ;
        RECT 754.500 38.700 756.300 45.600 ;
        RECT 775.500 38.700 777.300 48.600 ;
        RECT 796.500 38.700 798.300 48.600 ;
        RECT 814.800 38.700 816.600 43.800 ;
        RECT 835.800 38.700 837.600 43.800 ;
        RECT 853.800 38.700 855.600 42.600 ;
        RECT 858.450 38.700 867.450 108.300 ;
        RECT 0.600 36.300 867.450 38.700 ;
        RECT 13.800 32.400 15.600 36.300 ;
        RECT 23.700 26.400 25.500 36.300 ;
        RECT 52.800 31.200 54.600 36.300 ;
        RECT 68.400 31.200 70.200 36.300 ;
        RECT 86.700 26.400 88.500 36.300 ;
        RECT 107.700 26.400 109.500 36.300 ;
        RECT 128.700 26.400 130.500 36.300 ;
        RECT 149.400 32.400 151.200 36.300 ;
        RECT 175.500 26.400 177.300 36.300 ;
        RECT 186.000 29.400 187.800 36.300 ;
        RECT 193.500 32.400 195.300 36.300 ;
        RECT 209.100 32.400 211.200 36.300 ;
        RECT 215.400 32.400 217.200 36.300 ;
        RECT 242.400 31.200 244.200 36.300 ;
        RECT 260.400 32.400 262.200 36.300 ;
        RECT 283.800 31.200 285.600 36.300 ;
        RECT 296.400 32.400 298.200 36.300 ;
        RECT 314.400 31.200 316.200 36.300 ;
        RECT 332.700 29.400 334.500 36.300 ;
        RECT 358.800 31.200 360.600 36.300 ;
        RECT 379.500 29.400 381.300 36.300 ;
        RECT 394.800 32.400 396.600 36.300 ;
        RECT 407.700 29.400 409.500 36.300 ;
        RECT 427.800 32.400 429.600 36.300 ;
        RECT 435.150 32.400 436.950 36.300 ;
        RECT 444.450 32.400 446.250 36.300 ;
        RECT 451.350 32.400 453.150 36.300 ;
        RECT 460.350 32.400 462.150 36.300 ;
        RECT 478.500 29.400 480.300 36.300 ;
        RECT 496.500 29.400 498.300 36.300 ;
        RECT 514.800 32.400 516.600 36.300 ;
        RECT 532.500 29.400 534.300 36.300 ;
        RECT 550.500 29.400 552.300 36.300 ;
        RECT 571.500 26.400 573.300 36.300 ;
        RECT 589.800 31.200 591.600 36.300 ;
        RECT 607.500 29.400 609.300 36.300 ;
        RECT 627.300 29.400 629.100 36.300 ;
        RECT 641.700 29.400 643.500 36.300 ;
        RECT 659.700 29.400 661.500 36.300 ;
        RECT 688.500 26.400 690.300 36.300 ;
        RECT 703.800 32.400 705.600 36.300 ;
        RECT 724.500 26.400 726.300 36.300 ;
        RECT 734.700 29.400 736.500 36.300 ;
        RECT 749.850 32.400 751.650 36.300 ;
        RECT 758.850 32.400 760.650 36.300 ;
        RECT 765.750 32.400 767.550 36.300 ;
        RECT 775.050 32.400 776.850 36.300 ;
        RECT 789.000 29.400 790.800 36.300 ;
        RECT 796.500 32.400 798.300 36.300 ;
        RECT 812.400 31.200 814.200 36.300 ;
        RECT 833.700 29.400 835.500 36.300 ;
        RECT 848.400 32.400 850.200 36.300 ;
        RECT 858.450 0.300 867.450 36.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 864.300 857.400 866.700 ;
        RECT -9.450 794.700 -0.450 864.300 ;
        RECT 13.800 858.000 15.600 864.300 ;
        RECT 19.800 857.400 21.600 864.300 ;
        RECT 29.400 857.400 31.200 864.300 ;
        RECT 35.400 858.000 37.200 864.300 ;
        RECT 53.400 853.200 55.200 864.300 ;
        RECT 72.300 851.400 74.100 864.300 ;
        RECT 79.800 857.400 81.600 864.300 ;
        RECT 95.400 857.400 97.200 864.300 ;
        RECT 102.900 851.400 104.700 864.300 ;
        RECT 118.800 857.400 120.600 864.300 ;
        RECT 133.800 858.000 135.600 864.300 ;
        RECT 139.800 857.400 141.600 864.300 ;
        RECT 150.300 851.400 152.100 864.300 ;
        RECT 157.800 857.400 159.600 864.300 ;
        RECT 173.400 853.200 175.200 864.300 ;
        RECT 196.800 857.400 198.600 864.300 ;
        RECT 206.400 857.400 208.200 864.300 ;
        RECT 212.400 858.000 214.200 864.300 ;
        RECT 232.800 858.000 234.600 864.300 ;
        RECT 238.800 857.400 240.600 864.300 ;
        RECT 251.400 857.400 253.200 864.300 ;
        RECT 258.900 851.400 260.700 864.300 ;
        RECT 274.800 857.400 276.600 864.300 ;
        RECT 287.400 857.400 289.200 864.300 ;
        RECT 294.900 851.400 296.700 864.300 ;
        RECT 305.400 857.400 307.200 864.300 ;
        RECT 327.300 851.400 329.100 864.300 ;
        RECT 349.800 851.400 351.600 864.300 ;
        RECT 362.400 857.400 364.200 864.300 ;
        RECT 369.900 851.400 371.700 864.300 ;
        RECT 385.800 857.400 387.600 864.300 ;
        RECT 396.300 851.400 398.100 864.300 ;
        RECT 403.800 857.400 405.600 864.300 ;
        RECT 424.800 853.200 426.600 864.300 ;
        RECT 437.400 857.400 439.200 864.300 ;
        RECT 443.400 857.400 445.200 864.300 ;
        RECT 459.900 851.400 461.700 864.300 ;
        RECT 481.800 858.000 483.600 864.300 ;
        RECT 487.800 857.400 489.600 864.300 ;
        RECT 502.800 857.400 504.600 864.300 ;
        RECT 514.800 857.400 516.600 864.300 ;
        RECT 520.800 857.400 522.600 864.300 ;
        RECT 530.400 851.400 532.200 864.300 ;
        RECT 536.400 851.400 538.200 864.300 ;
        RECT 542.400 851.400 544.200 864.300 ;
        RECT 548.400 851.400 550.200 864.300 ;
        RECT 554.400 851.400 556.200 864.300 ;
        RECT 562.200 857.400 564.000 864.300 ;
        RECT 568.800 857.400 570.600 864.300 ;
        RECT 574.800 857.400 576.600 864.300 ;
        RECT 580.800 857.400 582.600 864.300 ;
        RECT 597.000 857.400 598.800 864.300 ;
        RECT 603.900 857.400 605.700 864.300 ;
        RECT 616.500 859.950 618.300 864.300 ;
        RECT 622.500 857.400 624.300 864.300 ;
        RECT 628.500 858.450 630.300 864.300 ;
        RECT 628.500 857.550 633.450 858.450 ;
        RECT 628.500 857.400 630.300 857.550 ;
        RECT 632.550 850.050 633.450 857.550 ;
        RECT 640.800 857.400 642.600 864.300 ;
        RECT 646.800 857.400 648.600 864.300 ;
        RECT 652.200 857.400 654.000 864.300 ;
        RECT 658.800 857.400 660.600 864.300 ;
        RECT 664.800 857.400 666.600 864.300 ;
        RECT 670.800 857.400 672.600 864.300 ;
        RECT 687.000 857.400 688.800 864.300 ;
        RECT 693.900 857.400 695.700 864.300 ;
        RECT 706.500 859.950 708.300 864.300 ;
        RECT 712.500 859.050 714.300 864.300 ;
        RECT 712.350 856.950 714.450 859.050 ;
        RECT 718.500 857.400 720.300 864.300 ;
        RECT 731.400 857.400 733.200 864.300 ;
        RECT 738.900 851.400 740.700 864.300 ;
        RECT 757.800 851.400 759.600 864.300 ;
        RECT 767.400 857.400 769.200 864.300 ;
        RECT 787.800 857.400 789.600 864.300 ;
        RECT 794.550 860.400 796.350 864.300 ;
        RECT 803.250 857.400 805.050 864.300 ;
        RECT 809.850 857.400 811.650 864.300 ;
        RECT 820.050 857.400 821.850 864.300 ;
        RECT 833.400 851.400 835.200 864.300 ;
        RECT 631.950 847.950 634.050 850.050 ;
        RECT 16.800 794.700 18.600 805.800 ;
        RECT 34.800 794.700 36.600 801.000 ;
        RECT 40.800 794.700 42.600 801.600 ;
        RECT 53.400 794.700 55.200 801.600 ;
        RECT 60.900 794.700 62.700 807.600 ;
        RECT 74.400 794.700 76.200 801.600 ;
        RECT 81.900 794.700 83.700 807.600 ;
        RECT 97.800 794.700 99.600 801.600 ;
        RECT 107.400 794.700 109.200 801.600 ;
        RECT 113.400 794.700 115.200 801.000 ;
        RECT 136.800 794.700 138.600 805.800 ;
        RECT 156.300 794.700 158.100 807.600 ;
        RECT 170.400 794.700 172.200 801.600 ;
        RECT 176.400 794.700 178.200 801.600 ;
        RECT 199.800 794.700 201.600 805.500 ;
        RECT 212.400 794.700 214.200 801.600 ;
        RECT 218.400 794.700 220.200 801.600 ;
        RECT 230.400 794.700 232.200 801.600 ;
        RECT 236.400 794.700 238.200 801.000 ;
        RECT 251.400 794.700 253.200 801.600 ;
        RECT 257.400 794.700 259.200 801.000 ;
        RECT 274.800 794.700 276.600 801.600 ;
        RECT 280.800 794.700 282.600 801.600 ;
        RECT 295.800 794.700 297.600 801.000 ;
        RECT 301.800 794.700 303.600 801.600 ;
        RECT 311.400 794.700 313.200 801.600 ;
        RECT 317.400 794.700 319.200 801.000 ;
        RECT 332.400 794.700 334.200 801.600 ;
        RECT 338.400 794.700 340.200 801.600 ;
        RECT 355.800 794.700 357.600 801.600 ;
        RECT 365.400 794.700 367.200 801.600 ;
        RECT 371.400 794.700 373.200 801.000 ;
        RECT 386.400 794.700 388.200 801.600 ;
        RECT 406.800 794.700 408.600 801.000 ;
        RECT 412.800 794.700 414.600 801.600 ;
        RECT 427.800 794.700 429.600 801.000 ;
        RECT 433.800 794.700 435.600 801.600 ;
        RECT 445.800 794.700 447.600 801.600 ;
        RECT 451.800 794.700 453.600 801.600 ;
        RECT 468.300 794.700 470.100 807.600 ;
        RECT 482.400 794.700 484.200 801.600 ;
        RECT 488.400 794.700 490.200 801.600 ;
        RECT 503.400 794.700 505.200 801.600 ;
        RECT 510.900 794.700 512.700 807.600 ;
        RECT 523.800 794.700 525.600 801.600 ;
        RECT 529.800 794.700 531.600 801.600 ;
        RECT 542.400 794.700 544.200 801.600 ;
        RECT 549.900 794.700 551.700 807.600 ;
        RECT 562.800 794.700 564.600 801.600 ;
        RECT 568.800 794.700 570.600 801.600 ;
        RECT 586.800 794.700 588.600 805.800 ;
        RECT 604.800 794.700 606.600 801.600 ;
        RECT 619.800 794.700 621.600 801.600 ;
        RECT 629.400 794.700 631.200 801.600 ;
        RECT 635.400 794.700 637.200 801.000 ;
        RECT 655.800 794.700 657.600 801.600 ;
        RECT 666.300 794.700 668.100 807.600 ;
        RECT 673.800 794.700 675.600 801.600 ;
        RECT 687.300 794.700 689.100 807.600 ;
        RECT 694.800 794.700 696.600 801.600 ;
        RECT 708.300 794.700 710.100 807.600 ;
        RECT 715.800 794.700 717.600 801.600 ;
        RECT 733.200 794.700 735.000 807.600 ;
        RECT 739.800 794.700 741.600 801.600 ;
        RECT 749.400 794.700 751.200 807.600 ;
        RECT 767.400 794.700 769.200 807.600 ;
        RECT 789.900 794.700 791.700 807.600 ;
        RECT 806.400 794.700 808.200 807.600 ;
        RECT 816.900 794.700 818.700 807.600 ;
        RECT 841.800 794.700 843.600 805.500 ;
        RECT -9.450 792.300 857.400 794.700 ;
        RECT -9.450 722.700 -0.450 792.300 ;
        RECT 16.800 779.400 18.600 792.300 ;
        RECT 28.800 785.400 30.600 792.300 ;
        RECT 34.800 785.400 36.600 792.300 ;
        RECT 52.800 781.200 54.600 792.300 ;
        RECT 65.400 785.400 67.200 792.300 ;
        RECT 71.400 786.000 73.200 792.300 ;
        RECT 91.200 779.400 93.000 792.300 ;
        RECT 97.800 785.400 99.600 792.300 ;
        RECT 110.400 785.400 112.200 792.300 ;
        RECT 117.900 779.400 119.700 792.300 ;
        RECT 129.300 779.400 131.100 792.300 ;
        RECT 136.800 785.400 138.600 792.300 ;
        RECT 154.200 779.400 156.000 792.300 ;
        RECT 160.800 785.400 162.600 792.300 ;
        RECT 170.400 779.400 172.200 792.300 ;
        RECT 196.800 781.200 198.600 792.300 ;
        RECT 214.800 786.000 216.600 792.300 ;
        RECT 220.800 785.400 222.600 792.300 ;
        RECT 230.400 785.400 232.200 792.300 ;
        RECT 236.400 785.400 238.200 792.300 ;
        RECT 253.200 779.400 255.000 792.300 ;
        RECT 259.800 785.400 261.600 792.300 ;
        RECT 274.800 786.000 276.600 792.300 ;
        RECT 280.800 785.400 282.600 792.300 ;
        RECT 290.400 785.400 292.200 792.300 ;
        RECT 296.400 785.400 298.200 792.300 ;
        RECT 311.400 785.400 313.200 792.300 ;
        RECT 318.900 779.400 320.700 792.300 ;
        RECT 332.400 785.400 334.200 792.300 ;
        RECT 339.900 779.400 341.700 792.300 ;
        RECT 350.400 779.400 352.200 792.300 ;
        RECT 368.400 785.400 370.200 792.300 ;
        RECT 375.000 779.400 376.800 792.300 ;
        RECT 394.800 786.000 396.600 792.300 ;
        RECT 400.800 785.400 402.600 792.300 ;
        RECT 410.400 785.400 412.200 792.300 ;
        RECT 425.400 785.400 427.200 792.300 ;
        RECT 431.400 785.400 433.200 792.300 ;
        RECT 443.400 785.400 445.200 792.300 ;
        RECT 449.400 785.400 451.200 792.300 ;
        RECT 461.400 785.400 463.200 792.300 ;
        RECT 467.400 786.000 469.200 792.300 ;
        RECT 487.800 786.000 489.600 792.300 ;
        RECT 493.800 785.400 495.600 792.300 ;
        RECT 506.400 781.200 508.200 792.300 ;
        RECT 527.400 785.400 529.200 792.300 ;
        RECT 534.900 779.400 536.700 792.300 ;
        RECT 548.400 785.400 550.200 792.300 ;
        RECT 555.900 779.400 557.700 792.300 ;
        RECT 571.200 779.400 573.000 792.300 ;
        RECT 577.800 785.400 579.600 792.300 ;
        RECT 592.800 785.400 594.600 792.300 ;
        RECT 602.400 779.400 604.200 792.300 ;
        RECT 620.400 779.400 622.200 792.300 ;
        RECT 630.900 779.400 632.700 792.300 ;
        RECT 652.800 781.200 654.600 792.300 ;
        RECT 665.400 785.400 667.200 792.300 ;
        RECT 683.400 781.500 685.200 792.300 ;
        RECT 705.300 779.400 707.100 792.300 ;
        RECT 712.800 785.400 714.600 792.300 ;
        RECT 728.400 781.200 730.200 792.300 ;
        RECT 747.300 779.400 749.100 792.300 ;
        RECT 754.800 785.400 756.600 792.300 ;
        RECT 761.700 785.400 763.500 792.300 ;
        RECT 767.700 787.050 769.500 792.300 ;
        RECT 773.700 787.950 775.500 792.300 ;
        RECT 767.550 784.950 769.650 787.050 ;
        RECT 786.300 785.400 788.100 792.300 ;
        RECT 793.200 785.400 795.000 792.300 ;
        RECT 809.400 785.400 811.200 792.300 ;
        RECT 815.400 785.400 817.200 792.300 ;
        RECT 821.400 785.400 823.200 792.300 ;
        RECT 828.000 785.400 829.800 792.300 ;
        RECT 839.400 785.400 841.200 792.300 ;
        RECT 10.800 722.700 12.600 729.600 ;
        RECT 16.800 722.700 18.600 729.600 ;
        RECT 29.400 722.700 31.200 729.600 ;
        RECT 36.900 722.700 38.700 735.600 ;
        RECT 48.300 722.700 50.100 735.600 ;
        RECT 55.800 722.700 57.600 729.600 ;
        RECT 76.800 722.700 78.600 733.800 ;
        RECT 94.800 722.700 96.600 729.000 ;
        RECT 100.800 722.700 102.600 729.600 ;
        RECT 110.400 722.700 112.200 729.600 ;
        RECT 116.400 722.700 118.200 729.600 ;
        RECT 128.400 722.700 130.200 729.600 ;
        RECT 143.400 722.700 145.200 729.600 ;
        RECT 149.400 722.700 151.200 729.000 ;
        RECT 164.400 722.700 166.200 729.600 ;
        RECT 170.400 722.700 172.200 729.600 ;
        RECT 186.900 722.700 188.700 735.600 ;
        RECT 205.800 722.700 207.600 729.600 ;
        RECT 211.800 722.700 213.600 729.600 ;
        RECT 229.800 722.700 231.600 735.600 ;
        RECT 241.800 722.700 243.600 729.600 ;
        RECT 247.800 722.700 249.600 729.600 ;
        RECT 257.400 722.700 259.200 729.600 ;
        RECT 277.800 722.700 279.600 729.000 ;
        RECT 283.800 722.700 285.600 729.600 ;
        RECT 300.300 722.700 302.100 735.600 ;
        RECT 314.400 722.700 316.200 729.600 ;
        RECT 320.400 722.700 322.200 729.600 ;
        RECT 332.400 722.700 334.200 735.600 ;
        RECT 353.400 722.700 355.200 729.600 ;
        RECT 360.900 722.700 362.700 735.600 ;
        RECT 371.400 722.700 373.200 729.600 ;
        RECT 391.800 722.700 393.600 729.600 ;
        RECT 401.400 722.700 403.200 735.600 ;
        RECT 419.400 722.700 421.200 729.600 ;
        RECT 425.400 722.700 427.200 729.600 ;
        RECT 440.400 722.700 442.200 729.600 ;
        RECT 447.900 722.700 449.700 735.600 ;
        RECT 458.400 722.700 460.200 729.600 ;
        RECT 464.400 722.700 466.200 729.600 ;
        RECT 479.400 722.700 481.200 729.600 ;
        RECT 486.900 722.700 488.700 735.600 ;
        RECT 502.800 722.700 504.600 729.600 ;
        RECT 516.300 722.700 518.100 735.600 ;
        RECT 526.800 722.700 528.600 735.600 ;
        RECT 536.400 722.700 538.200 729.600 ;
        RECT 542.400 722.700 544.200 729.600 ;
        RECT 556.800 722.700 558.600 735.600 ;
        RECT 562.800 722.700 564.600 735.600 ;
        RECT 572.400 722.700 574.200 735.600 ;
        RECT 590.400 722.700 592.200 735.600 ;
        RECT 611.400 722.700 613.200 729.600 ;
        RECT 618.900 722.700 620.700 735.600 ;
        RECT 629.400 722.700 631.200 729.600 ;
        RECT 649.800 722.700 651.600 729.600 ;
        RECT 659.400 722.700 661.200 735.600 ;
        RECT 677.400 722.700 679.200 735.600 ;
        RECT 697.800 722.700 699.600 729.600 ;
        RECT 703.800 722.700 705.600 729.600 ;
        RECT 710.550 722.700 712.350 726.600 ;
        RECT 719.250 722.700 721.050 729.600 ;
        RECT 725.850 722.700 727.650 729.600 ;
        RECT 736.050 722.700 737.850 729.600 ;
        RECT 749.400 722.700 751.200 729.600 ;
        RECT 755.400 722.700 757.200 729.600 ;
        RECT 770.400 722.700 772.200 729.600 ;
        RECT 777.900 722.700 779.700 735.600 ;
        RECT 793.800 722.700 795.600 729.600 ;
        RECT 806.700 722.700 808.500 735.600 ;
        RECT 822.300 722.700 824.100 735.600 ;
        RECT 829.800 722.700 831.600 729.600 ;
        RECT 842.400 722.700 844.200 729.600 ;
        RECT 848.400 722.700 850.200 729.600 ;
        RECT -9.450 720.300 857.400 722.700 ;
        RECT -9.450 650.700 -0.450 720.300 ;
        RECT 13.800 714.000 15.600 720.300 ;
        RECT 19.800 713.400 21.600 720.300 ;
        RECT 32.400 709.200 34.200 720.300 ;
        RECT 51.300 707.400 53.100 720.300 ;
        RECT 58.800 713.400 60.600 720.300 ;
        RECT 72.300 707.400 74.100 720.300 ;
        RECT 79.800 713.400 81.600 720.300 ;
        RECT 92.400 713.400 94.200 720.300 ;
        RECT 98.400 714.000 100.200 720.300 ;
        RECT 113.400 713.400 115.200 720.300 ;
        RECT 119.400 714.000 121.200 720.300 ;
        RECT 137.400 709.200 139.200 720.300 ;
        RECT 156.300 707.400 158.100 720.300 ;
        RECT 163.800 713.400 165.600 720.300 ;
        RECT 178.800 713.400 180.600 720.300 ;
        RECT 184.800 713.400 186.600 720.300 ;
        RECT 194.400 713.400 196.200 720.300 ;
        RECT 200.400 714.000 202.200 720.300 ;
        RECT 223.800 707.400 225.600 720.300 ;
        RECT 238.800 714.000 240.600 720.300 ;
        RECT 244.800 713.400 246.600 720.300 ;
        RECT 254.400 707.400 256.200 720.300 ;
        RECT 264.900 707.400 266.700 720.300 ;
        RECT 283.800 714.000 285.600 720.300 ;
        RECT 289.800 713.400 291.600 720.300 ;
        RECT 307.800 709.200 309.600 720.300 ;
        RECT 320.400 713.400 322.200 720.300 ;
        RECT 335.400 713.400 337.200 720.300 ;
        RECT 351.300 707.400 353.100 720.300 ;
        RECT 358.800 713.400 360.600 720.300 ;
        RECT 376.800 707.400 378.600 720.300 ;
        RECT 386.400 713.400 388.200 720.300 ;
        RECT 392.400 713.400 394.200 720.300 ;
        RECT 408.300 707.400 410.100 720.300 ;
        RECT 418.800 707.400 420.600 720.300 ;
        RECT 430.800 713.400 432.600 720.300 ;
        RECT 436.800 713.400 438.600 720.300 ;
        RECT 450.900 707.400 452.700 720.300 ;
        RECT 472.800 713.400 474.600 720.300 ;
        RECT 482.400 713.400 484.200 720.300 ;
        RECT 488.400 714.000 490.200 720.300 ;
        RECT 503.400 713.400 505.200 720.300 ;
        RECT 509.400 713.400 511.200 720.300 ;
        RECT 526.800 707.400 528.600 720.300 ;
        RECT 536.400 713.400 538.200 720.300 ;
        RECT 551.400 707.400 553.200 720.300 ;
        RECT 571.800 713.400 573.600 720.300 ;
        RECT 577.800 713.400 579.600 720.300 ;
        RECT 587.400 707.400 589.200 720.300 ;
        RECT 605.400 707.400 607.200 720.300 ;
        RECT 623.400 713.400 625.200 720.300 ;
        RECT 629.400 713.400 631.200 720.300 ;
        RECT 639.150 713.400 640.950 720.300 ;
        RECT 649.350 713.400 651.150 720.300 ;
        RECT 655.950 713.400 657.750 720.300 ;
        RECT 664.650 716.400 666.450 720.300 ;
        RECT 677.400 713.400 679.200 720.300 ;
        RECT 683.400 713.400 685.200 720.300 ;
        RECT 695.400 713.400 697.200 720.300 ;
        RECT 707.550 716.400 709.350 720.300 ;
        RECT 716.250 713.400 718.050 720.300 ;
        RECT 722.850 713.400 724.650 720.300 ;
        RECT 733.050 713.400 734.850 720.300 ;
        RECT 746.400 713.400 748.200 720.300 ;
        RECT 752.400 713.400 754.200 720.300 ;
        RECT 767.400 713.400 769.200 720.300 ;
        RECT 774.900 707.400 776.700 720.300 ;
        RECT 790.500 707.400 792.300 720.300 ;
        RECT 808.800 713.400 810.600 720.300 ;
        RECT 816.150 713.400 817.950 720.300 ;
        RECT 826.350 713.400 828.150 720.300 ;
        RECT 832.950 713.400 834.750 720.300 ;
        RECT 841.650 716.400 843.450 720.300 ;
        RECT 11.400 650.700 13.200 657.600 ;
        RECT 18.900 650.700 20.700 663.600 ;
        RECT 37.800 650.700 39.600 661.800 ;
        RECT 58.800 650.700 60.600 663.600 ;
        RECT 70.800 650.700 72.600 657.600 ;
        RECT 76.800 650.700 78.600 657.600 ;
        RECT 91.800 650.700 93.600 657.000 ;
        RECT 97.800 650.700 99.600 657.600 ;
        RECT 107.400 650.700 109.200 657.600 ;
        RECT 113.400 650.700 115.200 657.000 ;
        RECT 128.400 650.700 130.200 657.600 ;
        RECT 143.400 650.700 145.200 657.600 ;
        RECT 149.400 650.700 151.200 657.000 ;
        RECT 164.400 650.700 166.200 657.600 ;
        RECT 170.400 650.700 172.200 657.000 ;
        RECT 185.400 650.700 187.200 657.600 ;
        RECT 191.400 650.700 193.200 657.000 ;
        RECT 206.400 650.700 208.200 657.600 ;
        RECT 212.400 650.700 214.200 657.600 ;
        RECT 224.400 650.700 226.200 657.600 ;
        RECT 241.800 650.700 243.600 657.600 ;
        RECT 247.800 650.700 249.600 657.600 ;
        RECT 257.400 650.700 259.200 663.600 ;
        RECT 280.800 650.700 282.600 661.800 ;
        RECT 298.800 650.700 300.600 657.000 ;
        RECT 304.800 650.700 306.600 657.600 ;
        RECT 314.400 650.700 316.200 657.600 ;
        RECT 320.400 650.700 322.200 657.600 ;
        RECT 335.400 650.700 337.200 657.600 ;
        RECT 342.900 650.700 344.700 663.600 ;
        RECT 355.800 650.700 357.600 657.600 ;
        RECT 361.800 650.700 363.600 657.600 ;
        RECT 376.200 650.700 378.000 663.600 ;
        RECT 382.800 650.700 384.600 657.600 ;
        RECT 403.800 650.700 405.600 661.500 ;
        RECT 416.400 650.700 418.200 657.600 ;
        RECT 422.400 650.700 424.200 657.600 ;
        RECT 437.400 650.700 439.200 663.600 ;
        RECT 458.700 650.700 460.500 663.600 ;
        RECT 473.400 650.700 475.200 657.600 ;
        RECT 479.400 650.700 481.200 657.600 ;
        RECT 491.400 650.700 493.200 663.600 ;
        RECT 507.300 650.700 509.100 663.600 ;
        RECT 514.800 650.700 516.600 657.600 ;
        RECT 531.900 650.700 533.700 663.600 ;
        RECT 549.300 650.700 551.100 663.600 ;
        RECT 556.800 650.700 558.600 657.600 ;
        RECT 571.800 650.700 573.600 657.600 ;
        RECT 577.800 650.700 579.600 657.600 ;
        RECT 592.500 650.700 594.300 663.600 ;
        RECT 608.700 650.700 610.500 663.600 ;
        RECT 625.800 650.700 627.600 657.600 ;
        RECT 631.800 650.700 633.600 657.600 ;
        RECT 644.400 650.700 646.200 657.600 ;
        RECT 651.900 650.700 653.700 663.600 ;
        RECT 662.400 650.700 664.200 663.600 ;
        RECT 668.400 650.700 670.200 663.600 ;
        RECT 674.400 650.700 676.200 663.600 ;
        RECT 680.400 650.700 682.200 663.600 ;
        RECT 686.400 650.700 688.200 663.600 ;
        RECT 695.550 650.700 697.350 654.600 ;
        RECT 704.250 650.700 706.050 657.600 ;
        RECT 710.850 650.700 712.650 657.600 ;
        RECT 721.050 650.700 722.850 657.600 ;
        RECT 737.400 650.700 739.200 657.600 ;
        RECT 744.900 650.700 746.700 663.600 ;
        RECT 755.400 650.700 757.200 657.600 ;
        RECT 761.400 650.700 763.200 657.600 ;
        RECT 776.700 650.700 778.500 663.600 ;
        RECT 788.550 650.700 790.350 654.600 ;
        RECT 797.250 650.700 799.050 657.600 ;
        RECT 803.850 650.700 805.650 657.600 ;
        RECT 814.050 650.700 815.850 657.600 ;
        RECT 828.300 650.700 830.100 663.600 ;
        RECT 835.800 650.700 837.600 657.600 ;
        RECT -9.450 648.300 857.400 650.700 ;
        RECT -9.450 578.700 -0.450 648.300 ;
        RECT 16.800 637.200 18.600 648.300 ;
        RECT 34.800 642.000 36.600 648.300 ;
        RECT 40.800 641.400 42.600 648.300 ;
        RECT 52.800 641.400 54.600 648.300 ;
        RECT 58.800 641.400 60.600 648.300 ;
        RECT 73.800 642.000 75.600 648.300 ;
        RECT 79.800 641.400 81.600 648.300 ;
        RECT 92.400 641.400 94.200 648.300 ;
        RECT 99.900 635.400 101.700 648.300 ;
        RECT 121.800 637.500 123.600 648.300 ;
        RECT 134.400 641.400 136.200 648.300 ;
        RECT 140.400 641.400 142.200 648.300 ;
        RECT 152.400 641.400 154.200 648.300 ;
        RECT 159.000 635.400 160.800 648.300 ;
        RECT 178.800 642.000 180.600 648.300 ;
        RECT 184.800 641.400 186.600 648.300 ;
        RECT 199.800 641.400 201.600 648.300 ;
        RECT 214.800 641.400 216.600 648.300 ;
        RECT 227.400 641.400 229.200 648.300 ;
        RECT 234.900 635.400 236.700 648.300 ;
        RECT 250.800 642.000 252.600 648.300 ;
        RECT 256.800 641.400 258.600 648.300 ;
        RECT 266.400 641.400 268.200 648.300 ;
        RECT 272.400 641.400 274.200 648.300 ;
        RECT 287.400 641.400 289.200 648.300 ;
        RECT 294.900 635.400 296.700 648.300 ;
        RECT 305.400 641.400 307.200 648.300 ;
        RECT 311.400 641.400 313.200 648.300 ;
        RECT 326.400 641.400 328.200 648.300 ;
        RECT 333.900 635.400 335.700 648.300 ;
        RECT 345.300 635.400 347.100 648.300 ;
        RECT 352.800 641.400 354.600 648.300 ;
        RECT 370.200 635.400 372.000 648.300 ;
        RECT 376.800 641.400 378.600 648.300 ;
        RECT 389.400 637.500 391.200 648.300 ;
        RECT 413.400 637.500 415.200 648.300 ;
        RECT 434.400 641.400 436.200 648.300 ;
        RECT 451.800 641.400 453.600 648.300 ;
        RECT 457.800 641.400 459.600 648.300 ;
        RECT 472.200 635.400 474.000 648.300 ;
        RECT 478.800 641.400 480.600 648.300 ;
        RECT 491.400 641.400 493.200 648.300 ;
        RECT 498.900 635.400 500.700 648.300 ;
        RECT 510.300 635.400 512.100 648.300 ;
        RECT 517.800 641.400 519.600 648.300 ;
        RECT 535.800 641.400 537.600 648.300 ;
        RECT 547.800 641.400 549.600 648.300 ;
        RECT 553.800 641.400 555.600 648.300 ;
        RECT 563.400 641.400 565.200 648.300 ;
        RECT 569.400 641.400 571.200 648.300 ;
        RECT 583.800 641.400 585.600 648.300 ;
        RECT 589.800 641.400 591.600 648.300 ;
        RECT 599.400 641.400 601.200 648.300 ;
        RECT 617.700 635.400 619.500 648.300 ;
        RECT 632.400 641.400 634.200 648.300 ;
        RECT 638.400 641.400 640.200 648.300 ;
        RECT 653.400 641.400 655.200 648.300 ;
        RECT 660.900 635.400 662.700 648.300 ;
        RECT 668.550 644.400 670.350 648.300 ;
        RECT 677.250 641.400 679.050 648.300 ;
        RECT 683.850 641.400 685.650 648.300 ;
        RECT 694.050 641.400 695.850 648.300 ;
        RECT 712.500 635.400 714.300 648.300 ;
        RECT 723.150 641.400 724.950 648.300 ;
        RECT 733.350 641.400 735.150 648.300 ;
        RECT 739.950 641.400 741.750 648.300 ;
        RECT 748.650 644.400 750.450 648.300 ;
        RECT 764.700 635.400 766.500 648.300 ;
        RECT 780.300 635.400 782.100 648.300 ;
        RECT 787.800 641.400 789.600 648.300 ;
        RECT 800.400 641.400 802.200 648.300 ;
        RECT 806.400 641.400 808.200 648.300 ;
        RECT 820.800 641.400 822.600 648.300 ;
        RECT 826.800 641.400 828.600 648.300 ;
        RECT 837.300 635.400 839.100 648.300 ;
        RECT 844.800 641.400 846.600 648.300 ;
        RECT 13.800 578.700 15.600 585.000 ;
        RECT 19.800 578.700 21.600 585.600 ;
        RECT 32.400 578.700 34.200 589.800 ;
        RECT 50.400 578.700 52.200 585.600 ;
        RECT 56.400 578.700 58.200 585.000 ;
        RECT 72.300 578.700 74.100 591.600 ;
        RECT 79.800 578.700 81.600 585.600 ;
        RECT 92.400 578.700 94.200 585.600 ;
        RECT 98.400 578.700 100.200 585.600 ;
        RECT 110.400 578.700 112.200 591.600 ;
        RECT 128.400 578.700 130.200 585.600 ;
        RECT 134.400 578.700 136.200 585.600 ;
        RECT 148.800 578.700 150.600 585.600 ;
        RECT 154.800 578.700 156.600 585.600 ;
        RECT 169.800 578.700 171.600 585.000 ;
        RECT 175.800 578.700 177.600 585.600 ;
        RECT 188.400 578.700 190.200 589.800 ;
        RECT 214.800 578.700 216.600 589.800 ;
        RECT 228.300 578.700 230.100 591.600 ;
        RECT 235.800 578.700 237.600 585.600 ;
        RECT 248.400 578.700 250.200 585.600 ;
        RECT 263.400 578.700 265.200 585.600 ;
        RECT 269.400 578.700 271.200 585.600 ;
        RECT 286.200 578.700 288.000 591.600 ;
        RECT 292.800 578.700 294.600 585.600 ;
        RECT 302.400 578.700 304.200 591.600 ;
        RECT 328.800 578.700 330.600 589.500 ;
        RECT 346.500 578.700 348.300 591.600 ;
        RECT 362.700 578.700 364.500 591.600 ;
        RECT 382.500 578.700 384.300 591.600 ;
        RECT 397.800 578.700 399.600 585.600 ;
        RECT 403.800 578.700 405.600 585.600 ;
        RECT 420.300 578.700 422.100 591.600 ;
        RECT 441.300 578.700 443.100 591.600 ;
        RECT 463.800 578.700 465.600 589.800 ;
        RECT 481.800 578.700 483.600 585.000 ;
        RECT 487.800 578.700 489.600 585.600 ;
        RECT 502.800 578.700 504.600 585.600 ;
        RECT 517.800 578.700 519.600 585.000 ;
        RECT 523.800 578.700 525.600 585.600 ;
        RECT 536.400 578.700 538.200 589.800 ;
        RECT 555.300 578.700 557.100 591.600 ;
        RECT 562.800 578.700 564.600 585.600 ;
        RECT 575.400 578.700 577.200 591.600 ;
        RECT 594.300 578.700 596.100 591.600 ;
        RECT 601.800 578.700 603.600 585.600 ;
        RECT 614.400 578.700 616.200 591.600 ;
        RECT 620.400 578.700 622.200 591.600 ;
        RECT 626.400 578.700 628.200 591.600 ;
        RECT 632.400 578.700 634.200 591.600 ;
        RECT 638.400 578.700 640.200 591.600 ;
        RECT 652.800 578.700 654.600 585.600 ;
        RECT 658.800 578.700 660.600 585.600 ;
        RECT 671.400 578.700 673.200 585.600 ;
        RECT 678.900 578.700 680.700 591.600 ;
        RECT 689.400 578.700 691.200 585.600 ;
        RECT 695.400 578.700 697.200 585.600 ;
        RECT 710.400 578.700 712.200 585.600 ;
        RECT 717.900 578.700 719.700 591.600 ;
        RECT 729.300 578.700 731.100 591.600 ;
        RECT 736.800 578.700 738.600 585.600 ;
        RECT 749.400 578.700 751.200 585.600 ;
        RECT 755.400 578.700 757.200 585.600 ;
        RECT 768.300 578.700 770.100 591.600 ;
        RECT 775.800 578.700 777.600 585.600 ;
        RECT 788.400 578.700 790.200 585.600 ;
        RECT 794.400 578.700 796.200 585.600 ;
        RECT 811.800 578.700 813.600 585.600 ;
        RECT 821.400 578.700 823.200 591.600 ;
        RECT 827.400 578.700 829.200 591.600 ;
        RECT 842.700 578.700 844.500 591.600 ;
        RECT -9.450 576.300 857.400 578.700 ;
        RECT -9.450 506.700 -0.450 576.300 ;
        RECT 13.500 563.400 15.300 576.300 ;
        RECT 29.400 569.400 31.200 576.300 ;
        RECT 36.900 563.400 38.700 576.300 ;
        RECT 50.400 569.400 52.200 576.300 ;
        RECT 57.900 563.400 59.700 576.300 ;
        RECT 71.400 566.400 73.200 576.300 ;
        RECT 109.800 565.200 111.600 576.300 ;
        RECT 127.800 570.000 129.600 576.300 ;
        RECT 133.800 569.400 135.600 576.300 ;
        RECT 154.800 565.500 156.600 576.300 ;
        RECT 172.200 563.400 174.000 576.300 ;
        RECT 178.800 569.400 180.600 576.300 ;
        RECT 193.800 570.000 195.600 576.300 ;
        RECT 199.800 569.400 201.600 576.300 ;
        RECT 214.800 569.400 216.600 576.300 ;
        RECT 227.400 569.400 229.200 576.300 ;
        RECT 234.900 563.400 236.700 576.300 ;
        RECT 248.400 569.400 250.200 576.300 ;
        RECT 255.900 563.400 257.700 576.300 ;
        RECT 273.300 563.400 275.100 576.300 ;
        RECT 287.400 563.400 289.200 576.300 ;
        RECT 305.400 569.400 307.200 576.300 ;
        RECT 311.400 569.400 313.200 576.300 ;
        RECT 323.400 569.400 325.200 576.300 ;
        RECT 330.000 563.400 331.800 576.300 ;
        RECT 352.800 563.400 354.600 576.300 ;
        RECT 362.400 569.400 364.200 576.300 ;
        RECT 368.400 569.400 370.200 576.300 ;
        RECT 380.400 569.400 382.200 576.300 ;
        RECT 397.800 569.400 399.600 576.300 ;
        RECT 403.800 569.400 405.600 576.300 ;
        RECT 421.800 565.200 423.600 576.300 ;
        RECT 436.800 569.400 438.600 576.300 ;
        RECT 442.800 569.400 444.600 576.300 ;
        RECT 455.400 565.500 457.200 576.300 ;
        RECT 476.400 563.400 478.200 576.300 ;
        RECT 495.300 563.400 497.100 576.300 ;
        RECT 502.800 569.400 504.600 576.300 ;
        RECT 523.800 563.400 525.600 576.300 ;
        RECT 533.400 569.400 535.200 576.300 ;
        RECT 539.400 570.000 541.200 576.300 ;
        RECT 554.400 569.400 556.200 576.300 ;
        RECT 560.400 570.000 562.200 576.300 ;
        RECT 575.400 569.400 577.200 576.300 ;
        RECT 581.400 570.000 583.200 576.300 ;
        RECT 596.400 569.400 598.200 576.300 ;
        RECT 603.000 563.400 604.800 576.300 ;
        RECT 618.300 563.400 620.100 576.300 ;
        RECT 625.800 569.400 627.600 576.300 ;
        RECT 635.550 572.400 637.350 576.300 ;
        RECT 644.250 569.400 646.050 576.300 ;
        RECT 650.850 569.400 652.650 576.300 ;
        RECT 661.050 569.400 662.850 576.300 ;
        RECT 671.550 572.400 673.350 576.300 ;
        RECT 680.250 569.400 682.050 576.300 ;
        RECT 686.850 569.400 688.650 576.300 ;
        RECT 697.050 569.400 698.850 576.300 ;
        RECT 707.550 572.400 709.350 576.300 ;
        RECT 716.250 569.400 718.050 576.300 ;
        RECT 722.850 569.400 724.650 576.300 ;
        RECT 733.050 569.400 734.850 576.300 ;
        RECT 747.300 563.400 749.100 576.300 ;
        RECT 754.800 569.400 756.600 576.300 ;
        RECT 767.400 569.400 769.200 576.300 ;
        RECT 773.400 569.400 775.200 576.300 ;
        RECT 785.400 569.400 787.200 576.300 ;
        RECT 797.550 572.400 799.350 576.300 ;
        RECT 806.250 569.400 808.050 576.300 ;
        RECT 812.850 569.400 814.650 576.300 ;
        RECT 823.050 569.400 824.850 576.300 ;
        RECT 836.400 569.400 838.200 576.300 ;
        RECT 16.800 506.700 18.600 517.800 ;
        RECT 29.400 506.700 31.200 513.600 ;
        RECT 35.400 506.700 37.200 513.000 ;
        RECT 50.400 506.700 52.200 513.600 ;
        RECT 56.400 506.700 58.200 513.000 ;
        RECT 74.400 506.700 76.200 517.800 ;
        RECT 93.300 506.700 95.100 519.600 ;
        RECT 100.800 506.700 102.600 513.600 ;
        RECT 113.400 506.700 115.200 513.600 ;
        RECT 119.400 506.700 121.200 513.000 ;
        RECT 137.400 506.700 139.200 517.800 ;
        RECT 160.800 506.700 162.600 513.600 ;
        RECT 173.400 506.700 175.200 517.500 ;
        RECT 194.400 506.700 196.200 513.600 ;
        RECT 200.400 506.700 202.200 513.000 ;
        RECT 217.800 506.700 219.600 513.600 ;
        RECT 223.800 506.700 225.600 513.600 ;
        RECT 238.200 506.700 240.000 519.600 ;
        RECT 244.800 506.700 246.600 513.600 ;
        RECT 257.400 506.700 259.200 517.500 ;
        RECT 280.800 506.700 282.600 513.600 ;
        RECT 286.800 506.700 288.600 513.600 ;
        RECT 296.400 506.700 298.200 519.600 ;
        RECT 317.400 506.700 319.200 513.600 ;
        RECT 324.900 506.700 326.700 519.600 ;
        RECT 335.400 506.700 337.200 513.600 ;
        RECT 350.400 506.700 352.200 513.600 ;
        RECT 356.400 506.700 358.200 513.600 ;
        RECT 371.400 506.700 373.200 517.800 ;
        RECT 389.400 506.700 391.200 513.600 ;
        RECT 404.400 506.700 406.200 519.600 ;
        RECT 423.300 506.700 425.100 519.600 ;
        RECT 430.800 506.700 432.600 513.600 ;
        RECT 443.400 506.700 445.200 513.600 ;
        RECT 458.400 506.700 460.200 513.600 ;
        RECT 464.400 506.700 466.200 513.000 ;
        RECT 482.400 506.700 484.200 517.800 ;
        RECT 500.400 506.700 502.200 513.600 ;
        RECT 518.400 506.700 520.200 517.800 ;
        RECT 536.400 506.700 538.200 513.600 ;
        RECT 542.400 506.700 544.200 513.000 ;
        RECT 558.300 506.700 560.100 519.600 ;
        RECT 565.800 506.700 567.600 513.600 ;
        RECT 580.800 506.700 582.600 519.600 ;
        RECT 586.800 506.700 588.600 519.600 ;
        RECT 592.800 506.700 594.600 519.600 ;
        RECT 598.800 506.700 600.600 519.600 ;
        RECT 604.800 506.700 606.600 519.600 ;
        RECT 616.800 506.700 618.600 519.600 ;
        RECT 622.800 506.700 624.600 519.600 ;
        RECT 628.800 506.700 630.600 519.600 ;
        RECT 634.800 506.700 636.600 519.600 ;
        RECT 640.800 506.700 642.600 519.600 ;
        RECT 651.300 506.700 653.100 519.600 ;
        RECT 658.800 506.700 660.600 513.600 ;
        RECT 671.400 506.700 673.200 513.600 ;
        RECT 677.400 506.700 679.200 513.600 ;
        RECT 690.300 506.700 692.100 519.600 ;
        RECT 697.800 506.700 699.600 513.600 ;
        RECT 710.400 506.700 712.200 513.600 ;
        RECT 716.400 506.700 718.200 513.600 ;
        RECT 725.550 506.700 727.350 510.600 ;
        RECT 734.250 506.700 736.050 513.600 ;
        RECT 740.850 506.700 742.650 513.600 ;
        RECT 751.050 506.700 752.850 513.600 ;
        RECT 767.400 506.700 769.200 517.800 ;
        RECT 786.300 506.700 788.100 519.600 ;
        RECT 793.800 506.700 795.600 513.600 ;
        RECT 806.400 506.700 808.200 513.600 ;
        RECT 822.300 506.700 824.100 519.600 ;
        RECT 829.800 506.700 831.600 513.600 ;
        RECT 842.400 506.700 844.200 513.600 ;
        RECT 848.400 506.700 850.200 513.600 ;
        RECT -9.450 504.300 857.400 506.700 ;
        RECT -9.450 434.700 -0.450 504.300 ;
        RECT 11.400 497.400 13.200 504.300 ;
        RECT 18.900 491.400 20.700 504.300 ;
        RECT 30.300 491.400 32.100 504.300 ;
        RECT 37.800 497.400 39.600 504.300 ;
        RECT 50.400 497.400 52.200 504.300 ;
        RECT 56.400 498.000 58.200 504.300 ;
        RECT 76.800 498.000 78.600 504.300 ;
        RECT 82.800 497.400 84.600 504.300 ;
        RECT 95.400 493.200 97.200 504.300 ;
        RECT 118.800 497.400 120.600 504.300 ;
        RECT 131.400 493.200 133.200 504.300 ;
        RECT 150.300 491.400 152.100 504.300 ;
        RECT 157.800 497.400 159.600 504.300 ;
        RECT 170.400 497.400 172.200 504.300 ;
        RECT 176.400 498.000 178.200 504.300 ;
        RECT 194.400 497.400 196.200 504.300 ;
        RECT 201.900 491.400 203.700 504.300 ;
        RECT 217.800 497.400 219.600 504.300 ;
        RECT 232.500 491.400 234.300 504.300 ;
        RECT 250.800 498.000 252.600 504.300 ;
        RECT 256.800 497.400 258.600 504.300 ;
        RECT 271.800 497.400 273.600 504.300 ;
        RECT 281.400 497.400 283.200 504.300 ;
        RECT 288.000 491.400 289.800 504.300 ;
        RECT 302.400 497.400 304.200 504.300 ;
        RECT 308.400 497.400 310.200 504.300 ;
        RECT 322.800 497.400 324.600 504.300 ;
        RECT 328.800 497.400 330.600 504.300 ;
        RECT 340.800 497.400 342.600 504.300 ;
        RECT 346.800 497.400 348.600 504.300 ;
        RECT 356.400 497.400 358.200 504.300 ;
        RECT 362.400 498.000 364.200 504.300 ;
        RECT 380.400 493.200 382.200 504.300 ;
        RECT 401.400 497.400 403.200 504.300 ;
        RECT 408.900 491.400 410.700 504.300 ;
        RECT 427.800 491.400 429.600 504.300 ;
        RECT 442.800 497.400 444.600 504.300 ;
        RECT 455.400 493.200 457.200 504.300 ;
        RECT 476.400 494.400 478.200 504.300 ;
        RECT 511.800 497.400 513.600 504.300 ;
        RECT 522.300 491.400 524.100 504.300 ;
        RECT 529.800 497.400 531.600 504.300 ;
        RECT 539.550 500.400 541.350 504.300 ;
        RECT 548.250 497.400 550.050 504.300 ;
        RECT 554.850 497.400 556.650 504.300 ;
        RECT 565.050 497.400 566.850 504.300 ;
        RECT 575.550 500.400 577.350 504.300 ;
        RECT 584.250 497.400 586.050 504.300 ;
        RECT 590.850 497.400 592.650 504.300 ;
        RECT 601.050 497.400 602.850 504.300 ;
        RECT 616.800 497.400 618.600 504.300 ;
        RECT 622.800 497.400 624.600 504.300 ;
        RECT 635.400 497.400 637.200 504.300 ;
        RECT 642.900 491.400 644.700 504.300 ;
        RECT 653.400 497.400 655.200 504.300 ;
        RECT 673.800 497.400 675.600 504.300 ;
        RECT 685.800 497.400 687.600 504.300 ;
        RECT 691.800 497.400 693.600 504.300 ;
        RECT 703.800 497.400 705.600 504.300 ;
        RECT 709.800 497.400 711.600 504.300 ;
        RECT 722.400 493.500 724.200 504.300 ;
        RECT 746.400 497.400 748.200 504.300 ;
        RECT 753.900 491.400 755.700 504.300 ;
        RECT 769.800 497.400 771.600 504.300 ;
        RECT 787.800 491.400 789.600 504.300 ;
        RECT 798.300 491.400 800.100 504.300 ;
        RECT 805.800 497.400 807.600 504.300 ;
        RECT 821.400 497.400 823.200 504.300 ;
        RECT 828.900 491.400 830.700 504.300 ;
        RECT 847.800 491.400 849.600 504.300 ;
        RECT 13.200 434.700 15.000 447.600 ;
        RECT 19.800 434.700 21.600 441.600 ;
        RECT 29.400 434.700 31.200 441.600 ;
        RECT 35.400 434.700 37.200 441.600 ;
        RECT 52.800 434.700 54.600 441.000 ;
        RECT 58.800 434.700 60.600 441.600 ;
        RECT 76.800 434.700 78.600 445.800 ;
        RECT 94.800 434.700 96.600 441.000 ;
        RECT 100.800 434.700 102.600 441.600 ;
        RECT 110.400 434.700 112.200 441.600 ;
        RECT 128.400 434.700 130.200 441.600 ;
        RECT 135.900 434.700 137.700 447.600 ;
        RECT 154.800 434.700 156.600 447.600 ;
        RECT 164.400 434.700 166.200 441.600 ;
        RECT 170.400 434.700 172.200 441.600 ;
        RECT 187.800 434.700 189.600 441.000 ;
        RECT 193.800 434.700 195.600 441.600 ;
        RECT 203.400 434.700 205.200 441.600 ;
        RECT 209.400 434.700 211.200 441.600 ;
        RECT 224.400 434.700 226.200 445.500 ;
        RECT 250.500 434.700 252.300 447.600 ;
        RECT 268.800 434.700 270.600 441.000 ;
        RECT 274.800 434.700 276.600 441.600 ;
        RECT 285.300 434.700 287.100 447.600 ;
        RECT 292.800 434.700 294.600 441.600 ;
        RECT 308.400 434.700 310.200 441.600 ;
        RECT 315.900 434.700 317.700 447.600 ;
        RECT 326.400 434.700 328.200 441.600 ;
        RECT 333.000 434.700 334.800 447.600 ;
        RECT 347.400 434.700 349.200 441.600 ;
        RECT 354.000 434.700 355.800 447.600 ;
        RECT 370.800 434.700 372.600 441.600 ;
        RECT 376.800 434.700 378.600 441.600 ;
        RECT 389.400 434.700 391.200 441.600 ;
        RECT 396.900 434.700 398.700 447.600 ;
        RECT 408.300 434.700 410.100 447.600 ;
        RECT 415.800 434.700 417.600 441.600 ;
        RECT 429.300 434.700 431.100 447.600 ;
        RECT 436.800 434.700 438.600 441.600 ;
        RECT 454.800 434.700 456.600 441.600 ;
        RECT 465.300 434.700 467.100 447.600 ;
        RECT 472.800 434.700 474.600 441.600 ;
        RECT 486.300 434.700 488.100 447.600 ;
        RECT 493.800 434.700 495.600 441.600 ;
        RECT 507.300 434.700 509.100 447.600 ;
        RECT 514.800 434.700 516.600 441.600 ;
        RECT 532.500 434.700 534.300 447.600 ;
        RECT 547.800 434.700 549.600 447.600 ;
        RECT 553.800 434.700 555.600 447.600 ;
        RECT 566.700 434.700 568.500 447.600 ;
        RECT 581.400 434.700 583.200 441.600 ;
        RECT 604.800 434.700 606.600 447.600 ;
        RECT 614.400 434.700 616.200 441.600 ;
        RECT 637.800 434.700 639.600 447.600 ;
        RECT 648.300 434.700 650.100 447.600 ;
        RECT 655.800 434.700 657.600 441.600 ;
        RECT 670.800 434.700 672.600 441.600 ;
        RECT 676.800 434.700 678.600 441.600 ;
        RECT 689.400 434.700 691.200 445.500 ;
        RECT 711.300 434.700 713.100 447.600 ;
        RECT 718.800 434.700 720.600 441.600 ;
        RECT 731.400 434.700 733.200 441.600 ;
        RECT 737.400 434.700 739.200 441.600 ;
        RECT 749.400 434.700 751.200 441.600 ;
        RECT 755.400 434.700 757.200 441.000 ;
        RECT 770.400 434.700 772.200 441.600 ;
        RECT 776.400 434.700 778.200 441.000 ;
        RECT 794.400 434.700 796.200 441.600 ;
        RECT 801.900 434.700 803.700 447.600 ;
        RECT 815.400 434.700 817.200 441.600 ;
        RECT 822.900 434.700 824.700 447.600 ;
        RECT 837.900 434.700 839.700 447.600 ;
        RECT -9.450 432.300 857.400 434.700 ;
        RECT -9.450 362.700 -0.450 432.300 ;
        RECT 11.400 425.400 13.200 432.300 ;
        RECT 18.900 419.400 20.700 432.300 ;
        RECT 34.800 426.000 36.600 432.300 ;
        RECT 40.800 425.400 42.600 432.300 ;
        RECT 58.800 421.200 60.600 432.300 ;
        RECT 74.400 425.400 76.200 432.300 ;
        RECT 81.900 419.400 83.700 432.300 ;
        RECT 97.800 425.400 99.600 432.300 ;
        RECT 110.400 425.400 112.200 432.300 ;
        RECT 117.900 419.400 119.700 432.300 ;
        RECT 129.300 419.400 131.100 432.300 ;
        RECT 136.800 425.400 138.600 432.300 ;
        RECT 151.800 425.400 153.600 432.300 ;
        RECT 157.800 425.400 159.600 432.300 ;
        RECT 167.400 425.400 169.200 432.300 ;
        RECT 173.400 425.400 175.200 432.300 ;
        RECT 185.400 425.400 187.200 432.300 ;
        RECT 191.400 425.400 193.200 432.300 ;
        RECT 208.200 419.400 210.000 432.300 ;
        RECT 214.800 425.400 216.600 432.300 ;
        RECT 227.400 421.500 229.200 432.300 ;
        RECT 251.700 419.400 253.500 432.300 ;
        RECT 269.700 419.400 271.500 432.300 ;
        RECT 286.800 425.400 288.600 432.300 ;
        RECT 292.800 425.400 294.600 432.300 ;
        RECT 305.400 425.400 307.200 432.300 ;
        RECT 312.900 419.400 314.700 432.300 ;
        RECT 323.400 425.400 325.200 432.300 ;
        RECT 329.400 425.400 331.200 432.300 ;
        RECT 346.200 419.400 348.000 432.300 ;
        RECT 352.800 425.400 354.600 432.300 ;
        RECT 362.400 425.400 364.200 432.300 ;
        RECT 368.400 425.400 370.200 432.300 ;
        RECT 383.400 421.200 385.200 432.300 ;
        RECT 406.500 419.400 408.300 432.300 ;
        RECT 420.300 419.400 422.100 432.300 ;
        RECT 427.800 425.400 429.600 432.300 ;
        RECT 441.300 419.400 443.100 432.300 ;
        RECT 448.800 425.400 450.600 432.300 ;
        RECT 466.800 425.400 468.600 432.300 ;
        RECT 473.550 428.400 475.350 432.300 ;
        RECT 482.250 425.400 484.050 432.300 ;
        RECT 488.850 425.400 490.650 432.300 ;
        RECT 499.050 425.400 500.850 432.300 ;
        RECT 513.300 419.400 515.100 432.300 ;
        RECT 520.800 425.400 522.600 432.300 ;
        RECT 533.400 425.400 535.200 432.300 ;
        RECT 539.400 425.400 541.200 432.300 ;
        RECT 559.800 419.400 561.600 432.300 ;
        RECT 574.500 419.400 576.300 432.300 ;
        RECT 589.800 425.400 591.600 432.300 ;
        RECT 595.800 425.400 597.600 432.300 ;
        RECT 606.300 419.400 608.100 432.300 ;
        RECT 613.800 425.400 615.600 432.300 ;
        RECT 637.800 421.500 639.600 432.300 ;
        RECT 651.300 419.400 653.100 432.300 ;
        RECT 658.800 425.400 660.600 432.300 ;
        RECT 673.800 425.400 675.600 432.300 ;
        RECT 679.800 425.400 681.600 432.300 ;
        RECT 690.300 419.400 692.100 432.300 ;
        RECT 697.800 425.400 699.600 432.300 ;
        RECT 713.400 425.400 715.200 432.300 ;
        RECT 720.900 419.400 722.700 432.300 ;
        RECT 734.400 424.200 736.200 432.300 ;
        RECT 743.400 419.400 745.200 432.300 ;
        RECT 755.400 425.400 757.200 432.300 ;
        RECT 761.400 425.400 763.200 432.300 ;
        RECT 778.800 419.400 780.600 432.300 ;
        RECT 793.800 419.400 795.600 432.300 ;
        RECT 805.800 425.400 807.600 432.300 ;
        RECT 811.800 425.400 813.600 432.300 ;
        RECT 821.400 425.400 823.200 432.300 ;
        RECT 827.400 425.400 829.200 432.300 ;
        RECT 839.400 425.400 841.200 432.300 ;
        RECT 846.000 419.400 847.800 432.300 ;
        RECT 13.800 362.700 15.600 369.000 ;
        RECT 19.800 362.700 21.600 369.600 ;
        RECT 32.400 362.700 34.200 373.800 ;
        RECT 55.800 362.700 57.600 369.000 ;
        RECT 61.800 362.700 63.600 369.600 ;
        RECT 82.800 362.700 84.600 373.500 ;
        RECT 103.800 362.700 105.600 373.800 ;
        RECT 121.800 362.700 123.600 369.600 ;
        RECT 133.800 362.700 135.600 369.600 ;
        RECT 139.800 362.700 141.600 369.600 ;
        RECT 154.800 362.700 156.600 369.000 ;
        RECT 160.800 362.700 162.600 369.600 ;
        RECT 170.400 362.700 172.200 375.600 ;
        RECT 190.800 362.700 192.600 369.600 ;
        RECT 196.800 362.700 198.600 369.600 ;
        RECT 211.800 362.700 213.600 369.600 ;
        RECT 226.800 362.700 228.600 369.600 ;
        RECT 241.800 362.700 243.600 369.000 ;
        RECT 247.800 362.700 249.600 369.600 ;
        RECT 268.800 362.700 270.600 373.500 ;
        RECT 286.800 362.700 288.600 369.600 ;
        RECT 301.800 362.700 303.600 369.000 ;
        RECT 307.800 362.700 309.600 369.600 ;
        RECT 318.300 362.700 320.100 375.600 ;
        RECT 325.800 362.700 327.600 369.600 ;
        RECT 343.200 362.700 345.000 375.600 ;
        RECT 349.800 362.700 351.600 369.600 ;
        RECT 364.500 362.700 366.300 375.600 ;
        RECT 377.400 362.700 379.200 369.600 ;
        RECT 384.000 362.700 385.800 375.600 ;
        RECT 403.500 362.700 405.300 375.600 ;
        RECT 416.400 362.700 418.200 369.600 ;
        RECT 434.400 362.700 436.200 373.500 ;
        RECT 452.550 362.700 454.350 366.600 ;
        RECT 461.250 362.700 463.050 369.600 ;
        RECT 467.850 362.700 469.650 369.600 ;
        RECT 478.050 362.700 479.850 369.600 ;
        RECT 492.300 362.700 494.100 375.600 ;
        RECT 499.800 362.700 501.600 369.600 ;
        RECT 515.400 362.700 517.200 373.800 ;
        RECT 536.400 362.700 538.200 369.600 ;
        RECT 543.900 362.700 545.700 375.600 ;
        RECT 557.400 362.700 559.200 369.600 ;
        RECT 564.900 362.700 566.700 375.600 ;
        RECT 577.800 362.700 579.600 375.600 ;
        RECT 586.800 362.700 588.600 370.800 ;
        RECT 599.400 362.700 601.200 369.600 ;
        RECT 605.400 362.700 607.200 369.600 ;
        RECT 618.300 362.700 620.100 375.600 ;
        RECT 625.800 362.700 627.600 369.600 ;
        RECT 641.400 362.700 643.200 373.500 ;
        RECT 667.800 362.700 669.600 369.000 ;
        RECT 673.800 362.700 675.600 369.600 ;
        RECT 686.700 362.700 688.500 375.600 ;
        RECT 703.800 362.700 705.600 369.600 ;
        RECT 709.800 362.700 711.600 369.600 ;
        RECT 719.400 362.700 721.200 369.600 ;
        RECT 739.800 362.700 741.600 369.600 ;
        RECT 755.700 362.700 757.500 375.600 ;
        RECT 770.400 362.700 772.200 369.600 ;
        RECT 776.400 362.700 778.200 369.600 ;
        RECT 791.400 362.700 793.200 369.600 ;
        RECT 798.900 362.700 800.700 375.600 ;
        RECT 812.400 362.700 814.200 373.500 ;
        RECT 833.400 362.700 835.200 369.600 ;
        RECT 839.400 362.700 841.200 369.600 ;
        RECT -9.450 360.300 857.400 362.700 ;
        RECT -9.450 290.700 -0.450 360.300 ;
        RECT 13.800 354.000 15.600 360.300 ;
        RECT 19.800 353.400 21.600 360.300 ;
        RECT 32.400 353.400 34.200 360.300 ;
        RECT 39.900 347.400 41.700 360.300 ;
        RECT 51.300 347.400 53.100 360.300 ;
        RECT 58.800 353.400 60.600 360.300 ;
        RECT 76.800 354.000 78.600 360.300 ;
        RECT 82.800 353.400 84.600 360.300 ;
        RECT 95.400 353.400 97.200 360.300 ;
        RECT 102.900 347.400 104.700 360.300 ;
        RECT 113.400 353.400 115.200 360.300 ;
        RECT 119.400 354.000 121.200 360.300 ;
        RECT 135.300 347.400 137.100 360.300 ;
        RECT 142.800 353.400 144.600 360.300 ;
        RECT 160.800 354.000 162.600 360.300 ;
        RECT 166.800 353.400 168.600 360.300 ;
        RECT 181.800 354.000 183.600 360.300 ;
        RECT 187.800 353.400 189.600 360.300 ;
        RECT 197.400 353.400 199.200 360.300 ;
        RECT 203.400 353.400 205.200 360.300 ;
        RECT 218.400 353.400 220.200 360.300 ;
        RECT 225.900 347.400 227.700 360.300 ;
        RECT 236.400 347.400 238.200 360.300 ;
        RECT 257.400 353.400 259.200 360.300 ;
        RECT 264.900 347.400 266.700 360.300 ;
        RECT 278.400 353.400 280.200 360.300 ;
        RECT 285.900 347.400 287.700 360.300 ;
        RECT 297.300 347.400 299.100 360.300 ;
        RECT 304.800 353.400 306.600 360.300 ;
        RECT 319.800 353.400 321.600 360.300 ;
        RECT 325.800 353.400 327.600 360.300 ;
        RECT 340.200 347.400 342.000 360.300 ;
        RECT 346.800 353.400 348.600 360.300 ;
        RECT 358.800 353.400 360.600 360.300 ;
        RECT 364.800 353.400 366.600 360.300 ;
        RECT 374.400 347.400 376.200 360.300 ;
        RECT 389.400 353.400 391.200 360.300 ;
        RECT 395.400 353.400 397.200 360.300 ;
        RECT 410.700 347.400 412.500 360.300 ;
        RECT 430.800 353.400 432.600 360.300 ;
        RECT 448.800 347.400 450.600 360.300 ;
        RECT 469.800 349.500 471.600 360.300 ;
        RECT 490.800 347.400 492.600 360.300 ;
        RECT 508.800 347.400 510.600 360.300 ;
        RECT 526.800 349.200 528.600 360.300 ;
        RECT 544.800 353.400 546.600 360.300 ;
        RECT 555.300 347.400 557.100 360.300 ;
        RECT 562.800 353.400 564.600 360.300 ;
        RECT 577.800 353.400 579.600 360.300 ;
        RECT 583.800 353.400 585.600 360.300 ;
        RECT 594.300 347.400 596.100 360.300 ;
        RECT 601.800 353.400 603.600 360.300 ;
        RECT 617.400 353.400 619.200 360.300 ;
        RECT 624.900 347.400 626.700 360.300 ;
        RECT 635.400 347.400 637.200 360.300 ;
        RECT 655.800 353.400 657.600 360.300 ;
        RECT 661.800 353.400 663.600 360.300 ;
        RECT 682.800 349.500 684.600 360.300 ;
        RECT 698.400 349.500 700.200 360.300 ;
        RECT 721.800 353.400 723.600 360.300 ;
        RECT 727.800 353.400 729.600 360.300 ;
        RECT 742.200 347.400 744.000 360.300 ;
        RECT 748.800 353.400 750.600 360.300 ;
        RECT 761.400 349.500 763.200 360.300 ;
        RECT 785.400 349.500 787.200 360.300 ;
        RECT 809.400 353.400 811.200 360.300 ;
        RECT 816.900 347.400 818.700 360.300 ;
        RECT 828.300 347.400 830.100 360.300 ;
        RECT 835.800 353.400 837.600 360.300 ;
        RECT 16.800 290.700 18.600 301.800 ;
        RECT 29.400 290.700 31.200 297.600 ;
        RECT 35.400 290.700 37.200 297.000 ;
        RECT 58.800 290.700 60.600 301.800 ;
        RECT 74.400 290.700 76.200 297.600 ;
        RECT 81.900 290.700 83.700 303.600 ;
        RECT 97.200 290.700 99.000 303.600 ;
        RECT 103.800 290.700 105.600 297.600 ;
        RECT 113.400 290.700 115.200 297.600 ;
        RECT 119.400 290.700 121.200 297.600 ;
        RECT 131.400 290.700 133.200 297.600 ;
        RECT 137.400 290.700 139.200 297.600 ;
        RECT 151.800 290.700 153.600 297.600 ;
        RECT 157.800 290.700 159.600 297.600 ;
        RECT 172.800 290.700 174.600 297.000 ;
        RECT 178.800 290.700 180.600 297.600 ;
        RECT 193.800 290.700 195.600 297.000 ;
        RECT 199.800 290.700 201.600 297.600 ;
        RECT 214.800 290.700 216.600 297.600 ;
        RECT 235.800 290.700 237.600 301.500 ;
        RECT 250.800 290.700 252.600 297.600 ;
        RECT 256.800 290.700 258.600 297.600 ;
        RECT 277.800 290.700 279.600 301.500 ;
        RECT 295.800 290.700 297.600 297.000 ;
        RECT 301.800 290.700 303.600 297.600 ;
        RECT 312.300 290.700 314.100 303.600 ;
        RECT 319.800 290.700 321.600 297.600 ;
        RECT 334.800 290.700 336.600 297.600 ;
        RECT 340.800 290.700 342.600 297.600 ;
        RECT 355.800 290.700 357.600 297.000 ;
        RECT 361.800 290.700 363.600 297.600 ;
        RECT 372.300 290.700 374.100 303.600 ;
        RECT 379.800 290.700 381.600 297.600 ;
        RECT 392.400 290.700 394.200 297.600 ;
        RECT 399.000 290.700 400.800 303.600 ;
        RECT 413.400 290.700 415.200 297.600 ;
        RECT 428.400 290.700 430.200 297.600 ;
        RECT 434.400 290.700 436.200 297.600 ;
        RECT 446.400 290.700 448.200 297.600 ;
        RECT 452.400 290.700 454.200 297.600 ;
        RECT 465.300 290.700 467.100 303.600 ;
        RECT 472.800 290.700 474.600 297.600 ;
        RECT 485.400 290.700 487.200 297.600 ;
        RECT 491.400 290.700 493.200 297.600 ;
        RECT 506.400 290.700 508.200 301.800 ;
        RECT 525.300 290.700 527.100 303.600 ;
        RECT 532.800 290.700 534.600 297.600 ;
        RECT 545.400 290.700 547.200 303.600 ;
        RECT 568.800 290.700 570.600 297.000 ;
        RECT 574.800 290.700 576.600 297.600 ;
        RECT 584.400 290.700 586.200 297.600 ;
        RECT 590.400 290.700 592.200 297.600 ;
        RECT 607.800 290.700 609.600 297.000 ;
        RECT 613.800 290.700 615.600 297.600 ;
        RECT 626.400 290.700 628.200 297.600 ;
        RECT 633.900 290.700 635.700 303.600 ;
        RECT 647.400 290.700 649.200 297.600 ;
        RECT 654.900 290.700 656.700 303.600 ;
        RECT 670.200 290.700 672.000 303.600 ;
        RECT 676.800 290.700 678.600 297.600 ;
        RECT 687.300 290.700 689.100 303.600 ;
        RECT 694.800 290.700 696.600 297.600 ;
        RECT 707.400 290.700 709.200 297.600 ;
        RECT 713.400 290.700 715.200 297.600 ;
        RECT 727.800 290.700 729.600 297.600 ;
        RECT 733.800 290.700 735.600 297.600 ;
        RECT 746.400 290.700 748.200 297.600 ;
        RECT 753.900 290.700 755.700 303.600 ;
        RECT 765.300 290.700 767.100 303.600 ;
        RECT 772.800 290.700 774.600 297.600 ;
        RECT 786.300 290.700 788.100 303.600 ;
        RECT 793.800 290.700 795.600 297.600 ;
        RECT 811.200 290.700 813.000 303.600 ;
        RECT 817.800 290.700 819.600 297.600 ;
        RECT 827.400 290.700 829.200 297.600 ;
        RECT 834.000 290.700 835.800 303.600 ;
        RECT -9.450 288.300 857.400 290.700 ;
        RECT -9.450 218.700 -0.450 288.300 ;
        RECT 16.800 277.200 18.600 288.300 ;
        RECT 29.400 281.400 31.200 288.300 ;
        RECT 35.400 282.000 37.200 288.300 ;
        RECT 51.300 275.400 53.100 288.300 ;
        RECT 58.800 281.400 60.600 288.300 ;
        RECT 72.300 275.400 74.100 288.300 ;
        RECT 79.800 281.400 81.600 288.300 ;
        RECT 92.400 281.400 94.200 288.300 ;
        RECT 98.400 282.000 100.200 288.300 ;
        RECT 113.400 281.400 115.200 288.300 ;
        RECT 119.400 282.000 121.200 288.300 ;
        RECT 134.400 281.400 136.200 288.300 ;
        RECT 140.400 282.000 142.200 288.300 ;
        RECT 158.400 277.200 160.200 288.300 ;
        RECT 177.300 275.400 179.100 288.300 ;
        RECT 184.800 281.400 186.600 288.300 ;
        RECT 205.800 277.200 207.600 288.300 ;
        RECT 223.800 281.400 225.600 288.300 ;
        RECT 238.200 275.400 240.000 288.300 ;
        RECT 244.800 281.400 246.600 288.300 ;
        RECT 254.400 281.400 256.200 288.300 ;
        RECT 260.400 281.400 262.200 288.300 ;
        RECT 279.300 275.400 281.100 288.300 ;
        RECT 293.400 281.400 295.200 288.300 ;
        RECT 299.400 281.400 301.200 288.300 ;
        RECT 314.400 281.400 316.200 288.300 ;
        RECT 321.900 275.400 323.700 288.300 ;
        RECT 340.800 275.400 342.600 288.300 ;
        RECT 351.300 275.400 353.100 288.300 ;
        RECT 358.800 281.400 360.600 288.300 ;
        RECT 371.400 275.400 373.200 288.300 ;
        RECT 389.400 281.400 391.200 288.300 ;
        RECT 395.400 281.400 397.200 288.300 ;
        RECT 412.800 281.400 414.600 288.300 ;
        RECT 424.800 281.400 426.600 288.300 ;
        RECT 430.800 281.400 432.600 288.300 ;
        RECT 448.800 277.200 450.600 288.300 ;
        RECT 472.800 277.500 474.600 288.300 ;
        RECT 485.400 281.400 487.200 288.300 ;
        RECT 491.400 281.400 493.200 288.300 ;
        RECT 503.400 275.400 505.200 288.300 ;
        RECT 521.400 275.400 523.200 288.300 ;
        RECT 542.400 281.400 544.200 288.300 ;
        RECT 549.900 275.400 551.700 288.300 ;
        RECT 571.800 277.500 573.600 288.300 ;
        RECT 587.400 277.200 589.200 288.300 ;
        RECT 608.400 281.400 610.200 288.300 ;
        RECT 615.900 275.400 617.700 288.300 ;
        RECT 629.400 281.400 631.200 288.300 ;
        RECT 636.900 275.400 638.700 288.300 ;
        RECT 647.400 281.400 649.200 288.300 ;
        RECT 662.400 281.400 664.200 288.300 ;
        RECT 680.400 281.400 682.200 288.300 ;
        RECT 687.900 275.400 689.700 288.300 ;
        RECT 701.400 277.200 703.200 288.300 ;
        RECT 722.700 275.400 724.500 288.300 ;
        RECT 738.300 275.400 740.100 288.300 ;
        RECT 745.800 281.400 747.600 288.300 ;
        RECT 761.400 277.200 763.200 288.300 ;
        RECT 782.700 275.400 784.500 288.300 ;
        RECT 805.800 275.400 807.600 288.300 ;
        RECT 820.500 275.400 822.300 288.300 ;
        RECT 836.400 281.400 838.200 288.300 ;
        RECT 843.900 275.400 845.700 288.300 ;
        RECT 11.400 218.700 13.200 225.600 ;
        RECT 18.900 218.700 20.700 231.600 ;
        RECT 37.800 218.700 39.600 229.800 ;
        RECT 58.800 218.700 60.600 229.800 ;
        RECT 71.400 218.700 73.200 225.600 ;
        RECT 77.400 218.700 79.200 225.000 ;
        RECT 97.800 218.700 99.600 225.000 ;
        RECT 103.800 218.700 105.600 225.600 ;
        RECT 121.800 218.700 123.600 229.800 ;
        RECT 135.300 218.700 137.100 231.600 ;
        RECT 142.800 218.700 144.600 225.600 ;
        RECT 158.400 218.700 160.200 229.800 ;
        RECT 176.400 218.700 178.200 225.600 ;
        RECT 182.400 218.700 184.200 225.000 ;
        RECT 198.300 218.700 200.100 231.600 ;
        RECT 205.800 218.700 207.600 225.600 ;
        RECT 219.300 218.700 221.100 231.600 ;
        RECT 226.800 218.700 228.600 225.600 ;
        RECT 239.400 218.700 241.200 225.600 ;
        RECT 245.400 218.700 247.200 225.000 ;
        RECT 263.400 218.700 265.200 229.800 ;
        RECT 281.400 218.700 283.200 225.600 ;
        RECT 287.400 218.700 289.200 225.000 ;
        RECT 305.400 218.700 307.200 229.800 ;
        RECT 323.400 218.700 325.200 225.600 ;
        RECT 329.400 218.700 331.200 225.000 ;
        RECT 352.800 218.700 354.600 229.800 ;
        RECT 365.400 218.700 367.200 225.600 ;
        RECT 371.400 218.700 373.200 225.000 ;
        RECT 391.800 218.700 393.600 225.600 ;
        RECT 404.400 218.700 406.200 225.600 ;
        RECT 411.900 218.700 413.700 231.600 ;
        RECT 423.300 218.700 425.100 231.600 ;
        RECT 430.800 218.700 432.600 225.600 ;
        RECT 443.400 218.700 445.200 225.600 ;
        RECT 449.400 218.700 451.200 225.600 ;
        RECT 463.800 218.700 465.600 225.600 ;
        RECT 469.800 218.700 471.600 225.600 ;
        RECT 479.400 218.700 481.200 225.600 ;
        RECT 486.000 218.700 487.800 231.600 ;
        RECT 501.300 218.700 503.100 231.600 ;
        RECT 508.800 218.700 510.600 225.600 ;
        RECT 522.300 218.700 524.100 231.600 ;
        RECT 529.800 218.700 531.600 225.600 ;
        RECT 542.400 218.700 544.200 225.600 ;
        RECT 548.400 218.700 550.200 225.600 ;
        RECT 565.800 218.700 567.600 225.600 ;
        RECT 580.800 218.700 582.600 225.600 ;
        RECT 587.550 218.700 589.350 222.600 ;
        RECT 596.250 218.700 598.050 225.600 ;
        RECT 602.850 218.700 604.650 225.600 ;
        RECT 613.050 218.700 614.850 225.600 ;
        RECT 626.400 218.700 628.200 225.600 ;
        RECT 641.400 218.700 643.200 225.600 ;
        RECT 647.400 218.700 649.200 225.600 ;
        RECT 661.800 218.700 663.600 225.600 ;
        RECT 667.800 218.700 669.600 225.600 ;
        RECT 680.400 218.700 682.200 226.800 ;
        RECT 689.400 218.700 691.200 231.600 ;
        RECT 704.400 218.700 706.200 225.600 ;
        RECT 711.900 218.700 713.700 231.600 ;
        RECT 723.300 218.700 725.100 231.600 ;
        RECT 730.800 218.700 732.600 225.600 ;
        RECT 744.300 218.700 746.100 231.600 ;
        RECT 751.800 218.700 753.600 225.600 ;
        RECT 765.300 218.700 767.100 231.600 ;
        RECT 772.800 218.700 774.600 225.600 ;
        RECT 788.400 218.700 790.200 229.800 ;
        RECT 814.800 218.700 816.600 229.800 ;
        RECT 828.300 218.700 830.100 231.600 ;
        RECT 835.800 218.700 837.600 225.600 ;
        RECT -9.450 216.300 857.400 218.700 ;
        RECT -9.450 146.700 -0.450 216.300 ;
        RECT 11.400 209.400 13.200 216.300 ;
        RECT 18.900 203.400 20.700 216.300 ;
        RECT 29.400 209.400 31.200 216.300 ;
        RECT 35.400 210.000 37.200 216.300 ;
        RECT 50.400 209.400 52.200 216.300 ;
        RECT 56.400 210.000 58.200 216.300 ;
        RECT 79.800 205.200 81.600 216.300 ;
        RECT 95.400 209.400 97.200 216.300 ;
        RECT 102.900 203.400 104.700 216.300 ;
        RECT 116.400 209.400 118.200 216.300 ;
        RECT 123.900 203.400 125.700 216.300 ;
        RECT 134.400 209.400 136.200 216.300 ;
        RECT 140.400 210.000 142.200 216.300 ;
        RECT 160.200 203.400 162.000 216.300 ;
        RECT 166.800 209.400 168.600 216.300 ;
        RECT 176.400 209.400 178.200 216.300 ;
        RECT 182.400 209.400 184.200 216.300 ;
        RECT 196.800 209.400 198.600 216.300 ;
        RECT 202.800 209.400 204.600 216.300 ;
        RECT 212.400 209.400 214.200 216.300 ;
        RECT 218.400 209.400 220.200 216.300 ;
        RECT 232.800 209.400 234.600 216.300 ;
        RECT 238.800 209.400 240.600 216.300 ;
        RECT 251.400 206.400 253.200 216.300 ;
        RECT 281.400 209.400 283.200 216.300 ;
        RECT 297.300 203.400 299.100 216.300 ;
        RECT 304.800 209.400 306.600 216.300 ;
        RECT 322.800 209.400 324.600 216.300 ;
        RECT 335.400 205.200 337.200 216.300 ;
        RECT 355.800 209.400 357.600 216.300 ;
        RECT 361.800 209.400 363.600 216.300 ;
        RECT 373.800 209.400 375.600 216.300 ;
        RECT 379.800 209.400 381.600 216.300 ;
        RECT 397.800 203.400 399.600 216.300 ;
        RECT 407.400 203.400 409.200 216.300 ;
        RECT 417.900 203.400 419.700 216.300 ;
        RECT 436.800 203.400 438.600 216.300 ;
        RECT 446.400 203.400 448.200 216.300 ;
        RECT 475.800 205.500 477.600 216.300 ;
        RECT 493.800 209.400 495.600 216.300 ;
        RECT 500.550 212.400 502.350 216.300 ;
        RECT 509.250 209.400 511.050 216.300 ;
        RECT 515.850 209.400 517.650 216.300 ;
        RECT 526.050 209.400 527.850 216.300 ;
        RECT 544.800 209.400 546.600 216.300 ;
        RECT 562.800 205.200 564.600 216.300 ;
        RECT 578.400 209.400 580.200 216.300 ;
        RECT 585.900 203.400 587.700 216.300 ;
        RECT 604.800 203.400 606.600 216.300 ;
        RECT 619.200 203.400 621.000 216.300 ;
        RECT 625.800 209.400 627.600 216.300 ;
        RECT 640.800 210.000 642.600 216.300 ;
        RECT 646.800 209.400 648.600 216.300 ;
        RECT 656.400 209.400 658.200 216.300 ;
        RECT 662.400 209.400 664.200 216.300 ;
        RECT 674.400 203.400 676.200 216.300 ;
        RECT 693.300 203.400 695.100 216.300 ;
        RECT 700.800 209.400 702.600 216.300 ;
        RECT 714.300 203.400 716.100 216.300 ;
        RECT 721.800 209.400 723.600 216.300 ;
        RECT 734.400 209.400 736.200 216.300 ;
        RECT 749.400 203.400 751.200 216.300 ;
        RECT 759.900 203.400 761.700 216.300 ;
        RECT 781.800 203.400 783.600 216.300 ;
        RECT 793.800 209.400 795.600 216.300 ;
        RECT 799.800 209.400 801.600 216.300 ;
        RECT 817.800 205.200 819.600 216.300 ;
        RECT 830.400 209.400 832.200 216.300 ;
        RECT 836.400 209.400 838.200 216.300 ;
        RECT 853.800 209.400 855.600 216.300 ;
        RECT 11.400 146.700 13.200 153.600 ;
        RECT 18.900 146.700 20.700 159.600 ;
        RECT 34.800 146.700 36.600 153.000 ;
        RECT 40.800 146.700 42.600 153.600 ;
        RECT 53.400 146.700 55.200 157.800 ;
        RECT 74.400 146.700 76.200 157.800 ;
        RECT 92.400 146.700 94.200 153.600 ;
        RECT 98.400 146.700 100.200 153.000 ;
        RECT 114.300 146.700 116.100 159.600 ;
        RECT 121.800 146.700 123.600 153.600 ;
        RECT 134.400 146.700 136.200 153.600 ;
        RECT 140.400 146.700 142.200 153.000 ;
        RECT 166.800 146.700 168.600 157.500 ;
        RECT 179.400 146.700 181.200 153.600 ;
        RECT 185.400 146.700 187.200 153.000 ;
        RECT 203.400 146.700 205.200 157.800 ;
        RECT 221.400 146.700 223.200 153.600 ;
        RECT 227.400 146.700 229.200 153.600 ;
        RECT 239.400 146.700 241.200 153.600 ;
        RECT 245.400 146.700 247.200 153.000 ;
        RECT 261.300 146.700 263.100 159.600 ;
        RECT 268.800 146.700 270.600 153.600 ;
        RECT 281.400 146.700 283.200 153.600 ;
        RECT 296.400 146.700 298.200 153.600 ;
        RECT 302.400 146.700 304.200 153.000 ;
        RECT 320.400 146.700 322.200 157.800 ;
        RECT 339.300 146.700 341.100 159.600 ;
        RECT 346.800 146.700 348.600 153.600 ;
        RECT 360.300 146.700 362.100 159.600 ;
        RECT 367.800 146.700 369.600 153.600 ;
        RECT 380.400 146.700 382.200 153.600 ;
        RECT 386.400 146.700 388.200 153.000 ;
        RECT 401.400 146.700 403.200 153.600 ;
        RECT 407.400 146.700 409.200 153.600 ;
        RECT 419.400 146.700 421.200 159.600 ;
        RECT 437.400 146.700 439.200 153.600 ;
        RECT 455.400 146.700 457.200 153.600 ;
        RECT 462.900 146.700 464.700 159.600 ;
        RECT 476.400 146.700 478.200 157.800 ;
        RECT 495.300 146.700 497.100 159.600 ;
        RECT 502.800 146.700 504.600 153.600 ;
        RECT 526.800 146.700 528.600 157.500 ;
        RECT 544.800 146.700 546.600 153.600 ;
        RECT 551.550 146.700 553.350 150.600 ;
        RECT 560.250 146.700 562.050 153.600 ;
        RECT 566.850 146.700 568.650 153.600 ;
        RECT 577.050 146.700 578.850 153.600 ;
        RECT 598.800 146.700 600.600 159.600 ;
        RECT 612.900 146.700 614.700 159.600 ;
        RECT 634.800 146.700 636.600 153.000 ;
        RECT 640.800 146.700 642.600 153.600 ;
        RECT 650.400 146.700 652.200 153.600 ;
        RECT 656.400 146.700 658.200 153.600 ;
        RECT 668.400 146.700 670.200 153.600 ;
        RECT 684.300 146.700 686.100 159.600 ;
        RECT 691.800 146.700 693.600 153.600 ;
        RECT 709.800 146.700 711.600 153.600 ;
        RECT 719.400 146.700 721.200 153.600 ;
        RECT 737.400 146.700 739.200 157.800 ;
        RECT 755.400 146.700 757.200 153.600 ;
        RECT 771.300 146.700 773.100 159.600 ;
        RECT 778.800 146.700 780.600 153.600 ;
        RECT 792.300 146.700 794.100 159.600 ;
        RECT 799.800 146.700 801.600 153.600 ;
        RECT 812.400 146.700 814.200 159.600 ;
        RECT 831.300 146.700 833.100 159.600 ;
        RECT 838.800 146.700 840.600 153.600 ;
        RECT -9.450 144.300 857.400 146.700 ;
        RECT -9.450 74.700 -0.450 144.300 ;
        RECT 13.800 137.400 15.600 144.300 ;
        RECT 26.400 133.200 28.200 144.300 ;
        RECT 44.400 137.400 46.200 144.300 ;
        RECT 50.400 138.000 52.200 144.300 ;
        RECT 65.400 137.400 67.200 144.300 ;
        RECT 71.400 138.000 73.200 144.300 ;
        RECT 89.400 137.400 91.200 144.300 ;
        RECT 96.900 131.400 98.700 144.300 ;
        RECT 107.400 137.400 109.200 144.300 ;
        RECT 113.400 138.000 115.200 144.300 ;
        RECT 131.400 133.200 133.200 144.300 ;
        RECT 152.400 137.400 154.200 144.300 ;
        RECT 159.900 131.400 161.700 144.300 ;
        RECT 178.800 131.400 180.600 144.300 ;
        RECT 191.400 137.400 193.200 144.300 ;
        RECT 198.900 131.400 200.700 144.300 ;
        RECT 214.800 137.400 216.600 144.300 ;
        RECT 231.300 131.400 233.100 144.300 ;
        RECT 245.400 131.400 247.200 144.300 ;
        RECT 271.800 131.400 273.600 144.300 ;
        RECT 285.900 131.400 287.700 144.300 ;
        RECT 310.800 133.200 312.600 144.300 ;
        RECT 323.400 137.400 325.200 144.300 ;
        RECT 329.400 138.000 331.200 144.300 ;
        RECT 344.400 137.400 346.200 144.300 ;
        RECT 351.000 131.400 352.800 144.300 ;
        RECT 370.800 137.400 372.600 144.300 ;
        RECT 381.300 131.400 383.100 144.300 ;
        RECT 388.800 137.400 390.600 144.300 ;
        RECT 402.300 131.400 404.100 144.300 ;
        RECT 409.800 137.400 411.600 144.300 ;
        RECT 424.800 137.400 426.600 144.300 ;
        RECT 430.800 137.400 432.600 144.300 ;
        RECT 443.400 133.200 445.200 144.300 ;
        RECT 461.400 137.400 463.200 144.300 ;
        RECT 467.400 138.000 469.200 144.300 ;
        RECT 484.800 131.400 486.600 144.300 ;
        RECT 490.800 131.400 492.600 144.300 ;
        RECT 503.400 133.200 505.200 144.300 ;
        RECT 529.800 133.200 531.600 144.300 ;
        RECT 547.800 137.400 549.600 144.300 ;
        RECT 557.400 137.400 559.200 144.300 ;
        RECT 563.400 137.400 565.200 144.300 ;
        RECT 576.300 131.400 578.100 144.300 ;
        RECT 583.800 137.400 585.600 144.300 ;
        RECT 598.800 137.400 600.600 144.300 ;
        RECT 604.800 137.400 606.600 144.300 ;
        RECT 616.800 137.400 618.600 144.300 ;
        RECT 622.800 137.400 624.600 144.300 ;
        RECT 635.400 133.200 637.200 144.300 ;
        RECT 658.800 137.400 660.600 144.300 ;
        RECT 671.400 137.400 673.200 144.300 ;
        RECT 678.900 131.400 680.700 144.300 ;
        RECT 694.200 131.400 696.000 144.300 ;
        RECT 700.800 137.400 702.600 144.300 ;
        RECT 715.800 138.000 717.600 144.300 ;
        RECT 721.800 137.400 723.600 144.300 ;
        RECT 736.800 137.400 738.600 144.300 ;
        RECT 751.800 137.400 753.600 144.300 ;
        RECT 764.400 137.400 766.200 144.300 ;
        RECT 771.900 131.400 773.700 144.300 ;
        RECT 784.800 137.400 786.600 144.300 ;
        RECT 790.800 137.400 792.600 144.300 ;
        RECT 803.400 137.400 805.200 144.300 ;
        RECT 810.900 131.400 812.700 144.300 ;
        RECT 824.400 137.400 826.200 144.300 ;
        RECT 831.900 131.400 833.700 144.300 ;
        RECT 843.300 131.400 845.100 144.300 ;
        RECT 850.800 137.400 852.600 144.300 ;
        RECT 13.800 74.700 15.600 81.600 ;
        RECT 26.400 74.700 28.200 81.600 ;
        RECT 33.900 74.700 35.700 87.600 ;
        RECT 49.800 74.700 51.600 81.000 ;
        RECT 55.800 74.700 57.600 81.600 ;
        RECT 68.400 74.700 70.200 85.800 ;
        RECT 94.800 74.700 96.600 85.800 ;
        RECT 112.800 74.700 114.600 81.000 ;
        RECT 118.800 74.700 120.600 81.600 ;
        RECT 133.800 74.700 135.600 81.000 ;
        RECT 139.800 74.700 141.600 81.600 ;
        RECT 152.400 74.700 154.200 81.600 ;
        RECT 159.900 74.700 161.700 87.600 ;
        RECT 171.300 74.700 173.100 87.600 ;
        RECT 178.800 74.700 180.600 81.600 ;
        RECT 194.400 74.700 196.200 81.600 ;
        RECT 201.900 74.700 203.700 87.600 ;
        RECT 217.800 74.700 219.600 81.000 ;
        RECT 223.800 74.700 225.600 81.600 ;
        RECT 241.800 74.700 243.600 85.800 ;
        RECT 257.400 74.700 259.200 81.600 ;
        RECT 264.900 74.700 266.700 87.600 ;
        RECT 275.400 74.700 277.200 81.600 ;
        RECT 290.400 74.700 292.200 81.600 ;
        RECT 296.400 74.700 298.200 81.000 ;
        RECT 316.800 74.700 318.600 81.000 ;
        RECT 322.800 74.700 324.600 81.600 ;
        RECT 335.400 74.700 337.200 85.800 ;
        RECT 356.400 74.700 358.200 81.600 ;
        RECT 363.900 74.700 365.700 87.600 ;
        RECT 374.400 74.700 376.200 81.600 ;
        RECT 392.400 74.700 394.200 81.600 ;
        RECT 399.900 74.700 401.700 87.600 ;
        RECT 411.300 74.700 413.100 87.600 ;
        RECT 418.800 74.700 420.600 81.600 ;
        RECT 436.800 74.700 438.600 81.000 ;
        RECT 442.800 74.700 444.600 81.600 ;
        RECT 455.400 74.700 457.200 85.800 ;
        RECT 475.800 74.700 477.600 81.600 ;
        RECT 481.800 74.700 483.600 81.600 ;
        RECT 491.400 74.700 493.200 81.600 ;
        RECT 508.800 74.700 510.600 81.600 ;
        RECT 514.800 74.700 516.600 81.600 ;
        RECT 532.800 74.700 534.600 85.800 ;
        RECT 546.300 74.700 548.100 87.600 ;
        RECT 553.800 74.700 555.600 81.600 ;
        RECT 568.800 74.700 570.600 81.600 ;
        RECT 574.800 74.700 576.600 81.600 ;
        RECT 589.200 74.700 591.000 87.600 ;
        RECT 595.800 74.700 597.600 81.600 ;
        RECT 605.400 74.700 607.200 87.600 ;
        RECT 631.800 74.700 633.600 87.600 ;
        RECT 641.400 74.700 643.200 87.600 ;
        RECT 659.400 74.700 661.200 87.600 ;
        RECT 680.400 74.700 682.200 85.800 ;
        RECT 699.300 74.700 701.100 87.600 ;
        RECT 706.800 74.700 708.600 81.600 ;
        RECT 719.400 74.700 721.200 81.600 ;
        RECT 725.400 74.700 727.200 81.600 ;
        RECT 742.800 74.700 744.600 81.600 ;
        RECT 753.300 74.700 755.100 87.600 ;
        RECT 760.800 74.700 762.600 81.600 ;
        RECT 778.800 74.700 780.600 81.000 ;
        RECT 784.800 74.700 786.600 81.600 ;
        RECT 797.400 74.700 799.200 85.800 ;
        RECT 815.400 74.700 817.200 81.600 ;
        RECT 830.400 74.700 832.200 81.600 ;
        RECT 836.400 74.700 838.200 81.600 ;
        RECT 853.800 74.700 855.600 81.600 ;
        RECT -9.450 72.300 857.400 74.700 ;
        RECT -9.450 2.700 -0.450 72.300 ;
        RECT 13.800 66.000 15.600 72.300 ;
        RECT 19.800 65.400 21.600 72.300 ;
        RECT 32.400 61.200 34.200 72.300 ;
        RECT 51.300 59.400 53.100 72.300 ;
        RECT 58.800 65.400 60.600 72.300 ;
        RECT 76.800 66.000 78.600 72.300 ;
        RECT 82.800 65.400 84.600 72.300 ;
        RECT 103.800 61.500 105.600 72.300 ;
        RECT 119.400 65.400 121.200 72.300 ;
        RECT 126.900 59.400 128.700 72.300 ;
        RECT 142.800 66.000 144.600 72.300 ;
        RECT 148.800 65.400 150.600 72.300 ;
        RECT 161.400 61.200 163.200 72.300 ;
        RECT 182.400 65.400 184.200 72.300 ;
        RECT 189.900 59.400 191.700 72.300 ;
        RECT 205.800 66.000 207.600 72.300 ;
        RECT 211.800 65.400 213.600 72.300 ;
        RECT 229.800 61.200 231.600 72.300 ;
        RECT 247.200 59.400 249.000 72.300 ;
        RECT 253.800 65.400 255.600 72.300 ;
        RECT 263.400 65.400 265.200 72.300 ;
        RECT 269.400 65.400 271.200 72.300 ;
        RECT 284.400 61.200 286.200 72.300 ;
        RECT 302.400 65.400 304.200 72.300 ;
        RECT 308.400 66.000 310.200 72.300 ;
        RECT 323.400 65.400 325.200 72.300 ;
        RECT 329.400 65.400 331.200 72.300 ;
        RECT 346.800 65.400 348.600 72.300 ;
        RECT 356.400 65.400 358.200 72.300 ;
        RECT 362.400 66.000 364.200 72.300 ;
        RECT 382.800 66.000 384.600 72.300 ;
        RECT 388.800 65.400 390.600 72.300 ;
        RECT 398.400 65.400 400.200 72.300 ;
        RECT 404.400 65.400 406.200 72.300 ;
        RECT 419.400 61.200 421.200 72.300 ;
        RECT 440.400 61.500 442.200 72.300 ;
        RECT 458.550 68.400 460.350 72.300 ;
        RECT 467.250 65.400 469.050 72.300 ;
        RECT 473.850 65.400 475.650 72.300 ;
        RECT 484.050 65.400 485.850 72.300 ;
        RECT 497.400 65.400 499.200 72.300 ;
        RECT 515.400 61.500 517.200 72.300 ;
        RECT 539.700 59.400 541.500 72.300 ;
        RECT 559.500 59.400 561.300 72.300 ;
        RECT 577.800 66.000 579.600 72.300 ;
        RECT 583.800 65.400 585.600 72.300 ;
        RECT 596.400 65.400 598.200 72.300 ;
        RECT 603.900 59.400 605.700 72.300 ;
        RECT 614.400 65.400 616.200 72.300 ;
        RECT 634.800 66.000 636.600 72.300 ;
        RECT 640.800 65.400 642.600 72.300 ;
        RECT 650.400 65.400 652.200 72.300 ;
        RECT 656.400 65.400 658.200 72.300 ;
        RECT 670.800 65.400 672.600 72.300 ;
        RECT 676.800 65.400 678.600 72.300 ;
        RECT 688.800 65.400 690.600 72.300 ;
        RECT 694.800 65.400 696.600 72.300 ;
        RECT 709.800 66.000 711.600 72.300 ;
        RECT 715.800 65.400 717.600 72.300 ;
        RECT 728.400 61.200 730.200 72.300 ;
        RECT 748.800 65.400 750.600 72.300 ;
        RECT 754.800 65.400 756.600 72.300 ;
        RECT 769.800 66.000 771.600 72.300 ;
        RECT 775.800 65.400 777.600 72.300 ;
        RECT 790.800 66.000 792.600 72.300 ;
        RECT 796.800 65.400 798.600 72.300 ;
        RECT 809.400 65.400 811.200 72.300 ;
        RECT 816.900 59.400 818.700 72.300 ;
        RECT 830.400 65.400 832.200 72.300 ;
        RECT 837.900 59.400 839.700 72.300 ;
        RECT 853.800 65.400 855.600 72.300 ;
        RECT 13.800 2.700 15.600 9.600 ;
        RECT 23.400 2.700 25.200 9.600 ;
        RECT 29.400 2.700 31.200 9.000 ;
        RECT 47.400 2.700 49.200 9.600 ;
        RECT 54.900 2.700 56.700 15.600 ;
        RECT 66.300 2.700 68.100 15.600 ;
        RECT 73.800 2.700 75.600 9.600 ;
        RECT 86.400 2.700 88.200 9.600 ;
        RECT 92.400 2.700 94.200 9.000 ;
        RECT 107.400 2.700 109.200 9.600 ;
        RECT 113.400 2.700 115.200 9.000 ;
        RECT 128.400 2.700 130.200 9.600 ;
        RECT 134.400 2.700 136.200 9.000 ;
        RECT 149.400 2.700 151.200 9.600 ;
        RECT 169.800 2.700 171.600 9.000 ;
        RECT 175.800 2.700 177.600 9.600 ;
        RECT 188.400 2.700 190.200 13.800 ;
        RECT 209.400 2.700 211.200 12.600 ;
        RECT 240.300 2.700 242.100 15.600 ;
        RECT 247.800 2.700 249.600 9.600 ;
        RECT 260.400 2.700 262.200 9.600 ;
        RECT 278.400 2.700 280.200 9.600 ;
        RECT 285.900 2.700 287.700 15.600 ;
        RECT 296.400 2.700 298.200 9.600 ;
        RECT 312.300 2.700 314.100 15.600 ;
        RECT 319.800 2.700 321.600 9.600 ;
        RECT 332.400 2.700 334.200 9.600 ;
        RECT 338.400 2.700 340.200 9.600 ;
        RECT 353.400 2.700 355.200 9.600 ;
        RECT 360.900 2.700 362.700 15.600 ;
        RECT 373.800 2.700 375.600 9.600 ;
        RECT 379.800 2.700 381.600 9.600 ;
        RECT 394.800 2.700 396.600 9.600 ;
        RECT 407.700 2.700 409.500 15.600 ;
        RECT 427.800 2.700 429.600 9.600 ;
        RECT 435.150 2.700 436.950 9.600 ;
        RECT 445.350 2.700 447.150 9.600 ;
        RECT 451.950 2.700 453.750 9.600 ;
        RECT 460.650 2.700 462.450 6.600 ;
        RECT 478.500 2.700 480.300 15.600 ;
        RECT 496.500 2.700 498.300 15.600 ;
        RECT 514.800 2.700 516.600 9.600 ;
        RECT 526.800 2.700 528.600 9.600 ;
        RECT 532.800 2.700 534.600 9.600 ;
        RECT 544.800 2.700 546.600 9.600 ;
        RECT 550.800 2.700 552.600 9.600 ;
        RECT 565.800 2.700 567.600 9.000 ;
        RECT 571.800 2.700 573.600 9.600 ;
        RECT 584.400 2.700 586.200 9.600 ;
        RECT 591.900 2.700 593.700 15.600 ;
        RECT 607.500 2.700 609.300 15.600 ;
        RECT 625.200 2.700 627.000 15.600 ;
        RECT 631.800 2.700 633.600 9.600 ;
        RECT 641.400 2.700 643.200 9.600 ;
        RECT 647.400 2.700 649.200 9.600 ;
        RECT 659.400 2.700 661.200 9.600 ;
        RECT 665.400 2.700 667.200 9.600 ;
        RECT 682.800 2.700 684.600 9.000 ;
        RECT 688.800 2.700 690.600 9.600 ;
        RECT 703.800 2.700 705.600 9.600 ;
        RECT 718.800 2.700 720.600 9.000 ;
        RECT 724.800 2.700 726.600 9.600 ;
        RECT 734.400 2.700 736.200 9.600 ;
        RECT 740.400 2.700 742.200 9.600 ;
        RECT 749.550 2.700 751.350 6.600 ;
        RECT 758.250 2.700 760.050 9.600 ;
        RECT 764.850 2.700 766.650 9.600 ;
        RECT 775.050 2.700 776.850 9.600 ;
        RECT 791.400 2.700 793.200 13.800 ;
        RECT 810.300 2.700 812.100 15.600 ;
        RECT 817.800 2.700 819.600 9.600 ;
        RECT 833.700 2.700 835.500 15.600 ;
        RECT 848.400 2.700 850.200 9.600 ;
        RECT -9.450 0.300 857.400 2.700 ;
      LAYER metal2 ;
        RECT 709.950 856.950 714.450 859.050 ;
        RECT 625.950 849.450 628.050 850.050 ;
        RECT 630.000 849.450 634.050 850.050 ;
        RECT 625.950 848.400 634.050 849.450 ;
        RECT 625.950 847.950 628.050 848.400 ;
        RECT 630.000 847.950 634.050 848.400 ;
        RECT 709.950 844.950 712.050 847.050 ;
        RECT 767.550 784.950 772.050 787.050 ;
        RECT 769.950 772.950 772.050 775.050 ;
      LAYER metal3 ;
        RECT 709.950 856.950 712.050 859.050 ;
        RECT 710.400 847.050 711.600 856.950 ;
        RECT 709.950 844.950 712.050 847.050 ;
        RECT 769.950 784.950 772.050 787.050 ;
        RECT 770.400 775.050 771.600 784.950 ;
        RECT 769.950 772.950 772.050 775.050 ;
    END
  END vdd
  PIN ABCmd_i[7]
    PORT
      LAYER metal1 ;
        RECT 565.950 523.950 568.050 526.050 ;
        RECT 529.950 484.950 532.050 487.050 ;
        RECT 415.950 451.950 418.050 454.050 ;
        RECT 436.950 448.950 439.050 454.050 ;
        RECT 472.950 451.950 475.200 454.050 ;
        RECT 478.950 451.950 481.050 454.050 ;
        RECT 479.550 442.050 480.450 451.950 ;
        RECT 478.950 439.950 481.050 442.050 ;
        RECT 562.950 379.950 565.050 382.050 ;
        RECT 544.950 310.950 547.050 313.050 ;
        RECT 502.950 265.950 505.050 268.050 ;
        RECT 517.950 265.950 523.050 268.050 ;
        RECT 508.950 235.950 511.050 238.050 ;
        RECT 607.950 169.950 610.050 172.050 ;
        RECT 502.950 163.950 505.050 166.050 ;
        RECT 388.800 124.950 391.050 127.050 ;
        RECT 490.950 124.950 493.200 127.050 ;
      LAYER metal2 ;
        RECT 646.950 864.450 649.050 865.050 ;
        RECT 646.950 863.400 744.450 864.450 ;
        RECT 646.950 862.950 649.050 863.400 ;
        RECT 743.400 861.450 744.450 863.400 ;
        RECT 757.950 861.450 760.050 862.200 ;
        RECT 743.400 860.400 760.050 861.450 ;
        RECT 757.950 860.100 760.050 860.400 ;
        RECT 628.950 687.450 631.050 688.050 ;
        RECT 643.950 687.450 646.050 688.050 ;
        RECT 628.950 686.400 646.050 687.450 ;
        RECT 628.950 685.950 631.050 686.400 ;
        RECT 643.950 685.950 646.050 686.400 ;
        RECT 571.950 618.450 574.050 619.050 ;
        RECT 628.950 618.450 631.050 619.200 ;
        RECT 571.950 617.400 631.050 618.450 ;
        RECT 571.950 616.950 574.050 617.400 ;
        RECT 628.950 617.100 631.050 617.400 ;
        RECT 535.950 576.450 538.050 577.050 ;
        RECT 571.950 576.450 574.050 577.050 ;
        RECT 535.950 575.400 574.050 576.450 ;
        RECT 535.950 574.950 538.050 575.400 ;
        RECT 571.950 574.950 574.050 575.400 ;
        RECT 563.100 523.950 568.050 526.050 ;
        RECT 529.950 513.450 532.050 514.050 ;
        RECT 535.950 513.450 538.050 514.050 ;
        RECT 565.800 513.450 567.900 514.050 ;
        RECT 529.950 512.400 567.900 513.450 ;
        RECT 529.950 511.950 532.050 512.400 ;
        RECT 535.950 511.950 538.050 512.400 ;
        RECT 565.800 511.950 567.900 512.400 ;
        RECT 475.950 495.450 478.050 496.050 ;
        RECT 529.950 495.450 532.050 496.050 ;
        RECT 475.950 494.400 532.050 495.450 ;
        RECT 475.950 493.950 478.050 494.400 ;
        RECT 529.950 493.950 532.050 494.400 ;
        RECT 529.950 484.950 532.050 490.050 ;
        RECT 415.950 450.450 418.050 454.050 ;
        RECT 436.950 453.450 439.050 454.050 ;
        RECT 448.950 453.450 451.050 454.050 ;
        RECT 436.950 452.400 451.050 453.450 ;
        RECT 436.950 451.950 439.050 452.400 ;
        RECT 448.950 451.950 451.050 452.400 ;
        RECT 473.100 453.450 475.200 454.050 ;
        RECT 475.950 453.450 481.050 454.050 ;
        RECT 473.100 452.400 481.050 453.450 ;
        RECT 473.100 451.950 475.200 452.400 ;
        RECT 475.950 451.950 481.050 452.400 ;
        RECT 436.950 450.450 439.050 451.050 ;
        RECT 415.950 450.000 439.050 450.450 ;
        RECT 416.400 449.400 439.050 450.000 ;
        RECT 436.950 448.950 439.050 449.400 ;
        RECT 448.950 441.450 451.050 442.050 ;
        RECT 478.950 441.450 481.050 442.050 ;
        RECT 505.950 441.450 508.050 442.050 ;
        RECT 448.950 440.400 508.050 441.450 ;
        RECT 448.950 439.950 451.050 440.400 ;
        RECT 478.950 439.950 481.050 440.400 ;
        RECT 505.950 439.950 508.050 440.400 ;
        RECT 562.950 381.450 565.050 382.050 ;
        RECT 568.950 381.450 571.050 382.050 ;
        RECT 562.950 380.400 571.050 381.450 ;
        RECT 562.950 379.950 565.050 380.400 ;
        RECT 568.950 379.950 571.050 380.400 ;
        RECT 505.950 348.450 508.050 349.050 ;
        RECT 505.950 347.400 534.450 348.450 ;
        RECT 505.950 346.950 508.050 347.400 ;
        RECT 533.400 345.450 534.450 347.400 ;
        RECT 541.950 345.450 544.050 346.050 ;
        RECT 533.400 344.400 544.050 345.450 ;
        RECT 541.950 343.950 544.050 344.400 ;
        RECT 514.950 315.450 517.050 316.050 ;
        RECT 540.000 315.450 544.050 316.050 ;
        RECT 514.950 314.400 544.050 315.450 ;
        RECT 514.950 313.950 517.050 314.400 ;
        RECT 539.400 313.950 544.050 314.400 ;
        RECT 539.400 312.450 540.450 313.950 ;
        RECT 544.950 312.450 547.050 313.050 ;
        RECT 568.800 312.450 570.900 313.050 ;
        RECT 539.400 311.400 570.900 312.450 ;
        RECT 544.950 310.950 547.050 311.400 ;
        RECT 568.800 310.950 570.900 311.400 ;
        RECT 514.950 270.450 517.050 271.050 ;
        RECT 503.400 270.000 517.050 270.450 ;
        RECT 502.950 269.400 517.050 270.000 ;
        RECT 502.950 265.950 505.050 269.400 ;
        RECT 514.950 268.950 517.050 269.400 ;
        RECT 515.400 268.050 516.450 268.950 ;
        RECT 515.400 265.950 520.050 268.050 ;
        RECT 515.400 265.050 516.450 265.950 ;
        RECT 513.000 264.900 516.450 265.050 ;
        RECT 511.950 263.400 516.450 264.900 ;
        RECT 511.950 262.950 516.000 263.400 ;
        RECT 511.950 262.800 514.050 262.950 ;
        RECT 508.950 235.950 514.050 238.050 ;
        RECT 496.950 216.450 499.050 217.050 ;
        RECT 511.950 216.450 514.050 217.200 ;
        RECT 496.950 215.400 514.050 216.450 ;
        RECT 496.950 214.950 499.050 215.400 ;
        RECT 511.950 215.100 514.050 215.400 ;
        RECT 604.950 169.950 610.050 172.050 ;
        RECT 493.950 162.450 496.050 163.050 ;
        RECT 502.950 162.450 505.050 166.050 ;
        RECT 547.950 162.450 550.050 163.050 ;
        RECT 493.950 161.400 550.050 162.450 ;
        RECT 493.950 160.950 496.050 161.400 ;
        RECT 547.950 160.950 550.050 161.400 ;
        RECT 551.100 150.450 553.200 151.050 ;
        RECT 604.950 150.450 607.050 151.050 ;
        RECT 551.100 149.400 607.050 150.450 ;
        RECT 551.100 148.950 553.200 149.400 ;
        RECT 604.950 148.950 607.050 149.400 ;
        RECT 394.950 138.450 397.050 139.050 ;
        RECT 490.950 138.450 493.050 139.050 ;
        RECT 394.950 137.400 493.050 138.450 ;
        RECT 394.950 136.950 397.050 137.400 ;
        RECT 490.950 136.950 493.050 137.400 ;
        RECT 394.950 129.450 397.050 130.050 ;
        RECT 492.000 129.450 495.900 130.050 ;
        RECT 389.250 129.000 397.050 129.450 ;
        RECT 491.550 129.000 495.900 129.450 ;
        RECT 388.950 128.400 397.050 129.000 ;
        RECT 388.950 127.050 391.050 128.400 ;
        RECT 394.950 127.950 397.050 128.400 ;
        RECT 490.950 127.950 495.900 129.000 ;
        RECT 388.800 126.000 391.050 127.050 ;
        RECT 490.950 127.050 493.050 127.950 ;
        RECT 490.950 126.000 493.200 127.050 ;
        RECT 388.800 124.950 390.900 126.000 ;
        RECT 491.100 124.950 493.200 126.000 ;
      LAYER metal3 ;
        RECT 646.950 862.950 649.050 865.050 ;
        RECT 647.400 717.600 648.600 862.950 ;
        RECT 758.400 862.200 759.600 873.600 ;
        RECT 757.950 860.100 760.050 862.200 ;
        RECT 644.400 716.400 648.600 717.600 ;
        RECT 644.400 688.050 645.600 716.400 ;
        RECT 628.950 685.950 631.050 688.050 ;
        RECT 643.950 685.950 646.050 688.050 ;
        RECT 629.400 619.200 630.600 685.950 ;
        RECT 571.950 616.950 574.050 619.050 ;
        RECT 628.950 617.100 631.050 619.200 ;
        RECT 572.400 577.050 573.600 616.950 ;
        RECT 535.950 574.950 538.050 577.050 ;
        RECT 571.950 574.950 574.050 577.050 ;
        RECT 536.400 514.050 537.600 574.950 ;
        RECT 563.100 525.600 567.000 526.050 ;
        RECT 563.100 523.950 567.600 525.600 ;
        RECT 566.400 514.050 567.600 523.950 ;
        RECT 529.950 511.950 532.050 514.050 ;
        RECT 535.950 511.950 538.050 514.050 ;
        RECT 565.800 511.950 567.900 514.050 ;
        RECT 530.400 496.050 531.600 511.950 ;
        RECT 475.950 493.950 478.050 496.050 ;
        RECT 529.950 493.950 532.050 496.050 ;
        RECT 476.400 454.050 477.600 493.950 ;
        RECT 530.400 490.050 531.600 493.950 ;
        RECT 529.950 487.950 532.050 490.050 ;
        RECT 448.950 451.950 451.050 454.050 ;
        RECT 475.950 451.950 478.050 454.050 ;
        RECT 449.400 442.050 450.600 451.950 ;
        RECT 448.950 439.950 451.050 442.050 ;
        RECT 505.950 439.950 508.050 442.050 ;
        RECT 506.400 349.050 507.600 439.950 ;
        RECT 568.950 379.950 571.050 382.050 ;
        RECT 505.950 346.950 508.050 349.050 ;
        RECT 541.950 343.950 544.050 346.050 ;
        RECT 542.400 316.050 543.600 343.950 ;
        RECT 514.950 313.950 517.050 316.050 ;
        RECT 541.950 313.950 544.050 316.050 ;
        RECT 515.400 271.050 516.600 313.950 ;
        RECT 569.400 313.050 570.600 379.950 ;
        RECT 568.800 310.950 570.900 313.050 ;
        RECT 514.950 268.950 517.050 271.050 ;
        RECT 511.950 262.800 514.050 264.900 ;
        RECT 512.400 238.050 513.600 262.800 ;
        RECT 511.950 235.950 514.050 238.050 ;
        RECT 512.400 217.200 513.600 235.950 ;
        RECT 496.950 214.950 499.050 217.050 ;
        RECT 511.950 215.100 514.050 217.200 ;
        RECT 497.400 195.600 498.600 214.950 ;
        RECT 494.400 194.400 498.600 195.600 ;
        RECT 494.400 163.050 495.600 194.400 ;
        RECT 604.950 169.950 607.050 172.050 ;
        RECT 493.950 162.600 496.050 163.050 ;
        RECT 491.400 161.400 496.050 162.600 ;
        RECT 491.400 139.050 492.600 161.400 ;
        RECT 493.950 160.950 496.050 161.400 ;
        RECT 547.950 160.950 550.050 163.050 ;
        RECT 548.400 153.600 549.600 160.950 ;
        RECT 548.400 153.000 552.600 153.600 ;
        RECT 548.400 152.400 553.050 153.000 ;
        RECT 550.950 151.050 553.050 152.400 ;
        RECT 605.400 151.050 606.600 169.950 ;
        RECT 550.950 150.000 553.200 151.050 ;
        RECT 551.100 148.950 553.200 150.000 ;
        RECT 604.950 148.950 607.050 151.050 ;
        RECT 394.950 136.950 397.050 139.050 ;
        RECT 490.950 136.950 493.050 139.050 ;
        RECT 395.400 130.050 396.600 136.950 ;
        RECT 491.400 135.600 492.600 136.950 ;
        RECT 491.400 134.400 495.600 135.600 ;
        RECT 494.400 130.050 495.600 134.400 ;
        RECT 394.950 127.950 397.050 130.050 ;
        RECT 493.800 127.950 495.900 130.050 ;
    END
  END ABCmd_i[7]
  PIN ABCmd_i[6]
    PORT
      LAYER metal1 ;
        RECT 694.950 694.950 697.050 697.050 ;
        RECT 544.950 187.950 547.050 193.050 ;
        RECT 556.950 127.950 559.050 130.050 ;
        RECT 583.950 52.950 586.050 55.050 ;
        RECT 595.950 52.950 598.050 55.050 ;
      LAYER metal2 ;
        RECT 745.950 864.450 748.050 865.050 ;
        RECT 763.950 864.450 766.050 865.050 ;
        RECT 745.950 863.400 766.050 864.450 ;
        RECT 745.950 862.950 748.050 863.400 ;
        RECT 763.950 862.950 766.050 863.400 ;
        RECT 724.950 834.450 727.050 835.050 ;
        RECT 745.950 834.450 748.050 835.050 ;
        RECT 724.950 833.400 748.050 834.450 ;
        RECT 724.950 832.950 727.050 833.400 ;
        RECT 745.950 832.950 748.050 833.400 ;
        RECT 706.950 756.450 709.050 757.050 ;
        RECT 724.950 756.450 727.050 757.050 ;
        RECT 706.950 755.400 727.050 756.450 ;
        RECT 706.950 754.950 709.050 755.400 ;
        RECT 724.950 754.950 727.050 755.400 ;
        RECT 691.950 750.450 694.050 751.050 ;
        RECT 706.950 750.450 709.050 751.050 ;
        RECT 691.950 749.400 709.050 750.450 ;
        RECT 691.950 748.950 694.050 749.400 ;
        RECT 706.950 748.950 709.050 749.400 ;
        RECT 670.950 696.450 673.050 697.050 ;
        RECT 691.950 696.450 697.050 697.050 ;
        RECT 670.950 695.400 697.050 696.450 ;
        RECT 670.950 694.950 673.050 695.400 ;
        RECT 691.950 694.950 697.050 695.400 ;
        RECT 664.950 657.450 667.050 658.050 ;
        RECT 670.950 657.450 673.050 658.050 ;
        RECT 664.950 656.400 673.050 657.450 ;
        RECT 664.950 655.950 667.050 656.400 ;
        RECT 670.950 655.950 673.050 656.400 ;
        RECT 569.100 513.450 571.200 514.050 ;
        RECT 661.950 513.450 664.050 514.050 ;
        RECT 569.100 512.400 664.050 513.450 ;
        RECT 569.100 511.950 571.200 512.400 ;
        RECT 661.950 511.950 664.050 512.400 ;
        RECT 523.950 462.450 526.050 463.050 ;
        RECT 568.950 462.450 571.050 463.050 ;
        RECT 523.950 461.400 571.050 462.450 ;
        RECT 523.950 460.950 526.050 461.400 ;
        RECT 568.950 460.950 571.050 461.400 ;
        RECT 523.950 363.450 526.050 364.050 ;
        RECT 562.950 363.450 565.050 364.050 ;
        RECT 523.950 362.400 565.050 363.450 ;
        RECT 523.950 361.950 526.050 362.400 ;
        RECT 562.950 361.950 565.050 362.400 ;
        RECT 562.950 327.450 565.050 328.050 ;
        RECT 616.950 327.450 619.050 328.050 ;
        RECT 562.950 326.400 619.050 327.450 ;
        RECT 562.950 325.950 565.050 326.400 ;
        RECT 616.950 325.950 619.050 326.400 ;
        RECT 616.950 297.450 619.050 298.200 ;
        RECT 625.950 297.450 628.050 297.900 ;
        RECT 616.950 296.400 628.050 297.450 ;
        RECT 616.950 296.100 619.050 296.400 ;
        RECT 625.950 295.800 628.050 296.400 ;
        RECT 604.950 216.450 607.050 217.050 ;
        RECT 625.950 216.450 628.050 217.050 ;
        RECT 604.950 215.400 628.050 216.450 ;
        RECT 604.950 214.950 607.050 215.400 ;
        RECT 625.950 214.950 628.050 215.400 ;
        RECT 544.950 189.450 547.050 190.050 ;
        RECT 553.950 189.450 556.050 190.050 ;
        RECT 604.950 189.450 607.050 190.050 ;
        RECT 544.950 188.400 607.050 189.450 ;
        RECT 544.950 187.950 547.050 188.400 ;
        RECT 553.950 187.950 556.050 188.400 ;
        RECT 604.950 187.950 607.050 188.400 ;
        RECT 553.950 127.950 559.050 130.050 ;
        RECT 556.950 63.450 559.050 64.050 ;
        RECT 583.950 63.450 586.050 64.050 ;
        RECT 556.950 62.400 586.050 63.450 ;
        RECT 556.950 61.950 559.050 62.400 ;
        RECT 583.950 61.950 586.050 62.400 ;
        RECT 583.950 54.450 589.050 55.050 ;
        RECT 595.950 54.450 598.050 55.050 ;
        RECT 583.950 53.400 598.050 54.450 ;
        RECT 583.950 52.950 589.050 53.400 ;
        RECT 595.950 52.950 598.050 53.400 ;
      LAYER metal3 ;
        RECT 764.400 865.050 765.600 873.600 ;
        RECT 745.950 862.950 748.050 865.050 ;
        RECT 763.950 862.950 766.050 865.050 ;
        RECT 746.400 835.050 747.600 862.950 ;
        RECT 724.950 832.950 727.050 835.050 ;
        RECT 745.950 832.950 748.050 835.050 ;
        RECT 725.400 757.050 726.600 832.950 ;
        RECT 706.950 754.950 709.050 757.050 ;
        RECT 724.950 754.950 727.050 757.050 ;
        RECT 707.400 751.050 708.600 754.950 ;
        RECT 691.950 748.950 694.050 751.050 ;
        RECT 706.950 748.950 709.050 751.050 ;
        RECT 692.400 697.050 693.600 748.950 ;
        RECT 670.950 694.950 673.050 697.050 ;
        RECT 691.950 694.950 694.050 697.050 ;
        RECT 671.400 658.050 672.600 694.950 ;
        RECT 664.950 655.950 667.050 658.050 ;
        RECT 670.950 655.950 673.050 658.050 ;
        RECT 665.400 615.600 666.600 655.950 ;
        RECT 662.400 614.400 666.600 615.600 ;
        RECT 662.400 514.050 663.600 614.400 ;
        RECT 569.100 511.950 571.200 514.050 ;
        RECT 661.950 511.950 664.050 514.050 ;
        RECT 569.400 463.050 570.600 511.950 ;
        RECT 523.950 460.950 526.050 463.050 ;
        RECT 568.950 460.950 571.050 463.050 ;
        RECT 524.400 364.050 525.600 460.950 ;
        RECT 523.950 361.950 526.050 364.050 ;
        RECT 562.950 361.950 565.050 364.050 ;
        RECT 563.400 328.050 564.600 361.950 ;
        RECT 562.950 325.950 565.050 328.050 ;
        RECT 616.950 325.950 619.050 328.050 ;
        RECT 617.400 298.200 618.600 325.950 ;
        RECT 616.950 296.100 619.050 298.200 ;
        RECT 625.950 295.800 628.050 297.900 ;
        RECT 626.400 217.050 627.600 295.800 ;
        RECT 604.950 214.950 607.050 217.050 ;
        RECT 625.950 214.950 628.050 217.050 ;
        RECT 605.400 190.050 606.600 214.950 ;
        RECT 553.950 187.950 556.050 190.050 ;
        RECT 604.950 187.950 607.050 190.050 ;
        RECT 554.400 130.050 555.600 187.950 ;
        RECT 553.950 127.950 556.050 130.050 ;
        RECT 554.400 102.600 555.600 127.950 ;
        RECT 554.400 101.400 558.600 102.600 ;
        RECT 557.400 64.050 558.600 101.400 ;
        RECT 556.950 61.950 559.050 64.050 ;
        RECT 583.950 61.950 586.050 64.050 ;
        RECT 584.400 55.050 585.600 61.950 ;
        RECT 584.400 53.400 589.050 55.050 ;
        RECT 585.000 52.950 589.050 53.400 ;
    END
  END ABCmd_i[6]
  PIN ABCmd_i[5]
    PORT
      LAYER metal1 ;
        RECT 832.950 844.950 835.050 847.050 ;
        RECT 793.950 745.950 796.050 748.050 ;
        RECT 841.950 520.950 844.050 523.050 ;
        RECT 853.950 499.950 856.050 502.050 ;
        RECT 703.950 487.950 706.050 490.050 ;
        RECT 829.950 483.450 832.050 484.050 ;
        RECT 834.000 483.450 838.050 484.050 ;
        RECT 829.950 482.550 838.050 483.450 ;
        RECT 829.950 481.950 832.050 482.550 ;
        RECT 834.000 481.950 838.050 482.550 ;
        RECT 847.950 483.450 850.050 484.050 ;
        RECT 854.550 483.450 855.450 499.950 ;
        RECT 847.950 482.550 855.450 483.450 ;
        RECT 847.950 481.950 850.050 482.550 ;
        RECT 679.950 420.000 682.050 424.050 ;
        RECT 748.950 421.950 751.050 424.050 ;
        RECT 680.550 418.050 681.450 420.000 ;
        RECT 679.950 415.950 682.050 418.050 ;
        RECT 749.550 406.050 750.450 421.950 ;
        RECT 748.950 403.950 751.050 406.050 ;
        RECT 709.950 376.950 712.050 379.050 ;
        RECT 769.800 376.950 772.050 379.050 ;
        RECT 649.950 352.950 652.050 355.050 ;
        RECT 650.550 334.050 651.450 352.950 ;
        RECT 649.950 331.950 652.050 334.050 ;
        RECT 706.950 304.950 709.050 307.050 ;
        RECT 733.800 304.950 736.050 307.050 ;
      LAYER metal2 ;
        RECT 790.950 861.450 793.050 862.050 ;
        RECT 829.950 861.450 832.050 862.050 ;
        RECT 790.950 860.400 832.050 861.450 ;
        RECT 790.950 859.950 793.050 860.400 ;
        RECT 829.950 859.950 832.050 860.400 ;
        RECT 829.950 844.950 835.050 847.050 ;
        RECT 799.950 750.450 802.050 751.050 ;
        RECT 856.950 750.450 859.050 751.050 ;
        RECT 799.950 749.400 859.050 750.450 ;
        RECT 799.950 748.950 802.050 749.400 ;
        RECT 856.950 748.950 859.050 749.400 ;
        RECT 793.950 747.450 796.050 748.050 ;
        RECT 800.400 747.450 801.450 748.950 ;
        RECT 793.950 746.400 801.450 747.450 ;
        RECT 793.950 745.950 796.050 746.400 ;
        RECT 838.950 564.450 841.050 565.050 ;
        RECT 856.950 564.450 859.050 565.050 ;
        RECT 838.950 563.400 859.050 564.450 ;
        RECT 838.950 562.950 841.050 563.400 ;
        RECT 856.950 562.950 859.050 563.400 ;
        RECT 838.950 520.950 844.050 523.050 ;
        RECT 838.950 501.450 841.050 502.050 ;
        RECT 853.950 501.450 856.050 502.050 ;
        RECT 838.950 500.400 856.050 501.450 ;
        RECT 838.950 499.950 841.050 500.400 ;
        RECT 853.950 499.950 856.050 500.400 ;
        RECT 662.100 498.450 664.200 499.050 ;
        RECT 662.100 497.400 687.450 498.450 ;
        RECT 662.100 496.950 664.200 497.400 ;
        RECT 686.400 495.450 687.450 497.400 ;
        RECT 694.800 495.450 696.900 496.050 ;
        RECT 686.400 494.400 696.900 495.450 ;
        RECT 694.800 493.950 696.900 494.400 ;
        RECT 702.000 489.450 706.050 490.050 ;
        RECT 701.400 487.950 706.050 489.450 ;
        RECT 694.950 486.450 697.050 487.050 ;
        RECT 701.400 486.450 702.450 487.950 ;
        RECT 694.950 485.400 702.450 486.450 ;
        RECT 694.950 484.950 697.050 485.400 ;
        RECT 835.950 481.950 840.900 484.050 ;
        RECT 751.950 468.450 754.050 469.050 ;
        RECT 751.950 467.400 792.450 468.450 ;
        RECT 751.950 466.950 754.050 467.400 ;
        RECT 791.400 465.450 792.450 467.400 ;
        RECT 838.950 465.450 841.050 466.050 ;
        RECT 791.400 464.400 841.050 465.450 ;
        RECT 838.950 463.950 841.050 464.400 ;
        RECT 658.950 423.450 661.050 424.050 ;
        RECT 679.950 423.450 682.050 424.050 ;
        RECT 658.950 422.400 682.050 423.450 ;
        RECT 658.950 421.950 661.050 422.400 ;
        RECT 679.950 421.950 682.050 422.400 ;
        RECT 748.950 423.450 751.050 424.050 ;
        RECT 754.950 423.450 757.050 424.050 ;
        RECT 748.950 422.400 757.050 423.450 ;
        RECT 748.950 421.950 751.050 422.400 ;
        RECT 754.950 421.950 757.050 422.400 ;
        RECT 679.950 417.450 682.050 418.050 ;
        RECT 685.950 417.450 688.050 418.050 ;
        RECT 679.950 416.400 688.050 417.450 ;
        RECT 679.950 415.950 682.050 416.400 ;
        RECT 685.950 415.950 688.050 416.400 ;
        RECT 727.950 405.450 730.050 406.050 ;
        RECT 748.950 405.450 751.050 406.050 ;
        RECT 763.950 405.450 766.050 406.050 ;
        RECT 727.950 404.400 766.050 405.450 ;
        RECT 727.950 403.950 730.050 404.400 ;
        RECT 748.950 403.950 751.050 404.400 ;
        RECT 763.950 403.950 766.050 404.400 ;
        RECT 664.950 396.450 667.050 397.050 ;
        RECT 685.950 396.450 688.050 397.050 ;
        RECT 727.950 396.450 730.050 397.050 ;
        RECT 664.950 395.400 730.050 396.450 ;
        RECT 664.950 394.950 667.050 395.400 ;
        RECT 685.950 394.950 688.050 395.400 ;
        RECT 727.950 394.950 730.050 395.400 ;
        RECT 709.950 378.450 712.050 379.050 ;
        RECT 727.950 378.450 730.050 379.050 ;
        RECT 709.950 377.400 730.050 378.450 ;
        RECT 709.950 376.950 712.050 377.400 ;
        RECT 727.950 376.950 730.050 377.400 ;
        RECT 769.800 378.000 771.900 379.050 ;
        RECT 769.800 376.950 772.050 378.000 ;
        RECT 619.950 375.450 622.050 376.050 ;
        RECT 763.950 375.450 766.050 376.050 ;
        RECT 769.950 375.450 772.050 376.950 ;
        RECT 619.950 374.400 627.450 375.450 ;
        RECT 619.950 373.950 622.050 374.400 ;
        RECT 626.400 372.450 627.450 374.400 ;
        RECT 763.950 375.000 772.050 375.450 ;
        RECT 763.950 374.400 771.300 375.000 ;
        RECT 763.950 373.950 766.050 374.400 ;
        RECT 664.950 372.450 667.050 373.050 ;
        RECT 626.400 371.400 667.050 372.450 ;
        RECT 664.950 370.950 667.050 371.400 ;
        RECT 619.950 354.450 622.050 355.050 ;
        RECT 649.950 354.450 652.050 355.050 ;
        RECT 619.950 353.400 652.050 354.450 ;
        RECT 619.950 352.950 622.050 353.400 ;
        RECT 649.950 352.950 652.050 353.400 ;
        RECT 649.950 333.450 652.050 334.050 ;
        RECT 682.950 333.450 685.050 334.050 ;
        RECT 649.950 332.400 685.050 333.450 ;
        RECT 649.950 331.950 652.050 332.400 ;
        RECT 682.950 331.950 685.050 332.400 ;
        RECT 682.950 324.450 685.050 325.050 ;
        RECT 700.950 324.450 703.050 325.050 ;
        RECT 727.800 324.450 729.900 325.050 ;
        RECT 682.950 323.400 729.900 324.450 ;
        RECT 682.950 322.950 685.050 323.400 ;
        RECT 700.950 322.950 703.050 323.400 ;
        RECT 727.800 322.950 729.900 323.400 ;
        RECT 700.950 306.450 703.050 307.050 ;
        RECT 706.950 306.450 709.050 307.050 ;
        RECT 700.950 305.400 709.050 306.450 ;
        RECT 700.950 304.950 703.050 305.400 ;
        RECT 706.950 304.950 709.050 305.400 ;
        RECT 731.100 304.950 735.900 307.050 ;
      LAYER metal3 ;
        RECT 791.400 862.050 792.600 873.600 ;
        RECT 790.950 859.950 793.050 862.050 ;
        RECT 829.950 859.950 832.050 862.050 ;
        RECT 791.400 858.600 792.600 859.950 ;
        RECT 791.400 857.400 798.600 858.600 ;
        RECT 797.400 840.600 798.600 857.400 ;
        RECT 830.400 847.050 831.600 859.950 ;
        RECT 829.950 844.950 832.050 847.050 ;
        RECT 797.400 839.400 801.600 840.600 ;
        RECT 800.400 751.050 801.600 839.400 ;
        RECT 799.950 748.950 802.050 751.050 ;
        RECT 856.950 748.950 859.050 751.050 ;
        RECT 857.400 565.050 858.600 748.950 ;
        RECT 838.950 562.950 841.050 565.050 ;
        RECT 856.950 562.950 859.050 565.050 ;
        RECT 839.400 523.050 840.600 562.950 ;
        RECT 838.950 520.950 841.050 523.050 ;
        RECT 839.400 502.050 840.600 520.950 ;
        RECT 838.950 499.950 841.050 502.050 ;
        RECT 662.100 496.950 664.200 499.050 ;
        RECT 662.400 483.600 663.600 496.950 ;
        RECT 694.800 493.950 696.900 496.050 ;
        RECT 695.400 487.050 696.600 493.950 ;
        RECT 694.950 484.950 697.050 487.050 ;
        RECT 839.400 484.050 840.600 499.950 ;
        RECT 659.400 482.400 663.600 483.600 ;
        RECT 659.400 424.050 660.600 482.400 ;
        RECT 838.800 481.950 840.900 484.050 ;
        RECT 751.950 466.950 754.050 469.050 ;
        RECT 752.400 447.600 753.600 466.950 ;
        RECT 839.400 466.050 840.600 481.950 ;
        RECT 838.950 463.950 841.050 466.050 ;
        RECT 752.400 446.400 756.600 447.600 ;
        RECT 755.400 424.050 756.600 446.400 ;
        RECT 658.950 421.950 661.050 424.050 ;
        RECT 754.950 421.950 757.050 424.050 ;
        RECT 685.950 415.950 688.050 418.050 ;
        RECT 686.400 397.050 687.600 415.950 ;
        RECT 727.950 403.950 730.050 406.050 ;
        RECT 763.950 403.950 766.050 406.050 ;
        RECT 728.400 397.050 729.600 403.950 ;
        RECT 664.950 394.950 667.050 397.050 ;
        RECT 685.950 394.950 688.050 397.050 ;
        RECT 727.950 394.950 730.050 397.050 ;
        RECT 619.950 373.950 622.050 376.050 ;
        RECT 620.400 355.050 621.600 373.950 ;
        RECT 665.400 373.050 666.600 394.950 ;
        RECT 728.400 379.050 729.600 394.950 ;
        RECT 727.950 376.950 730.050 379.050 ;
        RECT 764.400 376.050 765.600 403.950 ;
        RECT 763.950 373.950 766.050 376.050 ;
        RECT 664.950 370.950 667.050 373.050 ;
        RECT 619.950 352.950 622.050 355.050 ;
        RECT 682.950 331.950 685.050 334.050 ;
        RECT 683.400 325.050 684.600 331.950 ;
        RECT 682.950 322.950 685.050 325.050 ;
        RECT 700.950 322.950 703.050 325.050 ;
        RECT 727.800 324.000 729.900 325.050 ;
        RECT 727.800 322.950 730.050 324.000 ;
        RECT 701.400 307.050 702.600 322.950 ;
        RECT 727.950 321.600 730.050 322.950 ;
        RECT 727.950 321.000 732.600 321.600 ;
        RECT 728.400 320.400 732.600 321.000 ;
        RECT 731.400 307.050 732.600 320.400 ;
        RECT 700.950 304.950 703.050 307.050 ;
        RECT 731.100 304.950 733.200 307.050 ;
    END
  END ABCmd_i[5]
  PIN ABCmd_i[4]
    PORT
      LAYER metal1 ;
        RECT 808.950 694.950 811.050 697.050 ;
        RECT 829.950 523.950 832.050 526.050 ;
        RECT 830.550 522.000 831.450 523.950 ;
        RECT 829.950 517.950 832.050 522.000 ;
        RECT 847.950 520.950 850.050 523.050 ;
      LAYER metal2 ;
        RECT 814.950 741.450 817.050 742.050 ;
        RECT 820.800 741.450 822.900 742.050 ;
        RECT 814.950 740.400 822.900 741.450 ;
        RECT 814.950 739.950 817.050 740.400 ;
        RECT 820.800 739.950 822.900 740.400 ;
        RECT 808.950 696.450 811.050 697.050 ;
        RECT 814.950 696.450 817.050 697.050 ;
        RECT 808.950 695.400 817.050 696.450 ;
        RECT 808.950 691.950 811.050 695.400 ;
        RECT 814.950 694.950 817.050 695.400 ;
        RECT 808.950 621.450 811.050 622.050 ;
        RECT 829.950 621.450 832.050 622.050 ;
        RECT 808.950 620.400 832.050 621.450 ;
        RECT 808.950 619.950 811.050 620.400 ;
        RECT 829.950 619.950 832.050 620.400 ;
        RECT 829.950 519.450 832.050 520.050 ;
        RECT 847.950 519.450 850.050 523.050 ;
        RECT 829.950 519.000 850.050 519.450 ;
        RECT 829.950 518.400 849.450 519.000 ;
        RECT 829.950 517.950 832.050 518.400 ;
      LAYER metal3 ;
        RECT 821.400 742.050 822.600 873.600 ;
        RECT 814.950 739.950 817.050 742.050 ;
        RECT 820.800 739.950 822.900 742.050 ;
        RECT 815.400 697.050 816.600 739.950 ;
        RECT 814.950 694.950 817.050 697.050 ;
        RECT 808.950 691.950 811.050 694.050 ;
        RECT 809.400 622.050 810.600 691.950 ;
        RECT 808.950 619.950 811.050 622.050 ;
        RECT 829.950 619.950 832.050 622.050 ;
        RECT 830.400 520.050 831.600 619.950 ;
        RECT 829.950 517.950 832.050 520.050 ;
    END
  END ABCmd_i[4]
  PIN ABCmd_i[3]
    PORT
      LAYER metal1 ;
        RECT 826.950 817.950 829.050 820.050 ;
        RECT 827.550 808.050 828.450 817.950 ;
        RECT 826.950 805.950 829.050 808.050 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 817.950 595.950 823.050 598.050 ;
      LAYER metal2 ;
        RECT 826.950 817.950 829.050 823.050 ;
        RECT 826.950 807.450 829.050 808.050 ;
        RECT 847.950 807.450 850.050 808.050 ;
        RECT 826.950 806.400 850.050 807.450 ;
        RECT 826.950 805.950 829.050 806.400 ;
        RECT 847.950 805.950 850.050 806.400 ;
        RECT 811.950 654.450 814.050 655.050 ;
        RECT 847.950 654.450 850.050 655.050 ;
        RECT 811.950 653.400 850.050 654.450 ;
        RECT 811.950 652.950 814.050 653.400 ;
        RECT 847.950 652.950 850.050 653.400 ;
        RECT 811.950 598.950 814.050 604.050 ;
        RECT 812.100 597.450 814.200 598.050 ;
        RECT 817.950 597.450 820.050 598.050 ;
        RECT 812.100 596.400 820.050 597.450 ;
        RECT 812.100 595.950 814.200 596.400 ;
        RECT 817.950 595.950 820.050 596.400 ;
      LAYER metal3 ;
        RECT 827.400 823.050 828.600 873.600 ;
        RECT 826.950 820.950 829.050 823.050 ;
        RECT 847.950 805.950 850.050 808.050 ;
        RECT 848.400 655.050 849.600 805.950 ;
        RECT 811.950 652.950 814.050 655.050 ;
        RECT 847.950 652.950 850.050 655.050 ;
        RECT 812.400 601.050 813.600 652.950 ;
        RECT 811.950 598.050 814.050 601.050 ;
        RECT 811.950 597.000 814.200 598.050 ;
        RECT 812.100 595.950 814.200 597.000 ;
    END
  END ABCmd_i[3]
  PIN ABCmd_i[2]
    PORT
      LAYER metal1 ;
        RECT 751.950 382.950 754.050 385.050 ;
        RECT 718.800 265.950 721.050 268.050 ;
        RECT 778.950 265.950 781.050 268.050 ;
        RECT 823.950 265.950 826.050 268.050 ;
      LAYER metal2 ;
        RECT 790.950 387.450 793.050 388.050 ;
        RECT 758.400 386.400 793.050 387.450 ;
        RECT 751.950 384.450 754.050 385.050 ;
        RECT 758.400 384.450 759.450 386.400 ;
        RECT 790.950 385.950 793.050 386.400 ;
        RECT 751.950 383.400 759.450 384.450 ;
        RECT 751.950 382.950 754.050 383.400 ;
        RECT 790.950 363.450 793.050 364.050 ;
        RECT 844.950 363.450 847.050 364.050 ;
        RECT 790.950 362.400 847.050 363.450 ;
        RECT 790.950 361.950 793.050 362.400 ;
        RECT 844.950 361.950 847.050 362.400 ;
        RECT 829.950 306.450 832.050 307.050 ;
        RECT 844.950 306.450 847.050 307.050 ;
        RECT 829.950 305.400 847.050 306.450 ;
        RECT 829.950 304.950 832.050 305.400 ;
        RECT 844.950 304.950 847.050 305.400 ;
        RECT 715.950 279.450 718.050 280.050 ;
        RECT 778.950 279.450 781.050 280.050 ;
        RECT 829.950 279.450 832.050 280.050 ;
        RECT 856.950 279.450 859.050 280.050 ;
        RECT 715.950 278.400 859.050 279.450 ;
        RECT 715.950 277.950 718.050 278.400 ;
        RECT 778.950 277.950 781.050 278.400 ;
        RECT 829.950 277.950 832.050 278.400 ;
        RECT 856.950 277.950 859.050 278.400 ;
        RECT 856.950 270.450 859.050 271.050 ;
        RECT 856.950 269.400 864.450 270.450 ;
        RECT 856.950 268.950 859.050 269.400 ;
        RECT 716.100 265.950 720.900 268.050 ;
        RECT 778.950 265.950 783.900 268.050 ;
        RECT 823.950 267.450 826.050 268.050 ;
        RECT 829.950 267.450 832.050 268.050 ;
        RECT 823.950 266.400 832.050 267.450 ;
        RECT 823.950 265.950 826.050 266.400 ;
        RECT 829.950 265.950 832.050 266.400 ;
      LAYER metal3 ;
        RECT 790.950 385.950 793.050 388.050 ;
        RECT 791.400 364.050 792.600 385.950 ;
        RECT 790.950 361.950 793.050 364.050 ;
        RECT 844.950 361.950 847.050 364.050 ;
        RECT 845.400 307.050 846.600 361.950 ;
        RECT 829.950 304.950 832.050 307.050 ;
        RECT 844.950 304.950 847.050 307.050 ;
        RECT 830.400 280.050 831.600 304.950 ;
        RECT 715.950 277.950 718.050 280.050 ;
        RECT 778.950 277.950 781.050 280.050 ;
        RECT 829.950 277.950 832.050 280.050 ;
        RECT 856.950 277.950 859.050 280.050 ;
        RECT 716.400 268.050 717.600 277.950 ;
        RECT 779.400 268.050 780.600 277.950 ;
        RECT 830.400 268.050 831.600 277.950 ;
        RECT 857.400 271.050 858.600 277.950 ;
        RECT 856.950 268.950 859.050 271.050 ;
        RECT 716.100 265.950 718.200 268.050 ;
        RECT 779.400 266.400 783.900 268.050 ;
        RECT 780.000 265.950 783.900 266.400 ;
        RECT 829.950 265.950 832.050 268.050 ;
    END
  END ABCmd_i[2]
  PIN ABCmd_i[1]
    PORT
      LAYER metal1 ;
        RECT 685.950 487.950 688.050 490.050 ;
        RECT 673.950 478.950 676.050 481.050 ;
        RECT 793.950 412.950 796.050 418.050 ;
        RECT 742.950 409.950 745.050 412.050 ;
      LAYER metal2 ;
        RECT 679.950 489.450 682.050 490.050 ;
        RECT 685.950 489.450 688.050 490.050 ;
        RECT 679.950 488.400 688.050 489.450 ;
        RECT 679.950 487.950 682.050 488.400 ;
        RECT 685.950 487.950 688.050 488.400 ;
        RECT 673.950 480.450 676.050 481.050 ;
        RECT 679.950 480.450 682.050 481.050 ;
        RECT 673.950 479.400 682.050 480.450 ;
        RECT 673.950 478.950 676.050 479.400 ;
        RECT 679.950 478.950 682.050 479.400 ;
        RECT 679.950 465.450 682.050 466.050 ;
        RECT 679.950 464.400 711.450 465.450 ;
        RECT 679.950 463.950 682.050 464.400 ;
        RECT 710.400 462.450 711.450 464.400 ;
        RECT 736.950 462.450 739.050 463.050 ;
        RECT 710.400 461.400 739.050 462.450 ;
        RECT 736.950 460.950 739.050 461.400 ;
        RECT 736.950 441.450 739.050 442.200 ;
        RECT 745.950 441.450 748.050 442.050 ;
        RECT 736.950 440.400 748.050 441.450 ;
        RECT 736.950 440.100 739.050 440.400 ;
        RECT 745.950 439.950 748.050 440.400 ;
        RECT 745.950 420.450 748.050 421.050 ;
        RECT 745.950 419.400 768.450 420.450 ;
        RECT 745.950 418.950 748.050 419.400 ;
        RECT 767.400 417.450 768.450 419.400 ;
        RECT 793.950 417.450 799.050 418.050 ;
        RECT 767.400 416.400 799.050 417.450 ;
        RECT 793.950 415.950 799.050 416.400 ;
        RECT 856.950 414.450 859.050 415.050 ;
        RECT 856.950 413.400 864.450 414.450 ;
        RECT 856.950 412.950 859.050 413.400 ;
        RECT 742.950 409.950 748.050 412.050 ;
        RECT 796.950 399.450 799.050 400.050 ;
        RECT 856.950 399.450 859.050 400.050 ;
        RECT 796.950 398.400 859.050 399.450 ;
        RECT 796.950 397.950 799.050 398.400 ;
        RECT 856.950 397.950 859.050 398.400 ;
      LAYER metal3 ;
        RECT 679.950 487.950 682.050 490.050 ;
        RECT 680.400 481.050 681.600 487.950 ;
        RECT 679.950 478.950 682.050 481.050 ;
        RECT 680.400 466.050 681.600 478.950 ;
        RECT 679.950 463.950 682.050 466.050 ;
        RECT 736.950 460.950 739.050 463.050 ;
        RECT 737.400 442.200 738.600 460.950 ;
        RECT 736.950 440.100 739.050 442.200 ;
        RECT 745.950 439.950 748.050 442.050 ;
        RECT 746.400 421.050 747.600 439.950 ;
        RECT 745.950 418.950 748.050 421.050 ;
        RECT 746.400 412.050 747.600 418.950 ;
        RECT 796.950 415.950 799.050 418.050 ;
        RECT 745.950 409.950 748.050 412.050 ;
        RECT 797.400 400.050 798.600 415.950 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 857.400 400.050 858.600 412.950 ;
        RECT 796.950 397.950 799.050 400.050 ;
        RECT 856.950 397.950 859.050 400.050 ;
    END
  END ABCmd_i[1]
  PIN ABCmd_i[0]
    PORT
      LAYER metal1 ;
        RECT 652.950 478.950 655.050 481.050 ;
        RECT 604.950 454.950 607.050 457.050 ;
        RECT 637.950 454.950 640.050 457.050 ;
        RECT 814.950 423.450 817.050 427.050 ;
        RECT 853.950 424.950 856.050 427.050 ;
        RECT 812.550 423.000 817.050 423.450 ;
        RECT 812.550 422.550 816.450 423.000 ;
        RECT 812.550 418.050 813.450 422.550 ;
        RECT 854.550 421.050 855.450 424.950 ;
        RECT 853.950 418.950 856.050 421.050 ;
        RECT 811.950 415.950 814.050 418.050 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 778.950 412.950 781.200 415.050 ;
        RECT 721.950 409.950 724.050 412.050 ;
      LAYER metal2 ;
        RECT 652.950 478.950 658.050 481.050 ;
        RECT 638.100 462.450 640.200 463.050 ;
        RECT 655.950 462.450 658.050 463.050 ;
        RECT 638.100 461.400 658.050 462.450 ;
        RECT 638.100 460.950 640.200 461.400 ;
        RECT 655.950 460.950 658.050 461.400 ;
        RECT 604.950 451.950 607.050 457.050 ;
        RECT 637.950 451.950 640.050 457.050 ;
        RECT 604.950 447.450 607.050 448.050 ;
        RECT 637.800 447.450 639.900 448.050 ;
        RECT 604.950 446.400 639.900 447.450 ;
        RECT 604.950 445.950 607.050 446.400 ;
        RECT 637.800 445.950 639.900 446.400 ;
        RECT 656.100 438.450 658.200 439.050 ;
        RECT 656.100 437.400 732.450 438.450 ;
        RECT 656.100 436.950 658.200 437.400 ;
        RECT 731.400 436.050 732.450 437.400 ;
        RECT 730.950 435.450 733.050 436.050 ;
        RECT 781.950 435.450 784.050 436.050 ;
        RECT 730.950 434.400 784.050 435.450 ;
        RECT 730.950 433.950 733.050 434.400 ;
        RECT 781.950 433.950 784.050 434.400 ;
        RECT 781.950 426.450 784.050 427.050 ;
        RECT 814.950 426.450 817.050 427.050 ;
        RECT 853.950 426.450 856.050 427.050 ;
        RECT 781.950 425.400 856.050 426.450 ;
        RECT 781.950 424.950 784.050 425.400 ;
        RECT 814.950 424.950 817.050 425.400 ;
        RECT 853.950 424.950 856.050 425.400 ;
        RECT 853.950 420.450 856.050 421.050 ;
        RECT 853.950 419.400 864.450 420.450 ;
        RECT 853.950 418.950 856.050 419.400 ;
        RECT 730.950 412.950 733.050 418.050 ;
        RECT 779.100 412.950 784.050 415.050 ;
        RECT 721.950 411.450 724.050 412.050 ;
        RECT 730.800 411.450 732.900 412.050 ;
        RECT 721.950 410.400 732.900 411.450 ;
        RECT 721.950 409.950 724.050 410.400 ;
        RECT 730.800 409.950 732.900 410.400 ;
      LAYER metal3 ;
        RECT 655.950 478.950 658.050 481.050 ;
        RECT 656.400 463.050 657.600 478.950 ;
        RECT 638.100 460.950 640.200 463.050 ;
        RECT 655.950 460.950 658.050 463.050 ;
        RECT 638.400 454.050 639.600 460.950 ;
        RECT 604.950 451.950 607.050 454.050 ;
        RECT 637.950 451.950 640.050 454.050 ;
        RECT 605.400 448.050 606.600 451.950 ;
        RECT 638.400 448.050 639.600 451.950 ;
        RECT 604.950 445.950 607.050 448.050 ;
        RECT 637.800 445.950 639.900 448.050 ;
        RECT 656.400 439.050 657.600 460.950 ;
        RECT 656.100 436.950 658.200 439.050 ;
        RECT 730.950 433.950 733.050 436.050 ;
        RECT 781.950 433.950 784.050 436.050 ;
        RECT 731.400 418.050 732.600 433.950 ;
        RECT 782.400 427.050 783.600 433.950 ;
        RECT 781.950 424.950 784.050 427.050 ;
        RECT 730.950 415.950 733.050 418.050 ;
        RECT 731.400 412.050 732.600 415.950 ;
        RECT 782.400 415.050 783.600 424.950 ;
        RECT 781.950 412.950 784.050 415.050 ;
        RECT 730.800 409.950 732.900 412.050 ;
    END
  END ABCmd_i[0]
  PIN ACC_o[7]
    PORT
      LAYER metal1 ;
        RECT 556.950 49.950 559.050 52.050 ;
      LAYER metal2 ;
        RECT 553.950 49.950 559.050 52.050 ;
      LAYER metal3 ;
        RECT 553.950 51.600 558.000 52.050 ;
        RECT 553.950 49.950 558.600 51.600 ;
        RECT 557.400 -3.600 558.600 49.950 ;
    END
  END ACC_o[7]
  PIN ACC_o[6]
    PORT
      LAYER metal1 ;
        RECT 493.950 24.450 496.050 25.050 ;
        RECT 488.550 23.550 496.050 24.450 ;
        RECT 488.550 10.050 489.450 23.550 ;
        RECT 493.950 22.950 496.050 23.550 ;
        RECT 487.950 7.950 490.050 10.050 ;
      LAYER metal2 ;
        RECT 487.950 9.450 490.050 10.050 ;
        RECT 544.950 9.450 547.050 9.900 ;
        RECT 487.950 8.400 547.050 9.450 ;
        RECT 487.950 7.950 490.050 8.400 ;
        RECT 544.950 7.800 547.050 8.400 ;
      LAYER metal3 ;
        RECT 544.950 7.800 547.050 9.900 ;
        RECT 545.400 -3.600 546.600 7.800 ;
    END
  END ACC_o[6]
  PIN ACC_o[5]
    PORT
      LAYER metal1 ;
        RECT 541.950 51.450 544.050 52.050 ;
        RECT 546.000 51.450 550.050 52.050 ;
        RECT 541.950 50.550 550.050 51.450 ;
        RECT 541.950 49.950 544.050 50.550 ;
        RECT 546.000 49.950 550.050 50.550 ;
      LAYER metal2 ;
        RECT 544.950 49.950 550.050 52.050 ;
        RECT 538.950 27.450 541.050 28.050 ;
        RECT 544.950 27.450 547.050 28.050 ;
        RECT 538.950 26.400 547.050 27.450 ;
        RECT 538.950 25.950 541.050 26.400 ;
        RECT 544.950 25.950 547.050 26.400 ;
      LAYER metal3 ;
        RECT 544.950 49.950 547.050 52.050 ;
        RECT 545.400 28.050 546.600 49.950 ;
        RECT 538.950 25.950 541.050 28.050 ;
        RECT 544.950 25.950 547.050 28.050 ;
        RECT 539.400 -3.600 540.600 25.950 ;
    END
  END ACC_o[5]
  PIN ACC_o[4]
    PORT
      LAYER metal1 ;
        RECT 475.950 22.950 478.050 25.050 ;
      LAYER metal2 ;
        RECT 472.950 22.950 478.050 25.050 ;
      LAYER metal3 ;
        RECT 472.950 24.600 477.000 25.050 ;
        RECT 472.950 22.950 477.600 24.600 ;
        RECT 476.400 -3.600 477.600 22.950 ;
    END
  END ACC_o[4]
  PIN ACC_o[3]
    PORT
      LAYER metal1 ;
        RECT 409.950 22.950 412.050 25.050 ;
      LAYER metal2 ;
        RECT 407.100 22.950 412.050 25.050 ;
      LAYER metal3 ;
        RECT 407.100 22.950 409.200 25.050 ;
        RECT 407.400 -3.600 408.600 22.950 ;
    END
  END ACC_o[3]
  PIN ACC_o[2]
    PORT
      LAYER metal1 ;
        RECT 7.950 553.950 13.050 556.050 ;
      LAYER metal2 ;
        RECT -3.600 555.450 -2.550 558.450 ;
        RECT 7.950 555.450 10.050 556.050 ;
        RECT -3.600 554.400 10.050 555.450 ;
        RECT 7.950 553.950 10.050 554.400 ;
    END
  END ACC_o[2]
  PIN ACC_o[1]
    PORT
      LAYER metal1 ;
        RECT 1.950 418.950 4.050 421.050 ;
        RECT 2.550 412.050 3.450 418.950 ;
        RECT 1.950 409.950 4.050 412.050 ;
        RECT 400.950 384.450 403.050 385.050 ;
        RECT 395.550 383.550 403.050 384.450 ;
        RECT 395.550 376.050 396.450 383.550 ;
        RECT 400.950 382.950 403.050 383.550 ;
        RECT 394.950 373.950 397.050 376.050 ;
      LAYER metal2 ;
        RECT 1.950 420.450 4.050 421.050 ;
        RECT -3.600 419.400 4.050 420.450 ;
        RECT 1.950 418.950 4.050 419.400 ;
        RECT 1.950 409.950 7.050 412.050 ;
        RECT 4.950 399.450 7.050 400.050 ;
        RECT 160.950 399.450 163.050 400.050 ;
        RECT 4.950 398.400 163.050 399.450 ;
        RECT 4.950 397.950 7.050 398.400 ;
        RECT 160.950 397.950 163.050 398.400 ;
        RECT 394.950 375.450 397.050 376.050 ;
        RECT 347.400 374.400 397.050 375.450 ;
        RECT 160.950 372.450 163.050 373.050 ;
        RECT 347.400 372.450 348.450 374.400 ;
        RECT 394.950 373.950 397.050 374.400 ;
        RECT 160.950 371.400 348.450 372.450 ;
        RECT 160.950 370.950 163.050 371.400 ;
      LAYER metal3 ;
        RECT 4.950 409.950 7.050 412.050 ;
        RECT 5.400 400.050 6.600 409.950 ;
        RECT 4.950 397.950 7.050 400.050 ;
        RECT 160.950 397.950 163.050 400.050 ;
        RECT 161.400 373.050 162.600 397.950 ;
        RECT 160.950 370.950 163.050 373.050 ;
    END
  END ACC_o[1]
  PIN ACC_o[0]
    PORT
      LAYER metal1 ;
        RECT 403.950 411.450 406.050 412.050 ;
        RECT 398.550 410.550 406.050 411.450 ;
        RECT 398.550 403.050 399.450 410.550 ;
        RECT 403.950 409.950 406.050 410.550 ;
        RECT 397.950 400.950 400.050 403.050 ;
      LAYER metal2 ;
        RECT 1.950 414.450 4.050 415.050 ;
        RECT -3.600 413.400 4.050 414.450 ;
        RECT 1.950 412.950 4.050 413.400 ;
        RECT 1.950 402.450 4.050 403.050 ;
        RECT 397.950 402.450 400.050 403.050 ;
        RECT 1.950 401.400 400.050 402.450 ;
        RECT 1.950 400.950 4.050 401.400 ;
        RECT 397.950 400.950 400.050 401.400 ;
      LAYER metal3 ;
        RECT 1.950 412.950 4.050 415.050 ;
        RECT 2.400 403.050 3.600 412.950 ;
        RECT 1.950 400.950 4.050 403.050 ;
    END
  END ACC_o[0]
  PIN Done_o
    PORT
      LAYER metal1 ;
        RECT 604.950 22.950 607.050 25.050 ;
      LAYER metal2 ;
        RECT 601.950 22.950 607.050 25.050 ;
      LAYER metal3 ;
        RECT 601.950 24.600 606.000 25.050 ;
        RECT 601.950 22.950 606.600 24.600 ;
        RECT 605.400 -3.600 606.600 22.950 ;
    END
  END Done_o
  PIN LoadA_i
    PORT
      LAYER metal1 ;
        RECT 619.950 817.950 622.050 823.050 ;
        RECT 664.800 814.950 667.050 817.050 ;
        RECT 748.950 814.950 751.050 817.050 ;
      LAYER metal2 ;
        RECT 616.950 867.450 619.050 868.050 ;
        RECT 622.950 867.450 625.050 868.050 ;
        RECT 616.950 866.400 625.050 867.450 ;
        RECT 616.950 865.950 619.050 866.400 ;
        RECT 622.950 865.950 625.050 866.400 ;
        RECT 661.950 831.450 664.050 832.050 ;
        RECT 721.950 831.450 724.050 832.050 ;
        RECT 661.950 830.400 724.050 831.450 ;
        RECT 661.950 829.950 664.050 830.400 ;
        RECT 721.950 829.950 724.050 830.400 ;
        RECT 661.950 825.450 664.050 826.050 ;
        RECT 623.400 824.400 664.050 825.450 ;
        RECT 623.400 823.050 624.450 824.400 ;
        RECT 661.950 823.950 664.050 824.400 ;
        RECT 619.950 820.950 625.050 823.050 ;
        RECT 721.950 819.450 724.050 820.050 ;
        RECT 721.950 818.400 747.450 819.450 ;
        RECT 721.950 817.950 724.050 818.400 ;
        RECT 746.400 817.050 747.450 818.400 ;
        RECT 661.950 814.950 666.900 817.050 ;
        RECT 746.400 815.400 751.050 817.050 ;
        RECT 747.000 814.950 751.050 815.400 ;
      LAYER metal3 ;
        RECT 617.400 868.050 618.600 873.600 ;
        RECT 616.950 865.950 619.050 868.050 ;
        RECT 622.950 865.950 625.050 868.050 ;
        RECT 623.400 823.050 624.600 865.950 ;
        RECT 661.950 829.950 664.050 832.050 ;
        RECT 721.950 829.950 724.050 832.050 ;
        RECT 662.400 826.050 663.600 829.950 ;
        RECT 661.950 823.950 664.050 826.050 ;
        RECT 622.950 820.950 625.050 823.050 ;
        RECT 662.400 817.050 663.600 823.950 ;
        RECT 722.400 820.050 723.600 829.950 ;
        RECT 721.950 817.950 724.050 820.050 ;
        RECT 661.950 814.950 664.050 817.050 ;
    END
  END LoadA_i
  PIN LoadB_i
    PORT
      LAYER metal1 ;
        RECT 724.950 846.450 729.000 847.050 ;
        RECT 730.950 846.450 733.050 847.050 ;
        RECT 724.950 845.550 733.050 846.450 ;
        RECT 724.950 844.950 729.000 845.550 ;
        RECT 730.950 844.950 733.050 845.550 ;
        RECT 655.950 817.950 658.050 820.050 ;
        RECT 766.950 814.950 769.050 817.050 ;
        RECT 667.950 811.950 670.050 814.050 ;
      LAYER metal2 ;
        RECT 724.950 846.450 730.050 847.050 ;
        RECT 733.800 846.450 735.900 847.050 ;
        RECT 724.950 845.400 735.900 846.450 ;
        RECT 724.950 844.950 730.050 845.400 ;
        RECT 733.800 844.950 735.900 845.400 ;
        RECT 667.950 822.450 670.050 823.050 ;
        RECT 733.950 822.450 736.050 823.050 ;
        RECT 763.950 822.450 766.050 823.050 ;
        RECT 656.400 822.000 766.050 822.450 ;
        RECT 655.950 821.400 766.050 822.000 ;
        RECT 655.950 817.950 658.050 821.400 ;
        RECT 667.950 820.950 670.050 821.400 ;
        RECT 733.950 820.950 736.050 821.400 ;
        RECT 763.950 820.950 766.050 821.400 ;
        RECT 667.800 816.000 669.900 817.050 ;
        RECT 667.800 814.950 670.050 816.000 ;
        RECT 763.950 814.950 769.050 817.050 ;
        RECT 667.950 811.950 670.050 814.950 ;
      LAYER metal3 ;
        RECT 728.400 847.050 729.600 873.600 ;
        RECT 727.950 844.950 730.050 847.050 ;
        RECT 733.800 844.950 735.900 847.050 ;
        RECT 734.400 823.050 735.600 844.950 ;
        RECT 667.950 820.950 670.050 823.050 ;
        RECT 733.950 820.950 736.050 823.050 ;
        RECT 763.950 820.950 766.050 823.050 ;
        RECT 668.400 817.050 669.600 820.950 ;
        RECT 764.400 817.050 765.600 820.950 ;
        RECT 667.800 814.950 669.900 817.050 ;
        RECT 763.950 814.950 766.050 817.050 ;
    END
  END LoadB_i
  PIN LoadCmd_i
    PORT
      LAYER metal1 ;
        RECT 757.950 841.950 763.050 844.050 ;
        RECT 766.950 838.950 769.050 841.050 ;
      LAYER metal2 ;
        RECT 751.950 858.450 754.050 859.050 ;
        RECT 757.950 858.450 760.050 858.900 ;
        RECT 751.950 857.400 760.050 858.450 ;
        RECT 751.950 856.950 754.050 857.400 ;
        RECT 757.950 856.800 760.050 857.400 ;
        RECT 757.950 843.450 763.050 844.050 ;
        RECT 757.950 843.000 768.450 843.450 ;
        RECT 757.950 842.400 769.050 843.000 ;
        RECT 757.950 841.950 763.050 842.400 ;
        RECT 766.950 838.950 769.050 842.400 ;
      LAYER metal3 ;
        RECT 752.400 859.050 753.600 873.600 ;
        RECT 751.950 856.950 754.050 859.050 ;
        RECT 757.950 856.800 760.050 858.900 ;
        RECT 758.400 844.050 759.600 856.800 ;
        RECT 757.950 841.950 760.050 844.050 ;
    END
  END LoadCmd_i
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 532.950 844.950 535.050 847.050 ;
        RECT 664.950 669.450 667.050 670.050 ;
        RECT 659.550 668.550 667.050 669.450 ;
        RECT 659.550 661.050 660.450 668.550 ;
        RECT 664.950 667.950 667.050 668.550 ;
        RECT 658.950 658.950 661.050 661.050 ;
        RECT 616.950 595.950 619.050 598.050 ;
        RECT 601.800 523.950 604.050 526.050 ;
        RECT 637.950 523.950 640.050 526.050 ;
      LAYER metal2 ;
        RECT 532.950 846.450 535.050 847.050 ;
        RECT 541.950 846.450 544.050 847.050 ;
        RECT 532.950 845.400 544.050 846.450 ;
        RECT 532.950 844.950 535.050 845.400 ;
        RECT 541.950 844.950 544.050 845.400 ;
        RECT 541.950 831.450 544.050 832.050 ;
        RECT 586.950 831.450 589.050 832.050 ;
        RECT 541.950 830.400 589.050 831.450 ;
        RECT 541.950 829.950 544.050 830.400 ;
        RECT 586.950 829.950 589.050 830.400 ;
        RECT 586.950 660.450 589.050 661.050 ;
        RECT 607.950 660.450 610.050 661.050 ;
        RECT 658.950 660.450 661.050 661.050 ;
        RECT 586.950 659.400 661.050 660.450 ;
        RECT 586.950 658.950 589.050 659.400 ;
        RECT 607.950 658.950 610.050 659.400 ;
        RECT 658.950 658.950 661.050 659.400 ;
        RECT 601.950 597.450 604.050 598.050 ;
        RECT 607.950 597.450 610.050 598.050 ;
        RECT 616.950 597.450 619.050 598.050 ;
        RECT 601.950 596.400 619.050 597.450 ;
        RECT 601.950 595.950 604.050 596.400 ;
        RECT 607.950 595.950 610.050 596.400 ;
        RECT 616.950 595.950 619.050 596.400 ;
        RECT 601.800 528.450 603.900 529.050 ;
        RECT 601.800 527.400 636.450 528.450 ;
        RECT 601.800 526.950 604.050 527.400 ;
        RECT 601.950 526.050 604.050 526.950 ;
        RECT 601.800 525.000 604.050 526.050 ;
        RECT 635.400 526.050 636.450 527.400 ;
        RECT 601.800 523.950 603.900 525.000 ;
        RECT 635.400 524.400 640.050 526.050 ;
        RECT 636.000 523.950 640.050 524.400 ;
      LAYER metal3 ;
        RECT 542.400 847.050 543.600 873.600 ;
        RECT 541.950 844.950 544.050 847.050 ;
        RECT 542.400 832.050 543.600 844.950 ;
        RECT 541.950 829.950 544.050 832.050 ;
        RECT 586.950 829.950 589.050 832.050 ;
        RECT 587.400 661.050 588.600 829.950 ;
        RECT 586.950 658.950 589.050 661.050 ;
        RECT 607.950 658.950 610.050 661.050 ;
        RECT 608.400 598.050 609.600 658.950 ;
        RECT 601.950 595.950 604.050 598.050 ;
        RECT 607.950 595.950 610.050 598.050 ;
        RECT 602.400 529.050 603.600 595.950 ;
        RECT 601.800 526.950 603.900 529.050 ;
    END
  END clk
  PIN reset
    PORT
      LAYER metal1 ;
        RECT 787.800 838.950 790.050 841.050 ;
      LAYER metal2 ;
        RECT 784.950 864.450 787.050 865.050 ;
        RECT 832.950 864.450 835.050 865.050 ;
        RECT 784.950 863.400 835.050 864.450 ;
        RECT 784.950 862.950 787.050 863.400 ;
        RECT 832.950 862.950 835.050 863.400 ;
        RECT 787.800 843.000 789.900 844.050 ;
        RECT 787.800 841.950 790.050 843.000 ;
        RECT 787.950 841.050 790.050 841.950 ;
        RECT 787.800 840.000 790.050 841.050 ;
        RECT 787.800 838.950 789.900 840.000 ;
      LAYER metal3 ;
        RECT 833.400 865.050 834.600 873.600 ;
        RECT 784.950 862.950 787.050 865.050 ;
        RECT 832.950 862.950 835.050 865.050 ;
        RECT 785.400 858.600 786.600 862.950 ;
        RECT 785.400 857.400 789.600 858.600 ;
        RECT 788.400 844.050 789.600 857.400 ;
        RECT 787.800 843.000 789.900 844.050 ;
        RECT 787.800 841.950 790.050 843.000 ;
        RECT 787.950 840.000 790.050 841.950 ;
        RECT 788.400 839.400 789.600 840.000 ;
    END
  END reset
  OBS
      LAYER metal1 ;
        RECT 10.800 857.400 12.600 863.400 ;
        RECT 11.700 857.100 12.600 857.400 ;
        RECT 16.800 857.400 18.600 863.400 ;
        RECT 32.400 857.400 34.200 863.400 ;
        RECT 16.800 857.100 18.300 857.400 ;
        RECT 11.700 856.200 18.300 857.100 ;
        RECT 32.700 857.100 34.200 857.400 ;
        RECT 38.400 857.400 40.200 863.400 ;
        RECT 38.400 857.100 39.300 857.400 ;
        RECT 32.700 856.200 39.300 857.100 ;
        RECT 11.700 851.100 12.600 856.200 ;
        RECT 17.100 851.100 18.900 851.850 ;
        RECT 32.100 851.100 33.900 851.850 ;
        RECT 38.400 851.100 39.300 856.200 ;
        RECT 50.400 852.300 52.200 863.400 ;
        RECT 56.400 852.300 58.200 863.400 ;
        RECT 50.400 851.400 58.200 852.300 ;
        RECT 59.400 851.400 61.200 863.400 ;
        RECT 76.500 851.400 78.300 863.400 ;
        RECT 98.700 851.400 100.500 863.400 ;
        RECT 115.800 857.400 117.600 863.400 ;
        RECT 130.800 857.400 132.600 863.400 ;
        RECT 10.950 849.450 13.050 850.050 ;
        RECT 5.550 848.550 13.050 849.450 ;
        RECT 5.550 835.050 6.450 848.550 ;
        RECT 10.950 847.950 13.050 848.550 ;
        RECT 16.950 847.950 19.050 850.050 ;
        RECT 31.950 847.950 34.050 850.050 ;
        RECT 37.950 849.450 40.050 850.050 ;
        RECT 37.950 848.550 45.450 849.450 ;
        RECT 37.950 847.950 40.050 848.550 ;
        RECT 11.700 841.650 12.600 846.900 ;
        RECT 13.950 844.950 16.050 847.050 ;
        RECT 19.950 844.950 22.050 847.050 ;
        RECT 28.950 844.950 31.050 847.050 ;
        RECT 34.950 844.950 37.050 847.050 ;
        RECT 14.100 843.150 15.900 843.900 ;
        RECT 20.100 843.150 21.900 843.900 ;
        RECT 29.100 843.150 30.900 843.900 ;
        RECT 35.100 843.150 36.900 843.900 ;
        RECT 38.400 841.650 39.300 846.900 ;
        RECT 11.700 840.000 15.900 841.650 ;
        RECT 4.950 832.950 7.050 835.050 ;
        RECT 14.100 831.600 15.900 840.000 ;
        RECT 35.100 840.000 39.300 841.650 ;
        RECT 44.550 841.050 45.450 848.550 ;
        RECT 49.950 844.950 52.050 847.050 ;
        RECT 53.100 845.100 54.900 845.850 ;
        RECT 55.950 844.950 58.050 847.050 ;
        RECT 59.700 845.100 60.600 851.400 ;
        RECT 76.950 848.100 78.150 851.400 ;
        RECT 71.100 845.100 72.900 845.850 ;
        RECT 73.800 844.950 76.050 847.050 ;
        RECT 77.100 845.100 78.150 848.100 ;
        RECT 98.850 848.100 100.050 851.400 ;
        RECT 116.400 848.100 117.600 857.400 ;
        RECT 131.700 857.100 132.600 857.400 ;
        RECT 136.800 857.400 138.600 863.400 ;
        RECT 136.800 857.100 138.300 857.400 ;
        RECT 131.700 856.200 138.300 857.100 ;
        RECT 124.950 849.450 127.050 853.050 ;
        RECT 131.700 851.100 132.600 856.200 ;
        RECT 137.100 851.100 138.900 851.850 ;
        RECT 154.500 851.400 156.300 863.400 ;
        RECT 170.400 852.300 172.200 863.400 ;
        RECT 176.400 852.300 178.200 863.400 ;
        RECT 170.400 851.400 178.200 852.300 ;
        RECT 179.400 851.400 181.200 863.400 ;
        RECT 184.950 859.950 187.050 862.050 ;
        RECT 130.950 849.450 133.050 850.050 ;
        RECT 124.950 849.000 133.050 849.450 ;
        RECT 125.550 848.550 133.050 849.000 ;
        RECT 79.950 844.950 82.050 847.050 ;
        RECT 94.950 844.950 97.050 847.050 ;
        RECT 98.850 845.100 99.900 848.100 ;
        RECT 130.950 847.950 133.050 848.550 ;
        RECT 136.950 847.950 139.050 850.050 ;
        RECT 154.950 848.100 156.150 851.400 ;
        RECT 100.950 844.950 103.050 847.050 ;
        RECT 104.100 845.100 105.900 845.850 ;
        RECT 112.950 844.950 118.050 847.050 ;
        RECT 50.100 843.150 51.900 843.900 ;
        RECT 52.950 841.950 55.050 844.050 ;
        RECT 56.100 843.150 57.900 843.900 ;
        RECT 58.950 841.950 64.050 844.050 ;
        RECT 70.950 841.950 73.050 844.050 ;
        RECT 74.100 843.150 75.900 843.900 ;
        RECT 76.950 841.950 79.200 844.050 ;
        RECT 80.100 843.150 81.900 843.900 ;
        RECT 95.100 843.150 96.900 843.900 ;
        RECT 97.950 841.950 100.200 844.050 ;
        RECT 101.100 843.150 102.900 843.900 ;
        RECT 103.950 841.950 106.050 844.050 ;
        RECT 35.100 831.600 36.900 840.000 ;
        RECT 43.950 838.950 46.050 841.050 ;
        RECT 59.700 837.600 60.600 840.900 ;
        RECT 77.850 840.750 79.050 840.900 ;
        RECT 97.950 840.750 99.150 840.900 ;
        RECT 77.850 839.700 81.600 840.750 ;
        RECT 55.200 835.950 60.600 837.600 ;
        RECT 71.400 836.700 79.200 838.050 ;
        RECT 55.200 831.600 57.000 835.950 ;
        RECT 71.400 831.600 73.200 836.700 ;
        RECT 77.400 831.600 79.200 836.700 ;
        RECT 80.400 837.600 81.600 839.700 ;
        RECT 95.400 839.700 99.150 840.750 ;
        RECT 95.400 837.600 96.600 839.700 ;
        RECT 80.400 831.600 82.200 837.600 ;
        RECT 94.800 831.600 96.600 837.600 ;
        RECT 97.800 836.700 105.600 838.050 ;
        RECT 97.800 831.600 99.600 836.700 ;
        RECT 103.800 831.600 105.600 836.700 ;
        RECT 116.400 834.600 117.600 843.900 ;
        RECT 119.100 842.100 120.900 842.850 ;
        RECT 131.700 841.650 132.600 846.900 ;
        RECT 133.950 844.950 136.200 847.050 ;
        RECT 139.950 844.950 142.050 847.050 ;
        RECT 149.100 845.100 150.900 845.850 ;
        RECT 151.950 844.950 154.050 847.050 ;
        RECT 155.100 845.100 156.150 848.100 ;
        RECT 157.950 844.950 160.050 847.050 ;
        RECT 169.950 844.950 172.050 847.050 ;
        RECT 173.100 845.100 174.900 845.850 ;
        RECT 175.950 844.950 178.050 847.050 ;
        RECT 179.700 845.100 180.600 851.400 ;
        RECT 134.100 843.150 135.900 843.900 ;
        RECT 140.100 843.150 141.900 843.900 ;
        RECT 148.950 841.950 151.050 844.050 ;
        RECT 152.100 843.150 153.900 843.900 ;
        RECT 154.950 841.950 157.050 844.050 ;
        RECT 158.100 843.150 159.900 843.900 ;
        RECT 170.100 843.150 171.900 843.900 ;
        RECT 172.950 841.950 175.050 844.050 ;
        RECT 176.100 843.150 177.900 843.900 ;
        RECT 178.950 843.450 181.050 844.050 ;
        RECT 185.550 843.450 186.450 859.950 ;
        RECT 193.800 857.400 195.600 863.400 ;
        RECT 209.400 857.400 211.200 863.400 ;
        RECT 194.400 848.100 195.600 857.400 ;
        RECT 209.700 857.100 211.200 857.400 ;
        RECT 215.400 857.400 217.200 863.400 ;
        RECT 229.800 857.400 231.600 863.400 ;
        RECT 215.400 857.100 216.300 857.400 ;
        RECT 209.700 856.200 216.300 857.100 ;
        RECT 209.100 851.100 210.900 851.850 ;
        RECT 215.400 851.100 216.300 856.200 ;
        RECT 230.700 857.100 231.600 857.400 ;
        RECT 235.800 857.400 237.600 863.400 ;
        RECT 235.800 857.100 237.300 857.400 ;
        RECT 230.700 856.200 237.300 857.100 ;
        RECT 230.700 851.100 231.600 856.200 ;
        RECT 236.100 851.100 237.900 851.850 ;
        RECT 254.700 851.400 256.500 863.400 ;
        RECT 271.800 857.400 273.600 863.400 ;
        RECT 208.950 847.950 211.050 850.050 ;
        RECT 214.950 847.950 220.050 850.050 ;
        RECT 226.950 847.950 232.050 850.050 ;
        RECT 235.950 847.950 238.050 850.050 ;
        RECT 254.850 848.100 256.050 851.400 ;
        RECT 265.950 850.950 268.050 853.050 ;
        RECT 193.950 844.950 199.050 847.050 ;
        RECT 205.950 844.950 208.050 847.050 ;
        RECT 211.950 844.950 214.050 847.050 ;
        RECT 178.950 842.550 186.450 843.450 ;
        RECT 178.950 841.950 181.050 842.550 ;
        RECT 118.950 838.950 121.050 841.050 ;
        RECT 131.700 840.000 135.900 841.650 ;
        RECT 115.800 831.600 117.600 834.600 ;
        RECT 134.100 831.600 135.900 840.000 ;
        RECT 155.850 840.750 157.050 840.900 ;
        RECT 155.850 839.700 159.600 840.750 ;
        RECT 149.400 836.700 157.200 838.050 ;
        RECT 149.400 831.600 151.200 836.700 ;
        RECT 155.400 831.600 157.200 836.700 ;
        RECT 158.400 837.600 159.600 839.700 ;
        RECT 179.700 837.600 180.600 840.900 ;
        RECT 158.400 831.600 160.200 837.600 ;
        RECT 175.200 835.950 180.600 837.600 ;
        RECT 175.200 831.600 177.000 835.950 ;
        RECT 194.400 834.600 195.600 843.900 ;
        RECT 206.100 843.150 207.900 843.900 ;
        RECT 212.100 843.150 213.900 843.900 ;
        RECT 197.100 842.100 198.900 842.850 ;
        RECT 215.400 841.650 216.300 846.900 ;
        RECT 196.950 838.950 199.050 841.050 ;
        RECT 212.100 840.000 216.300 841.650 ;
        RECT 230.700 841.650 231.600 846.900 ;
        RECT 232.950 844.950 235.050 847.050 ;
        RECT 238.950 844.950 241.050 847.050 ;
        RECT 245.100 844.950 247.200 847.050 ;
        RECT 250.950 844.950 253.050 847.050 ;
        RECT 254.850 845.100 255.900 848.100 ;
        RECT 256.950 844.950 259.050 847.050 ;
        RECT 266.550 846.450 267.450 850.950 ;
        RECT 272.400 848.100 273.600 857.400 ;
        RECT 290.700 851.400 292.500 863.400 ;
        RECT 308.400 857.400 310.200 863.400 ;
        RECT 290.850 848.100 292.050 851.400 ;
        RECT 308.400 848.100 309.600 857.400 ;
        RECT 324.300 852.900 326.100 863.400 ;
        RECT 323.700 851.400 326.100 852.900 ;
        RECT 331.800 851.400 333.600 863.400 ;
        RECT 323.700 848.100 325.050 851.400 ;
        RECT 326.400 850.200 327.300 850.350 ;
        RECT 332.400 850.200 333.600 851.400 ;
        RECT 345.600 851.400 347.400 863.400 ;
        RECT 365.700 851.400 367.500 863.400 ;
        RECT 382.800 857.400 384.600 863.400 ;
        RECT 345.600 850.350 348.300 851.400 ;
        RECT 326.400 849.000 333.600 850.200 ;
        RECT 326.400 848.400 328.200 849.000 ;
        RECT 271.950 846.450 274.050 847.050 ;
        RECT 260.100 845.100 261.900 845.850 ;
        RECT 266.550 845.550 274.050 846.450 ;
        RECT 271.950 844.950 274.050 845.550 ;
        RECT 286.950 844.950 289.050 847.050 ;
        RECT 290.850 845.100 291.900 848.100 ;
        RECT 292.950 844.950 295.050 847.050 ;
        RECT 296.100 845.100 297.900 845.850 ;
        RECT 304.950 844.950 310.050 847.050 ;
        RECT 322.950 844.950 325.200 847.050 ;
        RECT 233.100 843.150 234.900 843.900 ;
        RECT 239.100 843.150 240.900 843.900 ;
        RECT 230.700 840.000 234.900 841.650 ;
        RECT 193.800 831.600 195.600 834.600 ;
        RECT 212.100 831.600 213.900 840.000 ;
        RECT 233.100 831.600 234.900 840.000 ;
        RECT 245.550 835.050 246.450 844.950 ;
        RECT 251.100 843.150 252.900 843.900 ;
        RECT 253.950 841.950 256.050 844.050 ;
        RECT 257.100 843.150 258.900 843.900 ;
        RECT 259.950 841.950 262.050 844.050 ;
        RECT 253.950 840.750 255.150 840.900 ;
        RECT 251.400 839.700 255.150 840.750 ;
        RECT 251.400 837.600 252.600 839.700 ;
        RECT 244.950 832.950 247.050 835.050 ;
        RECT 250.800 831.600 252.600 837.600 ;
        RECT 253.800 836.700 261.600 838.050 ;
        RECT 253.800 831.600 255.600 836.700 ;
        RECT 259.800 831.600 261.600 836.700 ;
        RECT 272.400 834.600 273.600 843.900 ;
        RECT 287.100 843.150 288.900 843.900 ;
        RECT 275.100 842.100 276.900 842.850 ;
        RECT 289.950 841.950 292.050 844.050 ;
        RECT 293.100 843.150 294.900 843.900 ;
        RECT 295.950 841.950 298.050 844.050 ;
        RECT 305.100 842.100 306.900 842.850 ;
        RECT 274.950 838.950 277.050 841.050 ;
        RECT 289.950 840.750 291.150 840.900 ;
        RECT 287.400 839.700 291.150 840.750 ;
        RECT 287.400 837.600 288.600 839.700 ;
        RECT 304.950 838.950 307.050 841.050 ;
        RECT 271.800 831.600 273.600 834.600 ;
        RECT 286.800 831.600 288.600 837.600 ;
        RECT 289.800 836.700 297.600 838.050 ;
        RECT 289.800 831.600 291.600 836.700 ;
        RECT 295.800 831.600 297.600 836.700 ;
        RECT 308.400 834.600 309.600 843.900 ;
        RECT 322.950 837.600 324.000 843.900 ;
        RECT 326.400 840.600 327.300 848.400 ;
        RECT 329.100 845.100 330.900 845.850 ;
        RECT 344.100 845.100 345.900 845.850 ;
        RECT 346.950 845.100 348.300 850.350 ;
        RECT 365.850 848.100 367.050 851.400 ;
        RECT 350.100 845.100 351.900 845.850 ;
        RECT 328.950 841.950 331.050 844.050 ;
        RECT 332.100 842.100 333.900 842.850 ;
        RECT 343.950 841.950 346.050 844.050 ;
        RECT 347.100 842.100 348.300 845.100 ;
        RECT 361.950 844.950 364.050 847.050 ;
        RECT 365.850 845.100 366.900 848.100 ;
        RECT 376.950 847.950 379.050 850.050 ;
        RECT 383.400 848.100 384.600 857.400 ;
        RECT 400.500 851.400 402.300 863.400 ;
        RECT 418.800 851.400 420.600 863.400 ;
        RECT 421.800 852.300 423.600 863.400 ;
        RECT 427.800 852.300 429.600 863.400 ;
        RECT 421.800 851.400 429.600 852.300 ;
        RECT 440.400 857.400 442.200 863.400 ;
        RECT 400.950 848.100 402.150 851.400 ;
        RECT 367.950 844.950 370.200 847.050 ;
        RECT 371.100 845.100 372.900 845.850 ;
        RECT 377.550 844.050 378.450 847.950 ;
        RECT 382.950 844.950 388.050 847.050 ;
        RECT 395.100 845.100 396.900 845.850 ;
        RECT 397.950 844.950 400.050 847.050 ;
        RECT 401.100 845.100 402.150 848.100 ;
        RECT 412.950 847.950 415.050 850.050 ;
        RECT 403.950 844.950 406.050 847.050 ;
        RECT 349.950 841.950 352.050 844.050 ;
        RECT 362.100 843.150 363.900 843.900 ;
        RECT 364.950 841.950 367.050 844.050 ;
        RECT 368.100 843.150 369.900 843.900 ;
        RECT 370.950 841.950 373.050 844.050 ;
        RECT 376.950 841.950 379.050 844.050 ;
        RECT 326.250 839.700 328.050 840.600 ;
        RECT 326.250 838.800 329.700 839.700 ;
        RECT 331.950 838.950 334.200 841.050 ;
        RECT 346.950 838.950 349.200 841.050 ;
        RECT 364.950 840.750 366.150 840.900 ;
        RECT 362.400 839.700 366.150 840.750 ;
        RECT 308.400 831.600 310.200 834.600 ;
        RECT 322.800 831.600 324.600 837.600 ;
        RECT 328.800 834.600 329.700 838.800 ;
        RECT 347.400 834.600 348.600 837.900 ;
        RECT 362.400 837.600 363.600 839.700 ;
        RECT 328.800 831.600 330.600 834.600 ;
        RECT 346.800 831.600 348.600 834.600 ;
        RECT 361.800 831.600 363.600 837.600 ;
        RECT 364.800 836.700 372.600 838.050 ;
        RECT 364.800 831.600 366.600 836.700 ;
        RECT 370.800 831.600 372.600 836.700 ;
        RECT 383.400 834.600 384.600 843.900 ;
        RECT 386.100 842.100 387.900 842.850 ;
        RECT 394.950 841.950 397.050 844.050 ;
        RECT 398.100 843.150 399.900 843.900 ;
        RECT 400.950 841.950 403.050 844.050 ;
        RECT 404.100 843.150 405.900 843.900 ;
        RECT 413.550 843.450 414.450 847.950 ;
        RECT 419.400 845.100 420.300 851.400 ;
        RECT 436.950 847.950 439.050 850.050 ;
        RECT 440.400 848.100 441.600 857.400 ;
        RECT 455.400 851.400 457.200 863.400 ;
        RECT 462.900 852.900 464.700 863.400 ;
        RECT 478.800 857.400 480.600 863.400 ;
        RECT 479.700 857.100 480.600 857.400 ;
        RECT 484.800 857.400 486.600 863.400 ;
        RECT 499.800 857.400 501.600 863.400 ;
        RECT 517.800 857.400 519.600 863.400 ;
        RECT 484.800 857.100 486.300 857.400 ;
        RECT 479.700 856.200 486.300 857.100 ;
        RECT 462.900 851.400 465.300 852.900 ;
        RECT 455.400 850.200 456.600 851.400 ;
        RECT 461.700 850.200 462.600 850.350 ;
        RECT 442.950 847.950 445.050 850.050 ;
        RECT 448.950 847.950 451.050 850.050 ;
        RECT 455.400 849.000 462.600 850.200 ;
        RECT 460.800 848.400 462.600 849.000 ;
        RECT 421.950 844.950 424.050 847.050 ;
        RECT 425.100 845.100 426.900 845.850 ;
        RECT 427.950 844.950 430.050 847.050 ;
        RECT 437.100 846.150 438.900 846.900 ;
        RECT 439.950 844.950 442.050 847.050 ;
        RECT 443.100 846.150 444.900 846.900 ;
        RECT 418.950 843.450 421.050 844.050 ;
        RECT 413.550 842.550 421.050 843.450 ;
        RECT 422.100 843.150 423.900 843.900 ;
        RECT 418.950 841.950 421.050 842.550 ;
        RECT 424.950 841.950 427.050 844.050 ;
        RECT 428.100 843.150 429.900 843.900 ;
        RECT 385.950 838.950 388.050 841.050 ;
        RECT 401.850 840.750 403.050 840.900 ;
        RECT 401.850 839.700 405.600 840.750 ;
        RECT 382.800 831.600 384.600 834.600 ;
        RECT 395.400 836.700 403.200 838.050 ;
        RECT 395.400 831.600 397.200 836.700 ;
        RECT 401.400 831.600 403.200 836.700 ;
        RECT 404.400 837.600 405.600 839.700 ;
        RECT 419.400 837.600 420.300 840.900 ;
        RECT 440.400 839.700 441.600 843.900 ;
        RECT 440.400 838.800 444.000 839.700 ;
        RECT 404.400 831.600 406.200 837.600 ;
        RECT 419.400 835.950 424.800 837.600 ;
        RECT 423.000 831.600 424.800 835.950 ;
        RECT 442.200 831.600 444.000 838.800 ;
        RECT 449.550 838.050 450.450 847.950 ;
        RECT 458.100 845.100 459.900 845.850 ;
        RECT 455.100 842.100 456.900 842.850 ;
        RECT 457.950 841.950 460.050 844.050 ;
        RECT 454.950 838.950 457.050 841.050 ;
        RECT 461.700 840.600 462.600 848.400 ;
        RECT 463.950 848.100 465.300 851.400 ;
        RECT 479.700 851.100 480.600 856.200 ;
        RECT 485.100 851.100 486.900 851.850 ;
        RECT 478.950 849.450 481.050 850.050 ;
        RECT 473.550 848.550 481.050 849.450 ;
        RECT 463.950 844.950 469.050 847.050 ;
        RECT 460.950 839.700 462.750 840.600 ;
        RECT 459.300 838.800 462.750 839.700 ;
        RECT 448.950 835.950 451.050 838.050 ;
        RECT 459.300 834.600 460.200 838.800 ;
        RECT 465.000 837.600 466.050 843.900 ;
        RECT 473.550 841.050 474.450 848.550 ;
        RECT 478.950 847.950 481.050 848.550 ;
        RECT 484.950 847.950 487.050 850.050 ;
        RECT 500.400 848.100 501.600 857.400 ;
        RECT 514.950 847.950 517.050 850.050 ;
        RECT 518.400 848.100 519.600 857.400 ;
        RECT 533.400 850.500 535.200 863.400 ;
        RECT 539.400 850.500 541.200 863.400 ;
        RECT 545.400 850.500 547.200 863.400 ;
        RECT 551.400 850.500 553.200 863.400 ;
        RECT 565.200 857.400 567.000 863.400 ;
        RECT 559.950 850.950 562.050 853.050 ;
        RECT 520.950 847.950 523.050 850.050 ;
        RECT 526.950 847.950 529.050 850.050 ;
        RECT 533.400 849.300 537.300 850.500 ;
        RECT 539.400 849.300 543.300 850.500 ;
        RECT 545.400 849.300 549.300 850.500 ;
        RECT 551.400 849.300 554.100 850.500 ;
        RECT 479.700 841.650 480.600 846.900 ;
        RECT 481.950 844.950 484.050 847.050 ;
        RECT 487.950 844.950 490.050 847.050 ;
        RECT 496.950 844.950 502.050 847.050 ;
        RECT 515.100 846.150 516.900 846.900 ;
        RECT 517.950 844.950 520.050 847.050 ;
        RECT 521.100 846.150 522.900 846.900 ;
        RECT 482.100 843.150 483.900 843.900 ;
        RECT 488.100 843.150 489.900 843.900 ;
        RECT 472.950 838.950 475.050 841.050 ;
        RECT 479.700 840.000 483.900 841.650 ;
        RECT 458.400 831.600 460.200 834.600 ;
        RECT 464.400 831.600 466.200 837.600 ;
        RECT 482.100 831.600 483.900 840.000 ;
        RECT 500.400 834.600 501.600 843.900 ;
        RECT 503.100 842.100 504.900 842.850 ;
        RECT 502.950 838.950 505.050 841.050 ;
        RECT 518.400 839.700 519.600 843.900 ;
        RECT 499.800 831.600 501.600 834.600 ;
        RECT 516.000 838.800 519.600 839.700 ;
        RECT 516.000 831.600 517.800 838.800 ;
        RECT 527.550 835.050 528.450 847.950 ;
        RECT 533.100 843.150 534.900 843.900 ;
        RECT 536.100 841.800 537.300 849.300 ;
        RECT 538.500 841.800 540.300 842.400 ;
        RECT 536.100 840.600 540.300 841.800 ;
        RECT 542.100 841.800 543.300 849.300 ;
        RECT 544.500 841.800 546.300 842.400 ;
        RECT 542.100 840.600 546.300 841.800 ;
        RECT 548.100 841.800 549.300 849.300 ;
        RECT 553.200 848.100 554.100 849.300 ;
        RECT 553.950 846.450 556.050 847.050 ;
        RECT 560.550 846.450 561.450 850.950 ;
        RECT 565.500 847.050 567.000 857.400 ;
        RECT 571.800 857.400 573.600 863.400 ;
        RECT 571.800 852.750 573.000 857.400 ;
        RECT 577.800 856.500 579.600 863.400 ;
        RECT 584.400 860.400 586.200 863.400 ;
        RECT 587.400 860.400 589.200 863.400 ;
        RECT 590.400 860.400 592.200 863.400 ;
        RECT 584.850 859.200 586.050 860.400 ;
        RECT 583.950 857.100 586.050 859.200 ;
        RECT 587.400 857.400 589.050 860.400 ;
        RECT 590.850 857.400 592.050 860.400 ;
        RECT 594.000 857.400 595.800 863.400 ;
        RECT 600.000 857.400 601.800 863.400 ;
        RECT 606.900 860.400 608.850 863.400 ;
        RECT 609.900 860.400 612.000 863.400 ;
        RECT 612.900 860.400 615.150 863.400 ;
        RECT 607.650 859.050 608.850 860.400 ;
        RECT 610.950 859.050 612.000 860.400 ;
        RECT 614.250 859.050 615.150 860.400 ;
        RECT 573.900 855.300 579.600 856.500 ;
        RECT 580.500 856.050 582.300 856.500 ;
        RECT 586.950 856.050 589.050 857.400 ;
        RECT 573.900 854.700 575.700 855.300 ;
        RECT 580.500 854.850 589.050 856.050 ;
        RECT 589.950 855.300 592.050 857.400 ;
        RECT 593.850 855.150 595.950 857.400 ;
        RECT 600.000 856.500 601.050 857.400 ;
        RECT 607.650 856.950 610.050 859.050 ;
        RECT 610.950 856.950 613.050 859.050 ;
        RECT 613.950 856.950 616.050 859.050 ;
        RECT 580.500 854.700 582.300 854.850 ;
        RECT 593.100 853.350 595.950 855.150 ;
        RECT 598.950 854.400 601.050 856.500 ;
        RECT 619.500 854.700 621.300 863.400 ;
        RECT 625.500 857.400 627.300 863.400 ;
        RECT 643.800 857.400 645.600 863.400 ;
        RECT 655.200 857.400 657.000 863.400 ;
        RECT 626.250 856.500 627.300 857.400 ;
        RECT 626.250 855.600 630.300 856.500 ;
        RECT 608.100 853.650 625.800 854.700 ;
        RECT 583.950 852.750 586.050 853.350 ;
        RECT 569.100 851.850 586.050 852.750 ;
        RECT 553.950 845.550 561.450 846.450 ;
        RECT 553.950 844.950 556.050 845.550 ;
        RECT 565.050 844.950 567.150 847.050 ;
        RECT 550.500 841.800 552.300 842.400 ;
        RECT 548.100 840.600 552.300 841.800 ;
        RECT 536.100 839.700 537.300 840.600 ;
        RECT 542.100 839.700 543.300 840.600 ;
        RECT 548.100 839.700 549.300 840.600 ;
        RECT 553.200 839.700 554.100 843.900 ;
        RECT 533.400 838.500 537.300 839.700 ;
        RECT 539.400 838.500 543.300 839.700 ;
        RECT 545.400 838.500 549.300 839.700 ;
        RECT 551.400 838.500 554.100 839.700 ;
        RECT 526.950 832.950 529.050 835.050 ;
        RECT 533.400 831.600 535.200 838.500 ;
        RECT 539.400 831.600 541.200 838.500 ;
        RECT 545.400 831.600 547.200 838.500 ;
        RECT 551.400 831.600 553.200 838.500 ;
        RECT 565.500 834.600 567.000 844.950 ;
        RECT 565.200 831.600 567.000 834.600 ;
        RECT 569.100 837.600 570.000 851.850 ;
        RECT 583.950 851.250 586.050 851.850 ;
        RECT 589.950 852.300 592.050 853.350 ;
        RECT 608.100 852.300 610.050 853.650 ;
        RECT 624.000 852.900 625.800 853.650 ;
        RECT 589.950 851.250 610.050 852.300 ;
        RECT 610.950 852.150 613.050 852.750 ;
        RECT 610.950 850.950 622.500 852.150 ;
        RECT 570.900 850.350 572.700 850.950 ;
        RECT 610.950 850.650 613.050 850.950 ;
        RECT 620.700 850.350 622.500 850.950 ;
        RECT 570.900 849.450 610.050 850.350 ;
        RECT 570.900 849.150 622.050 849.450 ;
        RECT 608.100 848.550 622.050 849.150 ;
        RECT 572.850 845.100 574.950 847.050 ;
        RECT 578.100 846.000 585.150 847.800 ;
        RECT 598.950 847.650 601.050 848.250 ;
        RECT 572.850 844.050 583.200 845.100 ;
        RECT 570.900 842.700 572.700 843.000 ;
        RECT 575.700 842.700 577.500 843.000 ;
        RECT 570.900 841.200 578.700 842.700 ;
        RECT 582.150 842.250 583.200 844.050 ;
        RECT 584.250 844.350 585.150 846.000 ;
        RECT 586.500 847.500 601.050 847.650 ;
        RECT 607.800 847.500 609.600 847.650 ;
        RECT 586.500 846.450 609.600 847.500 ;
        RECT 618.150 847.350 622.050 848.550 ;
        RECT 586.500 845.250 588.300 846.450 ;
        RECT 598.950 846.150 601.050 846.450 ;
        RECT 607.800 845.850 609.600 846.450 ;
        RECT 610.500 846.450 617.250 847.350 ;
        RECT 619.950 847.050 622.050 847.350 ;
        RECT 594.750 845.250 596.850 845.550 ;
        RECT 584.250 843.300 593.850 844.350 ;
        RECT 594.750 843.450 598.650 845.250 ;
        RECT 610.500 844.950 611.550 846.450 ;
        RECT 599.550 844.050 611.550 844.950 ;
        RECT 592.950 842.550 593.850 843.300 ;
        RECT 599.550 842.550 600.600 844.050 ;
        RECT 612.450 843.750 614.250 845.550 ;
        RECT 616.050 844.050 617.250 846.450 ;
        RECT 625.950 845.850 628.050 847.950 ;
        RECT 626.100 844.050 627.900 845.850 ;
        RECT 582.150 841.200 592.050 842.250 ;
        RECT 592.950 841.200 600.600 842.550 ;
        RECT 601.950 841.350 605.850 843.150 ;
        RECT 577.200 837.600 578.700 841.200 ;
        RECT 591.000 840.300 592.050 841.200 ;
        RECT 601.950 841.050 604.050 841.350 ;
        RECT 609.150 840.300 610.950 840.750 ;
        RECT 612.450 840.300 613.500 843.750 ;
        RECT 616.050 843.000 627.900 844.050 ;
        RECT 629.100 842.100 630.300 855.600 ;
        RECT 640.800 847.950 643.050 850.050 ;
        RECT 644.400 848.100 645.600 857.400 ;
        RECT 646.950 847.950 649.050 850.050 ;
        RECT 655.500 847.050 657.000 857.400 ;
        RECT 661.800 857.400 663.600 863.400 ;
        RECT 661.800 852.750 663.000 857.400 ;
        RECT 667.800 856.500 669.600 863.400 ;
        RECT 674.400 860.400 676.200 863.400 ;
        RECT 677.400 860.400 679.200 863.400 ;
        RECT 680.400 860.400 682.200 863.400 ;
        RECT 674.850 859.200 676.050 860.400 ;
        RECT 673.950 857.100 676.050 859.200 ;
        RECT 677.400 857.400 679.050 860.400 ;
        RECT 680.850 857.400 682.050 860.400 ;
        RECT 684.000 857.400 685.800 863.400 ;
        RECT 690.000 857.400 691.800 863.400 ;
        RECT 696.900 860.400 698.850 863.400 ;
        RECT 699.900 860.400 702.000 863.400 ;
        RECT 702.900 860.400 705.150 863.400 ;
        RECT 697.650 859.050 698.850 860.400 ;
        RECT 700.950 859.050 702.000 860.400 ;
        RECT 704.250 859.050 705.150 860.400 ;
        RECT 663.900 855.300 669.600 856.500 ;
        RECT 670.500 856.050 672.300 856.500 ;
        RECT 676.950 856.050 679.050 857.400 ;
        RECT 663.900 854.700 665.700 855.300 ;
        RECT 670.500 854.850 679.050 856.050 ;
        RECT 679.950 855.300 682.050 857.400 ;
        RECT 683.850 855.150 685.950 857.400 ;
        RECT 690.000 856.500 691.050 857.400 ;
        RECT 697.650 856.950 700.050 859.050 ;
        RECT 700.950 856.950 703.050 859.050 ;
        RECT 703.950 856.950 706.050 859.050 ;
        RECT 670.500 854.700 672.300 854.850 ;
        RECT 683.100 853.350 685.950 855.150 ;
        RECT 688.950 854.400 691.050 856.500 ;
        RECT 709.500 854.700 711.300 863.400 ;
        RECT 715.500 857.400 717.300 863.400 ;
        RECT 716.250 856.500 717.300 857.400 ;
        RECT 716.250 855.600 720.300 856.500 ;
        RECT 698.100 853.650 715.800 854.700 ;
        RECT 673.950 852.750 676.050 853.350 ;
        RECT 659.100 851.850 676.050 852.750 ;
        RECT 641.100 846.150 642.900 846.900 ;
        RECT 643.950 844.950 646.050 847.050 ;
        RECT 647.100 846.150 648.900 846.900 ;
        RECT 655.050 844.950 657.150 847.050 ;
        RECT 583.500 838.500 590.100 840.300 ;
        RECT 591.000 838.500 597.900 840.300 ;
        RECT 609.150 839.850 613.500 840.300 ;
        RECT 605.850 839.100 613.500 839.850 ;
        RECT 615.000 841.200 630.300 842.100 ;
        RECT 605.850 838.950 610.950 839.100 ;
        RECT 605.850 837.600 606.750 838.950 ;
        RECT 615.000 838.050 616.050 841.200 ;
        RECT 624.300 839.700 626.100 840.300 ;
        RECT 569.100 831.600 570.900 837.600 ;
        RECT 577.200 836.400 581.400 837.600 ;
        RECT 579.600 831.600 581.400 836.400 ;
        RECT 583.950 835.500 586.050 837.600 ;
        RECT 586.950 835.500 589.050 837.600 ;
        RECT 589.950 835.500 592.050 837.600 ;
        RECT 593.850 835.500 595.950 837.600 ;
        RECT 598.950 835.500 601.050 837.600 ;
        RECT 602.700 836.250 606.750 837.600 ;
        RECT 602.700 835.800 604.500 836.250 ;
        RECT 607.950 835.950 610.050 838.050 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 613.950 835.950 616.050 838.050 ;
        RECT 617.700 838.500 626.100 839.700 ;
        RECT 617.700 837.600 619.200 838.500 ;
        RECT 629.100 837.600 630.300 841.200 ;
        RECT 644.400 839.700 645.600 843.900 ;
        RECT 584.400 834.600 585.750 835.500 ;
        RECT 587.400 834.600 589.050 835.500 ;
        RECT 590.400 834.600 592.050 835.500 ;
        RECT 594.000 834.600 595.650 835.500 ;
        RECT 600.000 834.600 601.050 835.500 ;
        RECT 607.950 834.600 609.300 835.950 ;
        RECT 610.950 834.600 612.300 835.950 ;
        RECT 613.950 834.600 615.300 835.950 ;
        RECT 584.400 831.600 586.200 834.600 ;
        RECT 587.400 831.600 589.200 834.600 ;
        RECT 590.400 831.600 592.200 834.600 ;
        RECT 594.000 831.600 595.800 834.600 ;
        RECT 600.000 831.600 601.800 834.600 ;
        RECT 607.500 831.600 609.300 834.600 ;
        RECT 610.500 831.600 612.300 834.600 ;
        RECT 613.500 831.600 615.300 834.600 ;
        RECT 617.700 831.600 619.500 837.600 ;
        RECT 628.500 831.600 630.300 837.600 ;
        RECT 642.000 838.800 645.600 839.700 ;
        RECT 642.000 831.600 643.800 838.800 ;
        RECT 655.500 834.600 657.000 844.950 ;
        RECT 655.200 831.600 657.000 834.600 ;
        RECT 659.100 837.600 660.000 851.850 ;
        RECT 673.950 851.250 676.050 851.850 ;
        RECT 679.950 852.300 682.050 853.350 ;
        RECT 698.100 852.300 700.050 853.650 ;
        RECT 714.000 852.900 715.800 853.650 ;
        RECT 679.950 851.250 700.050 852.300 ;
        RECT 700.950 852.150 703.050 852.750 ;
        RECT 700.950 850.950 712.500 852.150 ;
        RECT 660.900 850.350 662.700 850.950 ;
        RECT 700.950 850.650 703.050 850.950 ;
        RECT 710.700 850.350 712.500 850.950 ;
        RECT 660.900 849.450 700.050 850.350 ;
        RECT 660.900 849.150 712.050 849.450 ;
        RECT 698.100 848.550 712.050 849.150 ;
        RECT 662.850 845.100 664.950 847.050 ;
        RECT 668.100 846.000 675.150 847.800 ;
        RECT 688.950 847.650 691.050 848.250 ;
        RECT 662.850 844.050 673.200 845.100 ;
        RECT 660.900 842.700 662.700 843.000 ;
        RECT 665.700 842.700 667.500 843.000 ;
        RECT 660.900 841.200 668.700 842.700 ;
        RECT 672.150 842.250 673.200 844.050 ;
        RECT 674.250 844.350 675.150 846.000 ;
        RECT 676.500 847.500 691.050 847.650 ;
        RECT 697.800 847.500 699.600 847.650 ;
        RECT 676.500 846.450 699.600 847.500 ;
        RECT 708.150 847.350 712.050 848.550 ;
        RECT 676.500 845.250 678.300 846.450 ;
        RECT 688.950 846.150 691.050 846.450 ;
        RECT 697.800 845.850 699.600 846.450 ;
        RECT 700.500 846.450 707.250 847.350 ;
        RECT 709.950 847.050 712.050 847.350 ;
        RECT 684.750 845.250 686.850 845.550 ;
        RECT 674.250 843.300 683.850 844.350 ;
        RECT 684.750 843.450 688.650 845.250 ;
        RECT 700.500 844.950 701.550 846.450 ;
        RECT 689.550 844.050 701.550 844.950 ;
        RECT 682.950 842.550 683.850 843.300 ;
        RECT 689.550 842.550 690.600 844.050 ;
        RECT 702.450 843.750 704.250 845.550 ;
        RECT 706.050 844.050 707.250 846.450 ;
        RECT 715.950 845.850 718.050 847.950 ;
        RECT 716.100 844.050 717.900 845.850 ;
        RECT 672.150 841.200 682.050 842.250 ;
        RECT 682.950 841.200 690.600 842.550 ;
        RECT 691.950 841.350 695.850 843.150 ;
        RECT 667.200 837.600 668.700 841.200 ;
        RECT 681.000 840.300 682.050 841.200 ;
        RECT 691.950 841.050 694.050 841.350 ;
        RECT 699.150 840.300 700.950 840.750 ;
        RECT 702.450 840.300 703.500 843.750 ;
        RECT 706.050 843.000 717.900 844.050 ;
        RECT 719.100 842.100 720.300 855.600 ;
        RECT 734.700 851.400 736.500 863.400 ;
        RECT 753.600 851.400 755.400 863.400 ;
        RECT 770.400 857.400 772.200 863.400 ;
        RECT 784.800 857.400 786.600 863.400 ;
        RECT 734.850 848.100 736.050 851.400 ;
        RECT 753.600 850.350 756.300 851.400 ;
        RECT 734.850 845.100 735.900 848.100 ;
        RECT 736.800 844.950 739.050 847.050 ;
        RECT 740.100 845.100 741.900 845.850 ;
        RECT 752.100 845.100 753.900 845.850 ;
        RECT 754.950 845.100 756.300 850.350 ;
        RECT 770.400 848.100 771.600 857.400 ;
        RECT 785.400 848.100 786.600 857.400 ;
        RECT 791.550 851.400 793.350 863.400 ;
        RECT 799.050 857.400 800.850 863.400 ;
        RECT 796.950 855.300 800.850 857.400 ;
        RECT 806.850 856.500 808.650 863.400 ;
        RECT 814.650 857.400 816.450 863.400 ;
        RECT 815.250 856.500 816.450 857.400 ;
        RECT 805.950 855.450 812.550 856.500 ;
        RECT 805.950 854.700 807.750 855.450 ;
        RECT 810.750 854.700 812.550 855.450 ;
        RECT 815.250 854.400 820.050 856.500 ;
        RECT 798.150 852.600 800.850 854.400 ;
        RECT 801.750 853.800 803.550 854.400 ;
        RECT 801.750 852.900 808.050 853.800 ;
        RECT 815.250 853.500 816.450 854.400 ;
        RECT 801.750 852.600 803.550 852.900 ;
        RECT 799.950 851.700 800.850 852.600 ;
        RECT 769.950 846.450 772.050 847.050 ;
        RECT 774.000 846.450 778.050 847.050 ;
        RECT 758.100 845.100 759.900 845.850 ;
        RECT 769.950 845.550 778.050 846.450 ;
        RECT 731.100 843.150 732.900 843.900 ;
        RECT 673.500 838.500 680.100 840.300 ;
        RECT 681.000 838.500 687.900 840.300 ;
        RECT 699.150 839.850 703.500 840.300 ;
        RECT 695.850 839.100 703.500 839.850 ;
        RECT 705.000 841.200 720.300 842.100 ;
        RECT 733.950 841.950 736.050 844.050 ;
        RECT 737.100 843.150 738.900 843.900 ;
        RECT 739.950 841.950 742.050 844.050 ;
        RECT 751.950 841.950 754.050 844.050 ;
        RECT 755.100 842.100 756.300 845.100 ;
        RECT 769.950 844.950 772.050 845.550 ;
        RECT 774.000 844.950 778.050 845.550 ;
        RECT 784.950 844.950 787.050 847.050 ;
        RECT 791.550 844.050 792.750 851.400 ;
        RECT 796.950 850.800 799.050 851.700 ;
        RECT 799.950 850.800 805.950 851.700 ;
        RECT 794.850 849.600 799.050 850.800 ;
        RECT 793.950 847.800 795.750 849.600 ;
        RECT 805.050 845.100 805.950 850.800 ;
        RECT 807.150 850.800 808.050 852.900 ;
        RECT 808.950 852.300 816.450 853.500 ;
        RECT 808.950 851.700 810.750 852.300 ;
        RECT 823.050 851.400 824.850 863.400 ;
        RECT 813.750 850.800 824.850 851.400 ;
        RECT 807.150 850.200 824.850 850.800 ;
        RECT 807.150 849.900 815.550 850.200 ;
        RECT 813.750 849.600 815.550 849.900 ;
        RECT 818.100 844.800 819.900 845.100 ;
        RECT 767.100 842.100 768.900 842.850 ;
        RECT 695.850 838.950 700.950 839.100 ;
        RECT 695.850 837.600 696.750 838.950 ;
        RECT 705.000 838.050 706.050 841.200 ;
        RECT 714.300 839.700 716.100 840.300 ;
        RECT 659.100 831.600 660.900 837.600 ;
        RECT 667.200 836.400 671.400 837.600 ;
        RECT 669.600 831.600 671.400 836.400 ;
        RECT 673.950 835.500 676.050 837.600 ;
        RECT 676.950 835.500 679.050 837.600 ;
        RECT 679.950 835.500 682.050 837.600 ;
        RECT 683.850 835.500 685.950 837.600 ;
        RECT 688.950 835.500 691.050 837.600 ;
        RECT 692.700 836.250 696.750 837.600 ;
        RECT 692.700 835.800 694.500 836.250 ;
        RECT 697.950 835.950 700.050 838.050 ;
        RECT 700.950 835.950 703.050 838.050 ;
        RECT 703.950 835.950 706.050 838.050 ;
        RECT 707.700 838.500 716.100 839.700 ;
        RECT 707.700 837.600 709.200 838.500 ;
        RECT 719.100 837.600 720.300 841.200 ;
        RECT 733.950 840.750 735.150 840.900 ;
        RECT 731.400 839.700 735.150 840.750 ;
        RECT 731.400 837.600 732.600 839.700 ;
        RECT 754.950 838.950 757.050 841.050 ;
        RECT 674.400 834.600 675.750 835.500 ;
        RECT 677.400 834.600 679.050 835.500 ;
        RECT 680.400 834.600 682.050 835.500 ;
        RECT 684.000 834.600 685.650 835.500 ;
        RECT 690.000 834.600 691.050 835.500 ;
        RECT 697.950 834.600 699.300 835.950 ;
        RECT 700.950 834.600 702.300 835.950 ;
        RECT 703.950 834.600 705.300 835.950 ;
        RECT 674.400 831.600 676.200 834.600 ;
        RECT 677.400 831.600 679.200 834.600 ;
        RECT 680.400 831.600 682.200 834.600 ;
        RECT 684.000 831.600 685.800 834.600 ;
        RECT 690.000 831.600 691.800 834.600 ;
        RECT 697.500 831.600 699.300 834.600 ;
        RECT 700.500 831.600 702.300 834.600 ;
        RECT 703.500 831.600 705.300 834.600 ;
        RECT 707.700 831.600 709.500 837.600 ;
        RECT 718.500 831.600 720.300 837.600 ;
        RECT 730.800 831.600 732.600 837.600 ;
        RECT 733.800 836.700 741.600 838.050 ;
        RECT 733.800 831.600 735.600 836.700 ;
        RECT 739.800 831.600 741.600 836.700 ;
        RECT 755.400 834.600 756.600 837.900 ;
        RECT 754.800 831.600 756.600 834.600 ;
        RECT 770.400 834.600 771.600 843.900 ;
        RECT 785.400 834.600 786.600 843.900 ;
        RECT 788.100 842.100 789.900 842.850 ;
        RECT 770.400 831.600 772.200 834.600 ;
        RECT 784.800 831.600 786.600 834.600 ;
        RECT 791.550 841.950 792.900 844.050 ;
        RECT 793.950 841.950 796.050 844.050 ;
        RECT 797.100 841.950 797.850 843.750 ;
        RECT 805.800 841.950 808.050 844.050 ;
        RECT 811.950 841.950 814.050 844.050 ;
        RECT 815.100 843.900 819.900 844.800 ;
        RECT 818.100 843.300 819.900 843.900 ;
        RECT 821.100 843.150 822.900 844.950 ;
        RECT 815.100 842.400 816.900 843.000 ;
        RECT 821.100 842.400 822.000 843.150 ;
        RECT 791.550 837.600 792.750 841.950 ;
        RECT 815.100 841.200 822.000 842.400 ;
        RECT 805.050 840.000 805.950 840.900 ;
        RECT 815.100 840.000 816.150 841.200 ;
        RECT 805.050 839.100 816.150 840.000 ;
        RECT 805.050 838.800 805.950 839.100 ;
        RECT 791.550 831.600 793.350 837.600 ;
        RECT 796.950 836.700 799.050 837.600 ;
        RECT 804.150 837.000 805.950 838.800 ;
        RECT 815.100 838.200 816.150 839.100 ;
        RECT 811.350 837.450 813.150 838.200 ;
        RECT 796.950 835.500 800.700 836.700 ;
        RECT 799.650 834.600 800.700 835.500 ;
        RECT 808.200 836.400 813.150 837.450 ;
        RECT 814.650 836.400 816.450 838.200 ;
        RECT 823.950 837.600 824.850 850.200 ;
        RECT 836.400 851.400 838.200 863.400 ;
        RECT 836.400 845.100 837.600 851.400 ;
        RECT 833.100 843.150 834.900 843.900 ;
        RECT 835.950 841.950 838.050 844.050 ;
        RECT 808.200 834.600 809.250 836.400 ;
        RECT 817.950 835.500 820.050 837.600 ;
        RECT 817.950 834.600 819.000 835.500 ;
        RECT 799.650 831.600 801.450 834.600 ;
        RECT 807.450 831.600 809.250 834.600 ;
        RECT 815.250 833.700 819.000 834.600 ;
        RECT 815.250 831.600 817.050 833.700 ;
        RECT 823.050 831.600 824.850 837.600 ;
        RECT 836.400 837.600 837.600 840.900 ;
        RECT 836.400 831.600 838.200 837.600 ;
        RECT 15.000 823.050 16.800 827.400 ;
        RECT 11.400 821.400 16.800 823.050 ;
        RECT 11.400 818.100 12.300 821.400 ;
        RECT 35.100 819.000 36.900 827.400 ;
        RECT 52.800 821.400 54.600 827.400 ;
        RECT 32.700 817.350 36.900 819.000 ;
        RECT 53.400 819.300 54.600 821.400 ;
        RECT 55.800 822.300 57.600 827.400 ;
        RECT 61.800 822.300 63.600 827.400 ;
        RECT 55.800 820.950 63.600 822.300 ;
        RECT 67.950 820.950 70.050 823.050 ;
        RECT 73.800 821.400 75.600 827.400 ;
        RECT 53.400 818.250 57.150 819.300 ;
        RECT 55.950 818.100 57.150 818.250 ;
        RECT 4.950 816.450 9.000 817.050 ;
        RECT 10.950 816.450 13.050 817.050 ;
        RECT 4.950 815.550 13.050 816.450 ;
        RECT 4.950 814.950 9.000 815.550 ;
        RECT 10.950 814.950 13.050 815.550 ;
        RECT 14.100 815.100 15.900 815.850 ;
        RECT 16.950 814.950 19.050 817.050 ;
        RECT 20.100 815.100 21.900 815.850 ;
        RECT 11.400 807.600 12.300 813.900 ;
        RECT 13.950 811.950 16.050 814.050 ;
        RECT 17.100 813.150 18.900 813.900 ;
        RECT 19.950 811.950 22.050 814.050 ;
        RECT 32.700 812.100 33.600 817.350 ;
        RECT 35.100 815.100 36.900 815.850 ;
        RECT 41.100 815.100 42.900 815.850 ;
        RECT 46.950 814.950 49.050 817.050 ;
        RECT 53.100 815.100 54.900 815.850 ;
        RECT 55.950 814.950 58.050 817.050 ;
        RECT 59.100 815.100 60.900 815.850 ;
        RECT 61.950 814.950 64.050 817.050 ;
        RECT 34.950 811.950 37.050 814.050 ;
        RECT 40.950 811.950 43.050 814.050 ;
        RECT 47.550 811.050 48.450 814.950 ;
        RECT 68.550 814.050 69.450 820.950 ;
        RECT 74.400 819.300 75.600 821.400 ;
        RECT 76.800 822.300 78.600 827.400 ;
        RECT 82.800 822.300 84.600 827.400 ;
        RECT 88.950 823.950 91.050 826.050 ;
        RECT 94.800 824.400 96.600 827.400 ;
        RECT 76.800 820.950 84.600 822.300 ;
        RECT 74.400 818.250 78.150 819.300 ;
        RECT 76.950 818.100 78.150 818.250 ;
        RECT 74.100 815.100 75.900 815.850 ;
        RECT 76.950 814.950 79.050 817.050 ;
        RECT 80.100 815.100 81.900 815.850 ;
        RECT 82.950 814.950 85.200 817.050 ;
        RECT 52.950 811.950 55.050 814.050 ;
        RECT 31.950 810.450 34.050 811.050 ;
        RECT 26.550 809.550 34.050 810.450 ;
        RECT 10.800 795.600 12.600 807.600 ;
        RECT 13.800 806.700 21.600 807.600 ;
        RECT 13.800 795.600 15.600 806.700 ;
        RECT 19.800 795.600 21.600 806.700 ;
        RECT 26.550 805.050 27.450 809.550 ;
        RECT 31.950 808.950 34.050 809.550 ;
        RECT 37.950 808.950 40.050 811.050 ;
        RECT 46.950 808.950 49.050 811.050 ;
        RECT 56.850 810.900 57.900 813.900 ;
        RECT 58.950 811.950 61.050 814.050 ;
        RECT 62.100 813.150 63.900 813.900 ;
        RECT 67.950 811.950 70.050 814.050 ;
        RECT 73.950 811.950 76.050 814.050 ;
        RECT 77.850 810.900 78.900 813.900 ;
        RECT 79.950 811.950 82.050 814.050 ;
        RECT 83.100 813.150 84.900 813.900 ;
        RECT 89.550 813.450 90.450 823.950 ;
        RECT 95.400 815.100 96.600 824.400 ;
        RECT 97.950 817.950 100.050 820.050 ;
        RECT 113.100 819.000 114.900 827.400 ;
        RECT 135.000 823.050 136.800 827.400 ;
        RECT 124.950 820.950 127.050 823.050 ;
        RECT 131.400 821.400 136.800 823.050 ;
        RECT 151.800 821.400 153.600 827.400 ;
        RECT 157.800 824.400 159.600 827.400 ;
        RECT 113.100 817.350 117.300 819.000 ;
        RECT 98.100 816.150 99.900 816.900 ;
        RECT 107.100 815.100 108.900 815.850 ;
        RECT 113.100 815.100 114.900 815.850 ;
        RECT 94.950 813.450 97.050 814.050 ;
        RECT 89.550 812.550 97.050 813.450 ;
        RECT 94.950 811.950 97.050 812.550 ;
        RECT 106.950 811.950 109.050 814.050 ;
        RECT 112.950 811.950 115.050 814.050 ;
        RECT 116.400 812.100 117.300 817.350 ;
        RECT 125.550 816.450 126.450 820.950 ;
        RECT 131.400 818.100 132.300 821.400 ;
        RECT 130.950 816.450 133.050 817.050 ;
        RECT 125.550 815.550 133.050 816.450 ;
        RECT 130.950 814.950 133.050 815.550 ;
        RECT 134.100 815.100 135.900 815.850 ;
        RECT 136.950 814.950 139.050 817.050 ;
        RECT 140.100 815.100 141.900 815.850 ;
        RECT 151.950 815.100 153.000 821.400 ;
        RECT 157.800 820.200 158.700 824.400 ;
        RECT 175.200 820.200 177.000 827.400 ;
        RECT 155.250 819.300 158.700 820.200 ;
        RECT 155.250 818.400 157.050 819.300 ;
        RECT 25.950 802.950 28.050 805.050 ;
        RECT 32.700 802.800 33.600 807.900 ;
        RECT 38.100 807.150 39.900 807.900 ;
        RECT 56.850 807.600 58.050 810.900 ;
        RECT 77.850 807.600 79.050 810.900 ;
        RECT 32.700 801.900 39.300 802.800 ;
        RECT 32.700 801.600 33.600 801.900 ;
        RECT 31.800 795.600 33.600 801.600 ;
        RECT 37.800 801.600 39.300 801.900 ;
        RECT 37.800 795.600 39.600 801.600 ;
        RECT 56.700 795.600 58.500 807.600 ;
        RECT 77.700 795.600 79.500 807.600 ;
        RECT 95.400 801.600 96.600 810.900 ;
        RECT 109.950 808.950 112.050 811.050 ;
        RECT 115.950 810.450 118.050 811.050 ;
        RECT 115.950 809.550 123.450 810.450 ;
        RECT 115.950 808.950 118.050 809.550 ;
        RECT 110.100 807.150 111.900 807.900 ;
        RECT 116.400 802.800 117.300 807.900 ;
        RECT 110.700 801.900 117.300 802.800 ;
        RECT 122.550 802.050 123.450 809.550 ;
        RECT 131.400 807.600 132.300 813.900 ;
        RECT 133.950 811.950 136.050 814.050 ;
        RECT 137.100 813.150 138.900 813.900 ;
        RECT 139.950 811.950 142.050 814.050 ;
        RECT 148.950 811.950 154.050 814.050 ;
        RECT 152.700 807.600 154.050 810.900 ;
        RECT 155.400 810.600 156.300 818.400 ;
        RECT 160.950 817.950 163.050 820.050 ;
        RECT 173.400 819.300 177.000 820.200 ;
        RECT 198.000 821.400 199.800 827.400 ;
        RECT 157.950 814.950 160.050 817.050 ;
        RECT 161.100 816.150 162.900 816.900 ;
        RECT 173.400 815.100 174.600 819.300 ;
        RECT 198.000 818.100 199.050 821.400 ;
        RECT 217.200 820.200 219.000 827.400 ;
        RECT 215.400 819.300 219.000 820.200 ;
        RECT 190.950 814.950 193.050 817.050 ;
        RECT 194.250 815.100 195.900 815.850 ;
        RECT 196.950 814.950 199.050 817.050 ;
        RECT 200.100 815.100 201.750 815.850 ;
        RECT 202.950 814.950 205.050 817.050 ;
        RECT 215.400 815.100 216.600 819.300 ;
        RECT 236.100 819.000 237.900 827.400 ;
        RECT 257.100 819.000 258.900 827.400 ;
        RECT 276.000 820.200 277.800 827.400 ;
        RECT 276.000 819.300 279.600 820.200 ;
        RECT 236.100 817.350 240.300 819.000 ;
        RECT 257.100 817.350 261.300 819.000 ;
        RECT 230.100 815.100 231.900 815.850 ;
        RECT 236.100 815.100 237.900 815.850 ;
        RECT 158.100 813.150 159.900 813.900 ;
        RECT 170.100 812.100 171.900 812.850 ;
        RECT 172.950 811.950 175.050 814.050 ;
        RECT 191.100 813.150 192.900 813.900 ;
        RECT 176.100 812.100 177.900 812.850 ;
        RECT 193.950 811.950 196.050 814.050 ;
        RECT 155.400 810.000 157.200 810.600 ;
        RECT 155.400 808.800 162.600 810.000 ;
        RECT 169.950 808.950 172.050 811.050 ;
        RECT 155.400 808.650 156.300 808.800 ;
        RECT 161.400 807.600 162.600 808.800 ;
        RECT 110.700 801.600 112.200 801.900 ;
        RECT 94.800 795.600 96.600 801.600 ;
        RECT 110.400 795.600 112.200 801.600 ;
        RECT 116.400 801.600 117.300 801.900 ;
        RECT 116.400 795.600 118.200 801.600 ;
        RECT 121.950 799.950 124.050 802.050 ;
        RECT 130.800 795.600 132.600 807.600 ;
        RECT 133.800 806.700 141.600 807.600 ;
        RECT 133.800 795.600 135.600 806.700 ;
        RECT 139.800 795.600 141.600 806.700 ;
        RECT 152.700 806.100 155.100 807.600 ;
        RECT 153.300 795.600 155.100 806.100 ;
        RECT 160.800 795.600 162.600 807.600 ;
        RECT 173.400 801.600 174.600 810.900 ;
        RECT 175.950 808.950 178.050 811.050 ;
        RECT 197.100 810.900 197.850 813.900 ;
        RECT 199.950 811.950 202.050 814.050 ;
        RECT 203.100 813.150 204.750 813.900 ;
        RECT 212.100 812.100 213.900 812.850 ;
        RECT 214.950 811.950 217.050 814.050 ;
        RECT 218.100 812.100 219.900 812.850 ;
        RECT 229.950 811.950 232.050 814.050 ;
        RECT 235.950 811.950 238.050 814.050 ;
        RECT 239.400 812.100 240.300 817.350 ;
        RECT 251.100 815.100 252.900 815.850 ;
        RECT 257.100 815.100 258.900 815.850 ;
        RECT 250.950 811.950 253.050 814.050 ;
        RECT 256.950 811.950 259.050 814.050 ;
        RECT 260.400 812.100 261.300 817.350 ;
        RECT 278.400 815.100 279.600 819.300 ;
        RECT 296.100 819.000 297.900 827.400 ;
        RECT 293.700 817.350 297.900 819.000 ;
        RECT 317.100 819.000 318.900 827.400 ;
        RECT 337.200 820.200 339.000 827.400 ;
        RECT 352.800 824.400 354.600 827.400 ;
        RECT 335.400 819.300 339.000 820.200 ;
        RECT 317.100 817.350 321.300 819.000 ;
        RECT 275.100 812.100 276.900 812.850 ;
        RECT 277.950 811.950 280.050 814.050 ;
        RECT 281.100 812.100 282.900 812.850 ;
        RECT 293.700 812.100 294.600 817.350 ;
        RECT 296.100 815.100 297.900 815.850 ;
        RECT 302.100 815.100 303.900 815.850 ;
        RECT 311.100 815.100 312.900 815.850 ;
        RECT 317.100 815.100 318.900 815.850 ;
        RECT 295.950 811.950 298.050 814.050 ;
        RECT 301.950 811.950 304.050 814.050 ;
        RECT 310.950 811.950 313.200 814.050 ;
        RECT 316.950 811.950 319.050 814.050 ;
        RECT 320.400 812.100 321.300 817.350 ;
        RECT 335.400 815.100 336.600 819.300 ;
        RECT 353.400 815.100 354.600 824.400 ;
        RECT 355.950 817.950 358.050 820.050 ;
        RECT 371.100 819.000 372.900 827.400 ;
        RECT 389.400 824.400 391.200 827.400 ;
        RECT 371.100 817.350 375.300 819.000 ;
        RECT 385.950 817.950 388.050 820.050 ;
        RECT 356.100 816.150 357.900 816.900 ;
        RECT 365.100 815.100 366.900 815.850 ;
        RECT 371.100 815.100 372.900 815.850 ;
        RECT 332.100 812.100 333.900 812.850 ;
        RECT 334.950 811.950 337.050 814.050 ;
        RECT 352.950 813.450 355.050 814.050 ;
        RECT 357.000 813.450 360.900 814.050 ;
        RECT 338.100 812.100 339.900 812.850 ;
        RECT 352.950 812.550 360.900 813.450 ;
        RECT 352.950 811.950 355.050 812.550 ;
        RECT 357.000 811.950 360.900 812.550 ;
        RECT 364.950 811.950 367.050 814.050 ;
        RECT 370.950 811.950 373.050 814.050 ;
        RECT 374.400 812.100 375.300 817.350 ;
        RECT 386.100 816.150 387.900 816.900 ;
        RECT 389.400 815.100 390.600 824.400 ;
        RECT 407.100 819.000 408.900 827.400 ;
        RECT 428.100 819.000 429.900 827.400 ;
        RECT 447.000 820.200 448.800 827.400 ;
        RECT 463.800 821.400 465.600 827.400 ;
        RECT 469.800 824.400 471.600 827.400 ;
        RECT 447.000 819.300 450.600 820.200 ;
        RECT 404.700 817.350 408.900 819.000 ;
        RECT 425.700 817.350 429.900 819.000 ;
        RECT 388.950 811.950 394.050 814.050 ;
        RECT 404.700 812.100 405.600 817.350 ;
        RECT 407.100 815.100 408.900 815.850 ;
        RECT 413.100 815.100 414.900 815.850 ;
        RECT 406.950 811.950 409.050 814.050 ;
        RECT 412.950 811.950 415.050 814.050 ;
        RECT 425.700 812.100 426.600 817.350 ;
        RECT 428.100 815.100 429.900 815.850 ;
        RECT 434.100 815.100 435.900 815.850 ;
        RECT 449.400 815.100 450.600 819.300 ;
        RECT 457.950 817.950 460.050 820.050 ;
        RECT 427.950 811.950 430.050 814.050 ;
        RECT 433.950 811.950 436.050 814.050 ;
        RECT 446.100 812.100 447.900 812.850 ;
        RECT 448.950 811.950 451.050 814.050 ;
        RECT 458.550 813.450 459.450 817.950 ;
        RECT 463.950 815.100 465.000 821.400 ;
        RECT 469.800 820.200 470.700 824.400 ;
        RECT 487.200 820.200 489.000 827.400 ;
        RECT 502.800 821.400 504.600 827.400 ;
        RECT 467.250 819.300 470.700 820.200 ;
        RECT 467.250 818.400 469.050 819.300 ;
        RECT 463.950 813.450 466.050 814.050 ;
        RECT 452.100 812.100 453.900 812.850 ;
        RECT 458.550 812.550 466.050 813.450 ;
        RECT 463.950 811.950 466.050 812.550 ;
        RECT 196.950 809.400 197.850 810.900 ;
        RECT 193.800 808.500 197.850 809.400 ;
        RECT 211.950 808.950 214.050 811.050 ;
        RECT 184.950 805.950 187.050 808.050 ;
        RECT 185.550 802.050 186.450 805.950 ;
        RECT 173.400 795.600 175.200 801.600 ;
        RECT 184.950 799.950 187.050 802.050 ;
        RECT 190.800 796.500 192.600 807.600 ;
        RECT 193.800 797.400 195.600 808.500 ;
        RECT 196.800 806.400 204.600 807.300 ;
        RECT 196.800 796.500 198.600 806.400 ;
        RECT 190.800 795.600 198.600 796.500 ;
        RECT 202.800 795.600 204.600 806.400 ;
        RECT 215.400 801.600 216.600 810.900 ;
        RECT 217.950 808.950 220.050 811.050 ;
        RECT 232.950 808.950 235.050 811.050 ;
        RECT 238.950 810.450 241.050 811.050 ;
        RECT 238.950 809.550 246.450 810.450 ;
        RECT 238.950 808.950 241.050 809.550 ;
        RECT 233.100 807.150 234.900 807.900 ;
        RECT 239.400 802.800 240.300 807.900 ;
        RECT 233.700 801.900 240.300 802.800 ;
        RECT 233.700 801.600 235.200 801.900 ;
        RECT 215.400 795.600 217.200 801.600 ;
        RECT 233.400 795.600 235.200 801.600 ;
        RECT 239.400 801.600 240.300 801.900 ;
        RECT 239.400 795.600 241.200 801.600 ;
        RECT 245.550 799.050 246.450 809.550 ;
        RECT 253.950 808.950 256.050 811.050 ;
        RECT 259.950 810.450 262.050 811.050 ;
        RECT 259.950 809.550 267.450 810.450 ;
        RECT 259.950 808.950 262.050 809.550 ;
        RECT 254.100 807.150 255.900 807.900 ;
        RECT 260.400 802.800 261.300 807.900 ;
        RECT 266.550 805.050 267.450 809.550 ;
        RECT 274.950 808.950 277.050 811.050 ;
        RECT 265.950 802.950 268.050 805.050 ;
        RECT 254.700 801.900 261.300 802.800 ;
        RECT 254.700 801.600 256.200 801.900 ;
        RECT 244.950 796.950 247.050 799.050 ;
        RECT 254.400 795.600 256.200 801.600 ;
        RECT 260.400 801.600 261.300 801.900 ;
        RECT 278.400 801.600 279.600 810.900 ;
        RECT 280.950 805.950 283.050 811.050 ;
        RECT 289.950 808.950 295.050 811.050 ;
        RECT 298.950 808.950 301.050 811.050 ;
        RECT 313.950 808.950 316.050 811.050 ;
        RECT 319.950 810.450 322.050 811.050 ;
        RECT 324.000 810.450 327.900 811.050 ;
        RECT 319.950 809.550 327.900 810.450 ;
        RECT 319.950 808.950 322.050 809.550 ;
        RECT 324.000 808.950 327.900 809.550 ;
        RECT 331.950 808.950 334.050 811.050 ;
        RECT 293.700 802.800 294.600 807.900 ;
        RECT 299.100 807.150 300.900 807.900 ;
        RECT 314.100 807.150 315.900 807.900 ;
        RECT 320.400 802.800 321.300 807.900 ;
        RECT 293.700 801.900 300.300 802.800 ;
        RECT 293.700 801.600 294.600 801.900 ;
        RECT 260.400 795.600 262.200 801.600 ;
        RECT 277.800 795.600 279.600 801.600 ;
        RECT 292.800 795.600 294.600 801.600 ;
        RECT 298.800 801.600 300.300 801.900 ;
        RECT 314.700 801.900 321.300 802.800 ;
        RECT 314.700 801.600 316.200 801.900 ;
        RECT 298.800 795.600 300.600 801.600 ;
        RECT 314.400 795.600 316.200 801.600 ;
        RECT 320.400 801.600 321.300 801.900 ;
        RECT 335.400 801.600 336.600 810.900 ;
        RECT 337.950 808.950 340.050 811.050 ;
        RECT 353.400 801.600 354.600 810.900 ;
        RECT 367.950 808.950 370.050 811.050 ;
        RECT 373.950 810.450 376.050 811.050 ;
        RECT 373.950 809.550 381.450 810.450 ;
        RECT 373.950 808.950 376.050 809.550 ;
        RECT 368.100 807.150 369.900 807.900 ;
        RECT 374.400 802.800 375.300 807.900 ;
        RECT 380.550 805.050 381.450 809.550 ;
        RECT 379.950 802.950 382.050 805.050 ;
        RECT 368.700 801.900 375.300 802.800 ;
        RECT 368.700 801.600 370.200 801.900 ;
        RECT 320.400 795.600 322.200 801.600 ;
        RECT 335.400 795.600 337.200 801.600 ;
        RECT 352.800 795.600 354.600 801.600 ;
        RECT 368.400 795.600 370.200 801.600 ;
        RECT 374.400 801.600 375.300 801.900 ;
        RECT 389.400 801.600 390.600 810.900 ;
        RECT 400.950 808.950 406.050 811.050 ;
        RECT 409.950 808.950 412.050 811.050 ;
        RECT 418.950 810.450 423.000 811.050 ;
        RECT 424.950 810.450 427.050 811.050 ;
        RECT 418.950 809.550 427.050 810.450 ;
        RECT 418.950 808.950 423.000 809.550 ;
        RECT 424.950 808.950 427.050 809.550 ;
        RECT 430.800 808.950 433.050 811.050 ;
        RECT 445.950 808.950 448.050 811.050 ;
        RECT 404.700 802.800 405.600 807.900 ;
        RECT 410.100 807.150 411.900 807.900 ;
        RECT 425.700 802.800 426.600 807.900 ;
        RECT 431.100 807.150 432.900 807.900 ;
        RECT 404.700 801.900 411.300 802.800 ;
        RECT 404.700 801.600 405.600 801.900 ;
        RECT 374.400 795.600 376.200 801.600 ;
        RECT 389.400 795.600 391.200 801.600 ;
        RECT 403.800 795.600 405.600 801.600 ;
        RECT 409.800 801.600 411.300 801.900 ;
        RECT 425.700 801.900 432.300 802.800 ;
        RECT 425.700 801.600 426.600 801.900 ;
        RECT 409.800 795.600 411.600 801.600 ;
        RECT 424.800 795.600 426.600 801.600 ;
        RECT 430.800 801.600 432.300 801.900 ;
        RECT 449.400 801.600 450.600 810.900 ;
        RECT 451.950 808.950 454.050 811.050 ;
        RECT 457.950 805.950 460.050 808.050 ;
        RECT 464.700 807.600 466.050 810.900 ;
        RECT 467.400 810.600 468.300 818.400 ;
        RECT 472.950 817.950 475.050 820.050 ;
        RECT 485.400 819.300 489.000 820.200 ;
        RECT 503.400 819.300 504.600 821.400 ;
        RECT 505.800 822.300 507.600 827.400 ;
        RECT 511.800 822.300 513.600 827.400 ;
        RECT 505.800 820.950 513.600 822.300 ;
        RECT 525.000 820.200 526.800 827.400 ;
        RECT 541.800 821.400 543.600 827.400 ;
        RECT 525.000 819.300 528.600 820.200 ;
        RECT 469.950 814.950 472.050 817.050 ;
        RECT 473.100 816.150 474.900 816.900 ;
        RECT 485.400 815.100 486.600 819.300 ;
        RECT 503.400 818.250 507.150 819.300 ;
        RECT 505.950 818.100 507.150 818.250 ;
        RECT 503.100 815.100 504.900 815.850 ;
        RECT 505.950 814.950 508.200 817.050 ;
        RECT 509.100 815.100 510.900 815.850 ;
        RECT 511.950 814.950 514.050 817.050 ;
        RECT 527.400 815.100 528.600 819.300 ;
        RECT 542.400 819.300 543.600 821.400 ;
        RECT 544.800 822.300 546.600 827.400 ;
        RECT 550.800 822.300 552.600 827.400 ;
        RECT 544.800 820.950 552.600 822.300 ;
        RECT 564.000 820.200 565.800 827.400 ;
        RECT 585.000 823.050 586.800 827.400 ;
        RECT 601.800 824.400 603.600 827.400 ;
        RECT 616.800 824.400 618.600 827.400 ;
        RECT 581.400 821.400 586.800 823.050 ;
        RECT 564.000 819.300 567.600 820.200 ;
        RECT 542.400 818.250 546.150 819.300 ;
        RECT 544.950 818.100 546.150 818.250 ;
        RECT 535.950 814.950 538.050 817.050 ;
        RECT 542.100 815.100 543.900 815.850 ;
        RECT 544.950 814.950 547.050 817.050 ;
        RECT 548.100 815.100 549.900 815.850 ;
        RECT 550.950 814.950 553.050 817.050 ;
        RECT 566.400 815.100 567.600 819.300 ;
        RECT 581.400 818.100 582.300 821.400 ;
        RECT 580.950 816.450 583.050 817.050 ;
        RECT 575.550 815.550 583.050 816.450 ;
        RECT 470.100 813.150 471.900 813.900 ;
        RECT 475.950 811.950 478.050 814.050 ;
        RECT 482.100 812.100 483.900 812.850 ;
        RECT 484.950 811.950 487.050 814.050 ;
        RECT 488.100 812.100 489.900 812.850 ;
        RECT 502.950 811.950 505.050 814.050 ;
        RECT 467.400 810.000 469.200 810.600 ;
        RECT 467.400 808.800 474.600 810.000 ;
        RECT 467.400 808.650 468.300 808.800 ;
        RECT 473.400 807.600 474.600 808.800 ;
        RECT 476.550 808.050 477.450 811.950 ;
        RECT 481.800 808.950 484.050 811.050 ;
        RECT 464.700 806.100 467.100 807.600 ;
        RECT 430.800 795.600 432.600 801.600 ;
        RECT 448.800 795.600 450.600 801.600 ;
        RECT 458.550 799.050 459.450 805.950 ;
        RECT 457.950 796.950 460.050 799.050 ;
        RECT 465.300 795.600 467.100 806.100 ;
        RECT 472.800 795.600 474.600 807.600 ;
        RECT 475.950 805.950 478.050 808.050 ;
        RECT 485.400 801.600 486.600 810.900 ;
        RECT 487.950 808.950 490.050 811.050 ;
        RECT 506.850 810.900 507.900 813.900 ;
        RECT 508.950 811.950 511.050 814.050 ;
        RECT 512.100 813.150 513.900 813.900 ;
        RECT 524.100 812.100 525.900 812.850 ;
        RECT 526.950 811.950 529.050 814.050 ;
        RECT 530.100 812.100 531.900 812.850 ;
        RECT 536.550 811.050 537.450 814.950 ;
        RECT 541.800 811.950 544.050 814.050 ;
        RECT 506.850 807.600 508.050 810.900 ;
        RECT 523.950 808.950 526.050 811.050 ;
        RECT 485.400 795.600 487.200 801.600 ;
        RECT 506.700 795.600 508.500 807.600 ;
        RECT 527.400 801.600 528.600 810.900 ;
        RECT 529.950 808.950 532.050 811.050 ;
        RECT 535.950 808.950 538.050 811.050 ;
        RECT 545.850 810.900 546.900 813.900 ;
        RECT 547.950 811.950 550.050 814.050 ;
        RECT 551.100 813.150 552.900 813.900 ;
        RECT 563.100 812.100 564.900 812.850 ;
        RECT 565.800 811.950 568.050 814.050 ;
        RECT 569.100 812.100 570.900 812.850 ;
        RECT 545.850 807.600 547.050 810.900 ;
        RECT 562.800 808.950 565.050 811.050 ;
        RECT 526.800 795.600 528.600 801.600 ;
        RECT 545.700 795.600 547.500 807.600 ;
        RECT 566.400 801.600 567.600 810.900 ;
        RECT 568.950 808.950 571.200 811.050 ;
        RECT 565.800 795.600 567.600 801.600 ;
        RECT 575.550 799.050 576.450 815.550 ;
        RECT 580.950 814.950 583.050 815.550 ;
        RECT 584.100 815.100 585.900 815.850 ;
        RECT 586.950 814.950 589.050 817.050 ;
        RECT 590.100 815.100 591.900 815.850 ;
        RECT 595.950 814.950 598.050 817.050 ;
        RECT 602.400 815.100 603.600 824.400 ;
        RECT 604.950 817.950 607.050 820.050 ;
        RECT 605.100 816.150 606.900 816.900 ;
        RECT 617.400 815.100 618.600 824.400 ;
        RECT 635.100 819.000 636.900 827.400 ;
        RECT 652.800 824.400 654.600 827.400 ;
        RECT 635.100 817.350 639.300 819.000 ;
        RECT 620.100 816.150 621.900 816.900 ;
        RECT 629.100 815.100 630.900 815.850 ;
        RECT 635.100 815.100 636.900 815.850 ;
        RECT 581.400 807.600 582.300 813.900 ;
        RECT 583.950 811.950 586.050 814.050 ;
        RECT 587.100 813.150 588.900 813.900 ;
        RECT 589.950 811.950 592.050 814.050 ;
        RECT 596.550 808.050 597.450 814.950 ;
        RECT 601.950 811.950 604.050 814.050 ;
        RECT 616.950 811.950 622.050 814.050 ;
        RECT 628.950 811.950 631.050 814.050 ;
        RECT 634.950 811.950 637.200 814.050 ;
        RECT 638.400 812.100 639.300 817.350 ;
        RECT 653.400 815.100 654.600 824.400 ;
        RECT 665.400 822.300 667.200 827.400 ;
        RECT 671.400 822.300 673.200 827.400 ;
        RECT 665.400 820.950 673.200 822.300 ;
        RECT 674.400 821.400 676.200 827.400 ;
        RECT 686.400 822.300 688.200 827.400 ;
        RECT 692.400 822.300 694.200 827.400 ;
        RECT 674.400 819.300 675.600 821.400 ;
        RECT 686.400 820.950 694.200 822.300 ;
        RECT 695.400 821.400 697.200 827.400 ;
        RECT 707.400 822.300 709.200 827.400 ;
        RECT 713.400 822.300 715.200 827.400 ;
        RECT 695.400 819.300 696.600 821.400 ;
        RECT 707.400 820.950 715.200 822.300 ;
        RECT 716.400 821.400 718.200 827.400 ;
        RECT 732.300 823.200 734.100 827.400 ;
        RECT 732.150 821.400 734.100 823.200 ;
        RECT 716.400 819.300 717.600 821.400 ;
        RECT 671.850 818.250 675.600 819.300 ;
        RECT 692.850 818.250 696.600 819.300 ;
        RECT 713.850 818.250 717.600 819.300 ;
        RECT 671.850 818.100 673.050 818.250 ;
        RECT 692.850 818.100 694.050 818.250 ;
        RECT 713.850 818.100 715.050 818.250 ;
        RECT 732.150 818.100 733.050 821.400 ;
        RECT 734.100 819.900 735.900 820.500 ;
        RECT 739.800 819.900 741.600 827.400 ;
        RECT 752.400 824.400 754.200 827.400 ;
        RECT 752.400 821.100 753.600 824.400 ;
        RECT 760.950 823.950 763.050 826.050 ;
        RECT 770.400 824.400 772.200 827.400 ;
        RECT 788.400 824.400 790.200 827.400 ;
        RECT 734.100 818.700 741.600 819.900 ;
        RECT 656.100 816.150 657.900 816.900 ;
        RECT 668.100 815.100 669.900 815.850 ;
        RECT 670.950 814.950 673.200 817.050 ;
        RECT 674.100 815.100 675.900 815.850 ;
        RECT 685.950 814.950 688.050 817.050 ;
        RECT 689.100 815.100 690.900 815.850 ;
        RECT 691.950 814.950 694.050 817.050 ;
        RECT 695.100 815.100 696.900 815.850 ;
        RECT 706.950 814.950 709.050 817.050 ;
        RECT 710.100 815.100 711.900 815.850 ;
        RECT 712.950 814.950 715.200 817.050 ;
        RECT 716.100 815.100 717.900 815.850 ;
        RECT 727.950 814.950 733.050 817.050 ;
        RECT 734.100 815.100 735.900 815.850 ;
        RECT 652.950 813.450 655.050 814.050 ;
        RECT 647.550 812.550 655.050 813.450 ;
        RECT 665.100 813.150 666.900 813.900 ;
        RECT 574.800 796.950 576.900 799.050 ;
        RECT 580.800 795.600 582.600 807.600 ;
        RECT 583.800 806.700 591.600 807.600 ;
        RECT 583.800 795.600 585.600 806.700 ;
        RECT 589.800 795.600 591.600 806.700 ;
        RECT 595.950 805.950 598.050 808.050 ;
        RECT 602.400 801.600 603.600 810.900 ;
        RECT 617.400 801.600 618.600 810.900 ;
        RECT 631.950 808.950 634.050 811.050 ;
        RECT 637.950 810.450 640.050 811.050 ;
        RECT 637.950 809.550 645.450 810.450 ;
        RECT 637.950 808.950 640.050 809.550 ;
        RECT 632.100 807.150 633.900 807.900 ;
        RECT 638.400 802.800 639.300 807.900 ;
        RECT 632.700 801.900 639.300 802.800 ;
        RECT 644.550 802.050 645.450 809.550 ;
        RECT 647.550 808.050 648.450 812.550 ;
        RECT 652.950 811.950 655.050 812.550 ;
        RECT 671.100 810.900 672.150 813.900 ;
        RECT 673.950 811.950 676.050 814.050 ;
        RECT 686.100 813.150 687.900 813.900 ;
        RECT 688.950 811.950 691.050 814.050 ;
        RECT 692.100 810.900 693.150 813.900 ;
        RECT 694.950 811.950 697.200 814.050 ;
        RECT 700.950 811.950 703.050 814.050 ;
        RECT 707.100 813.150 708.900 813.900 ;
        RECT 709.950 811.950 712.050 814.050 ;
        RECT 646.950 805.950 649.050 808.050 ;
        RECT 632.700 801.600 634.200 801.900 ;
        RECT 601.800 795.600 603.600 801.600 ;
        RECT 616.800 795.600 618.600 801.600 ;
        RECT 632.400 795.600 634.200 801.600 ;
        RECT 638.400 801.600 639.300 801.900 ;
        RECT 638.400 795.600 640.200 801.600 ;
        RECT 643.950 799.950 646.050 802.050 ;
        RECT 653.400 801.600 654.600 810.900 ;
        RECT 670.950 807.600 672.150 810.900 ;
        RECT 691.950 807.600 693.150 810.900 ;
        RECT 652.800 795.600 654.600 801.600 ;
        RECT 670.500 795.600 672.300 807.600 ;
        RECT 691.500 795.600 693.300 807.600 ;
        RECT 701.550 805.050 702.450 811.950 ;
        RECT 713.100 810.900 714.150 813.900 ;
        RECT 715.950 811.950 718.050 814.050 ;
        RECT 712.950 807.600 714.150 810.900 ;
        RECT 730.950 807.600 732.000 813.900 ;
        RECT 733.950 811.950 736.050 814.050 ;
        RECT 700.950 802.950 703.050 805.050 ;
        RECT 712.500 795.600 714.300 807.600 ;
        RECT 730.200 795.600 732.000 807.600 ;
        RECT 737.550 801.600 738.600 818.700 ;
        RECT 751.950 817.950 754.050 820.050 ;
        RECT 739.950 814.950 742.050 817.050 ;
        RECT 752.700 813.900 753.900 816.900 ;
        RECT 754.950 814.950 757.050 817.050 ;
        RECT 740.100 813.150 741.900 813.900 ;
        RECT 749.100 813.150 750.900 813.900 ;
        RECT 752.700 808.650 754.050 813.900 ;
        RECT 755.100 813.150 756.900 813.900 ;
        RECT 752.700 807.600 755.400 808.650 ;
        RECT 736.800 795.600 738.600 801.600 ;
        RECT 753.600 795.600 755.400 807.600 ;
        RECT 761.550 799.050 762.450 823.950 ;
        RECT 770.400 821.100 771.600 824.400 ;
        RECT 789.300 820.200 790.200 824.400 ;
        RECT 794.400 821.400 796.200 827.400 ;
        RECT 806.400 822.000 808.200 827.400 ;
        RECT 812.400 826.500 820.200 827.400 ;
        RECT 812.400 822.000 814.200 826.500 ;
        RECT 769.950 817.950 772.050 820.050 ;
        RECT 784.800 817.950 787.050 820.050 ;
        RECT 789.300 819.300 792.750 820.200 ;
        RECT 790.950 818.400 792.750 819.300 ;
        RECT 770.700 813.900 771.900 816.900 ;
        RECT 772.950 814.950 775.050 817.050 ;
        RECT 785.100 816.150 786.900 816.900 ;
        RECT 787.950 814.950 790.050 817.050 ;
        RECT 767.100 813.150 768.900 813.900 ;
        RECT 770.700 808.650 772.050 813.900 ;
        RECT 773.100 813.150 774.900 813.900 ;
        RECT 788.100 813.150 789.900 813.900 ;
        RECT 791.700 810.600 792.600 818.400 ;
        RECT 795.000 815.100 796.050 821.400 ;
        RECT 806.400 821.100 814.200 822.000 ;
        RECT 815.400 821.400 817.200 825.600 ;
        RECT 818.400 821.400 820.200 826.500 ;
        RECT 840.000 821.400 841.800 827.400 ;
        RECT 815.700 819.900 816.600 821.400 ;
        RECT 806.250 818.100 808.050 818.850 ;
        RECT 812.400 818.700 816.600 819.900 ;
        RECT 812.400 818.100 813.600 818.700 ;
        RECT 817.500 818.100 819.300 818.850 ;
        RECT 840.000 818.100 841.050 821.400 ;
        RECT 805.950 814.950 808.050 817.050 ;
        RECT 809.100 815.100 810.900 815.850 ;
        RECT 811.950 814.950 814.050 817.050 ;
        RECT 815.100 815.100 816.750 815.850 ;
        RECT 817.950 814.950 820.050 817.050 ;
        RECT 832.950 814.950 835.050 817.050 ;
        RECT 836.250 815.100 837.900 815.850 ;
        RECT 838.950 814.950 841.050 817.050 ;
        RECT 842.100 815.100 843.750 815.850 ;
        RECT 844.950 814.950 847.050 817.050 ;
        RECT 793.950 811.950 796.050 814.050 ;
        RECT 808.950 811.950 811.050 814.050 ;
        RECT 790.800 810.000 792.600 810.600 ;
        RECT 785.400 808.800 792.600 810.000 ;
        RECT 770.700 807.600 773.400 808.650 ;
        RECT 760.950 796.950 763.050 799.050 ;
        RECT 771.600 795.600 773.400 807.600 ;
        RECT 785.400 807.600 786.600 808.800 ;
        RECT 791.700 808.650 792.600 808.800 ;
        RECT 793.950 807.600 795.300 810.900 ;
        RECT 812.400 807.600 813.600 813.900 ;
        RECT 814.950 811.950 817.050 814.050 ;
        RECT 833.100 813.150 834.900 813.900 ;
        RECT 835.950 811.950 838.200 814.050 ;
        RECT 839.100 810.900 839.850 813.900 ;
        RECT 841.800 811.950 844.050 814.050 ;
        RECT 845.100 813.150 846.750 813.900 ;
        RECT 838.950 809.400 839.850 810.900 ;
        RECT 835.800 808.500 839.850 809.400 ;
        RECT 785.400 795.600 787.200 807.600 ;
        RECT 792.900 806.100 795.300 807.600 ;
        RECT 792.900 795.600 794.700 806.100 ;
        RECT 810.900 795.600 814.200 807.600 ;
        RECT 832.800 796.500 834.600 807.600 ;
        RECT 835.800 797.400 837.600 808.500 ;
        RECT 838.800 806.400 846.600 807.300 ;
        RECT 838.800 796.500 840.600 806.400 ;
        RECT 832.800 795.600 840.600 796.500 ;
        RECT 844.800 795.600 846.600 806.400 ;
        RECT 12.600 779.400 14.400 791.400 ;
        RECT 22.950 787.950 25.050 790.050 ;
        RECT 12.600 778.350 15.300 779.400 ;
        RECT 11.100 773.100 12.900 773.850 ;
        RECT 13.950 773.100 15.300 778.350 ;
        RECT 17.100 773.100 18.900 773.850 ;
        RECT 10.950 769.950 13.050 772.050 ;
        RECT 14.100 770.100 15.300 773.100 ;
        RECT 16.950 769.950 19.050 772.050 ;
        RECT 23.550 769.050 24.450 787.950 ;
        RECT 31.800 785.400 33.600 791.400 ;
        RECT 28.950 775.950 31.050 778.050 ;
        RECT 32.400 776.100 33.600 785.400 ;
        RECT 40.950 784.950 43.050 787.050 ;
        RECT 41.550 781.050 42.450 784.950 ;
        RECT 40.950 778.950 43.050 781.050 ;
        RECT 46.800 779.400 48.600 791.400 ;
        RECT 49.800 780.300 51.600 791.400 ;
        RECT 55.800 780.300 57.600 791.400 ;
        RECT 68.400 785.400 70.200 791.400 ;
        RECT 68.700 785.100 70.200 785.400 ;
        RECT 74.400 785.400 76.200 791.400 ;
        RECT 74.400 785.100 75.300 785.400 ;
        RECT 68.700 784.200 75.300 785.100 ;
        RECT 49.800 779.400 57.600 780.300 ;
        RECT 34.950 775.950 37.050 778.050 ;
        RECT 41.550 775.050 42.450 778.950 ;
        RECT 29.100 774.150 30.900 774.900 ;
        RECT 31.950 772.950 34.050 775.050 ;
        RECT 35.100 774.150 36.900 774.900 ;
        RECT 40.950 772.950 43.050 775.050 ;
        RECT 47.400 773.100 48.300 779.400 ;
        RECT 68.100 779.100 69.900 779.850 ;
        RECT 74.400 779.100 75.300 784.200 ;
        RECT 88.200 779.400 90.000 791.400 ;
        RECT 94.800 785.400 96.600 791.400 ;
        RECT 67.950 775.950 70.050 778.050 ;
        RECT 73.950 775.950 79.050 778.050 ;
        RECT 49.950 772.950 52.050 775.050 ;
        RECT 53.100 773.100 54.900 773.850 ;
        RECT 55.950 772.950 58.050 775.050 ;
        RECT 64.950 772.950 67.050 775.050 ;
        RECT 70.950 772.950 73.050 775.050 ;
        RECT 13.950 766.950 16.050 769.050 ;
        RECT 22.950 766.950 25.050 769.050 ;
        RECT 32.400 767.700 33.600 771.900 ;
        RECT 46.950 769.950 49.050 772.050 ;
        RECT 50.100 771.150 51.900 771.900 ;
        RECT 52.950 769.950 55.050 772.050 ;
        RECT 56.100 771.150 57.900 771.900 ;
        RECT 65.100 771.150 66.900 771.900 ;
        RECT 71.100 771.150 72.900 771.900 ;
        RECT 74.400 769.650 75.300 774.900 ;
        RECT 88.950 773.100 90.000 779.400 ;
        RECT 91.950 772.950 94.050 775.050 ;
        RECT 85.950 769.950 91.050 772.050 ;
        RECT 92.100 771.150 93.900 771.900 ;
        RECT 30.000 766.800 33.600 767.700 ;
        RECT 14.400 762.600 15.600 765.900 ;
        RECT 13.800 759.600 15.600 762.600 ;
        RECT 30.000 759.600 31.800 766.800 ;
        RECT 47.400 765.600 48.300 768.900 ;
        RECT 71.100 768.000 75.300 769.650 ;
        RECT 47.400 763.950 52.800 765.600 ;
        RECT 51.000 759.600 52.800 763.950 ;
        RECT 71.100 759.600 72.900 768.000 ;
        RECT 90.150 765.600 91.050 768.900 ;
        RECT 95.550 768.300 96.600 785.400 ;
        RECT 113.700 779.400 115.500 791.400 ;
        RECT 133.500 779.400 135.300 791.400 ;
        RECT 103.950 775.950 106.050 778.050 ;
        RECT 113.850 776.100 115.050 779.400 ;
        RECT 133.950 776.100 135.150 779.400 ;
        RECT 145.950 778.950 148.050 781.050 ;
        RECT 151.200 779.400 153.000 791.400 ;
        RECT 157.800 785.400 159.600 791.400 ;
        RECT 98.100 773.100 99.900 773.850 ;
        RECT 104.550 772.050 105.450 775.950 ;
        RECT 109.950 772.950 112.050 775.050 ;
        RECT 113.850 773.100 114.900 776.100 ;
        RECT 115.950 772.950 118.200 775.050 ;
        RECT 119.100 773.100 120.900 773.850 ;
        RECT 128.100 773.100 129.900 773.850 ;
        RECT 130.800 772.950 133.050 775.050 ;
        RECT 134.100 773.100 135.150 776.100 ;
        RECT 136.950 772.950 139.200 775.050 ;
        RECT 97.950 769.950 100.050 772.050 ;
        RECT 104.100 769.950 106.200 772.050 ;
        RECT 110.100 771.150 111.900 771.900 ;
        RECT 112.950 769.950 115.050 772.050 ;
        RECT 116.100 771.150 117.900 771.900 ;
        RECT 118.950 769.950 121.050 772.050 ;
        RECT 127.950 769.950 130.050 772.050 ;
        RECT 131.100 771.150 132.900 771.900 ;
        RECT 133.800 769.950 136.050 772.050 ;
        RECT 137.100 771.150 138.900 771.900 ;
        RECT 146.550 771.450 147.450 778.950 ;
        RECT 151.950 773.100 153.000 779.400 ;
        RECT 154.950 772.950 157.050 775.050 ;
        RECT 151.950 771.450 154.050 772.050 ;
        RECT 146.550 770.550 154.050 771.450 ;
        RECT 155.100 771.150 156.900 771.900 ;
        RECT 151.950 769.950 154.050 770.550 ;
        RECT 112.950 768.750 114.150 768.900 ;
        RECT 92.100 767.100 99.600 768.300 ;
        RECT 92.100 766.500 93.900 767.100 ;
        RECT 90.150 763.800 92.100 765.600 ;
        RECT 90.300 759.600 92.100 763.800 ;
        RECT 97.800 759.600 99.600 767.100 ;
        RECT 110.400 767.700 114.150 768.750 ;
        RECT 134.850 768.750 136.050 768.900 ;
        RECT 134.850 767.700 138.600 768.750 ;
        RECT 110.400 765.600 111.600 767.700 ;
        RECT 109.800 759.600 111.600 765.600 ;
        RECT 112.800 764.700 120.600 766.050 ;
        RECT 112.800 759.600 114.600 764.700 ;
        RECT 118.800 759.600 120.600 764.700 ;
        RECT 128.400 764.700 136.200 766.050 ;
        RECT 128.400 759.600 130.200 764.700 ;
        RECT 134.400 759.600 136.200 764.700 ;
        RECT 137.400 765.600 138.600 767.700 ;
        RECT 153.150 765.600 154.050 768.900 ;
        RECT 158.550 768.300 159.600 785.400 ;
        RECT 174.600 779.400 176.400 791.400 ;
        RECT 190.800 779.400 192.600 791.400 ;
        RECT 193.800 780.300 195.600 791.400 ;
        RECT 199.800 780.300 201.600 791.400 ;
        RECT 211.800 785.400 213.600 791.400 ;
        RECT 193.800 779.400 201.600 780.300 ;
        RECT 212.700 785.100 213.600 785.400 ;
        RECT 217.800 785.400 219.600 791.400 ;
        RECT 233.400 785.400 235.200 791.400 ;
        RECT 217.800 785.100 219.300 785.400 ;
        RECT 212.700 784.200 219.300 785.100 ;
        RECT 173.700 778.350 176.400 779.400 ;
        RECT 161.100 773.100 162.900 773.850 ;
        RECT 170.100 773.100 171.900 773.850 ;
        RECT 173.700 773.100 175.050 778.350 ;
        RECT 176.100 773.100 177.900 773.850 ;
        RECT 191.400 773.100 192.300 779.400 ;
        RECT 212.700 779.100 213.600 784.200 ;
        RECT 218.100 779.100 219.900 779.850 ;
        RECT 208.950 775.950 214.050 778.050 ;
        RECT 217.950 775.950 220.050 778.050 ;
        RECT 229.950 775.950 232.050 778.050 ;
        RECT 233.400 776.100 234.600 785.400 ;
        RECT 250.200 779.400 252.000 791.400 ;
        RECT 256.800 785.400 258.600 791.400 ;
        RECT 265.950 787.950 268.050 790.050 ;
        RECT 235.950 775.950 238.050 778.050 ;
        RECT 160.950 769.950 163.050 772.050 ;
        RECT 169.950 769.950 172.050 772.050 ;
        RECT 173.700 770.100 174.900 773.100 ;
        RECT 193.950 772.950 196.050 775.050 ;
        RECT 197.100 773.100 198.900 773.850 ;
        RECT 199.950 772.950 202.050 775.050 ;
        RECT 175.800 769.950 178.050 772.050 ;
        RECT 187.950 769.950 193.050 772.050 ;
        RECT 194.100 771.150 195.900 771.900 ;
        RECT 196.950 769.950 199.050 772.050 ;
        RECT 200.100 771.150 201.900 771.900 ;
        RECT 212.700 769.650 213.600 774.900 ;
        RECT 214.950 772.950 217.050 775.050 ;
        RECT 220.950 772.950 223.050 775.050 ;
        RECT 230.100 774.150 231.900 774.900 ;
        RECT 232.800 772.950 235.050 775.050 ;
        RECT 236.100 774.150 237.900 774.900 ;
        RECT 250.950 773.100 252.000 779.400 ;
        RECT 253.950 772.950 256.050 775.050 ;
        RECT 215.100 771.150 216.900 771.900 ;
        RECT 221.100 771.150 222.900 771.900 ;
        RECT 155.100 767.100 162.600 768.300 ;
        RECT 155.100 766.500 156.900 767.100 ;
        RECT 137.400 759.600 139.200 765.600 ;
        RECT 153.150 763.800 155.100 765.600 ;
        RECT 153.300 759.600 155.100 763.800 ;
        RECT 160.800 759.600 162.600 767.100 ;
        RECT 172.800 766.950 175.050 769.050 ;
        RECT 173.400 762.600 174.600 765.900 ;
        RECT 191.400 765.600 192.300 768.900 ;
        RECT 212.700 768.000 216.900 769.650 ;
        RECT 191.400 763.950 196.800 765.600 ;
        RECT 173.400 759.600 175.200 762.600 ;
        RECT 195.000 759.600 196.800 763.950 ;
        RECT 215.100 759.600 216.900 768.000 ;
        RECT 233.400 767.700 234.600 771.900 ;
        RECT 247.950 769.950 253.050 772.050 ;
        RECT 254.100 771.150 255.900 771.900 ;
        RECT 233.400 766.800 237.000 767.700 ;
        RECT 235.200 759.600 237.000 766.800 ;
        RECT 252.150 765.600 253.050 768.900 ;
        RECT 257.550 768.300 258.600 785.400 ;
        RECT 266.550 777.450 267.450 787.950 ;
        RECT 271.800 785.400 273.600 791.400 ;
        RECT 272.700 785.100 273.600 785.400 ;
        RECT 277.800 785.400 279.600 791.400 ;
        RECT 293.400 785.400 295.200 791.400 ;
        RECT 277.800 785.100 279.300 785.400 ;
        RECT 272.700 784.200 279.300 785.100 ;
        RECT 272.700 779.100 273.600 784.200 ;
        RECT 278.100 779.100 279.900 779.850 ;
        RECT 271.950 777.450 274.050 778.050 ;
        RECT 266.550 776.550 274.050 777.450 ;
        RECT 271.950 775.950 274.050 776.550 ;
        RECT 277.800 775.950 280.050 778.050 ;
        RECT 289.950 775.950 292.050 778.050 ;
        RECT 293.400 776.100 294.600 785.400 ;
        RECT 314.700 779.400 316.500 791.400 ;
        RECT 335.700 779.400 337.500 791.400 ;
        RECT 354.600 779.400 356.400 791.400 ;
        RECT 295.950 775.950 298.050 778.050 ;
        RECT 314.850 776.100 316.050 779.400 ;
        RECT 335.850 776.100 337.050 779.400 ;
        RECT 353.700 778.350 356.400 779.400 ;
        RECT 371.400 785.400 373.200 791.400 ;
        RECT 260.100 773.100 261.900 773.850 ;
        RECT 259.950 769.950 262.050 772.050 ;
        RECT 272.700 769.650 273.600 774.900 ;
        RECT 274.950 772.950 277.050 775.050 ;
        RECT 280.950 772.950 283.050 775.050 ;
        RECT 290.100 774.150 291.900 774.900 ;
        RECT 292.950 772.950 295.050 775.050 ;
        RECT 296.100 774.150 297.900 774.900 ;
        RECT 310.950 772.950 313.050 775.050 ;
        RECT 314.850 773.100 315.900 776.100 ;
        RECT 316.950 772.950 319.050 775.050 ;
        RECT 320.100 773.100 321.900 773.850 ;
        RECT 331.950 772.950 334.050 775.050 ;
        RECT 335.850 773.100 336.900 776.100 ;
        RECT 337.950 772.950 340.050 775.050 ;
        RECT 341.100 773.100 342.900 773.850 ;
        RECT 350.100 773.100 351.900 773.850 ;
        RECT 353.700 773.100 355.050 778.350 ;
        RECT 356.100 773.100 357.900 773.850 ;
        RECT 368.100 773.100 369.900 773.850 ;
        RECT 275.100 771.150 276.900 771.900 ;
        RECT 281.100 771.150 282.900 771.900 ;
        RECT 254.100 767.100 261.600 768.300 ;
        RECT 272.700 768.000 276.900 769.650 ;
        RECT 254.100 766.500 255.900 767.100 ;
        RECT 252.150 763.800 254.100 765.600 ;
        RECT 252.300 759.600 254.100 763.800 ;
        RECT 259.800 759.600 261.600 767.100 ;
        RECT 275.100 759.600 276.900 768.000 ;
        RECT 293.400 767.700 294.600 771.900 ;
        RECT 311.100 771.150 312.900 771.900 ;
        RECT 313.950 769.950 316.050 772.050 ;
        RECT 317.100 771.150 318.900 771.900 ;
        RECT 319.950 769.950 322.050 772.050 ;
        RECT 332.100 771.150 333.900 771.900 ;
        RECT 334.950 769.950 337.050 772.050 ;
        RECT 338.100 771.150 339.900 771.900 ;
        RECT 340.950 769.950 343.050 772.050 ;
        RECT 349.800 769.950 352.050 772.050 ;
        RECT 353.700 770.100 354.900 773.100 ;
        RECT 355.950 769.950 358.200 772.050 ;
        RECT 367.950 769.950 370.050 772.050 ;
        RECT 313.950 768.750 315.150 768.900 ;
        RECT 334.950 768.750 336.150 768.900 ;
        RECT 311.400 767.700 315.150 768.750 ;
        RECT 332.400 767.700 336.150 768.750 ;
        RECT 293.400 766.800 297.000 767.700 ;
        RECT 295.200 759.600 297.000 766.800 ;
        RECT 311.400 765.600 312.600 767.700 ;
        RECT 310.800 759.600 312.600 765.600 ;
        RECT 313.800 764.700 321.600 766.050 ;
        RECT 332.400 765.600 333.600 767.700 ;
        RECT 352.800 766.950 355.050 769.050 ;
        RECT 371.400 768.300 372.450 785.400 ;
        RECT 378.000 779.400 379.800 791.400 ;
        RECT 391.800 785.400 393.600 791.400 ;
        RECT 392.700 785.100 393.600 785.400 ;
        RECT 397.800 785.400 399.600 791.400 ;
        RECT 413.400 785.400 415.200 791.400 ;
        RECT 428.400 785.400 430.200 791.400 ;
        RECT 446.400 785.400 448.200 791.400 ;
        RECT 464.400 785.400 466.200 791.400 ;
        RECT 397.800 785.100 399.300 785.400 ;
        RECT 392.700 784.200 399.300 785.100 ;
        RECT 373.950 772.950 376.050 775.050 ;
        RECT 378.000 773.100 379.050 779.400 ;
        RECT 392.700 779.100 393.600 784.200 ;
        RECT 398.100 779.100 399.900 779.850 ;
        RECT 388.950 775.950 394.050 778.050 ;
        RECT 397.950 775.950 400.050 778.050 ;
        RECT 413.400 776.100 414.600 785.400 ;
        RECT 424.950 775.950 427.050 778.050 ;
        RECT 428.400 776.100 429.600 785.400 ;
        RECT 430.950 775.950 433.050 778.050 ;
        RECT 436.950 775.950 439.050 778.050 ;
        RECT 442.800 775.950 445.050 778.050 ;
        RECT 446.400 776.100 447.600 785.400 ;
        RECT 464.700 785.100 466.200 785.400 ;
        RECT 470.400 785.400 472.200 791.400 ;
        RECT 478.950 787.950 481.050 790.050 ;
        RECT 470.400 785.100 471.300 785.400 ;
        RECT 464.700 784.200 471.300 785.100 ;
        RECT 464.100 779.100 465.900 779.850 ;
        RECT 470.400 779.100 471.300 784.200 ;
        RECT 448.950 775.950 451.050 778.050 ;
        RECT 463.950 775.950 466.050 778.050 ;
        RECT 469.950 775.950 475.050 778.050 ;
        RECT 479.550 777.450 480.450 787.950 ;
        RECT 484.800 785.400 486.600 791.400 ;
        RECT 485.700 785.100 486.600 785.400 ;
        RECT 490.800 785.400 492.600 791.400 ;
        RECT 490.800 785.100 492.300 785.400 ;
        RECT 485.700 784.200 492.300 785.100 ;
        RECT 485.700 779.100 486.600 784.200 ;
        RECT 503.400 780.300 505.200 791.400 ;
        RECT 509.400 780.300 511.200 791.400 ;
        RECT 491.100 779.100 492.900 779.850 ;
        RECT 503.400 779.400 511.200 780.300 ;
        RECT 512.400 779.400 514.200 791.400 ;
        RECT 517.950 781.950 520.050 784.050 ;
        RECT 484.950 777.450 487.050 778.050 ;
        RECT 479.550 776.550 487.050 777.450 ;
        RECT 484.950 775.950 487.050 776.550 ;
        RECT 490.950 775.950 493.050 778.050 ;
        RECT 374.100 771.150 375.900 771.900 ;
        RECT 376.950 769.950 379.050 772.050 ;
        RECT 392.700 769.650 393.600 774.900 ;
        RECT 394.950 772.950 397.050 775.050 ;
        RECT 400.950 772.950 403.050 775.050 ;
        RECT 409.950 772.950 415.050 775.050 ;
        RECT 425.100 774.150 426.900 774.900 ;
        RECT 427.950 772.950 430.050 775.050 ;
        RECT 431.100 774.150 432.900 774.900 ;
        RECT 437.550 772.050 438.450 775.950 ;
        RECT 443.100 774.150 444.900 774.900 ;
        RECT 445.950 772.950 448.050 775.050 ;
        RECT 449.100 774.150 450.900 774.900 ;
        RECT 460.950 772.950 463.050 775.050 ;
        RECT 466.950 772.950 469.050 775.050 ;
        RECT 395.100 771.150 396.900 771.900 ;
        RECT 401.100 771.150 402.900 771.900 ;
        RECT 410.100 770.100 411.900 770.850 ;
        RECT 368.400 767.100 375.900 768.300 ;
        RECT 313.800 759.600 315.600 764.700 ;
        RECT 319.800 759.600 321.600 764.700 ;
        RECT 331.800 759.600 333.600 765.600 ;
        RECT 334.800 764.700 342.600 766.050 ;
        RECT 334.800 759.600 336.600 764.700 ;
        RECT 340.800 759.600 342.600 764.700 ;
        RECT 353.400 762.600 354.600 765.900 ;
        RECT 353.400 759.600 355.200 762.600 ;
        RECT 368.400 759.600 370.200 767.100 ;
        RECT 374.100 766.500 375.900 767.100 ;
        RECT 376.950 765.600 377.850 768.900 ;
        RECT 392.700 768.000 396.900 769.650 ;
        RECT 375.900 763.800 377.850 765.600 ;
        RECT 375.900 759.600 377.700 763.800 ;
        RECT 395.100 759.600 396.900 768.000 ;
        RECT 409.950 766.950 412.050 769.050 ;
        RECT 413.400 762.600 414.600 771.900 ;
        RECT 428.400 767.700 429.600 771.900 ;
        RECT 436.950 769.950 439.050 772.050 ;
        RECT 446.400 767.700 447.600 771.900 ;
        RECT 461.100 771.150 462.900 771.900 ;
        RECT 467.100 771.150 468.900 771.900 ;
        RECT 470.400 769.650 471.300 774.900 ;
        RECT 467.100 768.000 471.300 769.650 ;
        RECT 485.700 769.650 486.600 774.900 ;
        RECT 487.950 772.950 490.050 775.050 ;
        RECT 493.950 772.950 496.050 775.050 ;
        RECT 502.950 772.950 505.050 775.050 ;
        RECT 506.100 773.100 507.900 773.850 ;
        RECT 508.950 772.950 511.050 775.050 ;
        RECT 512.700 773.100 513.600 779.400 ;
        RECT 488.100 771.150 489.900 771.900 ;
        RECT 494.100 771.150 495.900 771.900 ;
        RECT 503.100 771.150 504.900 771.900 ;
        RECT 505.800 769.950 508.050 772.050 ;
        RECT 509.100 771.150 510.900 771.900 ;
        RECT 511.950 769.950 514.050 772.050 ;
        RECT 485.700 768.000 489.900 769.650 ;
        RECT 428.400 766.800 432.000 767.700 ;
        RECT 446.400 766.800 450.000 767.700 ;
        RECT 413.400 759.600 415.200 762.600 ;
        RECT 430.200 759.600 432.000 766.800 ;
        RECT 448.200 759.600 450.000 766.800 ;
        RECT 467.100 759.600 468.900 768.000 ;
        RECT 488.100 759.600 489.900 768.000 ;
        RECT 512.700 765.600 513.600 768.900 ;
        RECT 508.200 763.950 513.600 765.600 ;
        RECT 508.200 759.600 510.000 763.950 ;
        RECT 518.550 763.050 519.450 781.950 ;
        RECT 530.700 779.400 532.500 791.400 ;
        RECT 551.700 779.400 553.500 791.400 ;
        RECT 530.850 776.100 532.050 779.400 ;
        RECT 551.850 776.100 553.050 779.400 ;
        RECT 562.950 778.950 565.050 781.050 ;
        RECT 568.200 779.400 570.000 791.400 ;
        RECT 574.800 785.400 576.600 791.400 ;
        RECT 589.800 785.400 591.600 791.400 ;
        RECT 526.950 772.950 529.050 775.050 ;
        RECT 530.850 773.100 531.900 776.100 ;
        RECT 532.950 772.950 535.050 775.050 ;
        RECT 536.100 773.100 537.900 773.850 ;
        RECT 541.950 772.950 544.050 775.050 ;
        RECT 547.950 772.950 550.050 775.050 ;
        RECT 551.850 773.100 552.900 776.100 ;
        RECT 553.800 772.950 556.050 775.050 ;
        RECT 557.100 773.100 558.900 773.850 ;
        RECT 527.100 771.150 528.900 771.900 ;
        RECT 529.950 769.950 532.050 772.050 ;
        RECT 533.100 771.150 534.900 771.900 ;
        RECT 535.950 769.950 538.050 772.050 ;
        RECT 542.550 769.050 543.450 772.950 ;
        RECT 548.100 771.150 549.900 771.900 ;
        RECT 550.950 769.950 553.050 772.050 ;
        RECT 554.100 771.150 555.900 771.900 ;
        RECT 556.950 769.950 559.200 772.050 ;
        RECT 563.550 771.450 564.450 778.950 ;
        RECT 568.950 773.100 570.000 779.400 ;
        RECT 571.950 772.950 574.050 775.050 ;
        RECT 568.950 771.450 571.050 772.050 ;
        RECT 563.550 770.550 571.050 771.450 ;
        RECT 572.100 771.150 573.900 771.900 ;
        RECT 568.950 769.950 571.050 770.550 ;
        RECT 529.950 768.750 531.150 768.900 ;
        RECT 527.400 767.700 531.150 768.750 ;
        RECT 527.400 765.600 528.600 767.700 ;
        RECT 541.950 766.950 544.050 769.050 ;
        RECT 550.950 768.750 552.150 768.900 ;
        RECT 548.400 767.700 552.150 768.750 ;
        RECT 517.950 760.950 520.050 763.050 ;
        RECT 526.800 759.600 528.600 765.600 ;
        RECT 529.800 764.700 537.600 766.050 ;
        RECT 548.400 765.600 549.600 767.700 ;
        RECT 529.800 759.600 531.600 764.700 ;
        RECT 535.800 759.600 537.600 764.700 ;
        RECT 547.800 759.600 549.600 765.600 ;
        RECT 550.800 764.700 558.600 766.050 ;
        RECT 550.800 759.600 552.600 764.700 ;
        RECT 556.800 759.600 558.600 764.700 ;
        RECT 570.150 765.600 571.050 768.900 ;
        RECT 575.550 768.300 576.600 785.400 ;
        RECT 590.400 776.100 591.600 785.400 ;
        RECT 606.600 779.400 608.400 791.400 ;
        RECT 624.900 779.400 628.200 791.400 ;
        RECT 640.800 784.950 642.900 787.050 ;
        RECT 605.700 778.350 608.400 779.400 ;
        RECT 578.100 773.100 579.900 773.850 ;
        RECT 586.950 772.950 592.050 775.050 ;
        RECT 602.100 773.100 603.900 773.850 ;
        RECT 605.700 773.100 607.050 778.350 ;
        RECT 608.100 773.100 609.900 773.850 ;
        RECT 577.950 769.950 580.050 772.050 ;
        RECT 572.100 767.100 579.600 768.300 ;
        RECT 572.100 766.500 573.900 767.100 ;
        RECT 570.150 763.800 572.100 765.600 ;
        RECT 570.300 759.600 572.100 763.800 ;
        RECT 577.800 759.600 579.600 767.100 ;
        RECT 590.400 762.600 591.600 771.900 ;
        RECT 593.100 770.100 594.900 770.850 ;
        RECT 601.950 769.950 604.050 772.050 ;
        RECT 605.700 770.100 606.900 773.100 ;
        RECT 622.950 772.950 625.050 775.050 ;
        RECT 626.400 773.100 627.600 779.400 ;
        RECT 638.100 778.950 640.200 781.050 ;
        RECT 628.950 772.950 631.200 775.050 ;
        RECT 607.950 769.950 610.050 772.050 ;
        RECT 619.800 769.950 622.050 772.050 ;
        RECT 623.100 771.150 624.900 771.900 ;
        RECT 625.950 769.950 628.050 772.050 ;
        RECT 629.100 771.150 630.750 771.900 ;
        RECT 631.950 769.950 634.050 772.050 ;
        RECT 592.950 766.950 595.050 769.050 ;
        RECT 604.950 766.950 607.050 769.050 ;
        RECT 620.250 768.150 622.050 768.900 ;
        RECT 626.400 768.300 627.600 768.900 ;
        RECT 626.400 767.100 630.600 768.300 ;
        RECT 631.500 768.150 633.300 768.900 ;
        RECT 589.800 759.600 591.600 762.600 ;
        RECT 605.400 762.600 606.600 765.900 ;
        RECT 620.400 765.000 628.200 765.900 ;
        RECT 629.700 765.600 630.600 767.100 ;
        RECT 638.550 766.050 639.450 778.950 ;
        RECT 641.550 771.450 642.450 784.950 ;
        RECT 646.800 779.400 648.600 791.400 ;
        RECT 649.800 780.300 651.600 791.400 ;
        RECT 655.800 780.300 657.600 791.400 ;
        RECT 661.950 787.950 664.050 790.050 ;
        RECT 649.800 779.400 657.600 780.300 ;
        RECT 647.400 773.100 648.300 779.400 ;
        RECT 649.800 772.950 652.050 775.050 ;
        RECT 653.100 773.100 654.900 773.850 ;
        RECT 655.950 772.950 658.050 775.050 ;
        RECT 662.550 774.450 663.450 787.950 ;
        RECT 668.400 785.400 670.200 791.400 ;
        RECT 668.400 776.100 669.600 785.400 ;
        RECT 673.950 784.950 676.050 787.050 ;
        RECT 667.950 774.450 670.050 775.050 ;
        RECT 662.550 773.550 670.050 774.450 ;
        RECT 667.950 772.950 670.050 773.550 ;
        RECT 646.950 771.450 649.050 772.050 ;
        RECT 641.550 770.550 649.050 771.450 ;
        RECT 650.100 771.150 651.900 771.900 ;
        RECT 646.950 769.950 649.050 770.550 ;
        RECT 605.400 759.600 607.200 762.600 ;
        RECT 620.400 759.600 622.200 765.000 ;
        RECT 626.400 760.500 628.200 765.000 ;
        RECT 629.400 761.400 631.200 765.600 ;
        RECT 632.400 760.500 634.200 765.600 ;
        RECT 637.950 763.950 640.050 766.050 ;
        RECT 647.400 765.600 648.300 768.900 ;
        RECT 652.950 766.950 655.050 772.050 ;
        RECT 656.100 771.150 657.900 771.900 ;
        RECT 665.100 770.100 666.900 770.850 ;
        RECT 664.950 766.950 667.050 769.050 ;
        RECT 647.400 763.950 652.800 765.600 ;
        RECT 626.400 759.600 634.200 760.500 ;
        RECT 651.000 759.600 652.800 763.950 ;
        RECT 668.400 762.600 669.600 771.900 ;
        RECT 674.550 769.050 675.450 784.950 ;
        RECT 680.400 780.600 682.200 791.400 ;
        RECT 686.400 790.500 694.200 791.400 ;
        RECT 686.400 780.600 688.200 790.500 ;
        RECT 680.400 779.700 688.200 780.600 ;
        RECT 689.400 778.500 691.200 789.600 ;
        RECT 692.400 779.400 694.200 790.500 ;
        RECT 709.500 779.400 711.300 791.400 ;
        RECT 725.400 780.300 727.200 791.400 ;
        RECT 731.400 780.300 733.200 791.400 ;
        RECT 725.400 779.400 733.200 780.300 ;
        RECT 734.400 779.400 736.200 791.400 ;
        RECT 751.500 779.400 753.300 791.400 ;
        RECT 764.700 785.400 766.500 791.400 ;
        RECT 764.700 784.500 765.750 785.400 ;
        RECT 761.700 783.600 765.750 784.500 ;
        RECT 687.150 777.600 691.200 778.500 ;
        RECT 687.150 776.100 688.050 777.600 ;
        RECT 709.950 776.100 711.150 779.400 ;
        RECT 680.250 773.100 681.900 773.850 ;
        RECT 682.800 772.950 685.050 775.050 ;
        RECT 687.150 773.100 687.900 776.100 ;
        RECT 688.950 772.950 691.050 775.050 ;
        RECT 692.100 773.100 693.900 773.850 ;
        RECT 704.100 773.100 705.900 773.850 ;
        RECT 706.950 772.950 709.050 775.050 ;
        RECT 710.100 773.100 711.150 776.100 ;
        RECT 712.950 772.950 715.050 775.050 ;
        RECT 724.950 772.950 727.050 775.050 ;
        RECT 728.100 773.100 729.900 773.850 ;
        RECT 730.950 772.950 733.050 775.050 ;
        RECT 734.700 773.100 735.600 779.400 ;
        RECT 751.950 776.100 753.150 779.400 ;
        RECT 746.100 773.100 747.900 773.850 ;
        RECT 748.950 772.950 751.050 775.050 ;
        RECT 752.100 773.100 753.150 776.100 ;
        RECT 754.950 772.950 757.050 775.050 ;
        RECT 679.950 769.950 682.050 772.050 ;
        RECT 683.250 771.150 684.900 771.900 ;
        RECT 685.950 769.950 688.050 772.050 ;
        RECT 689.100 771.150 690.750 771.900 ;
        RECT 691.950 769.950 694.050 772.050 ;
        RECT 703.950 769.950 706.050 772.050 ;
        RECT 707.100 771.150 708.900 771.900 ;
        RECT 709.950 769.950 712.050 772.050 ;
        RECT 713.100 771.150 714.900 771.900 ;
        RECT 725.100 771.150 726.900 771.900 ;
        RECT 727.950 769.950 730.050 772.050 ;
        RECT 731.100 771.150 732.900 771.900 ;
        RECT 733.950 769.950 736.050 772.050 ;
        RECT 745.950 769.950 748.050 772.050 ;
        RECT 749.100 771.150 750.900 771.900 ;
        RECT 751.950 769.950 754.050 772.050 ;
        RECT 755.100 771.150 756.900 771.900 ;
        RECT 761.700 770.100 762.900 783.600 ;
        RECT 770.700 782.700 772.500 791.400 ;
        RECT 776.850 788.400 779.100 791.400 ;
        RECT 780.000 788.400 782.100 791.400 ;
        RECT 783.150 788.400 785.100 791.400 ;
        RECT 776.850 787.050 777.750 788.400 ;
        RECT 780.000 787.050 781.050 788.400 ;
        RECT 783.150 787.050 784.350 788.400 ;
        RECT 775.950 784.950 778.050 787.050 ;
        RECT 778.950 784.950 781.050 787.050 ;
        RECT 781.950 784.950 784.350 787.050 ;
        RECT 790.200 785.400 792.000 791.400 ;
        RECT 796.200 785.400 798.000 791.400 ;
        RECT 799.800 788.400 801.600 791.400 ;
        RECT 802.800 788.400 804.600 791.400 ;
        RECT 805.800 788.400 807.600 791.400 ;
        RECT 799.950 785.400 801.150 788.400 ;
        RECT 802.950 785.400 804.600 788.400 ;
        RECT 805.950 787.200 807.150 788.400 ;
        RECT 790.950 784.500 792.000 785.400 ;
        RECT 766.200 781.650 783.900 782.700 ;
        RECT 790.950 782.400 793.050 784.500 ;
        RECT 796.050 783.150 798.150 785.400 ;
        RECT 799.950 783.300 802.050 785.400 ;
        RECT 802.950 784.050 805.050 785.400 ;
        RECT 805.950 785.100 808.050 787.200 ;
        RECT 812.400 784.500 814.200 791.400 ;
        RECT 818.400 785.400 820.200 791.400 ;
        RECT 809.700 784.050 811.500 784.500 ;
        RECT 766.200 780.900 768.000 781.650 ;
        RECT 778.950 780.150 781.050 780.750 ;
        RECT 769.500 778.950 781.050 780.150 ;
        RECT 781.950 780.300 783.900 781.650 ;
        RECT 796.050 781.350 798.900 783.150 ;
        RECT 802.950 782.850 811.500 784.050 ;
        RECT 812.400 783.300 818.100 784.500 ;
        RECT 809.700 782.700 811.500 782.850 ;
        RECT 816.300 782.700 818.100 783.300 ;
        RECT 799.950 780.300 802.050 781.350 ;
        RECT 781.950 779.250 802.050 780.300 ;
        RECT 805.950 780.750 808.050 781.350 ;
        RECT 819.000 780.750 820.200 785.400 ;
        RECT 825.000 785.400 826.800 791.400 ;
        RECT 842.400 785.400 844.200 791.400 ;
        RECT 805.950 779.850 822.900 780.750 ;
        RECT 805.950 779.250 808.050 779.850 ;
        RECT 769.500 778.350 771.300 778.950 ;
        RECT 778.950 778.650 781.050 778.950 ;
        RECT 819.300 778.350 821.100 778.950 ;
        RECT 781.950 777.450 821.100 778.350 ;
        RECT 769.950 777.150 821.100 777.450 ;
        RECT 769.950 776.550 783.900 777.150 ;
        RECT 763.950 773.850 766.050 775.950 ;
        RECT 769.950 775.350 773.850 776.550 ;
        RECT 790.950 775.650 793.050 776.250 ;
        RECT 782.400 775.500 784.200 775.650 ;
        RECT 790.950 775.500 805.500 775.650 ;
        RECT 769.950 775.050 772.050 775.350 ;
        RECT 774.750 774.450 781.500 775.350 ;
        RECT 764.100 772.050 765.900 773.850 ;
        RECT 774.750 772.050 775.950 774.450 ;
        RECT 764.100 771.000 775.950 772.050 ;
        RECT 777.750 771.750 779.550 773.550 ;
        RECT 780.450 772.950 781.500 774.450 ;
        RECT 782.400 774.450 805.500 775.500 ;
        RECT 782.400 773.850 784.200 774.450 ;
        RECT 790.950 774.150 793.050 774.450 ;
        RECT 795.150 773.250 797.250 773.550 ;
        RECT 803.700 773.250 805.500 774.450 ;
        RECT 806.850 774.000 813.900 775.800 ;
        RECT 780.450 772.050 792.450 772.950 ;
        RECT 761.700 769.200 777.000 770.100 ;
        RECT 673.950 766.950 676.050 769.050 ;
        RECT 685.950 765.600 687.000 768.900 ;
        RECT 710.850 768.750 712.050 768.900 ;
        RECT 710.850 767.700 714.600 768.750 ;
        RECT 668.400 759.600 670.200 762.600 ;
        RECT 685.200 759.600 687.000 765.600 ;
        RECT 704.400 764.700 712.200 766.050 ;
        RECT 704.400 759.600 706.200 764.700 ;
        RECT 710.400 759.600 712.200 764.700 ;
        RECT 713.400 765.600 714.600 767.700 ;
        RECT 734.700 765.600 735.600 768.900 ;
        RECT 752.850 768.750 754.050 768.900 ;
        RECT 752.850 767.700 756.600 768.750 ;
        RECT 713.400 759.600 715.200 765.600 ;
        RECT 730.200 763.950 735.600 765.600 ;
        RECT 746.400 764.700 754.200 766.050 ;
        RECT 730.200 759.600 732.000 763.950 ;
        RECT 746.400 759.600 748.200 764.700 ;
        RECT 752.400 759.600 754.200 764.700 ;
        RECT 755.400 765.600 756.600 767.700 ;
        RECT 761.700 765.600 762.900 769.200 ;
        RECT 765.900 767.700 767.700 768.300 ;
        RECT 765.900 766.500 774.300 767.700 ;
        RECT 772.800 765.600 774.300 766.500 ;
        RECT 755.400 759.600 757.200 765.600 ;
        RECT 761.700 759.600 763.500 765.600 ;
        RECT 772.500 759.600 774.300 765.600 ;
        RECT 775.950 766.050 777.000 769.200 ;
        RECT 778.500 768.300 779.550 771.750 ;
        RECT 786.150 769.350 790.050 771.150 ;
        RECT 787.950 769.050 790.050 769.350 ;
        RECT 791.400 770.550 792.450 772.050 ;
        RECT 793.350 771.450 797.250 773.250 ;
        RECT 806.850 772.350 807.750 774.000 ;
        RECT 817.050 773.100 819.150 775.050 ;
        RECT 798.150 771.300 807.750 772.350 ;
        RECT 808.800 772.050 819.150 773.100 ;
        RECT 798.150 770.550 799.050 771.300 ;
        RECT 791.400 769.200 799.050 770.550 ;
        RECT 808.800 770.250 809.850 772.050 ;
        RECT 814.500 770.700 816.300 771.000 ;
        RECT 819.300 770.700 821.100 771.000 ;
        RECT 799.950 769.200 809.850 770.250 ;
        RECT 813.300 769.200 821.100 770.700 ;
        RECT 781.050 768.300 782.850 768.750 ;
        RECT 799.950 768.300 801.000 769.200 ;
        RECT 778.500 767.850 782.850 768.300 ;
        RECT 778.500 767.100 786.150 767.850 ;
        RECT 781.050 766.950 786.150 767.100 ;
        RECT 775.950 763.950 778.050 766.050 ;
        RECT 778.950 763.950 781.050 766.050 ;
        RECT 781.950 763.950 784.050 766.050 ;
        RECT 785.250 765.600 786.150 766.950 ;
        RECT 794.100 766.500 801.000 768.300 ;
        RECT 801.900 766.500 808.500 768.300 ;
        RECT 813.300 765.600 814.800 769.200 ;
        RECT 822.000 765.600 822.900 779.850 ;
        RECT 825.000 775.050 826.500 785.400 ;
        RECT 829.950 781.950 832.050 784.050 ;
        RECT 824.850 772.950 826.950 775.050 ;
        RECT 785.250 764.250 789.300 765.600 ;
        RECT 776.700 762.600 778.050 763.950 ;
        RECT 779.700 762.600 781.050 763.950 ;
        RECT 782.700 762.600 784.050 763.950 ;
        RECT 787.500 763.800 789.300 764.250 ;
        RECT 790.950 763.500 793.050 765.600 ;
        RECT 796.050 763.500 798.150 765.600 ;
        RECT 799.950 763.500 802.050 765.600 ;
        RECT 802.950 763.500 805.050 765.600 ;
        RECT 805.950 763.500 808.050 765.600 ;
        RECT 810.600 764.400 814.800 765.600 ;
        RECT 790.950 762.600 792.000 763.500 ;
        RECT 796.350 762.600 798.000 763.500 ;
        RECT 799.950 762.600 801.600 763.500 ;
        RECT 802.950 762.600 804.600 763.500 ;
        RECT 806.250 762.600 807.600 763.500 ;
        RECT 776.700 759.600 778.500 762.600 ;
        RECT 779.700 759.600 781.500 762.600 ;
        RECT 782.700 759.600 784.500 762.600 ;
        RECT 790.200 759.600 792.000 762.600 ;
        RECT 796.200 759.600 798.000 762.600 ;
        RECT 799.800 759.600 801.600 762.600 ;
        RECT 802.800 759.600 804.600 762.600 ;
        RECT 805.800 759.600 807.600 762.600 ;
        RECT 810.600 759.600 812.400 764.400 ;
        RECT 821.100 759.600 822.900 765.600 ;
        RECT 825.000 762.600 826.500 772.950 ;
        RECT 830.550 769.050 831.450 781.950 ;
        RECT 842.400 776.100 843.600 785.400 ;
        RECT 841.950 774.450 844.050 775.050 ;
        RECT 846.000 774.450 850.050 775.050 ;
        RECT 841.950 773.550 850.050 774.450 ;
        RECT 841.950 772.950 844.050 773.550 ;
        RECT 846.000 772.950 850.050 773.550 ;
        RECT 839.100 770.100 840.900 770.850 ;
        RECT 829.950 766.950 832.050 769.050 ;
        RECT 838.950 766.950 841.050 769.050 ;
        RECT 842.400 762.600 843.600 771.900 ;
        RECT 825.000 759.600 826.800 762.600 ;
        RECT 842.400 759.600 844.200 762.600 ;
        RECT 12.000 748.200 13.800 755.400 ;
        RECT 22.950 751.950 25.050 754.050 ;
        RECT 12.000 747.300 15.600 748.200 ;
        RECT 14.400 743.100 15.600 747.300 ;
        RECT 11.100 740.100 12.900 740.850 ;
        RECT 13.950 739.950 16.050 742.050 ;
        RECT 17.100 740.100 18.900 740.850 ;
        RECT 10.950 736.950 13.050 739.050 ;
        RECT 14.400 729.600 15.600 738.900 ;
        RECT 16.950 736.950 19.050 739.050 ;
        RECT 23.550 730.050 24.450 751.950 ;
        RECT 28.800 749.400 30.600 755.400 ;
        RECT 29.400 747.300 30.600 749.400 ;
        RECT 31.800 750.300 33.600 755.400 ;
        RECT 37.800 750.300 39.600 755.400 ;
        RECT 31.800 748.950 39.600 750.300 ;
        RECT 47.400 750.300 49.200 755.400 ;
        RECT 53.400 750.300 55.200 755.400 ;
        RECT 47.400 748.950 55.200 750.300 ;
        RECT 56.400 749.400 58.200 755.400 ;
        RECT 75.000 751.050 76.800 755.400 ;
        RECT 85.950 751.950 88.050 754.050 ;
        RECT 56.400 747.300 57.600 749.400 ;
        RECT 64.950 748.950 67.050 751.050 ;
        RECT 71.400 749.400 76.800 751.050 ;
        RECT 29.400 746.250 33.150 747.300 ;
        RECT 31.950 746.100 33.150 746.250 ;
        RECT 53.850 746.250 57.600 747.300 ;
        RECT 53.850 746.100 55.050 746.250 ;
        RECT 29.100 743.100 30.900 743.850 ;
        RECT 31.950 742.950 34.050 745.050 ;
        RECT 35.100 743.100 36.900 743.850 ;
        RECT 37.950 742.950 40.050 745.050 ;
        RECT 46.950 742.950 49.050 745.050 ;
        RECT 50.100 743.100 51.900 743.850 ;
        RECT 52.950 742.950 55.200 745.050 ;
        RECT 56.100 743.100 57.900 743.850 ;
        RECT 28.950 739.950 31.050 742.050 ;
        RECT 32.850 738.900 33.900 741.900 ;
        RECT 34.950 739.950 37.200 742.050 ;
        RECT 38.100 741.150 39.900 741.900 ;
        RECT 47.100 741.150 48.900 741.900 ;
        RECT 49.950 739.950 52.050 742.050 ;
        RECT 53.100 738.900 54.150 741.900 ;
        RECT 55.950 739.950 58.050 742.050 ;
        RECT 32.850 735.600 34.050 738.900 ;
        RECT 52.950 735.600 54.150 738.900 ;
        RECT 13.800 723.600 15.600 729.600 ;
        RECT 22.950 727.950 25.050 730.050 ;
        RECT 32.700 723.600 34.500 735.600 ;
        RECT 52.500 723.600 54.300 735.600 ;
        RECT 65.550 730.050 66.450 748.950 ;
        RECT 71.400 746.100 72.300 749.400 ;
        RECT 67.950 742.950 73.050 745.050 ;
        RECT 74.100 743.100 75.900 743.850 ;
        RECT 76.950 742.950 79.050 745.050 ;
        RECT 80.100 743.100 81.900 743.850 ;
        RECT 71.400 735.600 72.300 741.900 ;
        RECT 73.950 739.950 76.050 742.050 ;
        RECT 77.100 741.150 78.900 741.900 ;
        RECT 79.950 739.950 82.050 742.050 ;
        RECT 64.950 727.950 67.050 730.050 ;
        RECT 70.800 723.600 72.600 735.600 ;
        RECT 73.800 734.700 81.600 735.600 ;
        RECT 73.800 723.600 75.600 734.700 ;
        RECT 79.800 723.600 81.600 734.700 ;
        RECT 86.550 730.050 87.450 751.950 ;
        RECT 95.100 747.000 96.900 755.400 ;
        RECT 115.200 748.200 117.000 755.400 ;
        RECT 92.700 745.350 96.900 747.000 ;
        RECT 113.400 747.300 117.000 748.200 ;
        RECT 131.400 752.400 133.200 755.400 ;
        RECT 92.700 740.100 93.600 745.350 ;
        RECT 95.100 743.100 96.900 743.850 ;
        RECT 101.100 743.100 102.900 743.850 ;
        RECT 113.400 743.100 114.600 747.300 ;
        RECT 127.950 745.950 130.050 748.050 ;
        RECT 128.100 744.150 129.900 744.900 ;
        RECT 131.400 743.100 132.600 752.400 ;
        RECT 149.100 747.000 150.900 755.400 ;
        RECT 169.200 748.200 171.000 755.400 ;
        RECT 177.000 753.450 181.050 754.050 ;
        RECT 167.400 747.300 171.000 748.200 ;
        RECT 176.550 751.950 181.050 753.450 ;
        RECT 185.400 752.400 187.200 755.400 ;
        RECT 176.550 748.050 177.450 751.950 ;
        RECT 186.300 748.200 187.200 752.400 ;
        RECT 191.400 749.400 193.200 755.400 ;
        RECT 149.100 745.350 153.300 747.000 ;
        RECT 143.100 743.100 144.900 743.850 ;
        RECT 149.100 743.100 150.900 743.850 ;
        RECT 94.950 739.950 97.050 742.050 ;
        RECT 100.950 739.950 103.050 742.050 ;
        RECT 110.100 740.100 111.900 740.850 ;
        RECT 112.950 739.950 115.050 742.050 ;
        RECT 116.100 740.100 117.900 740.850 ;
        RECT 130.950 739.950 136.050 742.050 ;
        RECT 142.800 739.950 145.050 742.050 ;
        RECT 148.950 739.950 151.200 742.050 ;
        RECT 152.400 740.100 153.300 745.350 ;
        RECT 167.400 743.100 168.600 747.300 ;
        RECT 175.950 745.950 178.050 748.050 ;
        RECT 181.950 745.950 184.050 748.050 ;
        RECT 186.300 747.300 189.750 748.200 ;
        RECT 187.950 746.400 189.750 747.300 ;
        RECT 164.100 740.100 165.900 740.850 ;
        RECT 166.950 739.950 169.050 742.050 ;
        RECT 170.100 740.100 171.900 740.850 ;
        RECT 176.550 739.050 177.450 745.950 ;
        RECT 182.100 744.150 183.900 744.900 ;
        RECT 184.950 742.950 187.050 745.050 ;
        RECT 185.100 741.150 186.900 741.900 ;
        RECT 88.950 736.950 94.050 739.050 ;
        RECT 97.800 736.950 100.050 739.050 ;
        RECT 109.950 736.950 112.050 739.050 ;
        RECT 92.700 730.800 93.600 735.900 ;
        RECT 98.100 735.150 99.900 735.900 ;
        RECT 103.950 733.950 106.050 736.050 ;
        RECT 85.950 727.950 88.050 730.050 ;
        RECT 92.700 729.900 99.300 730.800 ;
        RECT 104.550 730.050 105.450 733.950 ;
        RECT 92.700 729.600 93.600 729.900 ;
        RECT 91.800 723.600 93.600 729.600 ;
        RECT 97.800 729.600 99.300 729.900 ;
        RECT 97.800 723.600 99.600 729.600 ;
        RECT 103.950 727.950 106.050 730.050 ;
        RECT 113.400 729.600 114.600 738.900 ;
        RECT 115.950 736.950 118.050 739.050 ;
        RECT 131.400 729.600 132.600 738.900 ;
        RECT 145.950 736.950 148.050 739.050 ;
        RECT 151.950 736.950 154.050 739.050 ;
        RECT 163.950 736.950 166.050 739.050 ;
        RECT 146.100 735.150 147.900 735.900 ;
        RECT 152.400 730.800 153.300 735.900 ;
        RECT 146.700 729.900 153.300 730.800 ;
        RECT 146.700 729.600 148.200 729.900 ;
        RECT 113.400 723.600 115.200 729.600 ;
        RECT 131.400 723.600 133.200 729.600 ;
        RECT 146.400 723.600 148.200 729.600 ;
        RECT 152.400 729.600 153.300 729.900 ;
        RECT 167.400 729.600 168.600 738.900 ;
        RECT 169.950 736.950 172.050 739.050 ;
        RECT 175.950 736.950 178.050 739.050 ;
        RECT 188.700 738.600 189.600 746.400 ;
        RECT 192.000 743.100 193.050 749.400 ;
        RECT 202.950 748.950 205.050 751.050 ;
        RECT 203.550 745.050 204.450 748.950 ;
        RECT 207.000 748.200 208.800 755.400 ;
        RECT 226.800 752.400 228.600 755.400 ;
        RECT 227.400 749.100 228.600 752.400 ;
        RECT 243.000 748.200 244.800 755.400 ;
        RECT 260.400 752.400 262.200 755.400 ;
        RECT 207.000 747.300 210.600 748.200 ;
        RECT 202.950 742.950 205.050 745.050 ;
        RECT 209.400 743.100 210.600 747.300 ;
        RECT 226.950 745.950 229.050 748.050 ;
        RECT 243.000 747.300 246.600 748.200 ;
        RECT 223.950 742.950 226.050 745.050 ;
        RECT 190.950 739.950 193.050 742.050 ;
        RECT 206.100 740.100 207.900 740.850 ;
        RECT 208.950 739.950 211.050 742.050 ;
        RECT 227.100 741.900 228.300 744.900 ;
        RECT 229.950 742.950 232.050 745.050 ;
        RECT 245.400 743.100 246.600 747.300 ;
        RECT 256.950 745.950 259.050 748.050 ;
        RECT 257.100 744.150 258.900 744.900 ;
        RECT 260.400 743.100 261.600 752.400 ;
        RECT 278.100 747.000 279.900 755.400 ;
        RECT 295.800 749.400 297.600 755.400 ;
        RECT 301.800 752.400 303.600 755.400 ;
        RECT 275.700 745.350 279.900 747.000 ;
        RECT 224.100 741.150 225.900 741.900 ;
        RECT 212.100 740.100 213.900 740.850 ;
        RECT 187.800 738.000 189.600 738.600 ;
        RECT 182.400 736.800 189.600 738.000 ;
        RECT 182.400 735.600 183.600 736.800 ;
        RECT 188.700 736.650 189.600 736.800 ;
        RECT 190.950 735.600 192.300 738.900 ;
        RECT 205.950 736.950 208.050 739.050 ;
        RECT 152.400 723.600 154.200 729.600 ;
        RECT 167.400 723.600 169.200 729.600 ;
        RECT 182.400 723.600 184.200 735.600 ;
        RECT 189.900 734.100 192.300 735.600 ;
        RECT 189.900 723.600 191.700 734.100 ;
        RECT 209.400 729.600 210.600 738.900 ;
        RECT 211.950 736.950 214.050 739.050 ;
        RECT 226.950 736.650 228.300 741.900 ;
        RECT 230.100 741.150 231.900 741.900 ;
        RECT 242.100 740.100 243.900 740.850 ;
        RECT 244.950 739.950 247.050 742.050 ;
        RECT 248.100 740.100 249.900 740.850 ;
        RECT 259.950 739.950 265.050 742.050 ;
        RECT 275.700 740.100 276.600 745.350 ;
        RECT 278.100 743.100 279.900 743.850 ;
        RECT 284.100 743.100 285.900 743.850 ;
        RECT 295.950 743.100 297.000 749.400 ;
        RECT 301.800 748.200 302.700 752.400 ;
        RECT 319.200 748.200 321.000 755.400 ;
        RECT 335.400 752.400 337.200 755.400 ;
        RECT 335.400 749.100 336.600 752.400 ;
        RECT 352.800 749.400 354.600 755.400 ;
        RECT 299.250 747.300 302.700 748.200 ;
        RECT 299.250 746.400 301.050 747.300 ;
        RECT 277.950 739.950 280.050 742.050 ;
        RECT 283.950 739.950 286.050 742.050 ;
        RECT 295.950 741.450 298.050 742.050 ;
        RECT 290.550 740.550 298.050 741.450 ;
        RECT 241.950 736.950 244.050 739.050 ;
        RECT 208.800 723.600 210.600 729.600 ;
        RECT 225.600 735.600 228.300 736.650 ;
        RECT 225.600 723.600 227.400 735.600 ;
        RECT 245.400 729.600 246.600 738.900 ;
        RECT 247.950 736.950 250.050 739.050 ;
        RECT 244.800 723.600 246.600 729.600 ;
        RECT 260.400 729.600 261.600 738.900 ;
        RECT 271.950 736.950 277.050 739.050 ;
        RECT 280.950 736.950 283.200 739.050 ;
        RECT 290.550 736.050 291.450 740.550 ;
        RECT 295.950 739.950 298.050 740.550 ;
        RECT 275.700 730.800 276.600 735.900 ;
        RECT 281.100 735.150 282.900 735.900 ;
        RECT 289.950 733.950 292.050 736.050 ;
        RECT 296.700 735.600 298.050 738.900 ;
        RECT 299.400 738.600 300.300 746.400 ;
        RECT 304.950 745.950 307.050 748.050 ;
        RECT 317.400 747.300 321.000 748.200 ;
        RECT 301.950 742.950 304.050 745.050 ;
        RECT 305.100 744.150 306.900 744.900 ;
        RECT 317.400 743.100 318.600 747.300 ;
        RECT 334.950 745.950 337.050 748.050 ;
        RECT 353.400 747.300 354.600 749.400 ;
        RECT 355.800 750.300 357.600 755.400 ;
        RECT 361.800 750.300 363.600 755.400 ;
        RECT 355.800 748.950 363.600 750.300 ;
        RECT 374.400 752.400 376.200 755.400 ;
        RECT 353.400 746.250 357.150 747.300 ;
        RECT 355.950 746.100 357.150 746.250 ;
        RECT 370.950 745.950 373.050 748.050 ;
        RECT 331.800 742.950 334.050 745.050 ;
        RECT 302.100 741.150 303.900 741.900 ;
        RECT 314.100 740.100 315.900 740.850 ;
        RECT 316.950 739.950 319.050 742.050 ;
        RECT 335.700 741.900 336.900 744.900 ;
        RECT 337.800 742.950 340.050 745.050 ;
        RECT 353.100 743.100 354.900 743.850 ;
        RECT 355.800 742.950 358.050 745.050 ;
        RECT 359.100 743.100 360.900 743.850 ;
        RECT 361.950 742.950 364.200 745.050 ;
        RECT 371.100 744.150 372.900 744.900 ;
        RECT 374.400 743.100 375.600 752.400 ;
        RECT 379.950 751.950 382.050 754.050 ;
        RECT 388.800 752.400 390.600 755.400 ;
        RECT 332.100 741.150 333.900 741.900 ;
        RECT 320.100 740.100 321.900 740.850 ;
        RECT 299.400 738.000 301.200 738.600 ;
        RECT 299.400 736.800 306.600 738.000 ;
        RECT 313.950 736.950 316.050 739.050 ;
        RECT 299.400 736.650 300.300 736.800 ;
        RECT 305.400 735.600 306.600 736.800 ;
        RECT 296.700 734.100 299.100 735.600 ;
        RECT 275.700 729.900 282.300 730.800 ;
        RECT 275.700 729.600 276.600 729.900 ;
        RECT 260.400 723.600 262.200 729.600 ;
        RECT 274.800 723.600 276.600 729.600 ;
        RECT 280.800 729.600 282.300 729.900 ;
        RECT 280.800 723.600 282.600 729.600 ;
        RECT 297.300 723.600 299.100 734.100 ;
        RECT 304.800 723.600 306.600 735.600 ;
        RECT 317.400 729.600 318.600 738.900 ;
        RECT 319.950 736.950 322.050 739.050 ;
        RECT 335.700 736.650 337.050 741.900 ;
        RECT 338.100 741.150 339.900 741.900 ;
        RECT 352.950 739.950 355.050 742.050 ;
        RECT 356.850 738.900 357.900 741.900 ;
        RECT 358.950 739.950 361.050 742.050 ;
        RECT 362.100 741.150 363.900 741.900 ;
        RECT 373.950 741.450 376.050 742.050 ;
        RECT 380.550 741.450 381.450 751.950 ;
        RECT 389.400 743.100 390.600 752.400 ;
        RECT 404.400 752.400 406.200 755.400 ;
        RECT 391.950 745.950 394.050 751.050 ;
        RECT 404.400 749.100 405.600 752.400 ;
        RECT 424.200 748.200 426.000 755.400 ;
        RECT 439.800 749.400 441.600 755.400 ;
        RECT 403.950 745.950 406.050 748.050 ;
        RECT 422.400 747.300 426.000 748.200 ;
        RECT 440.400 747.300 441.600 749.400 ;
        RECT 442.800 750.300 444.600 755.400 ;
        RECT 448.800 750.300 450.600 755.400 ;
        RECT 442.800 748.950 450.600 750.300 ;
        RECT 463.200 748.200 465.000 755.400 ;
        RECT 478.800 749.400 480.600 755.400 ;
        RECT 461.400 747.300 465.000 748.200 ;
        RECT 479.400 747.300 480.600 749.400 ;
        RECT 481.800 750.300 483.600 755.400 ;
        RECT 487.800 750.300 489.600 755.400 ;
        RECT 499.800 752.400 501.600 755.400 ;
        RECT 481.800 748.950 489.600 750.300 ;
        RECT 392.100 744.150 393.900 744.900 ;
        RECT 400.950 742.950 403.200 745.050 ;
        RECT 373.950 740.550 381.450 741.450 ;
        RECT 388.950 741.450 391.050 742.050 ;
        RECT 393.000 741.450 397.050 742.050 ;
        RECT 404.700 741.900 405.900 744.900 ;
        RECT 406.950 742.950 409.200 745.050 ;
        RECT 422.400 743.100 423.600 747.300 ;
        RECT 440.400 746.250 444.150 747.300 ;
        RECT 442.950 746.100 444.150 746.250 ;
        RECT 440.100 743.100 441.900 743.850 ;
        RECT 442.800 742.950 445.050 745.050 ;
        RECT 446.100 743.100 447.900 743.850 ;
        RECT 448.950 742.950 451.050 745.050 ;
        RECT 461.400 743.100 462.600 747.300 ;
        RECT 479.400 746.250 483.150 747.300 ;
        RECT 481.950 746.100 483.150 746.250 ;
        RECT 479.100 743.100 480.900 743.850 ;
        RECT 481.950 742.950 484.050 745.050 ;
        RECT 485.100 743.100 486.900 743.850 ;
        RECT 487.950 742.950 490.200 745.050 ;
        RECT 500.400 743.100 501.600 752.400 ;
        RECT 514.800 754.500 522.600 755.400 ;
        RECT 514.800 749.400 516.600 754.500 ;
        RECT 517.800 749.400 519.600 753.600 ;
        RECT 520.800 750.000 522.600 754.500 ;
        RECT 526.800 750.000 528.600 755.400 ;
        RECT 502.950 745.950 505.050 748.050 ;
        RECT 518.400 747.900 519.300 749.400 ;
        RECT 520.800 749.100 528.600 750.000 ;
        RECT 541.200 748.200 543.000 755.400 ;
        RECT 559.800 749.400 561.600 755.400 ;
        RECT 575.400 752.400 577.200 755.400 ;
        RECT 593.400 752.400 595.200 755.400 ;
        RECT 515.700 746.100 517.500 746.850 ;
        RECT 518.400 746.700 522.600 747.900 ;
        RECT 539.400 747.300 543.000 748.200 ;
        RECT 521.400 746.100 522.600 746.700 ;
        RECT 526.950 746.100 528.750 746.850 ;
        RECT 503.100 744.150 504.900 744.900 ;
        RECT 514.950 742.950 517.050 745.050 ;
        RECT 518.250 743.100 519.900 743.850 ;
        RECT 520.950 742.950 523.050 745.050 ;
        RECT 524.100 743.100 525.900 743.850 ;
        RECT 526.950 742.950 529.050 745.050 ;
        RECT 539.400 743.100 540.600 747.300 ;
        RECT 559.950 743.100 561.300 749.400 ;
        RECT 575.400 749.100 576.600 752.400 ;
        RECT 593.400 749.100 594.600 752.400 ;
        RECT 601.950 751.950 604.050 754.050 ;
        RECT 574.950 745.950 577.050 748.050 ;
        RECT 592.950 745.950 595.050 748.050 ;
        RECT 602.550 745.050 603.450 751.950 ;
        RECT 610.800 749.400 612.600 755.400 ;
        RECT 611.400 747.300 612.600 749.400 ;
        RECT 613.800 750.300 615.600 755.400 ;
        RECT 619.800 750.300 621.600 755.400 ;
        RECT 613.800 748.950 621.600 750.300 ;
        RECT 632.400 752.400 634.200 755.400 ;
        RECT 646.800 752.400 648.600 755.400 ;
        RECT 611.400 746.250 615.150 747.300 ;
        RECT 613.950 746.100 615.150 746.250 ;
        RECT 628.950 745.950 631.200 748.050 ;
        RECT 563.100 743.100 564.900 743.850 ;
        RECT 388.950 740.550 397.050 741.450 ;
        RECT 401.100 741.150 402.900 741.900 ;
        RECT 373.950 739.950 376.050 740.550 ;
        RECT 388.950 739.950 391.050 740.550 ;
        RECT 393.000 739.950 397.050 740.550 ;
        RECT 335.700 735.600 338.400 736.650 ;
        RECT 356.850 735.600 358.050 738.900 ;
        RECT 317.400 723.600 319.200 729.600 ;
        RECT 336.600 723.600 338.400 735.600 ;
        RECT 356.700 723.600 358.500 735.600 ;
        RECT 374.400 729.600 375.600 738.900 ;
        RECT 389.400 729.600 390.600 738.900 ;
        RECT 404.700 736.650 406.050 741.900 ;
        RECT 407.100 741.150 408.900 741.900 ;
        RECT 419.100 740.100 420.900 740.850 ;
        RECT 421.950 739.950 424.050 742.050 ;
        RECT 425.100 740.100 426.900 740.850 ;
        RECT 430.950 739.950 433.050 742.050 ;
        RECT 439.950 739.950 442.050 742.050 ;
        RECT 418.950 736.950 421.050 739.050 ;
        RECT 404.700 735.600 407.400 736.650 ;
        RECT 374.400 723.600 376.200 729.600 ;
        RECT 388.800 723.600 390.600 729.600 ;
        RECT 405.600 723.600 407.400 735.600 ;
        RECT 422.400 729.600 423.600 738.900 ;
        RECT 424.950 736.950 427.050 739.050 ;
        RECT 431.550 730.050 432.450 739.950 ;
        RECT 443.850 738.900 444.900 741.900 ;
        RECT 445.950 739.950 448.050 742.050 ;
        RECT 449.100 741.150 450.900 741.900 ;
        RECT 458.100 740.100 459.900 740.850 ;
        RECT 460.950 739.950 463.050 742.050 ;
        RECT 464.100 740.100 465.900 740.850 ;
        RECT 478.950 739.950 481.050 742.050 ;
        RECT 443.850 735.600 445.050 738.900 ;
        RECT 457.950 736.950 460.050 739.050 ;
        RECT 422.400 723.600 424.200 729.600 ;
        RECT 430.950 727.950 433.050 730.050 ;
        RECT 443.700 723.600 445.500 735.600 ;
        RECT 461.400 729.600 462.600 738.900 ;
        RECT 463.950 736.950 466.050 739.050 ;
        RECT 482.850 738.900 483.900 741.900 ;
        RECT 484.950 739.950 487.050 742.050 ;
        RECT 488.100 741.150 489.900 741.900 ;
        RECT 499.950 741.450 502.050 742.050 ;
        RECT 504.000 741.450 508.050 742.050 ;
        RECT 499.950 740.550 508.050 741.450 ;
        RECT 499.950 739.950 502.050 740.550 ;
        RECT 504.000 739.950 508.050 740.550 ;
        RECT 517.950 739.950 520.050 742.050 ;
        RECT 482.850 735.600 484.050 738.900 ;
        RECT 461.400 723.600 463.200 729.600 ;
        RECT 482.700 723.600 484.500 735.600 ;
        RECT 500.400 729.600 501.600 738.900 ;
        RECT 521.400 735.600 522.600 741.900 ;
        RECT 523.950 739.950 526.050 742.050 ;
        RECT 536.100 740.100 537.900 740.850 ;
        RECT 538.950 739.950 541.050 742.050 ;
        RECT 542.100 740.100 543.900 740.850 ;
        RECT 556.950 739.950 559.050 742.050 ;
        RECT 535.950 736.950 538.050 739.050 ;
        RECT 499.800 723.600 501.600 729.600 ;
        RECT 520.800 723.600 524.100 735.600 ;
        RECT 539.400 729.600 540.600 738.900 ;
        RECT 541.950 736.950 544.050 739.050 ;
        RECT 560.100 738.900 561.300 743.100 ;
        RECT 571.950 742.950 574.050 745.050 ;
        RECT 562.950 739.950 568.050 742.050 ;
        RECT 575.700 741.900 576.900 744.900 ;
        RECT 577.950 742.950 580.050 745.050 ;
        RECT 589.950 742.950 592.050 745.050 ;
        RECT 593.700 741.900 594.900 744.900 ;
        RECT 595.950 742.950 598.050 745.050 ;
        RECT 601.950 742.950 604.050 745.050 ;
        RECT 611.100 743.100 612.900 743.850 ;
        RECT 613.950 742.950 616.050 745.050 ;
        RECT 617.100 743.100 618.900 743.850 ;
        RECT 619.950 742.950 622.200 745.050 ;
        RECT 629.100 744.150 630.900 744.900 ;
        RECT 632.400 743.100 633.600 752.400 ;
        RECT 647.400 743.100 648.600 752.400 ;
        RECT 662.400 752.400 664.200 755.400 ;
        RECT 680.400 752.400 682.200 755.400 ;
        RECT 662.400 749.100 663.600 752.400 ;
        RECT 680.400 749.100 681.600 752.400 ;
        RECT 699.000 748.200 700.800 755.400 ;
        RECT 707.550 749.400 709.350 755.400 ;
        RECT 715.650 752.400 717.450 755.400 ;
        RECT 723.450 752.400 725.250 755.400 ;
        RECT 731.250 753.300 733.050 755.400 ;
        RECT 731.250 752.400 735.000 753.300 ;
        RECT 715.650 751.500 716.700 752.400 ;
        RECT 712.950 750.300 716.700 751.500 ;
        RECT 724.200 750.600 725.250 752.400 ;
        RECT 733.950 751.500 735.000 752.400 ;
        RECT 712.950 749.400 715.050 750.300 ;
        RECT 649.950 745.950 652.050 748.050 ;
        RECT 661.950 745.950 664.200 748.050 ;
        RECT 679.950 745.950 682.200 748.050 ;
        RECT 699.000 747.300 702.600 748.200 ;
        RECT 650.100 744.150 651.900 744.900 ;
        RECT 658.950 742.950 661.050 745.050 ;
        RECT 572.100 741.150 573.900 741.900 ;
        RECT 559.950 735.600 561.300 738.900 ;
        RECT 575.700 736.650 577.050 741.900 ;
        RECT 578.100 741.150 579.900 741.900 ;
        RECT 590.100 741.150 591.900 741.900 ;
        RECT 593.700 736.650 595.050 741.900 ;
        RECT 596.100 741.150 597.900 741.900 ;
        RECT 575.700 735.600 578.400 736.650 ;
        RECT 593.700 735.600 596.400 736.650 ;
        RECT 539.400 723.600 541.200 729.600 ;
        RECT 559.800 723.600 561.600 735.600 ;
        RECT 576.600 723.600 578.400 735.600 ;
        RECT 594.600 723.600 596.400 735.600 ;
        RECT 602.550 730.050 603.450 742.950 ;
        RECT 610.950 739.950 613.050 742.050 ;
        RECT 614.850 738.900 615.900 741.900 ;
        RECT 616.950 739.950 619.050 742.050 ;
        RECT 620.100 741.150 621.900 741.900 ;
        RECT 631.950 741.450 634.050 742.050 ;
        RECT 631.950 740.550 639.450 741.450 ;
        RECT 631.950 739.950 634.050 740.550 ;
        RECT 614.850 735.600 616.050 738.900 ;
        RECT 601.950 727.950 604.050 730.050 ;
        RECT 614.700 723.600 616.500 735.600 ;
        RECT 632.400 729.600 633.600 738.900 ;
        RECT 638.550 733.050 639.450 740.550 ;
        RECT 646.950 739.950 649.050 742.050 ;
        RECT 662.700 741.900 663.900 744.900 ;
        RECT 664.950 742.950 667.050 745.050 ;
        RECT 676.950 742.950 679.200 745.050 ;
        RECT 680.700 741.900 681.900 744.900 ;
        RECT 682.950 742.950 685.050 745.050 ;
        RECT 691.950 742.950 694.050 745.050 ;
        RECT 701.400 743.100 702.600 747.300 ;
        RECT 707.550 745.050 708.750 749.400 ;
        RECT 720.150 748.200 721.950 750.000 ;
        RECT 724.200 749.550 729.150 750.600 ;
        RECT 727.350 748.800 729.150 749.550 ;
        RECT 730.650 748.800 732.450 750.600 ;
        RECT 733.950 749.400 736.050 751.500 ;
        RECT 739.050 749.400 740.850 755.400 ;
        RECT 721.050 747.900 721.950 748.200 ;
        RECT 731.100 747.900 732.150 748.800 ;
        RECT 721.050 747.000 732.150 747.900 ;
        RECT 721.050 746.100 721.950 747.000 ;
        RECT 731.100 745.800 732.150 747.000 ;
        RECT 707.550 742.950 708.900 745.050 ;
        RECT 709.950 742.950 712.050 745.050 ;
        RECT 713.100 743.250 713.850 745.050 ;
        RECT 721.950 742.950 724.050 745.050 ;
        RECT 727.950 742.950 730.050 745.050 ;
        RECT 731.100 744.600 738.000 745.800 ;
        RECT 731.100 744.000 732.900 744.600 ;
        RECT 737.100 743.850 738.000 744.600 ;
        RECT 734.100 743.100 735.900 743.700 ;
        RECT 659.100 741.150 660.900 741.900 ;
        RECT 637.950 730.950 640.050 733.050 ;
        RECT 647.400 729.600 648.600 738.900 ;
        RECT 662.700 736.650 664.050 741.900 ;
        RECT 665.100 741.150 666.900 741.900 ;
        RECT 677.100 741.150 678.900 741.900 ;
        RECT 680.700 736.650 682.050 741.900 ;
        RECT 683.100 741.150 684.900 741.900 ;
        RECT 662.700 735.600 665.400 736.650 ;
        RECT 632.400 723.600 634.200 729.600 ;
        RECT 646.800 723.600 648.600 729.600 ;
        RECT 663.600 723.600 665.400 735.600 ;
        RECT 670.950 733.950 673.050 736.050 ;
        RECT 680.700 735.600 683.400 736.650 ;
        RECT 692.550 736.050 693.450 742.950 ;
        RECT 698.100 740.100 699.900 740.850 ;
        RECT 700.950 739.950 703.050 742.050 ;
        RECT 704.100 740.100 705.900 740.850 ;
        RECT 697.950 736.950 700.050 739.050 ;
        RECT 671.550 730.050 672.450 733.950 ;
        RECT 670.950 727.950 673.050 730.050 ;
        RECT 681.600 723.600 683.400 735.600 ;
        RECT 691.950 733.950 694.050 736.050 ;
        RECT 701.400 729.600 702.600 738.900 ;
        RECT 703.950 736.950 706.050 739.050 ;
        RECT 700.800 723.600 702.600 729.600 ;
        RECT 707.550 735.600 708.750 742.950 ;
        RECT 731.100 742.200 735.900 743.100 ;
        RECT 734.100 741.900 735.900 742.200 ;
        RECT 737.100 742.050 738.900 743.850 ;
        RECT 709.950 737.400 711.750 739.200 ;
        RECT 710.850 736.200 715.050 737.400 ;
        RECT 721.050 736.200 721.950 741.900 ;
        RECT 729.750 737.100 731.550 737.400 ;
        RECT 707.550 723.600 709.350 735.600 ;
        RECT 712.950 735.300 715.050 736.200 ;
        RECT 715.950 735.300 721.950 736.200 ;
        RECT 723.150 736.800 731.550 737.100 ;
        RECT 739.950 736.800 740.850 749.400 ;
        RECT 754.200 748.200 756.000 755.400 ;
        RECT 769.800 749.400 771.600 755.400 ;
        RECT 752.400 747.300 756.000 748.200 ;
        RECT 770.400 747.300 771.600 749.400 ;
        RECT 772.800 750.300 774.600 755.400 ;
        RECT 778.800 750.300 780.600 755.400 ;
        RECT 790.800 752.400 792.600 755.400 ;
        RECT 803.400 752.400 805.200 755.400 ;
        RECT 772.800 748.950 780.600 750.300 ;
        RECT 752.400 743.100 753.600 747.300 ;
        RECT 770.400 746.250 774.150 747.300 ;
        RECT 772.950 746.100 774.150 746.250 ;
        RECT 770.100 743.100 771.900 743.850 ;
        RECT 772.950 742.950 775.050 745.050 ;
        RECT 776.100 743.100 777.900 743.850 ;
        RECT 778.950 742.950 781.050 745.050 ;
        RECT 791.400 743.100 792.600 752.400 ;
        RECT 804.000 748.500 805.200 752.400 ;
        RECT 809.700 749.400 811.500 755.400 ;
        RECT 821.400 750.300 823.200 755.400 ;
        RECT 827.400 750.300 829.200 755.400 ;
        RECT 804.000 747.600 809.100 748.500 ;
        RECT 807.150 746.700 809.100 747.600 ;
        RECT 807.150 746.100 808.050 746.700 ;
        RECT 810.000 746.100 811.200 749.400 ;
        RECT 821.400 748.950 829.200 750.300 ;
        RECT 830.400 749.400 832.200 755.400 ;
        RECT 830.400 747.300 831.600 749.400 ;
        RECT 847.200 748.200 849.000 755.400 ;
        RECT 827.850 746.250 831.600 747.300 ;
        RECT 845.400 747.300 849.000 748.200 ;
        RECT 827.850 746.100 829.050 746.250 ;
        RECT 794.100 744.150 795.900 744.900 ;
        RECT 799.950 742.950 805.050 745.050 ;
        RECT 749.100 740.100 750.900 740.850 ;
        RECT 751.950 739.950 754.050 742.050 ;
        RECT 755.100 740.100 756.900 740.850 ;
        RECT 769.950 739.950 772.050 742.050 ;
        RECT 742.950 736.950 745.050 739.050 ;
        RECT 748.950 736.950 751.050 739.050 ;
        RECT 723.150 736.200 740.850 736.800 ;
        RECT 715.950 734.400 716.850 735.300 ;
        RECT 714.150 732.600 716.850 734.400 ;
        RECT 717.750 734.100 719.550 734.400 ;
        RECT 723.150 734.100 724.050 736.200 ;
        RECT 729.750 735.600 740.850 736.200 ;
        RECT 717.750 733.200 724.050 734.100 ;
        RECT 724.950 734.700 726.750 735.300 ;
        RECT 724.950 733.500 732.450 734.700 ;
        RECT 717.750 732.600 719.550 733.200 ;
        RECT 731.250 732.600 732.450 733.500 ;
        RECT 712.950 729.600 716.850 731.700 ;
        RECT 721.950 731.550 723.750 732.300 ;
        RECT 726.750 731.550 728.550 732.300 ;
        RECT 721.950 730.500 728.550 731.550 ;
        RECT 731.250 730.500 736.050 732.600 ;
        RECT 715.050 723.600 716.850 729.600 ;
        RECT 722.850 723.600 724.650 730.500 ;
        RECT 731.250 729.600 732.450 730.500 ;
        RECT 730.650 723.600 732.450 729.600 ;
        RECT 739.050 723.600 740.850 735.600 ;
        RECT 743.550 727.050 744.450 736.950 ;
        RECT 752.400 729.600 753.600 738.900 ;
        RECT 754.950 736.950 757.050 739.050 ;
        RECT 773.850 738.900 774.900 741.900 ;
        RECT 775.800 739.950 778.050 742.050 ;
        RECT 779.100 741.150 780.900 741.900 ;
        RECT 790.950 739.950 793.050 742.050 ;
        RECT 807.150 741.900 807.900 746.100 ;
        RECT 808.950 742.950 811.050 745.050 ;
        RECT 820.950 744.450 823.050 745.050 ;
        RECT 815.550 743.550 823.050 744.450 ;
        RECT 803.100 741.150 804.900 741.900 ;
        RECT 773.850 735.600 775.050 738.900 ;
        RECT 742.950 724.950 745.050 727.050 ;
        RECT 752.400 723.600 754.200 729.600 ;
        RECT 773.700 723.600 775.500 735.600 ;
        RECT 791.400 729.600 792.600 738.900 ;
        RECT 807.150 738.300 808.050 741.900 ;
        RECT 807.150 737.400 809.100 738.300 ;
        RECT 790.800 723.600 792.600 729.600 ;
        RECT 803.400 736.500 809.100 737.400 ;
        RECT 803.400 729.600 804.600 736.500 ;
        RECT 810.000 735.600 811.200 741.900 ;
        RECT 803.400 723.600 805.200 729.600 ;
        RECT 809.700 723.600 811.500 735.600 ;
        RECT 815.550 727.050 816.450 743.550 ;
        RECT 820.950 742.950 823.050 743.550 ;
        RECT 824.100 743.100 825.900 743.850 ;
        RECT 826.950 742.950 829.050 745.050 ;
        RECT 830.100 743.100 831.900 743.850 ;
        RECT 845.400 743.100 846.600 747.300 ;
        RECT 821.100 741.150 822.900 741.900 ;
        RECT 823.950 739.950 826.200 742.050 ;
        RECT 827.100 738.900 828.150 741.900 ;
        RECT 829.950 739.950 832.050 742.050 ;
        RECT 842.100 740.100 843.900 740.850 ;
        RECT 844.950 739.950 847.050 742.050 ;
        RECT 848.100 740.100 849.900 740.850 ;
        RECT 826.950 735.600 828.150 738.900 ;
        RECT 841.950 736.950 844.050 739.050 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 826.500 723.600 828.300 735.600 ;
        RECT 845.400 729.600 846.600 738.900 ;
        RECT 847.950 736.950 850.050 739.050 ;
        RECT 845.400 723.600 847.200 729.600 ;
        RECT 10.800 713.400 12.600 719.400 ;
        RECT 11.700 713.100 12.600 713.400 ;
        RECT 16.800 713.400 18.600 719.400 ;
        RECT 16.800 713.100 18.300 713.400 ;
        RECT 11.700 712.200 18.300 713.100 ;
        RECT 11.700 707.100 12.600 712.200 ;
        RECT 29.400 708.300 31.200 719.400 ;
        RECT 35.400 708.300 37.200 719.400 ;
        RECT 17.100 707.100 18.900 707.850 ;
        RECT 29.400 707.400 37.200 708.300 ;
        RECT 38.400 707.400 40.200 719.400 ;
        RECT 55.500 707.400 57.300 719.400 ;
        RECT 58.950 709.950 61.050 712.050 ;
        RECT 10.950 705.450 13.050 706.050 ;
        RECT 5.550 704.550 13.050 705.450 ;
        RECT 5.550 697.050 6.450 704.550 ;
        RECT 10.950 703.950 13.050 704.550 ;
        RECT 16.950 703.950 19.050 706.050 ;
        RECT 11.700 697.650 12.600 702.900 ;
        RECT 13.950 700.950 16.050 703.050 ;
        RECT 19.950 700.950 22.050 703.050 ;
        RECT 28.800 700.950 31.050 703.050 ;
        RECT 32.100 701.100 33.900 701.850 ;
        RECT 34.950 700.950 37.050 703.050 ;
        RECT 38.700 701.100 39.600 707.400 ;
        RECT 55.950 704.100 57.150 707.400 ;
        RECT 50.100 701.100 51.900 701.850 ;
        RECT 52.950 700.950 55.050 703.050 ;
        RECT 56.100 701.100 57.150 704.100 ;
        RECT 59.550 703.050 60.450 709.950 ;
        RECT 76.500 707.400 78.300 719.400 ;
        RECT 95.400 713.400 97.200 719.400 ;
        RECT 95.700 713.100 97.200 713.400 ;
        RECT 101.400 713.400 103.200 719.400 ;
        RECT 116.400 713.400 118.200 719.400 ;
        RECT 101.400 713.100 102.300 713.400 ;
        RECT 95.700 712.200 102.300 713.100 ;
        RECT 116.700 713.100 118.200 713.400 ;
        RECT 122.400 713.400 124.200 719.400 ;
        RECT 122.400 713.100 123.300 713.400 ;
        RECT 116.700 712.200 123.300 713.100 ;
        RECT 76.950 704.100 78.150 707.400 ;
        RECT 95.100 707.100 96.900 707.850 ;
        RECT 101.400 707.100 102.300 712.200 ;
        RECT 116.100 707.100 117.900 707.850 ;
        RECT 122.400 707.100 123.300 712.200 ;
        RECT 134.400 708.300 136.200 719.400 ;
        RECT 140.400 708.300 142.200 719.400 ;
        RECT 134.400 707.400 142.200 708.300 ;
        RECT 143.400 707.400 145.200 719.400 ;
        RECT 160.500 707.400 162.300 719.400 ;
        RECT 181.800 713.400 183.600 719.400 ;
        RECT 197.400 713.400 199.200 719.400 ;
        RECT 58.950 700.950 61.200 703.050 ;
        RECT 71.100 701.100 72.900 701.850 ;
        RECT 73.950 700.950 76.050 703.050 ;
        RECT 77.100 701.100 78.150 704.100 ;
        RECT 94.950 703.950 97.200 706.050 ;
        RECT 100.950 705.450 103.050 706.050 ;
        RECT 100.950 704.550 108.450 705.450 ;
        RECT 100.950 703.950 103.050 704.550 ;
        RECT 79.950 700.950 82.050 703.050 ;
        RECT 91.950 700.950 94.050 703.050 ;
        RECT 97.950 700.950 100.050 703.050 ;
        RECT 14.100 699.150 15.900 699.900 ;
        RECT 20.100 699.150 21.900 699.900 ;
        RECT 29.100 699.150 30.900 699.900 ;
        RECT 31.950 697.950 34.050 700.050 ;
        RECT 35.100 699.150 36.900 699.900 ;
        RECT 37.950 697.950 43.050 700.050 ;
        RECT 49.950 697.950 52.050 700.050 ;
        RECT 53.100 699.150 54.900 699.900 ;
        RECT 55.950 697.950 58.050 700.050 ;
        RECT 59.100 699.150 60.900 699.900 ;
        RECT 70.950 697.950 73.050 700.050 ;
        RECT 74.100 699.150 75.900 699.900 ;
        RECT 76.950 697.950 79.050 700.050 ;
        RECT 80.100 699.150 81.900 699.900 ;
        RECT 92.100 699.150 93.900 699.900 ;
        RECT 98.100 699.150 99.900 699.900 ;
        RECT 101.400 697.650 102.300 702.900 ;
        RECT 4.950 694.950 7.050 697.050 ;
        RECT 11.700 696.000 15.900 697.650 ;
        RECT 14.100 687.600 15.900 696.000 ;
        RECT 38.700 693.600 39.600 696.900 ;
        RECT 56.850 696.750 58.050 696.900 ;
        RECT 77.850 696.750 79.050 696.900 ;
        RECT 56.850 695.700 60.600 696.750 ;
        RECT 77.850 695.700 81.600 696.750 ;
        RECT 34.200 691.950 39.600 693.600 ;
        RECT 50.400 692.700 58.200 694.050 ;
        RECT 34.200 687.600 36.000 691.950 ;
        RECT 50.400 687.600 52.200 692.700 ;
        RECT 56.400 687.600 58.200 692.700 ;
        RECT 59.400 693.600 60.600 695.700 ;
        RECT 59.400 687.600 61.200 693.600 ;
        RECT 71.400 692.700 79.200 694.050 ;
        RECT 71.400 687.600 73.200 692.700 ;
        RECT 77.400 687.600 79.200 692.700 ;
        RECT 80.400 693.600 81.600 695.700 ;
        RECT 98.100 696.000 102.300 697.650 ;
        RECT 80.400 687.600 82.200 693.600 ;
        RECT 98.100 687.600 99.900 696.000 ;
        RECT 107.550 691.050 108.450 704.550 ;
        RECT 115.950 703.950 118.050 706.050 ;
        RECT 121.950 705.450 124.050 706.050 ;
        RECT 121.950 704.550 129.450 705.450 ;
        RECT 121.950 703.950 124.050 704.550 ;
        RECT 112.950 700.950 115.050 703.050 ;
        RECT 118.950 700.950 121.050 703.050 ;
        RECT 113.100 699.150 114.900 699.900 ;
        RECT 119.100 699.150 120.900 699.900 ;
        RECT 122.400 697.650 123.300 702.900 ;
        RECT 119.100 696.000 123.300 697.650 ;
        RECT 106.950 688.950 109.050 691.050 ;
        RECT 119.100 687.600 120.900 696.000 ;
        RECT 128.550 691.050 129.450 704.550 ;
        RECT 133.950 700.950 136.050 703.050 ;
        RECT 137.100 701.100 138.900 701.850 ;
        RECT 139.950 700.950 142.050 703.050 ;
        RECT 143.700 701.100 144.600 707.400 ;
        RECT 148.950 703.950 151.050 706.050 ;
        RECT 160.950 704.100 162.150 707.400 ;
        RECT 134.100 699.150 135.900 699.900 ;
        RECT 136.800 697.950 139.050 700.050 ;
        RECT 140.100 699.150 141.900 699.900 ;
        RECT 142.950 699.450 145.050 700.050 ;
        RECT 149.550 699.450 150.450 703.950 ;
        RECT 155.100 701.100 156.900 701.850 ;
        RECT 157.950 700.950 160.050 703.050 ;
        RECT 161.100 701.100 162.150 704.100 ;
        RECT 178.950 703.950 181.050 706.050 ;
        RECT 182.400 704.100 183.600 713.400 ;
        RECT 197.700 713.100 199.200 713.400 ;
        RECT 203.400 713.400 205.200 719.400 ;
        RECT 203.400 713.100 204.300 713.400 ;
        RECT 197.700 712.200 204.300 713.100 ;
        RECT 197.100 707.100 198.900 707.850 ;
        RECT 203.400 707.100 204.300 712.200 ;
        RECT 219.600 707.400 221.400 719.400 ;
        RECT 235.800 713.400 237.600 719.400 ;
        RECT 236.700 713.100 237.600 713.400 ;
        RECT 241.800 713.400 243.600 719.400 ;
        RECT 241.800 713.100 243.300 713.400 ;
        RECT 236.700 712.200 243.300 713.100 ;
        RECT 219.600 706.350 222.300 707.400 ;
        RECT 236.700 707.100 237.600 712.200 ;
        RECT 242.100 707.100 243.900 707.850 ;
        RECT 258.900 707.400 262.200 719.400 ;
        RECT 280.800 713.400 282.600 719.400 ;
        RECT 281.700 713.100 282.600 713.400 ;
        RECT 286.800 713.400 288.600 719.400 ;
        RECT 286.800 713.100 288.300 713.400 ;
        RECT 281.700 712.200 288.300 713.100 ;
        RECT 184.950 703.950 187.050 706.050 ;
        RECT 196.950 703.950 199.050 706.050 ;
        RECT 202.950 705.450 205.050 706.050 ;
        RECT 202.950 704.550 210.450 705.450 ;
        RECT 202.950 703.950 205.050 704.550 ;
        RECT 163.950 700.950 166.050 703.050 ;
        RECT 179.100 702.150 180.900 702.900 ;
        RECT 181.950 700.950 184.050 703.050 ;
        RECT 185.100 702.150 186.900 702.900 ;
        RECT 193.950 700.950 196.050 703.050 ;
        RECT 199.950 700.950 202.050 703.050 ;
        RECT 142.950 698.550 150.450 699.450 ;
        RECT 142.950 697.950 145.050 698.550 ;
        RECT 154.950 697.950 157.050 700.050 ;
        RECT 158.100 699.150 159.900 699.900 ;
        RECT 160.950 697.950 163.050 700.050 ;
        RECT 164.100 699.150 165.900 699.900 ;
        RECT 143.700 693.600 144.600 696.900 ;
        RECT 161.850 696.750 163.050 696.900 ;
        RECT 161.850 695.700 165.600 696.750 ;
        RECT 182.400 695.700 183.600 699.900 ;
        RECT 194.100 699.150 195.900 699.900 ;
        RECT 200.100 699.150 201.900 699.900 ;
        RECT 203.400 697.650 204.300 702.900 ;
        RECT 139.200 691.950 144.600 693.600 ;
        RECT 155.400 692.700 163.200 694.050 ;
        RECT 127.950 688.950 130.050 691.050 ;
        RECT 139.200 687.600 141.000 691.950 ;
        RECT 155.400 687.600 157.200 692.700 ;
        RECT 161.400 687.600 163.200 692.700 ;
        RECT 164.400 693.600 165.600 695.700 ;
        RECT 180.000 694.800 183.600 695.700 ;
        RECT 200.100 696.000 204.300 697.650 ;
        RECT 164.400 687.600 166.200 693.600 ;
        RECT 180.000 687.600 181.800 694.800 ;
        RECT 200.100 687.600 201.900 696.000 ;
        RECT 209.550 691.050 210.450 704.550 ;
        RECT 218.100 701.100 219.900 701.850 ;
        RECT 220.950 701.100 222.300 706.350 ;
        RECT 232.950 703.950 238.050 706.050 ;
        RECT 241.950 703.950 244.200 706.050 ;
        RECT 224.100 701.100 225.900 701.850 ;
        RECT 217.950 697.950 220.050 700.050 ;
        RECT 221.100 698.100 222.300 701.100 ;
        RECT 223.950 697.950 226.050 700.050 ;
        RECT 236.700 697.650 237.600 702.900 ;
        RECT 238.950 700.950 241.050 703.050 ;
        RECT 244.950 700.950 247.050 703.050 ;
        RECT 256.950 700.950 259.050 703.050 ;
        RECT 260.400 701.100 261.600 707.400 ;
        RECT 281.700 707.100 282.600 712.200 ;
        RECT 287.100 707.100 288.900 707.850 ;
        RECT 301.800 707.400 303.600 719.400 ;
        RECT 304.800 708.300 306.600 719.400 ;
        RECT 310.800 708.300 312.600 719.400 ;
        RECT 304.800 707.400 312.600 708.300 ;
        RECT 323.400 713.400 325.200 719.400 ;
        RECT 338.400 713.400 340.200 719.400 ;
        RECT 277.950 703.950 283.050 706.050 ;
        RECT 286.950 703.950 289.050 706.050 ;
        RECT 262.950 700.950 265.050 703.050 ;
        RECT 239.100 699.150 240.900 699.900 ;
        RECT 245.100 699.150 246.900 699.900 ;
        RECT 253.800 697.950 256.050 700.050 ;
        RECT 257.100 699.150 258.900 699.900 ;
        RECT 259.950 697.950 262.200 700.050 ;
        RECT 263.100 699.150 264.750 699.900 ;
        RECT 265.950 697.950 268.200 700.050 ;
        RECT 281.700 697.650 282.600 702.900 ;
        RECT 283.950 700.950 286.050 703.050 ;
        RECT 289.950 700.950 292.200 703.050 ;
        RECT 302.400 701.100 303.300 707.400 ;
        RECT 323.400 704.100 324.600 713.400 ;
        RECT 331.950 706.950 334.050 709.050 ;
        RECT 304.950 700.950 307.050 703.050 ;
        RECT 308.100 701.100 309.900 701.850 ;
        RECT 310.950 700.950 313.050 703.050 ;
        RECT 319.950 700.950 325.050 703.050 ;
        RECT 332.550 702.450 333.450 706.950 ;
        RECT 338.400 704.100 339.600 713.400 ;
        RECT 355.500 707.400 357.300 719.400 ;
        RECT 373.800 707.400 375.600 719.400 ;
        RECT 355.950 704.100 357.150 707.400 ;
        RECT 337.950 702.450 340.050 703.050 ;
        RECT 332.550 701.550 340.050 702.450 ;
        RECT 337.950 700.950 340.050 701.550 ;
        RECT 350.100 701.100 351.900 701.850 ;
        RECT 352.950 700.950 355.050 703.050 ;
        RECT 356.100 701.100 357.150 704.100 ;
        RECT 358.950 700.950 361.050 703.050 ;
        RECT 374.400 701.100 375.600 707.400 ;
        RECT 389.400 713.400 391.200 719.400 ;
        RECT 397.950 715.950 400.050 718.050 ;
        RECT 385.950 703.950 388.050 706.050 ;
        RECT 389.400 704.100 390.600 713.400 ;
        RECT 391.950 708.000 394.050 712.050 ;
        RECT 392.550 706.050 393.450 708.000 ;
        RECT 391.950 703.950 394.050 706.050 ;
        RECT 376.950 700.950 379.050 703.050 ;
        RECT 386.100 702.150 387.900 702.900 ;
        RECT 388.800 700.950 391.050 703.050 ;
        RECT 392.100 702.150 393.900 702.900 ;
        RECT 398.550 700.050 399.450 715.950 ;
        RECT 412.800 707.400 416.100 719.400 ;
        RECT 433.800 713.400 435.600 719.400 ;
        RECT 409.950 700.950 412.050 703.050 ;
        RECT 413.400 701.100 414.600 707.400 ;
        RECT 430.950 703.950 433.050 709.050 ;
        RECT 434.400 704.100 435.600 713.400 ;
        RECT 446.400 707.400 448.200 719.400 ;
        RECT 453.900 708.900 455.700 719.400 ;
        RECT 469.800 713.400 471.600 719.400 ;
        RECT 485.400 713.400 487.200 719.400 ;
        RECT 453.900 707.400 456.300 708.900 ;
        RECT 446.400 706.200 447.600 707.400 ;
        RECT 452.700 706.200 453.600 706.350 ;
        RECT 436.950 703.950 439.050 706.050 ;
        RECT 446.400 705.000 453.600 706.200 ;
        RECT 451.800 704.400 453.600 705.000 ;
        RECT 415.950 700.950 418.050 703.050 ;
        RECT 431.100 702.150 432.900 702.900 ;
        RECT 433.950 700.950 436.050 703.050 ;
        RECT 437.100 702.150 438.900 702.900 ;
        RECT 449.100 701.100 450.900 701.850 ;
        RECT 284.100 699.150 285.900 699.900 ;
        RECT 290.100 699.150 291.900 699.900 ;
        RECT 298.800 697.950 304.050 700.050 ;
        RECT 305.100 699.150 306.900 699.900 ;
        RECT 307.800 697.950 310.050 700.050 ;
        RECT 311.100 699.150 312.900 699.900 ;
        RECT 320.100 698.100 321.900 698.850 ;
        RECT 220.800 694.950 223.050 697.050 ;
        RECT 236.700 696.000 240.900 697.650 ;
        RECT 254.250 696.150 256.050 696.900 ;
        RECT 260.400 696.300 261.600 696.900 ;
        RECT 208.950 688.950 211.050 691.050 ;
        RECT 221.400 690.600 222.600 693.900 ;
        RECT 220.800 687.600 222.600 690.600 ;
        RECT 239.100 687.600 240.900 696.000 ;
        RECT 260.400 695.100 264.600 696.300 ;
        RECT 265.500 696.150 267.300 696.900 ;
        RECT 281.700 696.000 285.900 697.650 ;
        RECT 254.400 693.000 262.200 693.900 ;
        RECT 263.700 693.600 264.600 695.100 ;
        RECT 254.400 687.600 256.200 693.000 ;
        RECT 260.400 688.500 262.200 693.000 ;
        RECT 263.400 689.400 265.200 693.600 ;
        RECT 266.400 688.500 268.200 693.600 ;
        RECT 260.400 687.600 268.200 688.500 ;
        RECT 284.100 687.600 285.900 696.000 ;
        RECT 302.400 693.600 303.300 696.900 ;
        RECT 319.950 694.950 322.050 697.050 ;
        RECT 302.400 691.950 307.800 693.600 ;
        RECT 306.000 687.600 307.800 691.950 ;
        RECT 323.400 690.600 324.600 699.900 ;
        RECT 335.100 698.100 336.900 698.850 ;
        RECT 334.950 694.950 337.050 697.050 ;
        RECT 338.400 690.600 339.600 699.900 ;
        RECT 349.800 697.950 352.050 700.050 ;
        RECT 353.100 699.150 354.900 699.900 ;
        RECT 355.950 697.950 358.200 700.050 ;
        RECT 359.100 699.150 360.900 699.900 ;
        RECT 373.950 697.950 376.050 700.050 ;
        RECT 377.100 699.150 378.900 699.900 ;
        RECT 356.850 696.750 358.050 696.900 ;
        RECT 356.850 695.700 360.600 696.750 ;
        RECT 350.400 692.700 358.200 694.050 ;
        RECT 323.400 687.600 325.200 690.600 ;
        RECT 338.400 687.600 340.200 690.600 ;
        RECT 350.400 687.600 352.200 692.700 ;
        RECT 356.400 687.600 358.200 692.700 ;
        RECT 359.400 693.600 360.600 695.700 ;
        RECT 374.400 693.600 375.600 696.900 ;
        RECT 389.400 695.700 390.600 699.900 ;
        RECT 397.950 697.950 400.050 700.050 ;
        RECT 406.950 697.950 409.050 700.050 ;
        RECT 410.250 699.150 411.900 699.900 ;
        RECT 412.800 697.950 415.050 700.050 ;
        RECT 416.100 699.150 417.900 699.900 ;
        RECT 418.950 697.950 421.050 700.050 ;
        RECT 407.700 696.150 409.500 696.900 ;
        RECT 413.400 696.300 414.600 696.900 ;
        RECT 389.400 694.800 393.000 695.700 ;
        RECT 359.400 687.600 361.200 693.600 ;
        RECT 373.800 687.600 375.600 693.600 ;
        RECT 391.200 687.600 393.000 694.800 ;
        RECT 410.400 695.100 414.600 696.300 ;
        RECT 418.950 696.150 420.750 696.900 ;
        RECT 434.400 695.700 435.600 699.900 ;
        RECT 446.100 698.100 447.900 698.850 ;
        RECT 448.950 697.950 451.050 700.050 ;
        RECT 410.400 693.600 411.300 695.100 ;
        RECT 432.000 694.800 435.600 695.700 ;
        RECT 445.950 694.950 448.050 697.050 ;
        RECT 452.700 696.600 453.600 704.400 ;
        RECT 454.950 704.100 456.300 707.400 ;
        RECT 470.400 704.100 471.600 713.400 ;
        RECT 485.700 713.100 487.200 713.400 ;
        RECT 491.400 713.400 493.200 719.400 ;
        RECT 506.400 713.400 508.200 719.400 ;
        RECT 491.400 713.100 492.300 713.400 ;
        RECT 485.700 712.200 492.300 713.100 ;
        RECT 485.100 707.100 486.900 707.850 ;
        RECT 491.400 707.100 492.300 712.200 ;
        RECT 484.950 703.950 487.050 706.050 ;
        RECT 490.950 703.950 495.900 706.050 ;
        RECT 502.950 703.950 505.050 706.050 ;
        RECT 506.400 704.100 507.600 713.400 ;
        RECT 523.800 707.400 525.600 719.400 ;
        RECT 508.950 703.950 511.050 706.050 ;
        RECT 454.950 700.950 460.050 703.050 ;
        RECT 469.950 700.950 475.050 703.050 ;
        RECT 481.950 700.950 484.050 703.050 ;
        RECT 487.950 700.950 490.050 703.050 ;
        RECT 451.950 695.700 453.750 696.600 ;
        RECT 450.300 694.800 453.750 695.700 ;
        RECT 406.800 688.500 408.600 693.600 ;
        RECT 409.800 689.400 411.600 693.600 ;
        RECT 412.800 693.000 420.600 693.900 ;
        RECT 412.800 688.500 414.600 693.000 ;
        RECT 406.800 687.600 414.600 688.500 ;
        RECT 418.800 687.600 420.600 693.000 ;
        RECT 432.000 687.600 433.800 694.800 ;
        RECT 450.300 690.600 451.200 694.800 ;
        RECT 456.000 693.600 457.050 699.900 ;
        RECT 449.400 687.600 451.200 690.600 ;
        RECT 455.400 687.600 457.200 693.600 ;
        RECT 470.400 690.600 471.600 699.900 ;
        RECT 482.100 699.150 483.900 699.900 ;
        RECT 488.100 699.150 489.900 699.900 ;
        RECT 473.100 698.100 474.900 698.850 ;
        RECT 491.400 697.650 492.300 702.900 ;
        RECT 503.100 702.150 504.900 702.900 ;
        RECT 505.950 700.950 508.050 703.050 ;
        RECT 509.100 702.150 510.900 702.900 ;
        RECT 524.400 701.100 525.600 707.400 ;
        RECT 539.400 713.400 541.200 719.400 ;
        RECT 539.400 704.100 540.600 713.400 ;
        RECT 555.600 707.400 557.400 719.400 ;
        RECT 574.800 713.400 576.600 719.400 ;
        RECT 554.700 706.350 557.400 707.400 ;
        RECT 565.950 706.950 568.050 709.050 ;
        RECT 526.950 700.950 529.050 703.050 ;
        RECT 538.950 700.950 544.050 703.050 ;
        RECT 551.100 701.100 552.900 701.850 ;
        RECT 554.700 701.100 556.050 706.350 ;
        RECT 557.100 701.100 558.900 701.850 ;
        RECT 472.950 694.950 475.050 697.050 ;
        RECT 488.100 696.000 492.300 697.650 ;
        RECT 469.800 687.600 471.600 690.600 ;
        RECT 488.100 687.600 489.900 696.000 ;
        RECT 506.400 695.700 507.600 699.900 ;
        RECT 520.950 697.950 526.050 700.050 ;
        RECT 527.100 699.150 528.900 699.900 ;
        RECT 536.100 698.100 537.900 698.850 ;
        RECT 506.400 694.800 510.000 695.700 ;
        RECT 508.200 687.600 510.000 694.800 ;
        RECT 524.400 693.600 525.600 696.900 ;
        RECT 535.950 694.950 538.050 697.050 ;
        RECT 523.800 687.600 525.600 693.600 ;
        RECT 539.400 690.600 540.600 699.900 ;
        RECT 550.950 697.950 553.050 700.050 ;
        RECT 554.700 698.100 555.900 701.100 ;
        RECT 566.550 700.050 567.450 706.950 ;
        RECT 571.950 703.950 574.050 706.050 ;
        RECT 575.400 704.100 576.600 713.400 ;
        RECT 591.600 707.400 593.400 719.400 ;
        RECT 609.600 707.400 611.400 719.400 ;
        RECT 590.700 706.350 593.400 707.400 ;
        RECT 608.700 706.350 611.400 707.400 ;
        RECT 626.400 713.400 628.200 719.400 ;
        RECT 577.950 703.950 580.050 706.050 ;
        RECT 572.100 702.150 573.900 702.900 ;
        RECT 574.950 700.950 577.050 703.050 ;
        RECT 578.100 702.150 579.900 702.900 ;
        RECT 587.100 701.100 588.900 701.850 ;
        RECT 590.700 701.100 592.050 706.350 ;
        RECT 593.100 701.100 594.900 701.850 ;
        RECT 605.100 701.100 606.900 701.850 ;
        RECT 608.700 701.100 610.050 706.350 ;
        RECT 622.950 703.950 625.050 706.050 ;
        RECT 626.400 704.100 627.600 713.400 ;
        RECT 636.150 707.400 637.950 719.400 ;
        RECT 644.550 713.400 646.350 719.400 ;
        RECT 644.550 712.500 645.750 713.400 ;
        RECT 652.350 712.500 654.150 719.400 ;
        RECT 660.150 713.400 661.950 719.400 ;
        RECT 640.950 710.400 645.750 712.500 ;
        RECT 648.450 711.450 655.050 712.500 ;
        RECT 648.450 710.700 650.250 711.450 ;
        RECT 653.250 710.700 655.050 711.450 ;
        RECT 660.150 711.300 664.050 713.400 ;
        RECT 644.550 709.500 645.750 710.400 ;
        RECT 657.450 709.800 659.250 710.400 ;
        RECT 644.550 708.300 652.050 709.500 ;
        RECT 650.250 707.700 652.050 708.300 ;
        RECT 652.950 708.900 659.250 709.800 ;
        RECT 636.150 706.800 647.250 707.400 ;
        RECT 652.950 706.800 653.850 708.900 ;
        RECT 657.450 708.600 659.250 708.900 ;
        RECT 660.150 708.600 662.850 710.400 ;
        RECT 660.150 707.700 661.050 708.600 ;
        RECT 636.150 706.200 653.850 706.800 ;
        RECT 628.950 703.950 631.050 706.050 ;
        RECT 623.100 702.150 624.900 702.900 ;
        RECT 611.100 701.100 612.900 701.850 ;
        RECT 556.950 697.950 559.050 700.050 ;
        RECT 565.950 697.950 568.050 700.050 ;
        RECT 553.950 694.950 556.050 697.050 ;
        RECT 575.400 695.700 576.600 699.900 ;
        RECT 586.800 697.950 589.050 700.050 ;
        RECT 590.700 698.100 591.900 701.100 ;
        RECT 592.950 697.950 595.200 700.050 ;
        RECT 598.950 697.950 601.050 700.050 ;
        RECT 604.950 697.950 607.050 700.050 ;
        RECT 608.700 698.100 609.900 701.100 ;
        RECT 625.950 700.950 628.050 703.050 ;
        RECT 629.100 702.150 630.900 702.900 ;
        RECT 610.950 697.950 613.050 700.050 ;
        RECT 573.000 694.800 576.600 695.700 ;
        RECT 589.800 694.950 592.050 697.050 ;
        RECT 554.400 690.600 555.600 693.900 ;
        RECT 539.400 687.600 541.200 690.600 ;
        RECT 554.400 687.600 556.200 690.600 ;
        RECT 573.000 687.600 574.800 694.800 ;
        RECT 590.400 690.600 591.600 693.900 ;
        RECT 599.550 691.050 600.450 697.950 ;
        RECT 607.950 694.950 610.050 697.050 ;
        RECT 626.400 695.700 627.600 699.900 ;
        RECT 626.400 694.800 630.000 695.700 ;
        RECT 590.400 687.600 592.200 690.600 ;
        RECT 598.950 688.950 601.050 691.050 ;
        RECT 608.400 690.600 609.600 693.900 ;
        RECT 608.400 687.600 610.200 690.600 ;
        RECT 628.200 687.600 630.000 694.800 ;
        RECT 636.150 693.600 637.050 706.200 ;
        RECT 645.450 705.900 653.850 706.200 ;
        RECT 655.050 706.800 661.050 707.700 ;
        RECT 661.950 706.800 664.050 707.700 ;
        RECT 667.650 707.400 669.450 719.400 ;
        RECT 645.450 705.600 647.250 705.900 ;
        RECT 655.050 701.100 655.950 706.800 ;
        RECT 661.950 705.600 666.150 706.800 ;
        RECT 665.250 703.800 667.050 705.600 ;
        RECT 638.100 699.150 639.900 700.950 ;
        RECT 641.100 700.800 642.900 701.100 ;
        RECT 641.100 699.900 645.900 700.800 ;
        RECT 668.250 700.050 669.450 707.400 ;
        RECT 680.400 713.400 682.200 719.400 ;
        RECT 698.400 713.400 700.200 719.400 ;
        RECT 676.950 703.950 679.050 706.050 ;
        RECT 680.400 704.100 681.600 713.400 ;
        RECT 682.950 703.950 685.050 706.050 ;
        RECT 698.400 704.100 699.600 713.400 ;
        RECT 704.550 707.400 706.350 719.400 ;
        RECT 712.050 713.400 713.850 719.400 ;
        RECT 709.950 711.300 713.850 713.400 ;
        RECT 719.850 712.500 721.650 719.400 ;
        RECT 727.650 713.400 729.450 719.400 ;
        RECT 728.250 712.500 729.450 713.400 ;
        RECT 718.950 711.450 725.550 712.500 ;
        RECT 718.950 710.700 720.750 711.450 ;
        RECT 723.750 710.700 725.550 711.450 ;
        RECT 728.250 710.400 733.050 712.500 ;
        RECT 711.150 708.600 713.850 710.400 ;
        RECT 714.750 709.800 716.550 710.400 ;
        RECT 714.750 708.900 721.050 709.800 ;
        RECT 728.250 709.500 729.450 710.400 ;
        RECT 714.750 708.600 716.550 708.900 ;
        RECT 712.950 707.700 713.850 708.600 ;
        RECT 677.100 702.150 678.900 702.900 ;
        RECT 679.950 700.950 682.050 703.050 ;
        RECT 683.100 702.150 684.900 702.900 ;
        RECT 697.950 700.950 700.050 703.050 ;
        RECT 641.100 699.300 642.900 699.900 ;
        RECT 639.000 698.400 639.900 699.150 ;
        RECT 644.100 698.400 645.900 699.000 ;
        RECT 639.000 697.200 645.900 698.400 ;
        RECT 646.950 697.950 649.050 700.050 ;
        RECT 652.950 697.950 655.050 700.050 ;
        RECT 663.150 697.950 663.900 699.750 ;
        RECT 664.950 697.950 667.050 700.050 ;
        RECT 668.100 697.950 669.450 700.050 ;
        RECT 704.550 700.050 705.750 707.400 ;
        RECT 709.950 706.800 712.050 707.700 ;
        RECT 712.950 706.800 718.950 707.700 ;
        RECT 707.850 705.600 712.050 706.800 ;
        RECT 706.950 703.800 708.750 705.600 ;
        RECT 718.050 701.100 718.950 706.800 ;
        RECT 720.150 706.800 721.050 708.900 ;
        RECT 721.950 708.300 729.450 709.500 ;
        RECT 721.950 707.700 723.750 708.300 ;
        RECT 736.050 707.400 737.850 719.400 ;
        RECT 726.750 706.800 737.850 707.400 ;
        RECT 720.150 706.200 737.850 706.800 ;
        RECT 720.150 705.900 728.550 706.200 ;
        RECT 726.750 705.600 728.550 705.900 ;
        RECT 731.100 700.800 732.900 701.100 ;
        RECT 644.850 696.000 645.900 697.200 ;
        RECT 655.050 696.000 655.950 696.900 ;
        RECT 644.850 695.100 655.950 696.000 ;
        RECT 644.850 694.200 645.900 695.100 ;
        RECT 655.050 694.800 655.950 695.100 ;
        RECT 636.150 687.600 637.950 693.600 ;
        RECT 640.950 691.500 643.050 693.600 ;
        RECT 644.550 692.400 646.350 694.200 ;
        RECT 647.850 693.450 649.650 694.200 ;
        RECT 647.850 692.400 652.800 693.450 ;
        RECT 655.050 693.000 656.850 694.800 ;
        RECT 668.250 693.600 669.450 697.950 ;
        RECT 680.400 695.700 681.600 699.900 ;
        RECT 695.100 698.100 696.900 698.850 ;
        RECT 680.400 694.800 684.000 695.700 ;
        RECT 661.950 692.700 664.050 693.600 ;
        RECT 642.000 690.600 643.050 691.500 ;
        RECT 651.750 690.600 652.800 692.400 ;
        RECT 660.300 691.500 664.050 692.700 ;
        RECT 660.300 690.600 661.350 691.500 ;
        RECT 642.000 689.700 645.750 690.600 ;
        RECT 643.950 687.600 645.750 689.700 ;
        RECT 651.750 687.600 653.550 690.600 ;
        RECT 659.550 687.600 661.350 690.600 ;
        RECT 667.650 687.600 669.450 693.600 ;
        RECT 682.200 687.600 684.000 694.800 ;
        RECT 698.400 690.600 699.600 699.900 ;
        RECT 704.550 697.950 705.900 700.050 ;
        RECT 706.950 697.950 709.050 700.050 ;
        RECT 710.100 697.950 710.850 699.750 ;
        RECT 718.950 697.950 721.050 700.050 ;
        RECT 724.950 697.950 727.050 700.050 ;
        RECT 728.100 699.900 732.900 700.800 ;
        RECT 731.100 699.300 732.900 699.900 ;
        RECT 734.100 699.150 735.900 700.950 ;
        RECT 728.100 698.400 729.900 699.000 ;
        RECT 734.100 698.400 735.000 699.150 ;
        RECT 704.550 693.600 705.750 697.950 ;
        RECT 728.100 697.200 735.000 698.400 ;
        RECT 718.050 696.000 718.950 696.900 ;
        RECT 728.100 696.000 729.150 697.200 ;
        RECT 718.050 695.100 729.150 696.000 ;
        RECT 718.050 694.800 718.950 695.100 ;
        RECT 698.400 687.600 700.200 690.600 ;
        RECT 704.550 687.600 706.350 693.600 ;
        RECT 709.950 692.700 712.050 693.600 ;
        RECT 717.150 693.000 718.950 694.800 ;
        RECT 728.100 694.200 729.150 695.100 ;
        RECT 724.350 693.450 726.150 694.200 ;
        RECT 709.950 691.500 713.700 692.700 ;
        RECT 712.650 690.600 713.700 691.500 ;
        RECT 721.200 692.400 726.150 693.450 ;
        RECT 727.650 692.400 729.450 694.200 ;
        RECT 736.950 693.600 737.850 706.200 ;
        RECT 749.400 713.400 751.200 719.400 ;
        RECT 745.950 703.950 748.050 706.050 ;
        RECT 749.400 704.100 750.600 713.400 ;
        RECT 770.700 707.400 772.500 719.400 ;
        RECT 787.500 707.400 789.300 719.400 ;
        RECT 793.800 713.400 795.600 719.400 ;
        RECT 805.800 713.400 807.600 719.400 ;
        RECT 751.950 703.950 754.050 706.050 ;
        RECT 770.850 704.100 772.050 707.400 ;
        RECT 746.100 702.150 747.900 702.900 ;
        RECT 748.950 700.950 751.050 703.050 ;
        RECT 752.100 702.150 753.900 702.900 ;
        RECT 766.950 700.950 769.050 703.050 ;
        RECT 770.850 701.100 771.900 704.100 ;
        RECT 772.950 700.950 775.050 703.050 ;
        RECT 776.100 701.100 777.900 701.850 ;
        RECT 787.800 701.100 789.000 707.400 ;
        RECT 794.400 706.500 795.600 713.400 ;
        RECT 789.900 705.600 795.600 706.500 ;
        RECT 789.900 704.700 791.850 705.600 ;
        RECT 790.950 701.100 791.850 704.700 ;
        RECT 806.400 704.100 807.600 713.400 ;
        RECT 813.150 707.400 814.950 719.400 ;
        RECT 821.550 713.400 823.350 719.400 ;
        RECT 821.550 712.500 822.750 713.400 ;
        RECT 829.350 712.500 831.150 719.400 ;
        RECT 837.150 713.400 838.950 719.400 ;
        RECT 817.950 710.400 822.750 712.500 ;
        RECT 825.450 711.450 832.050 712.500 ;
        RECT 825.450 710.700 827.250 711.450 ;
        RECT 830.250 710.700 832.050 711.450 ;
        RECT 837.150 711.300 841.050 713.400 ;
        RECT 821.550 709.500 822.750 710.400 ;
        RECT 834.450 709.800 836.250 710.400 ;
        RECT 821.550 708.300 829.050 709.500 ;
        RECT 827.250 707.700 829.050 708.300 ;
        RECT 829.950 708.900 836.250 709.800 ;
        RECT 813.150 706.800 824.250 707.400 ;
        RECT 829.950 706.800 830.850 708.900 ;
        RECT 834.450 708.600 836.250 708.900 ;
        RECT 837.150 708.600 839.850 710.400 ;
        RECT 837.150 707.700 838.050 708.600 ;
        RECT 813.150 706.200 830.850 706.800 ;
        RECT 794.100 701.100 795.900 701.850 ;
        RECT 749.400 695.700 750.600 699.900 ;
        RECT 767.100 699.150 768.900 699.900 ;
        RECT 769.950 697.950 772.050 700.050 ;
        RECT 773.100 699.150 774.900 699.900 ;
        RECT 775.950 697.950 781.050 700.050 ;
        RECT 784.950 697.950 790.050 700.050 ;
        RECT 791.100 696.900 791.850 701.100 ;
        RECT 805.950 700.950 808.050 703.050 ;
        RECT 793.950 697.950 796.050 700.050 ;
        RECT 769.950 696.750 771.150 696.900 ;
        RECT 767.400 695.700 771.150 696.750 ;
        RECT 749.400 694.800 753.000 695.700 ;
        RECT 721.200 690.600 722.250 692.400 ;
        RECT 730.950 691.500 733.050 693.600 ;
        RECT 730.950 690.600 732.000 691.500 ;
        RECT 712.650 687.600 714.450 690.600 ;
        RECT 720.450 687.600 722.250 690.600 ;
        RECT 728.250 689.700 732.000 690.600 ;
        RECT 728.250 687.600 730.050 689.700 ;
        RECT 736.050 687.600 737.850 693.600 ;
        RECT 751.200 687.600 753.000 694.800 ;
        RECT 767.400 693.600 768.600 695.700 ;
        RECT 766.800 687.600 768.600 693.600 ;
        RECT 769.800 692.700 777.600 694.050 ;
        RECT 787.800 693.600 789.000 696.900 ;
        RECT 790.950 696.300 791.850 696.900 ;
        RECT 789.900 695.400 791.850 696.300 ;
        RECT 789.900 694.500 795.000 695.400 ;
        RECT 769.800 687.600 771.600 692.700 ;
        RECT 775.800 687.600 777.600 692.700 ;
        RECT 787.500 687.600 789.300 693.600 ;
        RECT 793.800 690.600 795.000 694.500 ;
        RECT 806.400 690.600 807.600 699.900 ;
        RECT 809.100 698.100 810.900 698.850 ;
        RECT 793.800 687.600 795.600 690.600 ;
        RECT 805.800 687.600 807.600 690.600 ;
        RECT 813.150 693.600 814.050 706.200 ;
        RECT 822.450 705.900 830.850 706.200 ;
        RECT 832.050 706.800 838.050 707.700 ;
        RECT 838.950 706.800 841.050 707.700 ;
        RECT 844.650 707.400 846.450 719.400 ;
        RECT 822.450 705.600 824.250 705.900 ;
        RECT 832.050 701.100 832.950 706.800 ;
        RECT 838.950 705.600 843.150 706.800 ;
        RECT 842.250 703.800 844.050 705.600 ;
        RECT 815.100 699.150 816.900 700.950 ;
        RECT 818.100 700.800 819.900 701.100 ;
        RECT 818.100 699.900 822.900 700.800 ;
        RECT 845.250 700.050 846.450 707.400 ;
        RECT 818.100 699.300 819.900 699.900 ;
        RECT 816.000 698.400 816.900 699.150 ;
        RECT 821.100 698.400 822.900 699.000 ;
        RECT 816.000 697.200 822.900 698.400 ;
        RECT 823.800 697.950 826.050 700.050 ;
        RECT 829.950 697.950 832.050 700.050 ;
        RECT 840.150 697.950 840.900 699.750 ;
        RECT 841.950 697.950 844.050 700.050 ;
        RECT 845.100 697.950 846.450 700.050 ;
        RECT 821.850 696.000 822.900 697.200 ;
        RECT 832.050 696.000 832.950 696.900 ;
        RECT 821.850 695.100 832.950 696.000 ;
        RECT 821.850 694.200 822.900 695.100 ;
        RECT 832.050 694.800 832.950 695.100 ;
        RECT 813.150 687.600 814.950 693.600 ;
        RECT 817.950 691.500 820.050 693.600 ;
        RECT 821.550 692.400 823.350 694.200 ;
        RECT 824.850 693.450 826.650 694.200 ;
        RECT 824.850 692.400 829.800 693.450 ;
        RECT 832.050 693.000 833.850 694.800 ;
        RECT 845.250 693.600 846.450 697.950 ;
        RECT 838.950 692.700 841.050 693.600 ;
        RECT 819.000 690.600 820.050 691.500 ;
        RECT 828.750 690.600 829.800 692.400 ;
        RECT 837.300 691.500 841.050 692.700 ;
        RECT 837.300 690.600 838.350 691.500 ;
        RECT 819.000 689.700 822.750 690.600 ;
        RECT 820.950 687.600 822.750 689.700 ;
        RECT 828.750 687.600 830.550 690.600 ;
        RECT 836.550 687.600 838.350 690.600 ;
        RECT 844.650 687.600 846.450 693.600 ;
        RECT 10.800 677.400 12.600 683.400 ;
        RECT 11.400 675.300 12.600 677.400 ;
        RECT 13.800 678.300 15.600 683.400 ;
        RECT 19.800 678.300 21.600 683.400 ;
        RECT 25.950 679.950 28.050 682.050 ;
        RECT 13.800 676.950 21.600 678.300 ;
        RECT 11.400 674.250 15.150 675.300 ;
        RECT 13.950 674.100 15.150 674.250 ;
        RECT 11.100 671.100 12.900 671.850 ;
        RECT 13.950 670.950 16.050 673.050 ;
        RECT 17.100 671.100 18.900 671.850 ;
        RECT 19.950 670.950 22.050 673.050 ;
        RECT 26.550 672.450 27.450 679.950 ;
        RECT 36.000 679.050 37.800 683.400 ;
        RECT 55.800 680.400 57.600 683.400 ;
        RECT 32.400 677.400 37.800 679.050 ;
        RECT 32.400 674.100 33.300 677.400 ;
        RECT 56.400 677.100 57.600 680.400 ;
        RECT 72.000 676.200 73.800 683.400 ;
        RECT 55.950 673.950 58.050 676.050 ;
        RECT 72.000 675.300 75.600 676.200 ;
        RECT 31.950 672.450 34.050 673.050 ;
        RECT 26.550 671.550 34.050 672.450 ;
        RECT 31.950 670.950 34.050 671.550 ;
        RECT 35.100 671.100 36.900 671.850 ;
        RECT 37.950 670.950 40.050 673.050 ;
        RECT 41.100 671.100 42.900 671.850 ;
        RECT 52.950 670.950 55.050 673.050 ;
        RECT 10.950 667.950 13.050 670.050 ;
        RECT 14.850 666.900 15.900 669.900 ;
        RECT 16.950 667.950 19.050 670.050 ;
        RECT 20.100 669.150 21.900 669.900 ;
        RECT 14.850 663.600 16.050 666.900 ;
        RECT 32.400 663.600 33.300 669.900 ;
        RECT 34.950 667.950 37.200 670.050 ;
        RECT 38.100 669.150 39.900 669.900 ;
        RECT 40.950 667.950 43.050 670.050 ;
        RECT 56.100 669.900 57.300 672.900 ;
        RECT 58.950 670.950 61.050 673.050 ;
        RECT 74.400 671.100 75.600 675.300 ;
        RECT 92.100 675.000 93.900 683.400 ;
        RECT 89.700 673.350 93.900 675.000 ;
        RECT 113.100 675.000 114.900 683.400 ;
        RECT 131.400 680.400 133.200 683.400 ;
        RECT 113.100 673.350 117.300 675.000 ;
        RECT 127.950 673.950 130.050 676.050 ;
        RECT 53.100 669.150 54.900 669.900 ;
        RECT 55.950 664.650 57.300 669.900 ;
        RECT 59.100 669.150 60.900 669.900 ;
        RECT 71.100 668.100 72.900 668.850 ;
        RECT 73.950 667.950 76.050 670.050 ;
        RECT 77.100 668.100 78.900 668.850 ;
        RECT 89.700 668.100 90.600 673.350 ;
        RECT 92.100 671.100 93.900 671.850 ;
        RECT 98.100 671.100 99.900 671.850 ;
        RECT 107.100 671.100 108.900 671.850 ;
        RECT 113.100 671.100 114.900 671.850 ;
        RECT 91.950 667.950 94.050 670.050 ;
        RECT 97.950 667.950 100.050 670.050 ;
        RECT 106.950 667.950 109.050 670.050 ;
        RECT 112.950 667.950 115.050 670.050 ;
        RECT 116.400 668.100 117.300 673.350 ;
        RECT 128.100 672.150 129.900 672.900 ;
        RECT 131.400 671.100 132.600 680.400 ;
        RECT 149.100 675.000 150.900 683.400 ;
        RECT 170.100 675.000 171.900 683.400 ;
        RECT 191.100 675.000 192.900 683.400 ;
        RECT 211.200 676.200 213.000 683.400 ;
        RECT 209.400 675.300 213.000 676.200 ;
        RECT 227.400 680.400 229.200 683.400 ;
        RECT 149.100 673.350 153.300 675.000 ;
        RECT 170.100 673.350 174.300 675.000 ;
        RECT 191.100 673.350 195.300 675.000 ;
        RECT 143.100 671.100 144.900 671.850 ;
        RECT 149.100 671.100 150.900 671.850 ;
        RECT 130.950 667.950 136.050 670.050 ;
        RECT 142.950 667.950 145.050 670.050 ;
        RECT 148.950 667.950 151.050 670.050 ;
        RECT 152.400 668.100 153.300 673.350 ;
        RECT 164.100 671.100 165.900 671.850 ;
        RECT 170.100 671.100 171.900 671.850 ;
        RECT 163.950 667.950 166.050 670.050 ;
        RECT 169.950 667.950 172.050 670.050 ;
        RECT 173.400 668.100 174.300 673.350 ;
        RECT 185.100 671.100 186.900 671.850 ;
        RECT 191.100 671.100 192.900 671.850 ;
        RECT 184.950 667.950 187.050 670.050 ;
        RECT 190.950 667.950 193.050 670.050 ;
        RECT 194.400 668.100 195.300 673.350 ;
        RECT 199.950 670.950 202.050 673.050 ;
        RECT 209.400 671.100 210.600 675.300 ;
        RECT 223.950 673.950 226.050 676.050 ;
        RECT 217.950 670.950 220.050 673.050 ;
        RECT 224.100 672.150 225.900 672.900 ;
        RECT 227.400 671.100 228.600 680.400 ;
        RECT 243.000 676.200 244.800 683.400 ;
        RECT 260.400 677.400 262.200 683.400 ;
        RECT 279.000 679.050 280.800 683.400 ;
        RECT 275.400 677.400 280.800 679.050 ;
        RECT 243.000 675.300 246.600 676.200 ;
        RECT 245.400 671.100 246.600 675.300 ;
        RECT 260.400 674.100 261.600 677.400 ;
        RECT 275.400 674.100 276.300 677.400 ;
        RECT 299.100 675.000 300.900 683.400 ;
        RECT 319.200 676.200 321.000 683.400 ;
        RECT 322.950 679.950 325.050 682.050 ;
        RECT 296.700 673.350 300.900 675.000 ;
        RECT 317.400 675.300 321.000 676.200 ;
        RECT 257.100 671.100 258.900 671.850 ;
        RECT 259.950 670.950 262.050 673.050 ;
        RECT 271.950 670.950 277.050 673.050 ;
        RECT 278.100 671.100 279.900 671.850 ;
        RECT 280.950 670.950 283.200 673.050 ;
        RECT 284.100 671.100 285.900 671.850 ;
        RECT 70.950 664.950 73.050 667.050 ;
        RECT 54.600 663.600 57.300 664.650 ;
        RECT 14.700 651.600 16.500 663.600 ;
        RECT 31.800 651.600 33.600 663.600 ;
        RECT 34.800 662.700 42.600 663.600 ;
        RECT 34.800 651.600 36.600 662.700 ;
        RECT 40.800 651.600 42.600 662.700 ;
        RECT 54.600 651.600 56.400 663.600 ;
        RECT 74.400 657.600 75.600 666.900 ;
        RECT 76.950 664.950 79.050 667.050 ;
        RECT 88.950 666.450 91.050 667.050 ;
        RECT 83.550 665.550 91.050 666.450 ;
        RECT 73.800 651.600 75.600 657.600 ;
        RECT 83.550 655.050 84.450 665.550 ;
        RECT 88.950 664.950 91.050 665.550 ;
        RECT 94.950 664.950 97.050 667.050 ;
        RECT 109.950 664.950 112.050 667.050 ;
        RECT 115.950 666.450 118.050 667.050 ;
        RECT 115.950 665.550 123.450 666.450 ;
        RECT 115.950 664.950 118.050 665.550 ;
        RECT 89.700 658.800 90.600 663.900 ;
        RECT 95.100 663.150 96.900 663.900 ;
        RECT 110.100 663.150 111.900 663.900 ;
        RECT 116.400 658.800 117.300 663.900 ;
        RECT 122.550 661.050 123.450 665.550 ;
        RECT 121.950 658.950 124.050 661.050 ;
        RECT 89.700 657.900 96.300 658.800 ;
        RECT 89.700 657.600 90.600 657.900 ;
        RECT 82.950 652.950 85.050 655.050 ;
        RECT 88.800 651.600 90.600 657.600 ;
        RECT 94.800 657.600 96.300 657.900 ;
        RECT 110.700 657.900 117.300 658.800 ;
        RECT 110.700 657.600 112.200 657.900 ;
        RECT 94.800 651.600 96.600 657.600 ;
        RECT 110.400 651.600 112.200 657.600 ;
        RECT 116.400 657.600 117.300 657.900 ;
        RECT 131.400 657.600 132.600 666.900 ;
        RECT 145.950 664.950 148.050 667.050 ;
        RECT 151.950 666.450 154.050 667.050 ;
        RECT 151.950 665.550 159.450 666.450 ;
        RECT 151.950 664.950 154.050 665.550 ;
        RECT 146.100 663.150 147.900 663.900 ;
        RECT 152.400 658.800 153.300 663.900 ;
        RECT 146.700 657.900 153.300 658.800 ;
        RECT 146.700 657.600 148.200 657.900 ;
        RECT 116.400 651.600 118.200 657.600 ;
        RECT 131.400 651.600 133.200 657.600 ;
        RECT 146.400 651.600 148.200 657.600 ;
        RECT 152.400 657.600 153.300 657.900 ;
        RECT 152.400 651.600 154.200 657.600 ;
        RECT 158.550 655.050 159.450 665.550 ;
        RECT 166.950 664.950 169.050 667.050 ;
        RECT 172.950 664.950 178.050 667.050 ;
        RECT 187.950 664.950 190.050 667.050 ;
        RECT 193.950 666.450 196.050 667.050 ;
        RECT 200.550 666.450 201.450 670.950 ;
        RECT 206.100 668.100 207.900 668.850 ;
        RECT 208.950 667.950 211.050 670.050 ;
        RECT 212.100 668.100 213.900 668.850 ;
        RECT 193.950 665.550 201.450 666.450 ;
        RECT 193.950 664.950 196.050 665.550 ;
        RECT 205.950 664.950 208.050 667.050 ;
        RECT 167.100 663.150 168.900 663.900 ;
        RECT 173.400 658.800 174.300 663.900 ;
        RECT 188.100 663.150 189.900 663.900 ;
        RECT 194.400 658.800 195.300 663.900 ;
        RECT 167.700 657.900 174.300 658.800 ;
        RECT 167.700 657.600 169.200 657.900 ;
        RECT 157.950 652.950 160.050 655.050 ;
        RECT 167.400 651.600 169.200 657.600 ;
        RECT 173.400 657.600 174.300 657.900 ;
        RECT 188.700 657.900 195.300 658.800 ;
        RECT 188.700 657.600 190.200 657.900 ;
        RECT 173.400 651.600 175.200 657.600 ;
        RECT 188.400 651.600 190.200 657.600 ;
        RECT 194.400 657.600 195.300 657.900 ;
        RECT 209.400 657.600 210.600 666.900 ;
        RECT 211.950 664.950 214.200 667.050 ;
        RECT 218.550 664.050 219.450 670.950 ;
        RECT 224.100 667.950 229.050 670.050 ;
        RECT 242.100 668.100 243.900 668.850 ;
        RECT 244.800 667.950 247.050 670.050 ;
        RECT 248.100 668.100 249.900 668.850 ;
        RECT 256.950 667.950 259.050 670.050 ;
        RECT 217.950 661.950 220.050 664.050 ;
        RECT 227.400 657.600 228.600 666.900 ;
        RECT 241.950 664.950 244.050 667.050 ;
        RECT 245.400 657.600 246.600 666.900 ;
        RECT 247.950 664.950 250.050 667.050 ;
        RECT 194.400 651.600 196.200 657.600 ;
        RECT 209.400 651.600 211.200 657.600 ;
        RECT 227.400 651.600 229.200 657.600 ;
        RECT 244.800 651.600 246.600 657.600 ;
        RECT 260.400 663.600 261.600 669.900 ;
        RECT 275.400 663.600 276.300 669.900 ;
        RECT 277.950 667.950 280.050 670.050 ;
        RECT 281.100 669.150 282.900 669.900 ;
        RECT 283.950 667.950 286.050 670.050 ;
        RECT 296.700 668.100 297.600 673.350 ;
        RECT 299.100 671.100 300.900 671.850 ;
        RECT 305.100 671.100 306.900 671.850 ;
        RECT 317.400 671.100 318.600 675.300 ;
        RECT 323.550 673.050 324.450 679.950 ;
        RECT 334.800 677.400 336.600 683.400 ;
        RECT 335.400 675.300 336.600 677.400 ;
        RECT 337.800 678.300 339.600 683.400 ;
        RECT 343.800 678.300 345.600 683.400 ;
        RECT 349.950 679.950 352.050 682.050 ;
        RECT 337.800 676.950 345.600 678.300 ;
        RECT 335.400 674.250 339.150 675.300 ;
        RECT 337.950 674.100 339.150 674.250 ;
        RECT 322.950 670.950 325.050 673.050 ;
        RECT 335.100 671.100 336.900 671.850 ;
        RECT 337.950 670.950 340.050 673.050 ;
        RECT 341.100 671.100 342.900 671.850 ;
        RECT 343.950 670.950 346.050 673.050 ;
        RECT 298.950 667.950 301.050 670.050 ;
        RECT 304.950 667.950 307.050 670.050 ;
        RECT 314.100 668.100 315.900 668.850 ;
        RECT 316.950 667.950 319.050 670.050 ;
        RECT 320.100 668.100 321.900 668.850 ;
        RECT 334.800 667.950 337.050 670.050 ;
        RECT 289.950 666.450 294.000 667.050 ;
        RECT 295.950 666.450 298.050 667.050 ;
        RECT 289.950 665.550 298.050 666.450 ;
        RECT 289.950 664.950 294.000 665.550 ;
        RECT 295.950 664.950 298.050 665.550 ;
        RECT 301.950 664.950 304.200 667.050 ;
        RECT 313.950 664.950 316.050 667.050 ;
        RECT 260.400 651.600 262.200 663.600 ;
        RECT 274.800 651.600 276.600 663.600 ;
        RECT 277.800 662.700 285.600 663.600 ;
        RECT 277.800 651.600 279.600 662.700 ;
        RECT 283.800 651.600 285.600 662.700 ;
        RECT 296.700 658.800 297.600 663.900 ;
        RECT 302.100 663.150 303.900 663.900 ;
        RECT 296.700 657.900 303.300 658.800 ;
        RECT 296.700 657.600 297.600 657.900 ;
        RECT 295.800 651.600 297.600 657.600 ;
        RECT 301.800 657.600 303.300 657.900 ;
        RECT 317.400 657.600 318.600 666.900 ;
        RECT 319.950 664.950 322.050 667.050 ;
        RECT 338.850 666.900 339.900 669.900 ;
        RECT 340.950 667.950 343.050 670.050 ;
        RECT 344.100 669.150 345.900 669.900 ;
        RECT 338.850 663.600 340.050 666.900 ;
        RECT 301.800 651.600 303.600 657.600 ;
        RECT 317.400 651.600 319.200 657.600 ;
        RECT 338.700 651.600 340.500 663.600 ;
        RECT 350.550 658.050 351.450 679.950 ;
        RECT 357.000 676.200 358.800 683.400 ;
        RECT 375.300 679.200 377.100 683.400 ;
        RECT 375.150 677.400 377.100 679.200 ;
        RECT 357.000 675.300 360.600 676.200 ;
        RECT 359.400 671.100 360.600 675.300 ;
        RECT 375.150 674.100 376.050 677.400 ;
        RECT 377.100 675.900 378.900 676.500 ;
        RECT 382.800 675.900 384.600 683.400 ;
        RECT 377.100 674.700 384.600 675.900 ;
        RECT 402.000 677.400 403.800 683.400 ;
        RECT 373.950 672.450 376.050 673.050 ;
        RECT 368.550 671.550 376.050 672.450 ;
        RECT 356.100 668.100 357.900 668.850 ;
        RECT 358.950 667.950 361.050 670.050 ;
        RECT 362.100 668.100 363.900 668.850 ;
        RECT 368.550 667.050 369.450 671.550 ;
        RECT 373.950 670.950 376.050 671.550 ;
        RECT 377.100 671.100 378.900 671.850 ;
        RECT 355.950 664.950 358.050 667.050 ;
        RECT 349.950 655.950 352.050 658.050 ;
        RECT 359.400 657.600 360.600 666.900 ;
        RECT 361.950 664.950 364.050 667.050 ;
        RECT 367.950 664.950 370.050 667.050 ;
        RECT 362.550 663.000 363.450 664.950 ;
        RECT 373.950 663.600 375.000 669.900 ;
        RECT 376.950 667.950 379.050 670.050 ;
        RECT 361.950 658.950 364.050 663.000 ;
        RECT 358.800 651.600 360.600 657.600 ;
        RECT 373.200 651.600 375.000 663.600 ;
        RECT 380.550 657.600 381.600 674.700 ;
        RECT 402.000 674.100 403.050 677.400 ;
        RECT 421.200 676.200 423.000 683.400 ;
        RECT 440.400 680.400 442.200 683.400 ;
        RECT 455.400 680.400 457.200 683.400 ;
        RECT 440.400 677.100 441.600 680.400 ;
        RECT 419.400 675.300 423.000 676.200 ;
        RECT 456.000 676.500 457.200 680.400 ;
        RECT 461.700 677.400 463.500 683.400 ;
        RECT 382.950 670.950 385.050 673.050 ;
        RECT 394.950 670.950 397.050 673.050 ;
        RECT 398.250 671.100 399.900 671.850 ;
        RECT 400.950 670.950 403.050 673.050 ;
        RECT 404.100 671.100 405.750 671.850 ;
        RECT 406.950 670.950 409.200 673.050 ;
        RECT 419.400 671.100 420.600 675.300 ;
        RECT 439.950 673.950 442.200 676.050 ;
        RECT 456.000 675.600 461.100 676.500 ;
        RECT 459.150 674.700 461.100 675.600 ;
        RECT 459.150 674.100 460.050 674.700 ;
        RECT 462.000 674.100 463.200 677.400 ;
        RECT 478.200 676.200 480.000 683.400 ;
        RECT 476.400 675.300 480.000 676.200 ;
        RECT 494.400 677.400 496.200 683.400 ;
        RECT 506.400 678.300 508.200 683.400 ;
        RECT 512.400 678.300 514.200 683.400 ;
        RECT 436.950 670.950 439.050 673.050 ;
        RECT 383.100 669.150 384.900 669.900 ;
        RECT 395.100 669.150 396.900 669.900 ;
        RECT 397.950 667.950 400.200 670.050 ;
        RECT 401.100 666.900 401.850 669.900 ;
        RECT 403.950 667.950 406.050 670.050 ;
        RECT 407.100 669.150 408.750 669.900 ;
        RECT 416.100 668.100 417.900 668.850 ;
        RECT 418.950 667.950 421.050 670.050 ;
        RECT 440.700 669.900 441.900 672.900 ;
        RECT 442.950 670.950 445.050 673.050 ;
        RECT 454.950 670.950 457.050 673.050 ;
        RECT 459.150 669.900 459.900 674.100 ;
        RECT 460.950 670.950 466.050 673.050 ;
        RECT 476.400 671.100 477.600 675.300 ;
        RECT 494.400 674.100 495.600 677.400 ;
        RECT 506.400 676.950 514.200 678.300 ;
        RECT 515.400 677.400 517.200 683.400 ;
        RECT 530.400 680.400 532.200 683.400 ;
        RECT 515.400 675.300 516.600 677.400 ;
        RECT 531.300 676.200 532.200 680.400 ;
        RECT 536.400 677.400 538.200 683.400 ;
        RECT 548.400 678.300 550.200 683.400 ;
        RECT 554.400 678.300 556.200 683.400 ;
        RECT 512.850 674.250 516.600 675.300 ;
        RECT 512.850 674.100 514.050 674.250 ;
        RECT 526.950 673.950 529.050 676.050 ;
        RECT 531.300 675.300 534.750 676.200 ;
        RECT 532.950 674.400 534.750 675.300 ;
        RECT 485.100 670.950 487.200 673.050 ;
        RECT 491.100 671.100 492.900 671.850 ;
        RECT 493.950 670.950 499.050 673.050 ;
        RECT 505.950 670.950 508.050 673.050 ;
        RECT 509.100 671.100 510.900 671.850 ;
        RECT 511.950 670.950 514.050 673.050 ;
        RECT 527.100 672.150 528.900 672.900 ;
        RECT 515.100 671.100 516.900 671.850 ;
        RECT 529.950 670.950 532.050 673.050 ;
        RECT 437.100 669.150 438.900 669.900 ;
        RECT 422.100 668.100 423.900 668.850 ;
        RECT 400.950 665.400 401.850 666.900 ;
        RECT 397.800 664.500 401.850 665.400 ;
        RECT 415.950 664.950 418.050 667.050 ;
        RECT 379.800 651.600 381.600 657.600 ;
        RECT 394.800 652.500 396.600 663.600 ;
        RECT 397.800 653.400 399.600 664.500 ;
        RECT 400.800 662.400 408.600 663.300 ;
        RECT 400.800 652.500 402.600 662.400 ;
        RECT 394.800 651.600 402.600 652.500 ;
        RECT 406.800 651.600 408.600 662.400 ;
        RECT 419.400 657.600 420.600 666.900 ;
        RECT 421.950 664.950 424.050 667.050 ;
        RECT 440.700 664.650 442.050 669.900 ;
        RECT 443.100 669.150 444.900 669.900 ;
        RECT 455.100 669.150 456.900 669.900 ;
        RECT 459.150 666.300 460.050 669.900 ;
        RECT 459.150 665.400 461.100 666.300 ;
        RECT 440.700 663.600 443.400 664.650 ;
        RECT 419.400 651.600 421.200 657.600 ;
        RECT 441.600 651.600 443.400 663.600 ;
        RECT 455.400 664.500 461.100 665.400 ;
        RECT 455.400 657.600 456.600 664.500 ;
        RECT 462.000 663.600 463.200 669.900 ;
        RECT 473.100 668.100 474.900 668.850 ;
        RECT 475.950 667.950 478.200 670.050 ;
        RECT 479.100 668.100 480.900 668.850 ;
        RECT 485.550 667.050 486.450 670.950 ;
        RECT 490.950 667.950 493.050 670.050 ;
        RECT 472.950 664.950 475.050 667.050 ;
        RECT 455.400 651.600 457.200 657.600 ;
        RECT 461.700 651.600 463.500 663.600 ;
        RECT 473.550 663.000 474.450 664.950 ;
        RECT 472.950 658.950 475.050 663.000 ;
        RECT 476.400 657.600 477.600 666.900 ;
        RECT 478.950 664.950 481.050 667.050 ;
        RECT 484.950 664.950 487.050 667.050 ;
        RECT 494.400 663.600 495.600 669.900 ;
        RECT 506.100 669.150 507.900 669.900 ;
        RECT 508.950 667.950 511.050 670.050 ;
        RECT 512.100 666.900 513.150 669.900 ;
        RECT 514.950 667.950 517.050 670.050 ;
        RECT 530.100 669.150 531.900 669.900 ;
        RECT 511.950 663.600 513.150 666.900 ;
        RECT 533.700 666.600 534.600 674.400 ;
        RECT 537.000 671.100 538.050 677.400 ;
        RECT 548.400 676.950 556.200 678.300 ;
        RECT 557.400 677.400 559.200 683.400 ;
        RECT 557.400 675.300 558.600 677.400 ;
        RECT 573.000 676.200 574.800 683.400 ;
        RECT 589.500 677.400 591.300 683.400 ;
        RECT 595.800 680.400 597.600 683.400 ;
        RECT 605.400 680.400 607.200 683.400 ;
        RECT 573.000 675.300 576.600 676.200 ;
        RECT 554.850 674.250 558.600 675.300 ;
        RECT 554.850 674.100 556.050 674.250 ;
        RECT 547.950 670.950 550.050 673.050 ;
        RECT 551.100 671.100 552.900 671.850 ;
        RECT 553.950 670.950 556.200 673.050 ;
        RECT 557.100 671.100 558.900 671.850 ;
        RECT 575.400 671.100 576.600 675.300 ;
        RECT 589.800 674.100 591.000 677.400 ;
        RECT 595.800 676.500 597.000 680.400 ;
        RECT 591.900 675.600 597.000 676.500 ;
        RECT 606.000 676.500 607.200 680.400 ;
        RECT 611.700 677.400 613.500 683.400 ;
        RECT 606.000 675.600 611.100 676.500 ;
        RECT 591.900 674.700 593.850 675.600 ;
        RECT 592.950 674.100 593.850 674.700 ;
        RECT 589.950 670.950 592.050 673.050 ;
        RECT 535.950 667.950 538.050 670.050 ;
        RECT 548.100 669.150 549.900 669.900 ;
        RECT 550.950 667.950 553.050 670.050 ;
        RECT 554.100 666.900 555.150 669.900 ;
        RECT 556.950 667.950 559.050 670.050 ;
        RECT 572.100 668.100 573.900 668.850 ;
        RECT 574.950 667.950 577.050 670.050 ;
        RECT 593.100 669.900 593.850 674.100 ;
        RECT 609.150 674.700 611.100 675.600 ;
        RECT 609.150 674.100 610.050 674.700 ;
        RECT 612.000 674.100 613.200 677.400 ;
        RECT 627.000 676.200 628.800 683.400 ;
        RECT 643.800 677.400 645.600 683.400 ;
        RECT 627.000 675.300 630.600 676.200 ;
        RECT 595.950 670.950 598.200 673.050 ;
        RECT 604.950 670.950 607.050 673.050 ;
        RECT 609.150 669.900 609.900 674.100 ;
        RECT 610.950 672.450 613.050 673.050 ;
        RECT 616.950 672.450 619.050 673.050 ;
        RECT 610.950 671.550 619.050 672.450 ;
        RECT 610.950 670.950 613.050 671.550 ;
        RECT 616.950 670.950 619.050 671.550 ;
        RECT 629.400 671.100 630.600 675.300 ;
        RECT 644.400 675.300 645.600 677.400 ;
        RECT 646.800 678.300 648.600 683.400 ;
        RECT 652.800 678.300 654.600 683.400 ;
        RECT 646.800 676.950 654.600 678.300 ;
        RECT 665.400 676.500 667.200 683.400 ;
        RECT 671.400 676.500 673.200 683.400 ;
        RECT 677.400 676.500 679.200 683.400 ;
        RECT 683.400 676.500 685.200 683.400 ;
        RECT 692.550 677.400 694.350 683.400 ;
        RECT 700.650 680.400 702.450 683.400 ;
        RECT 708.450 680.400 710.250 683.400 ;
        RECT 716.250 681.300 718.050 683.400 ;
        RECT 716.250 680.400 720.000 681.300 ;
        RECT 700.650 679.500 701.700 680.400 ;
        RECT 697.950 678.300 701.700 679.500 ;
        RECT 709.200 678.600 710.250 680.400 ;
        RECT 718.950 679.500 720.000 680.400 ;
        RECT 697.950 677.400 700.050 678.300 ;
        RECT 665.400 675.300 669.300 676.500 ;
        RECT 671.400 675.300 675.300 676.500 ;
        RECT 677.400 675.300 681.300 676.500 ;
        RECT 683.400 675.300 686.100 676.500 ;
        RECT 644.400 674.250 648.150 675.300 ;
        RECT 646.950 674.100 648.150 674.250 ;
        RECT 668.100 674.400 669.300 675.300 ;
        RECT 674.100 674.400 675.300 675.300 ;
        RECT 680.100 674.400 681.300 675.300 ;
        RECT 668.100 673.200 672.300 674.400 ;
        RECT 644.100 671.100 645.900 671.850 ;
        RECT 646.950 670.950 649.200 673.050 ;
        RECT 650.100 671.100 651.900 671.850 ;
        RECT 652.950 670.950 655.050 673.050 ;
        RECT 665.100 671.100 666.900 671.850 ;
        RECT 578.100 668.100 579.900 668.850 ;
        RECT 532.800 666.000 534.600 666.600 ;
        RECT 527.400 664.800 534.600 666.000 ;
        RECT 527.400 663.600 528.600 664.800 ;
        RECT 533.700 664.650 534.600 664.800 ;
        RECT 535.950 663.600 537.300 666.900 ;
        RECT 553.950 663.600 555.150 666.900 ;
        RECT 571.950 664.950 574.050 667.050 ;
        RECT 476.400 651.600 478.200 657.600 ;
        RECT 494.400 651.600 496.200 663.600 ;
        RECT 511.500 651.600 513.300 663.600 ;
        RECT 527.400 651.600 529.200 663.600 ;
        RECT 534.900 662.100 537.300 663.600 ;
        RECT 534.900 651.600 536.700 662.100 ;
        RECT 553.500 651.600 555.300 663.600 ;
        RECT 575.400 657.600 576.600 666.900 ;
        RECT 577.950 664.950 580.200 667.050 ;
        RECT 589.800 663.600 591.000 669.900 ;
        RECT 592.950 666.300 593.850 669.900 ;
        RECT 596.100 669.150 597.900 669.900 ;
        RECT 605.100 669.150 606.900 669.900 ;
        RECT 591.900 665.400 593.850 666.300 ;
        RECT 609.150 666.300 610.050 669.900 ;
        RECT 609.150 665.400 611.100 666.300 ;
        RECT 591.900 664.500 597.600 665.400 ;
        RECT 574.800 651.600 576.600 657.600 ;
        RECT 589.500 651.600 591.300 663.600 ;
        RECT 596.400 657.600 597.600 664.500 ;
        RECT 595.800 651.600 597.600 657.600 ;
        RECT 605.400 664.500 611.100 665.400 ;
        RECT 605.400 657.600 606.600 664.500 ;
        RECT 612.000 663.600 613.200 669.900 ;
        RECT 617.550 667.050 618.450 670.950 ;
        RECT 626.100 668.100 627.900 668.850 ;
        RECT 628.950 667.950 631.050 670.050 ;
        RECT 632.100 668.100 633.900 668.850 ;
        RECT 643.800 667.950 646.050 670.050 ;
        RECT 616.950 664.950 619.050 667.050 ;
        RECT 625.950 664.950 628.050 667.050 ;
        RECT 605.400 651.600 607.200 657.600 ;
        RECT 611.700 651.600 613.500 663.600 ;
        RECT 629.400 657.600 630.600 666.900 ;
        RECT 631.950 664.950 634.050 667.050 ;
        RECT 647.850 666.900 648.900 669.900 ;
        RECT 649.950 667.950 652.050 670.050 ;
        RECT 653.100 669.150 654.900 669.900 ;
        RECT 647.850 663.600 649.050 666.900 ;
        RECT 668.100 665.700 669.300 673.200 ;
        RECT 670.500 672.600 672.300 673.200 ;
        RECT 674.100 673.200 678.300 674.400 ;
        RECT 674.100 665.700 675.300 673.200 ;
        RECT 676.500 672.600 678.300 673.200 ;
        RECT 680.100 673.200 684.300 674.400 ;
        RECT 680.100 665.700 681.300 673.200 ;
        RECT 682.500 672.600 684.300 673.200 ;
        RECT 685.200 671.100 686.100 675.300 ;
        RECT 692.550 673.050 693.750 677.400 ;
        RECT 705.150 676.200 706.950 678.000 ;
        RECT 709.200 677.550 714.150 678.600 ;
        RECT 712.350 676.800 714.150 677.550 ;
        RECT 715.650 676.800 717.450 678.600 ;
        RECT 718.950 677.400 721.050 679.500 ;
        RECT 724.050 677.400 725.850 683.400 ;
        RECT 736.800 677.400 738.600 683.400 ;
        RECT 706.050 675.900 706.950 676.200 ;
        RECT 716.100 675.900 717.150 676.800 ;
        RECT 706.050 675.000 717.150 675.900 ;
        RECT 706.050 674.100 706.950 675.000 ;
        RECT 716.100 673.800 717.150 675.000 ;
        RECT 692.550 670.950 693.900 673.050 ;
        RECT 694.950 670.950 697.200 673.050 ;
        RECT 698.100 671.250 698.850 673.050 ;
        RECT 706.800 670.950 709.050 673.050 ;
        RECT 712.950 670.950 715.050 673.050 ;
        RECT 716.100 672.600 723.000 673.800 ;
        RECT 716.100 672.000 717.900 672.600 ;
        RECT 722.100 671.850 723.000 672.600 ;
        RECT 719.100 671.100 720.900 671.700 ;
        RECT 685.950 667.950 688.050 670.050 ;
        RECT 685.200 665.700 686.100 666.900 ;
        RECT 665.400 664.500 669.300 665.700 ;
        RECT 671.400 664.500 675.300 665.700 ;
        RECT 677.400 664.500 681.300 665.700 ;
        RECT 683.400 664.500 686.100 665.700 ;
        RECT 628.800 651.600 630.600 657.600 ;
        RECT 647.700 651.600 649.500 663.600 ;
        RECT 665.400 651.600 667.200 664.500 ;
        RECT 671.400 651.600 673.200 664.500 ;
        RECT 677.400 651.600 679.200 664.500 ;
        RECT 683.400 651.600 685.200 664.500 ;
        RECT 692.550 663.600 693.750 670.950 ;
        RECT 716.100 670.200 720.900 671.100 ;
        RECT 719.100 669.900 720.900 670.200 ;
        RECT 722.100 670.050 723.900 671.850 ;
        RECT 694.950 665.400 696.750 667.200 ;
        RECT 695.850 664.200 700.050 665.400 ;
        RECT 706.050 664.200 706.950 669.900 ;
        RECT 714.750 665.100 716.550 665.400 ;
        RECT 692.550 651.600 694.350 663.600 ;
        RECT 697.950 663.300 700.050 664.200 ;
        RECT 700.950 663.300 706.950 664.200 ;
        RECT 708.150 664.800 716.550 665.100 ;
        RECT 724.950 664.800 725.850 677.400 ;
        RECT 737.400 675.300 738.600 677.400 ;
        RECT 739.800 678.300 741.600 683.400 ;
        RECT 745.800 678.300 747.600 683.400 ;
        RECT 739.800 676.950 747.600 678.300 ;
        RECT 760.200 676.200 762.000 683.400 ;
        RECT 773.400 680.400 775.200 683.400 ;
        RECT 758.400 675.300 762.000 676.200 ;
        RECT 774.000 676.500 775.200 680.400 ;
        RECT 779.700 677.400 781.500 683.400 ;
        RECT 785.550 677.400 787.350 683.400 ;
        RECT 793.650 680.400 795.450 683.400 ;
        RECT 801.450 680.400 803.250 683.400 ;
        RECT 809.250 681.300 811.050 683.400 ;
        RECT 809.250 680.400 813.000 681.300 ;
        RECT 793.650 679.500 794.700 680.400 ;
        RECT 790.950 678.300 794.700 679.500 ;
        RECT 802.200 678.600 803.250 680.400 ;
        RECT 811.950 679.500 813.000 680.400 ;
        RECT 790.950 677.400 793.050 678.300 ;
        RECT 774.000 675.600 779.100 676.500 ;
        RECT 737.400 674.250 741.150 675.300 ;
        RECT 739.950 674.100 741.150 674.250 ;
        RECT 737.100 671.100 738.900 671.850 ;
        RECT 739.950 670.950 742.050 673.050 ;
        RECT 743.100 671.100 744.900 671.850 ;
        RECT 745.950 670.950 748.050 673.050 ;
        RECT 758.400 671.100 759.600 675.300 ;
        RECT 777.150 674.700 779.100 675.600 ;
        RECT 777.150 674.100 778.050 674.700 ;
        RECT 780.000 674.100 781.200 677.400 ;
        RECT 772.950 670.950 775.050 673.050 ;
        RECT 736.950 667.950 739.050 670.050 ;
        RECT 708.150 664.200 725.850 664.800 ;
        RECT 700.950 662.400 701.850 663.300 ;
        RECT 699.150 660.600 701.850 662.400 ;
        RECT 702.750 662.100 704.550 662.400 ;
        RECT 708.150 662.100 709.050 664.200 ;
        RECT 714.750 663.600 725.850 664.200 ;
        RECT 740.850 666.900 741.900 669.900 ;
        RECT 742.950 667.950 745.050 670.050 ;
        RECT 746.100 669.150 747.900 669.900 ;
        RECT 755.100 668.100 756.900 668.850 ;
        RECT 757.800 667.950 760.050 670.050 ;
        RECT 777.150 669.900 777.900 674.100 ;
        RECT 785.550 673.050 786.750 677.400 ;
        RECT 798.150 676.200 799.950 678.000 ;
        RECT 802.200 677.550 807.150 678.600 ;
        RECT 805.350 676.800 807.150 677.550 ;
        RECT 808.650 676.800 810.450 678.600 ;
        RECT 811.950 677.400 814.050 679.500 ;
        RECT 817.050 677.400 818.850 683.400 ;
        RECT 799.050 675.900 799.950 676.200 ;
        RECT 809.100 675.900 810.150 676.800 ;
        RECT 799.050 675.000 810.150 675.900 ;
        RECT 799.050 674.100 799.950 675.000 ;
        RECT 809.100 673.800 810.150 675.000 ;
        RECT 778.950 670.950 784.050 673.050 ;
        RECT 785.550 670.950 786.900 673.050 ;
        RECT 787.950 670.950 790.050 673.050 ;
        RECT 791.100 671.250 791.850 673.050 ;
        RECT 799.950 670.950 802.050 673.050 ;
        RECT 805.950 670.950 808.050 673.050 ;
        RECT 809.100 672.600 816.000 673.800 ;
        RECT 809.100 672.000 810.900 672.600 ;
        RECT 815.100 671.850 816.000 672.600 ;
        RECT 812.100 671.100 813.900 671.700 ;
        RECT 773.100 669.150 774.900 669.900 ;
        RECT 761.100 668.100 762.900 668.850 ;
        RECT 740.850 663.600 742.050 666.900 ;
        RECT 754.950 664.950 757.050 667.050 ;
        RECT 702.750 661.200 709.050 662.100 ;
        RECT 709.950 662.700 711.750 663.300 ;
        RECT 709.950 661.500 717.450 662.700 ;
        RECT 702.750 660.600 704.550 661.200 ;
        RECT 716.250 660.600 717.450 661.500 ;
        RECT 697.950 657.600 701.850 659.700 ;
        RECT 706.950 659.550 708.750 660.300 ;
        RECT 711.750 659.550 713.550 660.300 ;
        RECT 706.950 658.500 713.550 659.550 ;
        RECT 716.250 658.500 721.050 660.600 ;
        RECT 700.050 651.600 701.850 657.600 ;
        RECT 707.850 651.600 709.650 658.500 ;
        RECT 716.250 657.600 717.450 658.500 ;
        RECT 715.650 651.600 717.450 657.600 ;
        RECT 724.050 651.600 725.850 663.600 ;
        RECT 740.700 651.600 742.500 663.600 ;
        RECT 758.400 657.600 759.600 666.900 ;
        RECT 760.950 664.950 763.050 667.050 ;
        RECT 777.150 666.300 778.050 669.900 ;
        RECT 777.150 665.400 779.100 666.300 ;
        RECT 773.400 664.500 779.100 665.400 ;
        RECT 773.400 657.600 774.600 664.500 ;
        RECT 780.000 663.600 781.200 669.900 ;
        RECT 785.550 663.600 786.750 670.950 ;
        RECT 809.100 670.200 813.900 671.100 ;
        RECT 812.100 669.900 813.900 670.200 ;
        RECT 815.100 670.050 816.900 671.850 ;
        RECT 787.950 665.400 789.750 667.200 ;
        RECT 788.850 664.200 793.050 665.400 ;
        RECT 799.050 664.200 799.950 669.900 ;
        RECT 807.750 665.100 809.550 665.400 ;
        RECT 758.400 651.600 760.200 657.600 ;
        RECT 773.400 651.600 775.200 657.600 ;
        RECT 779.700 651.600 781.500 663.600 ;
        RECT 785.550 651.600 787.350 663.600 ;
        RECT 790.950 663.300 793.050 664.200 ;
        RECT 793.950 663.300 799.950 664.200 ;
        RECT 801.150 664.800 809.550 665.100 ;
        RECT 817.950 664.800 818.850 677.400 ;
        RECT 827.400 678.300 829.200 683.400 ;
        RECT 833.400 678.300 835.200 683.400 ;
        RECT 827.400 676.950 835.200 678.300 ;
        RECT 836.400 677.400 838.200 683.400 ;
        RECT 836.400 675.300 837.600 677.400 ;
        RECT 833.850 674.250 837.600 675.300 ;
        RECT 833.850 674.100 835.050 674.250 ;
        RECT 826.950 670.950 829.050 673.050 ;
        RECT 830.100 671.100 831.900 671.850 ;
        RECT 832.950 670.950 835.050 673.050 ;
        RECT 836.100 671.100 837.900 671.850 ;
        RECT 827.100 669.150 828.900 669.900 ;
        RECT 829.950 667.950 832.050 670.050 ;
        RECT 833.100 666.900 834.150 669.900 ;
        RECT 835.950 667.950 838.050 670.050 ;
        RECT 801.150 664.200 818.850 664.800 ;
        RECT 793.950 662.400 794.850 663.300 ;
        RECT 792.150 660.600 794.850 662.400 ;
        RECT 795.750 662.100 797.550 662.400 ;
        RECT 801.150 662.100 802.050 664.200 ;
        RECT 807.750 663.600 818.850 664.200 ;
        RECT 832.950 663.600 834.150 666.900 ;
        RECT 795.750 661.200 802.050 662.100 ;
        RECT 802.950 662.700 804.750 663.300 ;
        RECT 802.950 661.500 810.450 662.700 ;
        RECT 795.750 660.600 797.550 661.200 ;
        RECT 809.250 660.600 810.450 661.500 ;
        RECT 790.950 657.600 794.850 659.700 ;
        RECT 799.950 659.550 801.750 660.300 ;
        RECT 804.750 659.550 806.550 660.300 ;
        RECT 799.950 658.500 806.550 659.550 ;
        RECT 809.250 658.500 814.050 660.600 ;
        RECT 793.050 651.600 794.850 657.600 ;
        RECT 800.850 651.600 802.650 658.500 ;
        RECT 809.250 657.600 810.450 658.500 ;
        RECT 808.650 651.600 810.450 657.600 ;
        RECT 817.050 651.600 818.850 663.600 ;
        RECT 832.500 651.600 834.300 663.600 ;
        RECT 10.800 635.400 12.600 647.400 ;
        RECT 13.800 636.300 15.600 647.400 ;
        RECT 19.800 636.300 21.600 647.400 ;
        RECT 31.800 641.400 33.600 647.400 ;
        RECT 13.800 635.400 21.600 636.300 ;
        RECT 32.700 641.100 33.600 641.400 ;
        RECT 37.800 641.400 39.600 647.400 ;
        RECT 55.800 641.400 57.600 647.400 ;
        RECT 70.800 641.400 72.600 647.400 ;
        RECT 37.800 641.100 39.300 641.400 ;
        RECT 32.700 640.200 39.300 641.100 ;
        RECT 11.400 629.100 12.300 635.400 ;
        RECT 32.700 635.100 33.600 640.200 ;
        RECT 38.100 635.100 39.900 635.850 ;
        RECT 28.950 631.950 34.050 634.050 ;
        RECT 37.950 631.950 40.050 634.050 ;
        RECT 52.950 631.950 55.050 634.050 ;
        RECT 56.400 632.100 57.600 641.400 ;
        RECT 71.700 641.100 72.600 641.400 ;
        RECT 76.800 641.400 78.600 647.400 ;
        RECT 85.950 643.950 88.050 646.050 ;
        RECT 76.800 641.100 78.300 641.400 ;
        RECT 71.700 640.200 78.300 641.100 ;
        RECT 71.700 635.100 72.600 640.200 ;
        RECT 77.100 635.100 78.900 635.850 ;
        RECT 58.950 631.950 61.050 634.050 ;
        RECT 64.950 633.450 69.000 634.050 ;
        RECT 70.950 633.450 73.050 634.050 ;
        RECT 64.950 632.550 73.050 633.450 ;
        RECT 64.950 631.950 69.000 632.550 ;
        RECT 70.950 631.950 73.050 632.550 ;
        RECT 76.950 631.950 79.050 634.050 ;
        RECT 13.950 628.950 16.050 631.050 ;
        RECT 17.100 629.100 18.900 629.850 ;
        RECT 19.950 628.950 22.050 631.050 ;
        RECT 10.950 625.950 13.050 628.050 ;
        RECT 14.100 627.150 15.900 627.900 ;
        RECT 16.950 625.050 19.050 628.050 ;
        RECT 20.100 627.150 21.900 627.900 ;
        RECT 11.400 621.600 12.300 624.900 ;
        RECT 16.800 623.550 19.050 625.050 ;
        RECT 32.700 625.650 33.600 630.900 ;
        RECT 34.950 628.950 37.050 631.050 ;
        RECT 40.950 628.950 43.050 631.050 ;
        RECT 53.100 630.150 54.900 630.900 ;
        RECT 55.800 628.950 58.050 631.050 ;
        RECT 59.100 630.150 60.900 630.900 ;
        RECT 35.100 627.150 36.900 627.900 ;
        RECT 41.100 627.150 42.900 627.900 ;
        RECT 32.700 624.000 36.900 625.650 ;
        RECT 16.800 622.950 18.900 623.550 ;
        RECT 11.400 619.950 16.800 621.600 ;
        RECT 15.000 615.600 16.800 619.950 ;
        RECT 35.100 615.600 36.900 624.000 ;
        RECT 56.400 623.700 57.600 627.900 ;
        RECT 71.700 625.650 72.600 630.900 ;
        RECT 73.950 628.950 76.050 631.050 ;
        RECT 79.950 628.950 82.050 631.050 ;
        RECT 86.550 628.050 87.450 643.950 ;
        RECT 95.700 635.400 97.500 647.400 ;
        RECT 112.800 646.500 120.600 647.400 ;
        RECT 112.800 635.400 114.600 646.500 ;
        RECT 95.850 632.100 97.050 635.400 ;
        RECT 115.800 634.500 117.600 645.600 ;
        RECT 118.800 636.600 120.600 646.500 ;
        RECT 124.800 636.600 126.600 647.400 ;
        RECT 118.800 635.700 126.600 636.600 ;
        RECT 137.400 641.400 139.200 647.400 ;
        RECT 155.400 641.400 157.200 647.400 ;
        RECT 115.800 633.600 119.850 634.500 ;
        RECT 118.950 632.100 119.850 633.600 ;
        RECT 91.950 628.950 94.050 631.050 ;
        RECT 95.850 629.100 96.900 632.100 ;
        RECT 97.950 628.950 100.200 631.050 ;
        RECT 101.100 629.100 102.900 629.850 ;
        RECT 106.950 628.950 109.050 631.050 ;
        RECT 113.100 629.100 114.900 629.850 ;
        RECT 115.950 628.950 118.050 631.050 ;
        RECT 119.100 629.100 119.850 632.100 ;
        RECT 133.950 631.950 136.050 634.050 ;
        RECT 137.400 632.100 138.600 641.400 ;
        RECT 139.950 631.950 142.050 634.050 ;
        RECT 121.950 628.950 124.050 631.050 ;
        RECT 134.100 630.150 135.900 630.900 ;
        RECT 125.100 629.100 126.750 629.850 ;
        RECT 136.800 628.950 139.050 631.050 ;
        RECT 140.100 630.150 141.900 630.900 ;
        RECT 152.100 629.100 153.900 629.850 ;
        RECT 74.100 627.150 75.900 627.900 ;
        RECT 80.100 627.150 81.900 627.900 ;
        RECT 85.950 625.950 88.050 628.050 ;
        RECT 92.100 627.150 93.900 627.900 ;
        RECT 94.950 625.950 97.050 628.050 ;
        RECT 98.100 627.150 99.900 627.900 ;
        RECT 100.950 625.950 103.200 628.050 ;
        RECT 71.700 624.000 75.900 625.650 ;
        RECT 94.950 624.750 96.150 624.900 ;
        RECT 54.000 622.800 57.600 623.700 ;
        RECT 54.000 615.600 55.800 622.800 ;
        RECT 74.100 615.600 75.900 624.000 ;
        RECT 92.400 623.700 96.150 624.750 ;
        RECT 92.400 621.600 93.600 623.700 ;
        RECT 91.800 615.600 93.600 621.600 ;
        RECT 94.800 620.700 102.600 622.050 ;
        RECT 94.800 615.600 96.600 620.700 ;
        RECT 100.800 615.600 102.600 620.700 ;
        RECT 107.550 619.050 108.450 628.950 ;
        RECT 112.800 625.950 115.050 628.050 ;
        RECT 116.250 627.150 117.900 627.900 ;
        RECT 118.950 625.950 121.200 628.050 ;
        RECT 122.100 627.150 123.750 627.900 ;
        RECT 124.950 625.950 127.200 628.050 ;
        RECT 120.000 621.600 121.050 624.900 ;
        RECT 137.400 623.700 138.600 627.900 ;
        RECT 151.950 625.950 154.050 628.050 ;
        RECT 155.400 624.300 156.450 641.400 ;
        RECT 162.000 635.400 163.800 647.400 ;
        RECT 166.950 643.950 169.050 646.050 ;
        RECT 157.950 628.950 160.050 631.050 ;
        RECT 162.000 629.100 163.050 635.400 ;
        RECT 158.100 627.150 159.900 627.900 ;
        RECT 160.950 627.450 163.050 628.050 ;
        RECT 167.550 627.450 168.450 643.950 ;
        RECT 175.800 641.400 177.600 647.400 ;
        RECT 176.700 641.100 177.600 641.400 ;
        RECT 181.800 641.400 183.600 647.400 ;
        RECT 196.800 641.400 198.600 647.400 ;
        RECT 211.800 641.400 213.600 647.400 ;
        RECT 181.800 641.100 183.300 641.400 ;
        RECT 176.700 640.200 183.300 641.100 ;
        RECT 176.700 635.100 177.600 640.200 ;
        RECT 182.100 635.100 183.900 635.850 ;
        RECT 172.950 631.950 178.050 634.050 ;
        RECT 181.800 631.950 184.050 634.050 ;
        RECT 197.400 632.100 198.600 641.400 ;
        RECT 205.950 634.950 208.050 637.050 ;
        RECT 160.950 626.550 168.450 627.450 ;
        RECT 160.950 625.950 163.050 626.550 ;
        RECT 176.700 625.650 177.600 630.900 ;
        RECT 178.950 628.950 181.050 631.050 ;
        RECT 184.950 628.950 187.050 631.050 ;
        RECT 193.950 628.950 199.050 631.050 ;
        RECT 206.550 630.450 207.450 634.950 ;
        RECT 212.400 632.100 213.600 641.400 ;
        RECT 230.700 635.400 232.500 647.400 ;
        RECT 247.800 641.400 249.600 647.400 ;
        RECT 248.700 641.100 249.600 641.400 ;
        RECT 253.800 641.400 255.600 647.400 ;
        RECT 269.400 641.400 271.200 647.400 ;
        RECT 253.800 641.100 255.300 641.400 ;
        RECT 248.700 640.200 255.300 641.100 ;
        RECT 241.950 637.950 244.050 640.050 ;
        RECT 230.850 632.100 232.050 635.400 ;
        RECT 211.950 630.450 214.050 631.050 ;
        RECT 206.550 629.550 214.050 630.450 ;
        RECT 211.950 628.950 214.050 629.550 ;
        RECT 226.950 628.950 229.050 631.050 ;
        RECT 230.850 629.100 231.900 632.100 ;
        RECT 232.950 628.950 235.050 631.050 ;
        RECT 236.100 629.100 237.900 629.850 ;
        RECT 179.100 627.150 180.900 627.900 ;
        RECT 185.100 627.150 186.900 627.900 ;
        RECT 137.400 622.800 141.000 623.700 ;
        RECT 106.950 616.950 109.050 619.050 ;
        RECT 120.000 615.600 121.800 621.600 ;
        RECT 139.200 615.600 141.000 622.800 ;
        RECT 152.400 623.100 159.900 624.300 ;
        RECT 152.400 615.600 154.200 623.100 ;
        RECT 158.100 622.500 159.900 623.100 ;
        RECT 160.950 621.600 161.850 624.900 ;
        RECT 176.700 624.000 180.900 625.650 ;
        RECT 159.900 619.800 161.850 621.600 ;
        RECT 159.900 615.600 161.700 619.800 ;
        RECT 179.100 615.600 180.900 624.000 ;
        RECT 197.400 618.600 198.600 627.900 ;
        RECT 200.100 626.100 201.900 626.850 ;
        RECT 199.950 622.950 202.050 625.050 ;
        RECT 212.400 618.600 213.600 627.900 ;
        RECT 227.100 627.150 228.900 627.900 ;
        RECT 215.100 626.100 216.900 626.850 ;
        RECT 229.950 625.950 232.050 628.050 ;
        RECT 233.100 627.150 234.900 627.900 ;
        RECT 235.950 625.950 238.050 628.050 ;
        RECT 214.950 622.950 217.050 625.050 ;
        RECT 229.950 624.750 231.150 624.900 ;
        RECT 227.400 623.700 231.150 624.750 ;
        RECT 227.400 621.600 228.600 623.700 ;
        RECT 242.550 622.050 243.450 637.950 ;
        RECT 248.700 635.100 249.600 640.200 ;
        RECT 254.100 635.100 255.900 635.850 ;
        RECT 244.950 631.950 250.050 634.050 ;
        RECT 253.950 631.950 256.050 634.050 ;
        RECT 265.950 631.950 268.050 634.050 ;
        RECT 269.400 632.100 270.600 641.400 ;
        RECT 290.700 635.400 292.500 647.400 ;
        RECT 308.400 641.400 310.200 647.400 ;
        RECT 271.950 631.950 274.200 634.050 ;
        RECT 290.850 632.100 292.050 635.400 ;
        RECT 248.700 625.650 249.600 630.900 ;
        RECT 250.950 628.950 253.050 631.050 ;
        RECT 256.950 628.950 259.200 631.050 ;
        RECT 266.100 630.150 267.900 630.900 ;
        RECT 268.800 628.950 271.050 631.050 ;
        RECT 272.100 630.150 273.900 630.900 ;
        RECT 286.800 628.950 289.050 631.050 ;
        RECT 290.850 629.100 291.900 632.100 ;
        RECT 304.950 631.950 307.050 634.050 ;
        RECT 308.400 632.100 309.600 641.400 ;
        RECT 329.700 635.400 331.500 647.400 ;
        RECT 349.500 635.400 351.300 647.400 ;
        RECT 358.950 640.950 361.050 643.050 ;
        RECT 310.950 631.950 313.050 634.050 ;
        RECT 329.850 632.100 331.050 635.400 ;
        RECT 349.950 632.100 351.150 635.400 ;
        RECT 292.950 628.950 295.050 631.050 ;
        RECT 305.100 630.150 306.900 630.900 ;
        RECT 296.100 629.100 297.900 629.850 ;
        RECT 307.800 628.950 310.050 631.050 ;
        RECT 311.100 630.150 312.900 630.900 ;
        RECT 325.950 628.950 328.050 631.050 ;
        RECT 329.850 629.100 330.900 632.100 ;
        RECT 331.950 628.950 334.050 631.050 ;
        RECT 335.100 629.100 336.900 629.850 ;
        RECT 344.100 629.100 345.900 629.850 ;
        RECT 346.950 628.950 349.200 631.050 ;
        RECT 350.100 629.100 351.150 632.100 ;
        RECT 359.550 631.050 360.450 640.950 ;
        RECT 361.950 634.950 364.050 637.050 ;
        RECT 367.200 635.400 369.000 647.400 ;
        RECT 373.800 641.400 375.600 647.400 ;
        RECT 352.950 628.950 355.050 631.050 ;
        RECT 358.950 628.950 361.050 631.050 ;
        RECT 251.100 627.150 252.900 627.900 ;
        RECT 257.100 627.150 258.900 627.900 ;
        RECT 248.700 624.000 252.900 625.650 ;
        RECT 196.800 615.600 198.600 618.600 ;
        RECT 211.800 615.600 213.600 618.600 ;
        RECT 226.800 615.600 228.600 621.600 ;
        RECT 229.800 620.700 237.600 622.050 ;
        RECT 229.800 615.600 231.600 620.700 ;
        RECT 235.800 615.600 237.600 620.700 ;
        RECT 242.550 620.550 247.050 622.050 ;
        RECT 243.000 619.950 247.050 620.550 ;
        RECT 251.100 615.600 252.900 624.000 ;
        RECT 269.400 623.700 270.600 627.900 ;
        RECT 287.100 627.150 288.900 627.900 ;
        RECT 289.950 625.950 292.050 628.050 ;
        RECT 293.100 627.150 294.900 627.900 ;
        RECT 295.950 625.950 298.050 628.050 ;
        RECT 289.950 624.750 291.150 624.900 ;
        RECT 287.400 623.700 291.150 624.750 ;
        RECT 308.400 623.700 309.600 627.900 ;
        RECT 320.100 625.950 322.200 628.050 ;
        RECT 326.100 627.150 327.900 627.900 ;
        RECT 328.950 625.950 331.050 628.050 ;
        RECT 332.100 627.150 333.900 627.900 ;
        RECT 334.950 625.950 337.050 628.050 ;
        RECT 343.950 625.950 346.050 628.050 ;
        RECT 347.100 627.150 348.900 627.900 ;
        RECT 349.950 625.950 352.050 628.050 ;
        RECT 353.100 627.150 354.900 627.900 ;
        RECT 269.400 622.800 273.000 623.700 ;
        RECT 271.200 615.600 273.000 622.800 ;
        RECT 287.400 621.600 288.600 623.700 ;
        RECT 308.400 622.800 312.000 623.700 ;
        RECT 286.800 615.600 288.600 621.600 ;
        RECT 289.800 620.700 297.600 622.050 ;
        RECT 289.800 615.600 291.600 620.700 ;
        RECT 295.800 615.600 297.600 620.700 ;
        RECT 310.200 615.600 312.000 622.800 ;
        RECT 320.550 622.050 321.450 625.950 ;
        RECT 362.550 625.050 363.450 634.950 ;
        RECT 367.950 629.100 369.000 635.400 ;
        RECT 370.950 628.950 373.050 631.050 ;
        RECT 364.950 625.950 370.050 628.050 ;
        RECT 371.100 627.150 372.900 627.900 ;
        RECT 328.950 624.750 330.150 624.900 ;
        RECT 326.400 623.700 330.150 624.750 ;
        RECT 350.850 624.750 352.050 624.900 ;
        RECT 350.850 623.700 354.600 624.750 ;
        RECT 319.950 619.950 322.050 622.050 ;
        RECT 326.400 621.600 327.600 623.700 ;
        RECT 325.800 615.600 327.600 621.600 ;
        RECT 328.800 620.700 336.600 622.050 ;
        RECT 328.800 615.600 330.600 620.700 ;
        RECT 334.800 615.600 336.600 620.700 ;
        RECT 344.400 620.700 352.200 622.050 ;
        RECT 344.400 615.600 346.200 620.700 ;
        RECT 350.400 615.600 352.200 620.700 ;
        RECT 353.400 621.600 354.600 623.700 ;
        RECT 361.950 622.950 364.050 625.050 ;
        RECT 369.150 621.600 370.050 624.900 ;
        RECT 374.550 624.300 375.600 641.400 ;
        RECT 386.400 636.600 388.200 647.400 ;
        RECT 392.400 646.500 400.200 647.400 ;
        RECT 392.400 636.600 394.200 646.500 ;
        RECT 386.400 635.700 394.200 636.600 ;
        RECT 395.400 634.500 397.200 645.600 ;
        RECT 398.400 635.400 400.200 646.500 ;
        RECT 403.950 643.950 406.050 646.050 ;
        RECT 393.150 633.600 397.200 634.500 ;
        RECT 393.150 632.100 394.050 633.600 ;
        RECT 377.100 629.100 378.900 629.850 ;
        RECT 386.250 629.100 387.900 629.850 ;
        RECT 388.950 628.950 391.050 631.050 ;
        RECT 393.150 629.100 393.900 632.100 ;
        RECT 394.950 628.950 397.200 631.050 ;
        RECT 398.100 629.100 399.900 629.850 ;
        RECT 404.550 628.050 405.450 643.950 ;
        RECT 410.400 636.600 412.200 647.400 ;
        RECT 416.400 646.500 424.200 647.400 ;
        RECT 416.400 636.600 418.200 646.500 ;
        RECT 410.400 635.700 418.200 636.600 ;
        RECT 419.400 634.500 421.200 645.600 ;
        RECT 422.400 635.400 424.200 646.500 ;
        RECT 437.400 641.400 439.200 647.400 ;
        RECT 454.800 641.400 456.600 647.400 ;
        RECT 417.150 633.600 421.200 634.500 ;
        RECT 417.150 632.100 418.050 633.600 ;
        RECT 437.400 632.100 438.600 641.400 ;
        RECT 410.250 629.100 411.900 629.850 ;
        RECT 412.950 628.950 415.050 631.050 ;
        RECT 417.150 629.100 417.900 632.100 ;
        RECT 451.950 631.950 454.050 634.050 ;
        RECT 455.400 632.100 456.600 641.400 ;
        RECT 463.950 640.950 466.050 643.050 ;
        RECT 457.950 631.950 460.050 634.050 ;
        RECT 418.950 628.950 421.050 631.050 ;
        RECT 436.950 630.450 439.050 631.050 ;
        RECT 422.100 629.100 423.900 629.850 ;
        RECT 436.950 629.550 444.450 630.450 ;
        RECT 452.100 630.150 453.900 630.900 ;
        RECT 436.950 628.950 439.050 629.550 ;
        RECT 376.950 625.950 379.050 628.050 ;
        RECT 385.950 625.950 388.050 628.050 ;
        RECT 389.250 627.150 390.900 627.900 ;
        RECT 391.950 625.950 394.050 628.050 ;
        RECT 395.100 627.150 396.750 627.900 ;
        RECT 397.950 625.950 400.050 628.050 ;
        RECT 404.100 625.950 406.200 628.050 ;
        RECT 409.800 625.950 412.050 628.050 ;
        RECT 413.250 627.150 414.900 627.900 ;
        RECT 415.800 625.950 418.050 628.050 ;
        RECT 419.100 627.150 420.750 627.900 ;
        RECT 421.950 625.950 424.200 628.050 ;
        RECT 434.100 626.100 435.900 626.850 ;
        RECT 371.100 623.100 378.600 624.300 ;
        RECT 371.100 622.500 372.900 623.100 ;
        RECT 353.400 615.600 355.200 621.600 ;
        RECT 369.150 619.800 371.100 621.600 ;
        RECT 369.300 615.600 371.100 619.800 ;
        RECT 376.800 615.600 378.600 623.100 ;
        RECT 391.950 621.600 393.000 624.900 ;
        RECT 404.550 622.050 405.450 625.950 ;
        RECT 391.200 615.600 393.000 621.600 ;
        RECT 403.950 619.950 406.050 622.050 ;
        RECT 415.950 621.600 417.000 624.900 ;
        RECT 433.950 622.950 436.050 625.050 ;
        RECT 415.200 615.600 417.000 621.600 ;
        RECT 437.400 618.600 438.600 627.900 ;
        RECT 443.550 619.050 444.450 629.550 ;
        RECT 454.950 628.950 457.050 631.050 ;
        RECT 458.100 630.150 459.900 630.900 ;
        RECT 455.400 623.700 456.600 627.900 ;
        RECT 464.550 627.450 465.450 640.950 ;
        RECT 469.200 635.400 471.000 647.400 ;
        RECT 475.800 641.400 477.600 647.400 ;
        RECT 469.950 629.100 471.000 635.400 ;
        RECT 472.950 628.950 475.050 631.050 ;
        RECT 469.950 627.450 472.050 628.050 ;
        RECT 464.550 626.550 472.050 627.450 ;
        RECT 473.100 627.150 474.900 627.900 ;
        RECT 469.950 625.950 472.050 626.550 ;
        RECT 453.000 622.800 456.600 623.700 ;
        RECT 437.400 615.600 439.200 618.600 ;
        RECT 442.950 616.950 445.050 619.050 ;
        RECT 453.000 615.600 454.800 622.800 ;
        RECT 471.150 621.600 472.050 624.900 ;
        RECT 476.550 624.300 477.600 641.400 ;
        RECT 484.950 640.950 487.050 643.050 ;
        RECT 479.100 629.100 480.900 629.850 ;
        RECT 478.950 625.950 481.050 628.050 ;
        RECT 485.550 625.050 486.450 640.950 ;
        RECT 494.700 635.400 496.500 647.400 ;
        RECT 514.500 635.400 516.300 647.400 ;
        RECT 532.800 641.400 534.600 647.400 ;
        RECT 550.800 641.400 552.600 647.400 ;
        RECT 494.850 632.100 496.050 635.400 ;
        RECT 514.950 632.100 516.150 635.400 ;
        RECT 533.400 632.100 534.600 641.400 ;
        RECT 490.800 628.950 493.050 631.050 ;
        RECT 494.850 629.100 495.900 632.100 ;
        RECT 496.950 628.950 499.200 631.050 ;
        RECT 500.100 629.100 501.900 629.850 ;
        RECT 509.100 629.100 510.900 629.850 ;
        RECT 511.950 628.950 514.050 631.050 ;
        RECT 515.100 629.100 516.150 632.100 ;
        RECT 547.950 631.950 550.050 634.050 ;
        RECT 551.400 632.100 552.600 641.400 ;
        RECT 566.400 641.400 568.200 647.400 ;
        RECT 586.800 641.400 588.600 647.400 ;
        RECT 553.950 631.950 556.050 634.050 ;
        RECT 562.950 631.950 565.050 634.050 ;
        RECT 566.400 632.100 567.600 641.400 ;
        RECT 568.950 631.950 571.050 634.050 ;
        RECT 583.950 631.950 586.050 634.050 ;
        RECT 587.400 632.100 588.600 641.400 ;
        RECT 602.400 641.400 604.200 647.400 ;
        RECT 589.950 631.950 592.050 634.050 ;
        RECT 602.400 632.100 603.600 641.400 ;
        RECT 607.950 640.950 610.050 643.050 ;
        RECT 614.400 641.400 616.200 647.400 ;
        RECT 517.950 628.950 520.050 631.050 ;
        RECT 529.950 628.950 535.050 631.050 ;
        RECT 548.100 630.150 549.900 630.900 ;
        RECT 550.950 628.950 553.050 631.050 ;
        RECT 554.100 630.150 555.900 630.900 ;
        RECT 563.100 630.150 564.900 630.900 ;
        RECT 565.950 628.950 568.050 631.050 ;
        RECT 569.100 630.150 570.900 630.900 ;
        RECT 584.100 630.150 585.900 630.900 ;
        RECT 586.950 628.950 589.050 631.050 ;
        RECT 590.100 630.150 591.900 630.900 ;
        RECT 601.950 628.950 604.050 631.050 ;
        RECT 491.100 627.150 492.900 627.900 ;
        RECT 493.950 625.950 496.200 628.050 ;
        RECT 497.100 627.150 498.900 627.900 ;
        RECT 499.950 625.950 502.050 628.050 ;
        RECT 508.800 625.950 511.050 628.050 ;
        RECT 512.100 627.150 513.900 627.900 ;
        RECT 514.950 625.950 517.050 628.050 ;
        RECT 518.100 627.150 519.900 627.900 ;
        RECT 473.100 623.100 480.600 624.300 ;
        RECT 473.100 622.500 474.900 623.100 ;
        RECT 471.150 619.800 473.100 621.600 ;
        RECT 471.300 615.600 473.100 619.800 ;
        RECT 478.800 615.600 480.600 623.100 ;
        RECT 484.950 622.950 487.050 625.050 ;
        RECT 493.950 624.750 495.150 624.900 ;
        RECT 491.400 623.700 495.150 624.750 ;
        RECT 515.850 624.750 517.050 624.900 ;
        RECT 515.850 623.700 519.600 624.750 ;
        RECT 491.400 621.600 492.600 623.700 ;
        RECT 490.800 615.600 492.600 621.600 ;
        RECT 493.800 620.700 501.600 622.050 ;
        RECT 493.800 615.600 495.600 620.700 ;
        RECT 499.800 615.600 501.600 620.700 ;
        RECT 509.400 620.700 517.200 622.050 ;
        RECT 509.400 615.600 511.200 620.700 ;
        RECT 515.400 615.600 517.200 620.700 ;
        RECT 518.400 621.600 519.600 623.700 ;
        RECT 518.400 615.600 520.200 621.600 ;
        RECT 533.400 618.600 534.600 627.900 ;
        RECT 536.100 626.100 537.900 626.850 ;
        RECT 535.950 622.950 538.050 625.050 ;
        RECT 551.400 623.700 552.600 627.900 ;
        RECT 532.800 615.600 534.600 618.600 ;
        RECT 549.000 622.800 552.600 623.700 ;
        RECT 566.400 623.700 567.600 627.900 ;
        RECT 587.400 623.700 588.600 627.900 ;
        RECT 599.100 626.100 600.900 626.850 ;
        RECT 566.400 622.800 570.000 623.700 ;
        RECT 549.000 615.600 550.800 622.800 ;
        RECT 568.200 615.600 570.000 622.800 ;
        RECT 585.000 622.800 588.600 623.700 ;
        RECT 598.950 622.950 601.050 625.050 ;
        RECT 585.000 615.600 586.800 622.800 ;
        RECT 602.400 618.600 603.600 627.900 ;
        RECT 608.550 622.050 609.450 640.950 ;
        RECT 614.400 634.500 615.600 641.400 ;
        RECT 620.700 635.400 622.500 647.400 ;
        RECT 635.400 641.400 637.200 647.400 ;
        RECT 625.950 637.950 628.050 640.050 ;
        RECT 614.400 633.600 620.100 634.500 ;
        RECT 618.150 632.700 620.100 633.600 ;
        RECT 614.100 629.100 615.900 629.850 ;
        RECT 618.150 629.100 619.050 632.700 ;
        RECT 621.000 629.100 622.200 635.400 ;
        RECT 626.550 634.050 627.450 637.950 ;
        RECT 625.950 631.950 628.050 634.050 ;
        RECT 631.950 631.950 634.050 634.050 ;
        RECT 635.400 632.100 636.600 641.400 ;
        RECT 656.700 635.400 658.500 647.400 ;
        RECT 665.550 635.400 667.350 647.400 ;
        RECT 673.050 641.400 674.850 647.400 ;
        RECT 670.950 639.300 674.850 641.400 ;
        RECT 680.850 640.500 682.650 647.400 ;
        RECT 688.650 641.400 690.450 647.400 ;
        RECT 689.250 640.500 690.450 641.400 ;
        RECT 679.950 639.450 686.550 640.500 ;
        RECT 679.950 638.700 681.750 639.450 ;
        RECT 684.750 638.700 686.550 639.450 ;
        RECT 689.250 638.400 694.050 640.500 ;
        RECT 672.150 636.600 674.850 638.400 ;
        RECT 675.750 637.800 677.550 638.400 ;
        RECT 675.750 636.900 682.050 637.800 ;
        RECT 689.250 637.500 690.450 638.400 ;
        RECT 675.750 636.600 677.550 636.900 ;
        RECT 673.950 635.700 674.850 636.600 ;
        RECT 637.950 631.950 640.050 634.050 ;
        RECT 656.850 632.100 658.050 635.400 ;
        RECT 613.950 625.950 616.050 628.050 ;
        RECT 618.150 624.900 618.900 629.100 ;
        RECT 619.950 627.450 622.050 628.050 ;
        RECT 626.550 627.450 627.450 631.950 ;
        RECT 632.100 630.150 633.900 630.900 ;
        RECT 634.950 628.950 637.050 631.050 ;
        RECT 638.100 630.150 639.900 630.900 ;
        RECT 652.800 628.950 655.050 631.050 ;
        RECT 656.850 629.100 657.900 632.100 ;
        RECT 658.800 628.950 661.050 631.050 ;
        RECT 662.100 629.100 663.900 629.850 ;
        RECT 665.550 628.050 666.750 635.400 ;
        RECT 670.950 634.800 673.050 635.700 ;
        RECT 673.950 634.800 679.950 635.700 ;
        RECT 668.850 633.600 673.050 634.800 ;
        RECT 667.950 631.800 669.750 633.600 ;
        RECT 679.050 629.100 679.950 634.800 ;
        RECT 681.150 634.800 682.050 636.900 ;
        RECT 682.950 636.300 690.450 637.500 ;
        RECT 682.950 635.700 684.750 636.300 ;
        RECT 697.050 635.400 698.850 647.400 ;
        RECT 709.500 635.400 711.300 647.400 ;
        RECT 715.800 641.400 717.600 647.400 ;
        RECT 687.750 634.800 698.850 635.400 ;
        RECT 681.150 634.200 698.850 634.800 ;
        RECT 681.150 633.900 689.550 634.200 ;
        RECT 687.750 633.600 689.550 633.900 ;
        RECT 619.950 626.550 627.450 627.450 ;
        RECT 619.950 625.950 622.050 626.550 ;
        RECT 618.150 624.300 619.050 624.900 ;
        RECT 618.150 623.400 620.100 624.300 ;
        RECT 615.000 622.500 620.100 623.400 ;
        RECT 607.950 619.950 610.050 622.050 ;
        RECT 615.000 618.600 616.200 622.500 ;
        RECT 621.000 621.600 622.200 624.900 ;
        RECT 635.400 623.700 636.600 627.900 ;
        RECT 653.100 627.150 654.900 627.900 ;
        RECT 655.950 625.950 658.050 628.050 ;
        RECT 659.100 627.150 660.900 627.900 ;
        RECT 661.950 625.950 664.050 628.050 ;
        RECT 665.550 625.950 666.900 628.050 ;
        RECT 667.950 625.950 670.050 628.050 ;
        RECT 671.100 625.950 671.850 627.750 ;
        RECT 679.950 625.950 682.050 628.050 ;
        RECT 685.950 625.950 688.050 631.050 ;
        RECT 692.100 628.800 693.900 629.100 ;
        RECT 689.100 627.900 693.900 628.800 ;
        RECT 692.100 627.300 693.900 627.900 ;
        RECT 695.100 627.150 696.900 628.950 ;
        RECT 689.100 626.400 690.900 627.000 ;
        RECT 695.100 626.400 696.000 627.150 ;
        RECT 655.950 624.750 657.150 624.900 ;
        RECT 653.400 623.700 657.150 624.750 ;
        RECT 635.400 622.800 639.000 623.700 ;
        RECT 602.400 615.600 604.200 618.600 ;
        RECT 614.400 615.600 616.200 618.600 ;
        RECT 620.700 615.600 622.500 621.600 ;
        RECT 637.200 615.600 639.000 622.800 ;
        RECT 653.400 621.600 654.600 623.700 ;
        RECT 652.800 615.600 654.600 621.600 ;
        RECT 655.800 620.700 663.600 622.050 ;
        RECT 655.800 615.600 657.600 620.700 ;
        RECT 661.800 615.600 663.600 620.700 ;
        RECT 665.550 621.600 666.750 625.950 ;
        RECT 689.100 625.200 696.000 626.400 ;
        RECT 679.050 624.000 679.950 624.900 ;
        RECT 689.100 624.000 690.150 625.200 ;
        RECT 679.050 623.100 690.150 624.000 ;
        RECT 679.050 622.800 679.950 623.100 ;
        RECT 665.550 615.600 667.350 621.600 ;
        RECT 670.950 620.700 673.050 621.600 ;
        RECT 678.150 621.000 679.950 622.800 ;
        RECT 689.100 622.200 690.150 623.100 ;
        RECT 685.350 621.450 687.150 622.200 ;
        RECT 670.950 619.500 674.700 620.700 ;
        RECT 673.650 618.600 674.700 619.500 ;
        RECT 682.200 620.400 687.150 621.450 ;
        RECT 688.650 620.400 690.450 622.200 ;
        RECT 697.950 621.600 698.850 634.200 ;
        RECT 709.800 629.100 711.000 635.400 ;
        RECT 716.400 634.500 717.600 641.400 ;
        RECT 711.900 633.600 717.600 634.500 ;
        RECT 720.150 635.400 721.950 647.400 ;
        RECT 728.550 641.400 730.350 647.400 ;
        RECT 728.550 640.500 729.750 641.400 ;
        RECT 736.350 640.500 738.150 647.400 ;
        RECT 744.150 641.400 745.950 647.400 ;
        RECT 724.950 638.400 729.750 640.500 ;
        RECT 732.450 639.450 739.050 640.500 ;
        RECT 732.450 638.700 734.250 639.450 ;
        RECT 737.250 638.700 739.050 639.450 ;
        RECT 744.150 639.300 748.050 641.400 ;
        RECT 728.550 637.500 729.750 638.400 ;
        RECT 741.450 637.800 743.250 638.400 ;
        RECT 728.550 636.300 736.050 637.500 ;
        RECT 734.250 635.700 736.050 636.300 ;
        RECT 736.950 636.900 743.250 637.800 ;
        RECT 720.150 634.800 731.250 635.400 ;
        RECT 736.950 634.800 737.850 636.900 ;
        RECT 741.450 636.600 743.250 636.900 ;
        RECT 744.150 636.600 746.850 638.400 ;
        RECT 744.150 635.700 745.050 636.600 ;
        RECT 720.150 634.200 737.850 634.800 ;
        RECT 711.900 632.700 713.850 633.600 ;
        RECT 712.950 629.100 713.850 632.700 ;
        RECT 716.100 629.100 717.900 629.850 ;
        RECT 706.800 625.950 712.050 628.050 ;
        RECT 713.100 624.900 713.850 629.100 ;
        RECT 715.950 625.950 718.050 628.050 ;
        RECT 709.800 621.600 711.000 624.900 ;
        RECT 712.950 624.300 713.850 624.900 ;
        RECT 711.900 623.400 713.850 624.300 ;
        RECT 711.900 622.500 717.000 623.400 ;
        RECT 682.200 618.600 683.250 620.400 ;
        RECT 691.950 619.500 694.050 621.600 ;
        RECT 691.950 618.600 693.000 619.500 ;
        RECT 673.650 615.600 675.450 618.600 ;
        RECT 681.450 615.600 683.250 618.600 ;
        RECT 689.250 617.700 693.000 618.600 ;
        RECT 689.250 615.600 691.050 617.700 ;
        RECT 697.050 615.600 698.850 621.600 ;
        RECT 709.500 615.600 711.300 621.600 ;
        RECT 715.800 618.600 717.000 622.500 ;
        RECT 720.150 621.600 721.050 634.200 ;
        RECT 729.450 633.900 737.850 634.200 ;
        RECT 739.050 634.800 745.050 635.700 ;
        RECT 745.950 634.800 748.050 635.700 ;
        RECT 751.650 635.400 753.450 647.400 ;
        RECT 729.450 633.600 731.250 633.900 ;
        RECT 739.050 629.100 739.950 634.800 ;
        RECT 745.950 633.600 750.150 634.800 ;
        RECT 749.250 631.800 751.050 633.600 ;
        RECT 722.100 627.150 723.900 628.950 ;
        RECT 725.100 628.800 726.900 629.100 ;
        RECT 725.100 627.900 729.900 628.800 ;
        RECT 752.250 628.050 753.450 635.400 ;
        RECT 761.400 641.400 763.200 647.400 ;
        RECT 761.400 634.500 762.600 641.400 ;
        RECT 767.700 635.400 769.500 647.400 ;
        RECT 784.500 635.400 786.300 647.400 ;
        RECT 803.400 641.400 805.200 647.400 ;
        RECT 823.800 641.400 825.600 647.400 ;
        RECT 761.400 633.600 767.100 634.500 ;
        RECT 765.150 632.700 767.100 633.600 ;
        RECT 761.100 629.100 762.900 629.850 ;
        RECT 765.150 629.100 766.050 632.700 ;
        RECT 768.000 629.100 769.200 635.400 ;
        RECT 784.950 632.100 786.150 635.400 ;
        RECT 779.100 629.100 780.900 629.850 ;
        RECT 725.100 627.300 726.900 627.900 ;
        RECT 723.000 626.400 723.900 627.150 ;
        RECT 728.100 626.400 729.900 627.000 ;
        RECT 723.000 625.200 729.900 626.400 ;
        RECT 730.950 625.950 733.050 628.050 ;
        RECT 736.950 625.950 739.050 628.050 ;
        RECT 747.150 625.950 747.900 627.750 ;
        RECT 748.950 625.950 751.050 628.050 ;
        RECT 752.100 625.950 753.450 628.050 ;
        RECT 760.950 625.950 763.050 628.050 ;
        RECT 728.850 624.000 729.900 625.200 ;
        RECT 739.050 624.000 739.950 624.900 ;
        RECT 728.850 623.100 739.950 624.000 ;
        RECT 728.850 622.200 729.900 623.100 ;
        RECT 739.050 622.800 739.950 623.100 ;
        RECT 715.800 615.600 717.600 618.600 ;
        RECT 720.150 615.600 721.950 621.600 ;
        RECT 724.950 619.500 727.050 621.600 ;
        RECT 728.550 620.400 730.350 622.200 ;
        RECT 731.850 621.450 733.650 622.200 ;
        RECT 731.850 620.400 736.800 621.450 ;
        RECT 739.050 621.000 740.850 622.800 ;
        RECT 752.250 621.600 753.450 625.950 ;
        RECT 765.150 624.900 765.900 629.100 ;
        RECT 781.950 628.950 784.050 631.050 ;
        RECT 785.100 629.100 786.150 632.100 ;
        RECT 799.950 631.950 802.050 634.050 ;
        RECT 803.400 632.100 804.600 641.400 ;
        RECT 805.950 631.950 808.050 634.050 ;
        RECT 820.950 631.950 823.050 634.050 ;
        RECT 824.400 632.100 825.600 641.400 ;
        RECT 841.500 635.400 843.300 647.400 ;
        RECT 826.950 631.950 829.050 634.050 ;
        RECT 841.950 632.100 843.150 635.400 ;
        RECT 787.950 628.950 790.050 631.050 ;
        RECT 800.100 630.150 801.900 630.900 ;
        RECT 802.950 628.950 805.050 631.050 ;
        RECT 806.100 630.150 807.900 630.900 ;
        RECT 821.100 630.150 822.900 630.900 ;
        RECT 823.800 628.950 826.050 631.050 ;
        RECT 827.100 630.150 828.900 630.900 ;
        RECT 836.100 629.100 837.900 629.850 ;
        RECT 838.950 628.950 841.050 631.050 ;
        RECT 842.100 629.100 843.150 632.100 ;
        RECT 844.950 628.950 847.050 631.050 ;
        RECT 766.950 627.450 769.050 628.050 ;
        RECT 771.000 627.450 774.900 628.050 ;
        RECT 766.950 626.550 774.900 627.450 ;
        RECT 766.950 625.950 769.050 626.550 ;
        RECT 771.000 625.950 774.900 626.550 ;
        RECT 778.950 625.950 781.050 628.050 ;
        RECT 782.100 627.150 783.900 627.900 ;
        RECT 784.950 625.950 787.050 628.050 ;
        RECT 788.100 627.150 789.900 627.900 ;
        RECT 765.150 624.300 766.050 624.900 ;
        RECT 765.150 623.400 767.100 624.300 ;
        RECT 745.950 620.700 748.050 621.600 ;
        RECT 726.000 618.600 727.050 619.500 ;
        RECT 735.750 618.600 736.800 620.400 ;
        RECT 744.300 619.500 748.050 620.700 ;
        RECT 744.300 618.600 745.350 619.500 ;
        RECT 726.000 617.700 729.750 618.600 ;
        RECT 727.950 615.600 729.750 617.700 ;
        RECT 735.750 615.600 737.550 618.600 ;
        RECT 743.550 615.600 745.350 618.600 ;
        RECT 751.650 615.600 753.450 621.600 ;
        RECT 762.000 622.500 767.100 623.400 ;
        RECT 762.000 618.600 763.200 622.500 ;
        RECT 768.000 621.600 769.200 624.900 ;
        RECT 785.850 624.750 787.050 624.900 ;
        RECT 785.850 623.700 789.600 624.750 ;
        RECT 761.400 615.600 763.200 618.600 ;
        RECT 767.700 615.600 769.500 621.600 ;
        RECT 779.400 620.700 787.200 622.050 ;
        RECT 779.400 615.600 781.200 620.700 ;
        RECT 785.400 615.600 787.200 620.700 ;
        RECT 788.400 621.600 789.600 623.700 ;
        RECT 803.400 623.700 804.600 627.900 ;
        RECT 824.400 623.700 825.600 627.900 ;
        RECT 835.950 625.950 838.050 628.050 ;
        RECT 839.100 627.150 840.900 627.900 ;
        RECT 841.950 625.950 844.050 628.050 ;
        RECT 845.100 627.150 846.900 627.900 ;
        RECT 842.850 624.750 844.050 624.900 ;
        RECT 842.850 623.700 846.600 624.750 ;
        RECT 803.400 622.800 807.000 623.700 ;
        RECT 788.400 615.600 790.200 621.600 ;
        RECT 805.200 615.600 807.000 622.800 ;
        RECT 822.000 622.800 825.600 623.700 ;
        RECT 822.000 615.600 823.800 622.800 ;
        RECT 836.400 620.700 844.200 622.050 ;
        RECT 836.400 615.600 838.200 620.700 ;
        RECT 842.400 615.600 844.200 620.700 ;
        RECT 845.400 621.600 846.600 623.700 ;
        RECT 845.400 615.600 847.200 621.600 ;
        RECT 14.100 603.000 15.900 611.400 ;
        RECT 34.200 607.050 36.000 611.400 ;
        RECT 34.200 605.400 39.600 607.050 ;
        RECT 11.700 601.350 15.900 603.000 ;
        RECT 38.700 602.100 39.600 605.400 ;
        RECT 56.100 603.000 57.900 611.400 ;
        RECT 71.400 606.300 73.200 611.400 ;
        RECT 77.400 606.300 79.200 611.400 ;
        RECT 71.400 604.950 79.200 606.300 ;
        RECT 80.400 605.400 82.200 611.400 ;
        RECT 80.400 603.300 81.600 605.400 ;
        RECT 97.200 604.200 99.000 611.400 ;
        RECT 113.400 608.400 115.200 611.400 ;
        RECT 103.950 604.950 106.050 607.050 ;
        RECT 113.400 605.100 114.600 608.400 ;
        RECT 56.100 601.350 60.300 603.000 ;
        RECT 77.850 602.250 81.600 603.300 ;
        RECT 95.400 603.300 99.000 604.200 ;
        RECT 77.850 602.100 79.050 602.250 ;
        RECT 11.700 596.100 12.600 601.350 ;
        RECT 14.100 599.100 15.900 599.850 ;
        RECT 20.100 599.100 21.900 599.850 ;
        RECT 29.100 599.100 30.900 599.850 ;
        RECT 31.950 598.950 34.200 601.050 ;
        RECT 35.100 599.100 36.900 599.850 ;
        RECT 37.950 598.950 43.050 601.050 ;
        RECT 50.100 599.100 51.900 599.850 ;
        RECT 56.100 599.100 57.900 599.850 ;
        RECT 13.950 595.950 16.050 598.050 ;
        RECT 19.950 595.950 22.050 598.050 ;
        RECT 28.950 595.950 31.050 598.050 ;
        RECT 32.100 597.150 33.900 597.900 ;
        RECT 34.950 595.950 37.050 598.050 ;
        RECT 10.950 592.950 13.050 595.050 ;
        RECT 16.950 592.950 19.050 595.050 ;
        RECT 11.700 586.800 12.600 591.900 ;
        RECT 17.100 591.150 18.900 591.900 ;
        RECT 38.700 591.600 39.600 597.900 ;
        RECT 49.950 595.950 52.050 598.050 ;
        RECT 55.950 595.950 58.050 598.050 ;
        RECT 59.400 596.100 60.300 601.350 ;
        RECT 70.950 598.950 73.050 601.050 ;
        RECT 74.100 599.100 75.900 599.850 ;
        RECT 76.950 598.950 79.200 601.050 ;
        RECT 80.100 599.100 81.900 599.850 ;
        RECT 95.400 599.100 96.600 603.300 ;
        RECT 104.550 601.050 105.450 604.950 ;
        RECT 133.200 604.200 135.000 611.400 ;
        RECT 112.950 601.950 115.050 604.050 ;
        RECT 131.400 603.300 135.000 604.200 ;
        RECT 150.000 604.200 151.800 611.400 ;
        RECT 150.000 603.300 153.600 604.200 ;
        RECT 103.950 598.950 106.050 601.050 ;
        RECT 109.950 598.950 112.050 601.050 ;
        RECT 71.100 597.150 72.900 597.900 ;
        RECT 73.950 595.950 76.050 598.050 ;
        RECT 52.950 592.950 55.050 595.050 ;
        RECT 58.950 592.950 64.050 595.050 ;
        RECT 77.100 594.900 78.150 597.900 ;
        RECT 79.950 595.950 82.050 598.050 ;
        RECT 92.100 596.100 93.900 596.850 ;
        RECT 94.950 595.950 97.200 598.050 ;
        RECT 98.100 596.100 99.900 596.850 ;
        RECT 29.400 590.700 37.200 591.600 ;
        RECT 11.700 585.900 18.300 586.800 ;
        RECT 11.700 585.600 12.600 585.900 ;
        RECT 10.800 579.600 12.600 585.600 ;
        RECT 16.800 585.600 18.300 585.900 ;
        RECT 16.800 579.600 18.600 585.600 ;
        RECT 29.400 579.600 31.200 590.700 ;
        RECT 35.400 579.600 37.200 590.700 ;
        RECT 38.400 579.600 40.200 591.600 ;
        RECT 53.100 591.150 54.900 591.900 ;
        RECT 59.400 586.800 60.300 591.900 ;
        RECT 76.950 591.600 78.150 594.900 ;
        RECT 91.950 592.950 94.050 595.050 ;
        RECT 53.700 585.900 60.300 586.800 ;
        RECT 53.700 585.600 55.200 585.900 ;
        RECT 53.400 579.600 55.200 585.600 ;
        RECT 59.400 585.600 60.300 585.900 ;
        RECT 59.400 579.600 61.200 585.600 ;
        RECT 76.500 579.600 78.300 591.600 ;
        RECT 95.400 585.600 96.600 594.900 ;
        RECT 97.950 592.950 100.050 595.050 ;
        RECT 104.550 589.050 105.450 598.950 ;
        RECT 113.700 597.900 114.900 600.900 ;
        RECT 115.950 598.950 118.050 601.050 ;
        RECT 131.400 599.100 132.600 603.300 ;
        RECT 152.400 599.100 153.600 603.300 ;
        RECT 170.100 603.000 171.900 611.400 ;
        RECT 190.200 607.050 192.000 611.400 ;
        RECT 213.000 607.050 214.800 611.400 ;
        RECT 190.200 605.400 195.600 607.050 ;
        RECT 167.700 601.350 171.900 603.000 ;
        RECT 194.700 602.100 195.600 605.400 ;
        RECT 209.400 605.400 214.800 607.050 ;
        RECT 227.400 606.300 229.200 611.400 ;
        RECT 233.400 606.300 235.200 611.400 ;
        RECT 209.400 602.100 210.300 605.400 ;
        RECT 227.400 604.950 235.200 606.300 ;
        RECT 236.400 605.400 238.200 611.400 ;
        RECT 251.400 608.400 253.200 611.400 ;
        RECT 236.400 603.300 237.600 605.400 ;
        RECT 241.950 604.950 244.050 607.050 ;
        RECT 233.850 602.250 237.600 603.300 ;
        RECT 233.850 602.100 235.050 602.250 ;
        RECT 110.100 597.150 111.900 597.900 ;
        RECT 113.700 592.650 115.050 597.900 ;
        RECT 116.100 597.150 117.900 597.900 ;
        RECT 128.100 596.100 129.900 596.850 ;
        RECT 130.950 595.950 133.050 598.050 ;
        RECT 134.100 596.100 135.900 596.850 ;
        RECT 149.100 596.100 150.900 596.850 ;
        RECT 151.950 595.950 154.050 598.050 ;
        RECT 155.100 596.100 156.900 596.850 ;
        RECT 167.700 596.100 168.600 601.350 ;
        RECT 170.100 599.100 171.900 599.850 ;
        RECT 176.100 599.100 177.900 599.850 ;
        RECT 185.100 599.100 186.900 599.850 ;
        RECT 187.950 598.950 190.050 601.050 ;
        RECT 191.100 599.100 192.900 599.850 ;
        RECT 193.950 598.950 199.050 601.050 ;
        RECT 208.950 600.450 211.050 601.050 ;
        RECT 203.550 599.550 211.050 600.450 ;
        RECT 169.800 595.950 172.050 598.050 ;
        RECT 175.950 595.950 178.050 598.050 ;
        RECT 184.950 595.950 187.050 598.050 ;
        RECT 188.100 597.150 189.900 597.900 ;
        RECT 190.950 595.950 193.050 598.050 ;
        RECT 127.950 592.950 130.050 595.050 ;
        RECT 113.700 591.600 116.400 592.650 ;
        RECT 103.950 586.950 106.050 589.050 ;
        RECT 95.400 579.600 97.200 585.600 ;
        RECT 114.600 579.600 116.400 591.600 ;
        RECT 131.400 585.600 132.600 594.900 ;
        RECT 133.950 592.950 136.200 595.050 ;
        RECT 148.950 592.950 151.050 595.050 ;
        RECT 152.400 585.600 153.600 594.900 ;
        RECT 154.950 592.950 157.050 595.050 ;
        RECT 166.950 594.450 169.050 595.050 ;
        RECT 161.550 593.550 169.050 594.450 ;
        RECT 161.550 586.050 162.450 593.550 ;
        RECT 166.950 592.950 169.050 593.550 ;
        RECT 172.950 592.950 175.050 595.050 ;
        RECT 167.700 586.800 168.600 591.900 ;
        RECT 173.100 591.150 174.900 591.900 ;
        RECT 194.700 591.600 195.600 597.900 ;
        RECT 185.400 590.700 193.200 591.600 ;
        RECT 131.400 579.600 133.200 585.600 ;
        RECT 151.800 579.600 153.600 585.600 ;
        RECT 160.950 583.950 163.050 586.050 ;
        RECT 167.700 585.900 174.300 586.800 ;
        RECT 167.700 585.600 168.600 585.900 ;
        RECT 166.800 579.600 168.600 585.600 ;
        RECT 172.800 585.600 174.300 585.900 ;
        RECT 172.800 579.600 174.600 585.600 ;
        RECT 185.400 579.600 187.200 590.700 ;
        RECT 191.400 579.600 193.200 590.700 ;
        RECT 194.400 579.600 196.200 591.600 ;
        RECT 203.550 589.050 204.450 599.550 ;
        RECT 208.950 598.950 211.050 599.550 ;
        RECT 212.100 599.100 213.900 599.850 ;
        RECT 214.950 598.950 217.050 601.050 ;
        RECT 218.100 599.100 219.900 599.850 ;
        RECT 226.800 598.950 229.050 601.050 ;
        RECT 230.100 599.100 231.900 599.850 ;
        RECT 232.800 598.950 235.050 601.050 ;
        RECT 236.100 599.100 237.900 599.850 ;
        RECT 209.400 591.600 210.300 597.900 ;
        RECT 211.950 595.950 214.050 598.050 ;
        RECT 215.100 597.150 216.900 597.900 ;
        RECT 217.950 595.950 220.050 598.050 ;
        RECT 227.100 597.150 228.900 597.900 ;
        RECT 229.950 595.950 232.050 598.050 ;
        RECT 233.100 594.900 234.150 597.900 ;
        RECT 235.950 595.950 238.200 598.050 ;
        RECT 242.550 595.050 243.450 604.950 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 248.100 600.150 249.900 600.900 ;
        RECT 251.400 599.100 252.600 608.400 ;
        RECT 268.200 604.200 270.000 611.400 ;
        RECT 285.300 607.200 287.100 611.400 ;
        RECT 266.400 603.300 270.000 604.200 ;
        RECT 285.150 605.400 287.100 607.200 ;
        RECT 266.400 599.100 267.600 603.300 ;
        RECT 285.150 602.100 286.050 605.400 ;
        RECT 287.100 603.900 288.900 604.500 ;
        RECT 292.800 603.900 294.600 611.400 ;
        RECT 287.100 602.700 294.600 603.900 ;
        RECT 305.400 605.400 307.200 611.400 ;
        RECT 283.950 598.950 286.050 601.050 ;
        RECT 287.100 599.100 288.900 599.850 ;
        RECT 247.950 595.950 253.050 598.050 ;
        RECT 263.100 596.100 264.900 596.850 ;
        RECT 265.950 595.950 268.050 598.050 ;
        RECT 269.100 596.100 270.900 596.850 ;
        RECT 232.950 591.600 234.150 594.900 ;
        RECT 241.950 592.950 244.050 595.050 ;
        RECT 202.950 586.950 205.050 589.050 ;
        RECT 208.800 579.600 210.600 591.600 ;
        RECT 211.800 590.700 219.600 591.600 ;
        RECT 211.800 579.600 213.600 590.700 ;
        RECT 217.800 579.600 219.600 590.700 ;
        RECT 232.500 579.600 234.300 591.600 ;
        RECT 251.400 585.600 252.600 594.900 ;
        RECT 262.800 592.950 265.050 595.050 ;
        RECT 266.400 585.600 267.600 594.900 ;
        RECT 268.950 592.950 271.050 595.050 ;
        RECT 283.950 591.600 285.000 597.900 ;
        RECT 286.950 595.950 289.050 598.050 ;
        RECT 251.400 579.600 253.200 585.600 ;
        RECT 266.400 579.600 268.200 585.600 ;
        RECT 283.200 579.600 285.000 591.600 ;
        RECT 290.550 585.600 291.600 602.700 ;
        RECT 305.400 602.100 306.600 605.400 ;
        RECT 310.950 604.950 313.050 607.050 ;
        RECT 327.000 605.400 328.800 611.400 ;
        RECT 337.950 607.950 340.050 610.050 ;
        RECT 292.950 598.950 295.050 601.050 ;
        RECT 304.950 600.450 307.050 601.050 ;
        RECT 311.550 600.450 312.450 604.950 ;
        RECT 327.000 602.100 328.050 605.400 ;
        RECT 302.100 599.100 303.900 599.850 ;
        RECT 304.950 599.550 312.450 600.450 ;
        RECT 304.950 598.950 307.050 599.550 ;
        RECT 319.950 598.950 322.050 601.050 ;
        RECT 323.250 599.100 324.900 599.850 ;
        RECT 325.950 598.950 328.050 601.050 ;
        RECT 329.100 599.100 330.750 599.850 ;
        RECT 331.950 598.950 334.050 601.050 ;
        RECT 338.550 600.450 339.450 607.950 ;
        RECT 343.500 605.400 345.300 611.400 ;
        RECT 349.800 608.400 351.600 611.400 ;
        RECT 359.400 608.400 361.200 611.400 ;
        RECT 343.800 602.100 345.000 605.400 ;
        RECT 349.800 604.500 351.000 608.400 ;
        RECT 345.900 603.600 351.000 604.500 ;
        RECT 360.000 604.500 361.200 608.400 ;
        RECT 365.700 605.400 367.500 611.400 ;
        RECT 360.000 603.600 365.100 604.500 ;
        RECT 345.900 602.700 347.850 603.600 ;
        RECT 346.950 602.100 347.850 602.700 ;
        RECT 343.950 600.450 346.050 601.050 ;
        RECT 338.550 599.550 346.050 600.450 ;
        RECT 343.950 598.950 346.050 599.550 ;
        RECT 293.100 597.150 294.900 597.900 ;
        RECT 301.950 595.950 304.050 598.050 ;
        RECT 289.800 579.600 291.600 585.600 ;
        RECT 305.400 591.600 306.600 597.900 ;
        RECT 320.100 597.150 321.900 597.900 ;
        RECT 322.950 595.950 325.050 598.050 ;
        RECT 326.100 594.900 326.850 597.900 ;
        RECT 328.950 595.950 331.050 598.050 ;
        RECT 347.100 597.900 347.850 602.100 ;
        RECT 363.150 602.700 365.100 603.600 ;
        RECT 363.150 602.100 364.050 602.700 ;
        RECT 366.000 602.100 367.200 605.400 ;
        RECT 373.950 604.950 376.050 607.050 ;
        RECT 379.500 605.400 381.300 611.400 ;
        RECT 385.800 608.400 387.600 611.400 ;
        RECT 349.950 598.950 352.050 601.050 ;
        RECT 358.950 598.950 361.050 601.050 ;
        RECT 363.150 597.900 363.900 602.100 ;
        RECT 364.950 600.450 367.050 601.050 ;
        RECT 364.950 599.550 372.450 600.450 ;
        RECT 364.950 598.950 367.050 599.550 ;
        RECT 332.100 597.150 333.750 597.900 ;
        RECT 325.950 593.400 326.850 594.900 ;
        RECT 322.800 592.500 326.850 593.400 ;
        RECT 305.400 579.600 307.200 591.600 ;
        RECT 319.800 580.500 321.600 591.600 ;
        RECT 322.800 581.400 324.600 592.500 ;
        RECT 343.800 591.600 345.000 597.900 ;
        RECT 346.950 594.300 347.850 597.900 ;
        RECT 350.100 597.150 351.900 597.900 ;
        RECT 359.100 597.150 360.900 597.900 ;
        RECT 345.900 593.400 347.850 594.300 ;
        RECT 363.150 594.300 364.050 597.900 ;
        RECT 363.150 593.400 365.100 594.300 ;
        RECT 345.900 592.500 351.600 593.400 ;
        RECT 325.800 590.400 333.600 591.300 ;
        RECT 325.800 580.500 327.600 590.400 ;
        RECT 319.800 579.600 327.600 580.500 ;
        RECT 331.800 579.600 333.600 590.400 ;
        RECT 343.500 579.600 345.300 591.600 ;
        RECT 350.400 585.600 351.600 592.500 ;
        RECT 349.800 579.600 351.600 585.600 ;
        RECT 359.400 592.500 365.100 593.400 ;
        RECT 359.400 585.600 360.600 592.500 ;
        RECT 366.000 591.600 367.200 597.900 ;
        RECT 371.550 592.050 372.450 599.550 ;
        RECT 374.550 595.050 375.450 604.950 ;
        RECT 379.800 602.100 381.000 605.400 ;
        RECT 385.800 604.500 387.000 608.400 ;
        RECT 381.900 603.600 387.000 604.500 ;
        RECT 399.000 604.200 400.800 611.400 ;
        RECT 415.800 605.400 417.600 611.400 ;
        RECT 421.800 608.400 423.600 611.400 ;
        RECT 381.900 602.700 383.850 603.600 ;
        RECT 399.000 603.300 402.600 604.200 ;
        RECT 382.950 602.100 383.850 602.700 ;
        RECT 376.950 598.950 382.050 601.050 ;
        RECT 383.100 597.900 383.850 602.100 ;
        RECT 385.950 598.950 388.050 601.050 ;
        RECT 401.400 599.100 402.600 603.300 ;
        RECT 415.950 599.100 417.000 605.400 ;
        RECT 421.800 604.200 422.700 608.400 ;
        RECT 436.800 605.400 438.600 611.400 ;
        RECT 442.800 608.400 444.600 611.400 ;
        RECT 419.250 603.300 422.700 604.200 ;
        RECT 419.250 602.400 421.050 603.300 ;
        RECT 373.950 592.950 376.050 595.050 ;
        RECT 359.400 579.600 361.200 585.600 ;
        RECT 365.700 579.600 367.500 591.600 ;
        RECT 370.950 589.950 373.050 592.050 ;
        RECT 379.800 591.600 381.000 597.900 ;
        RECT 382.950 594.300 383.850 597.900 ;
        RECT 386.100 597.150 387.900 597.900 ;
        RECT 398.100 596.100 399.900 596.850 ;
        RECT 400.950 595.950 403.050 598.050 ;
        RECT 404.100 596.100 405.900 596.850 ;
        RECT 415.950 595.950 418.050 598.050 ;
        RECT 381.900 593.400 383.850 594.300 ;
        RECT 381.900 592.500 387.600 593.400 ;
        RECT 397.800 592.950 400.050 595.050 ;
        RECT 379.500 579.600 381.300 591.600 ;
        RECT 386.400 585.600 387.600 592.500 ;
        RECT 401.400 585.600 402.600 594.900 ;
        RECT 403.950 592.950 406.050 595.050 ;
        RECT 416.700 591.600 418.050 594.900 ;
        RECT 419.400 594.600 420.300 602.400 ;
        RECT 424.950 601.950 427.050 604.050 ;
        RECT 421.950 598.950 424.050 601.050 ;
        RECT 425.100 600.150 426.900 600.900 ;
        RECT 436.950 599.100 438.000 605.400 ;
        RECT 442.800 604.200 443.700 608.400 ;
        RECT 462.000 607.050 463.800 611.400 ;
        RECT 440.250 603.300 443.700 604.200 ;
        RECT 458.400 605.400 463.800 607.050 ;
        RECT 440.250 602.400 442.050 603.300 ;
        RECT 422.100 597.150 423.900 597.900 ;
        RECT 436.950 595.950 439.050 598.050 ;
        RECT 419.400 594.000 421.200 594.600 ;
        RECT 419.400 592.800 426.600 594.000 ;
        RECT 419.400 592.650 420.300 592.800 ;
        RECT 425.400 591.600 426.600 592.800 ;
        RECT 416.700 590.100 419.100 591.600 ;
        RECT 385.800 579.600 387.600 585.600 ;
        RECT 400.800 579.600 402.600 585.600 ;
        RECT 417.300 579.600 419.100 590.100 ;
        RECT 424.800 579.600 426.600 591.600 ;
        RECT 437.700 591.600 439.050 594.900 ;
        RECT 440.400 594.600 441.300 602.400 ;
        RECT 445.950 601.950 448.050 604.050 ;
        RECT 458.400 602.100 459.300 605.400 ;
        RECT 482.100 603.000 483.900 611.400 ;
        RECT 499.800 608.400 501.600 611.400 ;
        RECT 479.700 601.350 483.900 603.000 ;
        RECT 442.950 598.950 445.050 601.050 ;
        RECT 446.100 600.150 447.900 600.900 ;
        RECT 457.950 598.950 460.050 601.050 ;
        RECT 461.100 599.100 462.900 599.850 ;
        RECT 463.950 598.950 466.050 601.050 ;
        RECT 467.100 599.100 468.900 599.850 ;
        RECT 443.100 597.150 444.900 597.900 ;
        RECT 440.400 594.000 442.200 594.600 ;
        RECT 440.400 592.800 447.600 594.000 ;
        RECT 440.400 592.650 441.300 592.800 ;
        RECT 446.400 591.600 447.600 592.800 ;
        RECT 458.400 591.600 459.300 597.900 ;
        RECT 460.800 595.950 463.050 598.050 ;
        RECT 464.100 597.150 465.900 597.900 ;
        RECT 466.950 595.950 469.200 598.050 ;
        RECT 479.700 596.100 480.600 601.350 ;
        RECT 482.100 599.100 483.900 599.850 ;
        RECT 488.100 599.100 489.900 599.850 ;
        RECT 500.400 599.100 501.600 608.400 ;
        RECT 502.950 601.950 505.050 604.050 ;
        RECT 518.100 603.000 519.900 611.400 ;
        RECT 538.200 607.050 540.000 611.400 ;
        RECT 538.200 605.400 543.600 607.050 ;
        RECT 515.700 601.350 519.900 603.000 ;
        RECT 542.700 602.100 543.600 605.400 ;
        RECT 554.400 606.300 556.200 611.400 ;
        RECT 560.400 606.300 562.200 611.400 ;
        RECT 554.400 604.950 562.200 606.300 ;
        RECT 563.400 605.400 565.200 611.400 ;
        RECT 578.400 608.400 580.200 611.400 ;
        RECT 563.400 603.300 564.600 605.400 ;
        RECT 578.400 605.100 579.600 608.400 ;
        RECT 593.400 606.300 595.200 611.400 ;
        RECT 599.400 606.300 601.200 611.400 ;
        RECT 593.400 604.950 601.200 606.300 ;
        RECT 602.400 605.400 604.200 611.400 ;
        RECT 560.850 602.250 564.600 603.300 ;
        RECT 560.850 602.100 562.050 602.250 ;
        RECT 577.950 601.950 580.050 604.050 ;
        RECT 602.400 603.300 603.600 605.400 ;
        RECT 617.400 604.500 619.200 611.400 ;
        RECT 623.400 604.500 625.200 611.400 ;
        RECT 629.400 604.500 631.200 611.400 ;
        RECT 635.400 604.500 637.200 611.400 ;
        RECT 643.950 607.950 646.050 610.050 ;
        RECT 617.400 603.300 621.300 604.500 ;
        RECT 623.400 603.300 627.300 604.500 ;
        RECT 629.400 603.300 633.300 604.500 ;
        RECT 635.400 603.300 638.100 604.500 ;
        RECT 599.850 602.250 603.600 603.300 ;
        RECT 620.100 602.400 621.300 603.300 ;
        RECT 626.100 602.400 627.300 603.300 ;
        RECT 632.100 602.400 633.300 603.300 ;
        RECT 599.850 602.100 601.050 602.250 ;
        RECT 503.100 600.150 504.900 600.900 ;
        RECT 481.950 595.950 484.050 598.050 ;
        RECT 487.950 595.950 490.050 598.050 ;
        RECT 499.950 595.950 505.050 598.050 ;
        RECT 515.700 596.100 516.600 601.350 ;
        RECT 620.100 601.200 624.300 602.400 ;
        RECT 518.100 599.100 519.900 599.850 ;
        RECT 524.100 599.100 525.900 599.850 ;
        RECT 533.100 599.100 534.900 599.850 ;
        RECT 535.950 598.950 538.050 601.050 ;
        RECT 539.100 599.100 540.900 599.850 ;
        RECT 541.950 598.950 547.050 601.050 ;
        RECT 550.950 598.950 556.050 601.050 ;
        RECT 557.100 599.100 558.900 599.850 ;
        RECT 559.950 598.950 562.050 601.050 ;
        RECT 563.100 599.100 564.900 599.850 ;
        RECT 574.950 598.950 577.050 601.050 ;
        RECT 517.950 595.950 520.050 598.050 ;
        RECT 523.950 595.950 526.200 598.050 ;
        RECT 532.950 595.950 535.050 598.050 ;
        RECT 536.100 597.150 537.900 597.900 ;
        RECT 538.950 595.950 541.050 598.050 ;
        RECT 478.950 592.950 481.050 595.050 ;
        RECT 484.800 592.950 487.050 595.050 ;
        RECT 437.700 590.100 440.100 591.600 ;
        RECT 438.300 579.600 440.100 590.100 ;
        RECT 445.800 579.600 447.600 591.600 ;
        RECT 457.800 579.600 459.600 591.600 ;
        RECT 460.800 590.700 468.600 591.600 ;
        RECT 460.800 579.600 462.600 590.700 ;
        RECT 466.800 579.600 468.600 590.700 ;
        RECT 479.700 586.800 480.600 591.900 ;
        RECT 485.100 591.150 486.900 591.900 ;
        RECT 479.700 585.900 486.300 586.800 ;
        RECT 479.700 585.600 480.600 585.900 ;
        RECT 478.800 579.600 480.600 585.600 ;
        RECT 484.800 585.600 486.300 585.900 ;
        RECT 500.400 585.600 501.600 594.900 ;
        RECT 511.950 592.950 517.050 595.050 ;
        RECT 520.950 592.950 523.050 595.050 ;
        RECT 515.700 586.800 516.600 591.900 ;
        RECT 521.100 591.150 522.900 591.900 ;
        RECT 542.700 591.600 543.600 597.900 ;
        RECT 554.100 597.150 555.900 597.900 ;
        RECT 556.950 595.950 559.050 598.050 ;
        RECT 560.100 594.900 561.150 597.900 ;
        RECT 562.950 595.950 565.050 598.050 ;
        RECT 578.700 597.900 579.900 600.900 ;
        RECT 580.950 598.950 583.050 601.050 ;
        RECT 589.950 598.950 595.050 601.050 ;
        RECT 596.100 599.100 597.900 599.850 ;
        RECT 598.950 598.950 601.200 601.050 ;
        RECT 602.100 599.100 603.900 599.850 ;
        RECT 617.100 599.100 618.900 599.850 ;
        RECT 575.100 597.150 576.900 597.900 ;
        RECT 559.950 591.600 561.150 594.900 ;
        RECT 578.700 592.650 580.050 597.900 ;
        RECT 581.100 597.150 582.900 597.900 ;
        RECT 593.100 597.150 594.900 597.900 ;
        RECT 595.950 595.950 598.050 598.050 ;
        RECT 599.100 594.900 600.150 597.900 ;
        RECT 601.950 595.950 604.050 598.050 ;
        RECT 578.700 591.600 581.400 592.650 ;
        RECT 598.950 591.600 600.150 594.900 ;
        RECT 533.400 590.700 541.200 591.600 ;
        RECT 515.700 585.900 522.300 586.800 ;
        RECT 515.700 585.600 516.600 585.900 ;
        RECT 484.800 579.600 486.600 585.600 ;
        RECT 499.800 579.600 501.600 585.600 ;
        RECT 514.800 579.600 516.600 585.600 ;
        RECT 520.800 585.600 522.300 585.900 ;
        RECT 520.800 579.600 522.600 585.600 ;
        RECT 533.400 579.600 535.200 590.700 ;
        RECT 539.400 579.600 541.200 590.700 ;
        RECT 542.400 579.600 544.200 591.600 ;
        RECT 559.500 579.600 561.300 591.600 ;
        RECT 579.600 579.600 581.400 591.600 ;
        RECT 598.500 579.600 600.300 591.600 ;
        RECT 602.550 589.050 603.450 595.950 ;
        RECT 620.100 593.700 621.300 601.200 ;
        RECT 622.500 600.600 624.300 601.200 ;
        RECT 626.100 601.200 630.300 602.400 ;
        RECT 626.100 593.700 627.300 601.200 ;
        RECT 628.500 600.600 630.300 601.200 ;
        RECT 632.100 601.200 636.300 602.400 ;
        RECT 632.100 593.700 633.300 601.200 ;
        RECT 634.500 600.600 636.300 601.200 ;
        RECT 637.200 599.100 638.100 603.300 ;
        RECT 637.950 597.450 640.050 598.050 ;
        RECT 644.550 597.450 645.450 607.950 ;
        RECT 654.000 604.200 655.800 611.400 ;
        RECT 670.800 605.400 672.600 611.400 ;
        RECT 654.000 603.300 657.600 604.200 ;
        RECT 656.400 599.100 657.600 603.300 ;
        RECT 671.400 603.300 672.600 605.400 ;
        RECT 673.800 606.300 675.600 611.400 ;
        RECT 679.800 606.300 681.600 611.400 ;
        RECT 673.800 604.950 681.600 606.300 ;
        RECT 694.200 604.200 696.000 611.400 ;
        RECT 709.800 605.400 711.600 611.400 ;
        RECT 692.400 603.300 696.000 604.200 ;
        RECT 710.400 603.300 711.600 605.400 ;
        RECT 712.800 606.300 714.600 611.400 ;
        RECT 718.800 606.300 720.600 611.400 ;
        RECT 712.800 604.950 720.600 606.300 ;
        RECT 728.400 606.300 730.200 611.400 ;
        RECT 734.400 606.300 736.200 611.400 ;
        RECT 728.400 604.950 736.200 606.300 ;
        RECT 737.400 605.400 739.200 611.400 ;
        RECT 737.400 603.300 738.600 605.400 ;
        RECT 754.200 604.200 756.000 611.400 ;
        RECT 760.950 604.950 763.050 607.050 ;
        RECT 767.400 606.300 769.200 611.400 ;
        RECT 773.400 606.300 775.200 611.400 ;
        RECT 767.400 604.950 775.200 606.300 ;
        RECT 776.400 605.400 778.200 611.400 ;
        RECT 781.950 607.950 784.050 610.050 ;
        RECT 671.400 602.250 675.150 603.300 ;
        RECT 673.950 602.100 675.150 602.250 ;
        RECT 671.100 599.100 672.900 599.850 ;
        RECT 673.950 598.950 676.050 601.050 ;
        RECT 677.100 599.100 678.900 599.850 ;
        RECT 679.950 598.950 682.050 601.050 ;
        RECT 692.400 599.100 693.600 603.300 ;
        RECT 710.400 602.250 714.150 603.300 ;
        RECT 712.950 602.100 714.150 602.250 ;
        RECT 734.850 602.250 738.600 603.300 ;
        RECT 752.400 603.300 756.000 604.200 ;
        RECT 734.850 602.100 736.050 602.250 ;
        RECT 710.100 599.100 711.900 599.850 ;
        RECT 712.950 598.950 715.050 601.050 ;
        RECT 716.100 599.100 717.900 599.850 ;
        RECT 718.950 598.950 721.050 601.050 ;
        RECT 727.800 598.950 730.050 601.050 ;
        RECT 731.100 599.100 732.900 599.850 ;
        RECT 733.950 598.950 736.050 601.050 ;
        RECT 737.100 599.100 738.900 599.850 ;
        RECT 752.400 599.100 753.600 603.300 ;
        RECT 761.550 600.450 762.450 604.950 ;
        RECT 776.400 603.300 777.600 605.400 ;
        RECT 773.850 602.250 777.600 603.300 ;
        RECT 773.850 602.100 775.050 602.250 ;
        RECT 766.950 600.450 769.050 601.050 ;
        RECT 761.550 599.550 769.050 600.450 ;
        RECT 766.950 598.950 769.050 599.550 ;
        RECT 770.100 599.100 771.900 599.850 ;
        RECT 772.950 598.950 775.200 601.050 ;
        RECT 776.100 599.100 777.900 599.850 ;
        RECT 637.950 596.550 645.450 597.450 ;
        RECT 637.950 595.950 640.050 596.550 ;
        RECT 653.100 596.100 654.900 596.850 ;
        RECT 655.950 595.950 658.050 598.050 ;
        RECT 659.100 596.100 660.900 596.850 ;
        RECT 670.950 595.950 673.050 598.050 ;
        RECT 637.200 593.700 638.100 594.900 ;
        RECT 617.400 592.500 621.300 593.700 ;
        RECT 623.400 592.500 627.300 593.700 ;
        RECT 629.400 592.500 633.300 593.700 ;
        RECT 635.400 592.500 638.100 593.700 ;
        RECT 652.950 592.950 655.050 595.050 ;
        RECT 601.950 586.950 604.050 589.050 ;
        RECT 617.400 579.600 619.200 592.500 ;
        RECT 623.400 579.600 625.200 592.500 ;
        RECT 629.400 579.600 631.200 592.500 ;
        RECT 635.400 579.600 637.200 592.500 ;
        RECT 653.550 591.000 654.450 592.950 ;
        RECT 652.950 586.950 655.050 591.000 ;
        RECT 656.400 585.600 657.600 594.900 ;
        RECT 658.950 592.950 661.050 595.050 ;
        RECT 674.850 594.900 675.900 597.900 ;
        RECT 676.950 595.950 679.050 598.050 ;
        RECT 680.100 597.150 681.900 597.900 ;
        RECT 689.100 596.100 690.900 596.850 ;
        RECT 691.950 595.950 694.050 598.050 ;
        RECT 695.100 596.100 696.900 596.850 ;
        RECT 709.950 595.950 712.050 598.050 ;
        RECT 674.850 591.600 676.050 594.900 ;
        RECT 688.800 592.950 691.050 595.050 ;
        RECT 655.800 579.600 657.600 585.600 ;
        RECT 674.700 579.600 676.500 591.600 ;
        RECT 692.400 585.600 693.600 594.900 ;
        RECT 694.950 592.950 697.050 595.050 ;
        RECT 713.850 594.900 714.900 597.900 ;
        RECT 715.950 595.950 718.050 598.050 ;
        RECT 719.100 597.150 720.900 597.900 ;
        RECT 728.100 597.150 729.900 597.900 ;
        RECT 730.950 595.950 733.050 598.050 ;
        RECT 734.100 594.900 735.150 597.900 ;
        RECT 736.950 595.950 739.050 598.050 ;
        RECT 749.100 596.100 750.900 596.850 ;
        RECT 751.950 595.950 754.050 598.050 ;
        RECT 767.100 597.150 768.900 597.900 ;
        RECT 755.100 596.100 756.900 596.850 ;
        RECT 769.950 595.950 772.050 598.050 ;
        RECT 706.950 589.950 709.050 592.050 ;
        RECT 713.850 591.600 715.050 594.900 ;
        RECT 733.950 591.600 735.150 594.900 ;
        RECT 748.950 592.950 751.050 595.050 ;
        RECT 707.550 586.050 708.450 589.950 ;
        RECT 692.400 579.600 694.200 585.600 ;
        RECT 706.800 583.950 708.900 586.050 ;
        RECT 713.700 579.600 715.500 591.600 ;
        RECT 733.500 579.600 735.300 591.600 ;
        RECT 752.400 585.600 753.600 594.900 ;
        RECT 754.950 592.950 757.200 595.050 ;
        RECT 773.100 594.900 774.150 597.900 ;
        RECT 775.950 595.950 778.050 598.050 ;
        RECT 755.550 591.000 756.450 592.950 ;
        RECT 772.950 591.600 774.150 594.900 ;
        RECT 754.950 586.950 757.050 591.000 ;
        RECT 752.400 579.600 754.200 585.600 ;
        RECT 772.500 579.600 774.300 591.600 ;
        RECT 782.550 583.050 783.450 607.950 ;
        RECT 793.200 604.200 795.000 611.400 ;
        RECT 808.800 608.400 810.600 611.400 ;
        RECT 791.400 603.300 795.000 604.200 ;
        RECT 791.400 599.100 792.600 603.300 ;
        RECT 809.400 599.100 810.600 608.400 ;
        RECT 824.400 605.400 826.200 611.400 ;
        RECT 839.400 608.400 841.200 611.400 ;
        RECT 812.100 600.150 813.900 600.900 ;
        RECT 821.100 599.100 822.900 599.850 ;
        RECT 824.700 599.100 826.050 605.400 ;
        RECT 840.000 604.500 841.200 608.400 ;
        RECT 845.700 605.400 847.500 611.400 ;
        RECT 850.950 607.950 853.050 610.050 ;
        RECT 840.000 603.600 845.100 604.500 ;
        RECT 843.150 602.700 845.100 603.600 ;
        RECT 843.150 602.100 844.050 602.700 ;
        RECT 846.000 602.100 847.200 605.400 ;
        RECT 788.100 596.100 789.900 596.850 ;
        RECT 790.950 595.950 793.050 598.050 ;
        RECT 794.100 596.100 795.900 596.850 ;
        RECT 808.800 595.950 811.050 598.050 ;
        RECT 787.950 592.950 790.050 595.050 ;
        RECT 791.400 585.600 792.600 594.900 ;
        RECT 793.950 592.950 796.050 595.050 ;
        RECT 824.700 594.900 825.900 599.100 ;
        RECT 838.950 598.950 841.050 601.050 ;
        RECT 826.950 597.450 829.050 598.050 ;
        RECT 843.150 597.900 843.900 602.100 ;
        RECT 844.950 598.950 847.050 601.050 ;
        RECT 851.550 598.050 852.450 607.950 ;
        RECT 826.950 596.550 834.450 597.450 ;
        RECT 839.100 597.150 840.900 597.900 ;
        RECT 826.950 595.950 829.050 596.550 ;
        RECT 809.400 585.600 810.600 594.900 ;
        RECT 824.700 591.600 826.050 594.900 ;
        RECT 781.950 580.950 784.050 583.050 ;
        RECT 791.400 579.600 793.200 585.600 ;
        RECT 808.800 579.600 810.600 585.600 ;
        RECT 824.400 579.600 826.200 591.600 ;
        RECT 833.550 583.050 834.450 596.550 ;
        RECT 843.150 594.300 844.050 597.900 ;
        RECT 843.150 593.400 845.100 594.300 ;
        RECT 839.400 592.500 845.100 593.400 ;
        RECT 839.400 585.600 840.600 592.500 ;
        RECT 846.000 591.600 847.200 597.900 ;
        RECT 850.950 595.950 853.050 598.050 ;
        RECT 832.950 580.950 835.050 583.050 ;
        RECT 839.400 579.600 841.200 585.600 ;
        RECT 845.700 579.600 847.500 591.600 ;
        RECT 10.500 563.400 12.300 575.400 ;
        RECT 16.800 569.400 18.600 575.400 ;
        RECT 10.800 557.100 12.000 563.400 ;
        RECT 17.400 562.500 18.600 569.400 ;
        RECT 32.700 563.400 34.500 575.400 ;
        RECT 12.900 561.600 18.600 562.500 ;
        RECT 12.900 560.700 14.850 561.600 ;
        RECT 13.950 557.100 14.850 560.700 ;
        RECT 32.850 560.100 34.050 563.400 ;
        RECT 43.950 562.950 46.050 565.050 ;
        RECT 53.700 563.400 55.500 575.400 ;
        RECT 68.400 565.500 70.200 575.400 ;
        RECT 74.400 574.500 82.200 575.400 ;
        RECT 74.400 565.500 76.200 574.500 ;
        RECT 68.400 564.600 76.200 565.500 ;
        RECT 77.400 565.800 79.200 573.600 ;
        RECT 80.400 566.700 82.200 574.500 ;
        RECT 84.000 574.500 91.800 575.400 ;
        RECT 84.000 565.800 85.800 574.500 ;
        RECT 77.400 564.900 85.800 565.800 ;
        RECT 87.000 565.800 88.800 573.600 ;
        RECT 87.000 563.400 88.200 565.800 ;
        RECT 90.000 565.200 91.800 574.500 ;
        RECT 103.800 563.400 105.600 575.400 ;
        RECT 106.800 564.300 108.600 575.400 ;
        RECT 112.800 564.300 114.600 575.400 ;
        RECT 124.800 569.400 126.600 575.400 ;
        RECT 106.800 563.400 114.600 564.300 ;
        RECT 125.700 569.100 126.600 569.400 ;
        RECT 130.800 569.400 132.600 575.400 ;
        RECT 145.800 574.500 153.600 575.400 ;
        RECT 130.800 569.100 132.300 569.400 ;
        RECT 125.700 568.200 132.300 569.100 ;
        RECT 17.100 557.100 18.900 557.850 ;
        RECT 14.100 552.900 14.850 557.100 ;
        RECT 28.950 556.950 31.050 559.050 ;
        RECT 32.850 557.100 33.900 560.100 ;
        RECT 34.950 556.950 37.050 559.050 ;
        RECT 38.100 557.100 39.900 557.850 ;
        RECT 44.550 556.050 45.450 562.950 ;
        RECT 53.850 560.100 55.050 563.400 ;
        RECT 84.750 562.200 88.200 563.400 ;
        RECT 49.800 556.950 52.050 559.050 ;
        RECT 53.850 557.100 54.900 560.100 ;
        RECT 84.750 559.950 85.950 562.200 ;
        RECT 55.950 556.950 58.050 559.050 ;
        RECT 59.100 557.100 60.900 557.850 ;
        RECT 71.100 556.950 72.900 557.700 ;
        RECT 76.950 556.800 79.050 559.050 ;
        RECT 80.100 556.950 81.900 557.700 ;
        RECT 16.950 553.950 19.050 556.050 ;
        RECT 29.100 555.150 30.900 555.900 ;
        RECT 31.950 553.950 34.050 556.050 ;
        RECT 35.100 555.150 36.900 555.900 ;
        RECT 37.950 553.950 40.050 556.050 ;
        RECT 43.800 553.950 45.900 556.050 ;
        RECT 50.100 555.150 51.900 555.900 ;
        RECT 52.950 553.950 55.050 556.050 ;
        RECT 56.100 555.150 57.900 555.900 ;
        RECT 58.950 553.950 61.200 556.050 ;
        RECT 70.950 553.800 73.050 555.900 ;
        RECT 77.100 555.000 78.900 555.750 ;
        RECT 10.800 549.600 12.000 552.900 ;
        RECT 13.950 552.300 14.850 552.900 ;
        RECT 31.950 552.750 33.150 552.900 ;
        RECT 52.950 552.750 54.150 552.900 ;
        RECT 12.900 551.400 14.850 552.300 ;
        RECT 29.400 551.700 33.150 552.750 ;
        RECT 50.400 551.700 54.150 552.750 ;
        RECT 12.900 550.500 18.000 551.400 ;
        RECT 10.500 543.600 12.300 549.600 ;
        RECT 16.800 546.600 18.000 550.500 ;
        RECT 29.400 549.600 30.600 551.700 ;
        RECT 16.800 543.600 18.600 546.600 ;
        RECT 28.800 543.600 30.600 549.600 ;
        RECT 31.800 548.700 39.600 550.050 ;
        RECT 50.400 549.600 51.600 551.700 ;
        RECT 79.950 550.950 82.050 555.900 ;
        RECT 84.750 555.750 84.900 559.950 ;
        RECT 88.050 558.900 91.050 559.050 ;
        RECT 85.950 556.950 91.050 558.900 ;
        RECT 104.400 557.100 105.300 563.400 ;
        RECT 125.700 563.100 126.600 568.200 ;
        RECT 131.100 563.100 132.900 563.850 ;
        RECT 145.800 563.400 147.600 574.500 ;
        RECT 148.800 562.500 150.600 573.600 ;
        RECT 151.800 564.600 153.600 574.500 ;
        RECT 157.800 564.600 159.600 575.400 ;
        RECT 151.800 563.700 159.600 564.600 ;
        RECT 169.200 563.400 171.000 575.400 ;
        RECT 175.800 569.400 177.600 575.400 ;
        RECT 190.800 569.400 192.600 575.400 ;
        RECT 124.950 561.450 127.050 562.050 ;
        RECT 119.550 560.550 127.050 561.450 ;
        RECT 106.950 556.950 109.050 559.050 ;
        RECT 110.100 557.100 111.900 557.850 ;
        RECT 112.950 556.950 115.050 559.050 ;
        RECT 85.950 556.800 88.050 556.950 ;
        RECT 31.800 543.600 33.600 548.700 ;
        RECT 37.800 543.600 39.600 548.700 ;
        RECT 49.800 543.600 51.600 549.600 ;
        RECT 52.800 548.700 60.600 550.050 ;
        RECT 52.800 543.600 54.600 548.700 ;
        RECT 58.800 543.600 60.600 548.700 ;
        RECT 84.750 548.400 85.950 555.750 ;
        RECT 100.950 553.950 106.050 556.050 ;
        RECT 107.100 555.150 108.900 555.900 ;
        RECT 109.950 553.950 112.050 556.050 ;
        RECT 113.100 555.150 114.900 555.900 ;
        RECT 75.150 547.500 85.950 548.400 ;
        RECT 104.400 549.600 105.300 552.900 ;
        RECT 104.400 547.950 109.800 549.600 ;
        RECT 75.150 546.600 76.200 547.500 ;
        RECT 81.150 546.600 82.200 547.500 ;
        RECT 74.400 543.600 76.200 546.600 ;
        RECT 80.400 543.600 82.200 546.600 ;
        RECT 108.000 543.600 109.800 547.950 ;
        RECT 119.550 547.050 120.450 560.550 ;
        RECT 124.950 559.950 127.050 560.550 ;
        RECT 130.950 559.950 133.050 562.050 ;
        RECT 148.800 561.600 152.850 562.500 ;
        RECT 151.950 560.100 152.850 561.600 ;
        RECT 125.700 553.650 126.600 558.900 ;
        RECT 127.950 556.950 130.050 559.050 ;
        RECT 133.950 556.950 136.200 559.050 ;
        RECT 146.100 557.100 147.900 557.850 ;
        RECT 148.950 556.950 151.200 559.050 ;
        RECT 152.100 557.100 152.850 560.100 ;
        RECT 154.950 556.950 157.200 559.050 ;
        RECT 158.100 557.100 159.750 557.850 ;
        RECT 169.950 557.100 171.000 563.400 ;
        RECT 172.950 556.950 175.050 559.050 ;
        RECT 128.100 555.150 129.900 555.900 ;
        RECT 134.100 555.150 135.900 555.900 ;
        RECT 145.950 553.950 148.050 556.050 ;
        RECT 149.250 555.150 150.900 555.900 ;
        RECT 151.950 553.950 154.200 556.050 ;
        RECT 155.100 555.150 156.750 555.900 ;
        RECT 157.950 553.950 160.050 556.050 ;
        RECT 169.950 555.450 172.050 556.050 ;
        RECT 164.550 554.550 172.050 555.450 ;
        RECT 173.100 555.150 174.900 555.900 ;
        RECT 125.700 552.000 129.900 553.650 ;
        RECT 118.950 544.950 121.050 547.050 ;
        RECT 128.100 543.600 129.900 552.000 ;
        RECT 153.000 549.600 154.050 552.900 ;
        RECT 164.550 550.050 165.450 554.550 ;
        RECT 169.950 553.950 172.050 554.550 ;
        RECT 153.000 543.600 154.800 549.600 ;
        RECT 163.950 547.950 166.050 550.050 ;
        RECT 171.150 549.600 172.050 552.900 ;
        RECT 176.550 552.300 177.600 569.400 ;
        RECT 191.700 569.100 192.600 569.400 ;
        RECT 196.800 569.400 198.600 575.400 ;
        RECT 211.800 569.400 213.600 575.400 ;
        RECT 196.800 569.100 198.300 569.400 ;
        RECT 191.700 568.200 198.300 569.100 ;
        RECT 191.700 563.100 192.600 568.200 ;
        RECT 197.100 563.100 198.900 563.850 ;
        RECT 187.950 559.950 193.050 562.050 ;
        RECT 196.950 559.950 199.050 562.050 ;
        RECT 212.400 560.100 213.600 569.400 ;
        RECT 230.700 563.400 232.500 575.400 ;
        RECT 251.700 563.400 253.500 575.400 ;
        RECT 270.300 564.900 272.100 575.400 ;
        RECT 269.700 563.400 272.100 564.900 ;
        RECT 277.800 563.400 279.600 575.400 ;
        RECT 291.600 563.400 293.400 575.400 ;
        RECT 298.800 571.950 300.900 574.050 ;
        RECT 230.850 560.100 232.050 563.400 ;
        RECT 251.850 560.100 253.050 563.400 ;
        RECT 269.700 560.100 271.050 563.400 ;
        RECT 272.400 562.200 273.300 562.350 ;
        RECT 278.400 562.200 279.600 563.400 ;
        RECT 272.400 561.000 279.600 562.200 ;
        RECT 290.700 562.350 293.400 563.400 ;
        RECT 272.400 560.400 274.200 561.000 ;
        RECT 179.100 557.100 180.900 557.850 ;
        RECT 178.950 553.950 181.050 556.050 ;
        RECT 191.700 553.650 192.600 558.900 ;
        RECT 193.950 556.950 196.050 559.050 ;
        RECT 199.950 556.950 202.050 559.050 ;
        RECT 208.950 556.950 214.050 559.050 ;
        RECT 226.950 556.950 229.050 559.050 ;
        RECT 230.850 557.100 231.900 560.100 ;
        RECT 232.950 556.950 235.050 559.050 ;
        RECT 236.100 557.100 237.900 557.850 ;
        RECT 247.950 556.950 250.050 559.050 ;
        RECT 251.850 557.100 252.900 560.100 ;
        RECT 253.950 556.950 256.050 559.050 ;
        RECT 268.950 558.450 271.050 559.050 ;
        RECT 257.100 557.100 258.900 557.850 ;
        RECT 263.550 557.550 271.050 558.450 ;
        RECT 194.100 555.150 195.900 555.900 ;
        RECT 200.100 555.150 201.900 555.900 ;
        RECT 173.100 551.100 180.600 552.300 ;
        RECT 191.700 552.000 195.900 553.650 ;
        RECT 173.100 550.500 174.900 551.100 ;
        RECT 171.150 547.800 173.100 549.600 ;
        RECT 171.300 543.600 173.100 547.800 ;
        RECT 178.800 543.600 180.600 551.100 ;
        RECT 194.100 543.600 195.900 552.000 ;
        RECT 212.400 546.600 213.600 555.900 ;
        RECT 227.100 555.150 228.900 555.900 ;
        RECT 215.100 554.100 216.900 554.850 ;
        RECT 229.950 553.950 232.050 556.050 ;
        RECT 233.100 555.150 234.900 555.900 ;
        RECT 235.950 553.950 238.050 556.050 ;
        RECT 248.100 555.150 249.900 555.900 ;
        RECT 250.950 553.950 253.200 556.050 ;
        RECT 254.100 555.150 255.900 555.900 ;
        RECT 256.950 553.950 259.050 556.050 ;
        RECT 214.950 550.950 217.050 553.050 ;
        RECT 229.950 552.750 231.150 552.900 ;
        RECT 250.950 552.750 252.150 552.900 ;
        RECT 227.400 551.700 231.150 552.750 ;
        RECT 248.400 551.700 252.150 552.750 ;
        RECT 227.400 549.600 228.600 551.700 ;
        RECT 211.800 543.600 213.600 546.600 ;
        RECT 226.800 543.600 228.600 549.600 ;
        RECT 229.800 548.700 237.600 550.050 ;
        RECT 248.400 549.600 249.600 551.700 ;
        RECT 263.550 550.050 264.450 557.550 ;
        RECT 268.950 556.950 271.050 557.550 ;
        RECT 229.800 543.600 231.600 548.700 ;
        RECT 235.800 543.600 237.600 548.700 ;
        RECT 247.800 543.600 249.600 549.600 ;
        RECT 250.800 548.700 258.600 550.050 ;
        RECT 250.800 543.600 252.600 548.700 ;
        RECT 256.800 543.600 258.600 548.700 ;
        RECT 262.950 547.950 265.050 550.050 ;
        RECT 268.950 549.600 270.000 555.900 ;
        RECT 272.400 552.600 273.300 560.400 ;
        RECT 275.100 557.100 276.900 557.850 ;
        RECT 287.100 557.100 288.900 557.850 ;
        RECT 290.700 557.100 292.050 562.350 ;
        RECT 293.100 557.100 294.900 557.850 ;
        RECT 274.950 553.950 277.050 556.050 ;
        RECT 278.100 554.100 279.900 554.850 ;
        RECT 286.950 553.950 289.050 556.050 ;
        RECT 290.700 554.100 291.900 557.100 ;
        RECT 292.950 553.950 295.050 556.050 ;
        RECT 272.250 551.700 274.050 552.600 ;
        RECT 272.250 550.800 275.700 551.700 ;
        RECT 277.950 550.950 280.050 553.050 ;
        RECT 289.950 550.950 292.050 553.050 ;
        RECT 268.800 543.600 270.600 549.600 ;
        RECT 274.800 546.600 275.700 550.800 ;
        RECT 299.550 550.050 300.450 571.950 ;
        RECT 308.400 569.400 310.200 575.400 ;
        RECT 326.400 569.400 328.200 575.400 ;
        RECT 304.950 559.950 307.050 562.050 ;
        RECT 308.400 560.100 309.600 569.400 ;
        RECT 310.800 567.000 312.900 568.050 ;
        RECT 310.800 565.950 313.050 567.000 ;
        RECT 316.950 565.950 319.050 568.050 ;
        RECT 310.950 564.000 313.050 565.950 ;
        RECT 311.550 562.050 312.450 564.000 ;
        RECT 310.950 559.950 313.200 562.050 ;
        RECT 305.100 558.150 306.900 558.900 ;
        RECT 307.950 556.950 310.050 559.050 ;
        RECT 311.100 558.150 312.900 558.900 ;
        RECT 308.400 551.700 309.600 555.900 ;
        RECT 317.550 553.050 318.450 565.950 ;
        RECT 323.100 557.100 324.900 557.850 ;
        RECT 322.950 553.950 325.050 556.050 ;
        RECT 308.400 550.800 312.000 551.700 ;
        RECT 316.950 550.950 319.050 553.050 ;
        RECT 326.400 552.300 327.450 569.400 ;
        RECT 333.000 563.400 334.800 575.400 ;
        RECT 337.950 571.950 340.050 574.050 ;
        RECT 328.950 556.950 331.050 559.050 ;
        RECT 333.000 557.100 334.050 563.400 ;
        RECT 329.100 555.150 330.900 555.900 ;
        RECT 331.950 555.450 334.050 556.050 ;
        RECT 338.550 555.450 339.450 571.950 ;
        RECT 348.600 563.400 350.400 575.400 ;
        RECT 365.400 569.400 367.200 575.400 ;
        RECT 383.400 569.400 385.200 575.400 ;
        RECT 400.800 569.400 402.600 575.400 ;
        RECT 348.600 562.350 351.300 563.400 ;
        RECT 347.100 557.100 348.900 557.850 ;
        RECT 349.950 557.100 351.300 562.350 ;
        RECT 361.950 559.950 364.050 562.050 ;
        RECT 365.400 560.100 366.600 569.400 ;
        RECT 367.950 559.950 370.050 562.050 ;
        RECT 383.400 560.100 384.600 569.400 ;
        RECT 397.950 559.950 400.050 562.050 ;
        RECT 401.400 560.100 402.600 569.400 ;
        RECT 415.800 563.400 417.600 575.400 ;
        RECT 418.800 564.300 420.600 575.400 ;
        RECT 424.800 564.300 426.600 575.400 ;
        RECT 439.800 569.400 441.600 575.400 ;
        RECT 418.800 563.400 426.600 564.300 ;
        RECT 403.950 559.950 406.050 562.050 ;
        RECT 362.100 558.150 363.900 558.900 ;
        RECT 353.100 557.100 354.900 557.850 ;
        RECT 331.950 554.550 339.450 555.450 ;
        RECT 331.950 553.950 334.050 554.550 ;
        RECT 346.950 553.950 349.050 556.050 ;
        RECT 350.100 554.100 351.300 557.100 ;
        RECT 364.950 556.950 367.050 559.050 ;
        RECT 368.100 558.150 369.900 558.900 ;
        RECT 379.950 556.950 385.050 559.050 ;
        RECT 398.100 558.150 399.900 558.900 ;
        RECT 400.950 556.950 403.050 559.050 ;
        RECT 404.100 558.150 405.900 558.900 ;
        RECT 416.400 557.100 417.300 563.400 ;
        RECT 436.950 559.950 439.050 562.050 ;
        RECT 440.400 560.100 441.600 569.400 ;
        RECT 448.950 568.950 451.050 571.050 ;
        RECT 442.950 564.000 445.050 568.050 ;
        RECT 443.550 562.050 444.450 564.000 ;
        RECT 449.550 562.050 450.450 568.950 ;
        RECT 452.400 564.600 454.200 575.400 ;
        RECT 458.400 574.500 466.200 575.400 ;
        RECT 458.400 564.600 460.200 574.500 ;
        RECT 452.400 563.700 460.200 564.600 ;
        RECT 461.400 562.500 463.200 573.600 ;
        RECT 464.400 563.400 466.200 574.500 ;
        RECT 480.600 563.400 482.400 575.400 ;
        RECT 499.500 563.400 501.300 575.400 ;
        RECT 519.600 563.400 521.400 575.400 ;
        RECT 536.400 569.400 538.200 575.400 ;
        RECT 536.700 569.100 538.200 569.400 ;
        RECT 542.400 569.400 544.200 575.400 ;
        RECT 557.400 569.400 559.200 575.400 ;
        RECT 542.400 569.100 543.300 569.400 ;
        RECT 536.700 568.200 543.300 569.100 ;
        RECT 557.700 569.100 559.200 569.400 ;
        RECT 563.400 569.400 565.200 575.400 ;
        RECT 578.400 569.400 580.200 575.400 ;
        RECT 563.400 569.100 564.300 569.400 ;
        RECT 557.700 568.200 564.300 569.100 ;
        RECT 578.700 569.100 580.200 569.400 ;
        RECT 584.400 569.400 586.200 575.400 ;
        RECT 599.400 569.400 601.200 575.400 ;
        RECT 584.400 569.100 585.300 569.400 ;
        RECT 578.700 568.200 585.300 569.100 ;
        RECT 442.950 559.950 445.050 562.050 ;
        RECT 448.950 559.950 451.050 562.050 ;
        RECT 459.150 561.600 463.200 562.500 ;
        RECT 479.700 562.350 482.400 563.400 ;
        RECT 459.150 560.100 460.050 561.600 ;
        RECT 418.950 556.950 421.050 559.050 ;
        RECT 422.100 557.100 423.900 557.850 ;
        RECT 424.950 556.950 427.200 559.050 ;
        RECT 437.100 558.150 438.900 558.900 ;
        RECT 439.950 556.950 442.050 559.050 ;
        RECT 443.100 558.150 444.900 558.900 ;
        RECT 452.250 557.100 453.900 557.850 ;
        RECT 454.800 556.950 457.050 559.050 ;
        RECT 459.150 557.100 459.900 560.100 ;
        RECT 460.950 556.950 463.200 559.050 ;
        RECT 464.100 557.100 465.900 557.850 ;
        RECT 469.950 556.950 472.050 559.050 ;
        RECT 476.100 557.100 477.900 557.850 ;
        RECT 479.700 557.100 481.050 562.350 ;
        RECT 499.950 560.100 501.150 563.400 ;
        RECT 519.600 562.350 522.300 563.400 ;
        RECT 536.100 563.100 537.900 563.850 ;
        RECT 542.400 563.100 543.300 568.200 ;
        RECT 557.100 563.100 558.900 563.850 ;
        RECT 563.400 563.100 564.300 568.200 ;
        RECT 578.100 563.100 579.900 563.850 ;
        RECT 584.400 563.100 585.300 568.200 ;
        RECT 482.100 557.100 483.900 557.850 ;
        RECT 494.100 557.100 495.900 557.850 ;
        RECT 352.950 553.950 355.050 556.050 ;
        RECT 323.400 551.100 330.900 552.300 ;
        RECT 290.400 546.600 291.600 549.900 ;
        RECT 298.950 547.950 301.050 550.050 ;
        RECT 274.800 543.600 276.600 546.600 ;
        RECT 290.400 543.600 292.200 546.600 ;
        RECT 310.200 543.600 312.000 550.800 ;
        RECT 323.400 543.600 325.200 551.100 ;
        RECT 329.100 550.500 330.900 551.100 ;
        RECT 331.950 549.600 332.850 552.900 ;
        RECT 349.950 550.950 352.050 553.050 ;
        RECT 365.400 551.700 366.600 555.900 ;
        RECT 380.100 554.100 381.900 554.850 ;
        RECT 365.400 550.800 369.000 551.700 ;
        RECT 379.950 550.950 382.050 553.050 ;
        RECT 330.900 547.800 332.850 549.600 ;
        RECT 330.900 543.600 332.700 547.800 ;
        RECT 350.400 546.600 351.600 549.900 ;
        RECT 349.800 543.600 351.600 546.600 ;
        RECT 367.200 543.600 369.000 550.800 ;
        RECT 383.400 546.600 384.600 555.900 ;
        RECT 401.400 551.700 402.600 555.900 ;
        RECT 415.950 553.950 418.050 556.050 ;
        RECT 419.100 555.150 420.900 555.900 ;
        RECT 421.950 553.950 424.050 556.050 ;
        RECT 425.100 555.150 426.900 555.900 ;
        RECT 399.000 550.800 402.600 551.700 ;
        RECT 383.400 543.600 385.200 546.600 ;
        RECT 399.000 543.600 400.800 550.800 ;
        RECT 416.400 549.600 417.300 552.900 ;
        RECT 440.400 551.700 441.600 555.900 ;
        RECT 451.950 553.950 454.050 556.050 ;
        RECT 455.250 555.150 456.900 555.900 ;
        RECT 457.800 553.950 460.050 556.050 ;
        RECT 461.100 555.150 462.750 555.900 ;
        RECT 463.950 553.950 466.200 556.050 ;
        RECT 438.000 550.800 441.600 551.700 ;
        RECT 416.400 547.950 421.800 549.600 ;
        RECT 420.000 543.600 421.800 547.950 ;
        RECT 438.000 543.600 439.800 550.800 ;
        RECT 457.950 549.600 459.000 552.900 ;
        RECT 457.200 543.600 459.000 549.600 ;
        RECT 470.550 547.050 471.450 556.950 ;
        RECT 475.800 553.950 478.050 556.050 ;
        RECT 479.700 554.100 480.900 557.100 ;
        RECT 496.950 556.950 499.050 559.050 ;
        RECT 500.100 557.100 501.150 560.100 ;
        RECT 502.950 556.950 505.050 559.050 ;
        RECT 518.100 557.100 519.900 557.850 ;
        RECT 520.950 557.100 522.300 562.350 ;
        RECT 535.950 559.950 538.050 562.050 ;
        RECT 541.950 559.950 547.050 562.050 ;
        RECT 556.950 559.950 559.050 562.050 ;
        RECT 562.950 561.450 565.050 562.050 ;
        RECT 562.950 560.550 570.450 561.450 ;
        RECT 562.950 559.950 565.050 560.550 ;
        RECT 524.100 557.100 525.900 557.850 ;
        RECT 481.950 553.950 484.050 556.050 ;
        RECT 493.950 553.950 496.050 556.050 ;
        RECT 497.100 555.150 498.900 555.900 ;
        RECT 499.950 553.950 502.050 556.050 ;
        RECT 503.100 555.150 504.900 555.900 ;
        RECT 517.950 553.950 520.050 556.050 ;
        RECT 521.100 554.100 522.300 557.100 ;
        RECT 532.950 556.950 535.050 559.050 ;
        RECT 538.950 556.950 541.050 559.050 ;
        RECT 523.950 553.950 526.050 556.050 ;
        RECT 533.100 555.150 534.900 555.900 ;
        RECT 539.100 555.150 540.900 555.900 ;
        RECT 542.400 553.650 543.300 558.900 ;
        RECT 553.950 556.950 556.050 559.050 ;
        RECT 559.950 556.950 562.050 559.050 ;
        RECT 554.100 555.150 555.900 555.900 ;
        RECT 560.100 555.150 561.900 555.900 ;
        RECT 563.400 553.650 564.300 558.900 ;
        RECT 569.550 556.050 570.450 560.550 ;
        RECT 577.950 559.950 580.050 562.050 ;
        RECT 583.950 559.950 589.050 562.050 ;
        RECT 574.800 556.950 577.050 559.050 ;
        RECT 580.950 556.950 583.200 559.050 ;
        RECT 568.950 553.950 571.050 556.050 ;
        RECT 575.100 555.150 576.900 555.900 ;
        RECT 581.100 555.150 582.900 555.900 ;
        RECT 584.400 553.650 585.300 558.900 ;
        RECT 596.100 557.100 597.900 557.850 ;
        RECT 595.950 553.950 598.050 556.050 ;
        RECT 478.950 550.950 481.050 553.050 ;
        RECT 500.850 552.750 502.050 552.900 ;
        RECT 500.850 551.700 504.600 552.750 ;
        RECT 469.950 544.950 472.050 547.050 ;
        RECT 479.400 546.600 480.600 549.900 ;
        RECT 494.400 548.700 502.200 550.050 ;
        RECT 479.400 543.600 481.200 546.600 ;
        RECT 494.400 543.600 496.200 548.700 ;
        RECT 500.400 543.600 502.200 548.700 ;
        RECT 503.400 549.600 504.600 551.700 ;
        RECT 520.950 550.950 523.050 553.050 ;
        RECT 539.100 552.000 543.300 553.650 ;
        RECT 560.100 552.000 564.300 553.650 ;
        RECT 581.100 552.000 585.300 553.650 ;
        RECT 599.400 552.300 600.450 569.400 ;
        RECT 606.000 563.400 607.800 575.400 ;
        RECT 622.500 563.400 624.300 575.400 ;
        RECT 632.550 563.400 634.350 575.400 ;
        RECT 640.050 569.400 641.850 575.400 ;
        RECT 637.950 567.300 641.850 569.400 ;
        RECT 647.850 568.500 649.650 575.400 ;
        RECT 655.650 569.400 657.450 575.400 ;
        RECT 656.250 568.500 657.450 569.400 ;
        RECT 646.950 567.450 653.550 568.500 ;
        RECT 646.950 566.700 648.750 567.450 ;
        RECT 651.750 566.700 653.550 567.450 ;
        RECT 656.250 566.400 661.050 568.500 ;
        RECT 639.150 564.600 641.850 566.400 ;
        RECT 642.750 565.800 644.550 566.400 ;
        RECT 642.750 564.900 649.050 565.800 ;
        RECT 656.250 565.500 657.450 566.400 ;
        RECT 642.750 564.600 644.550 564.900 ;
        RECT 640.950 563.700 641.850 564.600 ;
        RECT 601.950 556.950 604.050 559.050 ;
        RECT 606.000 557.100 607.050 563.400 ;
        RECT 622.950 560.100 624.150 563.400 ;
        RECT 617.100 557.100 618.900 557.850 ;
        RECT 619.950 556.950 622.050 559.050 ;
        RECT 623.100 557.100 624.150 560.100 ;
        RECT 625.950 556.950 628.050 559.050 ;
        RECT 632.550 556.050 633.750 563.400 ;
        RECT 637.950 562.800 640.050 563.700 ;
        RECT 640.950 562.800 646.950 563.700 ;
        RECT 635.850 561.600 640.050 562.800 ;
        RECT 634.950 559.800 636.750 561.600 ;
        RECT 646.050 557.100 646.950 562.800 ;
        RECT 648.150 562.800 649.050 564.900 ;
        RECT 649.950 564.300 657.450 565.500 ;
        RECT 649.950 563.700 651.750 564.300 ;
        RECT 664.050 563.400 665.850 575.400 ;
        RECT 654.750 562.800 665.850 563.400 ;
        RECT 648.150 562.200 665.850 562.800 ;
        RECT 648.150 561.900 656.550 562.200 ;
        RECT 654.750 561.600 656.550 561.900 ;
        RECT 659.100 556.800 660.900 557.100 ;
        RECT 602.100 555.150 603.900 555.900 ;
        RECT 604.950 553.950 607.050 556.050 ;
        RECT 616.950 553.950 619.050 556.050 ;
        RECT 620.100 555.150 621.900 555.900 ;
        RECT 622.950 553.950 625.050 556.050 ;
        RECT 626.100 555.150 627.900 555.900 ;
        RECT 632.550 553.950 633.900 556.050 ;
        RECT 634.950 553.950 637.050 556.050 ;
        RECT 638.100 553.950 638.850 555.750 ;
        RECT 646.950 553.950 649.050 556.050 ;
        RECT 652.950 553.950 655.050 556.050 ;
        RECT 656.100 555.900 660.900 556.800 ;
        RECT 659.100 555.300 660.900 555.900 ;
        RECT 662.100 555.150 663.900 556.950 ;
        RECT 656.100 554.400 657.900 555.000 ;
        RECT 662.100 554.400 663.000 555.150 ;
        RECT 503.400 543.600 505.200 549.600 ;
        RECT 521.400 546.600 522.600 549.900 ;
        RECT 520.800 543.600 522.600 546.600 ;
        RECT 539.100 543.600 540.900 552.000 ;
        RECT 560.100 543.600 561.900 552.000 ;
        RECT 581.100 543.600 582.900 552.000 ;
        RECT 596.400 551.100 603.900 552.300 ;
        RECT 596.400 543.600 598.200 551.100 ;
        RECT 602.100 550.500 603.900 551.100 ;
        RECT 604.950 549.600 605.850 552.900 ;
        RECT 623.850 552.750 625.050 552.900 ;
        RECT 623.850 551.700 627.600 552.750 ;
        RECT 603.900 547.800 605.850 549.600 ;
        RECT 617.400 548.700 625.200 550.050 ;
        RECT 603.900 543.600 605.700 547.800 ;
        RECT 617.400 543.600 619.200 548.700 ;
        RECT 623.400 543.600 625.200 548.700 ;
        RECT 626.400 549.600 627.600 551.700 ;
        RECT 632.550 549.600 633.750 553.950 ;
        RECT 656.100 553.200 663.000 554.400 ;
        RECT 646.050 552.000 646.950 552.900 ;
        RECT 656.100 552.000 657.150 553.200 ;
        RECT 646.050 551.100 657.150 552.000 ;
        RECT 646.050 550.800 646.950 551.100 ;
        RECT 626.400 543.600 628.200 549.600 ;
        RECT 632.550 543.600 634.350 549.600 ;
        RECT 637.950 548.700 640.050 549.600 ;
        RECT 645.150 549.000 646.950 550.800 ;
        RECT 656.100 550.200 657.150 551.100 ;
        RECT 652.350 549.450 654.150 550.200 ;
        RECT 637.950 547.500 641.700 548.700 ;
        RECT 640.650 546.600 641.700 547.500 ;
        RECT 649.200 548.400 654.150 549.450 ;
        RECT 655.650 548.400 657.450 550.200 ;
        RECT 664.950 549.600 665.850 562.200 ;
        RECT 649.200 546.600 650.250 548.400 ;
        RECT 658.950 547.500 661.050 549.600 ;
        RECT 658.950 546.600 660.000 547.500 ;
        RECT 640.650 543.600 642.450 546.600 ;
        RECT 648.450 543.600 650.250 546.600 ;
        RECT 656.250 545.700 660.000 546.600 ;
        RECT 656.250 543.600 658.050 545.700 ;
        RECT 664.050 543.600 665.850 549.600 ;
        RECT 668.550 563.400 670.350 575.400 ;
        RECT 676.050 569.400 677.850 575.400 ;
        RECT 673.950 567.300 677.850 569.400 ;
        RECT 683.850 568.500 685.650 575.400 ;
        RECT 691.650 569.400 693.450 575.400 ;
        RECT 692.250 568.500 693.450 569.400 ;
        RECT 682.950 567.450 689.550 568.500 ;
        RECT 682.950 566.700 684.750 567.450 ;
        RECT 687.750 566.700 689.550 567.450 ;
        RECT 692.250 566.400 697.050 568.500 ;
        RECT 675.150 564.600 677.850 566.400 ;
        RECT 678.750 565.800 680.550 566.400 ;
        RECT 678.750 564.900 685.050 565.800 ;
        RECT 692.250 565.500 693.450 566.400 ;
        RECT 678.750 564.600 680.550 564.900 ;
        RECT 676.950 563.700 677.850 564.600 ;
        RECT 668.550 556.050 669.750 563.400 ;
        RECT 673.950 562.800 676.050 563.700 ;
        RECT 676.950 562.800 682.950 563.700 ;
        RECT 671.850 561.600 676.050 562.800 ;
        RECT 670.950 559.800 672.750 561.600 ;
        RECT 682.050 557.100 682.950 562.800 ;
        RECT 684.150 562.800 685.050 564.900 ;
        RECT 685.950 564.300 693.450 565.500 ;
        RECT 685.950 563.700 687.750 564.300 ;
        RECT 700.050 563.400 701.850 575.400 ;
        RECT 690.750 562.800 701.850 563.400 ;
        RECT 684.150 562.200 701.850 562.800 ;
        RECT 684.150 561.900 692.550 562.200 ;
        RECT 690.750 561.600 692.550 561.900 ;
        RECT 668.550 553.950 669.900 556.050 ;
        RECT 670.950 553.950 673.050 556.050 ;
        RECT 674.100 553.950 674.850 555.750 ;
        RECT 682.950 553.950 685.050 556.050 ;
        RECT 688.950 553.950 691.050 559.050 ;
        RECT 695.100 556.800 696.900 557.100 ;
        RECT 692.100 555.900 696.900 556.800 ;
        RECT 695.100 555.300 696.900 555.900 ;
        RECT 698.100 555.150 699.900 556.950 ;
        RECT 692.100 554.400 693.900 555.000 ;
        RECT 698.100 554.400 699.000 555.150 ;
        RECT 668.550 549.600 669.750 553.950 ;
        RECT 692.100 553.200 699.000 554.400 ;
        RECT 682.050 552.000 682.950 552.900 ;
        RECT 692.100 552.000 693.150 553.200 ;
        RECT 682.050 551.100 693.150 552.000 ;
        RECT 682.050 550.800 682.950 551.100 ;
        RECT 668.550 543.600 670.350 549.600 ;
        RECT 673.950 548.700 676.050 549.600 ;
        RECT 681.150 549.000 682.950 550.800 ;
        RECT 692.100 550.200 693.150 551.100 ;
        RECT 688.350 549.450 690.150 550.200 ;
        RECT 673.950 547.500 677.700 548.700 ;
        RECT 676.650 546.600 677.700 547.500 ;
        RECT 685.200 548.400 690.150 549.450 ;
        RECT 691.650 548.400 693.450 550.200 ;
        RECT 700.950 549.600 701.850 562.200 ;
        RECT 685.200 546.600 686.250 548.400 ;
        RECT 694.950 547.500 697.050 549.600 ;
        RECT 694.950 546.600 696.000 547.500 ;
        RECT 676.650 543.600 678.450 546.600 ;
        RECT 684.450 543.600 686.250 546.600 ;
        RECT 692.250 545.700 696.000 546.600 ;
        RECT 692.250 543.600 694.050 545.700 ;
        RECT 700.050 543.600 701.850 549.600 ;
        RECT 704.550 563.400 706.350 575.400 ;
        RECT 712.050 569.400 713.850 575.400 ;
        RECT 709.950 567.300 713.850 569.400 ;
        RECT 719.850 568.500 721.650 575.400 ;
        RECT 727.650 569.400 729.450 575.400 ;
        RECT 728.250 568.500 729.450 569.400 ;
        RECT 718.950 567.450 725.550 568.500 ;
        RECT 718.950 566.700 720.750 567.450 ;
        RECT 723.750 566.700 725.550 567.450 ;
        RECT 728.250 566.400 733.050 568.500 ;
        RECT 711.150 564.600 713.850 566.400 ;
        RECT 714.750 565.800 716.550 566.400 ;
        RECT 714.750 564.900 721.050 565.800 ;
        RECT 728.250 565.500 729.450 566.400 ;
        RECT 714.750 564.600 716.550 564.900 ;
        RECT 712.950 563.700 713.850 564.600 ;
        RECT 704.550 556.050 705.750 563.400 ;
        RECT 709.950 562.800 712.050 563.700 ;
        RECT 712.950 562.800 718.950 563.700 ;
        RECT 707.850 561.600 712.050 562.800 ;
        RECT 706.950 559.800 708.750 561.600 ;
        RECT 718.050 557.100 718.950 562.800 ;
        RECT 720.150 562.800 721.050 564.900 ;
        RECT 721.950 564.300 729.450 565.500 ;
        RECT 721.950 563.700 723.750 564.300 ;
        RECT 736.050 563.400 737.850 575.400 ;
        RECT 751.500 563.400 753.300 575.400 ;
        RECT 770.400 569.400 772.200 575.400 ;
        RECT 788.400 569.400 790.200 575.400 ;
        RECT 726.750 562.800 737.850 563.400 ;
        RECT 720.150 562.200 737.850 562.800 ;
        RECT 720.150 561.900 728.550 562.200 ;
        RECT 726.750 561.600 728.550 561.900 ;
        RECT 731.100 556.800 732.900 557.100 ;
        RECT 704.550 553.950 705.900 556.050 ;
        RECT 706.950 553.950 709.050 556.050 ;
        RECT 710.100 553.950 710.850 555.750 ;
        RECT 718.800 553.950 721.050 556.050 ;
        RECT 724.950 553.950 727.050 556.050 ;
        RECT 728.100 555.900 732.900 556.800 ;
        RECT 731.100 555.300 732.900 555.900 ;
        RECT 734.100 555.150 735.900 556.950 ;
        RECT 728.100 554.400 729.900 555.000 ;
        RECT 734.100 554.400 735.000 555.150 ;
        RECT 704.550 549.600 705.750 553.950 ;
        RECT 728.100 553.200 735.000 554.400 ;
        RECT 718.050 552.000 718.950 552.900 ;
        RECT 728.100 552.000 729.150 553.200 ;
        RECT 718.050 551.100 729.150 552.000 ;
        RECT 718.050 550.800 718.950 551.100 ;
        RECT 704.550 543.600 706.350 549.600 ;
        RECT 709.950 548.700 712.050 549.600 ;
        RECT 717.150 549.000 718.950 550.800 ;
        RECT 728.100 550.200 729.150 551.100 ;
        RECT 724.350 549.450 726.150 550.200 ;
        RECT 709.950 547.500 713.700 548.700 ;
        RECT 712.650 546.600 713.700 547.500 ;
        RECT 721.200 548.400 726.150 549.450 ;
        RECT 727.650 548.400 729.450 550.200 ;
        RECT 736.950 549.600 737.850 562.200 ;
        RECT 751.950 560.100 753.150 563.400 ;
        RECT 746.100 557.100 747.900 557.850 ;
        RECT 748.950 556.950 751.050 559.050 ;
        RECT 752.100 557.100 753.150 560.100 ;
        RECT 766.950 559.950 769.050 562.050 ;
        RECT 770.400 560.100 771.600 569.400 ;
        RECT 772.950 559.950 775.050 562.050 ;
        RECT 788.400 560.100 789.600 569.400 ;
        RECT 794.550 563.400 796.350 575.400 ;
        RECT 802.050 569.400 803.850 575.400 ;
        RECT 799.950 567.300 803.850 569.400 ;
        RECT 809.850 568.500 811.650 575.400 ;
        RECT 817.650 569.400 819.450 575.400 ;
        RECT 818.250 568.500 819.450 569.400 ;
        RECT 808.950 567.450 815.550 568.500 ;
        RECT 808.950 566.700 810.750 567.450 ;
        RECT 813.750 566.700 815.550 567.450 ;
        RECT 818.250 566.400 823.050 568.500 ;
        RECT 801.150 564.600 803.850 566.400 ;
        RECT 804.750 565.800 806.550 566.400 ;
        RECT 804.750 564.900 811.050 565.800 ;
        RECT 818.250 565.500 819.450 566.400 ;
        RECT 804.750 564.600 806.550 564.900 ;
        RECT 802.950 563.700 803.850 564.600 ;
        RECT 754.950 556.950 757.050 559.050 ;
        RECT 767.100 558.150 768.900 558.900 ;
        RECT 769.950 556.950 772.050 559.050 ;
        RECT 773.100 558.150 774.900 558.900 ;
        RECT 787.950 556.950 790.050 559.050 ;
        RECT 794.550 556.050 795.750 563.400 ;
        RECT 799.950 562.800 802.050 563.700 ;
        RECT 802.950 562.800 808.950 563.700 ;
        RECT 797.850 561.600 802.050 562.800 ;
        RECT 796.950 559.800 798.750 561.600 ;
        RECT 808.050 557.100 808.950 562.800 ;
        RECT 810.150 562.800 811.050 564.900 ;
        RECT 811.950 564.300 819.450 565.500 ;
        RECT 811.950 563.700 813.750 564.300 ;
        RECT 826.050 563.400 827.850 575.400 ;
        RECT 816.750 562.800 827.850 563.400 ;
        RECT 810.150 562.200 827.850 562.800 ;
        RECT 810.150 561.900 818.550 562.200 ;
        RECT 816.750 561.600 818.550 561.900 ;
        RECT 821.100 556.800 822.900 557.100 ;
        RECT 745.800 553.950 748.050 556.050 ;
        RECT 749.100 555.150 750.900 555.900 ;
        RECT 751.950 553.950 754.050 556.050 ;
        RECT 755.100 555.150 756.900 555.900 ;
        RECT 752.850 552.750 754.050 552.900 ;
        RECT 752.850 551.700 756.600 552.750 ;
        RECT 721.200 546.600 722.250 548.400 ;
        RECT 730.950 547.500 733.050 549.600 ;
        RECT 730.950 546.600 732.000 547.500 ;
        RECT 712.650 543.600 714.450 546.600 ;
        RECT 720.450 543.600 722.250 546.600 ;
        RECT 728.250 545.700 732.000 546.600 ;
        RECT 728.250 543.600 730.050 545.700 ;
        RECT 736.050 543.600 737.850 549.600 ;
        RECT 746.400 548.700 754.200 550.050 ;
        RECT 746.400 543.600 748.200 548.700 ;
        RECT 752.400 543.600 754.200 548.700 ;
        RECT 755.400 549.600 756.600 551.700 ;
        RECT 770.400 551.700 771.600 555.900 ;
        RECT 785.100 554.100 786.900 554.850 ;
        RECT 770.400 550.800 774.000 551.700 ;
        RECT 784.950 550.950 787.050 553.050 ;
        RECT 755.400 543.600 757.200 549.600 ;
        RECT 772.200 543.600 774.000 550.800 ;
        RECT 788.400 546.600 789.600 555.900 ;
        RECT 794.550 553.950 795.900 556.050 ;
        RECT 796.950 553.950 799.050 556.050 ;
        RECT 800.100 553.950 800.850 555.750 ;
        RECT 808.800 553.950 811.050 556.050 ;
        RECT 814.950 553.950 817.050 556.050 ;
        RECT 818.100 555.900 822.900 556.800 ;
        RECT 821.100 555.300 822.900 555.900 ;
        RECT 824.100 555.150 825.900 556.950 ;
        RECT 818.100 554.400 819.900 555.000 ;
        RECT 824.100 554.400 825.000 555.150 ;
        RECT 794.550 549.600 795.750 553.950 ;
        RECT 818.100 553.200 825.000 554.400 ;
        RECT 808.050 552.000 808.950 552.900 ;
        RECT 818.100 552.000 819.150 553.200 ;
        RECT 808.050 551.100 819.150 552.000 ;
        RECT 808.050 550.800 808.950 551.100 ;
        RECT 788.400 543.600 790.200 546.600 ;
        RECT 794.550 543.600 796.350 549.600 ;
        RECT 799.950 548.700 802.050 549.600 ;
        RECT 807.150 549.000 808.950 550.800 ;
        RECT 818.100 550.200 819.150 551.100 ;
        RECT 814.350 549.450 816.150 550.200 ;
        RECT 799.950 547.500 803.700 548.700 ;
        RECT 802.650 546.600 803.700 547.500 ;
        RECT 811.200 548.400 816.150 549.450 ;
        RECT 817.650 548.400 819.450 550.200 ;
        RECT 826.950 549.600 827.850 562.200 ;
        RECT 839.400 569.400 841.200 575.400 ;
        RECT 839.400 560.100 840.600 569.400 ;
        RECT 838.950 556.950 844.050 559.050 ;
        RECT 836.100 554.100 837.900 554.850 ;
        RECT 835.950 550.950 838.050 553.050 ;
        RECT 811.200 546.600 812.250 548.400 ;
        RECT 820.950 547.500 823.050 549.600 ;
        RECT 820.950 546.600 822.000 547.500 ;
        RECT 802.650 543.600 804.450 546.600 ;
        RECT 810.450 543.600 812.250 546.600 ;
        RECT 818.250 545.700 822.000 546.600 ;
        RECT 818.250 543.600 820.050 545.700 ;
        RECT 826.050 543.600 827.850 549.600 ;
        RECT 839.400 546.600 840.600 555.900 ;
        RECT 839.400 543.600 841.200 546.600 ;
        RECT 15.000 535.050 16.800 539.400 ;
        RECT 11.400 533.400 16.800 535.050 ;
        RECT 11.400 530.100 12.300 533.400 ;
        RECT 35.100 531.000 36.900 539.400 ;
        RECT 56.100 531.000 57.900 539.400 ;
        RECT 76.200 535.050 78.000 539.400 ;
        RECT 64.950 532.950 67.050 535.050 ;
        RECT 76.200 533.400 81.600 535.050 ;
        RECT 35.100 529.350 39.300 531.000 ;
        RECT 56.100 529.350 60.300 531.000 ;
        RECT 10.800 526.950 13.050 529.050 ;
        RECT 14.100 527.100 15.900 527.850 ;
        RECT 16.800 526.950 19.050 529.050 ;
        RECT 20.100 527.100 21.900 527.850 ;
        RECT 29.100 527.100 30.900 527.850 ;
        RECT 35.100 527.100 36.900 527.850 ;
        RECT 11.400 519.600 12.300 525.900 ;
        RECT 13.950 523.950 16.050 526.050 ;
        RECT 17.100 525.150 18.900 525.900 ;
        RECT 19.950 523.950 22.200 526.050 ;
        RECT 28.950 523.950 31.050 526.050 ;
        RECT 34.950 523.950 37.050 526.050 ;
        RECT 38.400 524.100 39.300 529.350 ;
        RECT 50.100 527.100 51.900 527.850 ;
        RECT 56.100 527.100 57.900 527.850 ;
        RECT 49.950 523.950 52.050 526.050 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 59.400 524.100 60.300 529.350 ;
        RECT 31.950 520.950 34.200 523.050 ;
        RECT 37.950 520.950 43.050 523.050 ;
        RECT 52.800 520.950 55.050 523.050 ;
        RECT 58.950 522.450 61.050 523.050 ;
        RECT 65.550 522.450 66.450 532.950 ;
        RECT 80.700 530.100 81.600 533.400 ;
        RECT 92.400 534.300 94.200 539.400 ;
        RECT 98.400 534.300 100.200 539.400 ;
        RECT 92.400 532.950 100.200 534.300 ;
        RECT 101.400 533.400 103.200 539.400 ;
        RECT 101.400 531.300 102.600 533.400 ;
        RECT 98.850 530.250 102.600 531.300 ;
        RECT 119.100 531.000 120.900 539.400 ;
        RECT 139.200 535.050 141.000 539.400 ;
        RECT 157.800 536.400 159.600 539.400 ;
        RECT 139.200 533.400 144.600 535.050 ;
        RECT 98.850 530.100 100.050 530.250 ;
        RECT 119.100 529.350 123.300 531.000 ;
        RECT 143.700 530.100 144.600 533.400 ;
        RECT 71.100 527.100 72.900 527.850 ;
        RECT 73.950 526.950 76.050 529.050 ;
        RECT 77.100 527.100 78.900 527.850 ;
        RECT 79.950 526.950 85.050 529.050 ;
        RECT 91.950 526.950 94.050 529.050 ;
        RECT 95.100 527.100 96.900 527.850 ;
        RECT 97.950 526.950 100.200 529.050 ;
        RECT 101.100 527.100 102.900 527.850 ;
        RECT 113.100 527.100 114.900 527.850 ;
        RECT 119.100 527.100 120.900 527.850 ;
        RECT 70.950 523.950 73.050 526.050 ;
        RECT 74.100 525.150 75.900 525.900 ;
        RECT 76.950 523.950 79.050 526.050 ;
        RECT 58.950 521.550 66.450 522.450 ;
        RECT 58.950 520.950 61.050 521.550 ;
        RECT 10.800 507.600 12.600 519.600 ;
        RECT 13.800 518.700 21.600 519.600 ;
        RECT 32.100 519.150 33.900 519.900 ;
        RECT 13.800 507.600 15.600 518.700 ;
        RECT 19.800 507.600 21.600 518.700 ;
        RECT 38.400 514.800 39.300 519.900 ;
        RECT 53.100 519.150 54.900 519.900 ;
        RECT 59.400 514.800 60.300 519.900 ;
        RECT 80.700 519.600 81.600 525.900 ;
        RECT 92.100 525.150 93.900 525.900 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 98.100 522.900 99.150 525.900 ;
        RECT 100.950 523.950 103.050 526.050 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 118.950 523.950 121.050 526.050 ;
        RECT 122.400 524.100 123.300 529.350 ;
        RECT 134.100 527.100 135.900 527.850 ;
        RECT 136.950 526.950 139.050 529.050 ;
        RECT 142.950 528.450 145.050 529.050 ;
        RECT 140.100 527.100 141.900 527.850 ;
        RECT 142.950 527.550 150.450 528.450 ;
        RECT 142.950 526.950 145.050 527.550 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 137.100 525.150 138.900 525.900 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 97.950 519.600 99.150 522.900 ;
        RECT 115.950 520.950 118.050 523.050 ;
        RECT 121.950 520.950 127.050 523.050 ;
        RECT 32.700 513.900 39.300 514.800 ;
        RECT 32.700 513.600 34.200 513.900 ;
        RECT 32.400 507.600 34.200 513.600 ;
        RECT 38.400 513.600 39.300 513.900 ;
        RECT 53.700 513.900 60.300 514.800 ;
        RECT 53.700 513.600 55.200 513.900 ;
        RECT 38.400 507.600 40.200 513.600 ;
        RECT 53.400 507.600 55.200 513.600 ;
        RECT 59.400 513.600 60.300 513.900 ;
        RECT 71.400 518.700 79.200 519.600 ;
        RECT 59.400 507.600 61.200 513.600 ;
        RECT 71.400 507.600 73.200 518.700 ;
        RECT 77.400 507.600 79.200 518.700 ;
        RECT 80.400 507.600 82.200 519.600 ;
        RECT 97.500 507.600 99.300 519.600 ;
        RECT 116.100 519.150 117.900 519.900 ;
        RECT 122.400 514.800 123.300 519.900 ;
        RECT 143.700 519.600 144.600 525.900 ;
        RECT 116.700 513.900 123.300 514.800 ;
        RECT 116.700 513.600 118.200 513.900 ;
        RECT 116.400 507.600 118.200 513.600 ;
        RECT 122.400 513.600 123.300 513.900 ;
        RECT 134.400 518.700 142.200 519.600 ;
        RECT 122.400 507.600 124.200 513.600 ;
        RECT 134.400 507.600 136.200 518.700 ;
        RECT 140.400 507.600 142.200 518.700 ;
        RECT 143.400 507.600 145.200 519.600 ;
        RECT 149.550 517.050 150.450 527.550 ;
        RECT 158.400 527.100 159.600 536.400 ;
        RECT 175.200 533.400 177.000 539.400 ;
        RECT 160.950 529.950 163.050 532.050 ;
        RECT 175.950 530.100 177.000 533.400 ;
        RECT 200.100 531.000 201.900 539.400 ;
        RECT 219.000 532.200 220.800 539.400 ;
        RECT 237.300 535.200 239.100 539.400 ;
        RECT 237.150 533.400 239.100 535.200 ;
        RECT 219.000 531.300 222.600 532.200 ;
        RECT 200.100 529.350 204.300 531.000 ;
        RECT 161.100 528.150 162.900 528.900 ;
        RECT 169.950 526.950 172.050 529.050 ;
        RECT 173.250 527.100 174.900 527.850 ;
        RECT 175.950 526.950 178.050 529.050 ;
        RECT 179.100 527.100 180.750 527.850 ;
        RECT 181.950 526.950 184.050 529.050 ;
        RECT 194.100 527.100 195.900 527.850 ;
        RECT 200.100 527.100 201.900 527.850 ;
        RECT 154.950 523.950 160.050 526.050 ;
        RECT 170.250 525.150 171.900 525.900 ;
        RECT 172.950 523.950 175.050 526.050 ;
        RECT 177.150 522.900 177.900 525.900 ;
        RECT 178.950 523.950 181.050 526.050 ;
        RECT 182.100 525.150 183.900 525.900 ;
        RECT 193.950 523.950 196.050 526.050 ;
        RECT 199.950 523.950 202.050 526.050 ;
        RECT 203.400 524.100 204.300 529.350 ;
        RECT 221.400 527.100 222.600 531.300 ;
        RECT 237.150 530.100 238.050 533.400 ;
        RECT 239.100 531.900 240.900 532.500 ;
        RECT 244.800 531.900 246.600 539.400 ;
        RECT 259.200 533.400 261.000 539.400 ;
        RECT 239.100 530.700 246.600 531.900 ;
        RECT 232.800 526.950 238.050 529.050 ;
        RECT 239.100 527.100 240.900 527.850 ;
        RECT 218.100 524.100 219.900 524.850 ;
        RECT 220.950 523.950 223.050 526.050 ;
        RECT 224.100 524.100 225.900 524.850 ;
        RECT 148.950 514.950 151.050 517.050 ;
        RECT 158.400 513.600 159.600 522.900 ;
        RECT 177.150 521.400 178.050 522.900 ;
        RECT 177.150 520.500 181.200 521.400 ;
        RECT 196.950 520.950 199.050 523.050 ;
        RECT 202.950 520.950 208.050 523.050 ;
        RECT 217.950 520.950 220.200 523.050 ;
        RECT 157.800 507.600 159.600 513.600 ;
        RECT 170.400 518.400 178.200 519.300 ;
        RECT 170.400 507.600 172.200 518.400 ;
        RECT 176.400 508.500 178.200 518.400 ;
        RECT 179.400 509.400 181.200 520.500 ;
        RECT 182.400 508.500 184.200 519.600 ;
        RECT 197.100 519.150 198.900 519.900 ;
        RECT 203.400 514.800 204.300 519.900 ;
        RECT 197.700 513.900 204.300 514.800 ;
        RECT 197.700 513.600 199.200 513.900 ;
        RECT 176.400 507.600 184.200 508.500 ;
        RECT 197.400 507.600 199.200 513.600 ;
        RECT 203.400 513.600 204.300 513.900 ;
        RECT 221.400 513.600 222.600 522.900 ;
        RECT 223.950 520.950 226.050 523.050 ;
        RECT 229.950 520.950 232.050 523.050 ;
        RECT 230.550 517.050 231.450 520.950 ;
        RECT 235.950 519.600 237.000 525.900 ;
        RECT 238.950 520.950 241.050 526.050 ;
        RECT 230.100 514.950 232.200 517.050 ;
        RECT 203.400 507.600 205.200 513.600 ;
        RECT 220.800 507.600 222.600 513.600 ;
        RECT 235.200 507.600 237.000 519.600 ;
        RECT 242.550 513.600 243.600 530.700 ;
        RECT 259.950 530.100 261.000 533.400 ;
        RECT 282.000 532.200 283.800 539.400 ;
        RECT 299.400 536.400 301.200 539.400 ;
        RECT 299.400 533.100 300.600 536.400 ;
        RECT 316.800 533.400 318.600 539.400 ;
        RECT 282.000 531.300 285.600 532.200 ;
        RECT 244.950 526.950 247.050 529.050 ;
        RECT 253.950 526.950 256.050 529.050 ;
        RECT 257.250 527.100 258.900 527.850 ;
        RECT 259.950 526.950 262.050 529.050 ;
        RECT 263.100 527.100 264.750 527.850 ;
        RECT 265.950 526.950 271.050 529.050 ;
        RECT 284.400 527.100 285.600 531.300 ;
        RECT 298.800 529.950 301.050 532.050 ;
        RECT 317.400 531.300 318.600 533.400 ;
        RECT 319.800 534.300 321.600 539.400 ;
        RECT 325.800 534.300 327.600 539.400 ;
        RECT 319.800 532.950 327.600 534.300 ;
        RECT 338.400 536.400 340.200 539.400 ;
        RECT 317.400 530.250 321.150 531.300 ;
        RECT 319.950 530.100 321.150 530.250 ;
        RECT 334.950 529.950 337.050 532.050 ;
        RECT 295.950 526.950 298.050 529.050 ;
        RECT 245.100 525.150 246.900 525.900 ;
        RECT 254.250 525.150 255.900 525.900 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 261.150 522.900 261.900 525.900 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 266.100 525.150 267.900 525.900 ;
        RECT 281.100 524.100 282.900 524.850 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 299.700 525.900 300.900 528.900 ;
        RECT 301.950 526.950 304.050 529.050 ;
        RECT 317.100 527.100 318.900 527.850 ;
        RECT 319.950 526.950 322.050 529.050 ;
        RECT 323.100 527.100 324.900 527.850 ;
        RECT 325.950 526.950 328.050 529.050 ;
        RECT 335.100 528.150 336.900 528.900 ;
        RECT 338.400 527.100 339.600 536.400 ;
        RECT 343.950 532.950 346.050 535.050 ;
        RECT 296.100 525.150 297.900 525.900 ;
        RECT 287.100 524.100 288.900 524.850 ;
        RECT 261.150 521.400 262.050 522.900 ;
        RECT 261.150 520.500 265.200 521.400 ;
        RECT 280.950 520.950 283.050 523.050 ;
        RECT 241.800 507.600 243.600 513.600 ;
        RECT 254.400 518.400 262.200 519.300 ;
        RECT 254.400 507.600 256.200 518.400 ;
        RECT 260.400 508.500 262.200 518.400 ;
        RECT 263.400 509.400 265.200 520.500 ;
        RECT 266.400 508.500 268.200 519.600 ;
        RECT 284.400 513.600 285.600 522.900 ;
        RECT 286.950 520.950 289.050 523.050 ;
        RECT 299.700 520.650 301.050 525.900 ;
        RECT 302.100 525.150 303.900 525.900 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 320.850 522.900 321.900 525.900 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 326.100 525.150 327.900 525.900 ;
        RECT 337.950 525.450 340.050 526.050 ;
        RECT 332.550 524.550 340.050 525.450 ;
        RECT 299.700 519.600 302.400 520.650 ;
        RECT 320.850 519.600 322.050 522.900 ;
        RECT 260.400 507.600 268.200 508.500 ;
        RECT 283.800 507.600 285.600 513.600 ;
        RECT 300.600 507.600 302.400 519.600 ;
        RECT 320.700 507.600 322.500 519.600 ;
        RECT 332.550 514.050 333.450 524.550 ;
        RECT 337.950 523.950 340.050 524.550 ;
        RECT 331.800 511.950 333.900 514.050 ;
        RECT 338.400 513.600 339.600 522.900 ;
        RECT 344.550 514.050 345.450 532.950 ;
        RECT 355.200 532.200 357.000 539.400 ;
        RECT 373.200 535.050 375.000 539.400 ;
        RECT 392.400 536.400 394.200 539.400 ;
        RECT 407.400 536.400 409.200 539.400 ;
        RECT 373.200 533.400 378.600 535.050 ;
        RECT 353.400 531.300 357.000 532.200 ;
        RECT 353.400 527.100 354.600 531.300 ;
        RECT 377.700 530.100 378.600 533.400 ;
        RECT 388.950 529.950 391.050 532.050 ;
        RECT 368.100 527.100 369.900 527.850 ;
        RECT 370.950 526.950 373.050 529.050 ;
        RECT 374.100 527.100 375.900 527.850 ;
        RECT 376.950 526.950 382.050 529.050 ;
        RECT 389.100 528.150 390.900 528.900 ;
        RECT 392.400 527.100 393.600 536.400 ;
        RECT 407.400 533.100 408.600 536.400 ;
        RECT 422.400 534.300 424.200 539.400 ;
        RECT 428.400 534.300 430.200 539.400 ;
        RECT 422.400 532.950 430.200 534.300 ;
        RECT 431.400 533.400 433.200 539.400 ;
        RECT 446.400 536.400 448.200 539.400 ;
        RECT 406.950 529.950 409.050 532.050 ;
        RECT 431.400 531.300 432.600 533.400 ;
        RECT 428.850 530.250 432.600 531.300 ;
        RECT 428.850 530.100 430.050 530.250 ;
        RECT 442.950 529.950 445.050 532.050 ;
        RECT 403.800 526.950 406.050 529.050 ;
        RECT 350.100 524.100 351.900 524.850 ;
        RECT 352.950 523.950 355.050 526.050 ;
        RECT 356.100 524.100 357.900 524.850 ;
        RECT 367.950 523.950 370.050 526.050 ;
        RECT 371.100 525.150 372.900 525.900 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 349.950 520.950 352.050 523.050 ;
        RECT 338.400 507.600 340.200 513.600 ;
        RECT 343.950 511.950 346.050 514.050 ;
        RECT 353.400 513.600 354.600 522.900 ;
        RECT 355.950 520.950 358.050 523.050 ;
        RECT 377.700 519.600 378.600 525.900 ;
        RECT 391.950 523.950 397.050 526.050 ;
        RECT 407.700 525.900 408.900 528.900 ;
        RECT 409.950 526.950 412.050 529.050 ;
        RECT 415.950 526.950 418.050 529.050 ;
        RECT 421.950 526.950 424.050 529.050 ;
        RECT 425.100 527.100 426.900 527.850 ;
        RECT 427.950 526.950 430.050 529.050 ;
        RECT 443.100 528.150 444.900 528.900 ;
        RECT 431.100 527.100 432.900 527.850 ;
        RECT 446.400 527.100 447.600 536.400 ;
        RECT 464.100 531.000 465.900 539.400 ;
        RECT 484.200 535.050 486.000 539.400 ;
        RECT 493.950 535.950 496.050 538.050 ;
        RECT 503.400 536.400 505.200 539.400 ;
        RECT 484.200 533.400 489.600 535.050 ;
        RECT 464.100 529.350 468.300 531.000 ;
        RECT 472.950 529.950 475.050 532.050 ;
        RECT 488.700 530.100 489.600 533.400 ;
        RECT 458.100 527.100 459.900 527.850 ;
        RECT 464.100 527.100 465.900 527.850 ;
        RECT 404.100 525.150 405.900 525.900 ;
        RECT 368.400 518.700 376.200 519.600 ;
        RECT 353.400 507.600 355.200 513.600 ;
        RECT 368.400 507.600 370.200 518.700 ;
        RECT 374.400 507.600 376.200 518.700 ;
        RECT 377.400 507.600 379.200 519.600 ;
        RECT 392.400 513.600 393.600 522.900 ;
        RECT 407.700 520.650 409.050 525.900 ;
        RECT 410.100 525.150 411.900 525.900 ;
        RECT 407.700 519.600 410.400 520.650 ;
        RECT 392.400 507.600 394.200 513.600 ;
        RECT 408.600 507.600 410.400 519.600 ;
        RECT 416.550 517.050 417.450 526.950 ;
        RECT 422.100 525.150 423.900 525.900 ;
        RECT 424.950 523.950 427.050 526.050 ;
        RECT 428.100 522.900 429.150 525.900 ;
        RECT 430.950 523.950 433.050 526.050 ;
        RECT 445.950 523.950 451.050 526.050 ;
        RECT 457.950 523.950 460.200 526.050 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 467.400 524.100 468.300 529.350 ;
        RECT 427.950 519.600 429.150 522.900 ;
        RECT 415.950 514.950 418.050 517.050 ;
        RECT 427.500 507.600 429.300 519.600 ;
        RECT 446.400 513.600 447.600 522.900 ;
        RECT 460.950 520.950 463.050 523.050 ;
        RECT 466.950 522.450 469.050 523.050 ;
        RECT 473.550 522.450 474.450 529.950 ;
        RECT 479.100 527.100 480.900 527.850 ;
        RECT 481.800 526.950 484.050 529.050 ;
        RECT 485.100 527.100 486.900 527.850 ;
        RECT 487.950 526.950 493.050 529.050 ;
        RECT 494.550 526.050 495.450 535.950 ;
        RECT 499.950 529.950 502.050 532.050 ;
        RECT 500.100 528.150 501.900 528.900 ;
        RECT 503.400 527.100 504.600 536.400 ;
        RECT 520.200 535.050 522.000 539.400 ;
        RECT 520.200 533.400 525.600 535.050 ;
        RECT 524.700 530.100 525.600 533.400 ;
        RECT 542.100 531.000 543.900 539.400 ;
        RECT 550.950 535.950 553.050 538.050 ;
        RECT 542.100 529.350 546.300 531.000 ;
        RECT 515.100 527.100 516.900 527.850 ;
        RECT 517.950 526.950 520.050 529.050 ;
        RECT 521.100 527.100 522.900 527.850 ;
        RECT 523.950 526.950 529.050 529.050 ;
        RECT 536.100 527.100 537.900 527.850 ;
        RECT 542.100 527.100 543.900 527.850 ;
        RECT 478.950 523.950 481.050 526.050 ;
        RECT 482.100 525.150 483.900 525.900 ;
        RECT 484.950 523.950 487.050 526.050 ;
        RECT 466.950 521.550 474.450 522.450 ;
        RECT 466.950 520.950 469.050 521.550 ;
        RECT 461.100 519.150 462.900 519.900 ;
        RECT 467.400 514.800 468.300 519.900 ;
        RECT 488.700 519.600 489.600 525.900 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 502.950 525.450 505.050 526.050 ;
        RECT 502.950 525.000 510.450 525.450 ;
        RECT 502.950 524.550 511.050 525.000 ;
        RECT 502.950 523.950 505.050 524.550 ;
        RECT 461.700 513.900 468.300 514.800 ;
        RECT 461.700 513.600 463.200 513.900 ;
        RECT 446.400 507.600 448.200 513.600 ;
        RECT 461.400 507.600 463.200 513.600 ;
        RECT 467.400 513.600 468.300 513.900 ;
        RECT 479.400 518.700 487.200 519.600 ;
        RECT 467.400 507.600 469.200 513.600 ;
        RECT 479.400 507.600 481.200 518.700 ;
        RECT 485.400 507.600 487.200 518.700 ;
        RECT 488.400 507.600 490.200 519.600 ;
        RECT 503.400 513.600 504.600 522.900 ;
        RECT 508.950 520.950 511.050 524.550 ;
        RECT 514.950 523.950 517.050 526.050 ;
        RECT 518.100 525.150 519.900 525.900 ;
        RECT 520.950 523.950 523.050 526.050 ;
        RECT 524.700 519.600 525.600 525.900 ;
        RECT 535.800 523.950 538.050 526.050 ;
        RECT 541.950 523.950 544.050 526.050 ;
        RECT 545.400 524.100 546.300 529.350 ;
        RECT 538.950 520.950 541.050 523.050 ;
        RECT 544.950 522.450 547.050 523.050 ;
        RECT 551.550 522.450 552.450 535.950 ;
        RECT 557.400 534.300 559.200 539.400 ;
        RECT 563.400 534.300 565.200 539.400 ;
        RECT 557.400 532.950 565.200 534.300 ;
        RECT 566.400 533.400 568.200 539.400 ;
        RECT 566.400 531.300 567.600 533.400 ;
        RECT 583.800 532.500 585.600 539.400 ;
        RECT 589.800 532.500 591.600 539.400 ;
        RECT 595.800 532.500 597.600 539.400 ;
        RECT 601.800 532.500 603.600 539.400 ;
        RECT 619.800 532.500 621.600 539.400 ;
        RECT 625.800 532.500 627.600 539.400 ;
        RECT 631.800 532.500 633.600 539.400 ;
        RECT 637.800 532.500 639.600 539.400 ;
        RECT 650.400 534.300 652.200 539.400 ;
        RECT 656.400 534.300 658.200 539.400 ;
        RECT 650.400 532.950 658.200 534.300 ;
        RECT 659.400 533.400 661.200 539.400 ;
        RECT 563.850 530.250 567.600 531.300 ;
        RECT 582.900 531.300 585.600 532.500 ;
        RECT 587.700 531.300 591.600 532.500 ;
        RECT 593.700 531.300 597.600 532.500 ;
        RECT 599.700 531.300 603.600 532.500 ;
        RECT 618.900 531.300 621.600 532.500 ;
        RECT 623.700 531.300 627.600 532.500 ;
        RECT 629.700 531.300 633.600 532.500 ;
        RECT 635.700 531.300 639.600 532.500 ;
        RECT 659.400 531.300 660.600 533.400 ;
        RECT 676.200 532.200 678.000 539.400 ;
        RECT 689.400 534.300 691.200 539.400 ;
        RECT 695.400 534.300 697.200 539.400 ;
        RECT 689.400 532.950 697.200 534.300 ;
        RECT 698.400 533.400 700.200 539.400 ;
        RECT 563.850 530.100 565.050 530.250 ;
        RECT 556.950 526.950 559.050 529.050 ;
        RECT 560.100 527.100 561.900 527.850 ;
        RECT 562.950 526.950 565.050 529.050 ;
        RECT 566.100 527.100 567.900 527.850 ;
        RECT 582.900 527.100 583.800 531.300 ;
        RECT 587.700 530.400 588.900 531.300 ;
        RECT 593.700 530.400 594.900 531.300 ;
        RECT 599.700 530.400 600.900 531.300 ;
        RECT 584.700 529.200 588.900 530.400 ;
        RECT 584.700 528.600 586.500 529.200 ;
        RECT 557.100 525.150 558.900 525.900 ;
        RECT 559.800 523.950 562.050 526.050 ;
        RECT 563.100 522.900 564.150 525.900 ;
        RECT 577.950 523.950 583.050 526.050 ;
        RECT 544.950 521.550 552.450 522.450 ;
        RECT 544.950 520.950 547.050 521.550 ;
        RECT 515.400 518.700 523.200 519.600 ;
        RECT 503.400 507.600 505.200 513.600 ;
        RECT 515.400 507.600 517.200 518.700 ;
        RECT 521.400 507.600 523.200 518.700 ;
        RECT 524.400 507.600 526.200 519.600 ;
        RECT 539.100 519.150 540.900 519.900 ;
        RECT 545.400 514.800 546.300 519.900 ;
        RECT 562.950 519.600 564.150 522.900 ;
        RECT 582.900 521.700 583.800 522.900 ;
        RECT 587.700 521.700 588.900 529.200 ;
        RECT 590.700 529.200 594.900 530.400 ;
        RECT 590.700 528.600 592.500 529.200 ;
        RECT 593.700 521.700 594.900 529.200 ;
        RECT 596.700 529.200 600.900 530.400 ;
        RECT 596.700 528.600 598.500 529.200 ;
        RECT 599.700 521.700 600.900 529.200 ;
        RECT 602.100 527.100 603.900 527.850 ;
        RECT 618.900 527.100 619.800 531.300 ;
        RECT 623.700 530.400 624.900 531.300 ;
        RECT 629.700 530.400 630.900 531.300 ;
        RECT 635.700 530.400 636.900 531.300 ;
        RECT 620.700 529.200 624.900 530.400 ;
        RECT 620.700 528.600 622.500 529.200 ;
        RECT 616.950 523.950 622.050 526.050 ;
        RECT 618.900 521.700 619.800 522.900 ;
        RECT 623.700 521.700 624.900 529.200 ;
        RECT 626.700 529.200 630.900 530.400 ;
        RECT 626.700 528.600 628.500 529.200 ;
        RECT 629.700 521.700 630.900 529.200 ;
        RECT 632.700 529.200 636.900 530.400 ;
        RECT 656.850 530.250 660.600 531.300 ;
        RECT 674.400 531.300 678.000 532.200 ;
        RECT 698.400 531.300 699.600 533.400 ;
        RECT 715.200 532.200 717.000 539.400 ;
        RECT 656.850 530.100 658.050 530.250 ;
        RECT 632.700 528.600 634.500 529.200 ;
        RECT 635.700 521.700 636.900 529.200 ;
        RECT 638.100 527.100 639.900 527.850 ;
        RECT 649.950 526.950 652.050 529.050 ;
        RECT 653.100 527.100 654.900 527.850 ;
        RECT 655.950 526.950 658.050 529.050 ;
        RECT 659.100 527.100 660.900 527.850 ;
        RECT 664.950 526.950 667.050 529.050 ;
        RECT 674.400 527.100 675.600 531.300 ;
        RECT 695.850 530.250 699.600 531.300 ;
        RECT 713.400 531.300 717.000 532.200 ;
        RECT 722.550 533.400 724.350 539.400 ;
        RECT 730.650 536.400 732.450 539.400 ;
        RECT 738.450 536.400 740.250 539.400 ;
        RECT 746.250 537.300 748.050 539.400 ;
        RECT 746.250 536.400 750.000 537.300 ;
        RECT 730.650 535.500 731.700 536.400 ;
        RECT 727.950 534.300 731.700 535.500 ;
        RECT 739.200 534.600 740.250 536.400 ;
        RECT 748.950 535.500 750.000 536.400 ;
        RECT 727.950 533.400 730.050 534.300 ;
        RECT 695.850 530.100 697.050 530.250 ;
        RECT 685.950 526.950 691.050 529.050 ;
        RECT 692.100 527.100 693.900 527.850 ;
        RECT 694.950 526.950 697.050 529.050 ;
        RECT 698.100 527.100 699.900 527.850 ;
        RECT 713.400 527.100 714.600 531.300 ;
        RECT 722.550 529.050 723.750 533.400 ;
        RECT 735.150 532.200 736.950 534.000 ;
        RECT 739.200 533.550 744.150 534.600 ;
        RECT 742.350 532.800 744.150 533.550 ;
        RECT 745.650 532.800 747.450 534.600 ;
        RECT 748.950 533.400 751.050 535.500 ;
        RECT 754.050 533.400 755.850 539.400 ;
        RECT 769.200 535.050 771.000 539.400 ;
        RECT 769.200 533.400 774.600 535.050 ;
        RECT 736.050 531.900 736.950 532.200 ;
        RECT 746.100 531.900 747.150 532.800 ;
        RECT 736.050 531.000 747.150 531.900 ;
        RECT 736.050 530.100 736.950 531.000 ;
        RECT 746.100 529.800 747.150 531.000 ;
        RECT 722.550 526.950 723.900 529.050 ;
        RECT 724.950 526.950 727.050 529.050 ;
        RECT 728.100 527.250 728.850 529.050 ;
        RECT 736.950 526.950 739.050 529.050 ;
        RECT 742.950 526.950 745.050 529.050 ;
        RECT 746.100 528.600 753.000 529.800 ;
        RECT 746.100 528.000 747.900 528.600 ;
        RECT 752.100 527.850 753.000 528.600 ;
        RECT 749.100 527.100 750.900 527.700 ;
        RECT 650.100 525.150 651.900 525.900 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 656.100 522.900 657.150 525.900 ;
        RECT 658.950 523.950 661.050 526.050 ;
        RECT 582.900 520.500 585.600 521.700 ;
        RECT 587.700 520.500 591.600 521.700 ;
        RECT 593.700 520.500 597.600 521.700 ;
        RECT 599.700 520.500 603.600 521.700 ;
        RECT 618.900 520.500 621.600 521.700 ;
        RECT 623.700 520.500 627.600 521.700 ;
        RECT 629.700 520.500 633.600 521.700 ;
        RECT 635.700 520.500 639.600 521.700 ;
        RECT 539.700 513.900 546.300 514.800 ;
        RECT 539.700 513.600 541.200 513.900 ;
        RECT 539.400 507.600 541.200 513.600 ;
        RECT 545.400 513.600 546.300 513.900 ;
        RECT 545.400 507.600 547.200 513.600 ;
        RECT 562.500 507.600 564.300 519.600 ;
        RECT 583.800 507.600 585.600 520.500 ;
        RECT 589.800 507.600 591.600 520.500 ;
        RECT 595.800 507.600 597.600 520.500 ;
        RECT 601.800 507.600 603.600 520.500 ;
        RECT 619.800 507.600 621.600 520.500 ;
        RECT 625.800 507.600 627.600 520.500 ;
        RECT 631.800 507.600 633.600 520.500 ;
        RECT 637.800 507.600 639.600 520.500 ;
        RECT 655.950 519.600 657.150 522.900 ;
        RECT 655.500 507.600 657.300 519.600 ;
        RECT 665.550 517.050 666.450 526.950 ;
        RECT 671.100 524.100 672.900 524.850 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 689.100 525.150 690.900 525.900 ;
        RECT 677.100 524.100 678.900 524.850 ;
        RECT 691.950 523.950 694.050 526.050 ;
        RECT 670.950 520.950 673.050 523.050 ;
        RECT 664.950 514.950 667.050 517.050 ;
        RECT 674.400 513.600 675.600 522.900 ;
        RECT 676.950 520.950 679.050 523.050 ;
        RECT 695.100 522.900 696.150 525.900 ;
        RECT 697.950 523.950 700.050 526.050 ;
        RECT 710.100 524.100 711.900 524.850 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 716.100 524.100 717.900 524.850 ;
        RECT 694.950 519.600 696.150 522.900 ;
        RECT 709.950 520.950 712.050 523.050 ;
        RECT 674.400 507.600 676.200 513.600 ;
        RECT 694.500 507.600 696.300 519.600 ;
        RECT 713.400 513.600 714.600 522.900 ;
        RECT 715.950 520.950 718.050 523.050 ;
        RECT 722.550 519.600 723.750 526.950 ;
        RECT 746.100 526.200 750.900 527.100 ;
        RECT 749.100 525.900 750.900 526.200 ;
        RECT 752.100 526.050 753.900 527.850 ;
        RECT 724.950 521.400 726.750 523.200 ;
        RECT 725.850 520.200 730.050 521.400 ;
        RECT 736.050 520.200 736.950 525.900 ;
        RECT 744.750 521.100 746.550 521.400 ;
        RECT 713.400 507.600 715.200 513.600 ;
        RECT 722.550 507.600 724.350 519.600 ;
        RECT 727.950 519.300 730.050 520.200 ;
        RECT 730.950 519.300 736.950 520.200 ;
        RECT 738.150 520.800 746.550 521.100 ;
        RECT 754.950 520.800 755.850 533.400 ;
        RECT 773.700 530.100 774.600 533.400 ;
        RECT 785.400 534.300 787.200 539.400 ;
        RECT 791.400 534.300 793.200 539.400 ;
        RECT 785.400 532.950 793.200 534.300 ;
        RECT 794.400 533.400 796.200 539.400 ;
        RECT 809.400 536.400 811.200 539.400 ;
        RECT 794.400 531.300 795.600 533.400 ;
        RECT 791.850 530.250 795.600 531.300 ;
        RECT 791.850 530.100 793.050 530.250 ;
        RECT 805.950 529.950 808.050 532.050 ;
        RECT 764.100 527.100 765.900 527.850 ;
        RECT 766.950 526.950 769.050 529.050 ;
        RECT 772.950 528.450 775.050 529.050 ;
        RECT 770.100 527.100 771.900 527.850 ;
        RECT 772.950 527.550 780.450 528.450 ;
        RECT 772.950 526.950 775.050 527.550 ;
        RECT 763.950 523.950 766.050 526.050 ;
        RECT 767.100 525.150 768.900 525.900 ;
        RECT 769.950 523.950 772.050 526.050 ;
        RECT 738.150 520.200 755.850 520.800 ;
        RECT 730.950 518.400 731.850 519.300 ;
        RECT 729.150 516.600 731.850 518.400 ;
        RECT 732.750 518.100 734.550 518.400 ;
        RECT 738.150 518.100 739.050 520.200 ;
        RECT 744.750 519.600 755.850 520.200 ;
        RECT 773.700 519.600 774.600 525.900 ;
        RECT 732.750 517.200 739.050 518.100 ;
        RECT 739.950 518.700 741.750 519.300 ;
        RECT 739.950 517.500 747.450 518.700 ;
        RECT 732.750 516.600 734.550 517.200 ;
        RECT 746.250 516.600 747.450 517.500 ;
        RECT 727.950 513.600 731.850 515.700 ;
        RECT 736.950 515.550 738.750 516.300 ;
        RECT 741.750 515.550 743.550 516.300 ;
        RECT 736.950 514.500 743.550 515.550 ;
        RECT 746.250 514.500 751.050 516.600 ;
        RECT 730.050 507.600 731.850 513.600 ;
        RECT 737.850 507.600 739.650 514.500 ;
        RECT 746.250 513.600 747.450 514.500 ;
        RECT 745.650 507.600 747.450 513.600 ;
        RECT 754.050 507.600 755.850 519.600 ;
        RECT 764.400 518.700 772.200 519.600 ;
        RECT 764.400 507.600 766.200 518.700 ;
        RECT 770.400 507.600 772.200 518.700 ;
        RECT 773.400 507.600 775.200 519.600 ;
        RECT 779.550 511.050 780.450 527.550 ;
        RECT 784.800 526.950 787.050 529.050 ;
        RECT 788.100 527.100 789.900 527.850 ;
        RECT 790.950 526.950 793.050 529.050 ;
        RECT 806.100 528.150 807.900 528.900 ;
        RECT 794.100 527.100 795.900 527.850 ;
        RECT 809.400 527.100 810.600 536.400 ;
        RECT 821.400 534.300 823.200 539.400 ;
        RECT 827.400 534.300 829.200 539.400 ;
        RECT 821.400 532.950 829.200 534.300 ;
        RECT 830.400 533.400 832.200 539.400 ;
        RECT 830.400 531.300 831.600 533.400 ;
        RECT 847.200 532.200 849.000 539.400 ;
        RECT 827.850 530.250 831.600 531.300 ;
        RECT 845.400 531.300 849.000 532.200 ;
        RECT 827.850 530.100 829.050 530.250 ;
        RECT 820.950 526.950 823.050 529.050 ;
        RECT 824.100 527.100 825.900 527.850 ;
        RECT 826.950 526.950 829.050 529.050 ;
        RECT 830.100 527.100 831.900 527.850 ;
        RECT 845.400 527.100 846.600 531.300 ;
        RECT 785.100 525.150 786.900 525.900 ;
        RECT 787.950 523.950 790.050 526.050 ;
        RECT 791.100 522.900 792.150 525.900 ;
        RECT 793.950 523.950 796.050 526.050 ;
        RECT 808.950 523.950 814.050 526.050 ;
        RECT 821.100 525.150 822.900 525.900 ;
        RECT 823.950 523.950 826.050 526.050 ;
        RECT 790.950 519.600 792.150 522.900 ;
        RECT 778.950 508.950 781.050 511.050 ;
        RECT 790.500 507.600 792.300 519.600 ;
        RECT 794.550 517.050 795.450 523.950 ;
        RECT 827.100 522.900 828.150 525.900 ;
        RECT 842.100 524.100 843.900 524.850 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 848.100 524.100 849.900 524.850 ;
        RECT 853.950 523.950 856.050 526.050 ;
        RECT 793.950 514.950 796.050 517.050 ;
        RECT 809.400 513.600 810.600 522.900 ;
        RECT 826.950 519.600 828.150 522.900 ;
        RECT 809.400 507.600 811.200 513.600 ;
        RECT 826.500 507.600 828.300 519.600 ;
        RECT 845.400 513.600 846.600 522.900 ;
        RECT 845.400 507.600 847.200 513.600 ;
        RECT 854.550 511.050 855.450 523.950 ;
        RECT 853.950 508.950 856.050 511.050 ;
        RECT 14.700 491.400 16.500 503.400 ;
        RECT 34.500 491.400 36.300 503.400 ;
        RECT 53.400 497.400 55.200 503.400 ;
        RECT 53.700 497.100 55.200 497.400 ;
        RECT 59.400 497.400 61.200 503.400 ;
        RECT 59.400 497.100 60.300 497.400 ;
        RECT 53.700 496.200 60.300 497.100 ;
        RECT 67.950 496.950 70.050 499.050 ;
        RECT 73.800 497.400 75.600 503.400 ;
        RECT 74.700 497.100 75.600 497.400 ;
        RECT 79.800 497.400 81.600 503.400 ;
        RECT 79.800 497.100 81.300 497.400 ;
        RECT 14.850 488.100 16.050 491.400 ;
        RECT 34.950 488.100 36.150 491.400 ;
        RECT 53.100 491.100 54.900 491.850 ;
        RECT 59.400 491.100 60.300 496.200 ;
        RECT 10.950 484.950 13.050 487.050 ;
        RECT 14.850 485.100 15.900 488.100 ;
        RECT 16.950 484.950 19.050 487.050 ;
        RECT 20.100 485.100 21.900 485.850 ;
        RECT 29.100 485.100 30.900 485.850 ;
        RECT 31.950 484.950 34.200 487.050 ;
        RECT 35.100 485.100 36.150 488.100 ;
        RECT 52.950 487.950 55.200 490.050 ;
        RECT 58.950 487.950 64.050 490.050 ;
        RECT 68.550 489.450 69.450 496.950 ;
        RECT 74.700 496.200 81.300 497.100 ;
        RECT 74.700 491.100 75.600 496.200 ;
        RECT 92.400 492.300 94.200 503.400 ;
        RECT 98.400 492.300 100.200 503.400 ;
        RECT 80.100 491.100 81.900 491.850 ;
        RECT 92.400 491.400 100.200 492.300 ;
        RECT 101.400 491.400 103.200 503.400 ;
        RECT 115.800 497.400 117.600 503.400 ;
        RECT 73.950 489.450 76.050 490.050 ;
        RECT 68.550 488.550 76.050 489.450 ;
        RECT 73.950 487.950 76.050 488.550 ;
        RECT 79.950 487.950 82.050 490.050 ;
        RECT 37.950 484.950 40.200 487.050 ;
        RECT 49.950 484.950 52.050 487.050 ;
        RECT 55.950 484.950 58.050 487.050 ;
        RECT 11.100 483.150 12.900 483.900 ;
        RECT 13.950 481.950 16.050 484.050 ;
        RECT 17.100 483.150 18.900 483.900 ;
        RECT 19.950 481.950 22.200 484.050 ;
        RECT 28.950 481.950 31.050 484.050 ;
        RECT 32.100 483.150 33.900 483.900 ;
        RECT 34.950 481.950 37.050 484.050 ;
        RECT 38.100 483.150 39.900 483.900 ;
        RECT 50.100 483.150 51.900 483.900 ;
        RECT 56.100 483.150 57.900 483.900 ;
        RECT 59.400 481.650 60.300 486.900 ;
        RECT 13.950 480.750 15.150 480.900 ;
        RECT 11.400 479.700 15.150 480.750 ;
        RECT 35.850 480.750 37.050 480.900 ;
        RECT 35.850 479.700 39.600 480.750 ;
        RECT 11.400 477.600 12.600 479.700 ;
        RECT 10.800 471.600 12.600 477.600 ;
        RECT 13.800 476.700 21.600 478.050 ;
        RECT 13.800 471.600 15.600 476.700 ;
        RECT 19.800 471.600 21.600 476.700 ;
        RECT 29.400 476.700 37.200 478.050 ;
        RECT 29.400 471.600 31.200 476.700 ;
        RECT 35.400 471.600 37.200 476.700 ;
        RECT 38.400 477.600 39.600 479.700 ;
        RECT 56.100 480.000 60.300 481.650 ;
        RECT 74.700 481.650 75.600 486.900 ;
        RECT 76.950 484.950 79.050 487.050 ;
        RECT 82.800 484.950 85.050 487.050 ;
        RECT 91.800 484.950 94.050 487.050 ;
        RECT 95.100 485.100 96.900 485.850 ;
        RECT 97.950 484.950 100.050 487.050 ;
        RECT 101.700 485.100 102.600 491.400 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 77.100 483.150 78.900 483.900 ;
        RECT 83.100 483.150 84.900 483.900 ;
        RECT 92.100 483.150 93.900 483.900 ;
        RECT 94.950 481.950 97.200 484.050 ;
        RECT 98.100 483.150 99.900 483.900 ;
        RECT 100.950 483.450 103.050 484.050 ;
        RECT 107.550 483.450 108.450 490.950 ;
        RECT 116.400 488.100 117.600 497.400 ;
        RECT 128.400 492.300 130.200 503.400 ;
        RECT 134.400 492.300 136.200 503.400 ;
        RECT 128.400 491.400 136.200 492.300 ;
        RECT 137.400 491.400 139.200 503.400 ;
        RECT 154.500 491.400 156.300 503.400 ;
        RECT 173.400 497.400 175.200 503.400 ;
        RECT 173.700 497.100 175.200 497.400 ;
        RECT 179.400 497.400 181.200 503.400 ;
        RECT 179.400 497.100 180.300 497.400 ;
        RECT 173.700 496.200 180.300 497.100 ;
        RECT 184.950 496.950 187.050 499.050 ;
        RECT 112.950 484.950 118.050 487.050 ;
        RECT 124.950 484.950 130.050 487.050 ;
        RECT 131.100 485.100 132.900 485.850 ;
        RECT 133.950 484.950 136.050 487.050 ;
        RECT 137.700 485.100 138.600 491.400 ;
        RECT 154.950 488.100 156.150 491.400 ;
        RECT 173.100 491.100 174.900 491.850 ;
        RECT 179.400 491.100 180.300 496.200 ;
        RECT 149.100 485.100 150.900 485.850 ;
        RECT 151.950 484.950 154.050 487.050 ;
        RECT 155.100 485.100 156.150 488.100 ;
        RECT 172.950 487.950 175.200 490.050 ;
        RECT 178.950 489.450 181.050 490.050 ;
        RECT 185.550 489.450 186.450 496.950 ;
        RECT 197.700 491.400 199.500 503.400 ;
        RECT 214.800 497.400 216.600 503.400 ;
        RECT 178.950 488.550 186.450 489.450 ;
        RECT 178.950 487.950 181.050 488.550 ;
        RECT 197.850 488.100 199.050 491.400 ;
        RECT 215.400 488.100 216.600 497.400 ;
        RECT 229.500 491.400 231.300 503.400 ;
        RECT 235.800 497.400 237.600 503.400 ;
        RECT 247.800 497.400 249.600 503.400 ;
        RECT 157.950 484.950 160.050 487.050 ;
        RECT 169.950 484.950 172.050 487.050 ;
        RECT 175.950 484.950 178.050 487.050 ;
        RECT 100.950 482.550 108.450 483.450 ;
        RECT 100.950 481.950 103.050 482.550 ;
        RECT 74.700 480.000 78.900 481.650 ;
        RECT 38.400 471.600 40.200 477.600 ;
        RECT 56.100 471.600 57.900 480.000 ;
        RECT 77.100 471.600 78.900 480.000 ;
        RECT 101.700 477.600 102.600 480.900 ;
        RECT 97.200 475.950 102.600 477.600 ;
        RECT 97.200 471.600 99.000 475.950 ;
        RECT 116.400 474.600 117.600 483.900 ;
        RECT 128.100 483.150 129.900 483.900 ;
        RECT 119.100 482.100 120.900 482.850 ;
        RECT 130.950 481.950 133.050 484.050 ;
        RECT 134.100 483.150 135.900 483.900 ;
        RECT 136.950 481.950 142.050 484.050 ;
        RECT 148.950 481.950 151.050 484.050 ;
        RECT 152.100 483.150 153.900 483.900 ;
        RECT 154.800 481.950 157.050 484.050 ;
        RECT 158.100 483.150 159.900 483.900 ;
        RECT 170.100 483.150 171.900 483.900 ;
        RECT 176.100 483.150 177.900 483.900 ;
        RECT 179.400 481.650 180.300 486.900 ;
        RECT 193.950 484.950 196.050 487.050 ;
        RECT 197.850 485.100 198.900 488.100 ;
        RECT 199.950 484.950 202.050 487.050 ;
        RECT 203.100 485.100 204.900 485.850 ;
        RECT 211.950 484.950 217.050 487.050 ;
        RECT 229.800 485.100 231.000 491.400 ;
        RECT 236.400 490.500 237.600 497.400 ;
        RECT 248.700 497.100 249.600 497.400 ;
        RECT 253.800 497.400 255.600 503.400 ;
        RECT 268.800 497.400 270.600 503.400 ;
        RECT 253.800 497.100 255.300 497.400 ;
        RECT 248.700 496.200 255.300 497.100 ;
        RECT 248.700 491.100 249.600 496.200 ;
        RECT 254.100 491.100 255.900 491.850 ;
        RECT 231.900 489.600 237.600 490.500 ;
        RECT 231.900 488.700 233.850 489.600 ;
        RECT 232.950 485.100 233.850 488.700 ;
        RECT 244.950 487.950 250.050 490.050 ;
        RECT 253.950 487.950 256.050 490.050 ;
        RECT 269.400 488.100 270.600 497.400 ;
        RECT 284.400 497.400 286.200 503.400 ;
        RECT 236.100 485.100 237.900 485.850 ;
        RECT 194.100 483.150 195.900 483.900 ;
        RECT 196.950 481.950 199.050 484.050 ;
        RECT 200.100 483.150 201.900 483.900 ;
        RECT 202.950 481.950 205.050 484.050 ;
        RECT 118.950 478.950 121.050 481.050 ;
        RECT 137.700 477.600 138.600 480.900 ;
        RECT 155.850 480.750 157.050 480.900 ;
        RECT 155.850 479.700 159.600 480.750 ;
        RECT 115.800 471.600 117.600 474.600 ;
        RECT 133.200 475.950 138.600 477.600 ;
        RECT 149.400 476.700 157.200 478.050 ;
        RECT 133.200 471.600 135.000 475.950 ;
        RECT 149.400 471.600 151.200 476.700 ;
        RECT 155.400 471.600 157.200 476.700 ;
        RECT 158.400 477.600 159.600 479.700 ;
        RECT 176.100 480.000 180.300 481.650 ;
        RECT 158.400 471.600 160.200 477.600 ;
        RECT 176.100 471.600 177.900 480.000 ;
        RECT 187.950 478.950 190.050 481.050 ;
        RECT 196.950 480.750 198.150 480.900 ;
        RECT 194.400 479.700 198.150 480.750 ;
        RECT 188.550 475.050 189.450 478.950 ;
        RECT 194.400 477.600 195.600 479.700 ;
        RECT 187.950 472.950 190.050 475.050 ;
        RECT 193.800 471.600 195.600 477.600 ;
        RECT 196.800 476.700 204.600 478.050 ;
        RECT 196.800 471.600 198.600 476.700 ;
        RECT 202.800 471.600 204.600 476.700 ;
        RECT 215.400 474.600 216.600 483.900 ;
        RECT 218.100 482.100 219.900 482.850 ;
        RECT 226.950 481.950 232.050 484.050 ;
        RECT 217.950 478.950 220.050 481.050 ;
        RECT 233.100 480.900 233.850 485.100 ;
        RECT 235.950 481.950 241.200 484.050 ;
        RECT 229.800 477.600 231.000 480.900 ;
        RECT 232.950 480.300 233.850 480.900 ;
        RECT 231.900 479.400 233.850 480.300 ;
        RECT 248.700 481.650 249.600 486.900 ;
        RECT 250.950 484.950 253.050 487.050 ;
        RECT 256.950 484.950 259.050 487.050 ;
        RECT 265.950 484.950 271.050 487.050 ;
        RECT 281.100 485.100 282.900 485.850 ;
        RECT 251.100 483.150 252.900 483.900 ;
        RECT 257.100 483.150 258.900 483.900 ;
        RECT 248.700 480.000 252.900 481.650 ;
        RECT 231.900 478.500 237.000 479.400 ;
        RECT 214.800 471.600 216.600 474.600 ;
        RECT 229.500 471.600 231.300 477.600 ;
        RECT 235.800 474.600 237.000 478.500 ;
        RECT 235.800 471.600 237.600 474.600 ;
        RECT 251.100 471.600 252.900 480.000 ;
        RECT 269.400 474.600 270.600 483.900 ;
        RECT 272.100 482.100 273.900 482.850 ;
        RECT 280.950 481.950 283.050 484.050 ;
        RECT 271.950 478.950 274.050 481.050 ;
        RECT 284.400 480.300 285.450 497.400 ;
        RECT 291.000 491.400 292.800 503.400 ;
        RECT 305.400 497.400 307.200 503.400 ;
        RECT 313.950 501.450 318.000 502.050 ;
        RECT 313.950 499.950 318.450 501.450 ;
        RECT 286.950 484.950 289.050 490.050 ;
        RECT 291.000 485.100 292.050 491.400 ;
        RECT 295.950 487.950 298.050 490.050 ;
        RECT 301.950 487.950 304.050 490.050 ;
        RECT 305.400 488.100 306.600 497.400 ;
        RECT 307.950 487.950 310.050 490.050 ;
        RECT 287.100 483.150 288.900 483.900 ;
        RECT 289.950 483.450 292.050 484.050 ;
        RECT 296.550 483.450 297.450 487.950 ;
        RECT 317.550 487.050 318.450 499.950 ;
        RECT 325.800 497.400 327.600 503.400 ;
        RECT 343.800 497.400 345.600 503.400 ;
        RECT 359.400 497.400 361.200 503.400 ;
        RECT 322.950 487.950 325.050 490.050 ;
        RECT 326.400 488.100 327.600 497.400 ;
        RECT 340.950 490.050 343.050 493.050 ;
        RECT 328.950 487.950 331.050 490.050 ;
        RECT 340.800 487.950 343.050 490.050 ;
        RECT 344.400 488.100 345.600 497.400 ;
        RECT 359.700 497.100 361.200 497.400 ;
        RECT 365.400 497.400 367.200 503.400 ;
        RECT 365.400 497.100 366.300 497.400 ;
        RECT 359.700 496.200 366.300 497.100 ;
        RECT 359.100 491.100 360.900 491.850 ;
        RECT 365.400 491.100 366.300 496.200 ;
        RECT 377.400 492.300 379.200 503.400 ;
        RECT 383.400 492.300 385.200 503.400 ;
        RECT 377.400 491.400 385.200 492.300 ;
        RECT 386.400 491.400 388.200 503.400 ;
        RECT 346.950 487.950 349.200 490.050 ;
        RECT 358.950 487.950 361.050 490.050 ;
        RECT 364.950 487.950 370.050 490.050 ;
        RECT 302.100 486.150 303.900 486.900 ;
        RECT 304.950 484.950 307.050 487.050 ;
        RECT 308.100 486.150 309.900 486.900 ;
        RECT 316.950 484.950 319.050 487.050 ;
        RECT 323.100 486.150 324.900 486.900 ;
        RECT 325.950 484.950 328.050 487.050 ;
        RECT 329.100 486.150 330.900 486.900 ;
        RECT 341.100 486.150 342.900 486.900 ;
        RECT 343.800 484.950 346.050 487.050 ;
        RECT 347.100 486.150 348.900 486.900 ;
        RECT 355.950 484.950 358.050 487.050 ;
        RECT 361.950 484.950 364.050 487.050 ;
        RECT 289.950 482.550 297.450 483.450 ;
        RECT 289.950 481.950 292.050 482.550 ;
        RECT 281.400 479.100 288.900 480.300 ;
        RECT 268.800 471.600 270.600 474.600 ;
        RECT 281.400 471.600 283.200 479.100 ;
        RECT 287.100 478.500 288.900 479.100 ;
        RECT 289.950 477.600 290.850 480.900 ;
        RECT 305.400 479.700 306.600 483.900 ;
        RECT 326.400 479.700 327.600 483.900 ;
        RECT 344.400 479.700 345.600 483.900 ;
        RECT 356.100 483.150 357.900 483.900 ;
        RECT 362.100 483.150 363.900 483.900 ;
        RECT 365.400 481.650 366.300 486.900 ;
        RECT 376.950 484.950 379.050 487.050 ;
        RECT 380.100 485.100 381.900 485.850 ;
        RECT 382.950 484.950 385.050 487.050 ;
        RECT 386.700 485.100 387.600 491.400 ;
        RECT 394.950 490.950 397.050 493.050 ;
        RECT 404.700 491.400 406.500 503.400 ;
        RECT 415.950 499.950 418.050 502.050 ;
        RECT 395.550 484.050 396.450 490.950 ;
        RECT 404.850 488.100 406.050 491.400 ;
        RECT 400.950 484.950 403.050 487.050 ;
        RECT 404.850 485.100 405.900 488.100 ;
        RECT 406.950 484.950 409.050 487.050 ;
        RECT 410.100 485.100 411.900 485.850 ;
        RECT 377.100 483.150 378.900 483.900 ;
        RECT 379.950 481.950 382.050 484.050 ;
        RECT 383.100 483.150 384.900 483.900 ;
        RECT 385.950 483.450 388.050 484.050 ;
        RECT 385.950 482.550 393.450 483.450 ;
        RECT 385.950 481.950 388.050 482.550 ;
        RECT 305.400 478.800 309.000 479.700 ;
        RECT 288.900 475.800 290.850 477.600 ;
        RECT 288.900 471.600 290.700 475.800 ;
        RECT 307.200 471.600 309.000 478.800 ;
        RECT 324.000 478.800 327.600 479.700 ;
        RECT 342.000 478.800 345.600 479.700 ;
        RECT 362.100 480.000 366.300 481.650 ;
        RECT 324.000 471.600 325.800 478.800 ;
        RECT 342.000 471.600 343.800 478.800 ;
        RECT 362.100 471.600 363.900 480.000 ;
        RECT 386.700 477.600 387.600 480.900 ;
        RECT 382.200 475.950 387.600 477.600 ;
        RECT 382.200 471.600 384.000 475.950 ;
        RECT 392.550 475.050 393.450 482.550 ;
        RECT 394.950 481.950 397.050 484.050 ;
        RECT 401.100 483.150 402.900 483.900 ;
        RECT 403.950 481.950 406.050 484.050 ;
        RECT 407.100 483.150 408.900 483.900 ;
        RECT 409.950 481.950 412.050 484.050 ;
        RECT 403.950 480.750 405.150 480.900 ;
        RECT 401.400 479.700 405.150 480.750 ;
        RECT 401.400 477.600 402.600 479.700 ;
        RECT 416.550 478.050 417.450 499.950 ;
        RECT 423.600 491.400 425.400 503.400 ;
        RECT 439.800 497.400 441.600 503.400 ;
        RECT 423.600 490.350 426.300 491.400 ;
        RECT 422.100 485.100 423.900 485.850 ;
        RECT 424.950 485.100 426.300 490.350 ;
        RECT 440.400 488.100 441.600 497.400 ;
        RECT 452.400 492.300 454.200 503.400 ;
        RECT 458.400 492.300 460.200 503.400 ;
        RECT 452.400 491.400 460.200 492.300 ;
        RECT 461.400 491.400 463.200 503.400 ;
        RECT 473.400 493.500 475.200 503.400 ;
        RECT 479.400 502.500 487.200 503.400 ;
        RECT 479.400 493.500 481.200 502.500 ;
        RECT 473.400 492.600 481.200 493.500 ;
        RECT 482.400 493.800 484.200 501.600 ;
        RECT 485.400 494.700 487.200 502.500 ;
        RECT 489.000 502.500 496.800 503.400 ;
        RECT 489.000 493.800 490.800 502.500 ;
        RECT 482.400 492.900 490.800 493.800 ;
        RECT 492.000 493.800 493.800 501.600 ;
        RECT 492.000 491.400 493.200 493.800 ;
        RECT 495.000 493.200 496.800 502.500 ;
        RECT 508.800 497.400 510.600 503.400 ;
        RECT 428.100 485.100 429.900 485.850 ;
        RECT 421.950 481.950 424.050 484.050 ;
        RECT 425.100 482.100 426.300 485.100 ;
        RECT 436.950 484.950 442.050 487.050 ;
        RECT 451.950 484.950 454.050 487.050 ;
        RECT 455.100 485.100 456.900 485.850 ;
        RECT 457.950 484.950 460.050 487.050 ;
        RECT 461.700 485.100 462.600 491.400 ;
        RECT 489.750 490.200 493.200 491.400 ;
        RECT 476.100 484.950 477.900 485.700 ;
        RECT 481.950 484.800 484.050 490.050 ;
        RECT 489.750 487.950 490.950 490.200 ;
        RECT 509.400 488.100 510.600 497.400 ;
        RECT 526.500 491.400 528.300 503.400 ;
        RECT 536.550 491.400 538.350 503.400 ;
        RECT 544.050 497.400 545.850 503.400 ;
        RECT 541.950 495.300 545.850 497.400 ;
        RECT 551.850 496.500 553.650 503.400 ;
        RECT 559.650 497.400 561.450 503.400 ;
        RECT 560.250 496.500 561.450 497.400 ;
        RECT 550.950 495.450 557.550 496.500 ;
        RECT 550.950 494.700 552.750 495.450 ;
        RECT 555.750 494.700 557.550 495.450 ;
        RECT 560.250 494.400 565.050 496.500 ;
        RECT 543.150 492.600 545.850 494.400 ;
        RECT 546.750 493.800 548.550 494.400 ;
        RECT 546.750 492.900 553.050 493.800 ;
        RECT 560.250 493.500 561.450 494.400 ;
        RECT 546.750 492.600 548.550 492.900 ;
        RECT 544.950 491.700 545.850 492.600 ;
        RECT 526.950 488.100 528.150 491.400 ;
        RECT 485.100 484.950 486.900 485.700 ;
        RECT 427.950 481.950 430.050 484.050 ;
        RECT 424.950 478.950 427.050 481.050 ;
        RECT 391.950 472.950 394.050 475.050 ;
        RECT 400.800 471.600 402.600 477.600 ;
        RECT 403.800 476.700 411.600 478.050 ;
        RECT 403.800 471.600 405.600 476.700 ;
        RECT 409.800 471.600 411.600 476.700 ;
        RECT 415.950 475.950 418.050 478.050 ;
        RECT 425.400 474.600 426.600 477.900 ;
        RECT 440.400 474.600 441.600 483.900 ;
        RECT 452.100 483.150 453.900 483.900 ;
        RECT 443.100 482.100 444.900 482.850 ;
        RECT 454.950 481.950 457.050 484.050 ;
        RECT 458.100 483.150 459.900 483.900 ;
        RECT 460.950 481.950 466.050 484.050 ;
        RECT 475.950 481.800 478.050 483.900 ;
        RECT 482.100 483.000 483.900 483.750 ;
        RECT 442.950 478.950 445.050 481.050 ;
        RECT 461.700 477.600 462.600 480.900 ;
        RECT 484.950 478.950 487.050 483.900 ;
        RECT 489.750 483.750 489.900 487.950 ;
        RECT 493.050 486.900 496.050 487.050 ;
        RECT 490.950 484.950 496.050 486.900 ;
        RECT 508.950 486.450 511.050 487.050 ;
        RECT 513.000 486.450 517.050 487.050 ;
        RECT 508.950 485.550 517.050 486.450 ;
        RECT 508.950 484.950 511.050 485.550 ;
        RECT 513.000 484.950 517.050 485.550 ;
        RECT 521.100 485.100 522.900 485.850 ;
        RECT 523.950 484.950 526.050 487.050 ;
        RECT 527.100 485.100 528.150 488.100 ;
        RECT 490.950 484.800 493.050 484.950 ;
        RECT 536.550 484.050 537.750 491.400 ;
        RECT 541.950 490.800 544.050 491.700 ;
        RECT 544.950 490.800 550.950 491.700 ;
        RECT 539.850 489.600 544.050 490.800 ;
        RECT 538.950 487.800 540.750 489.600 ;
        RECT 550.050 485.100 550.950 490.800 ;
        RECT 552.150 490.800 553.050 492.900 ;
        RECT 553.950 492.300 561.450 493.500 ;
        RECT 553.950 491.700 555.750 492.300 ;
        RECT 568.050 491.400 569.850 503.400 ;
        RECT 558.750 490.800 569.850 491.400 ;
        RECT 552.150 490.200 569.850 490.800 ;
        RECT 552.150 489.900 560.550 490.200 ;
        RECT 558.750 489.600 560.550 489.900 ;
        RECT 557.100 486.450 559.200 487.050 ;
        RECT 556.950 484.950 559.200 486.450 ;
        RECT 424.800 471.600 426.600 474.600 ;
        RECT 439.800 471.600 441.600 474.600 ;
        RECT 457.200 475.950 462.600 477.600 ;
        RECT 489.750 476.400 490.950 483.750 ;
        RECT 457.200 471.600 459.000 475.950 ;
        RECT 480.150 475.500 490.950 476.400 ;
        RECT 480.150 474.600 481.200 475.500 ;
        RECT 486.150 474.600 487.200 475.500 ;
        RECT 509.400 474.600 510.600 483.900 ;
        RECT 512.100 482.100 513.900 482.850 ;
        RECT 517.950 481.950 523.050 484.050 ;
        RECT 524.100 483.150 525.900 483.900 ;
        RECT 526.950 481.950 529.050 484.050 ;
        RECT 530.100 483.150 531.900 483.900 ;
        RECT 536.550 481.950 537.900 484.050 ;
        RECT 538.950 481.950 541.050 484.050 ;
        RECT 542.100 481.950 542.850 483.750 ;
        RECT 550.950 481.950 553.050 484.050 ;
        RECT 556.950 481.950 559.050 484.950 ;
        RECT 563.100 484.800 564.900 485.100 ;
        RECT 560.100 483.900 564.900 484.800 ;
        RECT 563.100 483.300 564.900 483.900 ;
        RECT 566.100 483.150 567.900 484.950 ;
        RECT 560.100 482.400 561.900 483.000 ;
        RECT 566.100 482.400 567.000 483.150 ;
        RECT 511.950 478.950 514.050 481.050 ;
        RECT 527.850 480.750 529.050 480.900 ;
        RECT 527.850 479.700 531.600 480.750 ;
        RECT 479.400 471.600 481.200 474.600 ;
        RECT 485.400 471.600 487.200 474.600 ;
        RECT 508.800 471.600 510.600 474.600 ;
        RECT 521.400 476.700 529.200 478.050 ;
        RECT 521.400 471.600 523.200 476.700 ;
        RECT 527.400 471.600 529.200 476.700 ;
        RECT 530.400 477.600 531.600 479.700 ;
        RECT 536.550 477.600 537.750 481.950 ;
        RECT 560.100 481.200 567.000 482.400 ;
        RECT 550.050 480.000 550.950 480.900 ;
        RECT 560.100 480.000 561.150 481.200 ;
        RECT 550.050 479.100 561.150 480.000 ;
        RECT 550.050 478.800 550.950 479.100 ;
        RECT 530.400 471.600 532.200 477.600 ;
        RECT 536.550 471.600 538.350 477.600 ;
        RECT 541.950 476.700 544.050 477.600 ;
        RECT 549.150 477.000 550.950 478.800 ;
        RECT 560.100 478.200 561.150 479.100 ;
        RECT 556.350 477.450 558.150 478.200 ;
        RECT 541.950 475.500 545.700 476.700 ;
        RECT 544.650 474.600 545.700 475.500 ;
        RECT 553.200 476.400 558.150 477.450 ;
        RECT 559.650 476.400 561.450 478.200 ;
        RECT 568.950 477.600 569.850 490.200 ;
        RECT 553.200 474.600 554.250 476.400 ;
        RECT 562.950 475.500 565.050 477.600 ;
        RECT 562.950 474.600 564.000 475.500 ;
        RECT 544.650 471.600 546.450 474.600 ;
        RECT 552.450 471.600 554.250 474.600 ;
        RECT 560.250 473.700 564.000 474.600 ;
        RECT 560.250 471.600 562.050 473.700 ;
        RECT 568.050 471.600 569.850 477.600 ;
        RECT 572.550 491.400 574.350 503.400 ;
        RECT 580.050 497.400 581.850 503.400 ;
        RECT 577.950 495.300 581.850 497.400 ;
        RECT 587.850 496.500 589.650 503.400 ;
        RECT 595.650 497.400 597.450 503.400 ;
        RECT 596.250 496.500 597.450 497.400 ;
        RECT 586.950 495.450 593.550 496.500 ;
        RECT 586.950 494.700 588.750 495.450 ;
        RECT 591.750 494.700 593.550 495.450 ;
        RECT 596.250 494.400 601.050 496.500 ;
        RECT 579.150 492.600 581.850 494.400 ;
        RECT 582.750 493.800 584.550 494.400 ;
        RECT 582.750 492.900 589.050 493.800 ;
        RECT 596.250 493.500 597.450 494.400 ;
        RECT 582.750 492.600 584.550 492.900 ;
        RECT 580.950 491.700 581.850 492.600 ;
        RECT 572.550 484.050 573.750 491.400 ;
        RECT 577.950 490.800 580.050 491.700 ;
        RECT 580.950 490.800 586.950 491.700 ;
        RECT 575.850 489.600 580.050 490.800 ;
        RECT 574.950 487.800 576.750 489.600 ;
        RECT 586.050 485.100 586.950 490.800 ;
        RECT 588.150 490.800 589.050 492.900 ;
        RECT 589.950 492.300 597.450 493.500 ;
        RECT 589.950 491.700 591.750 492.300 ;
        RECT 604.050 491.400 605.850 503.400 ;
        RECT 619.800 497.400 621.600 503.400 ;
        RECT 594.750 490.800 605.850 491.400 ;
        RECT 588.150 490.200 605.850 490.800 ;
        RECT 588.150 489.900 596.550 490.200 ;
        RECT 594.750 489.600 596.550 489.900 ;
        RECT 572.550 481.950 573.900 484.050 ;
        RECT 574.950 481.950 577.050 484.050 ;
        RECT 578.100 481.950 578.850 483.750 ;
        RECT 586.950 481.950 589.050 484.050 ;
        RECT 592.950 481.950 595.050 487.050 ;
        RECT 599.100 484.800 600.900 485.100 ;
        RECT 596.100 483.900 600.900 484.800 ;
        RECT 599.100 483.300 600.900 483.900 ;
        RECT 602.100 483.150 603.900 484.950 ;
        RECT 596.100 482.400 597.900 483.000 ;
        RECT 602.100 482.400 603.000 483.150 ;
        RECT 572.550 477.600 573.750 481.950 ;
        RECT 596.100 481.200 603.000 482.400 ;
        RECT 586.050 480.000 586.950 480.900 ;
        RECT 596.100 480.000 597.150 481.200 ;
        RECT 586.050 479.100 597.150 480.000 ;
        RECT 586.050 478.800 586.950 479.100 ;
        RECT 572.550 471.600 574.350 477.600 ;
        RECT 577.950 476.700 580.050 477.600 ;
        RECT 585.150 477.000 586.950 478.800 ;
        RECT 596.100 478.200 597.150 479.100 ;
        RECT 592.350 477.450 594.150 478.200 ;
        RECT 577.950 475.500 581.700 476.700 ;
        RECT 580.650 474.600 581.700 475.500 ;
        RECT 589.200 476.400 594.150 477.450 ;
        RECT 595.650 476.400 597.450 478.200 ;
        RECT 604.950 477.600 605.850 490.200 ;
        RECT 616.950 487.950 619.050 490.050 ;
        RECT 620.400 488.100 621.600 497.400 ;
        RECT 638.700 491.400 640.500 503.400 ;
        RECT 656.400 497.400 658.200 503.400 ;
        RECT 670.800 497.400 672.600 503.400 ;
        RECT 688.800 497.400 690.600 503.400 ;
        RECT 706.800 497.400 708.600 503.400 ;
        RECT 622.950 487.950 625.050 490.050 ;
        RECT 638.850 488.100 640.050 491.400 ;
        RECT 656.400 488.100 657.600 497.400 ;
        RECT 671.400 488.100 672.600 497.400 ;
        RECT 689.400 488.100 690.600 497.400 ;
        RECT 698.100 493.950 700.200 496.050 ;
        RECT 698.550 490.050 699.450 493.950 ;
        RECT 617.100 486.150 618.900 486.900 ;
        RECT 619.950 484.950 622.050 487.050 ;
        RECT 623.100 486.150 624.900 486.900 ;
        RECT 634.800 484.950 637.050 487.050 ;
        RECT 638.850 485.100 639.900 488.100 ;
        RECT 691.950 487.950 694.050 490.050 ;
        RECT 697.950 487.950 700.050 490.050 ;
        RECT 707.400 488.100 708.600 497.400 ;
        RECT 719.400 492.600 721.200 503.400 ;
        RECT 725.400 502.500 733.200 503.400 ;
        RECT 725.400 492.600 727.200 502.500 ;
        RECT 719.400 491.700 727.200 492.600 ;
        RECT 728.400 490.500 730.200 501.600 ;
        RECT 731.400 491.400 733.200 502.500 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 749.700 491.400 751.500 503.400 ;
        RECT 766.800 497.400 768.600 503.400 ;
        RECT 709.950 487.950 712.050 490.050 ;
        RECT 726.150 489.600 730.200 490.500 ;
        RECT 726.150 488.100 727.050 489.600 ;
        RECT 640.950 484.950 643.050 487.050 ;
        RECT 644.100 485.100 645.900 485.850 ;
        RECT 655.950 484.950 658.050 487.050 ;
        RECT 670.950 484.950 673.050 487.050 ;
        RECT 686.100 486.150 687.900 486.900 ;
        RECT 688.950 484.950 691.050 487.050 ;
        RECT 692.100 486.150 693.900 486.900 ;
        RECT 704.100 486.150 705.900 486.900 ;
        RECT 706.950 484.950 709.050 487.050 ;
        RECT 710.100 486.150 711.900 486.900 ;
        RECT 719.250 485.100 720.900 485.850 ;
        RECT 721.950 484.950 724.050 487.050 ;
        RECT 726.150 485.100 726.900 488.100 ;
        RECT 727.950 484.950 730.050 487.050 ;
        RECT 731.100 485.100 732.900 485.850 ;
        RECT 737.550 484.050 738.450 490.950 ;
        RECT 749.850 488.100 751.050 491.400 ;
        RECT 760.950 490.950 763.050 493.050 ;
        RECT 745.950 484.950 748.050 487.050 ;
        RECT 749.850 485.100 750.900 488.100 ;
        RECT 751.950 484.950 754.050 487.050 ;
        RECT 761.550 486.450 762.450 490.950 ;
        RECT 767.400 488.100 768.600 497.400 ;
        RECT 783.600 491.400 785.400 503.400 ;
        RECT 802.500 491.400 804.300 503.400 ;
        RECT 824.700 491.400 826.500 503.400 ;
        RECT 843.600 491.400 845.400 503.400 ;
        RECT 783.600 490.350 786.300 491.400 ;
        RECT 766.950 486.450 769.050 487.050 ;
        RECT 755.100 485.100 756.900 485.850 ;
        RECT 761.550 485.550 769.050 486.450 ;
        RECT 766.950 484.950 769.050 485.550 ;
        RECT 782.100 485.100 783.900 485.850 ;
        RECT 784.950 485.100 786.300 490.350 ;
        RECT 802.950 488.100 804.150 491.400 ;
        RECT 788.100 485.100 789.900 485.850 ;
        RECT 797.100 485.100 798.900 485.850 ;
        RECT 620.400 479.700 621.600 483.900 ;
        RECT 635.100 483.150 636.900 483.900 ;
        RECT 637.950 481.950 640.050 484.050 ;
        RECT 641.100 483.150 642.900 483.900 ;
        RECT 643.950 481.950 646.050 484.050 ;
        RECT 653.100 482.100 654.900 482.850 ;
        RECT 637.950 480.750 639.150 480.900 ;
        RECT 589.200 474.600 590.250 476.400 ;
        RECT 598.950 475.500 601.050 477.600 ;
        RECT 598.950 474.600 600.000 475.500 ;
        RECT 580.650 471.600 582.450 474.600 ;
        RECT 588.450 471.600 590.250 474.600 ;
        RECT 596.250 473.700 600.000 474.600 ;
        RECT 596.250 471.600 598.050 473.700 ;
        RECT 604.050 471.600 605.850 477.600 ;
        RECT 618.000 478.800 621.600 479.700 ;
        RECT 635.400 479.700 639.150 480.750 ;
        RECT 618.000 471.600 619.800 478.800 ;
        RECT 635.400 477.600 636.600 479.700 ;
        RECT 634.800 471.600 636.600 477.600 ;
        RECT 637.800 476.700 645.600 478.050 ;
        RECT 637.800 471.600 639.600 476.700 ;
        RECT 643.800 471.600 645.600 476.700 ;
        RECT 656.400 474.600 657.600 483.900 ;
        RECT 671.400 474.600 672.600 483.900 ;
        RECT 674.100 482.100 675.900 482.850 ;
        RECT 689.400 479.700 690.600 483.900 ;
        RECT 707.400 479.700 708.600 483.900 ;
        RECT 718.950 481.950 721.050 484.050 ;
        RECT 722.250 483.150 723.900 483.900 ;
        RECT 724.950 481.950 727.050 484.050 ;
        RECT 728.100 483.150 729.750 483.900 ;
        RECT 730.950 481.950 733.050 484.050 ;
        RECT 736.950 481.950 739.050 484.050 ;
        RECT 746.100 483.150 747.900 483.900 ;
        RECT 748.950 481.950 751.050 484.050 ;
        RECT 752.100 483.150 753.900 483.900 ;
        RECT 754.950 481.950 757.050 484.050 ;
        RECT 656.400 471.600 658.200 474.600 ;
        RECT 670.800 471.600 672.600 474.600 ;
        RECT 687.000 478.800 690.600 479.700 ;
        RECT 705.000 478.800 708.600 479.700 ;
        RECT 687.000 471.600 688.800 478.800 ;
        RECT 705.000 471.600 706.800 478.800 ;
        RECT 724.950 477.600 726.000 480.900 ;
        RECT 748.950 480.750 750.150 480.900 ;
        RECT 746.400 479.700 750.150 480.750 ;
        RECT 746.400 477.600 747.600 479.700 ;
        RECT 724.200 471.600 726.000 477.600 ;
        RECT 745.800 471.600 747.600 477.600 ;
        RECT 748.800 476.700 756.600 478.050 ;
        RECT 748.800 471.600 750.600 476.700 ;
        RECT 754.800 471.600 756.600 476.700 ;
        RECT 767.400 474.600 768.600 483.900 ;
        RECT 770.100 482.100 771.900 482.850 ;
        RECT 781.950 481.950 784.050 484.050 ;
        RECT 785.100 482.100 786.300 485.100 ;
        RECT 799.950 484.950 802.050 487.050 ;
        RECT 803.100 485.100 804.150 488.100 ;
        RECT 824.850 488.100 826.050 491.400 ;
        RECT 843.600 490.350 846.300 491.400 ;
        RECT 805.950 484.950 808.050 487.050 ;
        RECT 820.950 484.950 823.050 487.050 ;
        RECT 824.850 485.100 825.900 488.100 ;
        RECT 826.950 484.950 829.050 487.050 ;
        RECT 830.100 485.100 831.900 485.850 ;
        RECT 842.100 485.100 843.900 485.850 ;
        RECT 844.950 485.100 846.300 490.350 ;
        RECT 848.100 485.100 849.900 485.850 ;
        RECT 787.950 481.950 790.050 484.050 ;
        RECT 796.950 481.950 799.050 484.050 ;
        RECT 800.100 483.150 801.900 483.900 ;
        RECT 802.950 481.950 805.050 484.050 ;
        RECT 806.100 483.150 807.900 483.900 ;
        RECT 821.100 483.150 822.900 483.900 ;
        RECT 823.950 481.950 826.050 484.050 ;
        RECT 827.100 483.150 828.900 483.900 ;
        RECT 841.950 481.950 844.200 484.050 ;
        RECT 845.100 482.100 846.300 485.100 ;
        RECT 769.950 478.950 772.050 481.050 ;
        RECT 784.950 478.950 787.050 481.050 ;
        RECT 803.850 480.750 805.050 480.900 ;
        RECT 823.950 480.750 825.150 480.900 ;
        RECT 803.850 479.700 807.600 480.750 ;
        RECT 785.400 474.600 786.600 477.900 ;
        RECT 766.800 471.600 768.600 474.600 ;
        RECT 784.800 471.600 786.600 474.600 ;
        RECT 797.400 476.700 805.200 478.050 ;
        RECT 797.400 471.600 799.200 476.700 ;
        RECT 803.400 471.600 805.200 476.700 ;
        RECT 806.400 477.600 807.600 479.700 ;
        RECT 821.400 479.700 825.150 480.750 ;
        RECT 821.400 477.600 822.600 479.700 ;
        RECT 844.950 478.950 847.050 481.050 ;
        RECT 806.400 471.600 808.200 477.600 ;
        RECT 820.800 471.600 822.600 477.600 ;
        RECT 823.800 476.700 831.600 478.050 ;
        RECT 823.800 471.600 825.600 476.700 ;
        RECT 829.800 471.600 831.600 476.700 ;
        RECT 845.400 474.600 846.600 477.900 ;
        RECT 844.800 471.600 846.600 474.600 ;
        RECT 12.300 463.200 14.100 467.400 ;
        RECT 12.150 461.400 14.100 463.200 ;
        RECT 12.150 458.100 13.050 461.400 ;
        RECT 14.100 459.900 15.900 460.500 ;
        RECT 19.800 459.900 21.600 467.400 ;
        RECT 34.200 460.200 36.000 467.400 ;
        RECT 40.950 463.950 43.050 466.050 ;
        RECT 14.100 458.700 21.600 459.900 ;
        RECT 32.400 459.300 36.000 460.200 ;
        RECT 10.950 456.450 13.050 457.050 ;
        RECT 5.550 455.550 13.050 456.450 ;
        RECT 5.550 439.050 6.450 455.550 ;
        RECT 10.950 454.950 13.050 455.550 ;
        RECT 14.100 455.100 15.900 455.850 ;
        RECT 10.950 447.600 12.000 453.900 ;
        RECT 13.950 451.950 16.050 454.050 ;
        RECT 4.950 436.950 7.050 439.050 ;
        RECT 10.200 435.600 12.000 447.600 ;
        RECT 17.550 441.600 18.600 458.700 ;
        RECT 19.950 454.950 22.050 457.050 ;
        RECT 32.400 455.100 33.600 459.300 ;
        RECT 20.100 453.150 21.900 453.900 ;
        RECT 29.100 452.100 30.900 452.850 ;
        RECT 31.950 451.950 34.050 454.050 ;
        RECT 35.100 452.100 36.900 452.850 ;
        RECT 41.550 451.050 42.450 463.950 ;
        RECT 43.950 457.950 46.050 460.050 ;
        RECT 53.100 459.000 54.900 467.400 ;
        RECT 75.000 463.050 76.800 467.400 ;
        RECT 28.950 448.950 31.050 451.050 ;
        RECT 16.800 435.600 18.600 441.600 ;
        RECT 32.400 441.600 33.600 450.900 ;
        RECT 34.950 448.950 37.050 451.050 ;
        RECT 40.800 448.950 42.900 451.050 ;
        RECT 44.550 442.050 45.450 457.950 ;
        RECT 50.700 457.350 54.900 459.000 ;
        RECT 71.400 461.400 76.800 463.050 ;
        RECT 71.400 458.100 72.300 461.400 ;
        RECT 95.100 459.000 96.900 467.400 ;
        RECT 113.400 464.400 115.200 467.400 ;
        RECT 92.700 457.350 96.900 459.000 ;
        RECT 109.950 457.950 112.050 460.050 ;
        RECT 50.700 452.100 51.600 457.350 ;
        RECT 53.100 455.100 54.900 455.850 ;
        RECT 59.100 455.100 60.900 455.850 ;
        RECT 67.950 454.950 73.050 457.050 ;
        RECT 74.100 455.100 75.900 455.850 ;
        RECT 76.800 454.950 79.050 457.050 ;
        RECT 80.100 455.100 81.900 455.850 ;
        RECT 52.950 451.950 55.050 454.050 ;
        RECT 58.950 451.950 61.050 454.050 ;
        RECT 46.950 448.950 52.050 451.050 ;
        RECT 55.950 448.950 58.050 451.050 ;
        RECT 50.700 442.800 51.600 447.900 ;
        RECT 56.100 447.150 57.900 447.900 ;
        RECT 71.400 447.600 72.300 453.900 ;
        RECT 73.950 451.950 76.050 454.050 ;
        RECT 77.100 453.150 78.900 453.900 ;
        RECT 79.950 451.950 82.050 454.050 ;
        RECT 92.700 452.100 93.600 457.350 ;
        RECT 110.100 456.150 111.900 456.900 ;
        RECT 95.100 455.100 96.900 455.850 ;
        RECT 101.100 455.100 102.900 455.850 ;
        RECT 113.400 455.100 114.600 464.400 ;
        RECT 127.800 461.400 129.600 467.400 ;
        RECT 128.400 459.300 129.600 461.400 ;
        RECT 130.800 462.300 132.600 467.400 ;
        RECT 136.800 462.300 138.600 467.400 ;
        RECT 151.800 464.400 153.600 467.400 ;
        RECT 130.800 460.950 138.600 462.300 ;
        RECT 152.400 461.100 153.600 464.400 ;
        RECT 169.200 460.200 171.000 467.400 ;
        RECT 128.400 458.250 132.150 459.300 ;
        RECT 130.950 458.100 132.150 458.250 ;
        RECT 151.800 457.950 154.050 460.050 ;
        RECT 167.400 459.300 171.000 460.200 ;
        RECT 128.100 455.100 129.900 455.850 ;
        RECT 130.800 454.950 133.050 457.050 ;
        RECT 134.100 455.100 135.900 455.850 ;
        RECT 136.950 454.950 139.050 457.050 ;
        RECT 148.950 454.950 151.050 457.050 ;
        RECT 94.950 451.950 97.050 454.050 ;
        RECT 100.950 451.950 103.050 454.050 ;
        RECT 109.950 451.950 115.050 454.050 ;
        RECT 127.800 451.950 130.050 454.050 ;
        RECT 91.950 450.450 94.050 451.050 ;
        RECT 86.550 449.550 94.050 450.450 ;
        RECT 32.400 435.600 34.200 441.600 ;
        RECT 43.950 439.950 46.050 442.050 ;
        RECT 50.700 441.900 57.300 442.800 ;
        RECT 50.700 441.600 51.600 441.900 ;
        RECT 49.800 435.600 51.600 441.600 ;
        RECT 55.800 441.600 57.300 441.900 ;
        RECT 55.800 435.600 57.600 441.600 ;
        RECT 70.800 435.600 72.600 447.600 ;
        RECT 73.800 446.700 81.600 447.600 ;
        RECT 73.800 435.600 75.600 446.700 ;
        RECT 79.800 435.600 81.600 446.700 ;
        RECT 86.550 445.050 87.450 449.550 ;
        RECT 91.950 448.950 94.050 449.550 ;
        RECT 97.950 448.950 100.050 451.050 ;
        RECT 131.850 450.900 132.900 453.900 ;
        RECT 133.950 451.950 136.050 454.050 ;
        RECT 152.100 453.900 153.300 456.900 ;
        RECT 154.950 454.950 157.050 457.050 ;
        RECT 167.400 455.100 168.600 459.300 ;
        RECT 188.100 459.000 189.900 467.400 ;
        RECT 208.200 460.200 210.000 467.400 ;
        RECT 226.200 461.400 228.000 467.400 ;
        RECT 247.500 461.400 249.300 467.400 ;
        RECT 253.800 464.400 255.600 467.400 ;
        RECT 185.700 457.350 189.900 459.000 ;
        RECT 206.400 459.300 210.000 460.200 ;
        RECT 137.100 453.150 138.900 453.900 ;
        RECT 149.100 453.150 150.900 453.900 ;
        RECT 85.950 442.950 88.050 445.050 ;
        RECT 92.700 442.800 93.600 447.900 ;
        RECT 98.100 447.150 99.900 447.900 ;
        RECT 92.700 441.900 99.300 442.800 ;
        RECT 92.700 441.600 93.600 441.900 ;
        RECT 91.800 435.600 93.600 441.600 ;
        RECT 97.800 441.600 99.300 441.900 ;
        RECT 113.400 441.600 114.600 450.900 ;
        RECT 131.850 447.600 133.050 450.900 ;
        RECT 151.950 448.650 153.300 453.900 ;
        RECT 155.100 453.150 156.900 453.900 ;
        RECT 164.100 452.100 165.900 452.850 ;
        RECT 166.950 451.950 169.050 454.050 ;
        RECT 170.100 452.100 171.900 452.850 ;
        RECT 185.700 452.100 186.600 457.350 ;
        RECT 188.100 455.100 189.900 455.850 ;
        RECT 194.100 455.100 195.900 455.850 ;
        RECT 206.400 455.100 207.600 459.300 ;
        RECT 226.950 458.100 228.000 461.400 ;
        RECT 247.800 458.100 249.000 461.400 ;
        RECT 253.800 460.500 255.000 464.400 ;
        RECT 259.950 463.950 262.050 466.050 ;
        RECT 249.900 459.600 255.000 460.500 ;
        RECT 249.900 458.700 251.850 459.600 ;
        RECT 250.950 458.100 251.850 458.700 ;
        RECT 214.950 454.950 217.050 457.050 ;
        RECT 220.950 454.950 223.050 457.050 ;
        RECT 224.250 455.100 225.900 455.850 ;
        RECT 226.950 454.950 229.050 457.050 ;
        RECT 230.100 455.100 231.750 455.850 ;
        RECT 232.950 454.950 235.050 457.050 ;
        RECT 247.950 456.450 250.050 457.050 ;
        RECT 242.550 455.550 250.050 456.450 ;
        RECT 187.950 451.950 190.050 454.050 ;
        RECT 193.950 451.950 196.050 454.050 ;
        RECT 203.100 452.100 204.900 452.850 ;
        RECT 205.950 451.950 208.050 454.050 ;
        RECT 209.100 452.100 210.900 452.850 ;
        RECT 163.950 448.950 166.050 451.050 ;
        RECT 150.600 447.600 153.300 448.650 ;
        RECT 97.800 435.600 99.600 441.600 ;
        RECT 113.400 435.600 115.200 441.600 ;
        RECT 131.700 435.600 133.500 447.600 ;
        RECT 150.600 435.600 152.400 447.600 ;
        RECT 167.400 441.600 168.600 450.900 ;
        RECT 169.950 448.950 172.050 451.050 ;
        RECT 184.950 450.450 187.050 451.050 ;
        RECT 179.550 449.550 187.050 450.450 ;
        RECT 179.550 445.050 180.450 449.550 ;
        RECT 184.950 448.950 187.050 449.550 ;
        RECT 190.950 448.950 193.050 451.050 ;
        RECT 202.950 448.950 205.050 451.050 ;
        RECT 178.950 442.950 181.050 445.050 ;
        RECT 185.700 442.800 186.600 447.900 ;
        RECT 191.100 447.150 192.900 447.900 ;
        RECT 185.700 441.900 192.300 442.800 ;
        RECT 185.700 441.600 186.600 441.900 ;
        RECT 167.400 435.600 169.200 441.600 ;
        RECT 184.800 435.600 186.600 441.600 ;
        RECT 190.800 441.600 192.300 441.900 ;
        RECT 206.400 441.600 207.600 450.900 ;
        RECT 208.950 448.950 211.050 451.050 ;
        RECT 215.550 445.050 216.450 454.950 ;
        RECT 221.250 453.150 222.900 453.900 ;
        RECT 223.800 451.950 226.050 454.050 ;
        RECT 228.150 450.900 228.900 453.900 ;
        RECT 229.950 451.950 232.050 454.050 ;
        RECT 233.100 453.150 234.900 453.900 ;
        RECT 228.150 449.400 229.050 450.900 ;
        RECT 228.150 448.500 232.200 449.400 ;
        RECT 221.400 446.400 229.200 447.300 ;
        RECT 214.950 442.950 217.050 445.050 ;
        RECT 190.800 435.600 192.600 441.600 ;
        RECT 206.400 435.600 208.200 441.600 ;
        RECT 221.400 435.600 223.200 446.400 ;
        RECT 227.400 436.500 229.200 446.400 ;
        RECT 230.400 437.400 232.200 448.500 ;
        RECT 233.400 436.500 235.200 447.600 ;
        RECT 242.550 445.050 243.450 455.550 ;
        RECT 247.950 454.950 250.050 455.550 ;
        RECT 251.100 453.900 251.850 458.100 ;
        RECT 253.950 454.950 256.050 457.050 ;
        RECT 247.800 447.600 249.000 453.900 ;
        RECT 250.950 450.300 251.850 453.900 ;
        RECT 254.100 453.150 255.900 453.900 ;
        RECT 249.900 449.400 251.850 450.300 ;
        RECT 260.550 450.450 261.450 463.950 ;
        RECT 269.100 459.000 270.900 467.400 ;
        RECT 284.400 462.300 286.200 467.400 ;
        RECT 290.400 462.300 292.200 467.400 ;
        RECT 284.400 460.950 292.200 462.300 ;
        RECT 293.400 461.400 295.200 467.400 ;
        RECT 293.400 459.300 294.600 461.400 ;
        RECT 302.100 460.950 304.200 463.050 ;
        RECT 307.800 461.400 309.600 467.400 ;
        RECT 266.700 457.350 270.900 459.000 ;
        RECT 290.850 458.250 294.600 459.300 ;
        RECT 290.850 458.100 292.050 458.250 ;
        RECT 266.700 452.100 267.600 457.350 ;
        RECT 269.100 455.100 270.900 455.850 ;
        RECT 275.100 455.100 276.900 455.850 ;
        RECT 283.950 454.950 286.050 457.050 ;
        RECT 287.100 455.100 288.900 455.850 ;
        RECT 289.950 454.950 292.050 457.050 ;
        RECT 293.100 455.100 294.900 455.850 ;
        RECT 298.950 454.950 301.050 457.050 ;
        RECT 268.950 451.950 271.050 454.050 ;
        RECT 274.950 451.950 277.050 454.050 ;
        RECT 284.100 453.150 285.900 453.900 ;
        RECT 286.950 451.950 289.050 454.050 ;
        RECT 265.950 450.450 268.050 451.050 ;
        RECT 260.550 449.550 268.050 450.450 ;
        RECT 249.900 448.500 255.600 449.400 ;
        RECT 265.950 448.950 268.050 449.550 ;
        RECT 271.950 448.950 274.050 451.050 ;
        RECT 290.100 450.900 291.150 453.900 ;
        RECT 292.950 451.950 295.050 454.050 ;
        RECT 241.950 442.950 244.050 445.050 ;
        RECT 227.400 435.600 235.200 436.500 ;
        RECT 247.500 435.600 249.300 447.600 ;
        RECT 254.400 441.600 255.600 448.500 ;
        RECT 266.700 442.800 267.600 447.900 ;
        RECT 272.100 447.150 273.900 447.900 ;
        RECT 289.950 447.600 291.150 450.900 ;
        RECT 266.700 441.900 273.300 442.800 ;
        RECT 266.700 441.600 267.600 441.900 ;
        RECT 253.800 435.600 255.600 441.600 ;
        RECT 265.800 435.600 267.600 441.600 ;
        RECT 271.800 441.600 273.300 441.900 ;
        RECT 271.800 435.600 273.600 441.600 ;
        RECT 289.500 435.600 291.300 447.600 ;
        RECT 293.550 445.050 294.450 451.950 ;
        RECT 299.550 451.050 300.450 454.950 ;
        RECT 298.950 448.950 301.050 451.050 ;
        RECT 302.550 445.050 303.450 460.950 ;
        RECT 308.400 459.300 309.600 461.400 ;
        RECT 310.800 462.300 312.600 467.400 ;
        RECT 316.800 462.300 318.600 467.400 ;
        RECT 310.800 460.950 318.600 462.300 ;
        RECT 326.400 459.900 328.200 467.400 ;
        RECT 333.900 463.200 335.700 467.400 ;
        RECT 340.950 463.950 343.050 466.050 ;
        RECT 333.900 461.400 335.850 463.200 ;
        RECT 332.100 459.900 333.900 460.500 ;
        RECT 308.400 458.250 312.150 459.300 ;
        RECT 326.400 458.700 333.900 459.900 ;
        RECT 310.950 458.100 312.150 458.250 ;
        RECT 308.100 455.100 309.900 455.850 ;
        RECT 310.950 454.950 313.200 457.050 ;
        RECT 314.100 455.100 315.900 455.850 ;
        RECT 316.950 454.950 319.200 457.050 ;
        RECT 325.950 454.950 328.050 457.050 ;
        RECT 307.800 451.950 310.050 454.050 ;
        RECT 311.850 450.900 312.900 453.900 ;
        RECT 313.950 451.950 316.050 454.050 ;
        RECT 317.100 453.150 318.900 453.900 ;
        RECT 326.100 453.150 327.900 453.900 ;
        RECT 311.850 447.600 313.050 450.900 ;
        RECT 292.950 442.950 295.050 445.050 ;
        RECT 301.950 442.950 304.050 445.050 ;
        RECT 311.700 435.600 313.500 447.600 ;
        RECT 329.400 441.600 330.450 458.700 ;
        RECT 334.950 458.100 335.850 461.400 ;
        RECT 334.950 456.450 337.050 457.050 ;
        RECT 341.550 456.450 342.450 463.950 ;
        RECT 347.400 459.900 349.200 467.400 ;
        RECT 354.900 463.200 356.700 467.400 ;
        RECT 361.800 463.950 363.900 466.050 ;
        RECT 365.100 463.950 367.200 466.050 ;
        RECT 354.900 461.400 356.850 463.200 ;
        RECT 353.100 459.900 354.900 460.500 ;
        RECT 347.400 458.700 354.900 459.900 ;
        RECT 332.100 455.100 333.900 455.850 ;
        RECT 334.950 455.550 342.450 456.450 ;
        RECT 334.950 454.950 337.050 455.550 ;
        RECT 346.950 454.950 349.050 457.050 ;
        RECT 331.950 451.950 334.050 454.050 ;
        RECT 336.000 447.600 337.050 453.900 ;
        RECT 347.100 453.150 348.900 453.900 ;
        RECT 329.400 435.600 331.200 441.600 ;
        RECT 336.000 435.600 337.800 447.600 ;
        RECT 350.400 441.600 351.450 458.700 ;
        RECT 355.950 458.100 356.850 461.400 ;
        RECT 362.550 460.050 363.450 463.950 ;
        RECT 361.950 457.950 364.050 460.050 ;
        RECT 353.100 455.100 354.900 455.850 ;
        RECT 355.950 454.950 358.200 457.050 ;
        RECT 352.950 451.950 355.050 454.050 ;
        RECT 357.000 447.600 358.050 453.900 ;
        RECT 350.400 435.600 352.200 441.600 ;
        RECT 357.000 435.600 358.800 447.600 ;
        RECT 365.550 445.050 366.450 463.950 ;
        RECT 372.000 460.200 373.800 467.400 ;
        RECT 388.800 461.400 390.600 467.400 ;
        RECT 372.000 459.300 375.600 460.200 ;
        RECT 374.400 455.100 375.600 459.300 ;
        RECT 382.950 457.950 385.050 460.050 ;
        RECT 389.400 459.300 390.600 461.400 ;
        RECT 391.800 462.300 393.600 467.400 ;
        RECT 397.800 462.300 399.600 467.400 ;
        RECT 391.800 460.950 399.600 462.300 ;
        RECT 407.400 462.300 409.200 467.400 ;
        RECT 413.400 462.300 415.200 467.400 ;
        RECT 407.400 460.950 415.200 462.300 ;
        RECT 416.400 461.400 418.200 467.400 ;
        RECT 416.400 459.300 417.600 461.400 ;
        RECT 421.950 460.950 424.050 463.050 ;
        RECT 428.400 462.300 430.200 467.400 ;
        RECT 434.400 462.300 436.200 467.400 ;
        RECT 428.400 460.950 436.200 462.300 ;
        RECT 437.400 461.400 439.200 467.400 ;
        RECT 451.800 464.400 453.600 467.400 ;
        RECT 389.400 458.250 393.150 459.300 ;
        RECT 391.950 458.100 393.150 458.250 ;
        RECT 413.850 458.250 417.600 459.300 ;
        RECT 413.850 458.100 415.050 458.250 ;
        RECT 371.100 452.100 372.900 452.850 ;
        RECT 373.950 451.950 376.050 454.050 ;
        RECT 377.100 452.100 378.900 452.850 ;
        RECT 383.550 451.050 384.450 457.950 ;
        RECT 389.100 455.100 390.900 455.850 ;
        RECT 391.800 454.950 394.050 457.050 ;
        RECT 395.100 455.100 396.900 455.850 ;
        RECT 397.950 454.950 400.050 457.050 ;
        RECT 406.950 454.950 409.050 457.050 ;
        RECT 410.100 455.100 411.900 455.850 ;
        RECT 412.950 454.950 415.050 457.050 ;
        RECT 416.100 455.100 417.900 455.850 ;
        RECT 422.550 454.050 423.450 460.950 ;
        RECT 437.400 459.300 438.600 461.400 ;
        RECT 445.950 460.950 448.050 463.050 ;
        RECT 434.850 458.250 438.600 459.300 ;
        RECT 434.850 458.100 436.050 458.250 ;
        RECT 427.950 454.950 430.050 457.050 ;
        RECT 431.100 455.100 432.900 455.850 ;
        RECT 433.950 454.950 436.050 457.050 ;
        RECT 437.100 455.100 438.900 455.850 ;
        RECT 388.950 451.950 391.050 454.050 ;
        RECT 370.950 448.950 373.050 451.050 ;
        RECT 364.950 442.950 367.050 445.050 ;
        RECT 374.400 441.600 375.600 450.900 ;
        RECT 376.950 448.950 379.050 451.050 ;
        RECT 382.950 448.950 385.050 451.050 ;
        RECT 392.850 450.900 393.900 453.900 ;
        RECT 394.950 451.950 397.050 454.050 ;
        RECT 398.100 453.150 399.900 453.900 ;
        RECT 407.100 453.150 408.900 453.900 ;
        RECT 409.950 451.950 412.050 454.050 ;
        RECT 413.100 450.900 414.150 453.900 ;
        RECT 421.950 451.950 424.050 454.050 ;
        RECT 428.100 453.150 429.900 453.900 ;
        RECT 430.950 451.950 433.050 454.050 ;
        RECT 434.100 450.900 435.150 453.900 ;
        RECT 392.850 447.600 394.050 450.900 ;
        RECT 412.950 447.600 414.150 450.900 ;
        RECT 433.950 447.600 435.150 450.900 ;
        RECT 373.800 435.600 375.600 441.600 ;
        RECT 392.700 435.600 394.500 447.600 ;
        RECT 412.500 435.600 414.300 447.600 ;
        RECT 433.500 435.600 435.300 447.600 ;
        RECT 446.550 439.050 447.450 460.950 ;
        RECT 452.400 455.100 453.600 464.400 ;
        RECT 464.400 462.300 466.200 467.400 ;
        RECT 470.400 462.300 472.200 467.400 ;
        RECT 464.400 460.950 472.200 462.300 ;
        RECT 473.400 461.400 475.200 467.400 ;
        RECT 485.400 462.300 487.200 467.400 ;
        RECT 491.400 462.300 493.200 467.400 ;
        RECT 454.950 457.950 457.050 460.050 ;
        RECT 473.400 459.300 474.600 461.400 ;
        RECT 485.400 460.950 493.200 462.300 ;
        RECT 494.400 461.400 496.200 467.400 ;
        RECT 506.400 462.300 508.200 467.400 ;
        RECT 512.400 462.300 514.200 467.400 ;
        RECT 494.400 459.300 495.600 461.400 ;
        RECT 506.400 460.950 514.200 462.300 ;
        RECT 515.400 461.400 517.200 467.400 ;
        RECT 529.500 461.400 531.300 467.400 ;
        RECT 535.800 464.400 537.600 467.400 ;
        RECT 515.400 459.300 516.600 461.400 ;
        RECT 470.850 458.250 474.600 459.300 ;
        RECT 491.850 458.250 495.600 459.300 ;
        RECT 512.850 458.250 516.600 459.300 ;
        RECT 470.850 458.100 472.050 458.250 ;
        RECT 491.850 458.100 493.050 458.250 ;
        RECT 512.850 458.100 514.050 458.250 ;
        RECT 529.800 458.100 531.000 461.400 ;
        RECT 535.800 460.500 537.000 464.400 ;
        RECT 550.800 461.400 552.600 467.400 ;
        RECT 563.400 464.400 565.200 467.400 ;
        RECT 531.900 459.600 537.000 460.500 ;
        RECT 531.900 458.700 533.850 459.600 ;
        RECT 532.950 458.100 533.850 458.700 ;
        RECT 455.100 456.150 456.900 456.900 ;
        RECT 463.950 454.950 466.050 457.050 ;
        RECT 467.100 455.100 468.900 455.850 ;
        RECT 469.950 454.950 472.050 457.050 ;
        RECT 473.100 455.100 474.900 455.850 ;
        RECT 484.950 454.950 487.050 457.050 ;
        RECT 488.100 455.100 489.900 455.850 ;
        RECT 490.800 454.950 493.050 457.050 ;
        RECT 494.100 455.100 495.900 455.850 ;
        RECT 505.950 454.950 508.050 457.050 ;
        RECT 509.100 455.100 510.900 455.850 ;
        RECT 511.950 454.950 514.050 457.050 ;
        RECT 515.100 455.100 516.900 455.850 ;
        RECT 529.950 454.950 532.050 457.050 ;
        RECT 451.950 451.950 457.050 454.050 ;
        RECT 464.100 453.150 465.900 453.900 ;
        RECT 466.950 451.950 469.050 454.050 ;
        RECT 470.100 450.900 471.150 453.900 ;
        RECT 485.100 453.150 486.900 453.900 ;
        RECT 487.950 451.950 490.050 454.050 ;
        RECT 491.100 450.900 492.150 453.900 ;
        RECT 493.950 451.950 496.050 454.050 ;
        RECT 506.100 453.150 507.900 453.900 ;
        RECT 508.950 451.950 511.050 454.050 ;
        RECT 512.100 450.900 513.150 453.900 ;
        RECT 514.950 451.950 517.050 454.050 ;
        RECT 533.100 453.900 533.850 458.100 ;
        RECT 535.950 454.950 538.200 457.050 ;
        RECT 550.950 455.100 552.300 461.400 ;
        RECT 564.000 460.500 565.200 464.400 ;
        RECT 569.700 461.400 571.500 467.400 ;
        RECT 574.950 463.950 577.050 466.050 ;
        RECT 584.400 464.400 586.200 467.400 ;
        RECT 601.800 464.400 603.600 467.400 ;
        RECT 564.000 459.600 569.100 460.500 ;
        RECT 567.150 458.700 569.100 459.600 ;
        RECT 567.150 458.100 568.050 458.700 ;
        RECT 570.000 458.100 571.200 461.400 ;
        RECT 554.100 455.100 555.900 455.850 ;
        RECT 452.400 441.600 453.600 450.900 ;
        RECT 469.950 447.600 471.150 450.900 ;
        RECT 490.950 447.600 492.150 450.900 ;
        RECT 511.950 447.600 513.150 450.900 ;
        RECT 529.800 447.600 531.000 453.900 ;
        RECT 532.950 450.300 533.850 453.900 ;
        RECT 536.100 453.150 537.900 453.900 ;
        RECT 547.950 451.950 550.050 454.050 ;
        RECT 551.100 450.900 552.300 455.100 ;
        RECT 562.950 454.950 565.050 457.050 ;
        RECT 553.950 451.950 556.050 454.050 ;
        RECT 567.150 453.900 567.900 458.100 ;
        RECT 568.950 456.450 571.050 457.050 ;
        RECT 575.550 456.450 576.450 463.950 ;
        RECT 580.950 457.950 583.050 460.050 ;
        RECT 568.950 455.550 576.450 456.450 ;
        RECT 581.100 456.150 582.900 456.900 ;
        RECT 568.950 454.950 571.050 455.550 ;
        RECT 584.400 455.100 585.600 464.400 ;
        RECT 602.400 461.100 603.600 464.400 ;
        RECT 617.400 464.400 619.200 467.400 ;
        RECT 634.800 464.400 636.600 467.400 ;
        RECT 601.950 457.950 604.050 460.050 ;
        RECT 613.950 457.950 616.050 460.050 ;
        RECT 598.950 454.950 601.050 457.050 ;
        RECT 563.100 453.150 564.900 453.900 ;
        RECT 531.900 449.400 533.850 450.300 ;
        RECT 531.900 448.500 537.600 449.400 ;
        RECT 445.950 436.950 448.050 439.050 ;
        RECT 451.800 435.600 453.600 441.600 ;
        RECT 469.500 435.600 471.300 447.600 ;
        RECT 490.500 435.600 492.300 447.600 ;
        RECT 511.500 435.600 513.300 447.600 ;
        RECT 529.500 435.600 531.300 447.600 ;
        RECT 536.400 441.600 537.600 448.500 ;
        RECT 538.800 445.950 540.900 448.050 ;
        RECT 550.950 447.600 552.300 450.900 ;
        RECT 567.150 450.300 568.050 453.900 ;
        RECT 567.150 449.400 569.100 450.300 ;
        RECT 563.400 448.500 569.100 449.400 ;
        RECT 535.800 435.600 537.600 441.600 ;
        RECT 539.550 439.050 540.450 445.950 ;
        RECT 538.950 436.950 541.050 439.050 ;
        RECT 550.800 435.600 552.600 447.600 ;
        RECT 563.400 441.600 564.600 448.500 ;
        RECT 570.000 447.600 571.200 453.900 ;
        RECT 583.950 451.950 589.050 454.050 ;
        RECT 602.100 453.900 603.300 456.900 ;
        RECT 614.100 456.150 615.900 456.900 ;
        RECT 617.400 455.100 618.600 464.400 ;
        RECT 635.400 461.100 636.600 464.400 ;
        RECT 647.400 462.300 649.200 467.400 ;
        RECT 653.400 462.300 655.200 467.400 ;
        RECT 647.400 460.950 655.200 462.300 ;
        RECT 656.400 461.400 658.200 467.400 ;
        RECT 634.800 457.950 637.050 460.050 ;
        RECT 656.400 459.300 657.600 461.400 ;
        RECT 672.000 460.200 673.800 467.400 ;
        RECT 691.200 461.400 693.000 467.400 ;
        RECT 672.000 459.300 675.600 460.200 ;
        RECT 653.850 458.250 657.600 459.300 ;
        RECT 653.850 458.100 655.050 458.250 ;
        RECT 631.950 454.950 634.050 457.050 ;
        RECT 599.100 453.150 600.900 453.900 ;
        RECT 563.400 435.600 565.200 441.600 ;
        RECT 569.700 435.600 571.500 447.600 ;
        RECT 584.400 441.600 585.600 450.900 ;
        RECT 601.950 448.650 603.300 453.900 ;
        RECT 605.100 453.150 606.900 453.900 ;
        RECT 616.950 451.950 622.050 454.050 ;
        RECT 635.100 453.900 636.300 456.900 ;
        RECT 646.950 454.950 649.050 457.050 ;
        RECT 650.100 455.100 651.900 455.850 ;
        RECT 652.950 454.950 655.050 457.050 ;
        RECT 656.100 455.100 657.900 455.850 ;
        RECT 674.400 455.100 675.600 459.300 ;
        RECT 691.950 458.100 693.000 461.400 ;
        RECT 710.400 462.300 712.200 467.400 ;
        RECT 716.400 462.300 718.200 467.400 ;
        RECT 710.400 460.950 718.200 462.300 ;
        RECT 719.400 461.400 721.200 467.400 ;
        RECT 719.400 459.300 720.600 461.400 ;
        RECT 736.200 460.200 738.000 467.400 ;
        RECT 716.850 458.250 720.600 459.300 ;
        RECT 734.400 459.300 738.000 460.200 ;
        RECT 716.850 458.100 718.050 458.250 ;
        RECT 685.950 454.950 688.050 457.050 ;
        RECT 689.250 455.100 690.900 455.850 ;
        RECT 691.950 454.950 694.050 457.050 ;
        RECT 695.100 455.100 696.750 455.850 ;
        RECT 697.950 454.950 700.050 457.050 ;
        RECT 709.950 454.950 712.050 457.050 ;
        RECT 713.100 455.100 714.900 455.850 ;
        RECT 715.950 454.950 718.050 457.050 ;
        RECT 719.100 455.100 720.900 455.850 ;
        RECT 734.400 455.100 735.600 459.300 ;
        RECT 755.100 459.000 756.900 467.400 ;
        RECT 776.100 459.000 777.900 467.400 ;
        RECT 793.800 461.400 795.600 467.400 ;
        RECT 794.400 459.300 795.600 461.400 ;
        RECT 796.800 462.300 798.600 467.400 ;
        RECT 802.800 462.300 804.600 467.400 ;
        RECT 796.800 460.950 804.600 462.300 ;
        RECT 814.800 461.400 816.600 467.400 ;
        RECT 815.400 459.300 816.600 461.400 ;
        RECT 817.800 462.300 819.600 467.400 ;
        RECT 823.800 462.300 825.600 467.400 ;
        RECT 836.400 464.400 838.200 467.400 ;
        RECT 817.800 460.950 825.600 462.300 ;
        RECT 837.300 460.200 838.200 464.400 ;
        RECT 842.400 461.400 844.200 467.400 ;
        RECT 755.100 457.350 759.300 459.000 ;
        RECT 776.100 457.350 780.300 459.000 ;
        RECT 794.400 458.250 798.150 459.300 ;
        RECT 815.400 458.250 819.150 459.300 ;
        RECT 796.950 458.100 798.150 458.250 ;
        RECT 817.950 458.100 819.150 458.250 ;
        RECT 832.950 457.950 835.050 460.050 ;
        RECT 837.300 459.300 840.750 460.200 ;
        RECT 838.950 458.400 840.750 459.300 ;
        RECT 749.100 455.100 750.900 455.850 ;
        RECT 755.100 455.100 756.900 455.850 ;
        RECT 632.100 453.150 633.900 453.900 ;
        RECT 607.950 448.950 610.050 451.050 ;
        RECT 600.600 447.600 603.300 448.650 ;
        RECT 584.400 435.600 586.200 441.600 ;
        RECT 600.600 435.600 602.400 447.600 ;
        RECT 608.550 442.050 609.450 448.950 ;
        RECT 607.800 439.950 609.900 442.050 ;
        RECT 617.400 441.600 618.600 450.900 ;
        RECT 634.950 448.650 636.300 453.900 ;
        RECT 638.100 453.150 639.900 453.900 ;
        RECT 647.100 453.150 648.900 453.900 ;
        RECT 649.950 451.950 652.200 454.050 ;
        RECT 653.100 450.900 654.150 453.900 ;
        RECT 655.950 451.950 658.050 454.050 ;
        RECT 671.100 452.100 672.900 452.850 ;
        RECT 673.950 451.950 676.050 454.050 ;
        RECT 686.250 453.150 687.900 453.900 ;
        RECT 677.100 452.100 678.900 452.850 ;
        RECT 688.950 451.950 691.050 454.050 ;
        RECT 633.600 447.600 636.300 448.650 ;
        RECT 617.400 435.600 619.200 441.600 ;
        RECT 633.600 435.600 635.400 447.600 ;
        RECT 641.100 445.950 643.200 448.050 ;
        RECT 652.950 447.600 654.150 450.900 ;
        RECT 656.550 450.000 657.450 451.950 ;
        RECT 641.550 439.050 642.450 445.950 ;
        RECT 640.800 436.950 642.900 439.050 ;
        RECT 652.500 435.600 654.300 447.600 ;
        RECT 655.950 445.950 658.050 450.000 ;
        RECT 670.950 448.950 673.050 451.050 ;
        RECT 674.400 441.600 675.600 450.900 ;
        RECT 676.950 448.950 679.200 451.050 ;
        RECT 693.150 450.900 693.900 453.900 ;
        RECT 694.950 451.950 697.050 454.050 ;
        RECT 698.100 453.150 699.900 453.900 ;
        RECT 710.100 453.150 711.900 453.900 ;
        RECT 712.800 451.950 715.050 454.050 ;
        RECT 716.100 450.900 717.150 453.900 ;
        RECT 718.950 451.950 721.050 454.050 ;
        RECT 731.100 452.100 732.900 452.850 ;
        RECT 733.950 451.950 736.200 454.050 ;
        RECT 737.100 452.100 738.900 452.850 ;
        RECT 742.800 451.950 744.900 454.050 ;
        RECT 748.950 451.950 751.050 454.050 ;
        RECT 754.950 451.950 757.050 454.050 ;
        RECT 758.400 452.100 759.300 457.350 ;
        RECT 770.100 455.100 771.900 455.850 ;
        RECT 776.100 455.100 777.900 455.850 ;
        RECT 769.950 451.950 772.050 454.050 ;
        RECT 775.950 451.950 778.050 454.050 ;
        RECT 779.400 452.100 780.300 457.350 ;
        RECT 784.950 454.950 787.050 457.050 ;
        RECT 794.100 455.100 795.900 455.850 ;
        RECT 796.800 454.950 799.050 457.050 ;
        RECT 800.100 455.100 801.900 455.850 ;
        RECT 802.950 454.950 805.200 457.050 ;
        RECT 808.950 454.950 811.050 457.050 ;
        RECT 815.100 455.100 816.900 455.850 ;
        RECT 817.950 454.950 820.050 457.050 ;
        RECT 821.100 455.100 822.900 455.850 ;
        RECT 823.950 454.950 826.050 457.050 ;
        RECT 833.100 456.150 834.900 456.900 ;
        RECT 835.950 454.950 838.050 457.050 ;
        RECT 693.150 449.400 694.050 450.900 ;
        RECT 693.150 448.500 697.200 449.400 ;
        RECT 673.800 435.600 675.600 441.600 ;
        RECT 686.400 446.400 694.200 447.300 ;
        RECT 686.400 435.600 688.200 446.400 ;
        RECT 692.400 436.500 694.200 446.400 ;
        RECT 695.400 437.400 697.200 448.500 ;
        RECT 715.950 447.600 717.150 450.900 ;
        RECT 724.950 448.950 727.050 451.050 ;
        RECT 730.950 448.950 733.200 451.050 ;
        RECT 698.400 436.500 700.200 447.600 ;
        RECT 692.400 435.600 700.200 436.500 ;
        RECT 715.500 435.600 717.300 447.600 ;
        RECT 725.550 442.050 726.450 448.950 ;
        RECT 724.950 439.950 727.050 442.050 ;
        RECT 734.400 441.600 735.600 450.900 ;
        RECT 736.950 448.950 739.050 451.050 ;
        RECT 743.550 445.050 744.450 451.950 ;
        RECT 751.950 448.950 754.050 451.050 ;
        RECT 757.950 450.450 760.050 451.050 ;
        RECT 762.000 450.450 766.050 451.050 ;
        RECT 757.950 449.550 766.050 450.450 ;
        RECT 757.950 448.950 760.050 449.550 ;
        RECT 762.000 448.950 766.050 449.550 ;
        RECT 772.950 448.950 775.050 451.050 ;
        RECT 778.950 450.450 781.050 451.050 ;
        RECT 785.550 450.450 786.450 454.950 ;
        RECT 793.950 451.950 796.050 454.050 ;
        RECT 778.950 449.550 786.450 450.450 ;
        RECT 797.850 450.900 798.900 453.900 ;
        RECT 799.800 451.950 802.050 454.050 ;
        RECT 803.100 453.150 804.900 453.900 ;
        RECT 778.950 448.950 781.050 449.550 ;
        RECT 752.100 447.150 753.900 447.900 ;
        RECT 742.950 442.950 745.050 445.050 ;
        RECT 758.400 442.800 759.300 447.900 ;
        RECT 773.100 447.150 774.900 447.900 ;
        RECT 779.400 442.800 780.300 447.900 ;
        RECT 797.850 447.600 799.050 450.900 ;
        RECT 752.700 441.900 759.300 442.800 ;
        RECT 752.700 441.600 754.200 441.900 ;
        RECT 734.400 435.600 736.200 441.600 ;
        RECT 752.400 435.600 754.200 441.600 ;
        RECT 758.400 441.600 759.300 441.900 ;
        RECT 773.700 441.900 780.300 442.800 ;
        RECT 773.700 441.600 775.200 441.900 ;
        RECT 758.400 435.600 760.200 441.600 ;
        RECT 773.400 435.600 775.200 441.600 ;
        RECT 779.400 441.600 780.300 441.900 ;
        RECT 779.400 435.600 781.200 441.600 ;
        RECT 797.700 435.600 799.500 447.600 ;
        RECT 809.550 439.050 810.450 454.950 ;
        RECT 814.950 451.950 817.050 454.050 ;
        RECT 818.850 450.900 819.900 453.900 ;
        RECT 820.950 451.950 823.050 454.050 ;
        RECT 824.100 453.150 825.900 453.900 ;
        RECT 836.100 453.150 837.900 453.900 ;
        RECT 818.850 447.600 820.050 450.900 ;
        RECT 839.700 450.600 840.600 458.400 ;
        RECT 843.000 455.100 844.050 461.400 ;
        RECT 841.950 451.950 844.050 454.050 ;
        RECT 838.800 450.000 840.600 450.600 ;
        RECT 833.400 448.800 840.600 450.000 ;
        RECT 833.400 447.600 834.600 448.800 ;
        RECT 839.700 448.650 840.600 448.800 ;
        RECT 841.950 447.600 843.300 450.900 ;
        RECT 808.950 436.950 811.050 439.050 ;
        RECT 818.700 435.600 820.500 447.600 ;
        RECT 833.400 435.600 835.200 447.600 ;
        RECT 840.900 446.100 843.300 447.600 ;
        RECT 840.900 435.600 842.700 446.100 ;
        RECT 14.700 419.400 16.500 431.400 ;
        RECT 31.800 425.400 33.600 431.400 ;
        RECT 32.700 425.100 33.600 425.400 ;
        RECT 37.800 425.400 39.600 431.400 ;
        RECT 37.800 425.100 39.300 425.400 ;
        RECT 32.700 424.200 39.300 425.100 ;
        RECT 14.850 416.100 16.050 419.400 ;
        RECT 32.700 419.100 33.600 424.200 ;
        RECT 38.100 419.100 39.900 419.850 ;
        RECT 52.800 419.400 54.600 431.400 ;
        RECT 55.800 420.300 57.600 431.400 ;
        RECT 61.800 420.300 63.600 431.400 ;
        RECT 55.800 419.400 63.600 420.300 ;
        RECT 77.700 419.400 79.500 431.400 ;
        RECT 94.800 425.400 96.600 431.400 ;
        RECT 10.800 412.950 13.050 415.050 ;
        RECT 14.850 413.100 15.900 416.100 ;
        RECT 25.950 415.950 28.050 418.050 ;
        RECT 31.950 415.950 34.050 418.050 ;
        RECT 37.950 415.950 40.050 418.050 ;
        RECT 16.950 412.950 19.200 415.050 ;
        RECT 20.100 413.100 21.900 413.850 ;
        RECT 26.550 412.050 27.450 415.950 ;
        RECT 11.100 411.150 12.900 411.900 ;
        RECT 13.800 409.950 16.050 412.050 ;
        RECT 17.100 411.150 18.900 411.900 ;
        RECT 19.950 409.950 22.050 412.050 ;
        RECT 26.100 409.950 28.200 412.050 ;
        RECT 32.700 409.650 33.600 414.900 ;
        RECT 34.950 412.950 37.050 415.050 ;
        RECT 40.950 412.950 43.050 415.050 ;
        RECT 53.400 413.100 54.300 419.400 ;
        RECT 55.950 412.950 58.050 418.050 ;
        RECT 77.850 416.100 79.050 419.400 ;
        RECT 95.400 416.100 96.600 425.400 ;
        RECT 113.700 419.400 115.500 431.400 ;
        RECT 133.500 419.400 135.300 431.400 ;
        RECT 154.800 425.400 156.600 431.400 ;
        RECT 113.850 416.100 115.050 419.400 ;
        RECT 133.950 416.100 135.150 419.400 ;
        RECT 59.100 413.100 60.900 413.850 ;
        RECT 61.950 412.950 64.200 415.050 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 77.850 413.100 78.900 416.100 ;
        RECT 79.950 412.950 82.050 415.050 ;
        RECT 83.100 413.100 84.900 413.850 ;
        RECT 94.950 412.950 100.050 415.050 ;
        RECT 109.950 412.950 112.050 415.050 ;
        RECT 113.850 413.100 114.900 416.100 ;
        RECT 115.950 412.950 118.050 415.050 ;
        RECT 119.100 413.100 120.900 413.850 ;
        RECT 128.100 413.100 129.900 413.850 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 134.100 413.100 135.150 416.100 ;
        RECT 146.100 415.950 148.200 418.050 ;
        RECT 151.950 415.950 154.050 418.050 ;
        RECT 155.400 416.100 156.600 425.400 ;
        RECT 170.400 425.400 172.200 431.400 ;
        RECT 188.400 425.400 190.200 431.400 ;
        RECT 157.950 415.950 160.050 418.050 ;
        RECT 166.950 415.950 169.050 418.050 ;
        RECT 170.400 416.100 171.600 425.400 ;
        RECT 184.950 420.000 187.050 424.050 ;
        RECT 185.550 418.050 186.450 420.000 ;
        RECT 172.950 415.950 175.050 418.050 ;
        RECT 184.950 415.950 187.050 418.050 ;
        RECT 188.400 416.100 189.600 425.400 ;
        RECT 205.200 419.400 207.000 431.400 ;
        RECT 211.800 425.400 213.600 431.400 ;
        RECT 190.950 415.950 193.050 418.050 ;
        RECT 136.950 412.950 139.050 415.050 ;
        RECT 35.100 411.150 36.900 411.900 ;
        RECT 41.100 411.150 42.900 411.900 ;
        RECT 49.950 409.950 55.050 412.050 ;
        RECT 56.100 411.150 57.900 411.900 ;
        RECT 58.950 409.950 61.050 412.050 ;
        RECT 62.100 411.150 63.900 411.900 ;
        RECT 74.100 411.150 75.900 411.900 ;
        RECT 76.950 409.950 79.050 412.050 ;
        RECT 80.100 411.150 81.900 411.900 ;
        RECT 82.950 409.950 85.050 412.050 ;
        RECT 13.950 408.750 15.150 408.900 ;
        RECT 11.400 407.700 15.150 408.750 ;
        RECT 32.700 408.000 36.900 409.650 ;
        RECT 11.400 405.600 12.600 407.700 ;
        RECT 10.800 399.600 12.600 405.600 ;
        RECT 13.800 404.700 21.600 406.050 ;
        RECT 13.800 399.600 15.600 404.700 ;
        RECT 19.800 399.600 21.600 404.700 ;
        RECT 35.100 399.600 36.900 408.000 ;
        RECT 53.400 405.600 54.300 408.900 ;
        RECT 76.950 408.750 78.150 408.900 ;
        RECT 74.400 407.700 78.150 408.750 ;
        RECT 74.400 405.600 75.600 407.700 ;
        RECT 53.400 403.950 58.800 405.600 ;
        RECT 57.000 399.600 58.800 403.950 ;
        RECT 73.800 399.600 75.600 405.600 ;
        RECT 76.800 404.700 84.600 406.050 ;
        RECT 76.800 399.600 78.600 404.700 ;
        RECT 82.800 399.600 84.600 404.700 ;
        RECT 95.400 402.600 96.600 411.900 ;
        RECT 110.100 411.150 111.900 411.900 ;
        RECT 98.100 410.100 99.900 410.850 ;
        RECT 112.950 409.950 115.050 412.050 ;
        RECT 116.100 411.150 117.900 411.900 ;
        RECT 118.950 409.950 121.050 412.050 ;
        RECT 127.950 409.950 130.050 412.050 ;
        RECT 131.100 411.150 132.900 411.900 ;
        RECT 133.950 409.950 136.200 412.050 ;
        RECT 137.100 411.150 138.900 411.900 ;
        RECT 146.550 409.050 147.450 415.950 ;
        RECT 152.100 414.150 153.900 414.900 ;
        RECT 154.800 412.950 157.050 415.050 ;
        RECT 158.100 414.150 159.900 414.900 ;
        RECT 167.100 414.150 168.900 414.900 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 173.100 414.150 174.900 414.900 ;
        RECT 185.100 414.150 186.900 414.900 ;
        RECT 187.950 412.950 190.200 415.050 ;
        RECT 191.100 414.150 192.900 414.900 ;
        RECT 205.950 413.100 207.000 419.400 ;
        RECT 208.950 412.950 211.050 418.050 ;
        RECT 97.950 406.950 100.050 409.050 ;
        RECT 112.950 408.750 114.150 408.900 ;
        RECT 110.400 407.700 114.150 408.750 ;
        RECT 134.850 408.750 136.050 408.900 ;
        RECT 134.850 407.700 138.600 408.750 ;
        RECT 110.400 405.600 111.600 407.700 ;
        RECT 94.800 399.600 96.600 402.600 ;
        RECT 109.800 399.600 111.600 405.600 ;
        RECT 112.800 404.700 120.600 406.050 ;
        RECT 112.800 399.600 114.600 404.700 ;
        RECT 118.800 399.600 120.600 404.700 ;
        RECT 128.400 404.700 136.200 406.050 ;
        RECT 128.400 399.600 130.200 404.700 ;
        RECT 134.400 399.600 136.200 404.700 ;
        RECT 137.400 405.600 138.600 407.700 ;
        RECT 145.950 406.950 148.050 409.050 ;
        RECT 155.400 407.700 156.600 411.900 ;
        RECT 153.000 406.800 156.600 407.700 ;
        RECT 170.400 407.700 171.600 411.900 ;
        RECT 188.400 407.700 189.600 411.900 ;
        RECT 205.950 411.450 208.050 412.050 ;
        RECT 200.550 411.000 208.050 411.450 ;
        RECT 209.100 411.150 210.900 411.900 ;
        RECT 199.950 410.550 208.050 411.000 ;
        RECT 170.400 406.800 174.000 407.700 ;
        RECT 188.400 406.800 192.000 407.700 ;
        RECT 199.950 406.950 202.050 410.550 ;
        RECT 205.950 409.950 208.050 410.550 ;
        RECT 137.400 399.600 139.200 405.600 ;
        RECT 153.000 399.600 154.800 406.800 ;
        RECT 172.200 399.600 174.000 406.800 ;
        RECT 190.200 399.600 192.000 406.800 ;
        RECT 207.150 405.600 208.050 408.900 ;
        RECT 212.550 408.300 213.600 425.400 ;
        RECT 224.400 420.600 226.200 431.400 ;
        RECT 230.400 430.500 238.200 431.400 ;
        RECT 230.400 420.600 232.200 430.500 ;
        RECT 224.400 419.700 232.200 420.600 ;
        RECT 233.400 418.500 235.200 429.600 ;
        RECT 236.400 419.400 238.200 430.500 ;
        RECT 241.950 427.950 244.050 430.050 ;
        RECT 231.150 417.600 235.200 418.500 ;
        RECT 231.150 416.100 232.050 417.600 ;
        RECT 215.100 413.100 216.900 413.850 ;
        RECT 224.250 413.100 225.900 413.850 ;
        RECT 226.950 412.950 229.050 415.050 ;
        RECT 231.150 413.100 231.900 416.100 ;
        RECT 232.950 412.950 235.050 415.050 ;
        RECT 236.100 413.100 237.900 413.850 ;
        RECT 214.950 409.950 217.050 412.050 ;
        RECT 223.800 409.950 226.050 412.050 ;
        RECT 227.250 411.150 228.900 411.900 ;
        RECT 229.950 409.950 232.050 412.050 ;
        RECT 233.100 411.150 234.750 411.900 ;
        RECT 235.950 409.950 238.050 412.050 ;
        RECT 242.550 409.050 243.450 427.950 ;
        RECT 248.400 425.400 250.200 431.400 ;
        RECT 248.400 418.500 249.600 425.400 ;
        RECT 254.700 419.400 256.500 431.400 ;
        RECT 266.400 425.400 268.200 431.400 ;
        RECT 248.400 417.600 254.100 418.500 ;
        RECT 252.150 416.700 254.100 417.600 ;
        RECT 248.100 413.100 249.900 413.850 ;
        RECT 252.150 413.100 253.050 416.700 ;
        RECT 255.000 413.100 256.200 419.400 ;
        RECT 266.400 418.500 267.600 425.400 ;
        RECT 272.700 419.400 274.500 431.400 ;
        RECT 280.950 427.950 283.050 430.050 ;
        RECT 266.400 417.600 272.100 418.500 ;
        RECT 270.150 416.700 272.100 417.600 ;
        RECT 266.100 413.100 267.900 413.850 ;
        RECT 270.150 413.100 271.050 416.700 ;
        RECT 273.000 413.100 274.200 419.400 ;
        RECT 281.550 415.050 282.450 427.950 ;
        RECT 289.800 425.400 291.600 431.400 ;
        RECT 286.950 415.950 289.050 418.050 ;
        RECT 290.400 416.100 291.600 425.400 ;
        RECT 308.700 419.400 310.500 431.400 ;
        RECT 326.400 425.400 328.200 431.400 ;
        RECT 317.100 421.950 319.200 424.050 ;
        RECT 292.950 415.950 295.050 418.050 ;
        RECT 308.850 416.100 310.050 419.400 ;
        RECT 317.550 418.050 318.450 421.950 ;
        RECT 247.950 409.950 250.050 412.050 ;
        RECT 209.100 407.100 216.600 408.300 ;
        RECT 209.100 406.500 210.900 407.100 ;
        RECT 207.150 403.800 209.100 405.600 ;
        RECT 207.300 399.600 209.100 403.800 ;
        RECT 214.800 399.600 216.600 407.100 ;
        RECT 229.950 405.600 231.000 408.900 ;
        RECT 241.950 406.950 244.050 409.050 ;
        RECT 252.150 408.900 252.900 413.100 ;
        RECT 253.950 409.950 256.050 412.050 ;
        RECT 265.950 409.950 268.050 412.050 ;
        RECT 270.150 408.900 270.900 413.100 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 287.100 414.150 288.900 414.900 ;
        RECT 289.950 412.950 292.050 415.050 ;
        RECT 293.100 414.150 294.900 414.900 ;
        RECT 298.950 412.950 301.050 415.050 ;
        RECT 304.950 412.950 307.050 415.050 ;
        RECT 308.850 413.100 309.900 416.100 ;
        RECT 316.950 415.950 319.050 418.050 ;
        RECT 322.950 415.950 325.050 418.050 ;
        RECT 326.400 416.100 327.600 425.400 ;
        RECT 343.200 419.400 345.000 431.400 ;
        RECT 349.800 425.400 351.600 431.400 ;
        RECT 328.950 415.950 331.200 418.050 ;
        RECT 337.950 415.950 340.050 418.050 ;
        RECT 310.950 412.950 313.050 415.050 ;
        RECT 323.100 414.150 324.900 414.900 ;
        RECT 314.100 413.100 315.900 413.850 ;
        RECT 325.950 412.950 328.050 415.050 ;
        RECT 329.100 414.150 330.900 414.900 ;
        RECT 271.950 409.950 274.050 412.050 ;
        RECT 252.150 408.300 253.050 408.900 ;
        RECT 252.150 407.400 254.100 408.300 ;
        RECT 229.200 399.600 231.000 405.600 ;
        RECT 249.000 406.500 254.100 407.400 ;
        RECT 249.000 402.600 250.200 406.500 ;
        RECT 255.000 405.600 256.200 408.900 ;
        RECT 270.150 408.300 271.050 408.900 ;
        RECT 270.150 407.400 272.100 408.300 ;
        RECT 267.000 406.500 272.100 407.400 ;
        RECT 248.400 399.600 250.200 402.600 ;
        RECT 254.700 399.600 256.500 405.600 ;
        RECT 267.000 402.600 268.200 406.500 ;
        RECT 273.000 405.600 274.200 408.900 ;
        RECT 290.400 407.700 291.600 411.900 ;
        RECT 288.000 406.800 291.600 407.700 ;
        RECT 266.400 399.600 268.200 402.600 ;
        RECT 272.700 399.600 274.500 405.600 ;
        RECT 288.000 399.600 289.800 406.800 ;
        RECT 299.550 406.050 300.450 412.950 ;
        RECT 305.100 411.150 306.900 411.900 ;
        RECT 307.950 409.950 310.050 412.050 ;
        RECT 311.100 411.150 312.900 411.900 ;
        RECT 313.950 409.950 316.050 412.050 ;
        RECT 307.950 408.750 309.150 408.900 ;
        RECT 305.400 407.700 309.150 408.750 ;
        RECT 326.400 407.700 327.600 411.900 ;
        RECT 338.550 411.450 339.450 415.950 ;
        RECT 343.950 413.100 345.000 419.400 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 343.950 411.450 346.050 412.050 ;
        RECT 338.550 410.550 346.050 411.450 ;
        RECT 347.100 411.150 348.900 411.900 ;
        RECT 343.950 409.950 346.050 410.550 ;
        RECT 298.950 403.950 301.050 406.050 ;
        RECT 305.400 405.600 306.600 407.700 ;
        RECT 326.400 406.800 330.000 407.700 ;
        RECT 304.800 399.600 306.600 405.600 ;
        RECT 307.800 404.700 315.600 406.050 ;
        RECT 307.800 399.600 309.600 404.700 ;
        RECT 313.800 399.600 315.600 404.700 ;
        RECT 328.200 399.600 330.000 406.800 ;
        RECT 345.150 405.600 346.050 408.900 ;
        RECT 350.550 408.300 351.600 425.400 ;
        RECT 365.400 425.400 367.200 431.400 ;
        RECT 361.800 415.950 364.050 418.050 ;
        RECT 365.400 416.100 366.600 425.400 ;
        RECT 380.400 420.300 382.200 431.400 ;
        RECT 386.400 420.300 388.200 431.400 ;
        RECT 380.400 419.400 388.200 420.300 ;
        RECT 389.400 419.400 391.200 431.400 ;
        RECT 403.500 419.400 405.300 431.400 ;
        RECT 409.800 425.400 411.600 431.400 ;
        RECT 367.950 415.950 370.050 418.050 ;
        RECT 362.100 414.150 363.900 414.900 ;
        RECT 353.100 413.100 354.900 413.850 ;
        RECT 364.950 412.950 367.050 415.050 ;
        RECT 368.100 414.150 369.900 414.900 ;
        RECT 379.950 412.950 382.050 418.050 ;
        RECT 383.100 413.100 384.900 413.850 ;
        RECT 385.950 412.950 388.050 415.050 ;
        RECT 389.700 413.100 390.600 419.400 ;
        RECT 403.800 413.100 405.000 419.400 ;
        RECT 410.400 418.500 411.600 425.400 ;
        RECT 424.500 419.400 426.300 431.400 ;
        RECT 445.500 419.400 447.300 431.400 ;
        RECT 463.800 425.400 465.600 431.400 ;
        RECT 405.900 417.600 411.600 418.500 ;
        RECT 405.900 416.700 407.850 417.600 ;
        RECT 406.950 413.100 407.850 416.700 ;
        RECT 424.950 416.100 426.150 419.400 ;
        RECT 445.950 416.100 447.150 419.400 ;
        RECT 464.400 416.100 465.600 425.400 ;
        RECT 470.550 419.400 472.350 431.400 ;
        RECT 478.050 425.400 479.850 431.400 ;
        RECT 475.950 423.300 479.850 425.400 ;
        RECT 485.850 424.500 487.650 431.400 ;
        RECT 493.650 425.400 495.450 431.400 ;
        RECT 494.250 424.500 495.450 425.400 ;
        RECT 484.950 423.450 491.550 424.500 ;
        RECT 484.950 422.700 486.750 423.450 ;
        RECT 489.750 422.700 491.550 423.450 ;
        RECT 494.250 422.400 499.050 424.500 ;
        RECT 477.150 420.600 479.850 422.400 ;
        RECT 480.750 421.800 482.550 422.400 ;
        RECT 480.750 420.900 487.050 421.800 ;
        RECT 494.250 421.500 495.450 422.400 ;
        RECT 480.750 420.600 482.550 420.900 ;
        RECT 478.950 419.700 479.850 420.600 ;
        RECT 410.100 413.100 411.900 413.850 ;
        RECT 419.100 413.100 420.900 413.850 ;
        RECT 352.950 409.950 355.050 412.050 ;
        RECT 347.100 407.100 354.600 408.300 ;
        RECT 347.100 406.500 348.900 407.100 ;
        RECT 345.150 403.800 347.100 405.600 ;
        RECT 345.300 399.600 347.100 403.800 ;
        RECT 352.800 399.600 354.600 407.100 ;
        RECT 365.400 407.700 366.600 411.900 ;
        RECT 380.100 411.150 381.900 411.900 ;
        RECT 382.800 409.950 385.050 412.050 ;
        RECT 386.100 411.150 387.900 411.900 ;
        RECT 388.950 411.450 391.050 412.050 ;
        RECT 388.950 410.550 396.450 411.450 ;
        RECT 388.950 409.950 391.050 410.550 ;
        RECT 365.400 406.800 369.000 407.700 ;
        RECT 367.200 399.600 369.000 406.800 ;
        RECT 389.700 405.600 390.600 408.900 ;
        RECT 395.550 406.050 396.450 410.550 ;
        RECT 407.100 408.900 407.850 413.100 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 425.100 413.100 426.150 416.100 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 440.100 413.100 441.900 413.850 ;
        RECT 442.950 412.950 445.050 415.050 ;
        RECT 446.100 413.100 447.150 416.100 ;
        RECT 448.950 412.950 451.050 415.050 ;
        RECT 463.950 412.950 466.050 415.050 ;
        RECT 470.550 412.050 471.750 419.400 ;
        RECT 475.950 418.800 478.050 419.700 ;
        RECT 478.950 418.800 484.950 419.700 ;
        RECT 473.850 417.600 478.050 418.800 ;
        RECT 472.950 415.800 474.750 417.600 ;
        RECT 484.050 413.100 484.950 418.800 ;
        RECT 486.150 418.800 487.050 420.900 ;
        RECT 487.950 420.300 495.450 421.500 ;
        RECT 487.950 419.700 489.750 420.300 ;
        RECT 502.050 419.400 503.850 431.400 ;
        RECT 492.750 418.800 503.850 419.400 ;
        RECT 505.950 418.950 508.050 421.050 ;
        RECT 517.500 419.400 519.300 431.400 ;
        RECT 536.400 425.400 538.200 431.400 ;
        RECT 486.150 418.200 503.850 418.800 ;
        RECT 486.150 417.900 494.550 418.200 ;
        RECT 492.750 417.600 494.550 417.900 ;
        RECT 497.100 412.800 498.900 413.100 ;
        RECT 409.950 409.950 412.050 412.050 ;
        RECT 418.950 409.950 421.050 412.050 ;
        RECT 422.100 411.150 423.900 411.900 ;
        RECT 424.950 409.950 427.050 412.050 ;
        RECT 428.100 411.150 429.900 411.900 ;
        RECT 439.950 409.950 442.050 412.050 ;
        RECT 443.100 411.150 444.900 411.900 ;
        RECT 445.950 409.950 448.050 412.050 ;
        RECT 449.100 411.150 450.900 411.900 ;
        RECT 385.200 403.950 390.600 405.600 ;
        RECT 394.950 403.950 397.050 406.050 ;
        RECT 403.800 405.600 405.000 408.900 ;
        RECT 406.950 408.300 407.850 408.900 ;
        RECT 405.900 407.400 407.850 408.300 ;
        RECT 425.850 408.750 427.050 408.900 ;
        RECT 446.850 408.750 448.050 408.900 ;
        RECT 425.850 407.700 429.600 408.750 ;
        RECT 446.850 407.700 450.600 408.750 ;
        RECT 405.900 406.500 411.000 407.400 ;
        RECT 385.200 399.600 387.000 403.950 ;
        RECT 403.500 399.600 405.300 405.600 ;
        RECT 409.800 402.600 411.000 406.500 ;
        RECT 419.400 404.700 427.200 406.050 ;
        RECT 409.800 399.600 411.600 402.600 ;
        RECT 419.400 399.600 421.200 404.700 ;
        RECT 425.400 399.600 427.200 404.700 ;
        RECT 428.400 405.600 429.600 407.700 ;
        RECT 428.400 399.600 430.200 405.600 ;
        RECT 440.400 404.700 448.200 406.050 ;
        RECT 440.400 399.600 442.200 404.700 ;
        RECT 446.400 399.600 448.200 404.700 ;
        RECT 449.400 405.600 450.600 407.700 ;
        RECT 449.400 399.600 451.200 405.600 ;
        RECT 464.400 402.600 465.600 411.900 ;
        RECT 467.100 410.100 468.900 410.850 ;
        RECT 470.550 409.950 471.900 412.050 ;
        RECT 466.950 406.950 469.050 409.050 ;
        RECT 463.800 399.600 465.600 402.600 ;
        RECT 470.550 405.600 471.750 409.950 ;
        RECT 472.950 406.950 475.050 412.050 ;
        RECT 476.100 409.950 476.850 411.750 ;
        RECT 484.950 409.950 487.050 412.050 ;
        RECT 490.950 409.950 493.050 412.050 ;
        RECT 494.100 411.900 498.900 412.800 ;
        RECT 497.100 411.300 498.900 411.900 ;
        RECT 500.100 411.150 501.900 412.950 ;
        RECT 494.100 410.400 495.900 411.000 ;
        RECT 500.100 410.400 501.000 411.150 ;
        RECT 494.100 409.200 501.000 410.400 ;
        RECT 484.050 408.000 484.950 408.900 ;
        RECT 494.100 408.000 495.150 409.200 ;
        RECT 484.050 407.100 495.150 408.000 ;
        RECT 484.050 406.800 484.950 407.100 ;
        RECT 470.550 399.600 472.350 405.600 ;
        RECT 475.950 404.700 478.050 405.600 ;
        RECT 483.150 405.000 484.950 406.800 ;
        RECT 494.100 406.200 495.150 407.100 ;
        RECT 490.350 405.450 492.150 406.200 ;
        RECT 475.950 403.500 479.700 404.700 ;
        RECT 478.650 402.600 479.700 403.500 ;
        RECT 487.200 404.400 492.150 405.450 ;
        RECT 493.650 404.400 495.450 406.200 ;
        RECT 502.950 405.600 503.850 418.200 ;
        RECT 506.550 411.450 507.450 418.950 ;
        RECT 517.950 416.100 519.150 419.400 ;
        RECT 532.950 418.050 535.050 421.050 ;
        RECT 512.100 413.100 513.900 413.850 ;
        RECT 514.950 412.950 517.050 415.050 ;
        RECT 518.100 413.100 519.150 416.100 ;
        RECT 529.950 415.950 535.050 418.050 ;
        RECT 536.400 416.100 537.600 425.400 ;
        RECT 555.600 419.400 557.400 431.400 ;
        RECT 565.950 427.950 568.050 430.050 ;
        RECT 555.600 418.350 558.300 419.400 ;
        RECT 538.950 415.950 541.050 418.050 ;
        RECT 520.950 412.950 523.050 415.050 ;
        RECT 533.100 414.150 534.900 414.900 ;
        RECT 535.800 412.950 538.050 415.050 ;
        RECT 539.100 414.150 540.900 414.900 ;
        RECT 554.100 413.100 555.900 413.850 ;
        RECT 556.950 413.100 558.300 418.350 ;
        RECT 560.100 413.100 561.900 413.850 ;
        RECT 511.950 411.450 514.050 412.050 ;
        RECT 506.550 410.550 514.050 411.450 ;
        RECT 515.100 411.150 516.900 411.900 ;
        RECT 511.950 409.950 514.050 410.550 ;
        RECT 517.950 409.950 520.050 412.050 ;
        RECT 521.100 411.150 522.900 411.900 ;
        RECT 518.850 408.750 520.050 408.900 ;
        RECT 518.850 407.700 522.600 408.750 ;
        RECT 487.200 402.600 488.250 404.400 ;
        RECT 496.950 403.500 499.050 405.600 ;
        RECT 496.950 402.600 498.000 403.500 ;
        RECT 478.650 399.600 480.450 402.600 ;
        RECT 486.450 399.600 488.250 402.600 ;
        RECT 494.250 401.700 498.000 402.600 ;
        RECT 494.250 399.600 496.050 401.700 ;
        RECT 502.050 399.600 503.850 405.600 ;
        RECT 512.400 404.700 520.200 406.050 ;
        RECT 512.400 399.600 514.200 404.700 ;
        RECT 518.400 399.600 520.200 404.700 ;
        RECT 521.400 405.600 522.600 407.700 ;
        RECT 536.400 407.700 537.600 411.900 ;
        RECT 553.950 409.950 556.050 412.050 ;
        RECT 557.100 410.100 558.300 413.100 ;
        RECT 559.950 409.950 562.050 412.050 ;
        RECT 536.400 406.800 540.000 407.700 ;
        RECT 556.950 406.950 559.050 409.050 ;
        RECT 521.400 399.600 523.200 405.600 ;
        RECT 538.200 399.600 540.000 406.800 ;
        RECT 566.550 406.050 567.450 427.950 ;
        RECT 571.500 419.400 573.300 431.400 ;
        RECT 577.800 425.400 579.600 431.400 ;
        RECT 592.800 425.400 594.600 431.400 ;
        RECT 571.800 413.100 573.000 419.400 ;
        RECT 578.400 418.500 579.600 425.400 ;
        RECT 573.900 417.600 579.600 418.500 ;
        RECT 573.900 416.700 575.850 417.600 ;
        RECT 574.950 413.100 575.850 416.700 ;
        RECT 589.950 415.950 592.050 421.050 ;
        RECT 593.400 416.100 594.600 425.400 ;
        RECT 610.500 419.400 612.300 431.400 ;
        RECT 628.800 430.500 636.600 431.400 ;
        RECT 628.800 419.400 630.600 430.500 ;
        RECT 595.950 415.950 598.050 418.050 ;
        RECT 610.950 416.100 612.150 419.400 ;
        RECT 631.800 418.500 633.600 429.600 ;
        RECT 634.800 420.600 636.600 430.500 ;
        RECT 640.800 420.600 642.600 431.400 ;
        RECT 634.800 419.700 642.600 420.600 ;
        RECT 655.500 419.400 657.300 431.400 ;
        RECT 676.800 425.400 678.600 431.400 ;
        RECT 631.800 417.600 635.850 418.500 ;
        RECT 634.950 416.100 635.850 417.600 ;
        RECT 655.950 416.100 657.150 419.400 ;
        RECT 590.100 414.150 591.900 414.900 ;
        RECT 578.100 413.100 579.900 413.850 ;
        RECT 568.950 409.950 574.050 412.050 ;
        RECT 575.100 408.900 575.850 413.100 ;
        RECT 592.950 412.950 595.050 415.050 ;
        RECT 596.100 414.150 597.900 414.900 ;
        RECT 605.100 413.100 606.900 413.850 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 611.100 413.100 612.150 416.100 ;
        RECT 613.950 412.950 616.050 415.050 ;
        RECT 629.100 413.100 630.900 413.850 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 635.100 413.100 635.850 416.100 ;
        RECT 637.950 412.950 640.050 415.050 ;
        RECT 641.100 413.100 642.750 413.850 ;
        RECT 650.100 413.100 651.900 413.850 ;
        RECT 652.950 412.950 655.050 415.050 ;
        RECT 656.100 413.100 657.150 416.100 ;
        RECT 673.950 415.950 676.050 418.050 ;
        RECT 677.400 416.100 678.600 425.400 ;
        RECT 694.500 419.400 696.300 431.400 ;
        RECT 706.950 424.950 709.050 427.050 ;
        RECT 694.950 416.100 696.150 419.400 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 674.100 414.150 675.900 414.900 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 680.100 414.150 681.900 414.900 ;
        RECT 689.100 413.100 690.900 413.850 ;
        RECT 691.800 412.950 694.050 415.050 ;
        RECT 695.100 413.100 696.150 416.100 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 577.950 409.950 580.050 412.050 ;
        RECT 557.400 402.600 558.600 405.900 ;
        RECT 565.950 403.950 568.050 406.050 ;
        RECT 571.800 405.600 573.000 408.900 ;
        RECT 574.950 408.300 575.850 408.900 ;
        RECT 573.900 407.400 575.850 408.300 ;
        RECT 593.400 407.700 594.600 411.900 ;
        RECT 604.800 409.950 607.050 412.050 ;
        RECT 608.100 411.150 609.900 411.900 ;
        RECT 610.950 409.950 613.050 412.050 ;
        RECT 614.100 411.150 615.900 411.900 ;
        RECT 628.950 409.950 631.050 412.050 ;
        RECT 632.250 411.150 633.900 411.900 ;
        RECT 634.950 409.950 637.050 412.050 ;
        RECT 638.100 411.150 639.750 411.900 ;
        RECT 640.950 409.950 643.050 412.050 ;
        RECT 649.950 409.950 652.050 412.050 ;
        RECT 653.100 411.150 654.900 411.900 ;
        RECT 655.950 409.950 658.050 412.050 ;
        RECT 659.100 411.150 660.900 411.900 ;
        RECT 611.850 408.750 613.050 408.900 ;
        RECT 611.850 407.700 615.600 408.750 ;
        RECT 573.900 406.500 579.000 407.400 ;
        RECT 556.800 399.600 558.600 402.600 ;
        RECT 571.500 399.600 573.300 405.600 ;
        RECT 577.800 402.600 579.000 406.500 ;
        RECT 591.000 406.800 594.600 407.700 ;
        RECT 577.800 399.600 579.600 402.600 ;
        RECT 591.000 399.600 592.800 406.800 ;
        RECT 605.400 404.700 613.200 406.050 ;
        RECT 605.400 399.600 607.200 404.700 ;
        RECT 611.400 399.600 613.200 404.700 ;
        RECT 614.400 405.600 615.600 407.700 ;
        RECT 636.000 405.600 637.050 408.900 ;
        RECT 656.850 408.750 658.050 408.900 ;
        RECT 656.850 407.700 660.600 408.750 ;
        RECT 677.400 407.700 678.600 411.900 ;
        RECT 688.800 409.950 691.050 412.050 ;
        RECT 692.100 411.150 693.900 411.900 ;
        RECT 694.950 409.950 697.200 412.050 ;
        RECT 698.100 411.150 699.900 411.900 ;
        RECT 704.550 409.050 705.450 412.950 ;
        RECT 695.850 408.750 697.050 408.900 ;
        RECT 695.850 407.700 699.600 408.750 ;
        RECT 614.400 399.600 616.200 405.600 ;
        RECT 636.000 399.600 637.800 405.600 ;
        RECT 650.400 404.700 658.200 406.050 ;
        RECT 650.400 399.600 652.200 404.700 ;
        RECT 656.400 399.600 658.200 404.700 ;
        RECT 659.400 405.600 660.600 407.700 ;
        RECT 675.000 406.800 678.600 407.700 ;
        RECT 659.400 399.600 661.200 405.600 ;
        RECT 675.000 399.600 676.800 406.800 ;
        RECT 689.400 404.700 697.200 406.050 ;
        RECT 689.400 399.600 691.200 404.700 ;
        RECT 695.400 399.600 697.200 404.700 ;
        RECT 698.400 405.600 699.600 407.700 ;
        RECT 703.950 406.950 706.050 409.050 ;
        RECT 707.550 406.050 708.450 424.950 ;
        RECT 716.700 419.400 718.500 431.400 ;
        RECT 731.400 424.200 733.200 430.200 ;
        RECT 716.850 416.100 718.050 419.400 ;
        RECT 732.300 419.100 733.200 424.200 ;
        RECT 738.900 420.900 740.700 430.200 ;
        RECT 758.400 425.400 760.200 431.400 ;
        RECT 738.900 420.000 741.000 420.900 ;
        RECT 732.300 418.200 738.450 419.100 ;
        RECT 712.950 412.950 715.050 415.050 ;
        RECT 716.850 413.100 717.900 416.100 ;
        RECT 737.250 415.500 738.450 418.200 ;
        RECT 740.100 416.100 741.000 420.000 ;
        RECT 754.800 415.950 757.050 418.050 ;
        RECT 758.400 416.100 759.600 425.400 ;
        RECT 775.800 419.400 777.600 431.400 ;
        RECT 784.950 427.950 787.050 430.050 ;
        RECT 760.950 415.950 763.050 418.050 ;
        RECT 718.950 412.950 721.050 415.050 ;
        RECT 722.100 413.100 723.900 413.850 ;
        RECT 734.100 413.100 735.900 413.850 ;
        RECT 737.250 413.700 738.900 415.500 ;
        RECT 713.100 411.150 714.900 411.900 ;
        RECT 715.950 409.950 718.050 412.050 ;
        RECT 719.100 411.150 720.900 411.900 ;
        RECT 731.100 411.150 732.900 411.900 ;
        RECT 733.950 409.950 736.200 412.050 ;
        RECT 715.950 408.750 717.150 408.900 ;
        RECT 713.400 407.700 717.150 408.750 ;
        RECT 737.250 408.000 738.450 413.700 ;
        RECT 739.950 412.950 742.050 415.050 ;
        RECT 755.100 414.150 756.900 414.900 ;
        RECT 743.100 413.100 744.900 413.850 ;
        RECT 757.950 412.950 760.200 415.050 ;
        RECT 761.100 414.150 762.900 414.900 ;
        RECT 776.400 413.100 777.600 419.400 ;
        RECT 698.400 399.600 700.200 405.600 ;
        RECT 706.950 403.950 709.050 406.050 ;
        RECT 713.400 405.600 714.600 407.700 ;
        RECT 732.150 407.100 738.450 408.000 ;
        RECT 712.800 399.600 714.600 405.600 ;
        RECT 715.800 404.700 723.600 406.050 ;
        RECT 715.800 399.600 717.600 404.700 ;
        RECT 721.800 399.600 723.600 404.700 ;
        RECT 732.150 403.800 733.200 407.100 ;
        RECT 740.100 406.200 741.000 411.900 ;
        RECT 758.400 407.700 759.600 411.900 ;
        RECT 772.950 409.950 778.050 412.050 ;
        RECT 779.100 411.150 780.900 411.900 ;
        RECT 758.400 406.800 762.000 407.700 ;
        RECT 731.400 400.800 733.200 403.800 ;
        RECT 738.900 405.300 741.000 406.200 ;
        RECT 738.900 400.800 740.700 405.300 ;
        RECT 760.200 399.600 762.000 406.800 ;
        RECT 776.400 405.600 777.600 408.900 ;
        RECT 785.550 406.050 786.450 427.950 ;
        RECT 790.800 419.400 792.600 431.400 ;
        RECT 808.800 425.400 810.600 431.400 ;
        RECT 799.950 421.950 802.050 424.050 ;
        RECT 791.400 413.100 792.600 419.400 ;
        RECT 790.950 409.950 793.050 412.050 ;
        RECT 794.100 411.150 795.900 411.900 ;
        RECT 775.800 399.600 777.600 405.600 ;
        RECT 784.950 403.950 787.050 406.050 ;
        RECT 791.400 405.600 792.600 408.900 ;
        RECT 790.800 399.600 792.600 405.600 ;
        RECT 800.550 403.050 801.450 421.950 ;
        RECT 805.950 415.950 808.050 418.050 ;
        RECT 809.400 416.100 810.600 425.400 ;
        RECT 824.400 425.400 826.200 431.400 ;
        RECT 842.400 425.400 844.200 431.400 ;
        RECT 820.950 415.950 823.050 418.050 ;
        RECT 824.400 416.100 825.600 425.400 ;
        RECT 832.950 421.950 835.050 424.050 ;
        RECT 826.950 415.950 829.050 418.050 ;
        RECT 806.100 414.150 807.900 414.900 ;
        RECT 808.950 412.950 811.050 415.050 ;
        RECT 812.100 414.150 813.900 414.900 ;
        RECT 821.100 414.150 822.900 414.900 ;
        RECT 823.800 412.950 826.050 415.050 ;
        RECT 827.100 414.150 828.900 414.900 ;
        RECT 833.550 412.050 834.450 421.950 ;
        RECT 839.100 413.100 840.900 413.850 ;
        RECT 809.400 407.700 810.600 411.900 ;
        RECT 807.000 406.800 810.600 407.700 ;
        RECT 824.400 407.700 825.600 411.900 ;
        RECT 832.950 409.950 835.050 412.050 ;
        RECT 838.950 409.950 841.050 412.050 ;
        RECT 842.400 408.300 843.450 425.400 ;
        RECT 849.000 419.400 850.800 431.400 ;
        RECT 844.950 412.950 847.050 415.050 ;
        RECT 849.000 413.100 850.050 419.400 ;
        RECT 845.100 411.150 846.900 411.900 ;
        RECT 847.950 411.450 850.050 412.050 ;
        RECT 847.950 410.550 855.450 411.450 ;
        RECT 847.950 409.950 850.050 410.550 ;
        RECT 824.400 406.800 828.000 407.700 ;
        RECT 799.800 400.950 801.900 403.050 ;
        RECT 807.000 399.600 808.800 406.800 ;
        RECT 826.200 399.600 828.000 406.800 ;
        RECT 839.400 407.100 846.900 408.300 ;
        RECT 839.400 399.600 841.200 407.100 ;
        RECT 845.100 406.500 846.900 407.100 ;
        RECT 847.950 405.600 848.850 408.900 ;
        RECT 846.900 403.800 848.850 405.600 ;
        RECT 846.900 399.600 848.700 403.800 ;
        RECT 854.550 403.050 855.450 410.550 ;
        RECT 853.950 400.950 856.050 403.050 ;
        RECT 14.100 387.000 15.900 395.400 ;
        RECT 34.200 391.050 36.000 395.400 ;
        RECT 49.950 391.950 52.050 394.050 ;
        RECT 34.200 389.400 39.600 391.050 ;
        RECT 11.700 385.350 15.900 387.000 ;
        RECT 38.700 386.100 39.600 389.400 ;
        RECT 46.800 385.950 48.900 388.050 ;
        RECT 11.700 380.100 12.600 385.350 ;
        RECT 14.100 383.100 15.900 383.850 ;
        RECT 20.100 383.100 21.900 383.850 ;
        RECT 29.100 383.100 30.900 383.850 ;
        RECT 31.950 382.950 34.200 385.050 ;
        RECT 35.100 383.100 36.900 383.850 ;
        RECT 37.950 382.950 43.050 385.050 ;
        RECT 13.950 379.950 16.050 382.050 ;
        RECT 19.950 379.950 22.050 382.050 ;
        RECT 28.800 379.950 31.050 382.050 ;
        RECT 32.100 381.150 33.900 381.900 ;
        RECT 34.950 379.950 37.200 382.050 ;
        RECT 7.950 376.950 13.050 379.050 ;
        RECT 16.950 376.950 19.050 379.050 ;
        RECT 11.700 370.800 12.600 375.900 ;
        RECT 17.100 375.150 18.900 375.900 ;
        RECT 38.700 375.600 39.600 381.900 ;
        RECT 47.550 376.050 48.450 385.950 ;
        RECT 50.550 385.050 51.450 391.950 ;
        RECT 56.100 387.000 57.900 395.400 ;
        RECT 53.700 385.350 57.900 387.000 ;
        RECT 81.000 389.400 82.800 395.400 ;
        RECT 102.000 391.050 103.800 395.400 ;
        RECT 118.800 392.400 120.600 395.400 ;
        RECT 98.400 389.400 103.800 391.050 ;
        RECT 81.000 386.100 82.050 389.400 ;
        RECT 98.400 386.100 99.300 389.400 ;
        RECT 112.950 385.950 115.050 388.050 ;
        RECT 50.100 382.950 52.200 385.050 ;
        RECT 53.700 380.100 54.600 385.350 ;
        RECT 56.100 383.100 57.900 383.850 ;
        RECT 62.100 383.100 63.900 383.850 ;
        RECT 73.950 382.950 76.050 385.050 ;
        RECT 77.250 383.100 78.900 383.850 ;
        RECT 79.950 382.950 82.050 385.050 ;
        RECT 83.100 383.100 84.750 383.850 ;
        RECT 85.950 382.950 88.050 385.050 ;
        RECT 91.950 384.450 96.000 385.050 ;
        RECT 97.950 384.450 100.050 385.050 ;
        RECT 91.950 383.550 100.050 384.450 ;
        RECT 91.950 382.950 96.000 383.550 ;
        RECT 97.950 382.950 100.050 383.550 ;
        RECT 101.100 383.100 102.900 383.850 ;
        RECT 103.950 382.950 106.050 385.050 ;
        RECT 107.100 383.100 108.900 383.850 ;
        RECT 55.950 379.950 58.050 382.050 ;
        RECT 61.950 379.950 64.050 382.050 ;
        RECT 74.100 381.150 75.900 381.900 ;
        RECT 76.950 379.950 79.050 382.050 ;
        RECT 49.950 376.950 55.050 379.050 ;
        RECT 58.950 376.950 61.050 379.050 ;
        RECT 80.100 378.900 80.850 381.900 ;
        RECT 82.950 379.950 85.050 382.050 ;
        RECT 86.100 381.150 87.750 381.900 ;
        RECT 79.950 377.400 80.850 378.900 ;
        RECT 76.800 376.500 80.850 377.400 ;
        RECT 29.400 374.700 37.200 375.600 ;
        RECT 11.700 369.900 18.300 370.800 ;
        RECT 11.700 369.600 12.600 369.900 ;
        RECT 10.800 363.600 12.600 369.600 ;
        RECT 16.800 369.600 18.300 369.900 ;
        RECT 16.800 363.600 18.600 369.600 ;
        RECT 29.400 363.600 31.200 374.700 ;
        RECT 35.400 363.600 37.200 374.700 ;
        RECT 38.400 363.600 40.200 375.600 ;
        RECT 46.950 373.950 49.050 376.050 ;
        RECT 53.700 370.800 54.600 375.900 ;
        RECT 59.100 375.150 60.900 375.900 ;
        RECT 53.700 369.900 60.300 370.800 ;
        RECT 53.700 369.600 54.600 369.900 ;
        RECT 52.800 363.600 54.600 369.600 ;
        RECT 58.800 369.600 60.300 369.900 ;
        RECT 58.800 363.600 60.600 369.600 ;
        RECT 73.800 364.500 75.600 375.600 ;
        RECT 76.800 365.400 78.600 376.500 ;
        RECT 98.400 375.600 99.300 381.900 ;
        RECT 100.950 379.950 103.050 382.050 ;
        RECT 104.100 381.150 105.900 381.900 ;
        RECT 106.950 379.950 109.050 382.050 ;
        RECT 113.550 381.450 114.450 385.950 ;
        RECT 119.400 383.100 120.600 392.400 ;
        RECT 129.000 390.450 133.050 391.050 ;
        RECT 128.550 388.950 133.050 390.450 ;
        RECT 121.950 385.950 124.050 388.050 ;
        RECT 122.100 384.150 123.900 384.900 ;
        RECT 128.550 382.050 129.450 388.950 ;
        RECT 135.000 388.200 136.800 395.400 ;
        RECT 135.000 387.300 138.600 388.200 ;
        RECT 137.400 383.100 138.600 387.300 ;
        RECT 155.100 387.000 156.900 395.400 ;
        RECT 173.400 392.400 175.200 395.400 ;
        RECT 173.400 389.100 174.600 392.400 ;
        RECT 181.950 391.950 184.050 394.050 ;
        RECT 152.700 385.350 156.900 387.000 ;
        RECT 172.950 385.950 175.050 388.050 ;
        RECT 118.950 381.450 121.050 382.050 ;
        RECT 113.550 380.550 121.050 381.450 ;
        RECT 79.800 374.400 87.600 375.300 ;
        RECT 79.800 364.500 81.600 374.400 ;
        RECT 73.800 363.600 81.600 364.500 ;
        RECT 85.800 363.600 87.600 374.400 ;
        RECT 97.800 363.600 99.600 375.600 ;
        RECT 100.800 374.700 108.600 375.600 ;
        RECT 100.800 363.600 102.600 374.700 ;
        RECT 106.800 363.600 108.600 374.700 ;
        RECT 113.550 367.050 114.450 380.550 ;
        RECT 118.950 379.950 121.050 380.550 ;
        RECT 127.950 379.950 130.050 382.050 ;
        RECT 134.100 380.100 135.900 380.850 ;
        RECT 136.950 379.950 139.050 382.050 ;
        RECT 140.100 380.100 141.900 380.850 ;
        RECT 152.700 380.100 153.600 385.350 ;
        RECT 155.100 383.100 156.900 383.850 ;
        RECT 161.100 383.100 162.900 383.850 ;
        RECT 169.950 382.950 172.050 385.050 ;
        RECT 154.950 379.950 157.050 382.050 ;
        RECT 160.950 379.950 163.050 382.050 ;
        RECT 173.700 381.900 174.900 384.900 ;
        RECT 175.950 382.950 178.200 385.050 ;
        RECT 170.100 381.150 171.900 381.900 ;
        RECT 119.400 369.600 120.600 378.900 ;
        RECT 130.950 376.950 136.050 379.050 ;
        RECT 137.400 369.600 138.600 378.900 ;
        RECT 139.950 376.950 142.050 379.050 ;
        RECT 151.950 378.450 154.050 379.050 ;
        RECT 146.550 377.550 154.050 378.450 ;
        RECT 112.950 364.950 115.050 367.050 ;
        RECT 118.800 363.600 120.600 369.600 ;
        RECT 136.800 363.600 138.600 369.600 ;
        RECT 146.550 367.050 147.450 377.550 ;
        RECT 151.950 376.950 154.050 377.550 ;
        RECT 157.950 376.950 160.050 379.050 ;
        RECT 173.700 376.650 175.050 381.900 ;
        RECT 176.100 381.150 177.900 381.900 ;
        RECT 152.700 370.800 153.600 375.900 ;
        RECT 158.100 375.150 159.900 375.900 ;
        RECT 173.700 375.600 176.400 376.650 ;
        RECT 152.700 369.900 159.300 370.800 ;
        RECT 152.700 369.600 153.600 369.900 ;
        RECT 145.950 364.950 148.050 367.050 ;
        RECT 151.800 363.600 153.600 369.600 ;
        RECT 157.800 369.600 159.300 369.900 ;
        RECT 157.800 363.600 159.600 369.600 ;
        RECT 174.600 363.600 176.400 375.600 ;
        RECT 182.550 367.050 183.450 391.950 ;
        RECT 192.000 388.200 193.800 395.400 ;
        RECT 208.800 392.400 210.600 395.400 ;
        RECT 223.800 392.400 225.600 395.400 ;
        RECT 192.000 387.300 195.600 388.200 ;
        RECT 194.400 383.100 195.600 387.300 ;
        RECT 209.400 383.100 210.600 392.400 ;
        RECT 211.950 385.950 214.050 388.050 ;
        RECT 212.100 384.150 213.900 384.900 ;
        RECT 224.400 383.100 225.600 392.400 ;
        RECT 226.950 385.950 229.050 388.050 ;
        RECT 242.100 387.000 243.900 395.400 ;
        RECT 239.700 385.350 243.900 387.000 ;
        RECT 267.000 389.400 268.800 395.400 ;
        RECT 283.800 392.400 285.600 395.400 ;
        RECT 267.000 386.100 268.050 389.400 ;
        RECT 227.100 384.150 228.900 384.900 ;
        RECT 191.100 380.100 192.900 380.850 ;
        RECT 193.950 379.950 196.050 382.050 ;
        RECT 197.100 380.100 198.900 380.850 ;
        RECT 208.950 379.950 214.050 382.050 ;
        RECT 223.950 379.950 226.050 382.050 ;
        RECT 239.700 380.100 240.600 385.350 ;
        RECT 242.100 383.100 243.900 383.850 ;
        RECT 248.100 383.100 249.900 383.850 ;
        RECT 259.950 382.950 262.050 385.050 ;
        RECT 263.250 383.100 264.900 383.850 ;
        RECT 265.950 382.950 268.200 385.050 ;
        RECT 269.100 383.100 270.750 383.850 ;
        RECT 271.950 382.950 274.050 385.050 ;
        RECT 284.400 383.100 285.600 392.400 ;
        RECT 286.950 385.950 289.050 388.050 ;
        RECT 302.100 387.000 303.900 395.400 ;
        RECT 317.400 390.300 319.200 395.400 ;
        RECT 323.400 390.300 325.200 395.400 ;
        RECT 317.400 388.950 325.200 390.300 ;
        RECT 326.400 389.400 328.200 395.400 ;
        RECT 342.300 391.200 344.100 395.400 ;
        RECT 342.150 389.400 344.100 391.200 ;
        RECT 326.400 387.300 327.600 389.400 ;
        RECT 299.700 385.350 303.900 387.000 ;
        RECT 323.850 386.250 327.600 387.300 ;
        RECT 323.850 386.100 325.050 386.250 ;
        RECT 342.150 386.100 343.050 389.400 ;
        RECT 344.100 387.900 345.900 388.500 ;
        RECT 349.800 387.900 351.600 395.400 ;
        RECT 355.950 391.950 358.050 394.050 ;
        RECT 344.100 386.700 351.600 387.900 ;
        RECT 287.100 384.150 288.900 384.900 ;
        RECT 241.950 379.950 244.050 382.050 ;
        RECT 247.950 379.950 250.050 382.050 ;
        RECT 260.100 381.150 261.900 381.900 ;
        RECT 262.950 379.950 265.050 382.050 ;
        RECT 190.950 376.950 193.050 379.050 ;
        RECT 194.400 369.600 195.600 378.900 ;
        RECT 196.950 376.950 199.050 379.050 ;
        RECT 209.400 369.600 210.600 378.900 ;
        RECT 224.400 369.600 225.600 378.900 ;
        RECT 232.950 378.450 237.000 379.050 ;
        RECT 238.950 378.450 241.050 379.050 ;
        RECT 232.950 377.550 241.050 378.450 ;
        RECT 232.950 376.950 237.000 377.550 ;
        RECT 238.950 376.950 241.050 377.550 ;
        RECT 244.950 376.950 247.050 379.050 ;
        RECT 266.100 378.900 266.850 381.900 ;
        RECT 268.950 379.950 271.050 382.050 ;
        RECT 272.100 381.150 273.750 381.900 ;
        RECT 283.950 381.450 286.050 382.050 ;
        RECT 278.550 380.550 286.050 381.450 ;
        RECT 265.950 377.400 266.850 378.900 ;
        RECT 262.800 376.500 266.850 377.400 ;
        RECT 239.700 370.800 240.600 375.900 ;
        RECT 245.100 375.150 246.900 375.900 ;
        RECT 239.700 369.900 246.300 370.800 ;
        RECT 239.700 369.600 240.600 369.900 ;
        RECT 181.950 364.950 184.050 367.050 ;
        RECT 193.800 363.600 195.600 369.600 ;
        RECT 208.800 363.600 210.600 369.600 ;
        RECT 223.800 363.600 225.600 369.600 ;
        RECT 238.800 363.600 240.600 369.600 ;
        RECT 244.800 369.600 246.300 369.900 ;
        RECT 244.800 363.600 246.600 369.600 ;
        RECT 259.800 364.500 261.600 375.600 ;
        RECT 262.800 365.400 264.600 376.500 ;
        RECT 265.800 374.400 273.600 375.300 ;
        RECT 265.800 364.500 267.600 374.400 ;
        RECT 259.800 363.600 267.600 364.500 ;
        RECT 271.800 363.600 273.600 374.400 ;
        RECT 278.550 370.050 279.450 380.550 ;
        RECT 283.950 379.950 286.050 380.550 ;
        RECT 299.700 380.100 300.600 385.350 ;
        RECT 302.100 383.100 303.900 383.850 ;
        RECT 308.100 383.100 309.900 383.850 ;
        RECT 316.950 382.950 319.050 385.050 ;
        RECT 320.100 383.100 321.900 383.850 ;
        RECT 322.800 382.950 325.050 385.050 ;
        RECT 326.100 383.100 327.900 383.850 ;
        RECT 337.950 382.950 343.050 385.050 ;
        RECT 344.100 383.100 345.900 383.850 ;
        RECT 301.950 379.950 304.050 382.050 ;
        RECT 307.950 379.950 310.050 382.050 ;
        RECT 317.100 381.150 318.900 381.900 ;
        RECT 319.950 379.950 322.050 382.050 ;
        RECT 277.950 367.950 280.050 370.050 ;
        RECT 284.400 369.600 285.600 378.900 ;
        RECT 298.950 378.450 301.050 379.050 ;
        RECT 283.800 363.600 285.600 369.600 ;
        RECT 293.550 377.550 301.050 378.450 ;
        RECT 293.550 367.050 294.450 377.550 ;
        RECT 298.950 376.950 301.050 377.550 ;
        RECT 304.950 376.950 307.050 379.050 ;
        RECT 323.100 378.900 324.150 381.900 ;
        RECT 325.950 379.950 328.200 382.050 ;
        RECT 299.700 370.800 300.600 375.900 ;
        RECT 305.100 375.150 306.900 375.900 ;
        RECT 322.950 375.600 324.150 378.900 ;
        RECT 340.950 375.600 342.000 381.900 ;
        RECT 343.950 379.950 346.050 382.050 ;
        RECT 299.700 369.900 306.300 370.800 ;
        RECT 299.700 369.600 300.600 369.900 ;
        RECT 292.950 364.950 295.050 367.050 ;
        RECT 298.800 363.600 300.600 369.600 ;
        RECT 304.800 369.600 306.300 369.900 ;
        RECT 304.800 363.600 306.600 369.600 ;
        RECT 322.500 363.600 324.300 375.600 ;
        RECT 340.200 363.600 342.000 375.600 ;
        RECT 347.550 369.600 348.600 386.700 ;
        RECT 349.950 382.950 352.050 385.050 ;
        RECT 356.550 384.450 357.450 391.950 ;
        RECT 361.500 389.400 363.300 395.400 ;
        RECT 367.800 392.400 369.600 395.400 ;
        RECT 361.800 386.100 363.000 389.400 ;
        RECT 367.800 388.500 369.000 392.400 ;
        RECT 363.900 387.600 369.000 388.500 ;
        RECT 377.400 387.900 379.200 395.400 ;
        RECT 384.900 391.200 386.700 395.400 ;
        RECT 384.900 389.400 386.850 391.200 ;
        RECT 400.500 389.400 402.300 395.400 ;
        RECT 406.800 392.400 408.600 395.400 ;
        RECT 419.400 392.400 421.200 395.400 ;
        RECT 383.100 387.900 384.900 388.500 ;
        RECT 363.900 386.700 365.850 387.600 ;
        RECT 377.400 386.700 384.900 387.900 ;
        RECT 364.950 386.100 365.850 386.700 ;
        RECT 361.950 384.450 364.050 385.050 ;
        RECT 356.550 383.550 364.050 384.450 ;
        RECT 361.950 382.950 364.050 383.550 ;
        RECT 365.100 381.900 365.850 386.100 ;
        RECT 367.950 382.950 370.050 385.050 ;
        RECT 376.950 382.950 379.050 385.050 ;
        RECT 350.100 381.150 351.900 381.900 ;
        RECT 361.800 375.600 363.000 381.900 ;
        RECT 364.950 378.300 365.850 381.900 ;
        RECT 368.100 381.150 369.900 381.900 ;
        RECT 377.100 381.150 378.900 381.900 ;
        RECT 363.900 377.400 365.850 378.300 ;
        RECT 363.900 376.500 369.600 377.400 ;
        RECT 346.800 363.600 348.600 369.600 ;
        RECT 361.500 363.600 363.300 375.600 ;
        RECT 368.400 369.600 369.600 376.500 ;
        RECT 367.800 363.600 369.600 369.600 ;
        RECT 380.400 369.600 381.450 386.700 ;
        RECT 385.950 386.100 386.850 389.400 ;
        RECT 400.800 386.100 402.000 389.400 ;
        RECT 406.800 388.500 408.000 392.400 ;
        RECT 402.900 387.600 408.000 388.500 ;
        RECT 402.900 386.700 404.850 387.600 ;
        RECT 403.950 386.100 404.850 386.700 ;
        RECT 383.100 383.100 384.900 383.850 ;
        RECT 385.950 382.950 388.050 385.050 ;
        RECT 382.950 379.950 385.050 382.050 ;
        RECT 404.100 381.900 404.850 386.100 ;
        RECT 412.950 385.950 418.050 388.050 ;
        RECT 406.950 382.950 409.050 385.050 ;
        RECT 416.100 384.150 417.900 384.900 ;
        RECT 419.400 383.100 420.600 392.400 ;
        RECT 424.950 391.950 427.050 394.050 ;
        RECT 387.000 375.600 388.050 381.900 ;
        RECT 400.800 375.600 402.000 381.900 ;
        RECT 403.950 378.300 404.850 381.900 ;
        RECT 407.100 381.150 408.900 381.900 ;
        RECT 418.950 379.950 424.050 382.050 ;
        RECT 402.900 377.400 404.850 378.300 ;
        RECT 402.900 376.500 408.600 377.400 ;
        RECT 380.400 363.600 382.200 369.600 ;
        RECT 387.000 363.600 388.800 375.600 ;
        RECT 400.500 363.600 402.300 375.600 ;
        RECT 407.400 369.600 408.600 376.500 ;
        RECT 406.800 363.600 408.600 369.600 ;
        RECT 419.400 369.600 420.600 378.900 ;
        RECT 425.550 370.050 426.450 391.950 ;
        RECT 436.200 389.400 438.000 395.400 ;
        RECT 436.950 386.100 438.000 389.400 ;
        RECT 449.550 389.400 451.350 395.400 ;
        RECT 457.650 392.400 459.450 395.400 ;
        RECT 465.450 392.400 467.250 395.400 ;
        RECT 473.250 393.300 475.050 395.400 ;
        RECT 473.250 392.400 477.000 393.300 ;
        RECT 457.650 391.500 458.700 392.400 ;
        RECT 454.950 390.300 458.700 391.500 ;
        RECT 466.200 390.600 467.250 392.400 ;
        RECT 475.950 391.500 477.000 392.400 ;
        RECT 454.950 389.400 457.050 390.300 ;
        RECT 449.550 385.050 450.750 389.400 ;
        RECT 462.150 388.200 463.950 390.000 ;
        RECT 466.200 389.550 471.150 390.600 ;
        RECT 469.350 388.800 471.150 389.550 ;
        RECT 472.650 388.800 474.450 390.600 ;
        RECT 475.950 389.400 478.050 391.500 ;
        RECT 481.050 389.400 482.850 395.400 ;
        RECT 463.050 387.900 463.950 388.200 ;
        RECT 473.100 387.900 474.150 388.800 ;
        RECT 463.050 387.000 474.150 387.900 ;
        RECT 463.050 386.100 463.950 387.000 ;
        RECT 473.100 385.800 474.150 387.000 ;
        RECT 430.950 382.950 433.050 385.050 ;
        RECT 434.250 383.100 435.900 383.850 ;
        RECT 436.800 382.950 439.050 385.050 ;
        RECT 440.100 383.100 441.750 383.850 ;
        RECT 442.950 382.950 445.050 385.050 ;
        RECT 449.550 382.950 450.900 385.050 ;
        RECT 451.950 382.950 454.050 385.050 ;
        RECT 455.100 383.250 455.850 385.050 ;
        RECT 463.950 382.950 466.050 385.050 ;
        RECT 469.950 382.950 472.050 385.050 ;
        RECT 473.100 384.600 480.000 385.800 ;
        RECT 473.100 384.000 474.900 384.600 ;
        RECT 479.100 383.850 480.000 384.600 ;
        RECT 476.100 383.100 477.900 383.700 ;
        RECT 431.250 381.150 432.900 381.900 ;
        RECT 433.800 379.950 436.050 382.050 ;
        RECT 438.150 378.900 438.900 381.900 ;
        RECT 439.950 379.950 442.200 382.050 ;
        RECT 443.100 381.150 444.900 381.900 ;
        RECT 438.150 377.400 439.050 378.900 ;
        RECT 438.150 376.500 442.200 377.400 ;
        RECT 431.400 374.400 439.200 375.300 ;
        RECT 419.400 363.600 421.200 369.600 ;
        RECT 424.950 367.950 427.050 370.050 ;
        RECT 431.400 363.600 433.200 374.400 ;
        RECT 437.400 364.500 439.200 374.400 ;
        RECT 440.400 365.400 442.200 376.500 ;
        RECT 449.550 375.600 450.750 382.950 ;
        RECT 473.100 382.200 477.900 383.100 ;
        RECT 476.100 381.900 477.900 382.200 ;
        RECT 479.100 382.050 480.900 383.850 ;
        RECT 451.950 377.400 453.750 379.200 ;
        RECT 452.850 376.200 457.050 377.400 ;
        RECT 463.050 376.200 463.950 381.900 ;
        RECT 471.750 377.100 473.550 377.400 ;
        RECT 443.400 364.500 445.200 375.600 ;
        RECT 437.400 363.600 445.200 364.500 ;
        RECT 449.550 363.600 451.350 375.600 ;
        RECT 454.950 375.300 457.050 376.200 ;
        RECT 457.950 375.300 463.950 376.200 ;
        RECT 465.150 376.800 473.550 377.100 ;
        RECT 481.950 376.800 482.850 389.400 ;
        RECT 491.400 390.300 493.200 395.400 ;
        RECT 497.400 390.300 499.200 395.400 ;
        RECT 491.400 388.950 499.200 390.300 ;
        RECT 500.400 389.400 502.200 395.400 ;
        RECT 505.950 391.950 508.050 394.050 ;
        RECT 500.400 387.300 501.600 389.400 ;
        RECT 497.850 386.250 501.600 387.300 ;
        RECT 497.850 386.100 499.050 386.250 ;
        RECT 490.950 384.450 493.050 385.050 ;
        RECT 465.150 376.200 482.850 376.800 ;
        RECT 457.950 374.400 458.850 375.300 ;
        RECT 456.150 372.600 458.850 374.400 ;
        RECT 459.750 374.100 461.550 374.400 ;
        RECT 465.150 374.100 466.050 376.200 ;
        RECT 471.750 375.600 482.850 376.200 ;
        RECT 485.550 383.550 493.050 384.450 ;
        RECT 485.550 376.050 486.450 383.550 ;
        RECT 490.950 382.950 493.050 383.550 ;
        RECT 494.100 383.100 495.900 383.850 ;
        RECT 496.950 382.950 499.200 385.050 ;
        RECT 500.100 383.100 501.900 383.850 ;
        RECT 506.550 382.050 507.450 391.950 ;
        RECT 517.200 391.050 519.000 395.400 ;
        RECT 517.200 389.400 522.600 391.050 ;
        RECT 521.700 386.100 522.600 389.400 ;
        RECT 526.950 388.950 529.050 391.050 ;
        RECT 535.800 389.400 537.600 395.400 ;
        RECT 512.100 383.100 513.900 383.850 ;
        RECT 514.950 382.950 517.050 385.050 ;
        RECT 520.950 384.450 523.050 385.050 ;
        RECT 527.550 384.450 528.450 388.950 ;
        RECT 529.950 385.950 532.050 388.050 ;
        RECT 536.400 387.300 537.600 389.400 ;
        RECT 538.800 390.300 540.600 395.400 ;
        RECT 544.800 390.300 546.600 395.400 ;
        RECT 538.800 388.950 546.600 390.300 ;
        RECT 556.800 389.400 558.600 395.400 ;
        RECT 557.400 387.300 558.600 389.400 ;
        RECT 559.800 390.300 561.600 395.400 ;
        RECT 565.800 390.300 567.600 395.400 ;
        RECT 559.800 388.950 567.600 390.300 ;
        RECT 582.300 389.700 584.100 394.200 ;
        RECT 582.000 388.800 584.100 389.700 ;
        RECT 589.800 391.200 591.600 394.200 ;
        RECT 536.400 386.250 540.150 387.300 ;
        RECT 557.400 386.250 561.150 387.300 ;
        RECT 538.950 386.100 540.150 386.250 ;
        RECT 559.950 386.100 561.150 386.250 ;
        RECT 518.100 383.100 519.900 383.850 ;
        RECT 520.950 383.550 528.450 384.450 ;
        RECT 520.950 382.950 523.050 383.550 ;
        RECT 530.550 382.050 531.450 385.950 ;
        RECT 536.100 383.100 537.900 383.850 ;
        RECT 538.950 382.950 541.050 385.050 ;
        RECT 542.100 383.100 543.900 383.850 ;
        RECT 544.950 382.950 547.050 385.050 ;
        RECT 550.950 382.950 553.050 385.050 ;
        RECT 557.100 383.100 558.900 383.850 ;
        RECT 559.950 382.950 562.050 385.050 ;
        RECT 565.950 384.450 568.050 385.050 ;
        RECT 563.100 383.100 564.900 383.850 ;
        RECT 565.950 383.550 573.450 384.450 ;
        RECT 565.950 382.950 568.050 383.550 ;
        RECT 491.100 381.150 492.900 381.900 ;
        RECT 493.950 379.950 496.050 382.050 ;
        RECT 497.100 378.900 498.150 381.900 ;
        RECT 499.950 379.950 502.050 382.050 ;
        RECT 505.950 379.950 508.050 382.050 ;
        RECT 511.800 379.950 514.050 382.050 ;
        RECT 515.100 381.150 516.900 381.900 ;
        RECT 517.950 379.950 520.050 382.050 ;
        RECT 459.750 373.200 466.050 374.100 ;
        RECT 466.950 374.700 468.750 375.300 ;
        RECT 466.950 373.500 474.450 374.700 ;
        RECT 459.750 372.600 461.550 373.200 ;
        RECT 473.250 372.600 474.450 373.500 ;
        RECT 454.950 369.600 458.850 371.700 ;
        RECT 463.950 371.550 465.750 372.300 ;
        RECT 468.750 371.550 470.550 372.300 ;
        RECT 463.950 370.500 470.550 371.550 ;
        RECT 473.250 370.500 478.050 372.600 ;
        RECT 457.050 363.600 458.850 369.600 ;
        RECT 464.850 363.600 466.650 370.500 ;
        RECT 473.250 369.600 474.450 370.500 ;
        RECT 472.650 363.600 474.450 369.600 ;
        RECT 481.050 363.600 482.850 375.600 ;
        RECT 484.950 373.950 487.050 376.050 ;
        RECT 496.950 375.600 498.150 378.900 ;
        RECT 496.500 363.600 498.300 375.600 ;
        RECT 506.550 370.050 507.450 379.950 ;
        RECT 521.700 375.600 522.600 381.900 ;
        RECT 529.950 379.950 532.050 382.050 ;
        RECT 535.950 379.950 538.050 382.050 ;
        RECT 539.850 378.900 540.900 381.900 ;
        RECT 541.950 379.950 544.050 382.050 ;
        RECT 545.100 381.150 546.900 381.900 ;
        RECT 551.550 379.050 552.450 382.950 ;
        RECT 556.950 379.950 559.050 382.050 ;
        RECT 539.850 375.600 541.050 378.900 ;
        RECT 550.950 376.950 553.050 379.050 ;
        RECT 560.850 378.900 561.900 381.900 ;
        RECT 566.100 381.150 567.900 381.900 ;
        RECT 560.850 375.600 562.050 378.900 ;
        RECT 512.400 374.700 520.200 375.600 ;
        RECT 505.950 367.950 508.050 370.050 ;
        RECT 512.400 363.600 514.200 374.700 ;
        RECT 518.400 363.600 520.200 374.700 ;
        RECT 521.400 363.600 523.200 375.600 ;
        RECT 539.700 363.600 541.500 375.600 ;
        RECT 560.700 363.600 562.500 375.600 ;
        RECT 572.550 370.050 573.450 383.550 ;
        RECT 577.950 382.950 580.050 385.050 ;
        RECT 582.000 383.100 582.900 388.800 ;
        RECT 589.800 387.900 590.850 391.200 ;
        RECT 604.200 388.200 606.000 395.400 ;
        RECT 611.100 391.950 613.200 394.050 ;
        RECT 584.550 387.000 590.850 387.900 ;
        RECT 602.400 387.300 606.000 388.200 ;
        RECT 578.100 381.150 579.900 381.900 ;
        RECT 580.950 379.950 583.050 382.050 ;
        RECT 584.550 381.300 585.750 387.000 ;
        RECT 586.950 382.950 589.050 385.050 ;
        RECT 590.100 383.100 591.900 383.850 ;
        RECT 602.400 383.100 603.600 387.300 ;
        RECT 584.100 379.500 585.750 381.300 ;
        RECT 587.100 381.150 588.900 381.900 ;
        RECT 589.950 379.950 592.050 382.050 ;
        RECT 599.100 380.100 600.900 380.850 ;
        RECT 601.950 379.950 604.050 382.050 ;
        RECT 605.100 380.100 606.900 380.850 ;
        RECT 582.000 375.000 582.900 378.900 ;
        RECT 584.550 376.800 585.750 379.500 ;
        RECT 611.550 379.050 612.450 391.950 ;
        RECT 617.400 390.300 619.200 395.400 ;
        RECT 623.400 390.300 625.200 395.400 ;
        RECT 617.400 388.950 625.200 390.300 ;
        RECT 626.400 389.400 628.200 395.400 ;
        RECT 643.200 389.400 645.000 395.400 ;
        RECT 626.400 387.300 627.600 389.400 ;
        RECT 623.850 386.250 627.600 387.300 ;
        RECT 623.850 386.100 625.050 386.250 ;
        RECT 643.950 386.100 645.000 389.400 ;
        RECT 668.100 387.000 669.900 395.400 ;
        RECT 683.400 392.400 685.200 395.400 ;
        RECT 684.000 388.500 685.200 392.400 ;
        RECT 689.700 389.400 691.500 395.400 ;
        RECT 684.000 387.600 689.100 388.500 ;
        RECT 665.700 385.350 669.900 387.000 ;
        RECT 687.150 386.700 689.100 387.600 ;
        RECT 687.150 386.100 688.050 386.700 ;
        RECT 690.000 386.100 691.200 389.400 ;
        RECT 705.000 388.200 706.800 395.400 ;
        RECT 722.400 392.400 724.200 395.400 ;
        RECT 736.800 392.400 738.600 395.400 ;
        RECT 752.400 392.400 754.200 395.400 ;
        RECT 705.000 387.300 708.600 388.200 ;
        RECT 616.800 382.950 619.050 385.050 ;
        RECT 620.100 383.100 621.900 383.850 ;
        RECT 622.950 382.950 625.200 385.050 ;
        RECT 626.100 383.100 627.900 383.850 ;
        RECT 631.800 382.950 633.900 385.050 ;
        RECT 637.950 382.950 640.050 385.050 ;
        RECT 641.250 383.100 642.900 383.850 ;
        RECT 643.950 382.950 646.050 385.050 ;
        RECT 647.100 383.100 648.750 383.850 ;
        RECT 649.950 382.950 652.050 385.050 ;
        RECT 658.950 382.950 661.050 385.050 ;
        RECT 617.100 381.150 618.900 381.900 ;
        RECT 619.950 379.950 622.050 382.050 ;
        RECT 598.950 376.950 601.050 379.050 ;
        RECT 584.550 375.900 590.700 376.800 ;
        RECT 582.000 374.100 584.100 375.000 ;
        RECT 571.950 367.950 574.050 370.050 ;
        RECT 582.300 364.800 584.100 374.100 ;
        RECT 589.800 370.800 590.700 375.900 ;
        RECT 589.800 364.800 591.600 370.800 ;
        RECT 602.400 369.600 603.600 378.900 ;
        RECT 604.950 376.950 607.050 379.050 ;
        RECT 610.950 376.950 613.050 379.050 ;
        RECT 623.100 378.900 624.150 381.900 ;
        RECT 625.950 379.950 628.050 382.050 ;
        RECT 622.950 375.600 624.150 378.900 ;
        RECT 602.400 363.600 604.200 369.600 ;
        RECT 622.500 363.600 624.300 375.600 ;
        RECT 632.550 367.050 633.450 382.950 ;
        RECT 638.250 381.150 639.900 381.900 ;
        RECT 640.950 379.950 643.050 382.050 ;
        RECT 645.150 378.900 645.900 381.900 ;
        RECT 646.950 379.950 649.200 382.050 ;
        RECT 650.100 381.150 651.900 381.900 ;
        RECT 645.150 377.400 646.050 378.900 ;
        RECT 659.550 378.450 660.450 382.950 ;
        RECT 665.700 380.100 666.600 385.350 ;
        RECT 668.100 383.100 669.900 383.850 ;
        RECT 674.100 383.100 675.900 383.850 ;
        RECT 679.950 382.950 685.050 385.050 ;
        RECT 667.950 379.950 670.050 382.050 ;
        RECT 673.950 379.950 676.050 382.050 ;
        RECT 687.150 381.900 687.900 386.100 ;
        RECT 688.950 384.450 691.050 385.050 ;
        RECT 688.950 383.550 696.450 384.450 ;
        RECT 688.950 382.950 691.050 383.550 ;
        RECT 683.100 381.150 684.900 381.900 ;
        RECT 664.950 378.450 667.050 379.050 ;
        RECT 659.550 377.550 667.050 378.450 ;
        RECT 645.150 376.500 649.200 377.400 ;
        RECT 664.950 376.950 667.050 377.550 ;
        RECT 670.950 376.950 673.050 379.050 ;
        RECT 687.150 378.300 688.050 381.900 ;
        RECT 687.150 377.400 689.100 378.300 ;
        RECT 638.400 374.400 646.200 375.300 ;
        RECT 631.950 364.950 634.050 367.050 ;
        RECT 638.400 363.600 640.200 374.400 ;
        RECT 644.400 364.500 646.200 374.400 ;
        RECT 647.400 365.400 649.200 376.500 ;
        RECT 683.400 376.500 689.100 377.400 ;
        RECT 650.400 364.500 652.200 375.600 ;
        RECT 665.700 370.800 666.600 375.900 ;
        RECT 671.100 375.150 672.900 375.900 ;
        RECT 665.700 369.900 672.300 370.800 ;
        RECT 665.700 369.600 666.600 369.900 ;
        RECT 644.400 363.600 652.200 364.500 ;
        RECT 664.800 363.600 666.600 369.600 ;
        RECT 670.800 369.600 672.300 369.900 ;
        RECT 683.400 369.600 684.600 376.500 ;
        RECT 690.000 375.600 691.200 381.900 ;
        RECT 670.800 363.600 672.600 369.600 ;
        RECT 683.400 363.600 685.200 369.600 ;
        RECT 689.700 363.600 691.500 375.600 ;
        RECT 695.550 367.050 696.450 383.550 ;
        RECT 707.400 383.100 708.600 387.300 ;
        RECT 718.950 385.950 721.050 388.050 ;
        RECT 719.100 384.150 720.900 384.900 ;
        RECT 722.400 383.100 723.600 392.400 ;
        RECT 737.400 383.100 738.600 392.400 ;
        RECT 753.000 388.500 754.200 392.400 ;
        RECT 758.700 389.400 760.500 395.400 ;
        RECT 739.950 385.950 742.050 388.050 ;
        RECT 753.000 387.600 758.100 388.500 ;
        RECT 756.150 386.700 758.100 387.600 ;
        RECT 756.150 386.100 757.050 386.700 ;
        RECT 759.000 386.100 760.200 389.400 ;
        RECT 775.200 388.200 777.000 395.400 ;
        RECT 790.800 389.400 792.600 395.400 ;
        RECT 773.400 387.300 777.000 388.200 ;
        RECT 791.400 387.300 792.600 389.400 ;
        RECT 793.800 390.300 795.600 395.400 ;
        RECT 799.800 390.300 801.600 395.400 ;
        RECT 793.800 388.950 801.600 390.300 ;
        RECT 814.200 389.400 816.000 395.400 ;
        RECT 740.100 384.150 741.900 384.900 ;
        RECT 704.100 380.100 705.900 380.850 ;
        RECT 706.950 379.950 709.050 382.050 ;
        RECT 710.100 380.100 711.900 380.850 ;
        RECT 718.950 379.950 724.050 382.050 ;
        RECT 730.950 379.950 733.050 382.050 ;
        RECT 736.950 379.950 739.050 382.050 ;
        RECT 756.150 381.900 756.900 386.100 ;
        RECT 757.950 382.950 763.050 385.050 ;
        RECT 773.400 383.100 774.600 387.300 ;
        RECT 791.400 386.250 795.150 387.300 ;
        RECT 793.950 386.100 795.150 386.250 ;
        RECT 814.950 386.100 816.000 389.400 ;
        RECT 826.950 388.950 829.050 391.050 ;
        RECT 791.100 383.100 792.900 383.850 ;
        RECT 793.950 382.950 796.050 385.050 ;
        RECT 797.100 383.100 798.900 383.850 ;
        RECT 799.950 382.950 802.050 385.050 ;
        RECT 808.950 382.950 811.050 385.050 ;
        RECT 812.250 383.100 813.900 383.850 ;
        RECT 814.950 382.950 817.050 385.050 ;
        RECT 818.100 383.100 819.750 383.850 ;
        RECT 820.950 382.950 823.050 385.050 ;
        RECT 752.100 381.150 753.900 381.900 ;
        RECT 700.950 376.950 706.050 379.050 ;
        RECT 707.400 369.600 708.600 378.900 ;
        RECT 694.950 364.950 697.050 367.050 ;
        RECT 706.800 363.600 708.600 369.600 ;
        RECT 722.400 369.600 723.600 378.900 ;
        RECT 731.550 370.050 732.450 379.950 ;
        RECT 722.400 363.600 724.200 369.600 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 737.400 369.600 738.600 378.900 ;
        RECT 756.150 378.300 757.050 381.900 ;
        RECT 756.150 377.400 758.100 378.300 ;
        RECT 736.800 363.600 738.600 369.600 ;
        RECT 752.400 376.500 758.100 377.400 ;
        RECT 752.400 369.600 753.600 376.500 ;
        RECT 759.000 375.600 760.200 381.900 ;
        RECT 770.100 380.100 771.900 380.850 ;
        RECT 772.950 379.950 775.050 382.050 ;
        RECT 776.100 380.100 777.900 380.850 ;
        RECT 790.950 379.950 793.050 382.050 ;
        RECT 752.400 363.600 754.200 369.600 ;
        RECT 758.700 363.600 760.500 375.600 ;
        RECT 773.400 369.600 774.600 378.900 ;
        RECT 775.950 376.950 778.050 379.050 ;
        RECT 794.850 378.900 795.900 381.900 ;
        RECT 796.950 379.950 799.050 382.050 ;
        RECT 800.100 381.150 801.900 381.900 ;
        RECT 809.250 381.150 810.900 381.900 ;
        RECT 811.950 379.950 814.050 382.050 ;
        RECT 816.150 378.900 816.900 381.900 ;
        RECT 817.950 379.950 820.050 382.050 ;
        RECT 821.100 381.150 822.900 381.900 ;
        RECT 794.850 375.600 796.050 378.900 ;
        RECT 816.150 377.400 817.050 378.900 ;
        RECT 816.150 376.500 820.200 377.400 ;
        RECT 773.400 363.600 775.200 369.600 ;
        RECT 794.700 363.600 796.500 375.600 ;
        RECT 809.400 374.400 817.200 375.300 ;
        RECT 809.400 363.600 811.200 374.400 ;
        RECT 815.400 364.500 817.200 374.400 ;
        RECT 818.400 365.400 820.200 376.500 ;
        RECT 821.400 364.500 823.200 375.600 ;
        RECT 827.550 370.050 828.450 388.950 ;
        RECT 838.200 388.200 840.000 395.400 ;
        RECT 853.950 391.950 856.050 394.050 ;
        RECT 844.950 388.950 847.050 391.050 ;
        RECT 836.400 387.300 840.000 388.200 ;
        RECT 836.400 383.100 837.600 387.300 ;
        RECT 833.100 380.100 834.900 380.850 ;
        RECT 835.950 379.950 838.050 382.050 ;
        RECT 839.100 380.100 840.900 380.850 ;
        RECT 845.550 379.050 846.450 388.950 ;
        RECT 832.950 376.950 835.050 379.050 ;
        RECT 826.950 367.950 829.050 370.050 ;
        RECT 836.400 369.600 837.600 378.900 ;
        RECT 838.950 376.950 841.050 379.050 ;
        RECT 844.950 376.950 847.050 379.050 ;
        RECT 854.550 370.050 855.450 391.950 ;
        RECT 815.400 363.600 823.200 364.500 ;
        RECT 836.400 363.600 838.200 369.600 ;
        RECT 853.950 367.950 856.050 370.050 ;
        RECT 10.800 353.400 12.600 359.400 ;
        RECT 11.700 353.100 12.600 353.400 ;
        RECT 16.800 353.400 18.600 359.400 ;
        RECT 16.800 353.100 18.300 353.400 ;
        RECT 11.700 352.200 18.300 353.100 ;
        RECT 11.700 347.100 12.600 352.200 ;
        RECT 17.100 347.100 18.900 347.850 ;
        RECT 35.700 347.400 37.500 359.400 ;
        RECT 55.500 347.400 57.300 359.400 ;
        RECT 73.800 353.400 75.600 359.400 ;
        RECT 74.700 353.100 75.600 353.400 ;
        RECT 79.800 353.400 81.600 359.400 ;
        RECT 79.800 353.100 81.300 353.400 ;
        RECT 74.700 352.200 81.300 353.100 ;
        RECT 10.800 343.950 13.050 346.050 ;
        RECT 16.950 343.950 19.050 346.050 ;
        RECT 35.850 344.100 37.050 347.400 ;
        RECT 55.950 344.100 57.150 347.400 ;
        RECT 74.700 347.100 75.600 352.200 ;
        RECT 80.100 347.100 81.900 347.850 ;
        RECT 98.700 347.400 100.500 359.400 ;
        RECT 116.400 353.400 118.200 359.400 ;
        RECT 116.700 353.100 118.200 353.400 ;
        RECT 122.400 353.400 124.200 359.400 ;
        RECT 122.400 353.100 123.300 353.400 ;
        RECT 116.700 352.200 123.300 353.100 ;
        RECT 73.950 345.450 76.050 346.050 ;
        RECT 11.700 337.650 12.600 342.900 ;
        RECT 13.950 340.950 16.050 343.050 ;
        RECT 19.950 340.950 22.050 343.050 ;
        RECT 31.950 340.950 34.050 343.050 ;
        RECT 35.850 341.100 36.900 344.100 ;
        RECT 37.950 340.950 40.050 343.050 ;
        RECT 41.100 341.100 42.900 341.850 ;
        RECT 50.100 341.100 51.900 341.850 ;
        RECT 52.800 340.950 55.050 343.050 ;
        RECT 56.100 341.100 57.150 344.100 ;
        RECT 68.550 344.550 76.050 345.450 ;
        RECT 58.950 340.950 61.200 343.050 ;
        RECT 14.100 339.150 15.900 339.900 ;
        RECT 20.100 339.150 21.900 339.900 ;
        RECT 32.100 339.150 33.900 339.900 ;
        RECT 34.950 337.950 37.050 340.050 ;
        RECT 38.100 339.150 39.900 339.900 ;
        RECT 40.950 337.950 43.050 340.050 ;
        RECT 49.950 337.950 52.050 340.050 ;
        RECT 53.100 339.150 54.900 339.900 ;
        RECT 55.800 337.950 58.050 340.050 ;
        RECT 59.100 339.150 60.900 339.900 ;
        RECT 11.700 336.000 15.900 337.650 ;
        RECT 34.950 336.750 36.150 336.900 ;
        RECT 14.100 327.600 15.900 336.000 ;
        RECT 32.400 335.700 36.150 336.750 ;
        RECT 56.850 336.750 58.050 336.900 ;
        RECT 56.850 335.700 60.600 336.750 ;
        RECT 32.400 333.600 33.600 335.700 ;
        RECT 31.800 327.600 33.600 333.600 ;
        RECT 34.800 332.700 42.600 334.050 ;
        RECT 34.800 327.600 36.600 332.700 ;
        RECT 40.800 327.600 42.600 332.700 ;
        RECT 50.400 332.700 58.200 334.050 ;
        RECT 50.400 327.600 52.200 332.700 ;
        RECT 56.400 327.600 58.200 332.700 ;
        RECT 59.400 333.600 60.600 335.700 ;
        RECT 59.400 327.600 61.200 333.600 ;
        RECT 68.550 331.050 69.450 344.550 ;
        RECT 73.950 343.950 76.050 344.550 ;
        RECT 79.950 343.950 82.050 346.050 ;
        RECT 98.850 344.100 100.050 347.400 ;
        RECT 116.100 347.100 117.900 347.850 ;
        RECT 122.400 347.100 123.300 352.200 ;
        RECT 139.500 347.400 141.300 359.400 ;
        RECT 157.800 353.400 159.600 359.400 ;
        RECT 158.700 353.100 159.600 353.400 ;
        RECT 163.800 353.400 165.600 359.400 ;
        RECT 178.800 353.400 180.600 359.400 ;
        RECT 163.800 353.100 165.300 353.400 ;
        RECT 158.700 352.200 165.300 353.100 ;
        RECT 179.700 353.100 180.600 353.400 ;
        RECT 184.800 353.400 186.600 359.400 ;
        RECT 200.400 353.400 202.200 359.400 ;
        RECT 184.800 353.100 186.300 353.400 ;
        RECT 179.700 352.200 186.300 353.100 ;
        RECT 74.700 337.650 75.600 342.900 ;
        RECT 76.950 340.950 79.050 343.050 ;
        RECT 82.950 340.950 85.050 343.050 ;
        RECT 94.800 340.950 97.050 343.050 ;
        RECT 98.850 341.100 99.900 344.100 ;
        RECT 115.950 343.950 118.050 346.050 ;
        RECT 121.950 343.950 124.050 346.050 ;
        RECT 139.950 344.100 141.150 347.400 ;
        RECT 158.700 347.100 159.600 352.200 ;
        RECT 164.100 347.100 165.900 347.850 ;
        RECT 179.700 347.100 180.600 352.200 ;
        RECT 185.100 347.100 186.900 347.850 ;
        RECT 100.800 340.950 103.050 343.050 ;
        RECT 104.100 341.100 105.900 341.850 ;
        RECT 112.950 340.950 115.050 343.050 ;
        RECT 118.950 340.950 121.050 343.050 ;
        RECT 77.100 339.150 78.900 339.900 ;
        RECT 83.100 339.150 84.900 339.900 ;
        RECT 95.100 339.150 96.900 339.900 ;
        RECT 97.950 337.950 100.050 340.050 ;
        RECT 101.100 339.150 102.900 339.900 ;
        RECT 103.950 337.950 106.200 340.050 ;
        RECT 113.100 339.150 114.900 339.900 ;
        RECT 119.100 339.150 120.900 339.900 ;
        RECT 122.400 337.650 123.300 342.900 ;
        RECT 134.100 341.100 135.900 341.850 ;
        RECT 136.950 340.950 139.200 343.050 ;
        RECT 140.100 341.100 141.150 344.100 ;
        RECT 154.950 343.950 160.050 346.050 ;
        RECT 163.950 343.950 166.050 346.050 ;
        RECT 178.950 345.450 181.050 346.050 ;
        RECT 173.550 344.550 181.050 345.450 ;
        RECT 142.950 340.950 145.050 343.050 ;
        RECT 133.950 337.950 136.050 340.050 ;
        RECT 137.100 339.150 138.900 339.900 ;
        RECT 139.950 337.950 142.050 340.050 ;
        RECT 143.100 339.150 144.900 339.900 ;
        RECT 74.700 336.000 78.900 337.650 ;
        RECT 97.950 336.750 99.150 336.900 ;
        RECT 67.950 328.950 70.050 331.050 ;
        RECT 77.100 327.600 78.900 336.000 ;
        RECT 95.400 335.700 99.150 336.750 ;
        RECT 119.100 336.000 123.300 337.650 ;
        RECT 158.700 337.650 159.600 342.900 ;
        RECT 160.950 340.950 163.050 343.050 ;
        RECT 166.950 340.950 169.050 343.050 ;
        RECT 161.100 339.150 162.900 339.900 ;
        RECT 167.100 339.150 168.900 339.900 ;
        RECT 140.850 336.750 142.050 336.900 ;
        RECT 95.400 333.600 96.600 335.700 ;
        RECT 94.800 327.600 96.600 333.600 ;
        RECT 97.800 332.700 105.600 334.050 ;
        RECT 97.800 327.600 99.600 332.700 ;
        RECT 103.800 327.600 105.600 332.700 ;
        RECT 119.100 327.600 120.900 336.000 ;
        RECT 140.850 335.700 144.600 336.750 ;
        RECT 158.700 336.000 162.900 337.650 ;
        RECT 173.550 337.050 174.450 344.550 ;
        RECT 178.950 343.950 181.050 344.550 ;
        RECT 184.950 343.950 187.050 346.050 ;
        RECT 196.950 343.950 199.050 346.050 ;
        RECT 200.400 344.100 201.600 353.400 ;
        RECT 221.700 347.400 223.500 359.400 ;
        RECT 240.600 347.400 242.400 359.400 ;
        RECT 247.950 349.950 250.050 352.050 ;
        RECT 202.950 343.950 205.050 346.050 ;
        RECT 221.850 344.100 223.050 347.400 ;
        RECT 239.700 346.350 242.400 347.400 ;
        RECT 179.700 337.650 180.600 342.900 ;
        RECT 181.950 340.950 184.050 343.050 ;
        RECT 187.950 340.950 190.050 343.050 ;
        RECT 197.100 342.150 198.900 342.900 ;
        RECT 199.950 340.950 202.050 343.050 ;
        RECT 203.100 342.150 204.900 342.900 ;
        RECT 217.950 340.950 220.050 343.050 ;
        RECT 221.850 341.100 222.900 344.100 ;
        RECT 223.950 340.950 226.050 343.050 ;
        RECT 227.100 341.100 228.900 341.850 ;
        RECT 236.100 341.100 237.900 341.850 ;
        RECT 239.700 341.100 241.050 346.350 ;
        RECT 242.100 341.100 243.900 341.850 ;
        RECT 182.100 339.150 183.900 339.900 ;
        RECT 188.100 339.150 189.900 339.900 ;
        RECT 134.400 332.700 142.200 334.050 ;
        RECT 134.400 327.600 136.200 332.700 ;
        RECT 140.400 327.600 142.200 332.700 ;
        RECT 143.400 333.600 144.600 335.700 ;
        RECT 143.400 327.600 145.200 333.600 ;
        RECT 161.100 327.600 162.900 336.000 ;
        RECT 172.950 334.950 175.050 337.050 ;
        RECT 179.700 336.000 183.900 337.650 ;
        RECT 182.100 327.600 183.900 336.000 ;
        RECT 200.400 335.700 201.600 339.900 ;
        RECT 218.100 339.150 219.900 339.900 ;
        RECT 220.950 337.950 223.050 340.050 ;
        RECT 224.100 339.150 225.900 339.900 ;
        RECT 226.950 337.950 229.050 340.050 ;
        RECT 235.950 337.950 238.050 340.050 ;
        RECT 239.700 338.100 240.900 341.100 ;
        RECT 248.550 340.050 249.450 349.950 ;
        RECT 260.700 347.400 262.500 359.400 ;
        RECT 271.950 355.950 274.050 358.050 ;
        RECT 260.850 344.100 262.050 347.400 ;
        RECT 256.950 340.950 259.050 343.050 ;
        RECT 260.850 341.100 261.900 344.100 ;
        RECT 262.950 340.950 265.050 343.050 ;
        RECT 266.100 341.100 267.900 341.850 ;
        RECT 241.950 337.950 244.050 340.050 ;
        RECT 247.950 337.950 250.050 340.050 ;
        RECT 257.100 339.150 258.900 339.900 ;
        RECT 259.950 337.950 262.050 340.050 ;
        RECT 263.100 339.150 264.900 339.900 ;
        RECT 265.950 337.950 268.050 340.050 ;
        RECT 272.550 337.050 273.450 355.950 ;
        RECT 281.700 347.400 283.500 359.400 ;
        RECT 301.500 347.400 303.300 359.400 ;
        RECT 322.800 353.400 324.600 359.400 ;
        RECT 281.850 344.100 283.050 347.400 ;
        RECT 301.950 344.100 303.150 347.400 ;
        RECT 277.950 340.950 280.050 343.050 ;
        RECT 281.850 341.100 282.900 344.100 ;
        RECT 283.950 340.950 286.050 343.050 ;
        RECT 287.100 341.100 288.900 341.850 ;
        RECT 296.100 341.100 297.900 341.850 ;
        RECT 298.950 340.950 301.050 343.050 ;
        RECT 302.100 341.100 303.150 344.100 ;
        RECT 319.950 343.950 322.050 346.050 ;
        RECT 323.400 344.100 324.600 353.400 ;
        RECT 337.200 347.400 339.000 359.400 ;
        RECT 343.800 353.400 345.600 359.400 ;
        RECT 361.800 353.400 363.600 359.400 ;
        RECT 325.950 343.950 328.050 346.050 ;
        RECT 304.950 340.950 307.050 343.050 ;
        RECT 320.100 342.150 321.900 342.900 ;
        RECT 322.950 340.950 325.050 343.050 ;
        RECT 326.100 342.150 327.900 342.900 ;
        RECT 337.950 341.100 339.000 347.400 ;
        RECT 340.950 340.950 343.050 343.050 ;
        RECT 278.100 339.150 279.900 339.900 ;
        RECT 280.950 337.950 283.200 340.050 ;
        RECT 284.100 339.150 285.900 339.900 ;
        RECT 286.950 337.950 289.200 340.050 ;
        RECT 295.950 337.950 298.050 340.050 ;
        RECT 299.100 339.150 300.900 339.900 ;
        RECT 301.950 337.950 304.050 340.050 ;
        RECT 305.100 339.150 306.900 339.900 ;
        RECT 220.950 336.750 222.150 336.900 ;
        RECT 218.400 335.700 222.150 336.750 ;
        RECT 200.400 334.800 204.000 335.700 ;
        RECT 202.200 327.600 204.000 334.800 ;
        RECT 218.400 333.600 219.600 335.700 ;
        RECT 238.950 334.950 241.050 337.050 ;
        RECT 259.950 336.750 261.150 336.900 ;
        RECT 257.400 335.700 261.150 336.750 ;
        RECT 217.800 327.600 219.600 333.600 ;
        RECT 220.800 332.700 228.600 334.050 ;
        RECT 220.800 327.600 222.600 332.700 ;
        RECT 226.800 327.600 228.600 332.700 ;
        RECT 239.400 330.600 240.600 333.900 ;
        RECT 257.400 333.600 258.600 335.700 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 280.950 336.750 282.150 336.900 ;
        RECT 278.400 335.700 282.150 336.750 ;
        RECT 302.850 336.750 304.050 336.900 ;
        RECT 302.850 335.700 306.600 336.750 ;
        RECT 323.400 335.700 324.600 339.900 ;
        RECT 337.950 339.450 340.050 340.050 ;
        RECT 239.400 327.600 241.200 330.600 ;
        RECT 256.800 327.600 258.600 333.600 ;
        RECT 259.800 332.700 267.600 334.050 ;
        RECT 278.400 333.600 279.600 335.700 ;
        RECT 259.800 327.600 261.600 332.700 ;
        RECT 265.800 327.600 267.600 332.700 ;
        RECT 277.800 327.600 279.600 333.600 ;
        RECT 280.800 332.700 288.600 334.050 ;
        RECT 280.800 327.600 282.600 332.700 ;
        RECT 286.800 327.600 288.600 332.700 ;
        RECT 296.400 332.700 304.200 334.050 ;
        RECT 296.400 327.600 298.200 332.700 ;
        RECT 302.400 327.600 304.200 332.700 ;
        RECT 305.400 333.600 306.600 335.700 ;
        RECT 321.000 334.800 324.600 335.700 ;
        RECT 332.550 338.550 340.050 339.450 ;
        RECT 341.100 339.150 342.900 339.900 ;
        RECT 305.400 327.600 307.200 333.600 ;
        RECT 321.000 327.600 322.800 334.800 ;
        RECT 332.550 331.050 333.450 338.550 ;
        RECT 337.950 337.950 340.050 338.550 ;
        RECT 339.150 333.600 340.050 336.900 ;
        RECT 344.550 336.300 345.600 353.400 ;
        RECT 358.950 343.950 361.050 349.050 ;
        RECT 362.400 344.100 363.600 353.400 ;
        RECT 377.400 347.400 379.200 359.400 ;
        RECT 382.950 352.950 385.050 355.050 ;
        RECT 392.400 353.400 394.200 359.400 ;
        RECT 400.950 355.950 403.050 358.050 ;
        RECT 364.950 343.950 367.050 346.050 ;
        RECT 359.100 342.150 360.900 342.900 ;
        RECT 347.100 341.100 348.900 341.850 ;
        RECT 361.950 340.950 364.050 343.050 ;
        RECT 365.100 342.150 366.900 342.900 ;
        RECT 373.950 340.950 376.050 343.050 ;
        RECT 377.400 341.100 378.600 347.400 ;
        RECT 346.950 337.950 349.200 340.050 ;
        RECT 341.100 335.100 348.600 336.300 ;
        RECT 362.400 335.700 363.600 339.900 ;
        RECT 374.100 339.150 375.900 339.900 ;
        RECT 376.950 337.950 379.050 340.050 ;
        RECT 341.100 334.500 342.900 335.100 ;
        RECT 339.150 331.800 341.100 333.600 ;
        RECT 331.950 328.950 334.050 331.050 ;
        RECT 339.300 327.600 341.100 331.800 ;
        RECT 346.800 327.600 348.600 335.100 ;
        RECT 360.000 334.800 363.600 335.700 ;
        RECT 360.000 327.600 361.800 334.800 ;
        RECT 377.400 333.600 378.600 336.900 ;
        RECT 383.550 334.050 384.450 352.950 ;
        RECT 388.950 343.950 391.050 346.050 ;
        RECT 392.400 344.100 393.600 353.400 ;
        RECT 401.550 346.050 402.450 355.950 ;
        RECT 407.400 353.400 409.200 359.400 ;
        RECT 407.400 346.500 408.600 353.400 ;
        RECT 413.700 347.400 415.500 359.400 ;
        RECT 427.800 353.400 429.600 359.400 ;
        RECT 394.950 345.450 397.050 346.050 ;
        RECT 399.000 345.450 403.050 346.050 ;
        RECT 407.400 345.600 413.100 346.500 ;
        RECT 394.950 344.550 403.050 345.450 ;
        RECT 394.950 343.950 397.050 344.550 ;
        RECT 399.000 343.950 403.050 344.550 ;
        RECT 411.150 344.700 413.100 345.600 ;
        RECT 389.100 342.150 390.900 342.900 ;
        RECT 391.950 340.950 394.050 343.050 ;
        RECT 395.100 342.150 396.900 342.900 ;
        RECT 407.100 341.100 408.900 341.850 ;
        RECT 411.150 341.100 412.050 344.700 ;
        RECT 414.000 341.100 415.200 347.400 ;
        RECT 428.400 344.100 429.600 353.400 ;
        RECT 436.950 349.950 439.050 352.050 ;
        RECT 392.400 335.700 393.600 339.900 ;
        RECT 406.950 337.950 409.050 340.050 ;
        RECT 411.150 336.900 411.900 341.100 ;
        RECT 424.950 340.950 430.050 343.050 ;
        RECT 437.550 340.050 438.450 349.950 ;
        RECT 444.600 347.400 446.400 359.400 ;
        RECT 460.800 358.500 468.600 359.400 ;
        RECT 460.800 347.400 462.600 358.500 ;
        RECT 444.600 346.350 447.300 347.400 ;
        RECT 443.100 341.100 444.900 341.850 ;
        RECT 445.950 341.100 447.300 346.350 ;
        RECT 463.800 346.500 465.600 357.600 ;
        RECT 466.800 348.600 468.600 358.500 ;
        RECT 472.800 348.600 474.600 359.400 ;
        RECT 466.800 347.700 474.600 348.600 ;
        RECT 486.600 347.400 488.400 359.400 ;
        RECT 496.950 355.950 499.050 358.050 ;
        RECT 497.550 352.050 498.450 355.950 ;
        RECT 496.950 349.950 499.050 352.050 ;
        RECT 463.800 345.600 467.850 346.500 ;
        RECT 486.600 346.350 489.300 347.400 ;
        RECT 466.950 344.100 467.850 345.600 ;
        RECT 449.100 341.100 450.900 341.850 ;
        RECT 461.100 341.100 462.900 341.850 ;
        RECT 412.950 337.950 418.050 340.050 ;
        RECT 411.150 336.300 412.050 336.900 ;
        RECT 392.400 334.800 396.000 335.700 ;
        RECT 411.150 335.400 413.100 336.300 ;
        RECT 377.400 327.600 379.200 333.600 ;
        RECT 382.950 331.950 385.050 334.050 ;
        RECT 394.200 327.600 396.000 334.800 ;
        RECT 408.000 334.500 413.100 335.400 ;
        RECT 408.000 330.600 409.200 334.500 ;
        RECT 414.000 333.600 415.200 336.900 ;
        RECT 407.400 327.600 409.200 330.600 ;
        RECT 413.700 327.600 415.500 333.600 ;
        RECT 428.400 330.600 429.600 339.900 ;
        RECT 431.100 338.100 432.900 338.850 ;
        RECT 436.950 337.950 439.050 340.050 ;
        RECT 442.950 337.950 445.050 340.050 ;
        RECT 446.100 338.100 447.300 341.100 ;
        RECT 463.950 340.950 466.050 343.050 ;
        RECT 467.100 341.100 467.850 344.100 ;
        RECT 469.950 340.950 472.050 343.050 ;
        RECT 473.100 341.100 474.750 341.850 ;
        RECT 485.100 341.100 486.900 341.850 ;
        RECT 487.950 341.100 489.300 346.350 ;
        RECT 491.100 341.100 492.900 341.850 ;
        RECT 448.950 337.950 451.050 340.050 ;
        RECT 460.800 337.950 463.050 340.050 ;
        RECT 464.250 339.150 465.900 339.900 ;
        RECT 466.950 337.950 469.050 340.050 ;
        RECT 470.100 339.150 471.750 339.900 ;
        RECT 472.950 337.950 475.050 340.050 ;
        RECT 484.950 339.450 487.050 340.050 ;
        RECT 479.550 338.550 487.050 339.450 ;
        RECT 430.950 331.950 433.050 337.050 ;
        RECT 445.950 334.950 448.050 337.050 ;
        RECT 446.400 330.600 447.600 333.900 ;
        RECT 427.800 327.600 429.600 330.600 ;
        RECT 445.800 327.600 447.600 330.600 ;
        RECT 468.000 333.600 469.050 336.900 ;
        RECT 468.000 327.600 469.800 333.600 ;
        RECT 479.550 331.050 480.450 338.550 ;
        RECT 484.950 337.950 487.050 338.550 ;
        RECT 488.100 338.100 489.300 341.100 ;
        RECT 490.950 337.950 493.050 340.050 ;
        RECT 497.550 339.450 498.450 349.950 ;
        RECT 504.600 347.400 506.400 359.400 ;
        RECT 514.950 349.950 517.050 352.050 ;
        RECT 504.600 346.350 507.300 347.400 ;
        RECT 503.100 341.100 504.900 341.850 ;
        RECT 505.950 341.100 507.300 346.350 ;
        RECT 509.100 341.100 510.900 341.850 ;
        RECT 502.950 339.450 505.050 340.050 ;
        RECT 497.550 338.550 505.050 339.450 ;
        RECT 502.950 337.950 505.050 338.550 ;
        RECT 506.100 338.100 507.300 341.100 ;
        RECT 508.950 337.950 511.200 340.050 ;
        RECT 515.550 339.450 516.450 349.950 ;
        RECT 520.800 347.400 522.600 359.400 ;
        RECT 523.800 348.300 525.600 359.400 ;
        RECT 529.800 348.300 531.600 359.400 ;
        RECT 541.800 353.400 543.600 359.400 ;
        RECT 523.800 347.400 531.600 348.300 ;
        RECT 521.400 341.100 522.300 347.400 ;
        RECT 542.400 344.100 543.600 353.400 ;
        RECT 547.950 346.950 550.050 349.050 ;
        RECT 559.500 347.400 561.300 359.400 ;
        RECT 571.950 355.950 574.050 358.050 ;
        RECT 523.950 340.950 526.050 343.050 ;
        RECT 527.100 341.100 528.900 341.850 ;
        RECT 529.950 340.950 532.050 343.050 ;
        RECT 541.950 342.450 544.050 343.050 ;
        RECT 548.550 342.450 549.450 346.950 ;
        RECT 559.950 344.100 561.150 347.400 ;
        RECT 541.950 341.550 549.450 342.450 ;
        RECT 541.950 340.950 544.050 341.550 ;
        RECT 554.100 341.100 555.900 341.850 ;
        RECT 556.800 340.950 559.050 343.050 ;
        RECT 560.100 341.100 561.150 344.100 ;
        RECT 562.950 340.950 565.050 343.050 ;
        RECT 572.550 340.050 573.450 355.950 ;
        RECT 580.800 353.400 582.600 359.400 ;
        RECT 577.950 343.950 580.050 346.050 ;
        RECT 581.400 344.100 582.600 353.400 ;
        RECT 598.500 347.400 600.300 359.400 ;
        RECT 607.950 355.950 610.050 358.050 ;
        RECT 583.950 343.950 586.050 346.050 ;
        RECT 598.950 344.100 600.150 347.400 ;
        RECT 578.100 342.150 579.900 342.900 ;
        RECT 580.950 340.950 583.200 343.050 ;
        RECT 584.100 342.150 585.900 342.900 ;
        RECT 593.100 341.100 594.900 341.850 ;
        RECT 595.950 340.950 598.050 343.050 ;
        RECT 599.100 341.100 600.150 344.100 ;
        RECT 601.950 340.950 604.050 343.050 ;
        RECT 520.950 339.450 523.050 340.050 ;
        RECT 515.550 338.550 523.050 339.450 ;
        RECT 524.100 339.150 525.900 339.900 ;
        RECT 487.950 334.950 490.050 337.050 ;
        RECT 505.950 334.950 508.050 337.050 ;
        RECT 515.550 334.050 516.450 338.550 ;
        RECT 520.950 337.950 523.050 338.550 ;
        RECT 526.950 337.950 529.200 340.050 ;
        RECT 530.100 339.150 531.900 339.900 ;
        RECT 478.950 328.950 481.050 331.050 ;
        RECT 488.400 330.600 489.600 333.900 ;
        RECT 506.400 330.600 507.600 333.900 ;
        RECT 514.950 331.950 517.050 334.050 ;
        RECT 521.400 333.600 522.300 336.900 ;
        RECT 521.400 331.950 526.800 333.600 ;
        RECT 487.800 327.600 489.600 330.600 ;
        RECT 505.800 327.600 507.600 330.600 ;
        RECT 525.000 327.600 526.800 331.950 ;
        RECT 542.400 330.600 543.600 339.900 ;
        RECT 545.100 338.100 546.900 338.850 ;
        RECT 553.950 337.950 556.050 340.050 ;
        RECT 557.100 339.150 558.900 339.900 ;
        RECT 559.950 337.950 562.050 340.050 ;
        RECT 563.100 339.150 564.900 339.900 ;
        RECT 571.950 337.950 574.050 340.050 ;
        RECT 544.950 334.950 547.050 337.050 ;
        RECT 560.850 336.750 562.050 336.900 ;
        RECT 560.850 335.700 564.600 336.750 ;
        RECT 581.400 335.700 582.600 339.900 ;
        RECT 592.950 337.950 595.050 340.050 ;
        RECT 596.100 339.150 597.900 339.900 ;
        RECT 598.950 337.950 601.050 340.050 ;
        RECT 602.100 339.150 603.900 339.900 ;
        RECT 599.850 336.750 601.050 336.900 ;
        RECT 599.850 335.700 603.600 336.750 ;
        RECT 541.800 327.600 543.600 330.600 ;
        RECT 554.400 332.700 562.200 334.050 ;
        RECT 554.400 327.600 556.200 332.700 ;
        RECT 560.400 327.600 562.200 332.700 ;
        RECT 563.400 333.600 564.600 335.700 ;
        RECT 579.000 334.800 582.600 335.700 ;
        RECT 563.400 327.600 565.200 333.600 ;
        RECT 579.000 327.600 580.800 334.800 ;
        RECT 593.400 332.700 601.200 334.050 ;
        RECT 593.400 327.600 595.200 332.700 ;
        RECT 599.400 327.600 601.200 332.700 ;
        RECT 602.400 333.600 603.600 335.700 ;
        RECT 602.400 327.600 604.200 333.600 ;
        RECT 608.550 331.050 609.450 355.950 ;
        RECT 620.700 347.400 622.500 359.400 ;
        RECT 639.600 347.400 641.400 359.400 ;
        RECT 658.800 353.400 660.600 359.400 ;
        RECT 620.850 344.100 622.050 347.400 ;
        RECT 638.700 346.350 641.400 347.400 ;
        RECT 616.950 340.950 619.050 343.050 ;
        RECT 620.850 341.100 621.900 344.100 ;
        RECT 622.950 340.950 625.050 343.050 ;
        RECT 626.100 341.100 627.900 341.850 ;
        RECT 635.100 341.100 636.900 341.850 ;
        RECT 638.700 341.100 640.050 346.350 ;
        RECT 655.950 343.950 658.050 346.050 ;
        RECT 659.400 344.100 660.600 353.400 ;
        RECT 673.800 358.500 681.600 359.400 ;
        RECT 673.800 347.400 675.600 358.500 ;
        RECT 676.800 346.500 678.600 357.600 ;
        RECT 679.800 348.600 681.600 358.500 ;
        RECT 685.800 348.600 687.600 359.400 ;
        RECT 691.950 355.950 694.050 358.050 ;
        RECT 692.550 349.050 693.450 355.950 ;
        RECT 679.800 347.700 687.600 348.600 ;
        RECT 691.950 346.950 694.050 349.050 ;
        RECT 695.400 348.600 697.200 359.400 ;
        RECT 701.400 358.500 709.200 359.400 ;
        RECT 701.400 348.600 703.200 358.500 ;
        RECT 695.400 347.700 703.200 348.600 ;
        RECT 704.400 346.500 706.200 357.600 ;
        RECT 707.400 347.400 709.200 358.500 ;
        RECT 724.800 353.400 726.600 359.400 ;
        RECT 712.950 346.950 715.050 349.050 ;
        RECT 661.950 343.950 664.050 346.050 ;
        RECT 676.800 345.600 680.850 346.500 ;
        RECT 679.950 344.100 680.850 345.600 ;
        RECT 656.100 342.150 657.900 342.900 ;
        RECT 641.100 341.100 642.900 341.850 ;
        RECT 610.950 337.950 613.050 340.050 ;
        RECT 617.100 339.150 618.900 339.900 ;
        RECT 619.950 337.950 622.050 340.050 ;
        RECT 623.100 339.150 624.900 339.900 ;
        RECT 625.950 337.950 628.050 340.050 ;
        RECT 634.800 337.950 637.050 340.050 ;
        RECT 638.700 338.100 639.900 341.100 ;
        RECT 658.950 340.950 661.050 343.050 ;
        RECT 662.100 342.150 663.900 342.900 ;
        RECT 674.100 341.100 675.900 341.850 ;
        RECT 676.950 340.950 679.050 343.050 ;
        RECT 680.100 341.100 680.850 344.100 ;
        RECT 702.150 345.600 706.200 346.500 ;
        RECT 702.150 344.100 703.050 345.600 ;
        RECT 682.950 340.950 685.050 343.050 ;
        RECT 686.100 341.100 687.750 341.850 ;
        RECT 695.250 341.100 696.900 341.850 ;
        RECT 697.950 340.950 700.050 343.050 ;
        RECT 702.150 341.100 702.900 344.100 ;
        RECT 703.950 340.950 706.200 343.050 ;
        RECT 707.100 341.100 708.900 341.850 ;
        RECT 713.550 340.050 714.450 346.950 ;
        RECT 721.950 343.950 724.050 346.050 ;
        RECT 725.400 344.100 726.600 353.400 ;
        RECT 739.200 347.400 741.000 359.400 ;
        RECT 745.800 353.400 747.600 359.400 ;
        RECT 727.950 343.950 730.050 346.050 ;
        RECT 715.950 340.950 718.050 343.050 ;
        RECT 722.100 342.150 723.900 342.900 ;
        RECT 724.950 340.950 727.200 343.050 ;
        RECT 728.100 342.150 729.900 342.900 ;
        RECT 739.950 341.100 741.000 347.400 ;
        RECT 742.950 340.950 745.050 343.050 ;
        RECT 640.950 337.950 643.200 340.050 ;
        RECT 611.550 331.050 612.450 337.950 ;
        RECT 619.950 336.750 621.150 336.900 ;
        RECT 617.400 335.700 621.150 336.750 ;
        RECT 617.400 333.600 618.600 335.700 ;
        RECT 637.800 334.950 640.050 337.050 ;
        RECT 659.400 335.700 660.600 339.900 ;
        RECT 673.800 337.950 676.050 340.050 ;
        RECT 677.250 339.150 678.900 339.900 ;
        RECT 679.950 337.950 682.050 340.050 ;
        RECT 683.100 339.150 684.750 339.900 ;
        RECT 685.950 337.950 688.050 340.050 ;
        RECT 694.950 337.950 697.050 340.050 ;
        RECT 698.250 339.150 699.900 339.900 ;
        RECT 700.950 337.950 703.050 340.050 ;
        RECT 704.100 339.150 705.750 339.900 ;
        RECT 706.950 337.950 709.050 340.050 ;
        RECT 712.950 337.950 715.050 340.050 ;
        RECT 657.000 334.800 660.600 335.700 ;
        RECT 607.800 328.950 609.900 331.050 ;
        RECT 611.100 328.950 613.200 331.050 ;
        RECT 616.800 327.600 618.600 333.600 ;
        RECT 619.800 332.700 627.600 334.050 ;
        RECT 619.800 327.600 621.600 332.700 ;
        RECT 625.800 327.600 627.600 332.700 ;
        RECT 638.400 330.600 639.600 333.900 ;
        RECT 638.400 327.600 640.200 330.600 ;
        RECT 657.000 327.600 658.800 334.800 ;
        RECT 681.000 333.600 682.050 336.900 ;
        RECT 700.950 333.600 702.000 336.900 ;
        RECT 681.000 327.600 682.800 333.600 ;
        RECT 700.200 327.600 702.000 333.600 ;
        RECT 716.550 331.050 717.450 340.950 ;
        RECT 725.400 335.700 726.600 339.900 ;
        RECT 736.950 337.950 742.050 340.050 ;
        RECT 743.100 339.150 744.900 339.900 ;
        RECT 723.000 334.800 726.600 335.700 ;
        RECT 715.950 328.950 718.050 331.050 ;
        RECT 723.000 327.600 724.800 334.800 ;
        RECT 741.150 333.600 742.050 336.900 ;
        RECT 746.550 336.300 747.600 353.400 ;
        RECT 758.400 348.600 760.200 359.400 ;
        RECT 764.400 358.500 772.200 359.400 ;
        RECT 764.400 348.600 766.200 358.500 ;
        RECT 758.400 347.700 766.200 348.600 ;
        RECT 767.400 346.500 769.200 357.600 ;
        RECT 770.400 347.400 772.200 358.500 ;
        RECT 775.950 346.950 778.050 349.050 ;
        RECT 782.400 348.600 784.200 359.400 ;
        RECT 788.400 358.500 796.200 359.400 ;
        RECT 788.400 348.600 790.200 358.500 ;
        RECT 782.400 347.700 790.200 348.600 ;
        RECT 765.150 345.600 769.200 346.500 ;
        RECT 765.150 344.100 766.050 345.600 ;
        RECT 749.100 341.100 750.900 341.850 ;
        RECT 758.250 341.100 759.900 341.850 ;
        RECT 760.950 340.950 763.050 343.050 ;
        RECT 765.150 341.100 765.900 344.100 ;
        RECT 766.950 340.950 769.050 343.050 ;
        RECT 770.100 341.100 771.900 341.850 ;
        RECT 776.550 340.050 777.450 346.950 ;
        RECT 791.400 346.500 793.200 357.600 ;
        RECT 794.400 347.400 796.200 358.500 ;
        RECT 802.950 349.950 805.050 352.050 ;
        RECT 789.150 345.600 793.200 346.500 ;
        RECT 789.150 344.100 790.050 345.600 ;
        RECT 782.250 341.100 783.900 341.850 ;
        RECT 784.950 340.950 787.050 343.050 ;
        RECT 789.150 341.100 789.900 344.100 ;
        RECT 790.800 340.950 793.050 343.050 ;
        RECT 794.100 341.100 795.900 341.850 ;
        RECT 748.950 337.950 751.050 340.050 ;
        RECT 757.800 337.950 760.050 340.050 ;
        RECT 761.250 339.150 762.900 339.900 ;
        RECT 763.950 337.950 766.050 340.050 ;
        RECT 767.100 339.150 768.750 339.900 ;
        RECT 769.950 337.950 772.050 340.050 ;
        RECT 775.950 337.950 778.050 340.050 ;
        RECT 781.950 337.950 784.050 340.050 ;
        RECT 785.250 339.150 786.900 339.900 ;
        RECT 787.950 337.950 790.050 340.050 ;
        RECT 791.100 339.150 792.750 339.900 ;
        RECT 793.950 337.950 796.050 340.050 ;
        RECT 743.100 335.100 750.600 336.300 ;
        RECT 743.100 334.500 744.900 335.100 ;
        RECT 741.150 331.800 743.100 333.600 ;
        RECT 741.300 327.600 743.100 331.800 ;
        RECT 748.800 327.600 750.600 335.100 ;
        RECT 763.950 333.600 765.000 336.900 ;
        RECT 787.950 333.600 789.000 336.900 ;
        RECT 763.200 327.600 765.000 333.600 ;
        RECT 787.200 327.600 789.000 333.600 ;
        RECT 803.550 331.050 804.450 349.950 ;
        RECT 812.700 347.400 814.500 359.400 ;
        RECT 832.500 347.400 834.300 359.400 ;
        RECT 844.950 355.950 847.050 358.050 ;
        RECT 845.550 349.050 846.450 355.950 ;
        RECT 812.850 344.100 814.050 347.400 ;
        RECT 832.950 344.100 834.150 347.400 ;
        RECT 844.950 346.950 847.050 349.050 ;
        RECT 808.950 340.950 811.050 343.050 ;
        RECT 812.850 341.100 813.900 344.100 ;
        RECT 814.950 340.950 817.050 343.050 ;
        RECT 818.100 341.100 819.900 341.850 ;
        RECT 827.100 341.100 828.900 341.850 ;
        RECT 829.950 340.950 832.050 343.050 ;
        RECT 833.100 341.100 834.150 344.100 ;
        RECT 835.950 342.450 838.050 343.050 ;
        RECT 835.950 341.550 843.450 342.450 ;
        RECT 835.950 340.950 838.050 341.550 ;
        RECT 809.100 339.150 810.900 339.900 ;
        RECT 811.950 337.950 814.050 340.050 ;
        RECT 815.100 339.150 816.900 339.900 ;
        RECT 817.950 337.950 820.050 340.050 ;
        RECT 826.800 337.950 829.050 340.050 ;
        RECT 830.100 339.150 831.900 339.900 ;
        RECT 832.950 337.950 835.200 340.050 ;
        RECT 836.100 339.150 837.900 339.900 ;
        RECT 811.950 336.750 813.150 336.900 ;
        RECT 809.400 335.700 813.150 336.750 ;
        RECT 833.850 336.750 835.050 336.900 ;
        RECT 833.850 335.700 837.600 336.750 ;
        RECT 809.400 333.600 810.600 335.700 ;
        RECT 802.950 328.950 805.050 331.050 ;
        RECT 808.800 327.600 810.600 333.600 ;
        RECT 811.800 332.700 819.600 334.050 ;
        RECT 811.800 327.600 813.600 332.700 ;
        RECT 817.800 327.600 819.600 332.700 ;
        RECT 827.400 332.700 835.200 334.050 ;
        RECT 827.400 327.600 829.200 332.700 ;
        RECT 833.400 327.600 835.200 332.700 ;
        RECT 836.400 333.600 837.600 335.700 ;
        RECT 836.400 327.600 838.200 333.600 ;
        RECT 842.550 331.050 843.450 341.550 ;
        RECT 841.950 328.950 844.050 331.050 ;
        RECT 15.000 319.050 16.800 323.400 ;
        RECT 11.400 317.400 16.800 319.050 ;
        RECT 11.400 314.100 12.300 317.400 ;
        RECT 35.100 315.000 36.900 323.400 ;
        RECT 57.000 319.050 58.800 323.400 ;
        RECT 67.950 319.950 70.050 322.050 ;
        RECT 53.400 317.400 58.800 319.050 ;
        RECT 35.100 313.350 39.300 315.000 ;
        RECT 53.400 314.100 54.300 317.400 ;
        RECT 10.950 310.950 13.050 313.050 ;
        RECT 14.100 311.100 15.900 311.850 ;
        RECT 16.950 310.950 19.200 313.050 ;
        RECT 20.100 311.100 21.900 311.850 ;
        RECT 29.100 311.100 30.900 311.850 ;
        RECT 35.100 311.100 36.900 311.850 ;
        RECT 11.400 303.600 12.300 309.900 ;
        RECT 13.950 307.950 16.050 310.050 ;
        RECT 17.100 309.150 18.900 309.900 ;
        RECT 19.950 307.950 22.050 310.050 ;
        RECT 28.950 307.950 31.200 310.050 ;
        RECT 34.950 307.950 37.050 310.050 ;
        RECT 38.400 308.100 39.300 313.350 ;
        RECT 49.950 310.950 55.050 313.050 ;
        RECT 56.100 311.100 57.900 311.850 ;
        RECT 58.950 310.950 61.050 313.050 ;
        RECT 62.100 311.100 63.900 311.850 ;
        RECT 31.950 304.950 34.050 307.050 ;
        RECT 37.950 304.950 43.050 307.050 ;
        RECT 10.800 291.600 12.600 303.600 ;
        RECT 13.800 302.700 21.600 303.600 ;
        RECT 32.100 303.150 33.900 303.900 ;
        RECT 13.800 291.600 15.600 302.700 ;
        RECT 19.800 291.600 21.600 302.700 ;
        RECT 38.400 298.800 39.300 303.900 ;
        RECT 53.400 303.600 54.300 309.900 ;
        RECT 55.800 307.950 58.050 310.050 ;
        RECT 59.100 309.150 60.900 309.900 ;
        RECT 61.950 307.950 64.050 310.050 ;
        RECT 32.700 297.900 39.300 298.800 ;
        RECT 32.700 297.600 34.200 297.900 ;
        RECT 32.400 291.600 34.200 297.600 ;
        RECT 38.400 297.600 39.300 297.900 ;
        RECT 38.400 291.600 40.200 297.600 ;
        RECT 52.800 291.600 54.600 303.600 ;
        RECT 55.800 302.700 63.600 303.600 ;
        RECT 55.800 291.600 57.600 302.700 ;
        RECT 61.800 291.600 63.600 302.700 ;
        RECT 68.550 295.050 69.450 319.950 ;
        RECT 73.800 317.400 75.600 323.400 ;
        RECT 74.400 315.300 75.600 317.400 ;
        RECT 76.800 318.300 78.600 323.400 ;
        RECT 82.800 318.300 84.600 323.400 ;
        RECT 96.300 319.200 98.100 323.400 ;
        RECT 76.800 316.950 84.600 318.300 ;
        RECT 96.150 317.400 98.100 319.200 ;
        RECT 74.400 314.250 78.150 315.300 ;
        RECT 76.950 314.100 78.150 314.250 ;
        RECT 96.150 314.100 97.050 317.400 ;
        RECT 98.100 315.900 99.900 316.500 ;
        RECT 103.800 315.900 105.600 323.400 ;
        RECT 118.200 316.200 120.000 323.400 ;
        RECT 136.200 316.200 138.000 323.400 ;
        RECT 98.100 314.700 105.600 315.900 ;
        RECT 116.400 315.300 120.000 316.200 ;
        RECT 134.400 315.300 138.000 316.200 ;
        RECT 153.000 316.200 154.800 323.400 ;
        RECT 153.000 315.300 156.600 316.200 ;
        RECT 74.100 311.100 75.900 311.850 ;
        RECT 76.950 310.950 79.050 313.050 ;
        RECT 80.100 311.100 81.900 311.850 ;
        RECT 82.950 310.950 85.050 313.050 ;
        RECT 94.950 312.450 97.050 313.050 ;
        RECT 89.550 311.550 97.050 312.450 ;
        RECT 73.950 307.950 76.050 310.050 ;
        RECT 77.850 306.900 78.900 309.900 ;
        RECT 79.950 307.950 82.050 310.050 ;
        RECT 83.100 309.150 84.900 309.900 ;
        RECT 77.850 303.600 79.050 306.900 ;
        RECT 67.950 292.950 70.050 295.050 ;
        RECT 77.700 291.600 79.500 303.600 ;
        RECT 89.550 295.050 90.450 311.550 ;
        RECT 94.950 310.950 97.050 311.550 ;
        RECT 98.100 311.100 99.900 311.850 ;
        RECT 94.950 303.600 96.000 309.900 ;
        RECT 97.800 307.950 100.050 310.050 ;
        RECT 88.950 292.950 91.050 295.050 ;
        RECT 94.200 291.600 96.000 303.600 ;
        RECT 101.550 297.600 102.600 314.700 ;
        RECT 103.950 310.950 106.050 313.050 ;
        RECT 116.400 311.100 117.600 315.300 ;
        RECT 134.400 311.100 135.600 315.300 ;
        RECT 155.400 311.100 156.600 315.300 ;
        RECT 173.100 315.000 174.900 323.400 ;
        RECT 194.100 315.000 195.900 323.400 ;
        RECT 211.800 320.400 213.600 323.400 ;
        RECT 170.700 313.350 174.900 315.000 ;
        RECT 191.700 313.350 195.900 315.000 ;
        RECT 104.100 309.150 105.900 309.900 ;
        RECT 113.100 308.100 114.900 308.850 ;
        RECT 115.950 307.950 118.050 310.050 ;
        RECT 119.100 308.100 120.900 308.850 ;
        RECT 124.950 307.950 127.050 310.050 ;
        RECT 131.100 308.100 132.900 308.850 ;
        RECT 133.950 307.950 136.050 310.050 ;
        RECT 137.100 308.100 138.900 308.850 ;
        RECT 152.100 308.100 153.900 308.850 ;
        RECT 154.950 307.950 157.050 310.050 ;
        RECT 158.100 308.100 159.900 308.850 ;
        RECT 170.700 308.100 171.600 313.350 ;
        RECT 173.100 311.100 174.900 311.850 ;
        RECT 179.100 311.100 180.900 311.850 ;
        RECT 172.950 307.950 175.050 310.050 ;
        RECT 178.950 307.950 181.050 310.050 ;
        RECT 191.700 308.100 192.600 313.350 ;
        RECT 194.100 311.100 195.900 311.850 ;
        RECT 200.100 311.100 201.900 311.850 ;
        RECT 212.400 311.100 213.600 320.400 ;
        RECT 234.000 317.400 235.800 323.400 ;
        RECT 214.950 313.950 217.050 316.050 ;
        RECT 234.000 314.100 235.050 317.400 ;
        RECT 252.000 316.200 253.800 323.400 ;
        RECT 276.000 317.400 277.800 323.400 ;
        RECT 252.000 315.300 255.600 316.200 ;
        RECT 215.100 312.150 216.900 312.900 ;
        RECT 226.950 310.950 229.050 313.050 ;
        RECT 230.250 311.100 231.900 311.850 ;
        RECT 232.950 310.950 235.050 313.050 ;
        RECT 236.100 311.100 237.750 311.850 ;
        RECT 238.950 310.950 241.050 313.050 ;
        RECT 254.400 311.100 255.600 315.300 ;
        RECT 276.000 314.100 277.050 317.400 ;
        RECT 296.100 315.000 297.900 323.400 ;
        RECT 311.400 318.300 313.200 323.400 ;
        RECT 317.400 318.300 319.200 323.400 ;
        RECT 311.400 316.950 319.200 318.300 ;
        RECT 320.400 317.400 322.200 323.400 ;
        RECT 320.400 315.300 321.600 317.400 ;
        RECT 336.000 316.200 337.800 323.400 ;
        RECT 336.000 315.300 339.600 316.200 ;
        RECT 293.700 313.350 297.900 315.000 ;
        RECT 317.850 314.250 321.600 315.300 ;
        RECT 317.850 314.100 319.050 314.250 ;
        RECT 268.950 310.950 271.050 313.050 ;
        RECT 272.250 311.100 273.900 311.850 ;
        RECT 274.950 310.950 277.050 313.050 ;
        RECT 278.100 311.100 279.750 311.850 ;
        RECT 280.950 310.950 283.050 313.050 ;
        RECT 193.950 307.950 196.050 310.050 ;
        RECT 199.950 307.950 202.050 310.050 ;
        RECT 208.950 307.950 214.050 310.050 ;
        RECT 227.100 309.150 228.900 309.900 ;
        RECT 229.950 307.950 232.050 310.050 ;
        RECT 112.950 304.950 115.050 307.050 ;
        RECT 100.800 291.600 102.600 297.600 ;
        RECT 116.400 297.600 117.600 306.900 ;
        RECT 118.950 304.950 121.050 307.050 ;
        RECT 125.550 301.050 126.450 307.950 ;
        RECT 130.950 304.950 133.050 307.050 ;
        RECT 124.950 298.950 127.050 301.050 ;
        RECT 134.400 297.600 135.600 306.900 ;
        RECT 136.950 304.950 139.050 307.050 ;
        RECT 151.950 304.950 154.050 307.050 ;
        RECT 155.400 297.600 156.600 306.900 ;
        RECT 157.950 304.950 160.050 307.050 ;
        RECT 166.950 304.950 172.050 307.050 ;
        RECT 175.950 304.950 178.050 307.050 ;
        RECT 190.950 306.450 193.050 307.050 ;
        RECT 185.550 305.550 193.050 306.450 ;
        RECT 170.700 298.800 171.600 303.900 ;
        RECT 176.100 303.150 177.900 303.900 ;
        RECT 185.550 301.050 186.450 305.550 ;
        RECT 190.950 304.950 193.050 305.550 ;
        RECT 196.950 304.950 199.050 307.050 ;
        RECT 233.100 306.900 233.850 309.900 ;
        RECT 235.950 307.950 238.050 310.050 ;
        RECT 239.100 309.150 240.750 309.900 ;
        RECT 251.100 308.100 252.900 308.850 ;
        RECT 253.950 307.950 256.050 310.050 ;
        RECT 269.100 309.150 270.900 309.900 ;
        RECT 257.100 308.100 258.900 308.850 ;
        RECT 271.950 307.950 274.050 310.050 ;
        RECT 184.950 298.950 187.050 301.050 ;
        RECT 191.700 298.800 192.600 303.900 ;
        RECT 197.100 303.150 198.900 303.900 ;
        RECT 170.700 297.900 177.300 298.800 ;
        RECT 170.700 297.600 171.600 297.900 ;
        RECT 116.400 291.600 118.200 297.600 ;
        RECT 134.400 291.600 136.200 297.600 ;
        RECT 154.800 291.600 156.600 297.600 ;
        RECT 169.800 291.600 171.600 297.600 ;
        RECT 175.800 297.600 177.300 297.900 ;
        RECT 191.700 297.900 198.300 298.800 ;
        RECT 191.700 297.600 192.600 297.900 ;
        RECT 175.800 291.600 177.600 297.600 ;
        RECT 190.800 291.600 192.600 297.600 ;
        RECT 196.800 297.600 198.300 297.900 ;
        RECT 212.400 297.600 213.600 306.900 ;
        RECT 232.950 305.400 233.850 306.900 ;
        RECT 229.800 304.500 233.850 305.400 ;
        RECT 250.800 304.950 253.050 307.050 ;
        RECT 196.800 291.600 198.600 297.600 ;
        RECT 211.800 291.600 213.600 297.600 ;
        RECT 226.800 292.500 228.600 303.600 ;
        RECT 229.800 293.400 231.600 304.500 ;
        RECT 232.800 302.400 240.600 303.300 ;
        RECT 232.800 292.500 234.600 302.400 ;
        RECT 226.800 291.600 234.600 292.500 ;
        RECT 238.800 291.600 240.600 302.400 ;
        RECT 254.400 297.600 255.600 306.900 ;
        RECT 256.950 304.950 259.050 307.050 ;
        RECT 275.100 306.900 275.850 309.900 ;
        RECT 277.950 307.950 280.200 310.050 ;
        RECT 281.100 309.150 282.750 309.900 ;
        RECT 293.700 308.100 294.600 313.350 ;
        RECT 296.100 311.100 297.900 311.850 ;
        RECT 302.100 311.100 303.900 311.850 ;
        RECT 310.950 310.950 313.050 313.050 ;
        RECT 314.100 311.100 315.900 311.850 ;
        RECT 316.950 310.950 319.050 313.050 ;
        RECT 320.100 311.100 321.900 311.850 ;
        RECT 338.400 311.100 339.600 315.300 ;
        RECT 356.100 315.000 357.900 323.400 ;
        RECT 371.400 318.300 373.200 323.400 ;
        RECT 377.400 318.300 379.200 323.400 ;
        RECT 371.400 316.950 379.200 318.300 ;
        RECT 380.400 317.400 382.200 323.400 ;
        RECT 380.400 315.300 381.600 317.400 ;
        RECT 353.700 313.350 357.900 315.000 ;
        RECT 377.850 314.250 381.600 315.300 ;
        RECT 392.400 315.900 394.200 323.400 ;
        RECT 399.900 319.200 401.700 323.400 ;
        RECT 416.400 320.400 418.200 323.400 ;
        RECT 399.900 317.400 401.850 319.200 ;
        RECT 398.100 315.900 399.900 316.500 ;
        RECT 392.400 314.700 399.900 315.900 ;
        RECT 377.850 314.100 379.050 314.250 ;
        RECT 295.950 307.950 298.050 310.050 ;
        RECT 301.950 307.950 304.050 310.050 ;
        RECT 311.100 309.150 312.900 309.900 ;
        RECT 313.950 307.950 316.050 310.050 ;
        RECT 274.950 305.400 275.850 306.900 ;
        RECT 271.800 304.500 275.850 305.400 ;
        RECT 283.950 304.950 286.050 307.050 ;
        RECT 292.950 304.950 295.050 307.050 ;
        RECT 298.950 304.950 301.200 307.050 ;
        RECT 317.100 306.900 318.150 309.900 ;
        RECT 319.950 307.950 322.050 310.050 ;
        RECT 335.100 308.100 336.900 308.850 ;
        RECT 337.950 307.950 340.050 310.050 ;
        RECT 341.100 308.100 342.900 308.850 ;
        RECT 353.700 308.100 354.600 313.350 ;
        RECT 356.100 311.100 357.900 311.850 ;
        RECT 362.100 311.100 363.900 311.850 ;
        RECT 370.950 310.950 373.050 313.050 ;
        RECT 374.100 311.100 375.900 311.850 ;
        RECT 376.950 310.950 379.050 313.050 ;
        RECT 380.100 311.100 381.900 311.850 ;
        RECT 391.950 310.950 394.050 313.050 ;
        RECT 355.950 307.950 358.050 310.050 ;
        RECT 361.950 307.950 364.050 310.050 ;
        RECT 371.100 309.150 372.900 309.900 ;
        RECT 373.950 307.950 376.050 310.050 ;
        RECT 253.800 291.600 255.600 297.600 ;
        RECT 268.800 292.500 270.600 303.600 ;
        RECT 271.800 293.400 273.600 304.500 ;
        RECT 274.800 302.400 282.600 303.300 ;
        RECT 274.800 292.500 276.600 302.400 ;
        RECT 268.800 291.600 276.600 292.500 ;
        RECT 280.800 291.600 282.600 302.400 ;
        RECT 284.550 301.050 285.450 304.950 ;
        RECT 283.950 298.950 286.050 301.050 ;
        RECT 293.700 298.800 294.600 303.900 ;
        RECT 299.100 303.150 300.900 303.900 ;
        RECT 316.950 303.600 318.150 306.900 ;
        RECT 334.950 304.950 337.050 307.050 ;
        RECT 293.700 297.900 300.300 298.800 ;
        RECT 293.700 297.600 294.600 297.900 ;
        RECT 292.800 291.600 294.600 297.600 ;
        RECT 298.800 297.600 300.300 297.900 ;
        RECT 298.800 291.600 300.600 297.600 ;
        RECT 316.500 291.600 318.300 303.600 ;
        RECT 338.400 297.600 339.600 306.900 ;
        RECT 340.950 301.950 343.050 307.050 ;
        RECT 352.950 306.450 355.050 307.050 ;
        RECT 347.550 305.550 355.050 306.450 ;
        RECT 337.800 291.600 339.600 297.600 ;
        RECT 347.550 295.050 348.450 305.550 ;
        RECT 352.950 304.950 355.050 305.550 ;
        RECT 358.950 304.950 361.050 307.050 ;
        RECT 377.100 306.900 378.150 309.900 ;
        RECT 379.950 307.950 382.050 310.050 ;
        RECT 392.100 309.150 393.900 309.900 ;
        RECT 353.700 298.800 354.600 303.900 ;
        RECT 359.100 303.150 360.900 303.900 ;
        RECT 376.950 303.600 378.150 306.900 ;
        RECT 353.700 297.900 360.300 298.800 ;
        RECT 353.700 297.600 354.600 297.900 ;
        RECT 346.950 292.950 349.050 295.050 ;
        RECT 352.800 291.600 354.600 297.600 ;
        RECT 358.800 297.600 360.300 297.900 ;
        RECT 358.800 291.600 360.600 297.600 ;
        RECT 376.500 291.600 378.300 303.600 ;
        RECT 395.400 297.600 396.450 314.700 ;
        RECT 400.950 314.100 401.850 317.400 ;
        RECT 412.950 313.950 415.050 316.050 ;
        RECT 398.100 311.100 399.900 311.850 ;
        RECT 400.950 310.950 403.050 313.050 ;
        RECT 413.100 312.150 414.900 312.900 ;
        RECT 416.400 311.100 417.600 320.400 ;
        RECT 433.200 316.200 435.000 323.400 ;
        RECT 439.950 316.950 442.050 319.050 ;
        RECT 431.400 315.300 435.000 316.200 ;
        RECT 431.400 311.100 432.600 315.300 ;
        RECT 397.950 307.950 400.050 310.050 ;
        RECT 402.000 303.600 403.050 309.900 ;
        RECT 415.950 309.450 418.050 310.050 ;
        RECT 410.550 309.000 418.050 309.450 ;
        RECT 409.950 308.550 418.050 309.000 ;
        RECT 409.950 304.950 412.050 308.550 ;
        RECT 415.950 307.950 418.050 308.550 ;
        RECT 428.100 308.100 429.900 308.850 ;
        RECT 430.950 307.950 433.050 310.050 ;
        RECT 434.100 308.100 435.900 308.850 ;
        RECT 395.400 291.600 397.200 297.600 ;
        RECT 402.000 291.600 403.800 303.600 ;
        RECT 416.400 297.600 417.600 306.900 ;
        RECT 427.950 304.950 430.050 307.050 ;
        RECT 428.550 303.000 429.450 304.950 ;
        RECT 427.950 298.950 430.050 303.000 ;
        RECT 431.400 297.600 432.600 306.900 ;
        RECT 433.950 306.450 436.050 307.050 ;
        RECT 440.550 306.450 441.450 316.950 ;
        RECT 451.200 316.200 453.000 323.400 ;
        RECT 464.400 318.300 466.200 323.400 ;
        RECT 470.400 318.300 472.200 323.400 ;
        RECT 464.400 316.950 472.200 318.300 ;
        RECT 473.400 317.400 475.200 323.400 ;
        RECT 449.400 315.300 453.000 316.200 ;
        RECT 473.400 315.300 474.600 317.400 ;
        RECT 490.200 316.200 492.000 323.400 ;
        RECT 496.950 319.950 499.050 322.050 ;
        RECT 449.400 311.100 450.600 315.300 ;
        RECT 470.850 314.250 474.600 315.300 ;
        RECT 488.400 315.300 492.000 316.200 ;
        RECT 470.850 314.100 472.050 314.250 ;
        RECT 463.950 310.950 466.050 313.050 ;
        RECT 467.100 311.100 468.900 311.850 ;
        RECT 469.950 310.950 472.200 313.050 ;
        RECT 473.100 311.100 474.900 311.850 ;
        RECT 488.400 311.100 489.600 315.300 ;
        RECT 446.100 308.100 447.900 308.850 ;
        RECT 448.950 307.950 451.050 310.050 ;
        RECT 464.100 309.150 465.900 309.900 ;
        RECT 452.100 308.100 453.900 308.850 ;
        RECT 466.950 307.950 469.050 310.050 ;
        RECT 433.950 305.550 441.450 306.450 ;
        RECT 433.950 304.950 436.050 305.550 ;
        RECT 416.400 291.600 418.200 297.600 ;
        RECT 431.400 291.600 433.200 297.600 ;
        RECT 440.550 295.050 441.450 305.550 ;
        RECT 445.950 304.950 448.050 307.050 ;
        RECT 449.400 297.600 450.600 306.900 ;
        RECT 451.950 301.950 454.050 307.050 ;
        RECT 470.100 306.900 471.150 309.900 ;
        RECT 472.950 307.950 475.050 310.050 ;
        RECT 485.100 308.100 486.900 308.850 ;
        RECT 487.800 307.950 490.050 310.050 ;
        RECT 491.100 308.100 492.900 308.850 ;
        RECT 469.950 303.600 471.150 306.900 ;
        RECT 439.950 292.950 442.050 295.050 ;
        RECT 449.400 291.600 451.200 297.600 ;
        RECT 469.500 291.600 471.300 303.600 ;
        RECT 484.950 301.950 487.050 307.050 ;
        RECT 488.400 297.600 489.600 306.900 ;
        RECT 490.950 304.950 493.050 307.050 ;
        RECT 488.400 291.600 490.200 297.600 ;
        RECT 497.550 295.050 498.450 319.950 ;
        RECT 508.200 319.050 510.000 323.400 ;
        RECT 508.200 317.400 513.600 319.050 ;
        RECT 512.700 314.100 513.600 317.400 ;
        RECT 524.400 318.300 526.200 323.400 ;
        RECT 530.400 318.300 532.200 323.400 ;
        RECT 524.400 316.950 532.200 318.300 ;
        RECT 533.400 317.400 535.200 323.400 ;
        RECT 538.950 319.950 541.050 322.050 ;
        RECT 548.400 320.400 550.200 323.400 ;
        RECT 533.400 315.300 534.600 317.400 ;
        RECT 530.850 314.250 534.600 315.300 ;
        RECT 530.850 314.100 532.050 314.250 ;
        RECT 503.100 311.100 504.900 311.850 ;
        RECT 505.950 310.950 508.050 313.050 ;
        RECT 511.950 312.450 514.050 313.050 ;
        RECT 509.100 311.100 510.900 311.850 ;
        RECT 511.950 311.550 519.450 312.450 ;
        RECT 511.950 310.950 514.050 311.550 ;
        RECT 502.950 307.950 505.050 310.050 ;
        RECT 506.100 309.150 507.900 309.900 ;
        RECT 508.950 307.950 511.050 310.050 ;
        RECT 512.700 303.600 513.600 309.900 ;
        RECT 503.400 302.700 511.200 303.600 ;
        RECT 496.950 292.950 499.050 295.050 ;
        RECT 503.400 291.600 505.200 302.700 ;
        RECT 509.400 291.600 511.200 302.700 ;
        RECT 512.400 291.600 514.200 303.600 ;
        RECT 518.550 295.050 519.450 311.550 ;
        RECT 523.950 310.950 526.050 313.050 ;
        RECT 527.100 311.100 528.900 311.850 ;
        RECT 529.950 310.950 532.200 313.050 ;
        RECT 533.100 311.100 534.900 311.850 ;
        RECT 524.100 309.150 525.900 309.900 ;
        RECT 526.950 307.950 529.050 310.050 ;
        RECT 530.100 306.900 531.150 309.900 ;
        RECT 532.950 307.950 535.050 310.050 ;
        RECT 539.550 307.050 540.450 319.950 ;
        RECT 548.400 317.100 549.600 320.400 ;
        RECT 547.950 313.950 550.050 316.050 ;
        RECT 569.100 315.000 570.900 323.400 ;
        RECT 589.200 316.200 591.000 323.400 ;
        RECT 566.700 313.350 570.900 315.000 ;
        RECT 587.400 315.300 591.000 316.200 ;
        RECT 548.700 309.900 549.900 312.900 ;
        RECT 550.950 312.450 553.050 313.050 ;
        RECT 550.950 311.550 558.450 312.450 ;
        RECT 550.950 310.950 553.050 311.550 ;
        RECT 545.100 309.150 546.900 309.900 ;
        RECT 529.950 303.600 531.150 306.900 ;
        RECT 538.950 304.950 541.050 307.050 ;
        RECT 548.700 304.650 550.050 309.900 ;
        RECT 551.100 309.150 552.900 309.900 ;
        RECT 548.700 303.600 551.400 304.650 ;
        RECT 517.950 292.950 520.050 295.050 ;
        RECT 529.500 291.600 531.300 303.600 ;
        RECT 549.600 291.600 551.400 303.600 ;
        RECT 557.550 298.050 558.450 311.550 ;
        RECT 566.700 308.100 567.600 313.350 ;
        RECT 569.100 311.100 570.900 311.850 ;
        RECT 575.100 311.100 576.900 311.850 ;
        RECT 587.400 311.100 588.600 315.300 ;
        RECT 595.950 313.950 598.050 316.050 ;
        RECT 608.100 315.000 609.900 323.400 ;
        RECT 625.800 317.400 627.600 323.400 ;
        RECT 568.950 307.950 571.050 310.050 ;
        RECT 574.950 307.950 577.050 310.050 ;
        RECT 584.100 308.100 585.900 308.850 ;
        RECT 586.950 307.950 589.200 310.050 ;
        RECT 590.100 308.100 591.900 308.850 ;
        RECT 596.550 307.050 597.450 313.950 ;
        RECT 605.700 313.350 609.900 315.000 ;
        RECT 626.400 315.300 627.600 317.400 ;
        RECT 628.800 318.300 630.600 323.400 ;
        RECT 634.800 318.300 636.600 323.400 ;
        RECT 640.950 319.950 643.050 322.050 ;
        RECT 628.800 316.950 636.600 318.300 ;
        RECT 626.400 314.250 630.150 315.300 ;
        RECT 628.950 314.100 630.150 314.250 ;
        RECT 605.700 308.100 606.600 313.350 ;
        RECT 608.100 311.100 609.900 311.850 ;
        RECT 614.100 311.100 615.900 311.850 ;
        RECT 626.100 311.100 627.900 311.850 ;
        RECT 628.950 310.950 631.050 313.050 ;
        RECT 632.100 311.100 633.900 311.850 ;
        RECT 634.950 310.950 637.050 313.050 ;
        RECT 607.800 307.950 610.050 310.050 ;
        RECT 613.950 307.950 616.050 310.050 ;
        RECT 625.950 307.950 628.050 310.050 ;
        RECT 562.950 304.950 568.050 307.050 ;
        RECT 571.950 304.950 574.050 307.050 ;
        RECT 583.950 304.950 586.050 307.050 ;
        RECT 566.700 298.800 567.600 303.900 ;
        RECT 572.100 303.150 573.900 303.900 ;
        RECT 556.950 295.950 559.050 298.050 ;
        RECT 566.700 297.900 573.300 298.800 ;
        RECT 566.700 297.600 567.600 297.900 ;
        RECT 565.800 291.600 567.600 297.600 ;
        RECT 571.800 297.600 573.300 297.900 ;
        RECT 587.400 297.600 588.600 306.900 ;
        RECT 589.950 304.950 592.050 307.050 ;
        RECT 595.950 304.950 598.050 307.050 ;
        RECT 604.950 304.950 607.050 307.050 ;
        RECT 610.950 304.950 613.050 307.050 ;
        RECT 629.850 306.900 630.900 309.900 ;
        RECT 631.950 307.950 634.050 310.050 ;
        RECT 635.100 309.150 636.900 309.900 ;
        RECT 605.700 298.800 606.600 303.900 ;
        RECT 611.100 303.150 612.900 303.900 ;
        RECT 629.850 303.600 631.050 306.900 ;
        RECT 605.700 297.900 612.300 298.800 ;
        RECT 605.700 297.600 606.600 297.900 ;
        RECT 571.800 291.600 573.600 297.600 ;
        RECT 587.400 291.600 589.200 297.600 ;
        RECT 604.800 291.600 606.600 297.600 ;
        RECT 610.800 297.600 612.300 297.900 ;
        RECT 610.800 291.600 612.600 297.600 ;
        RECT 629.700 291.600 631.500 303.600 ;
        RECT 641.550 298.050 642.450 319.950 ;
        RECT 646.800 317.400 648.600 323.400 ;
        RECT 647.400 315.300 648.600 317.400 ;
        RECT 649.800 318.300 651.600 323.400 ;
        RECT 655.800 318.300 657.600 323.400 ;
        RECT 669.300 319.200 671.100 323.400 ;
        RECT 649.800 316.950 657.600 318.300 ;
        RECT 669.150 317.400 671.100 319.200 ;
        RECT 647.400 314.250 651.150 315.300 ;
        RECT 649.950 314.100 651.150 314.250 ;
        RECT 669.150 314.100 670.050 317.400 ;
        RECT 671.100 315.900 672.900 316.500 ;
        RECT 676.800 315.900 678.600 323.400 ;
        RECT 686.400 318.300 688.200 323.400 ;
        RECT 692.400 318.300 694.200 323.400 ;
        RECT 686.400 316.950 694.200 318.300 ;
        RECT 695.400 317.400 697.200 323.400 ;
        RECT 700.950 319.950 703.050 322.050 ;
        RECT 671.100 314.700 678.600 315.900 ;
        RECT 695.400 315.300 696.600 317.400 ;
        RECT 647.100 311.100 648.900 311.850 ;
        RECT 649.950 310.950 652.050 313.050 ;
        RECT 653.100 311.100 654.900 311.850 ;
        RECT 655.950 310.950 658.050 313.050 ;
        RECT 667.950 312.450 670.050 313.050 ;
        RECT 662.550 312.000 670.050 312.450 ;
        RECT 661.950 311.550 670.050 312.000 ;
        RECT 646.950 307.950 649.050 310.050 ;
        RECT 650.850 306.900 651.900 309.900 ;
        RECT 652.950 307.950 655.050 310.050 ;
        RECT 656.100 309.150 657.900 309.900 ;
        RECT 661.950 307.950 664.050 311.550 ;
        RECT 667.950 310.950 670.050 311.550 ;
        RECT 671.100 311.100 672.900 311.850 ;
        RECT 650.850 303.600 652.050 306.900 ;
        RECT 667.950 303.600 669.000 309.900 ;
        RECT 670.950 307.950 673.050 310.050 ;
        RECT 640.950 295.950 643.050 298.050 ;
        RECT 650.700 291.600 652.500 303.600 ;
        RECT 667.200 291.600 669.000 303.600 ;
        RECT 674.550 297.600 675.600 314.700 ;
        RECT 692.850 314.250 696.600 315.300 ;
        RECT 692.850 314.100 694.050 314.250 ;
        RECT 676.950 310.950 679.050 313.050 ;
        RECT 685.950 310.950 688.050 313.050 ;
        RECT 689.100 311.100 690.900 311.850 ;
        RECT 691.950 310.950 694.050 313.050 ;
        RECT 695.100 311.100 696.900 311.850 ;
        RECT 677.100 309.150 678.900 309.900 ;
        RECT 686.100 309.150 687.900 309.900 ;
        RECT 688.950 307.950 691.050 310.050 ;
        RECT 692.100 306.900 693.150 309.900 ;
        RECT 694.950 307.950 697.050 310.050 ;
        RECT 691.950 303.600 693.150 306.900 ;
        RECT 673.800 291.600 675.600 297.600 ;
        RECT 691.500 291.600 693.300 303.600 ;
        RECT 701.550 301.050 702.450 319.950 ;
        RECT 712.200 316.200 714.000 323.400 ;
        RECT 710.400 315.300 714.000 316.200 ;
        RECT 729.000 316.200 730.800 323.400 ;
        RECT 745.800 317.400 747.600 323.400 ;
        RECT 729.000 315.300 732.600 316.200 ;
        RECT 710.400 311.100 711.600 315.300 ;
        RECT 721.950 310.950 724.050 313.050 ;
        RECT 731.400 311.100 732.600 315.300 ;
        RECT 746.400 315.300 747.600 317.400 ;
        RECT 748.800 318.300 750.600 323.400 ;
        RECT 754.800 318.300 756.600 323.400 ;
        RECT 748.800 316.950 756.600 318.300 ;
        RECT 764.400 318.300 766.200 323.400 ;
        RECT 770.400 318.300 772.200 323.400 ;
        RECT 764.400 316.950 772.200 318.300 ;
        RECT 773.400 317.400 775.200 323.400 ;
        RECT 785.400 318.300 787.200 323.400 ;
        RECT 791.400 318.300 793.200 323.400 ;
        RECT 773.400 315.300 774.600 317.400 ;
        RECT 785.400 316.950 793.200 318.300 ;
        RECT 794.400 317.400 796.200 323.400 ;
        RECT 810.300 319.200 812.100 323.400 ;
        RECT 794.400 315.300 795.600 317.400 ;
        RECT 799.800 316.950 801.900 319.050 ;
        RECT 810.150 317.400 812.100 319.200 ;
        RECT 746.400 314.250 750.150 315.300 ;
        RECT 748.950 314.100 750.150 314.250 ;
        RECT 770.850 314.250 774.600 315.300 ;
        RECT 791.850 314.250 795.600 315.300 ;
        RECT 770.850 314.100 772.050 314.250 ;
        RECT 791.850 314.100 793.050 314.250 ;
        RECT 800.550 313.050 801.450 316.950 ;
        RECT 810.150 314.100 811.050 317.400 ;
        RECT 812.100 315.900 813.900 316.500 ;
        RECT 817.800 315.900 819.600 323.400 ;
        RECT 812.100 314.700 819.600 315.900 ;
        RECT 827.400 315.900 829.200 323.400 ;
        RECT 834.900 319.200 836.700 323.400 ;
        RECT 841.950 319.950 844.050 322.050 ;
        RECT 834.900 317.400 836.850 319.200 ;
        RECT 833.100 315.900 834.900 316.500 ;
        RECT 827.400 314.700 834.900 315.900 ;
        RECT 746.100 311.100 747.900 311.850 ;
        RECT 748.950 310.950 751.050 313.050 ;
        RECT 752.100 311.100 753.900 311.850 ;
        RECT 754.950 310.950 757.050 313.050 ;
        RECT 763.950 310.950 766.050 313.050 ;
        RECT 767.100 311.100 768.900 311.850 ;
        RECT 769.950 310.950 772.050 313.050 ;
        RECT 773.100 311.100 774.900 311.850 ;
        RECT 784.800 310.950 787.050 313.050 ;
        RECT 788.100 311.100 789.900 311.850 ;
        RECT 790.800 310.950 793.050 313.050 ;
        RECT 794.100 311.100 795.900 311.850 ;
        RECT 799.950 310.950 802.050 313.050 ;
        RECT 808.950 312.450 811.050 313.050 ;
        RECT 803.550 311.550 811.050 312.450 ;
        RECT 707.100 308.100 708.900 308.850 ;
        RECT 709.950 307.950 712.050 310.050 ;
        RECT 713.100 308.100 714.900 308.850 ;
        RECT 701.550 299.550 706.050 301.050 ;
        RECT 702.000 298.950 706.050 299.550 ;
        RECT 710.400 297.600 711.600 306.900 ;
        RECT 712.950 304.950 715.050 307.050 ;
        RECT 718.800 304.950 720.900 307.050 ;
        RECT 710.400 291.600 712.200 297.600 ;
        RECT 719.550 295.050 720.450 304.950 ;
        RECT 722.550 304.050 723.450 310.950 ;
        RECT 728.100 308.100 729.900 308.850 ;
        RECT 730.950 307.950 733.050 310.050 ;
        RECT 734.100 308.100 735.900 308.850 ;
        RECT 745.950 307.950 748.050 310.050 ;
        RECT 727.800 304.950 730.050 307.050 ;
        RECT 749.850 306.900 750.900 309.900 ;
        RECT 751.950 307.950 754.050 310.050 ;
        RECT 755.100 309.150 756.900 309.900 ;
        RECT 764.100 309.150 765.900 309.900 ;
        RECT 766.950 307.950 769.050 310.050 ;
        RECT 770.100 306.900 771.150 309.900 ;
        RECT 772.950 307.950 775.200 310.050 ;
        RECT 785.100 309.150 786.900 309.900 ;
        RECT 787.950 307.950 790.050 310.050 ;
        RECT 721.950 301.950 724.050 304.050 ;
        RECT 727.950 301.950 730.050 304.950 ;
        RECT 731.400 297.600 732.600 306.900 ;
        RECT 749.850 303.600 751.050 306.900 ;
        RECT 769.950 303.600 771.150 306.900 ;
        RECT 718.950 292.950 721.050 295.050 ;
        RECT 730.800 291.600 732.600 297.600 ;
        RECT 749.700 291.600 751.500 303.600 ;
        RECT 769.500 291.600 771.300 303.600 ;
        RECT 773.550 301.050 774.450 307.950 ;
        RECT 791.100 306.900 792.150 309.900 ;
        RECT 793.950 307.950 796.050 310.050 ;
        RECT 803.550 307.050 804.450 311.550 ;
        RECT 808.950 310.950 811.050 311.550 ;
        RECT 812.100 311.100 813.900 311.850 ;
        RECT 790.950 303.600 792.150 306.900 ;
        RECT 802.950 304.950 805.050 307.050 ;
        RECT 808.950 303.600 810.000 309.900 ;
        RECT 811.950 307.950 814.050 310.050 ;
        RECT 772.800 298.950 774.900 301.050 ;
        RECT 790.500 291.600 792.300 303.600 ;
        RECT 808.200 291.600 810.000 303.600 ;
        RECT 815.550 297.600 816.600 314.700 ;
        RECT 817.950 310.950 820.050 313.050 ;
        RECT 826.950 310.950 829.050 313.050 ;
        RECT 818.100 309.150 819.900 309.900 ;
        RECT 827.100 309.150 828.900 309.900 ;
        RECT 814.800 291.600 816.600 297.600 ;
        RECT 830.400 297.600 831.450 314.700 ;
        RECT 835.950 314.100 836.850 317.400 ;
        RECT 835.950 312.450 838.050 313.050 ;
        RECT 842.550 312.450 843.450 319.950 ;
        RECT 833.100 311.100 834.900 311.850 ;
        RECT 835.950 311.550 843.450 312.450 ;
        RECT 835.950 310.950 838.050 311.550 ;
        RECT 832.950 307.950 835.050 310.050 ;
        RECT 837.000 303.600 838.050 309.900 ;
        RECT 830.400 291.600 832.200 297.600 ;
        RECT 837.000 291.600 838.800 303.600 ;
        RECT 842.550 298.050 843.450 311.550 ;
        RECT 850.950 304.950 853.050 307.050 ;
        RECT 851.550 298.050 852.450 304.950 ;
        RECT 853.950 301.950 856.050 304.050 ;
        RECT 841.950 295.950 844.050 298.050 ;
        RECT 850.950 295.950 853.050 298.050 ;
        RECT 854.550 295.050 855.450 301.950 ;
        RECT 852.000 294.900 855.450 295.050 ;
        RECT 850.950 293.400 855.450 294.900 ;
        RECT 850.950 292.950 855.000 293.400 ;
        RECT 850.950 292.800 853.050 292.950 ;
        RECT 10.800 275.400 12.600 287.400 ;
        RECT 13.800 276.300 15.600 287.400 ;
        RECT 19.800 276.300 21.600 287.400 ;
        RECT 32.400 281.400 34.200 287.400 ;
        RECT 32.700 281.100 34.200 281.400 ;
        RECT 38.400 281.400 40.200 287.400 ;
        RECT 43.950 283.950 46.050 286.050 ;
        RECT 38.400 281.100 39.300 281.400 ;
        RECT 32.700 280.200 39.300 281.100 ;
        RECT 13.800 275.400 21.600 276.300 ;
        RECT 11.400 269.100 12.300 275.400 ;
        RECT 32.100 275.100 33.900 275.850 ;
        RECT 38.400 275.100 39.300 280.200 ;
        RECT 31.950 271.950 34.050 274.050 ;
        RECT 37.950 273.450 40.050 274.050 ;
        RECT 44.550 273.450 45.450 283.950 ;
        RECT 55.500 275.400 57.300 287.400 ;
        RECT 37.950 272.550 45.450 273.450 ;
        RECT 37.950 271.950 40.050 272.550 ;
        RECT 55.950 272.100 57.150 275.400 ;
        RECT 64.950 274.950 67.050 277.050 ;
        RECT 76.500 275.400 78.300 287.400 ;
        RECT 95.400 281.400 97.200 287.400 ;
        RECT 95.700 281.100 97.200 281.400 ;
        RECT 101.400 281.400 103.200 287.400 ;
        RECT 116.400 281.400 118.200 287.400 ;
        RECT 101.400 281.100 102.300 281.400 ;
        RECT 95.700 280.200 102.300 281.100 ;
        RECT 116.700 281.100 118.200 281.400 ;
        RECT 122.400 281.400 124.200 287.400 ;
        RECT 137.400 281.400 139.200 287.400 ;
        RECT 122.400 281.100 123.300 281.400 ;
        RECT 116.700 280.200 123.300 281.100 ;
        RECT 137.700 281.100 139.200 281.400 ;
        RECT 143.400 281.400 145.200 287.400 ;
        RECT 143.400 281.100 144.300 281.400 ;
        RECT 137.700 280.200 144.300 281.100 ;
        RECT 13.950 268.950 16.050 271.050 ;
        RECT 17.100 269.100 18.900 269.850 ;
        RECT 19.800 268.950 22.050 271.050 ;
        RECT 28.950 268.950 31.050 271.050 ;
        RECT 34.950 268.950 37.050 271.050 ;
        RECT 10.950 265.950 13.050 268.050 ;
        RECT 14.100 267.150 15.900 267.900 ;
        RECT 16.800 265.950 19.050 268.050 ;
        RECT 20.100 267.150 21.900 267.900 ;
        RECT 29.100 267.150 30.900 267.900 ;
        RECT 35.100 267.150 36.900 267.900 ;
        RECT 38.400 265.650 39.300 270.900 ;
        RECT 50.100 269.100 51.900 269.850 ;
        RECT 52.950 268.950 55.200 271.050 ;
        RECT 56.100 269.100 57.150 272.100 ;
        RECT 58.950 268.950 61.050 271.050 ;
        RECT 65.550 268.050 66.450 274.950 ;
        RECT 76.950 272.100 78.150 275.400 ;
        RECT 95.100 275.100 96.900 275.850 ;
        RECT 101.400 275.100 102.300 280.200 ;
        RECT 116.100 275.100 117.900 275.850 ;
        RECT 122.400 275.100 123.300 280.200 ;
        RECT 137.100 275.100 138.900 275.850 ;
        RECT 143.400 275.100 144.300 280.200 ;
        RECT 155.400 276.300 157.200 287.400 ;
        RECT 161.400 276.300 163.200 287.400 ;
        RECT 155.400 275.400 163.200 276.300 ;
        RECT 164.400 275.400 166.200 287.400 ;
        RECT 169.950 280.950 172.050 283.050 ;
        RECT 71.100 269.100 72.900 269.850 ;
        RECT 73.950 268.950 76.050 271.050 ;
        RECT 77.100 269.100 78.150 272.100 ;
        RECT 94.950 271.950 97.050 274.050 ;
        RECT 100.950 273.450 103.050 274.050 ;
        RECT 100.950 272.550 108.450 273.450 ;
        RECT 100.950 271.950 103.050 272.550 ;
        RECT 79.950 268.950 82.050 271.050 ;
        RECT 91.950 268.950 94.050 271.050 ;
        RECT 97.950 268.950 100.050 271.050 ;
        RECT 49.950 265.950 52.050 268.050 ;
        RECT 53.100 267.150 54.900 267.900 ;
        RECT 55.950 265.950 58.050 268.050 ;
        RECT 59.100 267.150 60.900 267.900 ;
        RECT 64.950 265.950 67.050 268.050 ;
        RECT 70.950 265.950 73.050 268.050 ;
        RECT 74.100 267.150 75.900 267.900 ;
        RECT 76.950 265.950 79.050 268.050 ;
        RECT 80.100 267.150 81.900 267.900 ;
        RECT 85.950 265.950 88.050 268.050 ;
        RECT 92.100 267.150 93.900 267.900 ;
        RECT 98.100 267.150 99.900 267.900 ;
        RECT 11.400 261.600 12.300 264.900 ;
        RECT 35.100 264.000 39.300 265.650 ;
        RECT 56.850 264.750 58.050 264.900 ;
        RECT 77.850 264.750 79.050 264.900 ;
        RECT 11.400 259.950 16.800 261.600 ;
        RECT 15.000 255.600 16.800 259.950 ;
        RECT 35.100 255.600 36.900 264.000 ;
        RECT 56.850 263.700 60.600 264.750 ;
        RECT 77.850 263.700 81.600 264.750 ;
        RECT 50.400 260.700 58.200 262.050 ;
        RECT 50.400 255.600 52.200 260.700 ;
        RECT 56.400 255.600 58.200 260.700 ;
        RECT 59.400 261.600 60.600 263.700 ;
        RECT 59.400 255.600 61.200 261.600 ;
        RECT 71.400 260.700 79.200 262.050 ;
        RECT 71.400 255.600 73.200 260.700 ;
        RECT 77.400 255.600 79.200 260.700 ;
        RECT 80.400 261.600 81.600 263.700 ;
        RECT 86.550 262.050 87.450 265.950 ;
        RECT 101.400 265.650 102.300 270.900 ;
        RECT 98.100 264.000 102.300 265.650 ;
        RECT 80.400 255.600 82.200 261.600 ;
        RECT 85.950 259.950 88.050 262.050 ;
        RECT 98.100 255.600 99.900 264.000 ;
        RECT 107.550 262.050 108.450 272.550 ;
        RECT 115.950 271.950 118.050 274.050 ;
        RECT 121.950 273.450 124.050 274.050 ;
        RECT 121.950 272.550 129.450 273.450 ;
        RECT 121.950 271.950 124.050 272.550 ;
        RECT 112.950 268.950 115.050 271.050 ;
        RECT 118.950 268.950 121.050 271.050 ;
        RECT 113.100 267.150 114.900 267.900 ;
        RECT 119.100 267.150 120.900 267.900 ;
        RECT 122.400 265.650 123.300 270.900 ;
        RECT 119.100 264.000 123.300 265.650 ;
        RECT 106.950 259.950 109.050 262.050 ;
        RECT 119.100 255.600 120.900 264.000 ;
        RECT 128.550 259.050 129.450 272.550 ;
        RECT 136.950 271.950 139.050 274.050 ;
        RECT 142.950 273.450 145.050 274.050 ;
        RECT 147.000 273.450 151.050 274.050 ;
        RECT 142.950 272.550 151.050 273.450 ;
        RECT 142.950 271.950 145.050 272.550 ;
        RECT 147.000 271.950 151.050 272.550 ;
        RECT 133.950 268.950 136.050 271.050 ;
        RECT 139.950 268.950 142.050 271.050 ;
        RECT 134.100 267.150 135.900 267.900 ;
        RECT 140.100 267.150 141.900 267.900 ;
        RECT 143.400 265.650 144.300 270.900 ;
        RECT 154.950 268.950 157.050 271.050 ;
        RECT 158.100 269.100 159.900 269.850 ;
        RECT 160.950 268.950 163.050 271.050 ;
        RECT 164.700 269.100 165.600 275.400 ;
        RECT 155.100 267.150 156.900 267.900 ;
        RECT 157.800 265.950 160.050 268.050 ;
        RECT 161.100 267.150 162.900 267.900 ;
        RECT 163.950 265.950 169.050 268.050 ;
        RECT 140.100 264.000 144.300 265.650 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 140.100 255.600 141.900 264.000 ;
        RECT 164.700 261.600 165.600 264.900 ;
        RECT 170.550 262.050 171.450 280.950 ;
        RECT 181.500 275.400 183.300 287.400 ;
        RECT 193.950 283.950 196.050 286.050 ;
        RECT 181.950 272.100 183.150 275.400 ;
        RECT 176.100 269.100 177.900 269.850 ;
        RECT 178.950 268.950 181.050 271.050 ;
        RECT 182.100 269.100 183.150 272.100 ;
        RECT 184.950 268.950 187.050 271.050 ;
        RECT 175.950 265.950 178.050 268.050 ;
        RECT 179.100 267.150 180.900 267.900 ;
        RECT 181.950 265.950 184.050 268.050 ;
        RECT 185.100 267.150 186.900 267.900 ;
        RECT 194.550 267.450 195.450 283.950 ;
        RECT 199.800 275.400 201.600 287.400 ;
        RECT 202.800 276.300 204.600 287.400 ;
        RECT 208.800 276.300 210.600 287.400 ;
        RECT 220.800 281.400 222.600 287.400 ;
        RECT 202.800 275.400 210.600 276.300 ;
        RECT 200.400 269.100 201.300 275.400 ;
        RECT 221.400 272.100 222.600 281.400 ;
        RECT 235.200 275.400 237.000 287.400 ;
        RECT 241.800 281.400 243.600 287.400 ;
        RECT 202.950 268.950 205.050 271.050 ;
        RECT 206.100 269.100 207.900 269.850 ;
        RECT 208.950 268.950 211.050 271.050 ;
        RECT 217.950 268.950 223.050 271.050 ;
        RECT 235.950 269.100 237.000 275.400 ;
        RECT 238.950 268.950 241.050 271.050 ;
        RECT 199.950 267.450 202.050 268.050 ;
        RECT 194.550 266.550 202.050 267.450 ;
        RECT 203.100 267.150 204.900 267.900 ;
        RECT 199.950 265.950 202.050 266.550 ;
        RECT 205.950 265.950 208.050 268.050 ;
        RECT 209.100 267.150 210.900 267.900 ;
        RECT 182.850 264.750 184.050 264.900 ;
        RECT 182.850 263.700 186.600 264.750 ;
        RECT 160.200 259.950 165.600 261.600 ;
        RECT 169.950 259.950 172.050 262.050 ;
        RECT 176.400 260.700 184.200 262.050 ;
        RECT 160.200 255.600 162.000 259.950 ;
        RECT 176.400 255.600 178.200 260.700 ;
        RECT 182.400 255.600 184.200 260.700 ;
        RECT 185.400 261.600 186.600 263.700 ;
        RECT 200.400 261.600 201.300 264.900 ;
        RECT 185.400 255.600 187.200 261.600 ;
        RECT 200.400 259.950 205.800 261.600 ;
        RECT 204.000 255.600 205.800 259.950 ;
        RECT 221.400 258.600 222.600 267.900 ;
        RECT 224.100 266.100 225.900 266.850 ;
        RECT 232.950 265.950 238.050 268.050 ;
        RECT 239.100 267.150 240.900 267.900 ;
        RECT 223.950 262.950 226.050 265.050 ;
        RECT 229.950 262.950 232.050 265.050 ;
        RECT 230.550 259.050 231.450 262.950 ;
        RECT 237.150 261.600 238.050 264.900 ;
        RECT 242.550 264.300 243.600 281.400 ;
        RECT 257.400 281.400 259.200 287.400 ;
        RECT 253.950 271.950 256.050 274.050 ;
        RECT 257.400 272.100 258.600 281.400 ;
        RECT 266.100 277.950 268.200 280.050 ;
        RECT 259.950 271.950 262.050 274.050 ;
        RECT 254.100 270.150 255.900 270.900 ;
        RECT 245.100 269.100 246.900 269.850 ;
        RECT 256.950 268.950 259.050 271.050 ;
        RECT 260.100 270.150 261.900 270.900 ;
        RECT 244.950 265.950 247.050 268.050 ;
        RECT 239.100 263.100 246.600 264.300 ;
        RECT 239.100 262.500 240.900 263.100 ;
        RECT 237.150 259.800 239.100 261.600 ;
        RECT 220.800 255.600 222.600 258.600 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 237.300 255.600 239.100 259.800 ;
        RECT 244.800 255.600 246.600 263.100 ;
        RECT 257.400 263.700 258.600 267.900 ;
        RECT 257.400 262.800 261.000 263.700 ;
        RECT 259.200 255.600 261.000 262.800 ;
        RECT 266.550 262.050 267.450 277.950 ;
        RECT 276.300 276.900 278.100 287.400 ;
        RECT 275.700 275.400 278.100 276.900 ;
        RECT 283.800 275.400 285.600 287.400 ;
        RECT 275.700 272.100 277.050 275.400 ;
        RECT 278.400 274.200 279.300 274.350 ;
        RECT 284.400 274.200 285.600 275.400 ;
        RECT 278.400 273.000 285.600 274.200 ;
        RECT 296.400 281.400 298.200 287.400 ;
        RECT 307.950 283.950 310.050 286.050 ;
        RECT 278.400 272.400 280.200 273.000 ;
        RECT 271.950 268.950 277.050 271.050 ;
        RECT 265.950 259.950 268.050 262.050 ;
        RECT 274.950 261.600 276.000 267.900 ;
        RECT 278.400 264.600 279.300 272.400 ;
        RECT 292.950 271.950 295.050 274.050 ;
        RECT 296.400 272.100 297.600 281.400 ;
        RECT 298.950 271.950 301.050 274.050 ;
        RECT 293.100 270.150 294.900 270.900 ;
        RECT 281.100 269.100 282.900 269.850 ;
        RECT 295.800 268.950 298.050 271.050 ;
        RECT 299.100 270.150 300.900 270.900 ;
        RECT 280.950 265.950 283.050 268.050 ;
        RECT 284.100 266.100 285.900 266.850 ;
        RECT 278.250 263.700 280.050 264.600 ;
        RECT 278.250 262.800 281.700 263.700 ;
        RECT 283.950 262.950 286.200 265.050 ;
        RECT 296.400 263.700 297.600 267.900 ;
        RECT 296.400 262.800 300.000 263.700 ;
        RECT 274.800 255.600 276.600 261.600 ;
        RECT 280.800 258.600 281.700 262.800 ;
        RECT 280.800 255.600 282.600 258.600 ;
        RECT 298.200 255.600 300.000 262.800 ;
        RECT 308.550 259.050 309.450 283.950 ;
        RECT 317.700 275.400 319.500 287.400 ;
        RECT 336.600 275.400 338.400 287.400 ;
        RECT 355.500 275.400 357.300 287.400 ;
        RECT 375.600 275.400 377.400 287.400 ;
        RECT 317.850 272.100 319.050 275.400 ;
        RECT 336.600 274.350 339.300 275.400 ;
        RECT 313.950 268.950 316.050 271.050 ;
        RECT 317.850 269.100 318.900 272.100 ;
        RECT 319.950 268.950 322.050 271.050 ;
        RECT 323.100 269.100 324.900 269.850 ;
        RECT 335.100 269.100 336.900 269.850 ;
        RECT 337.950 269.100 339.300 274.350 ;
        RECT 355.950 272.100 357.150 275.400 ;
        RECT 341.100 269.100 342.900 269.850 ;
        RECT 350.100 269.100 351.900 269.850 ;
        RECT 314.100 267.150 315.900 267.900 ;
        RECT 316.950 265.950 319.050 268.050 ;
        RECT 320.100 267.150 321.900 267.900 ;
        RECT 322.950 265.950 325.050 268.050 ;
        RECT 334.950 265.950 337.050 268.050 ;
        RECT 338.100 266.100 339.300 269.100 ;
        RECT 352.950 268.950 355.050 271.050 ;
        RECT 356.100 269.100 357.150 272.100 ;
        RECT 374.700 274.350 377.400 275.400 ;
        RECT 392.400 281.400 394.200 287.400 ;
        RECT 409.800 281.400 411.600 287.400 ;
        RECT 427.800 281.400 429.600 287.400 ;
        RECT 358.950 268.950 361.050 271.050 ;
        RECT 371.100 269.100 372.900 269.850 ;
        RECT 374.700 269.100 376.050 274.350 ;
        RECT 382.950 271.950 385.050 274.050 ;
        RECT 388.950 271.950 391.050 274.050 ;
        RECT 392.400 272.100 393.600 281.400 ;
        RECT 394.950 271.950 397.050 274.050 ;
        RECT 410.400 272.100 411.600 281.400 ;
        RECT 424.950 276.000 427.050 280.050 ;
        RECT 425.550 274.050 426.450 276.000 ;
        RECT 424.950 271.950 427.050 274.050 ;
        RECT 428.400 272.100 429.600 281.400 ;
        RECT 442.800 275.400 444.600 287.400 ;
        RECT 445.800 276.300 447.600 287.400 ;
        RECT 451.800 276.300 453.600 287.400 ;
        RECT 445.800 275.400 453.600 276.300 ;
        RECT 463.800 286.500 471.600 287.400 ;
        RECT 463.800 275.400 465.600 286.500 ;
        RECT 430.950 271.950 433.050 274.050 ;
        RECT 436.950 271.950 439.050 274.050 ;
        RECT 377.100 269.100 378.900 269.850 ;
        RECT 340.950 265.950 343.050 268.050 ;
        RECT 346.950 265.950 352.050 268.050 ;
        RECT 353.100 267.150 354.900 267.900 ;
        RECT 355.800 265.950 358.050 268.050 ;
        RECT 359.100 267.150 360.900 267.900 ;
        RECT 370.950 265.950 373.050 268.050 ;
        RECT 374.700 266.100 375.900 269.100 ;
        RECT 383.550 268.050 384.450 271.950 ;
        RECT 389.100 270.150 390.900 270.900 ;
        RECT 391.950 268.950 394.050 271.050 ;
        RECT 395.100 270.150 396.900 270.900 ;
        RECT 409.950 268.950 412.050 271.050 ;
        RECT 418.950 268.950 421.050 271.050 ;
        RECT 425.100 270.150 426.900 270.900 ;
        RECT 427.800 268.950 430.050 271.050 ;
        RECT 431.100 270.150 432.900 270.900 ;
        RECT 376.950 265.950 379.050 268.050 ;
        RECT 382.950 265.950 385.050 268.050 ;
        RECT 316.950 264.750 318.150 264.900 ;
        RECT 314.400 263.700 318.150 264.750 ;
        RECT 314.400 261.600 315.600 263.700 ;
        RECT 337.950 262.950 340.050 265.050 ;
        RECT 356.850 264.750 358.050 264.900 ;
        RECT 356.850 263.700 360.600 264.750 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 313.800 255.600 315.600 261.600 ;
        RECT 316.800 260.700 324.600 262.050 ;
        RECT 316.800 255.600 318.600 260.700 ;
        RECT 322.800 255.600 324.600 260.700 ;
        RECT 338.400 258.600 339.600 261.900 ;
        RECT 337.800 255.600 339.600 258.600 ;
        RECT 350.400 260.700 358.200 262.050 ;
        RECT 350.400 255.600 352.200 260.700 ;
        RECT 356.400 255.600 358.200 260.700 ;
        RECT 359.400 261.600 360.600 263.700 ;
        RECT 373.950 262.950 376.050 265.050 ;
        RECT 392.400 263.700 393.600 267.900 ;
        RECT 392.400 262.800 396.000 263.700 ;
        RECT 359.400 255.600 361.200 261.600 ;
        RECT 374.400 258.600 375.600 261.900 ;
        RECT 374.400 255.600 376.200 258.600 ;
        RECT 394.200 255.600 396.000 262.800 ;
        RECT 410.400 258.600 411.600 267.900 ;
        RECT 413.100 266.100 414.900 266.850 ;
        RECT 412.950 262.950 415.050 265.050 ;
        RECT 419.550 262.050 420.450 268.950 ;
        RECT 437.550 268.050 438.450 271.950 ;
        RECT 443.400 269.100 444.300 275.400 ;
        RECT 466.800 274.500 468.600 285.600 ;
        RECT 469.800 276.600 471.600 286.500 ;
        RECT 475.800 276.600 477.600 287.400 ;
        RECT 478.950 283.950 481.050 286.050 ;
        RECT 469.800 275.700 477.600 276.600 ;
        RECT 457.950 271.950 460.050 274.050 ;
        RECT 466.800 273.600 470.850 274.500 ;
        RECT 479.550 274.050 480.450 283.950 ;
        RECT 488.400 281.400 490.200 287.400 ;
        RECT 469.950 272.100 470.850 273.600 ;
        RECT 445.950 268.950 448.050 271.050 ;
        RECT 449.100 269.100 450.900 269.850 ;
        RECT 451.950 268.950 454.050 271.050 ;
        RECT 458.550 268.050 459.450 271.950 ;
        RECT 464.100 269.100 465.900 269.850 ;
        RECT 466.950 268.950 469.050 271.050 ;
        RECT 470.100 269.100 470.850 272.100 ;
        RECT 478.800 271.950 480.900 274.050 ;
        RECT 484.950 271.950 487.050 274.050 ;
        RECT 488.400 272.100 489.600 281.400 ;
        RECT 507.600 275.400 509.400 287.400 ;
        RECT 525.600 275.400 527.400 287.400 ;
        RECT 535.950 283.950 538.050 286.050 ;
        RECT 506.700 274.350 509.400 275.400 ;
        RECT 524.700 274.350 527.400 275.400 ;
        RECT 490.950 271.950 493.050 274.050 ;
        RECT 472.950 268.950 475.050 271.050 ;
        RECT 485.100 270.150 486.900 270.900 ;
        RECT 476.100 269.100 477.750 269.850 ;
        RECT 487.950 268.950 490.050 271.050 ;
        RECT 491.100 270.150 492.900 270.900 ;
        RECT 503.100 269.100 504.900 269.850 ;
        RECT 506.700 269.100 508.050 274.350 ;
        RECT 514.950 271.950 517.050 274.050 ;
        RECT 509.100 269.100 510.900 269.850 ;
        RECT 428.400 263.700 429.600 267.900 ;
        RECT 436.950 265.950 439.050 268.050 ;
        RECT 442.950 265.950 445.050 268.050 ;
        RECT 446.100 267.150 447.900 267.900 ;
        RECT 426.000 262.800 429.600 263.700 ;
        RECT 418.950 259.950 421.050 262.050 ;
        RECT 409.800 255.600 411.600 258.600 ;
        RECT 426.000 255.600 427.800 262.800 ;
        RECT 443.400 261.600 444.300 264.900 ;
        RECT 448.950 262.950 451.050 268.050 ;
        RECT 452.100 267.150 453.900 267.900 ;
        RECT 457.950 265.950 460.050 268.050 ;
        RECT 463.950 265.950 466.050 268.050 ;
        RECT 467.250 267.150 468.900 267.900 ;
        RECT 469.950 265.950 472.050 268.050 ;
        RECT 473.100 267.150 474.750 267.900 ;
        RECT 475.950 265.950 478.050 268.050 ;
        RECT 471.000 261.600 472.050 264.900 ;
        RECT 488.400 263.700 489.600 267.900 ;
        RECT 506.700 266.100 507.900 269.100 ;
        RECT 508.950 265.950 511.050 268.050 ;
        RECT 488.400 262.800 492.000 263.700 ;
        RECT 505.950 262.950 508.050 265.050 ;
        RECT 443.400 259.950 448.800 261.600 ;
        RECT 447.000 255.600 448.800 259.950 ;
        RECT 471.000 255.600 472.800 261.600 ;
        RECT 490.200 255.600 492.000 262.800 ;
        RECT 515.550 262.050 516.450 271.950 ;
        RECT 521.100 269.100 522.900 269.850 ;
        RECT 524.700 269.100 526.050 274.350 ;
        RECT 536.550 271.050 537.450 283.950 ;
        RECT 545.700 275.400 547.500 287.400 ;
        RECT 562.800 286.500 570.600 287.400 ;
        RECT 556.950 283.950 559.050 286.050 ;
        RECT 545.850 272.100 547.050 275.400 ;
        RECT 527.100 269.100 528.900 269.850 ;
        RECT 524.700 266.100 525.900 269.100 ;
        RECT 535.950 268.950 538.050 271.050 ;
        RECT 541.950 268.950 544.050 271.050 ;
        RECT 545.850 269.100 546.900 272.100 ;
        RECT 547.800 268.950 550.050 271.050 ;
        RECT 551.100 269.100 552.900 269.850 ;
        RECT 526.950 267.450 529.050 268.050 ;
        RECT 526.950 266.550 534.450 267.450 ;
        RECT 542.100 267.150 543.900 267.900 ;
        RECT 526.950 265.950 529.050 266.550 ;
        RECT 523.950 262.950 526.050 265.050 ;
        RECT 506.400 258.600 507.600 261.900 ;
        RECT 514.950 259.950 517.050 262.050 ;
        RECT 524.400 258.600 525.600 261.900 ;
        RECT 533.550 259.050 534.450 266.550 ;
        RECT 544.950 265.950 547.050 268.050 ;
        RECT 548.100 267.150 549.900 267.900 ;
        RECT 550.950 265.950 553.050 268.050 ;
        RECT 544.950 264.750 546.150 264.900 ;
        RECT 542.400 263.700 546.150 264.750 ;
        RECT 542.400 261.600 543.600 263.700 ;
        RECT 557.550 262.050 558.450 283.950 ;
        RECT 562.800 275.400 564.600 286.500 ;
        RECT 565.800 274.500 567.600 285.600 ;
        RECT 568.800 276.600 570.600 286.500 ;
        RECT 574.800 276.600 576.600 287.400 ;
        RECT 568.800 275.700 576.600 276.600 ;
        RECT 584.400 276.300 586.200 287.400 ;
        RECT 590.400 276.300 592.200 287.400 ;
        RECT 584.400 275.400 592.200 276.300 ;
        RECT 593.400 275.400 595.200 287.400 ;
        RECT 611.700 275.400 613.500 287.400 ;
        RECT 632.700 275.400 634.500 287.400 ;
        RECT 650.400 281.400 652.200 287.400 ;
        RECT 665.400 281.400 667.200 287.400 ;
        RECT 565.800 273.600 569.850 274.500 ;
        RECT 568.950 272.100 569.850 273.600 ;
        RECT 563.100 269.100 564.900 269.850 ;
        RECT 565.800 268.950 568.050 271.050 ;
        RECT 569.100 269.100 569.850 272.100 ;
        RECT 571.950 268.950 574.050 271.050 ;
        RECT 575.100 269.100 576.750 269.850 ;
        RECT 583.800 268.950 586.050 271.050 ;
        RECT 587.100 269.100 588.900 269.850 ;
        RECT 589.950 268.950 592.050 271.050 ;
        RECT 593.700 269.100 594.600 275.400 ;
        RECT 611.850 272.100 613.050 275.400 ;
        RECT 632.850 272.100 634.050 275.400 ;
        RECT 650.400 272.100 651.600 281.400 ;
        RECT 665.400 272.100 666.600 281.400 ;
        RECT 683.700 275.400 685.500 287.400 ;
        RECT 698.400 276.300 700.200 287.400 ;
        RECT 704.400 276.300 706.200 287.400 ;
        RECT 698.400 275.400 706.200 276.300 ;
        RECT 707.400 275.400 709.200 287.400 ;
        RECT 719.400 281.400 721.200 287.400 ;
        RECT 683.850 272.100 685.050 275.400 ;
        RECT 607.950 268.950 610.050 271.050 ;
        RECT 611.850 269.100 612.900 272.100 ;
        RECT 613.950 268.950 616.050 271.050 ;
        RECT 617.100 269.100 618.900 269.850 ;
        RECT 628.950 268.950 631.050 271.050 ;
        RECT 632.850 269.100 633.900 272.100 ;
        RECT 634.950 268.950 637.050 271.050 ;
        RECT 638.100 269.100 639.900 269.850 ;
        RECT 649.950 268.950 652.050 271.050 ;
        RECT 658.950 270.450 663.000 271.050 ;
        RECT 664.950 270.450 667.050 271.050 ;
        RECT 658.950 269.550 667.050 270.450 ;
        RECT 658.950 268.950 663.000 269.550 ;
        RECT 664.950 268.950 667.050 269.550 ;
        RECT 679.950 268.950 682.050 271.050 ;
        RECT 683.850 269.100 684.900 272.100 ;
        RECT 685.950 268.950 688.050 271.050 ;
        RECT 689.100 269.100 690.900 269.850 ;
        RECT 697.800 268.950 700.050 271.050 ;
        RECT 701.100 269.100 702.900 269.850 ;
        RECT 703.950 268.950 706.050 271.050 ;
        RECT 707.700 269.100 708.600 275.400 ;
        RECT 719.400 274.500 720.600 281.400 ;
        RECT 725.700 275.400 727.500 287.400 ;
        RECT 742.500 275.400 744.300 287.400 ;
        RECT 719.400 273.600 725.100 274.500 ;
        RECT 723.150 272.700 725.100 273.600 ;
        RECT 719.100 269.100 720.900 269.850 ;
        RECT 723.150 269.100 724.050 272.700 ;
        RECT 726.000 269.100 727.200 275.400 ;
        RECT 742.950 272.100 744.150 275.400 ;
        RECT 751.950 274.950 754.050 277.050 ;
        RECT 758.400 276.300 760.200 287.400 ;
        RECT 764.400 276.300 766.200 287.400 ;
        RECT 758.400 275.400 766.200 276.300 ;
        RECT 767.400 275.400 769.200 287.400 ;
        RECT 779.400 281.400 781.200 287.400 ;
        RECT 737.100 269.100 738.900 269.850 ;
        RECT 562.800 265.950 565.050 268.050 ;
        RECT 566.250 267.150 567.900 267.900 ;
        RECT 568.950 265.950 571.050 268.050 ;
        RECT 572.100 267.150 573.750 267.900 ;
        RECT 574.950 265.950 577.050 268.050 ;
        RECT 584.100 267.150 585.900 267.900 ;
        RECT 586.950 265.950 589.050 268.050 ;
        RECT 590.100 267.150 591.900 267.900 ;
        RECT 592.950 265.950 598.050 268.050 ;
        RECT 608.100 267.150 609.900 267.900 ;
        RECT 610.800 265.950 613.050 268.050 ;
        RECT 614.100 267.150 615.900 267.900 ;
        RECT 616.800 265.950 619.050 268.050 ;
        RECT 629.100 267.150 630.900 267.900 ;
        RECT 631.800 265.950 634.050 268.050 ;
        RECT 635.100 267.150 636.900 267.900 ;
        RECT 637.950 265.950 640.200 268.050 ;
        RECT 647.100 266.100 648.900 266.850 ;
        RECT 506.400 255.600 508.200 258.600 ;
        RECT 524.400 255.600 526.200 258.600 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 541.800 255.600 543.600 261.600 ;
        RECT 544.800 260.700 552.600 262.050 ;
        RECT 544.800 255.600 546.600 260.700 ;
        RECT 550.800 255.600 552.600 260.700 ;
        RECT 556.950 259.950 559.050 262.050 ;
        RECT 570.000 261.600 571.050 264.900 ;
        RECT 593.700 261.600 594.600 264.900 ;
        RECT 610.950 264.750 612.150 264.900 ;
        RECT 631.950 264.750 633.150 264.900 ;
        RECT 608.400 263.700 612.150 264.750 ;
        RECT 629.400 263.700 633.150 264.750 ;
        RECT 608.400 261.600 609.600 263.700 ;
        RECT 570.000 255.600 571.800 261.600 ;
        RECT 589.200 259.950 594.600 261.600 ;
        RECT 589.200 255.600 591.000 259.950 ;
        RECT 607.800 255.600 609.600 261.600 ;
        RECT 610.800 260.700 618.600 262.050 ;
        RECT 629.400 261.600 630.600 263.700 ;
        RECT 646.950 262.950 649.050 265.050 ;
        RECT 610.800 255.600 612.600 260.700 ;
        RECT 616.800 255.600 618.600 260.700 ;
        RECT 628.800 255.600 630.600 261.600 ;
        RECT 631.800 260.700 639.600 262.050 ;
        RECT 631.800 255.600 633.600 260.700 ;
        RECT 637.800 255.600 639.600 260.700 ;
        RECT 650.400 258.600 651.600 267.900 ;
        RECT 662.100 266.100 663.900 266.850 ;
        RECT 661.950 262.950 664.050 265.050 ;
        RECT 665.400 258.600 666.600 267.900 ;
        RECT 680.100 267.150 681.900 267.900 ;
        RECT 682.950 265.950 685.050 268.050 ;
        RECT 686.100 267.150 687.900 267.900 ;
        RECT 688.950 265.950 691.050 268.050 ;
        RECT 698.100 267.150 699.900 267.900 ;
        RECT 700.950 265.950 703.050 268.050 ;
        RECT 704.100 267.150 705.900 267.900 ;
        RECT 706.950 267.450 709.050 268.050 ;
        RECT 711.000 267.450 714.900 268.050 ;
        RECT 706.950 266.550 714.900 267.450 ;
        RECT 706.950 265.950 709.050 266.550 ;
        RECT 711.000 265.950 714.900 266.550 ;
        RECT 723.150 264.900 723.900 269.100 ;
        RECT 739.950 268.950 742.050 271.050 ;
        RECT 743.100 269.100 744.150 272.100 ;
        RECT 745.950 268.950 748.050 271.050 ;
        RECT 752.550 268.050 753.450 274.950 ;
        RECT 757.950 268.950 760.050 271.050 ;
        RECT 761.100 269.100 762.900 269.850 ;
        RECT 763.950 268.950 766.050 271.050 ;
        RECT 767.700 269.100 768.600 275.400 ;
        RECT 779.400 274.500 780.600 281.400 ;
        RECT 785.700 275.400 787.500 287.400 ;
        RECT 793.950 280.950 796.050 283.050 ;
        RECT 772.950 271.950 775.050 274.050 ;
        RECT 779.400 273.600 785.100 274.500 ;
        RECT 783.150 272.700 785.100 273.600 ;
        RECT 724.950 265.950 727.050 268.050 ;
        RECT 736.950 265.950 739.050 268.050 ;
        RECT 740.100 267.150 741.900 267.900 ;
        RECT 742.950 265.950 745.050 268.050 ;
        RECT 746.100 267.150 747.900 267.900 ;
        RECT 751.950 265.950 754.050 268.050 ;
        RECT 758.100 267.150 759.900 267.900 ;
        RECT 760.800 265.950 763.050 268.050 ;
        RECT 764.100 267.150 765.900 267.900 ;
        RECT 766.950 265.950 769.050 268.050 ;
        RECT 682.950 264.750 684.150 264.900 ;
        RECT 680.400 263.700 684.150 264.750 ;
        RECT 680.400 261.600 681.600 263.700 ;
        RECT 650.400 255.600 652.200 258.600 ;
        RECT 665.400 255.600 667.200 258.600 ;
        RECT 679.800 255.600 681.600 261.600 ;
        RECT 682.800 260.700 690.600 262.050 ;
        RECT 707.700 261.600 708.600 264.900 ;
        RECT 723.150 264.300 724.050 264.900 ;
        RECT 723.150 263.400 725.100 264.300 ;
        RECT 682.800 255.600 684.600 260.700 ;
        RECT 688.800 255.600 690.600 260.700 ;
        RECT 703.200 259.950 708.600 261.600 ;
        RECT 720.000 262.500 725.100 263.400 ;
        RECT 703.200 255.600 705.000 259.950 ;
        RECT 720.000 258.600 721.200 262.500 ;
        RECT 726.000 261.600 727.200 264.900 ;
        RECT 743.850 264.750 745.050 264.900 ;
        RECT 743.850 263.700 747.600 264.750 ;
        RECT 719.400 255.600 721.200 258.600 ;
        RECT 725.700 255.600 727.500 261.600 ;
        RECT 737.400 260.700 745.200 262.050 ;
        RECT 737.400 255.600 739.200 260.700 ;
        RECT 743.400 255.600 745.200 260.700 ;
        RECT 746.400 261.600 747.600 263.700 ;
        RECT 767.700 261.600 768.600 264.900 ;
        RECT 746.400 255.600 748.200 261.600 ;
        RECT 763.200 259.950 768.600 261.600 ;
        RECT 763.200 255.600 765.000 259.950 ;
        RECT 773.550 259.050 774.450 271.950 ;
        RECT 779.100 269.100 780.900 269.850 ;
        RECT 783.150 269.100 784.050 272.700 ;
        RECT 786.000 269.100 787.200 275.400 ;
        RECT 790.800 271.950 792.900 274.050 ;
        RECT 783.150 264.900 783.900 269.100 ;
        RECT 784.950 265.950 787.200 268.050 ;
        RECT 783.150 264.300 784.050 264.900 ;
        RECT 783.150 263.400 785.100 264.300 ;
        RECT 780.000 262.500 785.100 263.400 ;
        RECT 773.550 257.550 778.050 259.050 ;
        RECT 780.000 258.600 781.200 262.500 ;
        RECT 786.000 261.600 787.200 264.900 ;
        RECT 774.000 256.950 778.050 257.550 ;
        RECT 779.400 255.600 781.200 258.600 ;
        RECT 785.700 255.600 787.500 261.600 ;
        RECT 791.550 259.050 792.450 271.950 ;
        RECT 794.550 259.050 795.450 280.950 ;
        RECT 801.600 275.400 803.400 287.400 ;
        RECT 817.500 275.400 819.300 287.400 ;
        RECT 823.800 281.400 825.600 287.400 ;
        RECT 801.600 274.350 804.300 275.400 ;
        RECT 800.100 269.100 801.900 269.850 ;
        RECT 802.950 269.100 804.300 274.350 ;
        RECT 806.100 269.100 807.900 269.850 ;
        RECT 817.800 269.100 819.000 275.400 ;
        RECT 824.400 274.500 825.600 281.400 ;
        RECT 830.100 280.950 832.200 283.050 ;
        RECT 819.900 273.600 825.600 274.500 ;
        RECT 819.900 272.700 821.850 273.600 ;
        RECT 820.950 269.100 821.850 272.700 ;
        RECT 824.100 269.100 825.900 269.850 ;
        RECT 799.950 265.950 802.050 268.050 ;
        RECT 803.100 266.100 804.300 269.100 ;
        RECT 805.950 265.950 808.050 268.050 ;
        RECT 814.950 265.950 820.050 268.050 ;
        RECT 802.950 262.950 805.050 265.050 ;
        RECT 821.100 264.900 821.850 269.100 ;
        RECT 790.800 256.950 792.900 259.050 ;
        RECT 794.100 256.950 796.200 259.050 ;
        RECT 803.400 258.600 804.600 261.900 ;
        RECT 817.800 261.600 819.000 264.900 ;
        RECT 820.950 264.300 821.850 264.900 ;
        RECT 819.900 263.400 821.850 264.300 ;
        RECT 819.900 262.500 825.000 263.400 ;
        RECT 802.800 255.600 804.600 258.600 ;
        RECT 817.500 255.600 819.300 261.600 ;
        RECT 823.800 258.600 825.000 262.500 ;
        RECT 830.550 259.050 831.450 280.950 ;
        RECT 839.700 275.400 841.500 287.400 ;
        RECT 853.950 283.950 856.050 286.050 ;
        RECT 839.850 272.100 841.050 275.400 ;
        RECT 835.950 268.950 838.050 271.050 ;
        RECT 839.850 269.100 840.900 272.100 ;
        RECT 850.950 271.950 853.050 274.050 ;
        RECT 841.950 268.950 844.050 271.050 ;
        RECT 845.100 269.100 846.900 269.850 ;
        RECT 851.550 268.050 852.450 271.950 ;
        RECT 836.100 267.150 837.900 267.900 ;
        RECT 838.950 265.950 841.050 268.050 ;
        RECT 842.100 267.150 843.900 267.900 ;
        RECT 844.950 265.950 847.050 268.050 ;
        RECT 850.950 265.950 853.050 268.050 ;
        RECT 838.950 264.750 840.150 264.900 ;
        RECT 836.400 263.700 840.150 264.750 ;
        RECT 836.400 261.600 837.600 263.700 ;
        RECT 823.800 255.600 825.600 258.600 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 835.800 255.600 837.600 261.600 ;
        RECT 838.800 260.700 846.600 262.050 ;
        RECT 838.800 255.600 840.600 260.700 ;
        RECT 844.800 255.600 846.600 260.700 ;
        RECT 854.550 259.050 855.450 283.950 ;
        RECT 850.950 257.550 855.450 259.050 ;
        RECT 850.950 256.950 855.000 257.550 ;
        RECT 10.800 245.400 12.600 251.400 ;
        RECT 11.400 243.300 12.600 245.400 ;
        RECT 13.800 246.300 15.600 251.400 ;
        RECT 19.800 246.300 21.600 251.400 ;
        RECT 25.950 247.950 28.050 250.050 ;
        RECT 13.800 244.950 21.600 246.300 ;
        RECT 11.400 242.250 15.150 243.300 ;
        RECT 13.950 242.100 15.150 242.250 ;
        RECT 11.100 239.100 12.900 239.850 ;
        RECT 13.950 238.950 16.050 241.050 ;
        RECT 17.100 239.100 18.900 239.850 ;
        RECT 19.950 238.950 22.050 241.050 ;
        RECT 26.550 240.450 27.450 247.950 ;
        RECT 36.000 247.050 37.800 251.400 ;
        RECT 57.000 247.050 58.800 251.400 ;
        RECT 32.400 245.400 37.800 247.050 ;
        RECT 53.400 245.400 58.800 247.050 ;
        RECT 32.400 242.100 33.300 245.400 ;
        RECT 53.400 242.100 54.300 245.400 ;
        RECT 77.100 243.000 78.900 251.400 ;
        RECT 98.100 243.000 99.900 251.400 ;
        RECT 120.000 247.050 121.800 251.400 ;
        RECT 77.100 241.350 81.300 243.000 ;
        RECT 31.950 240.450 34.050 241.050 ;
        RECT 26.550 239.550 34.050 240.450 ;
        RECT 31.950 238.950 34.050 239.550 ;
        RECT 35.100 239.100 36.900 239.850 ;
        RECT 37.950 238.950 40.200 241.050 ;
        RECT 52.950 240.450 55.050 241.050 ;
        RECT 41.100 239.100 42.900 239.850 ;
        RECT 47.550 239.550 55.050 240.450 ;
        RECT 10.950 235.950 13.050 238.050 ;
        RECT 14.850 234.900 15.900 237.900 ;
        RECT 16.950 235.950 19.050 238.050 ;
        RECT 20.100 237.150 21.900 237.900 ;
        RECT 14.850 231.600 16.050 234.900 ;
        RECT 32.400 231.600 33.300 237.900 ;
        RECT 34.950 235.950 37.050 238.050 ;
        RECT 38.100 237.150 39.900 237.900 ;
        RECT 40.950 235.950 43.050 238.050 ;
        RECT 47.550 235.050 48.450 239.550 ;
        RECT 52.950 238.950 55.050 239.550 ;
        RECT 56.100 239.100 57.900 239.850 ;
        RECT 58.950 238.950 61.050 241.050 ;
        RECT 62.100 239.100 63.900 239.850 ;
        RECT 71.100 239.100 72.900 239.850 ;
        RECT 77.100 239.100 78.900 239.850 ;
        RECT 46.950 232.950 49.050 235.050 ;
        RECT 53.400 231.600 54.300 237.900 ;
        RECT 55.950 235.950 58.050 238.050 ;
        RECT 59.100 237.150 60.900 237.900 ;
        RECT 61.950 235.950 64.050 238.050 ;
        RECT 70.950 235.950 73.050 238.050 ;
        RECT 76.950 235.950 79.050 238.050 ;
        RECT 80.400 236.100 81.300 241.350 ;
        RECT 95.700 241.350 99.900 243.000 ;
        RECT 116.400 245.400 121.800 247.050 ;
        RECT 134.400 246.300 136.200 251.400 ;
        RECT 140.400 246.300 142.200 251.400 ;
        RECT 116.400 242.100 117.300 245.400 ;
        RECT 134.400 244.950 142.200 246.300 ;
        RECT 143.400 245.400 145.200 251.400 ;
        RECT 148.950 247.950 151.050 250.050 ;
        RECT 143.400 243.300 144.600 245.400 ;
        RECT 140.850 242.250 144.600 243.300 ;
        RECT 140.850 242.100 142.050 242.250 ;
        RECT 95.700 236.100 96.600 241.350 ;
        RECT 98.100 239.100 99.900 239.850 ;
        RECT 104.100 239.100 105.900 239.850 ;
        RECT 112.800 238.950 118.050 241.050 ;
        RECT 119.100 239.100 120.900 239.850 ;
        RECT 121.800 238.950 124.050 241.050 ;
        RECT 125.100 239.100 126.900 239.850 ;
        RECT 133.950 238.950 136.050 241.050 ;
        RECT 137.100 239.100 138.900 239.850 ;
        RECT 139.950 238.950 142.050 241.050 ;
        RECT 143.100 239.100 144.900 239.850 ;
        RECT 149.550 238.050 150.450 247.950 ;
        RECT 160.200 247.050 162.000 251.400 ;
        RECT 160.200 245.400 165.600 247.050 ;
        RECT 164.700 242.100 165.600 245.400 ;
        RECT 169.950 244.950 172.050 247.050 ;
        RECT 155.100 239.100 156.900 239.850 ;
        RECT 157.950 238.950 160.050 241.050 ;
        RECT 161.100 239.100 162.900 239.850 ;
        RECT 163.950 238.950 169.050 241.050 ;
        RECT 170.550 238.050 171.450 244.950 ;
        RECT 182.100 243.000 183.900 251.400 ;
        RECT 190.950 247.950 193.050 250.050 ;
        RECT 182.100 241.350 186.300 243.000 ;
        RECT 176.100 239.100 177.900 239.850 ;
        RECT 182.100 239.100 183.900 239.850 ;
        RECT 97.950 235.950 100.050 238.050 ;
        RECT 103.950 235.950 106.050 238.050 ;
        RECT 73.800 232.950 76.050 235.050 ;
        RECT 79.950 232.950 82.050 235.050 ;
        RECT 94.950 234.450 97.050 235.050 ;
        RECT 89.550 233.550 97.050 234.450 ;
        RECT 14.700 219.600 16.500 231.600 ;
        RECT 31.800 219.600 33.600 231.600 ;
        RECT 34.800 230.700 42.600 231.600 ;
        RECT 34.800 219.600 36.600 230.700 ;
        RECT 40.800 219.600 42.600 230.700 ;
        RECT 52.800 219.600 54.600 231.600 ;
        RECT 55.800 230.700 63.600 231.600 ;
        RECT 74.100 231.150 75.900 231.900 ;
        RECT 55.800 219.600 57.600 230.700 ;
        RECT 61.800 219.600 63.600 230.700 ;
        RECT 80.400 226.800 81.300 231.900 ;
        RECT 74.700 225.900 81.300 226.800 ;
        RECT 89.550 226.050 90.450 233.550 ;
        RECT 94.950 232.950 97.050 233.550 ;
        RECT 100.950 232.950 103.050 235.050 ;
        RECT 95.700 226.800 96.600 231.900 ;
        RECT 101.100 231.150 102.900 231.900 ;
        RECT 116.400 231.600 117.300 237.900 ;
        RECT 118.950 235.950 121.050 238.050 ;
        RECT 122.100 237.150 123.900 237.900 ;
        RECT 124.950 235.950 127.050 238.050 ;
        RECT 134.100 237.150 135.900 237.900 ;
        RECT 136.950 235.950 139.050 238.050 ;
        RECT 140.100 234.900 141.150 237.900 ;
        RECT 142.950 235.950 145.050 238.050 ;
        RECT 148.950 235.950 151.050 238.050 ;
        RECT 154.950 235.950 157.050 238.050 ;
        RECT 158.100 237.150 159.900 237.900 ;
        RECT 160.950 235.950 163.050 238.050 ;
        RECT 139.950 231.600 141.150 234.900 ;
        RECT 149.550 232.050 150.450 235.950 ;
        RECT 74.700 225.600 76.200 225.900 ;
        RECT 74.400 219.600 76.200 225.600 ;
        RECT 80.400 225.600 81.300 225.900 ;
        RECT 80.400 219.600 82.200 225.600 ;
        RECT 88.950 223.950 91.050 226.050 ;
        RECT 95.700 225.900 102.300 226.800 ;
        RECT 95.700 225.600 96.600 225.900 ;
        RECT 94.800 219.600 96.600 225.600 ;
        RECT 100.800 225.600 102.300 225.900 ;
        RECT 100.800 219.600 102.600 225.600 ;
        RECT 115.800 219.600 117.600 231.600 ;
        RECT 118.800 230.700 126.600 231.600 ;
        RECT 118.800 219.600 120.600 230.700 ;
        RECT 124.800 219.600 126.600 230.700 ;
        RECT 139.500 219.600 141.300 231.600 ;
        RECT 148.950 229.950 151.050 232.050 ;
        RECT 164.700 231.600 165.600 237.900 ;
        RECT 169.950 235.950 172.050 238.050 ;
        RECT 175.950 235.950 178.050 238.050 ;
        RECT 181.950 235.950 184.050 238.050 ;
        RECT 185.400 236.100 186.300 241.350 ;
        RECT 178.950 232.950 181.050 235.050 ;
        RECT 184.950 234.450 187.050 235.050 ;
        RECT 191.550 234.450 192.450 247.950 ;
        RECT 197.400 246.300 199.200 251.400 ;
        RECT 203.400 246.300 205.200 251.400 ;
        RECT 197.400 244.950 205.200 246.300 ;
        RECT 206.400 245.400 208.200 251.400 ;
        RECT 218.400 246.300 220.200 251.400 ;
        RECT 224.400 246.300 226.200 251.400 ;
        RECT 206.400 243.300 207.600 245.400 ;
        RECT 218.400 244.950 226.200 246.300 ;
        RECT 227.400 245.400 229.200 251.400 ;
        RECT 227.400 243.300 228.600 245.400 ;
        RECT 232.950 244.950 235.050 247.050 ;
        RECT 203.850 242.250 207.600 243.300 ;
        RECT 224.850 242.250 228.600 243.300 ;
        RECT 203.850 242.100 205.050 242.250 ;
        RECT 224.850 242.100 226.050 242.250 ;
        RECT 196.950 238.950 199.050 241.050 ;
        RECT 200.100 239.100 201.900 239.850 ;
        RECT 202.950 238.950 205.050 241.050 ;
        RECT 206.100 239.100 207.900 239.850 ;
        RECT 217.800 238.950 220.050 241.050 ;
        RECT 221.100 239.100 222.900 239.850 ;
        RECT 223.950 238.950 226.050 241.050 ;
        RECT 227.100 239.100 228.900 239.850 ;
        RECT 197.100 237.150 198.900 237.900 ;
        RECT 199.950 235.950 202.050 238.050 ;
        RECT 203.100 234.900 204.150 237.900 ;
        RECT 205.950 235.950 208.050 238.050 ;
        RECT 218.100 237.150 219.900 237.900 ;
        RECT 220.950 235.950 223.050 238.050 ;
        RECT 224.100 234.900 225.150 237.900 ;
        RECT 226.950 235.950 229.050 238.050 ;
        RECT 184.950 233.550 192.450 234.450 ;
        RECT 184.950 232.950 187.050 233.550 ;
        RECT 155.400 230.700 163.200 231.600 ;
        RECT 155.400 219.600 157.200 230.700 ;
        RECT 161.400 219.600 163.200 230.700 ;
        RECT 164.400 219.600 166.200 231.600 ;
        RECT 179.100 231.150 180.900 231.900 ;
        RECT 185.400 226.800 186.300 231.900 ;
        RECT 202.950 231.600 204.150 234.900 ;
        RECT 223.950 231.600 225.150 234.900 ;
        RECT 179.700 225.900 186.300 226.800 ;
        RECT 179.700 225.600 181.200 225.900 ;
        RECT 179.400 219.600 181.200 225.600 ;
        RECT 185.400 225.600 186.300 225.900 ;
        RECT 185.400 219.600 187.200 225.600 ;
        RECT 202.500 219.600 204.300 231.600 ;
        RECT 223.500 219.600 225.300 231.600 ;
        RECT 233.550 226.050 234.450 244.950 ;
        RECT 245.100 243.000 246.900 251.400 ;
        RECT 265.200 247.050 267.000 251.400 ;
        RECT 265.200 245.400 270.600 247.050 ;
        RECT 245.100 241.350 249.300 243.000 ;
        RECT 269.700 242.100 270.600 245.400 ;
        RECT 287.100 243.000 288.900 251.400 ;
        RECT 307.200 247.050 309.000 251.400 ;
        RECT 307.200 245.400 312.600 247.050 ;
        RECT 287.100 241.350 291.300 243.000 ;
        RECT 311.700 242.100 312.600 245.400 ;
        RECT 316.950 244.950 319.050 247.050 ;
        RECT 239.100 239.100 240.900 239.850 ;
        RECT 245.100 239.100 246.900 239.850 ;
        RECT 238.800 235.950 241.050 238.050 ;
        RECT 244.950 235.950 247.200 238.050 ;
        RECT 248.400 236.100 249.300 241.350 ;
        RECT 253.950 238.950 256.050 241.050 ;
        RECT 260.100 239.100 261.900 239.850 ;
        RECT 262.950 238.950 265.050 241.050 ;
        RECT 268.950 240.450 271.050 241.050 ;
        RECT 266.100 239.100 267.900 239.850 ;
        RECT 268.950 239.550 276.450 240.450 ;
        RECT 268.950 238.950 271.050 239.550 ;
        RECT 241.950 232.950 244.050 235.050 ;
        RECT 247.950 234.450 250.050 235.050 ;
        RECT 254.550 234.450 255.450 238.950 ;
        RECT 259.950 235.950 262.050 238.050 ;
        RECT 263.100 237.150 264.900 237.900 ;
        RECT 265.950 235.950 268.050 238.050 ;
        RECT 247.950 233.550 255.450 234.450 ;
        RECT 247.950 232.950 250.050 233.550 ;
        RECT 242.100 231.150 243.900 231.900 ;
        RECT 248.400 226.800 249.300 231.900 ;
        RECT 269.700 231.600 270.600 237.900 ;
        RECT 232.950 223.950 235.050 226.050 ;
        RECT 242.700 225.900 249.300 226.800 ;
        RECT 242.700 225.600 244.200 225.900 ;
        RECT 242.400 219.600 244.200 225.600 ;
        RECT 248.400 225.600 249.300 225.900 ;
        RECT 260.400 230.700 268.200 231.600 ;
        RECT 248.400 219.600 250.200 225.600 ;
        RECT 260.400 219.600 262.200 230.700 ;
        RECT 266.400 219.600 268.200 230.700 ;
        RECT 269.400 219.600 271.200 231.600 ;
        RECT 275.550 229.050 276.450 239.550 ;
        RECT 281.100 239.100 282.900 239.850 ;
        RECT 287.100 239.100 288.900 239.850 ;
        RECT 280.950 235.950 283.050 238.050 ;
        RECT 286.950 235.950 289.050 238.050 ;
        RECT 290.400 236.100 291.300 241.350 ;
        RECT 302.100 239.100 303.900 239.850 ;
        RECT 304.950 238.950 307.050 241.050 ;
        RECT 310.950 240.450 313.050 241.050 ;
        RECT 317.550 240.450 318.450 244.950 ;
        RECT 329.100 243.000 330.900 251.400 ;
        RECT 351.000 247.050 352.800 251.400 ;
        RECT 347.400 245.400 352.800 247.050 ;
        RECT 329.100 241.350 333.300 243.000 ;
        RECT 347.400 242.100 348.300 245.400 ;
        RECT 371.100 243.000 372.900 251.400 ;
        RECT 388.800 248.400 390.600 251.400 ;
        RECT 371.100 241.350 375.300 243.000 ;
        RECT 308.100 239.100 309.900 239.850 ;
        RECT 310.950 239.550 318.450 240.450 ;
        RECT 310.950 238.950 313.050 239.550 ;
        RECT 323.100 239.100 324.900 239.850 ;
        RECT 329.100 239.100 330.900 239.850 ;
        RECT 301.950 235.950 304.050 238.050 ;
        RECT 305.100 237.150 306.900 237.900 ;
        RECT 307.950 235.950 310.050 238.050 ;
        RECT 283.950 232.950 286.050 235.050 ;
        RECT 289.950 232.950 295.050 235.050 ;
        RECT 284.100 231.150 285.900 231.900 ;
        RECT 274.950 226.950 277.050 229.050 ;
        RECT 290.400 226.800 291.300 231.900 ;
        RECT 311.700 231.600 312.600 237.900 ;
        RECT 322.950 235.950 325.050 238.050 ;
        RECT 328.950 235.950 331.050 238.050 ;
        RECT 332.400 236.100 333.300 241.350 ;
        RECT 343.950 238.950 349.050 241.050 ;
        RECT 350.100 239.100 351.900 239.850 ;
        RECT 352.950 238.950 355.050 241.050 ;
        RECT 356.100 239.100 357.900 239.850 ;
        RECT 365.100 239.100 366.900 239.850 ;
        RECT 371.100 239.100 372.900 239.850 ;
        RECT 325.950 232.950 328.050 235.050 ;
        RECT 331.950 232.950 337.050 235.050 ;
        RECT 284.700 225.900 291.300 226.800 ;
        RECT 284.700 225.600 286.200 225.900 ;
        RECT 284.400 219.600 286.200 225.600 ;
        RECT 290.400 225.600 291.300 225.900 ;
        RECT 302.400 230.700 310.200 231.600 ;
        RECT 290.400 219.600 292.200 225.600 ;
        RECT 302.400 219.600 304.200 230.700 ;
        RECT 308.400 219.600 310.200 230.700 ;
        RECT 311.400 219.600 313.200 231.600 ;
        RECT 326.100 231.150 327.900 231.900 ;
        RECT 332.400 226.800 333.300 231.900 ;
        RECT 347.400 231.600 348.300 237.900 ;
        RECT 349.950 235.950 352.050 238.050 ;
        RECT 353.100 237.150 354.900 237.900 ;
        RECT 355.950 235.950 358.050 238.050 ;
        RECT 364.950 235.950 367.050 238.050 ;
        RECT 370.950 235.950 373.050 238.050 ;
        RECT 374.400 236.100 375.300 241.350 ;
        RECT 389.400 239.100 390.600 248.400 ;
        RECT 403.800 245.400 405.600 251.400 ;
        RECT 391.950 241.950 394.050 244.050 ;
        RECT 404.400 243.300 405.600 245.400 ;
        RECT 406.800 246.300 408.600 251.400 ;
        RECT 412.800 246.300 414.600 251.400 ;
        RECT 406.800 244.950 414.600 246.300 ;
        RECT 422.400 246.300 424.200 251.400 ;
        RECT 428.400 246.300 430.200 251.400 ;
        RECT 422.400 244.950 430.200 246.300 ;
        RECT 431.400 245.400 433.200 251.400 ;
        RECT 431.400 243.300 432.600 245.400 ;
        RECT 448.200 244.200 450.000 251.400 ;
        RECT 404.400 242.250 408.150 243.300 ;
        RECT 406.950 242.100 408.150 242.250 ;
        RECT 428.850 242.250 432.600 243.300 ;
        RECT 446.400 243.300 450.000 244.200 ;
        RECT 465.000 244.200 466.800 251.400 ;
        RECT 465.000 243.300 468.600 244.200 ;
        RECT 428.850 242.100 430.050 242.250 ;
        RECT 392.100 240.150 393.900 240.900 ;
        RECT 404.100 239.100 405.900 239.850 ;
        RECT 406.950 238.950 409.050 241.050 ;
        RECT 410.100 239.100 411.900 239.850 ;
        RECT 412.950 238.950 415.050 241.050 ;
        RECT 421.950 238.950 424.050 241.050 ;
        RECT 425.100 239.100 426.900 239.850 ;
        RECT 427.800 238.950 430.050 241.050 ;
        RECT 431.100 239.100 432.900 239.850 ;
        RECT 446.400 239.100 447.600 243.300 ;
        RECT 467.400 239.100 468.600 243.300 ;
        RECT 479.400 243.900 481.200 251.400 ;
        RECT 486.900 247.200 488.700 251.400 ;
        RECT 486.900 245.400 488.850 247.200 ;
        RECT 485.100 243.900 486.900 244.500 ;
        RECT 479.400 242.700 486.900 243.900 ;
        RECT 478.950 238.950 481.050 241.050 ;
        RECT 388.950 235.950 394.050 238.050 ;
        RECT 403.950 235.950 406.050 238.050 ;
        RECT 367.950 232.950 370.050 235.050 ;
        RECT 373.950 234.450 376.050 235.050 ;
        RECT 373.950 233.550 381.450 234.450 ;
        RECT 373.950 232.950 376.050 233.550 ;
        RECT 326.700 225.900 333.300 226.800 ;
        RECT 326.700 225.600 328.200 225.900 ;
        RECT 326.400 219.600 328.200 225.600 ;
        RECT 332.400 225.600 333.300 225.900 ;
        RECT 332.400 219.600 334.200 225.600 ;
        RECT 346.800 219.600 348.600 231.600 ;
        RECT 349.800 230.700 357.600 231.600 ;
        RECT 368.100 231.150 369.900 231.900 ;
        RECT 349.800 219.600 351.600 230.700 ;
        RECT 355.800 219.600 357.600 230.700 ;
        RECT 374.400 226.800 375.300 231.900 ;
        RECT 368.700 225.900 375.300 226.800 ;
        RECT 368.700 225.600 370.200 225.900 ;
        RECT 368.400 219.600 370.200 225.600 ;
        RECT 374.400 225.600 375.300 225.900 ;
        RECT 374.400 219.600 376.200 225.600 ;
        RECT 380.550 223.050 381.450 233.550 ;
        RECT 389.400 225.600 390.600 234.900 ;
        RECT 404.550 234.000 405.450 235.950 ;
        RECT 407.850 234.900 408.900 237.900 ;
        RECT 409.950 235.950 412.050 238.050 ;
        RECT 413.100 237.150 414.900 237.900 ;
        RECT 422.100 237.150 423.900 237.900 ;
        RECT 424.950 235.950 427.050 238.050 ;
        RECT 428.100 234.900 429.150 237.900 ;
        RECT 430.950 235.950 433.050 238.050 ;
        RECT 443.100 236.100 444.900 236.850 ;
        RECT 445.950 235.950 448.050 238.050 ;
        RECT 449.100 236.100 450.900 236.850 ;
        RECT 464.100 236.100 465.900 236.850 ;
        RECT 466.800 235.950 469.050 238.050 ;
        RECT 479.100 237.150 480.900 237.900 ;
        RECT 470.100 236.100 471.900 236.850 ;
        RECT 403.950 229.950 406.050 234.000 ;
        RECT 407.850 231.600 409.050 234.900 ;
        RECT 427.950 231.600 429.150 234.900 ;
        RECT 442.800 232.950 445.050 235.050 ;
        RECT 379.950 220.950 382.050 223.050 ;
        RECT 388.800 219.600 390.600 225.600 ;
        RECT 407.700 219.600 409.500 231.600 ;
        RECT 427.500 219.600 429.300 231.600 ;
        RECT 446.400 225.600 447.600 234.900 ;
        RECT 448.950 232.950 451.050 235.050 ;
        RECT 463.950 232.950 466.050 235.050 ;
        RECT 464.550 231.000 465.450 232.950 ;
        RECT 463.950 226.950 466.050 231.000 ;
        RECT 467.400 225.600 468.600 234.900 ;
        RECT 469.950 232.950 472.050 235.050 ;
        RECT 446.400 219.600 448.200 225.600 ;
        RECT 466.800 219.600 468.600 225.600 ;
        RECT 482.400 225.600 483.450 242.700 ;
        RECT 487.950 242.100 488.850 245.400 ;
        RECT 500.400 246.300 502.200 251.400 ;
        RECT 506.400 246.300 508.200 251.400 ;
        RECT 500.400 244.950 508.200 246.300 ;
        RECT 509.400 245.400 511.200 251.400 ;
        RECT 509.400 243.300 510.600 245.400 ;
        RECT 514.950 244.950 517.050 247.050 ;
        RECT 521.400 246.300 523.200 251.400 ;
        RECT 527.400 246.300 529.200 251.400 ;
        RECT 521.400 244.950 529.200 246.300 ;
        RECT 530.400 245.400 532.200 251.400 ;
        RECT 506.850 242.250 510.600 243.300 ;
        RECT 506.850 242.100 508.050 242.250 ;
        RECT 487.950 240.450 490.050 241.050 ;
        RECT 485.100 239.100 486.900 239.850 ;
        RECT 487.950 239.550 495.450 240.450 ;
        RECT 487.950 238.950 490.050 239.550 ;
        RECT 484.950 235.950 487.050 238.050 ;
        RECT 489.000 231.600 490.050 237.900 ;
        RECT 494.550 232.050 495.450 239.550 ;
        RECT 499.950 238.950 502.050 241.050 ;
        RECT 503.100 239.100 504.900 239.850 ;
        RECT 505.950 238.950 508.050 241.050 ;
        RECT 509.100 239.100 510.900 239.850 ;
        RECT 500.100 237.150 501.900 237.900 ;
        RECT 502.950 235.950 505.050 238.050 ;
        RECT 506.100 234.900 507.150 237.900 ;
        RECT 482.400 219.600 484.200 225.600 ;
        RECT 489.000 219.600 490.800 231.600 ;
        RECT 493.950 229.950 496.050 232.050 ;
        RECT 505.950 231.600 507.150 234.900 ;
        RECT 505.500 219.600 507.300 231.600 ;
        RECT 515.550 226.050 516.450 244.950 ;
        RECT 530.400 243.300 531.600 245.400 ;
        RECT 547.200 244.200 549.000 251.400 ;
        RECT 562.800 248.400 564.600 251.400 ;
        RECT 577.800 248.400 579.600 251.400 ;
        RECT 527.850 242.250 531.600 243.300 ;
        RECT 545.400 243.300 549.000 244.200 ;
        RECT 527.850 242.100 529.050 242.250 ;
        RECT 520.950 238.950 523.050 241.050 ;
        RECT 524.100 239.100 525.900 239.850 ;
        RECT 526.950 238.950 529.050 241.050 ;
        RECT 530.100 239.100 531.900 239.850 ;
        RECT 535.950 238.950 538.050 241.050 ;
        RECT 545.400 239.100 546.600 243.300 ;
        RECT 563.400 239.100 564.600 248.400 ;
        RECT 565.950 241.950 568.050 244.050 ;
        RECT 566.100 240.150 567.900 240.900 ;
        RECT 578.400 239.100 579.600 248.400 ;
        RECT 584.550 245.400 586.350 251.400 ;
        RECT 592.650 248.400 594.450 251.400 ;
        RECT 600.450 248.400 602.250 251.400 ;
        RECT 608.250 249.300 610.050 251.400 ;
        RECT 608.250 248.400 612.000 249.300 ;
        RECT 592.650 247.500 593.700 248.400 ;
        RECT 589.950 246.300 593.700 247.500 ;
        RECT 601.200 246.600 602.250 248.400 ;
        RECT 610.950 247.500 612.000 248.400 ;
        RECT 589.950 245.400 592.050 246.300 ;
        RECT 580.950 241.950 583.050 244.050 ;
        RECT 584.550 241.050 585.750 245.400 ;
        RECT 597.150 244.200 598.950 246.000 ;
        RECT 601.200 245.550 606.150 246.600 ;
        RECT 604.350 244.800 606.150 245.550 ;
        RECT 607.650 244.800 609.450 246.600 ;
        RECT 610.950 245.400 613.050 247.500 ;
        RECT 616.050 245.400 617.850 251.400 ;
        RECT 598.050 243.900 598.950 244.200 ;
        RECT 608.100 243.900 609.150 244.800 ;
        RECT 598.050 243.000 609.150 243.900 ;
        RECT 598.050 242.100 598.950 243.000 ;
        RECT 608.100 241.800 609.150 243.000 ;
        RECT 581.100 240.150 582.900 240.900 ;
        RECT 584.550 238.950 585.900 241.050 ;
        RECT 586.950 238.950 589.050 241.050 ;
        RECT 590.100 239.250 590.850 241.050 ;
        RECT 598.950 238.950 601.050 241.050 ;
        RECT 604.950 238.950 607.050 241.050 ;
        RECT 608.100 240.600 615.000 241.800 ;
        RECT 608.100 240.000 609.900 240.600 ;
        RECT 614.100 239.850 615.000 240.600 ;
        RECT 611.100 239.100 612.900 239.700 ;
        RECT 521.100 237.150 522.900 237.900 ;
        RECT 523.950 235.950 526.050 238.050 ;
        RECT 527.100 234.900 528.150 237.900 ;
        RECT 529.950 235.950 532.050 238.050 ;
        RECT 526.950 231.600 528.150 234.900 ;
        RECT 536.550 234.450 537.450 238.950 ;
        RECT 542.100 236.100 543.900 236.850 ;
        RECT 544.950 235.950 547.050 238.050 ;
        RECT 548.100 236.100 549.900 236.850 ;
        RECT 562.950 235.950 565.050 238.050 ;
        RECT 571.950 237.450 576.000 238.050 ;
        RECT 577.950 237.450 580.050 238.050 ;
        RECT 571.950 236.550 580.050 237.450 ;
        RECT 571.950 235.950 576.000 236.550 ;
        RECT 577.950 235.950 580.050 236.550 ;
        RECT 541.950 234.450 544.050 235.050 ;
        RECT 536.550 233.550 544.050 234.450 ;
        RECT 541.950 232.950 544.050 233.550 ;
        RECT 514.950 223.950 517.050 226.050 ;
        RECT 526.500 219.600 528.300 231.600 ;
        RECT 545.400 225.600 546.600 234.900 ;
        RECT 547.950 232.950 550.050 235.050 ;
        RECT 563.400 225.600 564.600 234.900 ;
        RECT 578.400 225.600 579.600 234.900 ;
        RECT 545.400 219.600 547.200 225.600 ;
        RECT 562.800 219.600 564.600 225.600 ;
        RECT 577.800 219.600 579.600 225.600 ;
        RECT 584.550 231.600 585.750 238.950 ;
        RECT 608.100 238.200 612.900 239.100 ;
        RECT 611.100 237.900 612.900 238.200 ;
        RECT 614.100 238.050 615.900 239.850 ;
        RECT 586.950 233.400 588.750 235.200 ;
        RECT 587.850 232.200 592.050 233.400 ;
        RECT 598.050 232.200 598.950 237.900 ;
        RECT 606.750 233.100 608.550 233.400 ;
        RECT 584.550 219.600 586.350 231.600 ;
        RECT 589.950 231.300 592.050 232.200 ;
        RECT 592.950 231.300 598.950 232.200 ;
        RECT 600.150 232.800 608.550 233.100 ;
        RECT 616.950 232.800 617.850 245.400 ;
        RECT 629.400 248.400 631.200 251.400 ;
        RECT 619.950 241.950 622.050 244.050 ;
        RECT 625.950 241.950 628.050 244.050 ;
        RECT 600.150 232.200 617.850 232.800 ;
        RECT 592.950 230.400 593.850 231.300 ;
        RECT 591.150 228.600 593.850 230.400 ;
        RECT 594.750 230.100 596.550 230.400 ;
        RECT 600.150 230.100 601.050 232.200 ;
        RECT 606.750 231.600 617.850 232.200 ;
        RECT 594.750 229.200 601.050 230.100 ;
        RECT 601.950 230.700 603.750 231.300 ;
        RECT 601.950 229.500 609.450 230.700 ;
        RECT 594.750 228.600 596.550 229.200 ;
        RECT 608.250 228.600 609.450 229.500 ;
        RECT 589.950 225.600 593.850 227.700 ;
        RECT 598.950 227.550 600.750 228.300 ;
        RECT 603.750 227.550 605.550 228.300 ;
        RECT 598.950 226.500 605.550 227.550 ;
        RECT 608.250 226.500 613.050 228.600 ;
        RECT 592.050 219.600 593.850 225.600 ;
        RECT 599.850 219.600 601.650 226.500 ;
        RECT 608.250 225.600 609.450 226.500 ;
        RECT 607.650 219.600 609.450 225.600 ;
        RECT 616.050 219.600 617.850 231.600 ;
        RECT 620.550 223.050 621.450 241.950 ;
        RECT 626.100 240.150 627.900 240.900 ;
        RECT 629.400 239.100 630.600 248.400 ;
        RECT 634.950 244.950 637.050 247.050 ;
        RECT 628.800 235.950 631.050 238.050 ;
        RECT 629.400 225.600 630.600 234.900 ;
        RECT 619.950 220.950 622.050 223.050 ;
        RECT 629.400 219.600 631.200 225.600 ;
        RECT 635.550 223.050 636.450 244.950 ;
        RECT 646.200 244.200 648.000 251.400 ;
        RECT 644.400 243.300 648.000 244.200 ;
        RECT 663.000 244.200 664.800 251.400 ;
        RECT 677.400 247.200 679.200 250.200 ;
        RECT 663.000 243.300 666.600 244.200 ;
        RECT 644.400 239.100 645.600 243.300 ;
        RECT 665.400 239.100 666.600 243.300 ;
        RECT 678.150 243.900 679.200 247.200 ;
        RECT 684.900 245.700 686.700 250.200 ;
        RECT 698.100 247.950 700.200 250.050 ;
        RECT 684.900 244.800 687.000 245.700 ;
        RECT 678.150 243.000 684.450 243.900 ;
        RECT 677.100 239.100 678.900 239.850 ;
        RECT 679.950 238.950 682.050 241.050 ;
        RECT 641.100 236.100 642.900 236.850 ;
        RECT 643.800 235.950 646.050 238.050 ;
        RECT 647.100 236.100 648.900 236.850 ;
        RECT 652.950 235.950 655.050 238.050 ;
        RECT 662.100 236.100 663.900 236.850 ;
        RECT 664.950 235.950 667.050 238.050 ;
        RECT 668.100 236.100 669.900 236.850 ;
        RECT 676.950 235.950 679.050 238.050 ;
        RECT 680.100 237.150 681.900 237.900 ;
        RECT 683.250 237.300 684.450 243.000 ;
        RECT 686.100 239.100 687.000 244.800 ;
        RECT 688.950 238.950 691.050 241.050 ;
        RECT 640.950 232.950 643.050 235.050 ;
        RECT 644.400 225.600 645.600 234.900 ;
        RECT 646.800 232.950 649.050 235.050 ;
        RECT 653.550 232.050 654.450 235.950 ;
        RECT 683.250 235.500 684.900 237.300 ;
        RECT 685.950 235.950 688.050 238.050 ;
        RECT 689.100 237.150 690.900 237.900 ;
        RECT 661.950 232.950 664.050 235.050 ;
        RECT 652.950 229.950 655.050 232.050 ;
        RECT 665.400 225.600 666.600 234.900 ;
        RECT 667.950 232.950 670.050 235.050 ;
        RECT 683.250 232.800 684.450 235.500 ;
        RECT 678.300 231.900 684.450 232.800 ;
        RECT 678.300 226.800 679.200 231.900 ;
        RECT 686.100 231.000 687.000 234.900 ;
        RECT 634.950 220.950 637.050 223.050 ;
        RECT 644.400 219.600 646.200 225.600 ;
        RECT 664.800 219.600 666.600 225.600 ;
        RECT 677.400 220.800 679.200 226.800 ;
        RECT 684.900 230.100 687.000 231.000 ;
        RECT 684.900 220.800 686.700 230.100 ;
        RECT 698.550 229.050 699.450 247.950 ;
        RECT 703.800 245.400 705.600 251.400 ;
        RECT 704.400 243.300 705.600 245.400 ;
        RECT 706.800 246.300 708.600 251.400 ;
        RECT 712.800 246.300 714.600 251.400 ;
        RECT 706.800 244.950 714.600 246.300 ;
        RECT 722.400 246.300 724.200 251.400 ;
        RECT 728.400 246.300 730.200 251.400 ;
        RECT 722.400 244.950 730.200 246.300 ;
        RECT 731.400 245.400 733.200 251.400 ;
        RECT 731.400 243.300 732.600 245.400 ;
        RECT 736.950 244.950 739.050 247.050 ;
        RECT 743.400 246.300 745.200 251.400 ;
        RECT 749.400 246.300 751.200 251.400 ;
        RECT 743.400 244.950 751.200 246.300 ;
        RECT 752.400 245.400 754.200 251.400 ;
        RECT 764.400 246.300 766.200 251.400 ;
        RECT 770.400 246.300 772.200 251.400 ;
        RECT 704.400 242.250 708.150 243.300 ;
        RECT 706.950 242.100 708.150 242.250 ;
        RECT 728.850 242.250 732.600 243.300 ;
        RECT 728.850 242.100 730.050 242.250 ;
        RECT 704.100 239.100 705.900 239.850 ;
        RECT 706.950 238.950 709.050 241.050 ;
        RECT 710.100 239.100 711.900 239.850 ;
        RECT 712.950 238.950 715.050 241.050 ;
        RECT 721.950 238.950 724.200 241.050 ;
        RECT 725.100 239.100 726.900 239.850 ;
        RECT 727.950 238.950 730.050 241.050 ;
        RECT 731.100 239.100 732.900 239.850 ;
        RECT 703.950 235.950 706.050 238.050 ;
        RECT 707.850 234.900 708.900 237.900 ;
        RECT 709.950 235.950 712.050 238.050 ;
        RECT 713.100 237.150 714.900 237.900 ;
        RECT 722.100 237.150 723.900 237.900 ;
        RECT 724.950 235.950 727.200 238.050 ;
        RECT 728.100 234.900 729.150 237.900 ;
        RECT 730.950 235.950 733.050 238.050 ;
        RECT 707.850 231.600 709.050 234.900 ;
        RECT 727.950 231.600 729.150 234.900 ;
        RECT 697.950 226.950 700.050 229.050 ;
        RECT 707.700 219.600 709.500 231.600 ;
        RECT 727.500 219.600 729.300 231.600 ;
        RECT 737.550 223.050 738.450 244.950 ;
        RECT 752.400 243.300 753.600 245.400 ;
        RECT 764.400 244.950 772.200 246.300 ;
        RECT 773.400 245.400 775.200 251.400 ;
        RECT 778.950 247.950 781.050 250.050 ;
        RECT 773.400 243.300 774.600 245.400 ;
        RECT 749.850 242.250 753.600 243.300 ;
        RECT 770.850 242.250 774.600 243.300 ;
        RECT 749.850 242.100 751.050 242.250 ;
        RECT 770.850 242.100 772.050 242.250 ;
        RECT 742.800 238.950 745.050 241.050 ;
        RECT 746.100 239.100 747.900 239.850 ;
        RECT 748.950 238.950 751.050 241.050 ;
        RECT 752.100 239.100 753.900 239.850 ;
        RECT 763.950 238.950 766.050 241.050 ;
        RECT 767.100 239.100 768.900 239.850 ;
        RECT 769.950 238.950 772.050 241.050 ;
        RECT 773.100 239.100 774.900 239.850 ;
        RECT 779.550 238.050 780.450 247.950 ;
        RECT 790.200 247.050 792.000 251.400 ;
        RECT 799.950 247.950 802.050 250.050 ;
        RECT 790.200 245.400 795.600 247.050 ;
        RECT 794.700 242.100 795.600 245.400 ;
        RECT 785.100 239.100 786.900 239.850 ;
        RECT 787.950 238.950 790.050 241.050 ;
        RECT 793.950 240.450 796.050 241.050 ;
        RECT 800.550 240.450 801.450 247.950 ;
        RECT 813.000 247.050 814.800 251.400 ;
        RECT 809.400 245.400 814.800 247.050 ;
        RECT 827.400 246.300 829.200 251.400 ;
        RECT 833.400 246.300 835.200 251.400 ;
        RECT 809.400 242.100 810.300 245.400 ;
        RECT 827.400 244.950 835.200 246.300 ;
        RECT 836.400 245.400 838.200 251.400 ;
        RECT 841.950 247.950 844.050 250.050 ;
        RECT 850.950 247.950 853.050 250.050 ;
        RECT 836.400 243.300 837.600 245.400 ;
        RECT 833.850 242.250 837.600 243.300 ;
        RECT 833.850 242.100 835.050 242.250 ;
        RECT 808.950 240.450 811.050 241.050 ;
        RECT 791.100 239.100 792.900 239.850 ;
        RECT 793.950 239.550 801.450 240.450 ;
        RECT 793.950 238.950 796.050 239.550 ;
        RECT 743.100 237.150 744.900 237.900 ;
        RECT 745.950 235.950 748.200 238.050 ;
        RECT 749.100 234.900 750.150 237.900 ;
        RECT 751.950 235.950 754.050 238.050 ;
        RECT 757.950 235.950 760.050 238.050 ;
        RECT 764.100 237.150 765.900 237.900 ;
        RECT 766.950 235.950 769.050 238.050 ;
        RECT 748.950 231.600 750.150 234.900 ;
        RECT 758.550 232.050 759.450 235.950 ;
        RECT 770.100 234.900 771.150 237.900 ;
        RECT 772.950 235.950 775.050 238.050 ;
        RECT 778.950 235.950 781.050 238.050 ;
        RECT 784.950 235.950 787.050 238.050 ;
        RECT 788.100 237.150 789.900 237.900 ;
        RECT 790.950 235.950 793.050 238.050 ;
        RECT 736.950 220.950 739.050 223.050 ;
        RECT 748.500 219.600 750.300 231.600 ;
        RECT 757.950 229.950 760.050 232.050 ;
        RECT 769.950 231.600 771.150 234.900 ;
        RECT 794.700 231.600 795.600 237.900 ;
        RECT 769.500 219.600 771.300 231.600 ;
        RECT 785.400 230.700 793.200 231.600 ;
        RECT 785.400 219.600 787.200 230.700 ;
        RECT 791.400 219.600 793.200 230.700 ;
        RECT 794.400 219.600 796.200 231.600 ;
        RECT 800.550 226.050 801.450 239.550 ;
        RECT 803.550 239.550 811.050 240.450 ;
        RECT 803.550 229.050 804.450 239.550 ;
        RECT 808.950 238.950 811.050 239.550 ;
        RECT 812.100 239.100 813.900 239.850 ;
        RECT 814.950 238.950 817.050 241.050 ;
        RECT 818.100 239.100 819.900 239.850 ;
        RECT 826.950 238.950 829.050 241.050 ;
        RECT 830.100 239.100 831.900 239.850 ;
        RECT 832.950 238.950 835.050 241.050 ;
        RECT 836.100 239.100 837.900 239.850 ;
        RECT 809.400 231.600 810.300 237.900 ;
        RECT 811.950 235.950 814.050 238.050 ;
        RECT 815.100 237.150 816.900 237.900 ;
        RECT 817.950 235.950 820.050 238.050 ;
        RECT 827.100 237.150 828.900 237.900 ;
        RECT 829.800 235.950 832.050 238.050 ;
        RECT 833.100 234.900 834.150 237.900 ;
        RECT 835.950 235.950 838.050 238.050 ;
        RECT 832.950 231.600 834.150 234.900 ;
        RECT 802.950 226.950 805.050 229.050 ;
        RECT 800.100 223.950 802.200 226.050 ;
        RECT 808.800 219.600 810.600 231.600 ;
        RECT 811.800 230.700 819.600 231.600 ;
        RECT 811.800 219.600 813.600 230.700 ;
        RECT 817.800 219.600 819.600 230.700 ;
        RECT 832.500 219.600 834.300 231.600 ;
        RECT 842.550 226.050 843.450 247.950 ;
        RECT 841.950 223.950 844.050 226.050 ;
        RECT 851.550 223.050 852.450 247.950 ;
        RECT 850.950 220.950 853.050 223.050 ;
        RECT 14.700 203.400 16.500 215.400 ;
        RECT 32.400 209.400 34.200 215.400 ;
        RECT 32.700 209.100 34.200 209.400 ;
        RECT 38.400 209.400 40.200 215.400 ;
        RECT 53.400 209.400 55.200 215.400 ;
        RECT 38.400 209.100 39.300 209.400 ;
        RECT 32.700 208.200 39.300 209.100 ;
        RECT 53.700 209.100 55.200 209.400 ;
        RECT 59.400 209.400 61.200 215.400 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 59.400 209.100 60.300 209.400 ;
        RECT 53.700 208.200 60.300 209.100 ;
        RECT 14.850 200.100 16.050 203.400 ;
        RECT 32.100 203.100 33.900 203.850 ;
        RECT 38.400 203.100 39.300 208.200 ;
        RECT 53.100 203.100 54.900 203.850 ;
        RECT 59.400 203.100 60.300 208.200 ;
        RECT 10.950 196.950 13.050 199.050 ;
        RECT 14.850 197.100 15.900 200.100 ;
        RECT 31.950 199.950 34.200 202.050 ;
        RECT 37.950 201.450 40.050 202.050 ;
        RECT 42.000 201.450 46.050 202.050 ;
        RECT 37.950 200.550 46.050 201.450 ;
        RECT 37.950 199.950 40.050 200.550 ;
        RECT 42.000 199.950 46.050 200.550 ;
        RECT 52.950 199.950 55.050 202.050 ;
        RECT 58.950 199.950 64.050 202.050 ;
        RECT 16.950 196.950 19.050 199.050 ;
        RECT 20.100 197.100 21.900 197.850 ;
        RECT 28.950 196.950 31.050 199.050 ;
        RECT 34.950 196.950 37.050 199.050 ;
        RECT 11.100 195.150 12.900 195.900 ;
        RECT 13.800 193.950 16.050 196.050 ;
        RECT 17.100 195.150 18.900 195.900 ;
        RECT 19.950 193.950 22.200 196.050 ;
        RECT 29.100 195.150 30.900 195.900 ;
        RECT 35.100 195.150 36.900 195.900 ;
        RECT 38.400 193.650 39.300 198.900 ;
        RECT 49.800 196.950 52.050 199.050 ;
        RECT 55.950 196.950 58.050 199.050 ;
        RECT 50.100 195.150 51.900 195.900 ;
        RECT 56.100 195.150 57.900 195.900 ;
        RECT 59.400 193.650 60.300 198.900 ;
        RECT 68.550 195.450 69.450 211.950 ;
        RECT 73.800 203.400 75.600 215.400 ;
        RECT 76.800 204.300 78.600 215.400 ;
        RECT 82.800 204.300 84.600 215.400 ;
        RECT 76.800 203.400 84.600 204.300 ;
        RECT 98.700 203.400 100.500 215.400 ;
        RECT 119.700 203.400 121.500 215.400 ;
        RECT 137.400 209.400 139.200 215.400 ;
        RECT 137.700 209.100 139.200 209.400 ;
        RECT 143.400 209.400 145.200 215.400 ;
        RECT 143.400 209.100 144.300 209.400 ;
        RECT 137.700 208.200 144.300 209.100 ;
        RECT 74.400 197.100 75.300 203.400 ;
        RECT 98.850 200.100 100.050 203.400 ;
        RECT 119.850 200.100 121.050 203.400 ;
        RECT 137.100 203.100 138.900 203.850 ;
        RECT 143.400 203.100 144.300 208.200 ;
        RECT 157.200 203.400 159.000 215.400 ;
        RECT 163.800 209.400 165.600 215.400 ;
        RECT 76.800 196.950 79.050 199.050 ;
        RECT 80.100 197.100 81.900 197.850 ;
        RECT 82.950 196.950 85.050 199.050 ;
        RECT 94.950 196.950 97.050 199.050 ;
        RECT 98.850 197.100 99.900 200.100 ;
        RECT 100.950 196.950 103.050 199.050 ;
        RECT 104.100 197.100 105.900 197.850 ;
        RECT 115.950 196.950 118.050 199.050 ;
        RECT 119.850 197.100 120.900 200.100 ;
        RECT 136.950 199.950 139.050 202.050 ;
        RECT 142.950 199.950 148.050 202.050 ;
        RECT 121.950 196.950 124.200 199.050 ;
        RECT 125.100 197.100 126.900 197.850 ;
        RECT 133.950 196.950 136.050 199.050 ;
        RECT 139.950 196.950 142.050 199.050 ;
        RECT 73.950 195.450 76.050 196.050 ;
        RECT 68.550 194.550 76.050 195.450 ;
        RECT 77.100 195.150 78.900 195.900 ;
        RECT 73.950 193.950 76.050 194.550 ;
        RECT 79.950 193.950 82.050 196.050 ;
        RECT 83.100 195.150 84.900 195.900 ;
        RECT 95.100 195.150 96.900 195.900 ;
        RECT 97.800 193.950 100.050 196.050 ;
        RECT 101.100 195.150 102.900 195.900 ;
        RECT 103.950 193.950 106.200 196.050 ;
        RECT 116.100 195.150 117.900 195.900 ;
        RECT 118.950 193.950 121.050 196.050 ;
        RECT 122.100 195.150 123.900 195.900 ;
        RECT 124.950 193.950 127.050 196.050 ;
        RECT 134.100 195.150 135.900 195.900 ;
        RECT 140.100 195.150 141.900 195.900 ;
        RECT 143.400 193.650 144.300 198.900 ;
        RECT 157.950 197.100 159.000 203.400 ;
        RECT 160.950 196.950 163.050 199.050 ;
        RECT 154.950 193.950 160.050 196.050 ;
        RECT 161.100 195.150 162.900 195.900 ;
        RECT 13.950 192.750 15.150 192.900 ;
        RECT 11.400 191.700 15.150 192.750 ;
        RECT 35.100 192.000 39.300 193.650 ;
        RECT 56.100 192.000 60.300 193.650 ;
        RECT 11.400 189.600 12.600 191.700 ;
        RECT 10.800 183.600 12.600 189.600 ;
        RECT 13.800 188.700 21.600 190.050 ;
        RECT 13.800 183.600 15.600 188.700 ;
        RECT 19.800 183.600 21.600 188.700 ;
        RECT 35.100 183.600 36.900 192.000 ;
        RECT 56.100 183.600 57.900 192.000 ;
        RECT 74.400 189.600 75.300 192.900 ;
        RECT 97.950 192.750 99.150 192.900 ;
        RECT 118.950 192.750 120.150 192.900 ;
        RECT 95.400 191.700 99.150 192.750 ;
        RECT 116.400 191.700 120.150 192.750 ;
        RECT 140.100 192.000 144.300 193.650 ;
        RECT 95.400 189.600 96.600 191.700 ;
        RECT 74.400 187.950 79.800 189.600 ;
        RECT 78.000 183.600 79.800 187.950 ;
        RECT 94.800 183.600 96.600 189.600 ;
        RECT 97.800 188.700 105.600 190.050 ;
        RECT 116.400 189.600 117.600 191.700 ;
        RECT 97.800 183.600 99.600 188.700 ;
        RECT 103.800 183.600 105.600 188.700 ;
        RECT 115.800 183.600 117.600 189.600 ;
        RECT 118.800 188.700 126.600 190.050 ;
        RECT 118.800 183.600 120.600 188.700 ;
        RECT 124.800 183.600 126.600 188.700 ;
        RECT 140.100 183.600 141.900 192.000 ;
        RECT 159.150 189.600 160.050 192.900 ;
        RECT 164.550 192.300 165.600 209.400 ;
        RECT 179.400 209.400 181.200 215.400 ;
        RECT 188.100 211.950 190.200 214.050 ;
        RECT 175.950 199.950 178.050 202.050 ;
        RECT 179.400 200.100 180.600 209.400 ;
        RECT 181.950 199.950 184.050 202.050 ;
        RECT 176.100 198.150 177.900 198.900 ;
        RECT 167.100 197.100 168.900 197.850 ;
        RECT 178.950 196.950 181.200 199.050 ;
        RECT 182.100 198.150 183.900 198.900 ;
        RECT 166.950 193.950 169.050 196.050 ;
        RECT 161.100 191.100 168.600 192.300 ;
        RECT 161.100 190.500 162.900 191.100 ;
        RECT 159.150 187.800 161.100 189.600 ;
        RECT 159.300 183.600 161.100 187.800 ;
        RECT 166.800 183.600 168.600 191.100 ;
        RECT 179.400 191.700 180.600 195.900 ;
        RECT 179.400 190.800 183.000 191.700 ;
        RECT 181.200 183.600 183.000 190.800 ;
        RECT 188.550 190.050 189.450 211.950 ;
        RECT 199.800 209.400 201.600 215.400 ;
        RECT 196.950 199.950 199.050 202.050 ;
        RECT 200.400 200.100 201.600 209.400 ;
        RECT 215.400 209.400 217.200 215.400 ;
        RECT 235.800 209.400 237.600 215.400 ;
        RECT 202.950 199.950 205.050 202.050 ;
        RECT 208.950 199.950 214.050 202.050 ;
        RECT 215.400 200.100 216.600 209.400 ;
        RECT 217.950 199.950 220.050 205.050 ;
        RECT 232.950 199.950 235.050 202.050 ;
        RECT 236.400 200.100 237.600 209.400 ;
        RECT 248.400 205.500 250.200 215.400 ;
        RECT 254.400 214.500 262.200 215.400 ;
        RECT 254.400 205.500 256.200 214.500 ;
        RECT 248.400 204.600 256.200 205.500 ;
        RECT 257.400 205.800 259.200 213.600 ;
        RECT 260.400 206.700 262.200 214.500 ;
        RECT 264.000 214.500 271.800 215.400 ;
        RECT 264.000 205.800 265.800 214.500 ;
        RECT 257.400 204.900 265.800 205.800 ;
        RECT 267.000 205.800 268.800 213.600 ;
        RECT 267.000 203.400 268.200 205.800 ;
        RECT 270.000 205.200 271.800 214.500 ;
        RECT 284.400 209.400 286.200 215.400 ;
        RECT 264.750 202.200 268.200 203.400 ;
        RECT 238.950 199.950 241.050 202.050 ;
        RECT 264.750 199.950 265.950 202.200 ;
        RECT 284.400 200.100 285.600 209.400 ;
        RECT 301.500 203.400 303.300 215.400 ;
        RECT 319.800 209.400 321.600 215.400 ;
        RECT 304.950 205.950 307.050 208.050 ;
        RECT 301.950 200.100 303.150 203.400 ;
        RECT 197.100 198.150 198.900 198.900 ;
        RECT 199.950 196.950 202.050 199.050 ;
        RECT 203.100 198.150 204.900 198.900 ;
        RECT 212.100 198.150 213.900 198.900 ;
        RECT 214.950 196.950 217.050 199.050 ;
        RECT 218.100 198.150 219.900 198.900 ;
        RECT 233.100 198.150 234.900 198.900 ;
        RECT 235.950 196.950 238.050 199.050 ;
        RECT 239.100 198.150 240.900 198.900 ;
        RECT 251.100 196.950 252.900 197.700 ;
        RECT 256.950 196.800 259.050 199.050 ;
        RECT 260.100 196.950 261.900 197.700 ;
        RECT 200.400 191.700 201.600 195.900 ;
        RECT 198.000 190.800 201.600 191.700 ;
        RECT 215.400 191.700 216.600 195.900 ;
        RECT 236.400 191.700 237.600 195.900 ;
        RECT 250.950 193.800 253.050 195.900 ;
        RECT 257.100 195.000 258.900 195.750 ;
        RECT 259.950 193.050 262.050 195.900 ;
        RECT 215.400 190.800 219.000 191.700 ;
        RECT 187.950 187.950 190.050 190.050 ;
        RECT 198.000 183.600 199.800 190.800 ;
        RECT 217.200 183.600 219.000 190.800 ;
        RECT 234.000 190.800 237.600 191.700 ;
        RECT 259.800 191.550 262.050 193.050 ;
        RECT 264.750 195.750 264.900 199.950 ;
        RECT 265.950 198.450 268.050 198.900 ;
        RECT 265.950 197.550 273.450 198.450 ;
        RECT 265.950 196.800 268.050 197.550 ;
        RECT 259.800 190.950 261.900 191.550 ;
        RECT 234.000 183.600 235.800 190.800 ;
        RECT 264.750 188.400 265.950 195.750 ;
        RECT 255.150 187.500 265.950 188.400 ;
        RECT 255.150 186.600 256.200 187.500 ;
        RECT 261.150 186.600 262.200 187.500 ;
        RECT 272.550 187.050 273.450 197.550 ;
        RECT 283.950 196.950 289.050 199.050 ;
        RECT 296.100 197.100 297.900 197.850 ;
        RECT 298.800 196.950 301.050 199.050 ;
        RECT 302.100 197.100 303.150 200.100 ;
        RECT 305.550 199.050 306.450 205.950 ;
        RECT 320.400 200.100 321.600 209.400 ;
        RECT 332.400 204.300 334.200 215.400 ;
        RECT 338.400 204.300 340.200 215.400 ;
        RECT 332.400 203.400 340.200 204.300 ;
        RECT 341.400 203.400 343.200 215.400 ;
        RECT 358.800 209.400 360.600 215.400 ;
        RECT 367.950 211.950 370.050 214.050 ;
        RECT 304.950 196.950 307.050 199.050 ;
        RECT 319.950 196.950 325.050 199.050 ;
        RECT 331.950 196.950 334.050 199.050 ;
        RECT 335.100 197.100 336.900 197.850 ;
        RECT 337.950 196.950 340.050 202.050 ;
        RECT 341.700 197.100 342.600 203.400 ;
        RECT 349.950 201.450 352.050 205.050 ;
        RECT 355.950 201.450 358.050 202.050 ;
        RECT 349.950 201.000 358.050 201.450 ;
        RECT 350.550 200.550 358.050 201.000 ;
        RECT 355.950 199.950 358.050 200.550 ;
        RECT 359.400 200.100 360.600 209.400 ;
        RECT 361.800 199.950 364.050 202.050 ;
        RECT 368.550 199.050 369.450 211.950 ;
        RECT 376.800 209.400 378.600 215.400 ;
        RECT 373.950 199.950 376.050 202.050 ;
        RECT 377.400 200.100 378.600 209.400 ;
        RECT 393.600 203.400 395.400 215.400 ;
        RECT 411.900 203.400 415.200 215.400 ;
        RECT 433.800 203.400 435.600 215.400 ;
        RECT 450.600 203.400 452.400 215.400 ;
        RECT 466.800 214.500 474.600 215.400 ;
        RECT 466.800 203.400 468.600 214.500 ;
        RECT 393.600 202.350 396.300 203.400 ;
        RECT 379.950 199.950 382.050 202.050 ;
        RECT 356.100 198.150 357.900 198.900 ;
        RECT 358.950 196.950 361.050 199.050 ;
        RECT 362.100 198.150 363.900 198.900 ;
        RECT 367.950 196.950 370.050 199.050 ;
        RECT 374.100 198.150 375.900 198.900 ;
        RECT 376.950 196.950 379.050 199.050 ;
        RECT 380.100 198.150 381.900 198.900 ;
        RECT 392.100 197.100 393.900 197.850 ;
        RECT 394.950 197.100 396.300 202.350 ;
        RECT 398.100 197.100 399.900 197.850 ;
        RECT 281.100 194.100 282.900 194.850 ;
        RECT 280.950 190.950 283.050 193.050 ;
        RECT 254.400 183.600 256.200 186.600 ;
        RECT 260.400 183.600 262.200 186.600 ;
        RECT 272.100 184.950 274.200 187.050 ;
        RECT 284.400 186.600 285.600 195.900 ;
        RECT 295.950 193.950 298.050 196.050 ;
        RECT 299.100 195.150 300.900 195.900 ;
        RECT 301.950 193.950 304.050 196.050 ;
        RECT 305.100 195.150 306.900 195.900 ;
        RECT 302.850 192.750 304.050 192.900 ;
        RECT 302.850 191.700 306.600 192.750 ;
        RECT 296.400 188.700 304.200 190.050 ;
        RECT 284.400 183.600 286.200 186.600 ;
        RECT 296.400 183.600 298.200 188.700 ;
        RECT 302.400 183.600 304.200 188.700 ;
        RECT 305.400 189.600 306.600 191.700 ;
        RECT 305.400 183.600 307.200 189.600 ;
        RECT 320.400 186.600 321.600 195.900 ;
        RECT 332.100 195.150 333.900 195.900 ;
        RECT 323.100 194.100 324.900 194.850 ;
        RECT 334.950 193.950 337.050 196.050 ;
        RECT 338.100 195.150 339.900 195.900 ;
        RECT 340.950 193.950 346.050 196.050 ;
        RECT 322.950 190.950 325.050 193.050 ;
        RECT 341.700 189.600 342.600 192.900 ;
        RECT 359.400 191.700 360.600 195.900 ;
        RECT 377.400 191.700 378.600 195.900 ;
        RECT 391.950 193.950 394.050 196.050 ;
        RECT 395.100 194.100 396.300 197.100 ;
        RECT 409.800 196.950 412.050 199.050 ;
        RECT 413.400 197.100 414.600 203.400 ;
        RECT 415.950 196.950 418.200 199.050 ;
        RECT 434.400 197.100 435.600 203.400 ;
        RECT 449.700 202.350 452.400 203.400 ;
        RECT 469.800 202.500 471.600 213.600 ;
        RECT 472.800 204.600 474.600 214.500 ;
        RECT 478.800 204.600 480.600 215.400 ;
        RECT 490.800 209.400 492.600 215.400 ;
        RECT 472.800 203.700 480.600 204.600 ;
        RECT 436.950 196.950 439.050 199.050 ;
        RECT 446.100 197.100 447.900 197.850 ;
        RECT 449.700 197.100 451.050 202.350 ;
        RECT 469.800 201.600 473.850 202.500 ;
        RECT 472.950 200.100 473.850 201.600 ;
        RECT 491.400 200.100 492.600 209.400 ;
        RECT 497.550 203.400 499.350 215.400 ;
        RECT 505.050 209.400 506.850 215.400 ;
        RECT 502.950 207.300 506.850 209.400 ;
        RECT 512.850 208.500 514.650 215.400 ;
        RECT 520.650 209.400 522.450 215.400 ;
        RECT 521.250 208.500 522.450 209.400 ;
        RECT 511.950 207.450 518.550 208.500 ;
        RECT 511.950 206.700 513.750 207.450 ;
        RECT 516.750 206.700 518.550 207.450 ;
        RECT 521.250 206.400 526.050 208.500 ;
        RECT 504.150 204.600 506.850 206.400 ;
        RECT 507.750 205.800 509.550 206.400 ;
        RECT 507.750 204.900 514.050 205.800 ;
        RECT 521.250 205.500 522.450 206.400 ;
        RECT 507.750 204.600 509.550 204.900 ;
        RECT 505.950 203.700 506.850 204.600 ;
        RECT 452.100 197.100 453.900 197.850 ;
        RECT 467.100 197.100 468.900 197.850 ;
        RECT 397.950 193.950 400.050 196.050 ;
        RECT 406.950 193.950 409.050 196.050 ;
        RECT 410.100 195.150 411.900 195.900 ;
        RECT 412.800 193.950 415.050 196.050 ;
        RECT 416.100 195.150 417.750 195.900 ;
        RECT 418.950 193.950 421.050 196.050 ;
        RECT 433.950 193.950 436.050 196.050 ;
        RECT 437.100 195.150 438.900 195.900 ;
        RECT 445.950 193.950 448.050 196.050 ;
        RECT 449.700 194.100 450.900 197.100 ;
        RECT 469.800 196.950 472.050 199.050 ;
        RECT 473.100 197.100 473.850 200.100 ;
        RECT 475.950 196.950 478.200 199.050 ;
        RECT 479.100 197.100 480.750 197.850 ;
        RECT 487.950 196.950 493.050 199.050 ;
        RECT 497.550 196.050 498.750 203.400 ;
        RECT 502.950 202.800 505.050 203.700 ;
        RECT 505.950 202.800 511.950 203.700 ;
        RECT 500.850 201.600 505.050 202.800 ;
        RECT 499.950 199.800 501.750 201.600 ;
        RECT 511.050 197.100 511.950 202.800 ;
        RECT 513.150 202.800 514.050 204.900 ;
        RECT 514.950 204.300 522.450 205.500 ;
        RECT 514.950 203.700 516.750 204.300 ;
        RECT 529.050 203.400 530.850 215.400 ;
        RECT 541.800 209.400 543.600 215.400 ;
        RECT 519.750 202.800 530.850 203.400 ;
        RECT 513.150 202.200 530.850 202.800 ;
        RECT 513.150 201.900 521.550 202.200 ;
        RECT 519.750 201.600 521.550 201.900 ;
        RECT 524.100 196.800 525.900 197.100 ;
        RECT 451.950 193.950 454.050 196.050 ;
        RECT 466.950 193.950 469.050 196.050 ;
        RECT 470.250 195.150 471.900 195.900 ;
        RECT 472.800 193.950 475.050 196.050 ;
        RECT 476.100 195.150 477.750 195.900 ;
        RECT 478.950 193.950 481.050 196.050 ;
        RECT 319.800 183.600 321.600 186.600 ;
        RECT 337.200 187.950 342.600 189.600 ;
        RECT 357.000 190.800 360.600 191.700 ;
        RECT 375.000 190.800 378.600 191.700 ;
        RECT 394.950 190.950 397.050 193.050 ;
        RECT 407.250 192.150 409.050 192.900 ;
        RECT 413.400 192.300 414.600 192.900 ;
        RECT 413.400 191.100 417.600 192.300 ;
        RECT 418.500 192.150 420.300 192.900 ;
        RECT 337.200 183.600 339.000 187.950 ;
        RECT 357.000 183.600 358.800 190.800 ;
        RECT 375.000 183.600 376.800 190.800 ;
        RECT 395.400 186.600 396.600 189.900 ;
        RECT 394.800 183.600 396.600 186.600 ;
        RECT 407.400 189.000 415.200 189.900 ;
        RECT 416.700 189.600 417.600 191.100 ;
        RECT 434.400 189.600 435.600 192.900 ;
        RECT 448.950 190.950 451.050 193.050 ;
        RECT 407.400 183.600 409.200 189.000 ;
        RECT 413.400 184.500 415.200 189.000 ;
        RECT 416.400 185.400 418.200 189.600 ;
        RECT 419.400 184.500 421.200 189.600 ;
        RECT 413.400 183.600 421.200 184.500 ;
        RECT 433.800 183.600 435.600 189.600 ;
        RECT 449.400 186.600 450.600 189.900 ;
        RECT 474.000 189.600 475.050 192.900 ;
        RECT 449.400 183.600 451.200 186.600 ;
        RECT 474.000 183.600 475.800 189.600 ;
        RECT 491.400 186.600 492.600 195.900 ;
        RECT 494.100 194.100 495.900 194.850 ;
        RECT 497.550 193.950 498.900 196.050 ;
        RECT 499.950 193.950 502.050 196.050 ;
        RECT 503.100 193.950 503.850 195.750 ;
        RECT 511.950 193.950 514.050 196.050 ;
        RECT 517.950 193.950 520.200 196.050 ;
        RECT 521.100 195.900 525.900 196.800 ;
        RECT 524.100 195.300 525.900 195.900 ;
        RECT 527.100 195.150 528.900 196.950 ;
        RECT 521.100 194.400 522.900 195.000 ;
        RECT 527.100 194.400 528.000 195.150 ;
        RECT 493.950 190.950 496.050 193.050 ;
        RECT 490.800 183.600 492.600 186.600 ;
        RECT 497.550 189.600 498.750 193.950 ;
        RECT 521.100 193.200 528.000 194.400 ;
        RECT 511.050 192.000 511.950 192.900 ;
        RECT 521.100 192.000 522.150 193.200 ;
        RECT 511.050 191.100 522.150 192.000 ;
        RECT 511.050 190.800 511.950 191.100 ;
        RECT 497.550 183.600 499.350 189.600 ;
        RECT 502.950 188.700 505.050 189.600 ;
        RECT 510.150 189.000 511.950 190.800 ;
        RECT 521.100 190.200 522.150 191.100 ;
        RECT 517.350 189.450 519.150 190.200 ;
        RECT 502.950 187.500 506.700 188.700 ;
        RECT 505.650 186.600 506.700 187.500 ;
        RECT 514.200 188.400 519.150 189.450 ;
        RECT 520.650 188.400 522.450 190.200 ;
        RECT 529.950 189.600 530.850 202.200 ;
        RECT 542.400 200.100 543.600 209.400 ;
        RECT 556.800 203.400 558.600 215.400 ;
        RECT 559.800 204.300 561.600 215.400 ;
        RECT 565.800 204.300 567.600 215.400 ;
        RECT 559.800 203.400 567.600 204.300 ;
        RECT 581.700 203.400 583.500 215.400 ;
        RECT 600.600 203.400 602.400 215.400 ;
        RECT 616.200 203.400 618.000 215.400 ;
        RECT 622.800 209.400 624.600 215.400 ;
        RECT 637.800 209.400 639.600 215.400 ;
        RECT 541.950 196.950 547.050 199.050 ;
        RECT 557.400 197.100 558.300 203.400 ;
        RECT 581.850 200.100 583.050 203.400 ;
        RECT 600.600 202.350 603.300 203.400 ;
        RECT 559.950 196.950 562.050 199.050 ;
        RECT 563.100 197.100 564.900 197.850 ;
        RECT 565.950 196.950 568.050 199.050 ;
        RECT 572.100 196.950 574.200 199.050 ;
        RECT 577.950 196.950 580.050 199.050 ;
        RECT 581.850 197.100 582.900 200.100 ;
        RECT 583.950 196.950 586.050 199.050 ;
        RECT 587.100 197.100 588.900 197.850 ;
        RECT 599.100 197.100 600.900 197.850 ;
        RECT 601.950 197.100 603.300 202.350 ;
        RECT 605.100 197.100 606.900 197.850 ;
        RECT 616.950 197.100 618.000 203.400 ;
        RECT 514.200 186.600 515.250 188.400 ;
        RECT 523.950 187.500 526.050 189.600 ;
        RECT 523.950 186.600 525.000 187.500 ;
        RECT 505.650 183.600 507.450 186.600 ;
        RECT 513.450 183.600 515.250 186.600 ;
        RECT 521.250 185.700 525.000 186.600 ;
        RECT 521.250 183.600 523.050 185.700 ;
        RECT 529.050 183.600 530.850 189.600 ;
        RECT 542.400 186.600 543.600 195.900 ;
        RECT 545.100 194.100 546.900 194.850 ;
        RECT 556.950 193.950 559.050 196.050 ;
        RECT 560.100 195.150 561.900 195.900 ;
        RECT 562.950 193.950 565.050 196.050 ;
        RECT 566.100 195.150 567.900 195.900 ;
        RECT 572.550 193.050 573.450 196.950 ;
        RECT 578.100 195.150 579.900 195.900 ;
        RECT 580.950 193.950 583.050 196.050 ;
        RECT 584.100 195.150 585.900 195.900 ;
        RECT 586.950 193.950 589.050 196.050 ;
        RECT 598.950 193.950 601.050 196.050 ;
        RECT 602.100 194.100 603.300 197.100 ;
        RECT 619.950 196.950 622.050 199.050 ;
        RECT 604.950 193.950 607.050 196.050 ;
        RECT 616.950 195.450 619.050 196.050 ;
        RECT 611.550 194.550 619.050 195.450 ;
        RECT 620.100 195.150 621.900 195.900 ;
        RECT 557.400 189.600 558.300 192.900 ;
        RECT 571.950 190.950 574.050 193.050 ;
        RECT 580.950 192.750 582.150 192.900 ;
        RECT 578.400 191.700 582.150 192.750 ;
        RECT 578.400 189.600 579.600 191.700 ;
        RECT 601.950 190.950 604.050 193.050 ;
        RECT 557.400 187.950 562.800 189.600 ;
        RECT 541.800 183.600 543.600 186.600 ;
        RECT 561.000 183.600 562.800 187.950 ;
        RECT 577.800 183.600 579.600 189.600 ;
        RECT 580.800 188.700 588.600 190.050 ;
        RECT 580.800 183.600 582.600 188.700 ;
        RECT 586.800 183.600 588.600 188.700 ;
        RECT 602.400 186.600 603.600 189.900 ;
        RECT 611.550 187.050 612.450 194.550 ;
        RECT 616.950 193.950 619.050 194.550 ;
        RECT 618.150 189.600 619.050 192.900 ;
        RECT 623.550 192.300 624.600 209.400 ;
        RECT 638.700 209.100 639.600 209.400 ;
        RECT 643.800 209.400 645.600 215.400 ;
        RECT 659.400 209.400 661.200 215.400 ;
        RECT 643.800 209.100 645.300 209.400 ;
        RECT 638.700 208.200 645.300 209.100 ;
        RECT 638.700 203.100 639.600 208.200 ;
        RECT 644.100 203.100 645.900 203.850 ;
        RECT 631.950 201.450 636.000 202.050 ;
        RECT 637.950 201.450 640.050 202.050 ;
        RECT 631.950 200.550 640.050 201.450 ;
        RECT 631.950 199.950 636.000 200.550 ;
        RECT 637.950 199.950 640.050 200.550 ;
        RECT 643.950 199.950 646.050 202.050 ;
        RECT 655.950 199.950 658.050 202.050 ;
        RECT 659.400 200.100 660.600 209.400 ;
        RECT 678.600 203.400 680.400 215.400 ;
        RECT 682.950 208.950 685.050 211.050 ;
        RECT 677.700 202.350 680.400 203.400 ;
        RECT 661.950 199.950 664.050 202.050 ;
        RECT 626.100 197.100 627.900 197.850 ;
        RECT 625.950 193.950 628.050 196.050 ;
        RECT 638.700 193.650 639.600 198.900 ;
        RECT 640.950 196.950 643.050 199.050 ;
        RECT 646.950 196.950 649.050 199.050 ;
        RECT 656.100 198.150 657.900 198.900 ;
        RECT 658.950 196.950 661.050 199.050 ;
        RECT 662.100 198.150 663.900 198.900 ;
        RECT 674.100 197.100 675.900 197.850 ;
        RECT 677.700 197.100 679.050 202.350 ;
        RECT 683.550 202.050 684.450 208.950 ;
        RECT 697.500 203.400 699.300 215.400 ;
        RECT 718.500 203.400 720.300 215.400 ;
        RECT 731.100 213.450 733.200 214.050 ;
        RECT 725.550 213.000 733.200 213.450 ;
        RECT 724.950 212.550 733.200 213.000 ;
        RECT 724.950 208.950 727.050 212.550 ;
        RECT 731.100 211.950 733.200 212.550 ;
        RECT 737.400 209.400 739.200 215.400 ;
        RECT 682.950 199.950 685.050 202.050 ;
        RECT 697.950 200.100 699.150 203.400 ;
        RECT 718.950 200.100 720.150 203.400 ;
        RECT 737.400 200.100 738.600 209.400 ;
        RECT 745.950 205.950 748.050 208.050 ;
        RECT 742.950 202.950 745.050 205.050 ;
        RECT 680.100 197.100 681.900 197.850 ;
        RECT 692.100 197.100 693.900 197.850 ;
        RECT 641.100 195.150 642.900 195.900 ;
        RECT 647.100 195.150 648.900 195.900 ;
        RECT 620.100 191.100 627.600 192.300 ;
        RECT 638.700 192.000 642.900 193.650 ;
        RECT 620.100 190.500 621.900 191.100 ;
        RECT 618.150 187.800 620.100 189.600 ;
        RECT 601.800 183.600 603.600 186.600 ;
        RECT 610.950 184.950 613.050 187.050 ;
        RECT 618.300 183.600 620.100 187.800 ;
        RECT 625.800 183.600 627.600 191.100 ;
        RECT 641.100 183.600 642.900 192.000 ;
        RECT 659.400 191.700 660.600 195.900 ;
        RECT 673.950 193.950 676.050 196.050 ;
        RECT 677.700 194.100 678.900 197.100 ;
        RECT 694.950 196.950 697.050 199.050 ;
        RECT 698.100 197.100 699.150 200.100 ;
        RECT 700.950 196.950 703.050 199.050 ;
        RECT 713.100 197.100 714.900 197.850 ;
        RECT 715.950 196.950 718.050 199.050 ;
        RECT 719.100 197.100 720.150 200.100 ;
        RECT 721.950 196.950 724.200 199.050 ;
        RECT 736.950 196.950 742.050 199.050 ;
        RECT 679.950 193.950 682.050 196.050 ;
        RECT 691.800 193.950 694.050 196.050 ;
        RECT 695.100 195.150 696.900 195.900 ;
        RECT 697.950 193.950 700.050 196.050 ;
        RECT 701.100 195.150 702.900 195.900 ;
        RECT 712.950 193.950 715.050 196.050 ;
        RECT 716.100 195.150 717.900 195.900 ;
        RECT 718.950 193.950 721.050 196.050 ;
        RECT 722.100 195.150 723.900 195.900 ;
        RECT 734.100 194.100 735.900 194.850 ;
        RECT 659.400 190.800 663.000 191.700 ;
        RECT 676.950 190.950 679.050 193.050 ;
        RECT 698.850 192.750 700.050 192.900 ;
        RECT 719.850 192.750 721.050 192.900 ;
        RECT 698.850 191.700 702.600 192.750 ;
        RECT 719.850 191.700 723.600 192.750 ;
        RECT 661.200 183.600 663.000 190.800 ;
        RECT 677.400 186.600 678.600 189.900 ;
        RECT 692.400 188.700 700.200 190.050 ;
        RECT 677.400 183.600 679.200 186.600 ;
        RECT 692.400 183.600 694.200 188.700 ;
        RECT 698.400 183.600 700.200 188.700 ;
        RECT 701.400 189.600 702.600 191.700 ;
        RECT 701.400 183.600 703.200 189.600 ;
        RECT 713.400 188.700 721.200 190.050 ;
        RECT 713.400 183.600 715.200 188.700 ;
        RECT 719.400 183.600 721.200 188.700 ;
        RECT 722.400 189.600 723.600 191.700 ;
        RECT 733.950 190.950 736.050 193.050 ;
        RECT 722.400 183.600 724.200 189.600 ;
        RECT 737.400 186.600 738.600 195.900 ;
        RECT 743.550 187.050 744.450 202.950 ;
        RECT 746.550 202.050 747.450 205.950 ;
        RECT 753.900 203.400 757.200 215.400 ;
        RECT 763.950 205.950 766.050 208.050 ;
        RECT 745.950 199.950 748.050 202.050 ;
        RECT 751.950 196.950 754.050 199.050 ;
        RECT 755.400 197.100 756.600 203.400 ;
        RECT 764.550 202.050 765.450 205.950 ;
        RECT 777.600 203.400 779.400 215.400 ;
        RECT 796.800 209.400 798.600 215.400 ;
        RECT 777.600 202.350 780.300 203.400 ;
        RECT 763.950 199.950 766.050 202.050 ;
        RECT 757.950 196.950 760.050 199.050 ;
        RECT 776.100 197.100 777.900 197.850 ;
        RECT 778.950 197.100 780.300 202.350 ;
        RECT 793.950 199.950 796.050 202.050 ;
        RECT 797.400 200.100 798.600 209.400 ;
        RECT 811.800 203.400 813.600 215.400 ;
        RECT 814.800 204.300 816.600 215.400 ;
        RECT 820.800 204.300 822.600 215.400 ;
        RECT 814.800 203.400 822.600 204.300 ;
        RECT 833.400 209.400 835.200 215.400 ;
        RECT 850.800 209.400 852.600 215.400 ;
        RECT 799.950 199.950 802.050 202.050 ;
        RECT 794.100 198.150 795.900 198.900 ;
        RECT 782.100 197.100 783.900 197.850 ;
        RECT 748.950 193.950 751.050 196.050 ;
        RECT 752.100 195.150 753.900 195.900 ;
        RECT 754.950 193.950 757.050 196.050 ;
        RECT 758.100 195.150 759.750 195.900 ;
        RECT 760.950 193.950 763.050 196.050 ;
        RECT 775.800 193.950 778.050 196.050 ;
        RECT 779.100 194.100 780.300 197.100 ;
        RECT 796.950 196.950 799.050 199.050 ;
        RECT 800.100 198.150 801.900 198.900 ;
        RECT 812.400 197.100 813.300 203.400 ;
        RECT 829.950 199.950 832.050 202.050 ;
        RECT 833.400 200.100 834.600 209.400 ;
        RECT 835.950 199.950 838.050 202.050 ;
        RECT 851.400 200.100 852.600 209.400 ;
        RECT 814.800 196.950 817.050 199.050 ;
        RECT 818.100 197.100 819.900 197.850 ;
        RECT 820.950 196.950 823.050 199.050 ;
        RECT 830.100 198.150 831.900 198.900 ;
        RECT 832.950 196.950 835.050 199.050 ;
        RECT 836.100 198.150 837.900 198.900 ;
        RECT 847.950 196.950 853.050 199.050 ;
        RECT 781.950 193.950 784.050 196.050 ;
        RECT 749.250 192.150 751.050 192.900 ;
        RECT 755.400 192.300 756.600 192.900 ;
        RECT 755.400 191.100 759.600 192.300 ;
        RECT 760.500 192.150 762.300 192.900 ;
        RECT 749.400 189.000 757.200 189.900 ;
        RECT 758.700 189.600 759.600 191.100 ;
        RECT 778.950 190.950 781.050 193.050 ;
        RECT 797.400 191.700 798.600 195.900 ;
        RECT 808.800 193.950 814.050 196.050 ;
        RECT 815.100 195.150 816.900 195.900 ;
        RECT 817.950 193.950 820.050 196.050 ;
        RECT 821.100 195.150 822.900 195.900 ;
        RECT 795.000 190.800 798.600 191.700 ;
        RECT 737.400 183.600 739.200 186.600 ;
        RECT 742.950 184.950 745.050 187.050 ;
        RECT 749.400 183.600 751.200 189.000 ;
        RECT 755.400 184.500 757.200 189.000 ;
        RECT 758.400 185.400 760.200 189.600 ;
        RECT 761.400 184.500 763.200 189.600 ;
        RECT 779.400 186.600 780.600 189.900 ;
        RECT 755.400 183.600 763.200 184.500 ;
        RECT 778.800 183.600 780.600 186.600 ;
        RECT 795.000 183.600 796.800 190.800 ;
        RECT 812.400 189.600 813.300 192.900 ;
        RECT 833.400 191.700 834.600 195.900 ;
        RECT 833.400 190.800 837.000 191.700 ;
        RECT 812.400 187.950 817.800 189.600 ;
        RECT 816.000 183.600 817.800 187.950 ;
        RECT 835.200 183.600 837.000 190.800 ;
        RECT 851.400 186.600 852.600 195.900 ;
        RECT 854.100 194.100 855.900 194.850 ;
        RECT 853.950 190.950 856.050 193.050 ;
        RECT 850.800 183.600 852.600 186.600 ;
        RECT 10.800 173.400 12.600 179.400 ;
        RECT 11.400 171.300 12.600 173.400 ;
        RECT 13.800 174.300 15.600 179.400 ;
        RECT 19.800 174.300 21.600 179.400 ;
        RECT 25.950 175.950 28.050 178.050 ;
        RECT 13.800 172.950 21.600 174.300 ;
        RECT 11.400 170.250 15.150 171.300 ;
        RECT 13.950 170.100 15.150 170.250 ;
        RECT 26.550 169.050 27.450 175.950 ;
        RECT 35.100 171.000 36.900 179.400 ;
        RECT 55.200 175.050 57.000 179.400 ;
        RECT 76.200 175.050 78.000 179.400 ;
        RECT 55.200 173.400 60.600 175.050 ;
        RECT 76.200 173.400 81.600 175.050 ;
        RECT 32.700 169.350 36.900 171.000 ;
        RECT 59.700 170.100 60.600 173.400 ;
        RECT 80.700 170.100 81.600 173.400 ;
        RECT 85.950 172.950 88.050 175.050 ;
        RECT 11.100 167.100 12.900 167.850 ;
        RECT 13.950 166.950 16.050 169.050 ;
        RECT 17.100 167.100 18.900 167.850 ;
        RECT 19.950 166.950 22.050 169.050 ;
        RECT 25.950 166.950 28.050 169.050 ;
        RECT 10.950 163.950 13.050 166.050 ;
        RECT 14.850 162.900 15.900 165.900 ;
        RECT 16.950 163.950 19.050 166.050 ;
        RECT 20.100 165.150 21.900 165.900 ;
        RECT 32.700 164.100 33.600 169.350 ;
        RECT 35.100 167.100 36.900 167.850 ;
        RECT 41.100 167.100 42.900 167.850 ;
        RECT 50.100 167.100 51.900 167.850 ;
        RECT 52.950 166.950 55.050 169.050 ;
        RECT 56.100 167.100 57.900 167.850 ;
        RECT 58.950 166.950 64.050 169.050 ;
        RECT 71.100 167.100 72.900 167.850 ;
        RECT 73.950 166.950 76.050 169.050 ;
        RECT 79.950 168.450 82.050 169.050 ;
        RECT 86.550 168.450 87.450 172.950 ;
        RECT 98.100 171.000 99.900 179.400 ;
        RECT 106.950 172.950 109.050 175.050 ;
        RECT 113.400 174.300 115.200 179.400 ;
        RECT 119.400 174.300 121.200 179.400 ;
        RECT 113.400 172.950 121.200 174.300 ;
        RECT 122.400 173.400 124.200 179.400 ;
        RECT 98.100 169.350 102.300 171.000 ;
        RECT 77.100 167.100 78.900 167.850 ;
        RECT 79.950 167.550 87.450 168.450 ;
        RECT 79.950 166.950 82.050 167.550 ;
        RECT 92.100 167.100 93.900 167.850 ;
        RECT 98.100 167.100 99.900 167.850 ;
        RECT 34.950 163.950 37.050 166.050 ;
        RECT 40.800 163.950 43.050 166.050 ;
        RECT 49.950 163.950 52.050 166.050 ;
        RECT 53.100 165.150 54.900 165.900 ;
        RECT 55.950 163.950 58.050 166.050 ;
        RECT 14.850 159.600 16.050 162.900 ;
        RECT 31.950 160.950 34.050 163.050 ;
        RECT 37.950 160.950 40.200 163.050 ;
        RECT 14.700 147.600 16.500 159.600 ;
        RECT 32.700 154.800 33.600 159.900 ;
        RECT 38.100 159.150 39.900 159.900 ;
        RECT 59.700 159.600 60.600 165.900 ;
        RECT 70.950 163.950 73.050 166.050 ;
        RECT 74.100 165.150 75.900 165.900 ;
        RECT 76.950 163.950 79.050 166.050 ;
        RECT 80.700 159.600 81.600 165.900 ;
        RECT 91.950 163.950 94.050 166.050 ;
        RECT 97.950 163.950 100.050 166.050 ;
        RECT 101.400 164.100 102.300 169.350 ;
        RECT 107.550 166.050 108.450 172.950 ;
        RECT 122.400 171.300 123.600 173.400 ;
        RECT 119.850 170.250 123.600 171.300 ;
        RECT 140.100 171.000 141.900 179.400 ;
        RECT 165.000 173.400 166.800 179.400 ;
        RECT 119.850 170.100 121.050 170.250 ;
        RECT 140.100 169.350 144.300 171.000 ;
        RECT 165.000 170.100 166.050 173.400 ;
        RECT 185.100 171.000 186.900 179.400 ;
        RECT 205.200 175.050 207.000 179.400 ;
        RECT 205.200 173.400 210.600 175.050 ;
        RECT 185.100 169.350 189.300 171.000 ;
        RECT 209.700 170.100 210.600 173.400 ;
        RECT 214.950 172.950 217.050 175.050 ;
        RECT 112.950 166.950 115.050 169.050 ;
        RECT 116.100 167.100 117.900 167.850 ;
        RECT 118.950 166.950 121.050 169.050 ;
        RECT 122.100 167.100 123.900 167.850 ;
        RECT 134.100 167.100 135.900 167.850 ;
        RECT 140.100 167.100 141.900 167.850 ;
        RECT 106.950 163.950 109.050 166.050 ;
        RECT 113.100 165.150 114.900 165.900 ;
        RECT 115.950 163.950 118.050 166.050 ;
        RECT 94.950 160.950 97.050 163.050 ;
        RECT 100.950 160.950 106.050 163.050 ;
        RECT 119.100 162.900 120.150 165.900 ;
        RECT 121.950 163.950 124.050 166.050 ;
        RECT 133.950 163.950 136.050 166.050 ;
        RECT 139.950 163.950 142.050 166.050 ;
        RECT 143.400 164.100 144.300 169.350 ;
        RECT 157.800 166.950 160.050 169.050 ;
        RECT 161.250 167.100 162.900 167.850 ;
        RECT 163.800 166.950 166.050 169.050 ;
        RECT 167.100 167.100 168.750 167.850 ;
        RECT 169.950 166.950 172.050 169.050 ;
        RECT 179.100 167.100 180.900 167.850 ;
        RECT 185.100 167.100 186.900 167.850 ;
        RECT 158.100 165.150 159.900 165.900 ;
        RECT 160.950 163.950 163.050 166.050 ;
        RECT 50.400 158.700 58.200 159.600 ;
        RECT 32.700 153.900 39.300 154.800 ;
        RECT 32.700 153.600 33.600 153.900 ;
        RECT 31.800 147.600 33.600 153.600 ;
        RECT 37.800 153.600 39.300 153.900 ;
        RECT 37.800 147.600 39.600 153.600 ;
        RECT 50.400 147.600 52.200 158.700 ;
        RECT 56.400 147.600 58.200 158.700 ;
        RECT 59.400 147.600 61.200 159.600 ;
        RECT 71.400 158.700 79.200 159.600 ;
        RECT 71.400 147.600 73.200 158.700 ;
        RECT 77.400 147.600 79.200 158.700 ;
        RECT 80.400 147.600 82.200 159.600 ;
        RECT 95.100 159.150 96.900 159.900 ;
        RECT 101.400 154.800 102.300 159.900 ;
        RECT 118.950 159.600 120.150 162.900 ;
        RECT 136.950 160.950 139.050 163.050 ;
        RECT 142.950 160.950 148.050 163.050 ;
        RECT 164.100 162.900 164.850 165.900 ;
        RECT 166.950 163.950 169.050 166.050 ;
        RECT 170.100 165.150 171.750 165.900 ;
        RECT 178.800 163.950 181.050 166.050 ;
        RECT 184.950 163.950 187.050 166.050 ;
        RECT 188.400 164.100 189.300 169.350 ;
        RECT 200.100 167.100 201.900 167.850 ;
        RECT 202.950 166.950 205.050 169.050 ;
        RECT 208.950 168.450 211.050 169.050 ;
        RECT 215.550 168.450 216.450 172.950 ;
        RECT 226.200 172.200 228.000 179.400 ;
        RECT 206.100 167.100 207.900 167.850 ;
        RECT 208.950 167.550 216.450 168.450 ;
        RECT 224.400 171.300 228.000 172.200 ;
        RECT 208.950 166.950 211.050 167.550 ;
        RECT 224.400 167.100 225.600 171.300 ;
        RECT 245.100 171.000 246.900 179.400 ;
        RECT 253.950 172.950 256.050 175.050 ;
        RECT 260.400 174.300 262.200 179.400 ;
        RECT 266.400 174.300 268.200 179.400 ;
        RECT 260.400 172.950 268.200 174.300 ;
        RECT 269.400 173.400 271.200 179.400 ;
        RECT 284.400 176.400 286.200 179.400 ;
        RECT 245.100 169.350 249.300 171.000 ;
        RECT 239.100 167.100 240.900 167.850 ;
        RECT 245.100 167.100 246.900 167.850 ;
        RECT 199.950 163.950 202.050 166.050 ;
        RECT 203.100 165.150 204.900 165.900 ;
        RECT 205.950 163.950 208.050 166.050 ;
        RECT 163.950 161.400 164.850 162.900 ;
        RECT 160.800 160.500 164.850 161.400 ;
        RECT 181.950 160.950 184.050 163.050 ;
        RECT 187.950 160.950 193.050 163.050 ;
        RECT 95.700 153.900 102.300 154.800 ;
        RECT 95.700 153.600 97.200 153.900 ;
        RECT 95.400 147.600 97.200 153.600 ;
        RECT 101.400 153.600 102.300 153.900 ;
        RECT 101.400 147.600 103.200 153.600 ;
        RECT 118.500 147.600 120.300 159.600 ;
        RECT 137.100 159.150 138.900 159.900 ;
        RECT 143.400 154.800 144.300 159.900 ;
        RECT 137.700 153.900 144.300 154.800 ;
        RECT 137.700 153.600 139.200 153.900 ;
        RECT 137.400 147.600 139.200 153.600 ;
        RECT 143.400 153.600 144.300 153.900 ;
        RECT 143.400 147.600 145.200 153.600 ;
        RECT 157.800 148.500 159.600 159.600 ;
        RECT 160.800 149.400 162.600 160.500 ;
        RECT 163.800 158.400 171.600 159.300 ;
        RECT 182.100 159.150 183.900 159.900 ;
        RECT 163.800 148.500 165.600 158.400 ;
        RECT 157.800 147.600 165.600 148.500 ;
        RECT 169.800 147.600 171.600 158.400 ;
        RECT 188.400 154.800 189.300 159.900 ;
        RECT 209.700 159.600 210.600 165.900 ;
        RECT 221.100 164.100 222.900 164.850 ;
        RECT 223.950 163.950 226.050 166.050 ;
        RECT 227.100 164.100 228.900 164.850 ;
        RECT 238.950 163.950 241.050 166.050 ;
        RECT 244.950 163.950 247.050 166.050 ;
        RECT 248.400 164.100 249.300 169.350 ;
        RECT 254.550 163.050 255.450 172.950 ;
        RECT 269.400 171.300 270.600 173.400 ;
        RECT 274.950 172.950 277.050 175.050 ;
        RECT 266.850 170.250 270.600 171.300 ;
        RECT 266.850 170.100 268.050 170.250 ;
        RECT 259.950 166.950 262.050 169.050 ;
        RECT 263.100 167.100 264.900 167.850 ;
        RECT 265.950 166.950 268.050 169.050 ;
        RECT 269.100 167.100 270.900 167.850 ;
        RECT 260.100 165.150 261.900 165.900 ;
        RECT 262.950 163.950 265.050 166.050 ;
        RECT 220.950 160.950 223.050 163.050 ;
        RECT 182.700 153.900 189.300 154.800 ;
        RECT 182.700 153.600 184.200 153.900 ;
        RECT 182.400 147.600 184.200 153.600 ;
        RECT 188.400 153.600 189.300 153.900 ;
        RECT 200.400 158.700 208.200 159.600 ;
        RECT 188.400 147.600 190.200 153.600 ;
        RECT 200.400 147.600 202.200 158.700 ;
        RECT 206.400 147.600 208.200 158.700 ;
        RECT 209.400 147.600 211.200 159.600 ;
        RECT 224.400 153.600 225.600 162.900 ;
        RECT 226.950 160.950 229.050 163.050 ;
        RECT 241.950 160.950 244.200 163.050 ;
        RECT 247.950 160.950 250.050 163.050 ;
        RECT 253.950 160.950 256.050 163.050 ;
        RECT 266.100 162.900 267.150 165.900 ;
        RECT 268.950 163.950 271.050 166.050 ;
        RECT 242.100 159.150 243.900 159.900 ;
        RECT 248.400 154.800 249.300 159.900 ;
        RECT 265.950 159.600 267.150 162.900 ;
        RECT 242.700 153.900 249.300 154.800 ;
        RECT 242.700 153.600 244.200 153.900 ;
        RECT 224.400 147.600 226.200 153.600 ;
        RECT 242.400 147.600 244.200 153.600 ;
        RECT 248.400 153.600 249.300 153.900 ;
        RECT 248.400 147.600 250.200 153.600 ;
        RECT 265.500 147.600 267.300 159.600 ;
        RECT 275.550 154.050 276.450 172.950 ;
        RECT 280.950 169.950 283.050 172.050 ;
        RECT 281.100 168.150 282.900 168.900 ;
        RECT 284.400 167.100 285.600 176.400 ;
        RECT 302.100 171.000 303.900 179.400 ;
        RECT 322.200 175.050 324.000 179.400 ;
        RECT 322.200 173.400 327.600 175.050 ;
        RECT 302.100 169.350 306.300 171.000 ;
        RECT 326.700 170.100 327.600 173.400 ;
        RECT 338.400 174.300 340.200 179.400 ;
        RECT 344.400 174.300 346.200 179.400 ;
        RECT 338.400 172.950 346.200 174.300 ;
        RECT 347.400 173.400 349.200 179.400 ;
        RECT 359.400 174.300 361.200 179.400 ;
        RECT 365.400 174.300 367.200 179.400 ;
        RECT 347.400 171.300 348.600 173.400 ;
        RECT 359.400 172.950 367.200 174.300 ;
        RECT 368.400 173.400 370.200 179.400 ;
        RECT 368.400 171.300 369.600 173.400 ;
        RECT 344.850 170.250 348.600 171.300 ;
        RECT 365.850 170.250 369.600 171.300 ;
        RECT 386.100 171.000 387.900 179.400 ;
        RECT 406.200 172.200 408.000 179.400 ;
        RECT 422.400 176.400 424.200 179.400 ;
        RECT 440.400 176.400 442.200 179.400 ;
        RECT 422.400 173.100 423.600 176.400 ;
        RECT 404.400 171.300 408.000 172.200 ;
        RECT 344.850 170.100 346.050 170.250 ;
        RECT 365.850 170.100 367.050 170.250 ;
        RECT 386.100 169.350 390.300 171.000 ;
        RECT 296.100 167.100 297.900 167.850 ;
        RECT 302.100 167.100 303.900 167.850 ;
        RECT 283.950 163.950 289.050 166.050 ;
        RECT 295.950 163.950 298.050 166.050 ;
        RECT 301.950 163.950 304.050 166.050 ;
        RECT 305.400 164.100 306.300 169.350 ;
        RECT 317.100 167.100 318.900 167.850 ;
        RECT 319.950 166.950 322.050 169.050 ;
        RECT 323.100 167.100 324.900 167.850 ;
        RECT 325.950 166.950 331.050 169.050 ;
        RECT 337.950 166.950 340.050 169.050 ;
        RECT 341.100 167.100 342.900 167.850 ;
        RECT 343.950 166.950 346.050 169.050 ;
        RECT 347.100 167.100 348.900 167.850 ;
        RECT 358.950 166.950 361.050 169.050 ;
        RECT 362.100 167.100 363.900 167.850 ;
        RECT 364.950 166.950 367.050 169.050 ;
        RECT 368.100 167.100 369.900 167.850 ;
        RECT 380.100 167.100 381.900 167.850 ;
        RECT 386.100 167.100 387.900 167.850 ;
        RECT 316.950 163.950 319.050 166.050 ;
        RECT 320.100 165.150 321.900 165.900 ;
        RECT 322.950 163.950 325.050 166.050 ;
        RECT 274.950 151.950 277.050 154.050 ;
        RECT 284.400 153.600 285.600 162.900 ;
        RECT 298.950 160.950 301.050 163.050 ;
        RECT 304.950 162.450 307.050 163.050 ;
        RECT 304.950 162.000 312.450 162.450 ;
        RECT 304.950 161.550 313.050 162.000 ;
        RECT 304.950 160.950 307.050 161.550 ;
        RECT 299.100 159.150 300.900 159.900 ;
        RECT 305.400 154.800 306.300 159.900 ;
        RECT 310.950 157.950 313.050 161.550 ;
        RECT 326.700 159.600 327.600 165.900 ;
        RECT 338.100 165.150 339.900 165.900 ;
        RECT 340.950 163.950 343.050 166.050 ;
        RECT 344.100 162.900 345.150 165.900 ;
        RECT 346.950 163.950 349.200 166.050 ;
        RECT 359.100 165.150 360.900 165.900 ;
        RECT 361.950 163.950 364.050 166.050 ;
        RECT 365.100 162.900 366.150 165.900 ;
        RECT 367.950 163.950 370.050 166.050 ;
        RECT 379.800 163.950 382.050 166.050 ;
        RECT 385.950 163.950 388.050 166.050 ;
        RECT 389.400 164.100 390.300 169.350 ;
        RECT 404.400 167.100 405.600 171.300 ;
        RECT 421.950 169.950 424.050 172.050 ;
        RECT 436.950 169.950 439.050 172.050 ;
        RECT 418.950 166.950 421.050 169.050 ;
        RECT 401.100 164.100 402.900 164.850 ;
        RECT 403.950 163.950 406.050 166.050 ;
        RECT 422.700 165.900 423.900 168.900 ;
        RECT 424.950 166.950 427.050 169.050 ;
        RECT 437.100 168.150 438.900 168.900 ;
        RECT 440.400 167.100 441.600 176.400 ;
        RECT 454.800 173.400 456.600 179.400 ;
        RECT 455.400 171.300 456.600 173.400 ;
        RECT 457.800 174.300 459.600 179.400 ;
        RECT 463.800 174.300 465.600 179.400 ;
        RECT 457.800 172.950 465.600 174.300 ;
        RECT 478.200 175.050 480.000 179.400 ;
        RECT 478.200 173.400 483.600 175.050 ;
        RECT 455.400 170.250 459.150 171.300 ;
        RECT 457.950 170.100 459.150 170.250 ;
        RECT 482.700 170.100 483.600 173.400 ;
        RECT 494.400 174.300 496.200 179.400 ;
        RECT 500.400 174.300 502.200 179.400 ;
        RECT 494.400 172.950 502.200 174.300 ;
        RECT 503.400 173.400 505.200 179.400 ;
        RECT 525.000 173.400 526.800 179.400 ;
        RECT 541.800 176.400 543.600 179.400 ;
        RECT 487.950 169.950 490.050 172.050 ;
        RECT 503.400 171.300 504.600 173.400 ;
        RECT 500.850 170.250 504.600 171.300 ;
        RECT 500.850 170.100 502.050 170.250 ;
        RECT 511.950 169.950 514.050 172.050 ;
        RECT 525.000 170.100 526.050 173.400 ;
        RECT 535.950 172.950 538.050 175.050 ;
        RECT 455.100 167.100 456.900 167.850 ;
        RECT 457.950 166.950 460.050 169.050 ;
        RECT 461.100 167.100 462.900 167.850 ;
        RECT 463.950 166.950 466.050 169.050 ;
        RECT 473.100 167.100 474.900 167.850 ;
        RECT 475.950 166.950 478.050 169.050 ;
        RECT 479.100 167.100 480.900 167.850 ;
        RECT 481.950 166.950 487.050 169.050 ;
        RECT 419.100 165.150 420.900 165.900 ;
        RECT 407.100 164.100 408.900 164.850 ;
        RECT 343.950 159.600 345.150 162.900 ;
        RECT 364.950 159.600 366.150 162.900 ;
        RECT 382.950 160.950 385.050 163.050 ;
        RECT 388.950 160.950 394.050 163.050 ;
        RECT 400.950 160.950 403.050 163.050 ;
        RECT 317.400 158.700 325.200 159.600 ;
        RECT 299.700 153.900 306.300 154.800 ;
        RECT 299.700 153.600 301.200 153.900 ;
        RECT 284.400 147.600 286.200 153.600 ;
        RECT 299.400 147.600 301.200 153.600 ;
        RECT 305.400 153.600 306.300 153.900 ;
        RECT 305.400 147.600 307.200 153.600 ;
        RECT 317.400 147.600 319.200 158.700 ;
        RECT 323.400 147.600 325.200 158.700 ;
        RECT 326.400 147.600 328.200 159.600 ;
        RECT 343.500 147.600 345.300 159.600 ;
        RECT 364.500 147.600 366.300 159.600 ;
        RECT 383.100 159.150 384.900 159.900 ;
        RECT 389.400 154.800 390.300 159.900 ;
        RECT 383.700 153.900 390.300 154.800 ;
        RECT 383.700 153.600 385.200 153.900 ;
        RECT 383.400 147.600 385.200 153.600 ;
        RECT 389.400 153.600 390.300 153.900 ;
        RECT 404.400 153.600 405.600 162.900 ;
        RECT 406.950 160.950 409.050 163.050 ;
        RECT 422.700 160.650 424.050 165.900 ;
        RECT 425.100 165.150 426.900 165.900 ;
        RECT 436.950 163.950 442.050 166.050 ;
        RECT 454.950 163.950 457.050 166.050 ;
        RECT 458.850 162.900 459.900 165.900 ;
        RECT 460.950 163.950 463.050 166.050 ;
        RECT 464.100 165.150 465.900 165.900 ;
        RECT 472.950 163.950 475.050 166.050 ;
        RECT 476.100 165.150 477.900 165.900 ;
        RECT 478.950 163.950 481.050 166.050 ;
        RECT 422.700 159.600 425.400 160.650 ;
        RECT 389.400 147.600 391.200 153.600 ;
        RECT 404.400 147.600 406.200 153.600 ;
        RECT 423.600 147.600 425.400 159.600 ;
        RECT 440.400 153.600 441.600 162.900 ;
        RECT 458.850 159.600 460.050 162.900 ;
        RECT 482.700 159.600 483.600 165.900 ;
        RECT 440.400 147.600 442.200 153.600 ;
        RECT 458.700 147.600 460.500 159.600 ;
        RECT 473.400 158.700 481.200 159.600 ;
        RECT 473.400 147.600 475.200 158.700 ;
        RECT 479.400 147.600 481.200 158.700 ;
        RECT 482.400 147.600 484.200 159.600 ;
        RECT 488.550 151.050 489.450 169.950 ;
        RECT 493.800 166.950 496.050 169.050 ;
        RECT 497.100 167.100 498.900 167.850 ;
        RECT 499.950 166.950 502.200 169.050 ;
        RECT 503.100 167.100 504.900 167.850 ;
        RECT 508.950 166.950 511.050 169.050 ;
        RECT 494.100 165.150 495.900 165.900 ;
        RECT 496.950 163.950 499.050 166.050 ;
        RECT 500.100 162.900 501.150 165.900 ;
        RECT 499.950 159.600 501.150 162.900 ;
        RECT 509.550 160.050 510.450 166.950 ;
        RECT 487.950 148.950 490.050 151.050 ;
        RECT 499.500 147.600 501.300 159.600 ;
        RECT 508.950 157.950 511.050 160.050 ;
        RECT 512.550 151.050 513.450 169.950 ;
        RECT 517.950 166.950 520.050 169.050 ;
        RECT 521.250 167.100 522.900 167.850 ;
        RECT 523.950 166.950 526.050 169.050 ;
        RECT 527.100 167.100 528.750 167.850 ;
        RECT 529.950 166.950 532.050 169.050 ;
        RECT 518.100 165.150 519.900 165.900 ;
        RECT 520.800 163.950 523.050 166.050 ;
        RECT 524.100 162.900 524.850 165.900 ;
        RECT 526.950 163.950 529.050 166.050 ;
        RECT 530.100 165.150 531.750 165.900 ;
        RECT 523.950 161.400 524.850 162.900 ;
        RECT 520.800 160.500 524.850 161.400 ;
        RECT 511.950 148.950 514.050 151.050 ;
        RECT 517.800 148.500 519.600 159.600 ;
        RECT 520.800 149.400 522.600 160.500 ;
        RECT 536.550 160.050 537.450 172.950 ;
        RECT 542.400 167.100 543.600 176.400 ;
        RECT 548.550 173.400 550.350 179.400 ;
        RECT 556.650 176.400 558.450 179.400 ;
        RECT 564.450 176.400 566.250 179.400 ;
        RECT 572.250 177.300 574.050 179.400 ;
        RECT 572.250 176.400 576.000 177.300 ;
        RECT 556.650 175.500 557.700 176.400 ;
        RECT 553.950 174.300 557.700 175.500 ;
        RECT 565.200 174.600 566.250 176.400 ;
        RECT 574.950 175.500 576.000 176.400 ;
        RECT 553.950 173.400 556.050 174.300 ;
        RECT 544.950 169.950 547.050 172.050 ;
        RECT 548.550 169.050 549.750 173.400 ;
        RECT 561.150 172.200 562.950 174.000 ;
        RECT 565.200 173.550 570.150 174.600 ;
        RECT 568.350 172.800 570.150 173.550 ;
        RECT 571.650 172.800 573.450 174.600 ;
        RECT 574.950 173.400 577.050 175.500 ;
        RECT 580.050 173.400 581.850 179.400 ;
        RECT 595.800 176.400 597.600 179.400 ;
        RECT 611.400 176.400 613.200 179.400 ;
        RECT 562.050 171.900 562.950 172.200 ;
        RECT 572.100 171.900 573.150 172.800 ;
        RECT 562.050 171.000 573.150 171.900 ;
        RECT 562.050 170.100 562.950 171.000 ;
        RECT 572.100 169.800 573.150 171.000 ;
        RECT 545.100 168.150 546.900 168.900 ;
        RECT 548.550 166.950 549.900 169.050 ;
        RECT 550.950 166.950 553.050 169.050 ;
        RECT 554.100 167.250 554.850 169.050 ;
        RECT 562.950 166.950 565.050 169.050 ;
        RECT 568.950 166.950 571.050 169.050 ;
        RECT 572.100 168.600 579.000 169.800 ;
        RECT 572.100 168.000 573.900 168.600 ;
        RECT 578.100 167.850 579.000 168.600 ;
        RECT 575.100 167.100 576.900 167.700 ;
        RECT 538.950 163.950 544.050 166.050 ;
        RECT 523.800 158.400 531.600 159.300 ;
        RECT 523.800 148.500 525.600 158.400 ;
        RECT 517.800 147.600 525.600 148.500 ;
        RECT 529.800 147.600 531.600 158.400 ;
        RECT 535.950 157.950 538.050 160.050 ;
        RECT 542.400 153.600 543.600 162.900 ;
        RECT 541.800 147.600 543.600 153.600 ;
        RECT 548.550 159.600 549.750 166.950 ;
        RECT 572.100 166.200 576.900 167.100 ;
        RECT 575.100 165.900 576.900 166.200 ;
        RECT 578.100 166.050 579.900 167.850 ;
        RECT 550.950 161.400 552.750 163.200 ;
        RECT 551.850 160.200 556.050 161.400 ;
        RECT 562.050 160.200 562.950 165.900 ;
        RECT 570.750 161.100 572.550 161.400 ;
        RECT 548.550 147.600 550.350 159.600 ;
        RECT 553.950 159.300 556.050 160.200 ;
        RECT 556.950 159.300 562.950 160.200 ;
        RECT 564.150 160.800 572.550 161.100 ;
        RECT 580.950 160.800 581.850 173.400 ;
        RECT 596.400 173.100 597.600 176.400 ;
        RECT 612.300 172.200 613.200 176.400 ;
        RECT 617.400 173.400 619.200 179.400 ;
        RECT 595.950 169.950 598.050 172.050 ;
        RECT 612.300 171.300 615.750 172.200 ;
        RECT 613.950 170.400 615.750 171.300 ;
        RECT 592.800 166.950 595.050 169.050 ;
        RECT 596.100 165.900 597.300 168.900 ;
        RECT 598.950 166.950 601.050 169.050 ;
        RECT 608.100 168.150 609.900 168.900 ;
        RECT 610.950 166.950 613.050 169.050 ;
        RECT 593.100 165.150 594.900 165.900 ;
        RECT 564.150 160.200 581.850 160.800 ;
        RECT 595.950 160.650 597.300 165.900 ;
        RECT 599.100 165.150 600.900 165.900 ;
        RECT 611.100 165.150 612.900 165.900 ;
        RECT 614.700 162.600 615.600 170.400 ;
        RECT 618.000 167.100 619.050 173.400 ;
        RECT 622.950 172.950 625.050 175.050 ;
        RECT 616.950 163.950 619.050 166.050 ;
        RECT 613.800 162.000 615.600 162.600 ;
        RECT 556.950 158.400 557.850 159.300 ;
        RECT 555.150 156.600 557.850 158.400 ;
        RECT 558.750 158.100 560.550 158.400 ;
        RECT 564.150 158.100 565.050 160.200 ;
        RECT 570.750 159.600 581.850 160.200 ;
        RECT 558.750 157.200 565.050 158.100 ;
        RECT 565.950 158.700 567.750 159.300 ;
        RECT 565.950 157.500 573.450 158.700 ;
        RECT 558.750 156.600 560.550 157.200 ;
        RECT 572.250 156.600 573.450 157.500 ;
        RECT 553.950 153.600 557.850 155.700 ;
        RECT 562.950 155.550 564.750 156.300 ;
        RECT 567.750 155.550 569.550 156.300 ;
        RECT 562.950 154.500 569.550 155.550 ;
        RECT 572.250 154.500 577.050 156.600 ;
        RECT 556.050 147.600 557.850 153.600 ;
        RECT 563.850 147.600 565.650 154.500 ;
        RECT 572.250 153.600 573.450 154.500 ;
        RECT 571.650 147.600 573.450 153.600 ;
        RECT 580.050 147.600 581.850 159.600 ;
        RECT 594.600 159.600 597.300 160.650 ;
        RECT 608.400 160.800 615.600 162.000 ;
        RECT 608.400 159.600 609.600 160.800 ;
        RECT 614.700 160.650 615.600 160.800 ;
        RECT 616.950 159.600 618.300 162.900 ;
        RECT 594.600 147.600 596.400 159.600 ;
        RECT 608.400 147.600 610.200 159.600 ;
        RECT 615.900 158.100 618.300 159.600 ;
        RECT 615.900 147.600 617.700 158.100 ;
        RECT 623.550 157.050 624.450 172.950 ;
        RECT 635.100 171.000 636.900 179.400 ;
        RECT 655.200 172.200 657.000 179.400 ;
        RECT 632.700 169.350 636.900 171.000 ;
        RECT 653.400 171.300 657.000 172.200 ;
        RECT 671.400 176.400 673.200 179.400 ;
        RECT 632.700 164.100 633.600 169.350 ;
        RECT 635.100 167.100 636.900 167.850 ;
        RECT 641.100 167.100 642.900 167.850 ;
        RECT 653.400 167.100 654.600 171.300 ;
        RECT 667.950 169.950 670.050 172.050 ;
        RECT 668.100 168.150 669.900 168.900 ;
        RECT 671.400 167.100 672.600 176.400 ;
        RECT 683.400 174.300 685.200 179.400 ;
        RECT 689.400 174.300 691.200 179.400 ;
        RECT 683.400 172.950 691.200 174.300 ;
        RECT 692.400 173.400 694.200 179.400 ;
        RECT 706.800 176.400 708.600 179.400 ;
        RECT 692.400 171.300 693.600 173.400 ;
        RECT 689.850 170.250 693.600 171.300 ;
        RECT 689.850 170.100 691.050 170.250 ;
        RECT 682.950 166.950 685.050 169.050 ;
        RECT 686.100 167.100 687.900 167.850 ;
        RECT 688.950 166.950 691.050 169.050 ;
        RECT 692.100 167.100 693.900 167.850 ;
        RECT 707.400 167.100 708.600 176.400 ;
        RECT 722.400 176.400 724.200 179.400 ;
        RECT 709.950 169.950 712.050 172.050 ;
        RECT 718.950 169.950 721.050 172.050 ;
        RECT 710.100 168.150 711.900 168.900 ;
        RECT 719.100 168.150 720.900 168.900 ;
        RECT 722.400 167.100 723.600 176.400 ;
        RECT 739.200 175.050 741.000 179.400 ;
        RECT 758.400 176.400 760.200 179.400 ;
        RECT 739.200 173.400 744.600 175.050 ;
        RECT 743.700 170.100 744.600 173.400 ;
        RECT 754.950 169.950 757.050 172.050 ;
        RECT 734.100 167.100 735.900 167.850 ;
        RECT 736.950 166.950 739.050 169.050 ;
        RECT 740.100 167.100 741.900 167.850 ;
        RECT 742.950 166.950 745.050 169.050 ;
        RECT 755.100 168.150 756.900 168.900 ;
        RECT 758.400 167.100 759.600 176.400 ;
        RECT 770.400 174.300 772.200 179.400 ;
        RECT 776.400 174.300 778.200 179.400 ;
        RECT 770.400 172.950 778.200 174.300 ;
        RECT 779.400 173.400 781.200 179.400 ;
        RECT 784.950 175.950 787.050 178.050 ;
        RECT 763.950 169.950 766.050 172.050 ;
        RECT 779.400 171.300 780.600 173.400 ;
        RECT 776.850 170.250 780.600 171.300 ;
        RECT 776.850 170.100 778.050 170.250 ;
        RECT 634.950 163.950 637.050 166.050 ;
        RECT 640.950 163.950 643.050 166.050 ;
        RECT 650.100 164.100 651.900 164.850 ;
        RECT 652.950 163.950 655.050 166.050 ;
        RECT 656.100 164.100 657.900 164.850 ;
        RECT 670.950 163.950 676.050 166.050 ;
        RECT 683.100 165.150 684.900 165.900 ;
        RECT 685.950 163.950 688.050 166.050 ;
        RECT 625.950 162.450 630.000 163.050 ;
        RECT 631.950 162.450 634.050 163.050 ;
        RECT 625.950 161.550 634.050 162.450 ;
        RECT 625.950 160.950 630.000 161.550 ;
        RECT 631.950 160.950 634.050 161.550 ;
        RECT 637.800 160.950 640.050 163.050 ;
        RECT 649.950 160.950 652.050 163.050 ;
        RECT 622.950 154.950 625.050 157.050 ;
        RECT 632.700 154.800 633.600 159.900 ;
        RECT 638.100 159.150 639.900 159.900 ;
        RECT 632.700 153.900 639.300 154.800 ;
        RECT 632.700 153.600 633.600 153.900 ;
        RECT 631.800 147.600 633.600 153.600 ;
        RECT 637.800 153.600 639.300 153.900 ;
        RECT 653.400 153.600 654.600 162.900 ;
        RECT 655.950 157.950 658.050 163.050 ;
        RECT 689.100 162.900 690.150 165.900 ;
        RECT 691.800 163.950 694.050 166.050 ;
        RECT 703.950 163.950 709.050 166.050 ;
        RECT 721.950 163.950 727.050 166.050 ;
        RECT 733.950 163.950 736.050 166.050 ;
        RECT 737.100 165.150 738.900 165.900 ;
        RECT 739.950 163.950 742.050 166.050 ;
        RECT 671.400 153.600 672.600 162.900 ;
        RECT 688.950 159.600 690.150 162.900 ;
        RECT 637.800 147.600 639.600 153.600 ;
        RECT 653.400 147.600 655.200 153.600 ;
        RECT 671.400 147.600 673.200 153.600 ;
        RECT 688.500 147.600 690.300 159.600 ;
        RECT 707.400 153.600 708.600 162.900 ;
        RECT 706.800 147.600 708.600 153.600 ;
        RECT 722.400 153.600 723.600 162.900 ;
        RECT 743.700 159.600 744.600 165.900 ;
        RECT 754.950 163.950 760.050 166.050 ;
        RECT 734.400 158.700 742.200 159.600 ;
        RECT 722.400 147.600 724.200 153.600 ;
        RECT 734.400 147.600 736.200 158.700 ;
        RECT 740.400 147.600 742.200 158.700 ;
        RECT 743.400 147.600 745.200 159.600 ;
        RECT 758.400 153.600 759.600 162.900 ;
        RECT 764.550 160.050 765.450 169.950 ;
        RECT 769.950 166.950 772.050 169.050 ;
        RECT 773.100 167.100 774.900 167.850 ;
        RECT 775.950 166.950 778.050 169.050 ;
        RECT 779.100 167.100 780.900 167.850 ;
        RECT 770.100 165.150 771.900 165.900 ;
        RECT 772.950 163.950 775.050 166.050 ;
        RECT 776.100 162.900 777.150 165.900 ;
        RECT 778.950 163.950 781.050 166.050 ;
        RECT 763.950 157.950 766.050 160.050 ;
        RECT 775.950 159.600 777.150 162.900 ;
        RECT 758.400 147.600 760.200 153.600 ;
        RECT 775.500 147.600 777.300 159.600 ;
        RECT 785.550 151.050 786.450 175.950 ;
        RECT 791.400 174.300 793.200 179.400 ;
        RECT 797.400 174.300 799.200 179.400 ;
        RECT 791.400 172.950 799.200 174.300 ;
        RECT 800.400 173.400 802.200 179.400 ;
        RECT 815.400 176.400 817.200 179.400 ;
        RECT 800.400 171.300 801.600 173.400 ;
        RECT 805.950 172.950 808.050 175.050 ;
        RECT 815.400 173.100 816.600 176.400 ;
        RECT 823.950 175.950 826.050 178.050 ;
        RECT 797.850 170.250 801.600 171.300 ;
        RECT 797.850 170.100 799.050 170.250 ;
        RECT 790.950 166.950 793.050 169.050 ;
        RECT 794.100 167.100 795.900 167.850 ;
        RECT 796.950 166.950 799.050 169.050 ;
        RECT 800.100 167.100 801.900 167.850 ;
        RECT 791.100 165.150 792.900 165.900 ;
        RECT 793.950 163.950 796.050 166.050 ;
        RECT 797.100 162.900 798.150 165.900 ;
        RECT 799.950 163.950 802.050 166.050 ;
        RECT 796.950 159.600 798.150 162.900 ;
        RECT 784.950 148.950 787.050 151.050 ;
        RECT 796.500 147.600 798.300 159.600 ;
        RECT 806.550 154.050 807.450 172.950 ;
        RECT 814.950 169.950 817.050 172.050 ;
        RECT 811.950 166.950 814.050 169.050 ;
        RECT 815.700 165.900 816.900 168.900 ;
        RECT 817.950 166.950 820.050 169.050 ;
        RECT 812.100 165.150 813.900 165.900 ;
        RECT 815.700 160.650 817.050 165.900 ;
        RECT 818.100 165.150 819.900 165.900 ;
        RECT 815.700 159.600 818.400 160.650 ;
        RECT 805.950 151.950 808.050 154.050 ;
        RECT 816.600 147.600 818.400 159.600 ;
        RECT 824.550 157.050 825.450 175.950 ;
        RECT 830.400 174.300 832.200 179.400 ;
        RECT 836.400 174.300 838.200 179.400 ;
        RECT 830.400 172.950 838.200 174.300 ;
        RECT 839.400 173.400 841.200 179.400 ;
        RECT 839.400 171.300 840.600 173.400 ;
        RECT 847.950 172.950 850.050 175.050 ;
        RECT 836.850 170.250 840.600 171.300 ;
        RECT 836.850 170.100 838.050 170.250 ;
        RECT 829.950 166.950 832.050 169.050 ;
        RECT 833.100 167.100 834.900 167.850 ;
        RECT 835.950 166.950 838.050 169.050 ;
        RECT 839.100 167.100 840.900 167.850 ;
        RECT 844.950 166.950 847.050 169.050 ;
        RECT 830.100 165.150 831.900 165.900 ;
        RECT 832.950 163.950 835.050 166.050 ;
        RECT 836.100 162.900 837.150 165.900 ;
        RECT 838.950 163.950 841.050 166.050 ;
        RECT 835.950 159.600 837.150 162.900 ;
        RECT 845.550 160.050 846.450 166.950 ;
        RECT 823.950 154.950 826.050 157.050 ;
        RECT 835.500 147.600 837.300 159.600 ;
        RECT 844.950 157.950 847.050 160.050 ;
        RECT 848.550 151.050 849.450 172.950 ;
        RECT 847.950 148.950 850.050 151.050 ;
        RECT 10.800 137.400 12.600 143.400 ;
        RECT 11.400 128.100 12.600 137.400 ;
        RECT 23.400 132.300 25.200 143.400 ;
        RECT 29.400 132.300 31.200 143.400 ;
        RECT 23.400 131.400 31.200 132.300 ;
        RECT 32.400 131.400 34.200 143.400 ;
        RECT 37.950 139.950 40.050 142.050 ;
        RECT 10.950 124.950 16.050 127.050 ;
        RECT 22.950 124.950 25.050 127.050 ;
        RECT 26.100 125.100 27.900 125.850 ;
        RECT 28.950 124.950 31.050 127.050 ;
        RECT 32.700 125.100 33.600 131.400 ;
        RECT 11.400 114.600 12.600 123.900 ;
        RECT 23.100 123.150 24.900 123.900 ;
        RECT 14.100 122.100 15.900 122.850 ;
        RECT 25.950 121.950 28.050 124.050 ;
        RECT 29.100 123.150 30.900 123.900 ;
        RECT 31.950 123.450 34.050 124.050 ;
        RECT 38.550 123.450 39.450 139.950 ;
        RECT 47.400 137.400 49.200 143.400 ;
        RECT 47.700 137.100 49.200 137.400 ;
        RECT 53.400 137.400 55.200 143.400 ;
        RECT 68.400 137.400 70.200 143.400 ;
        RECT 53.400 137.100 54.300 137.400 ;
        RECT 47.700 136.200 54.300 137.100 ;
        RECT 68.700 137.100 70.200 137.400 ;
        RECT 74.400 137.400 76.200 143.400 ;
        RECT 74.400 137.100 75.300 137.400 ;
        RECT 68.700 136.200 75.300 137.100 ;
        RECT 47.100 131.100 48.900 131.850 ;
        RECT 53.400 131.100 54.300 136.200 ;
        RECT 68.100 131.100 69.900 131.850 ;
        RECT 74.400 131.100 75.300 136.200 ;
        RECT 92.700 131.400 94.500 143.400 ;
        RECT 103.950 139.950 106.050 142.050 ;
        RECT 104.550 133.050 105.450 139.950 ;
        RECT 110.400 137.400 112.200 143.400 ;
        RECT 110.700 137.100 112.200 137.400 ;
        RECT 116.400 137.400 118.200 143.400 ;
        RECT 116.400 137.100 117.300 137.400 ;
        RECT 110.700 136.200 117.300 137.100 ;
        RECT 46.950 127.950 49.050 130.050 ;
        RECT 52.950 129.450 55.050 130.050 ;
        RECT 57.000 129.450 61.050 130.050 ;
        RECT 52.950 128.550 61.050 129.450 ;
        RECT 52.950 127.950 55.050 128.550 ;
        RECT 57.000 127.950 61.050 128.550 ;
        RECT 67.950 127.950 70.050 130.050 ;
        RECT 73.950 127.950 79.050 130.050 ;
        RECT 92.850 128.100 94.050 131.400 ;
        RECT 103.950 130.950 106.050 133.050 ;
        RECT 110.100 131.100 111.900 131.850 ;
        RECT 116.400 131.100 117.300 136.200 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 43.950 124.950 46.050 127.050 ;
        RECT 49.950 124.950 52.050 127.050 ;
        RECT 31.950 122.550 39.450 123.450 ;
        RECT 44.100 123.150 45.900 123.900 ;
        RECT 50.100 123.150 51.900 123.900 ;
        RECT 31.950 121.950 34.050 122.550 ;
        RECT 53.400 121.650 54.300 126.900 ;
        RECT 64.800 124.950 67.050 127.050 ;
        RECT 70.950 124.950 73.200 127.050 ;
        RECT 65.100 123.150 66.900 123.900 ;
        RECT 71.100 123.150 72.900 123.900 ;
        RECT 74.400 121.650 75.300 126.900 ;
        RECT 88.950 124.950 91.050 127.050 ;
        RECT 92.850 125.100 93.900 128.100 ;
        RECT 109.950 127.950 112.050 130.050 ;
        RECT 115.950 127.950 121.050 130.050 ;
        RECT 94.950 124.950 97.200 127.050 ;
        RECT 98.100 125.100 99.900 125.850 ;
        RECT 106.950 124.950 109.200 127.050 ;
        RECT 112.950 124.950 115.050 127.050 ;
        RECT 89.100 123.150 90.900 123.900 ;
        RECT 91.950 121.950 94.050 124.050 ;
        RECT 95.100 123.150 96.900 123.900 ;
        RECT 97.950 121.950 100.200 124.050 ;
        RECT 107.100 123.150 108.900 123.900 ;
        RECT 113.100 123.150 114.900 123.900 ;
        RECT 116.400 121.650 117.300 126.900 ;
        RECT 13.950 118.950 16.050 121.050 ;
        RECT 32.700 117.600 33.600 120.900 ;
        RECT 10.800 111.600 12.600 114.600 ;
        RECT 28.200 115.950 33.600 117.600 ;
        RECT 50.100 120.000 54.300 121.650 ;
        RECT 71.100 120.000 75.300 121.650 ;
        RECT 91.950 120.750 93.150 120.900 ;
        RECT 28.200 111.600 30.000 115.950 ;
        RECT 50.100 111.600 51.900 120.000 ;
        RECT 71.100 111.600 72.900 120.000 ;
        RECT 89.400 119.700 93.150 120.750 ;
        RECT 113.100 120.000 117.300 121.650 ;
        RECT 122.550 121.050 123.450 133.950 ;
        RECT 128.400 132.300 130.200 143.400 ;
        RECT 134.400 132.300 136.200 143.400 ;
        RECT 128.400 131.400 136.200 132.300 ;
        RECT 137.400 131.400 139.200 143.400 ;
        RECT 145.950 139.950 148.050 142.050 ;
        RECT 127.950 124.950 130.050 127.050 ;
        RECT 131.100 125.100 132.900 125.850 ;
        RECT 133.950 124.950 136.050 127.050 ;
        RECT 137.700 125.100 138.600 131.400 ;
        RECT 128.100 123.150 129.900 123.900 ;
        RECT 89.400 117.600 90.600 119.700 ;
        RECT 88.800 111.600 90.600 117.600 ;
        RECT 91.800 116.700 99.600 118.050 ;
        RECT 91.800 111.600 93.600 116.700 ;
        RECT 97.800 111.600 99.600 116.700 ;
        RECT 113.100 111.600 114.900 120.000 ;
        RECT 121.950 118.950 124.050 121.050 ;
        RECT 130.950 118.950 133.050 124.050 ;
        RECT 134.100 123.150 135.900 123.900 ;
        RECT 136.950 123.450 139.050 124.050 ;
        RECT 136.950 122.550 144.450 123.450 ;
        RECT 136.950 121.950 139.050 122.550 ;
        RECT 137.700 117.600 138.600 120.900 ;
        RECT 133.200 115.950 138.600 117.600 ;
        RECT 133.200 111.600 135.000 115.950 ;
        RECT 143.550 115.050 144.450 122.550 ;
        RECT 146.550 121.050 147.450 139.950 ;
        RECT 155.700 131.400 157.500 143.400 ;
        RECT 174.600 131.400 176.400 143.400 ;
        RECT 194.700 131.400 196.500 143.400 ;
        RECT 211.800 137.400 213.600 143.400 ;
        RECT 155.850 128.100 157.050 131.400 ;
        RECT 174.600 130.350 177.300 131.400 ;
        RECT 151.950 124.950 154.050 127.050 ;
        RECT 155.850 125.100 156.900 128.100 ;
        RECT 157.950 124.950 160.050 127.050 ;
        RECT 161.100 125.100 162.900 125.850 ;
        RECT 173.100 125.100 174.900 125.850 ;
        RECT 175.950 125.100 177.300 130.350 ;
        RECT 184.950 127.950 187.050 130.050 ;
        RECT 194.850 128.100 196.050 131.400 ;
        RECT 212.400 128.100 213.600 137.400 ;
        RECT 228.300 132.900 230.100 143.400 ;
        RECT 227.700 131.400 230.100 132.900 ;
        RECT 235.800 131.400 237.600 143.400 ;
        RECT 249.600 131.400 251.400 143.400 ;
        RECT 227.700 128.100 229.050 131.400 ;
        RECT 230.400 130.200 231.300 130.350 ;
        RECT 236.400 130.200 237.600 131.400 ;
        RECT 230.400 129.000 237.600 130.200 ;
        RECT 248.700 130.350 251.400 131.400 ;
        RECT 267.600 131.400 269.400 143.400 ;
        RECT 281.400 131.400 283.200 143.400 ;
        RECT 288.900 132.900 290.700 143.400 ;
        RECT 288.900 131.400 291.300 132.900 ;
        RECT 304.800 131.400 306.600 143.400 ;
        RECT 307.800 132.300 309.600 143.400 ;
        RECT 313.800 132.300 315.600 143.400 ;
        RECT 326.400 137.400 328.200 143.400 ;
        RECT 326.700 137.100 328.200 137.400 ;
        RECT 332.400 137.400 334.200 143.400 ;
        RECT 347.400 137.400 349.200 143.400 ;
        RECT 332.400 137.100 333.300 137.400 ;
        RECT 326.700 136.200 333.300 137.100 ;
        RECT 307.800 131.400 315.600 132.300 ;
        RECT 267.600 130.350 270.300 131.400 ;
        RECT 230.400 128.400 232.200 129.000 ;
        RECT 179.100 125.100 180.900 125.850 ;
        RECT 152.100 123.150 153.900 123.900 ;
        RECT 154.800 121.950 157.050 124.050 ;
        RECT 158.100 123.150 159.900 123.900 ;
        RECT 160.950 121.950 163.200 124.050 ;
        RECT 172.950 121.950 175.200 124.050 ;
        RECT 176.100 122.100 177.300 125.100 ;
        RECT 178.950 121.950 181.050 124.050 ;
        RECT 185.550 121.050 186.450 127.950 ;
        RECT 190.950 124.950 193.200 127.050 ;
        RECT 194.850 125.100 195.900 128.100 ;
        RECT 196.950 124.950 199.050 127.050 ;
        RECT 200.100 125.100 201.900 125.850 ;
        RECT 211.950 124.950 217.050 127.050 ;
        RECT 221.100 126.450 225.000 127.050 ;
        RECT 226.950 126.450 229.050 127.050 ;
        RECT 221.100 125.550 229.050 126.450 ;
        RECT 221.100 124.950 225.000 125.550 ;
        RECT 226.950 124.950 229.050 125.550 ;
        RECT 191.100 123.150 192.900 123.900 ;
        RECT 193.950 121.950 196.200 124.050 ;
        RECT 197.100 123.150 198.900 123.900 ;
        RECT 199.950 121.950 202.050 124.050 ;
        RECT 145.950 118.950 148.050 121.050 ;
        RECT 154.950 120.750 156.150 120.900 ;
        RECT 152.400 119.700 156.150 120.750 ;
        RECT 152.400 117.600 153.600 119.700 ;
        RECT 175.950 118.950 178.050 121.050 ;
        RECT 184.950 118.950 187.050 121.050 ;
        RECT 193.950 120.750 195.150 120.900 ;
        RECT 191.400 119.700 195.150 120.750 ;
        RECT 143.100 112.950 145.200 115.050 ;
        RECT 151.800 111.600 153.600 117.600 ;
        RECT 154.800 116.700 162.600 118.050 ;
        RECT 154.800 111.600 156.600 116.700 ;
        RECT 160.800 111.600 162.600 116.700 ;
        RECT 176.400 114.600 177.600 117.900 ;
        RECT 191.400 117.600 192.600 119.700 ;
        RECT 175.800 111.600 177.600 114.600 ;
        RECT 190.800 111.600 192.600 117.600 ;
        RECT 193.800 116.700 201.600 118.050 ;
        RECT 193.800 111.600 195.600 116.700 ;
        RECT 199.800 111.600 201.600 116.700 ;
        RECT 212.400 114.600 213.600 123.900 ;
        RECT 215.100 122.100 216.900 122.850 ;
        RECT 214.950 118.950 217.050 121.050 ;
        RECT 226.950 117.600 228.000 123.900 ;
        RECT 230.400 120.600 231.300 128.400 ;
        RECT 233.100 125.100 234.900 125.850 ;
        RECT 245.100 125.100 246.900 125.850 ;
        RECT 248.700 125.100 250.050 130.350 ;
        RECT 251.100 125.100 252.900 125.850 ;
        RECT 266.100 125.100 267.900 125.850 ;
        RECT 268.950 125.100 270.300 130.350 ;
        RECT 281.400 130.200 282.600 131.400 ;
        RECT 287.700 130.200 288.600 130.350 ;
        RECT 281.400 129.000 288.600 130.200 ;
        RECT 286.800 128.400 288.600 129.000 ;
        RECT 272.100 125.100 273.900 125.850 ;
        RECT 284.100 125.100 285.900 125.850 ;
        RECT 232.950 121.950 235.050 124.050 ;
        RECT 236.100 122.100 237.900 122.850 ;
        RECT 244.950 121.950 247.050 124.050 ;
        RECT 248.700 122.100 249.900 125.100 ;
        RECT 250.950 121.950 253.050 124.050 ;
        RECT 265.950 121.950 268.050 124.050 ;
        RECT 269.100 122.100 270.300 125.100 ;
        RECT 271.950 121.950 277.050 124.050 ;
        RECT 281.100 122.100 282.900 122.850 ;
        RECT 283.950 121.950 286.200 124.050 ;
        RECT 230.250 119.700 232.050 120.600 ;
        RECT 230.250 118.800 233.700 119.700 ;
        RECT 235.950 118.950 241.050 121.050 ;
        RECT 247.950 118.950 250.050 121.050 ;
        RECT 268.950 118.950 271.050 121.050 ;
        RECT 280.950 118.950 283.050 121.050 ;
        RECT 287.700 120.600 288.600 128.400 ;
        RECT 289.950 128.100 291.300 131.400 ;
        RECT 289.950 124.950 292.050 127.050 ;
        RECT 305.400 125.100 306.300 131.400 ;
        RECT 326.100 131.100 327.900 131.850 ;
        RECT 332.400 131.100 333.300 136.200 ;
        RECT 325.950 127.950 328.050 130.050 ;
        RECT 331.950 129.450 334.050 130.050 ;
        RECT 331.950 128.550 339.450 129.450 ;
        RECT 331.950 127.950 334.050 128.550 ;
        RECT 307.950 124.950 310.050 127.050 ;
        RECT 311.100 125.100 312.900 125.850 ;
        RECT 313.950 124.950 316.050 127.050 ;
        RECT 322.950 124.950 325.050 127.050 ;
        RECT 328.950 124.950 331.050 127.050 ;
        RECT 286.950 119.700 288.750 120.600 ;
        RECT 211.800 111.600 213.600 114.600 ;
        RECT 226.800 111.600 228.600 117.600 ;
        RECT 232.800 114.600 233.700 118.800 ;
        RECT 285.300 118.800 288.750 119.700 ;
        RECT 248.400 114.600 249.600 117.900 ;
        RECT 269.400 114.600 270.600 117.900 ;
        RECT 285.300 114.600 286.200 118.800 ;
        RECT 291.000 117.600 292.050 123.900 ;
        RECT 304.950 121.950 307.050 124.050 ;
        RECT 308.100 123.150 309.900 123.900 ;
        RECT 310.950 121.950 313.050 124.050 ;
        RECT 314.100 123.150 315.900 123.900 ;
        RECT 323.100 123.150 324.900 123.900 ;
        RECT 329.100 123.150 330.900 123.900 ;
        RECT 332.400 121.650 333.300 126.900 ;
        RECT 305.400 117.600 306.300 120.900 ;
        RECT 329.100 120.000 333.300 121.650 ;
        RECT 232.800 111.600 234.600 114.600 ;
        RECT 248.400 111.600 250.200 114.600 ;
        RECT 268.800 111.600 270.600 114.600 ;
        RECT 284.400 111.600 286.200 114.600 ;
        RECT 290.400 111.600 292.200 117.600 ;
        RECT 305.400 115.950 310.800 117.600 ;
        RECT 309.000 111.600 310.800 115.950 ;
        RECT 329.100 111.600 330.900 120.000 ;
        RECT 338.550 118.050 339.450 128.550 ;
        RECT 344.100 125.100 345.900 125.850 ;
        RECT 343.950 121.950 346.050 124.050 ;
        RECT 347.400 120.300 348.450 137.400 ;
        RECT 354.000 131.400 355.800 143.400 ;
        RECT 367.800 137.400 369.600 143.400 ;
        RECT 349.950 124.950 352.050 127.050 ;
        RECT 354.000 125.100 355.050 131.400 ;
        RECT 361.950 130.950 364.050 133.050 ;
        RECT 362.550 126.450 363.450 130.950 ;
        RECT 368.400 128.100 369.600 137.400 ;
        RECT 385.500 131.400 387.300 143.400 ;
        RECT 406.500 131.400 408.300 143.400 ;
        RECT 427.800 137.400 429.600 143.400 ;
        RECT 385.950 128.100 387.150 131.400 ;
        RECT 406.950 128.100 408.150 131.400 ;
        RECT 367.950 126.450 370.050 127.050 ;
        RECT 362.550 125.550 370.050 126.450 ;
        RECT 367.950 124.950 370.050 125.550 ;
        RECT 380.100 125.100 381.900 125.850 ;
        RECT 382.950 124.950 385.050 127.050 ;
        RECT 386.100 125.100 387.150 128.100 ;
        RECT 401.100 125.100 402.900 125.850 ;
        RECT 403.950 124.950 406.050 127.050 ;
        RECT 407.100 125.100 408.150 128.100 ;
        RECT 424.950 127.950 427.050 130.050 ;
        RECT 428.400 128.100 429.600 137.400 ;
        RECT 440.400 132.300 442.200 143.400 ;
        RECT 446.400 132.300 448.200 143.400 ;
        RECT 440.400 131.400 448.200 132.300 ;
        RECT 449.400 131.400 451.200 143.400 ;
        RECT 454.950 139.950 457.050 142.050 ;
        RECT 430.950 127.950 433.050 130.050 ;
        RECT 409.950 124.950 412.050 127.050 ;
        RECT 425.100 126.150 426.900 126.900 ;
        RECT 427.950 124.950 430.050 127.050 ;
        RECT 431.100 126.150 432.900 126.900 ;
        RECT 439.950 124.950 442.050 127.050 ;
        RECT 443.100 125.100 444.900 125.850 ;
        RECT 445.950 124.950 448.050 130.050 ;
        RECT 449.700 125.100 450.600 131.400 ;
        RECT 350.100 123.150 351.900 123.900 ;
        RECT 352.950 121.950 355.050 124.050 ;
        RECT 344.400 119.100 351.900 120.300 ;
        RECT 337.950 115.950 340.050 118.050 ;
        RECT 344.400 111.600 346.200 119.100 ;
        RECT 350.100 118.500 351.900 119.100 ;
        RECT 352.950 117.600 353.850 120.900 ;
        RECT 351.900 115.800 353.850 117.600 ;
        RECT 351.900 111.600 353.700 115.800 ;
        RECT 368.400 114.600 369.600 123.900 ;
        RECT 371.100 122.100 372.900 122.850 ;
        RECT 379.950 121.950 382.050 124.050 ;
        RECT 383.100 123.150 384.900 123.900 ;
        RECT 385.950 121.950 388.050 124.050 ;
        RECT 389.100 123.150 390.900 123.900 ;
        RECT 400.950 121.950 403.050 124.050 ;
        RECT 404.100 123.150 405.900 123.900 ;
        RECT 406.950 121.950 409.050 124.050 ;
        RECT 410.100 123.150 411.900 123.900 ;
        RECT 370.950 115.950 373.050 121.050 ;
        RECT 386.850 120.750 388.050 120.900 ;
        RECT 407.850 120.750 409.050 120.900 ;
        RECT 386.850 119.700 390.600 120.750 ;
        RECT 407.850 119.700 411.600 120.750 ;
        RECT 428.400 119.700 429.600 123.900 ;
        RECT 440.100 123.150 441.900 123.900 ;
        RECT 380.400 116.700 388.200 118.050 ;
        RECT 367.800 111.600 369.600 114.600 ;
        RECT 380.400 111.600 382.200 116.700 ;
        RECT 386.400 111.600 388.200 116.700 ;
        RECT 389.400 117.600 390.600 119.700 ;
        RECT 389.400 111.600 391.200 117.600 ;
        RECT 401.400 116.700 409.200 118.050 ;
        RECT 401.400 111.600 403.200 116.700 ;
        RECT 407.400 111.600 409.200 116.700 ;
        RECT 410.400 117.600 411.600 119.700 ;
        RECT 426.000 118.800 429.600 119.700 ;
        RECT 442.950 118.950 445.050 124.050 ;
        RECT 446.100 123.150 447.900 123.900 ;
        RECT 448.950 123.450 451.050 124.050 ;
        RECT 455.550 123.450 456.450 139.950 ;
        RECT 464.400 137.400 466.200 143.400 ;
        RECT 464.700 137.100 466.200 137.400 ;
        RECT 470.400 137.400 472.200 143.400 ;
        RECT 470.400 137.100 471.300 137.400 ;
        RECT 464.700 136.200 471.300 137.100 ;
        RECT 464.100 131.100 465.900 131.850 ;
        RECT 470.400 131.100 471.300 136.200 ;
        RECT 487.800 131.400 489.600 143.400 ;
        RECT 500.400 132.300 502.200 143.400 ;
        RECT 506.400 132.300 508.200 143.400 ;
        RECT 500.400 131.400 508.200 132.300 ;
        RECT 509.400 131.400 511.200 143.400 ;
        RECT 523.800 131.400 525.600 143.400 ;
        RECT 526.800 132.300 528.600 143.400 ;
        RECT 532.800 132.300 534.600 143.400 ;
        RECT 544.800 137.400 546.600 143.400 ;
        RECT 526.800 131.400 534.600 132.300 ;
        RECT 463.800 127.950 466.050 130.050 ;
        RECT 469.950 129.450 472.050 130.050 ;
        RECT 469.950 128.550 477.450 129.450 ;
        RECT 469.950 127.950 472.050 128.550 ;
        RECT 460.950 124.950 463.050 127.050 ;
        RECT 466.950 124.950 469.050 127.050 ;
        RECT 448.950 122.550 456.450 123.450 ;
        RECT 461.100 123.150 462.900 123.900 ;
        RECT 467.100 123.150 468.900 123.900 ;
        RECT 448.950 121.950 451.050 122.550 ;
        RECT 470.400 121.650 471.300 126.900 ;
        RECT 410.400 111.600 412.200 117.600 ;
        RECT 426.000 111.600 427.800 118.800 ;
        RECT 449.700 117.600 450.600 120.900 ;
        RECT 445.200 115.950 450.600 117.600 ;
        RECT 467.100 120.000 471.300 121.650 ;
        RECT 445.200 111.600 447.000 115.950 ;
        RECT 467.100 111.600 468.900 120.000 ;
        RECT 476.550 115.050 477.450 128.550 ;
        RECT 487.950 128.100 489.300 131.400 ;
        RECT 484.950 124.950 487.050 127.050 ;
        RECT 488.100 123.900 489.300 128.100 ;
        RECT 499.950 124.950 502.050 127.050 ;
        RECT 503.100 125.100 504.900 125.850 ;
        RECT 505.950 124.950 508.050 127.050 ;
        RECT 509.700 125.100 510.600 131.400 ;
        RECT 517.950 124.950 520.050 127.050 ;
        RECT 524.400 125.100 525.300 131.400 ;
        RECT 538.950 127.950 541.050 130.050 ;
        RECT 545.400 128.100 546.600 137.400 ;
        RECT 560.400 137.400 562.200 143.400 ;
        RECT 560.400 128.100 561.600 137.400 ;
        RECT 580.500 131.400 582.300 143.400 ;
        RECT 601.800 137.400 603.600 143.400 ;
        RECT 619.800 137.400 621.600 143.400 ;
        RECT 562.950 127.950 565.050 130.050 ;
        RECT 580.950 128.100 582.150 131.400 ;
        RECT 526.950 124.950 529.200 127.050 ;
        RECT 530.100 125.100 531.900 125.850 ;
        RECT 532.950 124.950 535.050 127.050 ;
        RECT 487.950 117.600 489.300 123.900 ;
        RECT 491.100 123.150 492.900 123.900 ;
        RECT 500.100 123.150 501.900 123.900 ;
        RECT 502.950 121.950 505.050 124.050 ;
        RECT 506.100 123.150 507.900 123.900 ;
        RECT 508.950 121.950 514.050 124.050 ;
        RECT 509.700 117.600 510.600 120.900 ;
        RECT 475.950 112.950 478.050 115.050 ;
        RECT 487.800 111.600 489.600 117.600 ;
        RECT 505.200 115.950 510.600 117.600 ;
        RECT 505.200 111.600 507.000 115.950 ;
        RECT 518.550 115.050 519.450 124.950 ;
        RECT 523.950 121.950 526.050 124.050 ;
        RECT 527.100 123.150 528.900 123.900 ;
        RECT 529.950 121.950 532.200 124.050 ;
        RECT 533.100 123.150 534.900 123.900 ;
        RECT 524.400 117.600 525.300 120.900 ;
        RECT 524.400 115.950 529.800 117.600 ;
        RECT 518.550 113.550 523.050 115.050 ;
        RECT 519.000 112.950 523.050 113.550 ;
        RECT 528.000 111.600 529.800 115.950 ;
        RECT 539.550 115.050 540.450 127.950 ;
        RECT 542.100 124.950 547.050 127.050 ;
        RECT 557.100 126.150 558.900 126.900 ;
        RECT 559.950 124.950 562.050 127.050 ;
        RECT 563.100 126.150 564.900 126.900 ;
        RECT 575.100 125.100 576.900 125.850 ;
        RECT 577.950 124.950 580.050 127.050 ;
        RECT 581.100 125.100 582.150 128.100 ;
        RECT 598.950 127.950 601.050 130.050 ;
        RECT 602.400 128.100 603.600 137.400 ;
        RECT 604.950 127.950 607.050 130.050 ;
        RECT 616.950 127.950 619.050 130.050 ;
        RECT 620.400 128.100 621.600 137.400 ;
        RECT 632.400 132.300 634.200 143.400 ;
        RECT 638.400 132.300 640.200 143.400 ;
        RECT 632.400 131.400 640.200 132.300 ;
        RECT 641.400 131.400 643.200 143.400 ;
        RECT 655.800 137.400 657.600 143.400 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 622.950 127.950 625.050 130.050 ;
        RECT 583.950 124.950 586.050 127.050 ;
        RECT 599.100 126.150 600.900 126.900 ;
        RECT 601.950 124.950 604.050 127.050 ;
        RECT 605.100 126.150 606.900 126.900 ;
        RECT 617.100 126.150 618.900 126.900 ;
        RECT 619.950 124.950 622.050 127.050 ;
        RECT 623.100 126.150 624.900 126.900 ;
        RECT 631.800 124.950 634.050 127.050 ;
        RECT 635.100 125.100 636.900 125.850 ;
        RECT 637.950 124.950 640.200 127.050 ;
        RECT 641.700 125.100 642.600 131.400 ;
        RECT 538.950 112.950 541.050 115.050 ;
        RECT 545.400 114.600 546.600 123.900 ;
        RECT 548.100 122.100 549.900 122.850 ;
        RECT 547.950 118.950 553.050 121.050 ;
        RECT 560.400 119.700 561.600 123.900 ;
        RECT 574.950 121.950 577.050 124.050 ;
        RECT 578.100 123.150 579.900 123.900 ;
        RECT 580.950 121.950 583.050 124.050 ;
        RECT 584.100 123.150 585.900 123.900 ;
        RECT 581.850 120.750 583.050 120.900 ;
        RECT 581.850 119.700 585.600 120.750 ;
        RECT 602.400 119.700 603.600 123.900 ;
        RECT 620.400 119.700 621.600 123.900 ;
        RECT 632.100 123.150 633.900 123.900 ;
        RECT 634.950 121.950 637.050 124.050 ;
        RECT 638.100 123.150 639.900 123.900 ;
        RECT 640.950 121.950 643.050 124.050 ;
        RECT 647.550 121.050 648.450 133.950 ;
        RECT 656.400 128.100 657.600 137.400 ;
        RECT 664.950 133.950 667.050 136.050 ;
        RECT 655.950 126.450 658.050 127.050 ;
        RECT 660.000 126.450 664.050 127.050 ;
        RECT 655.950 125.550 664.050 126.450 ;
        RECT 655.950 124.950 658.050 125.550 ;
        RECT 660.000 124.950 664.050 125.550 ;
        RECT 560.400 118.800 564.000 119.700 ;
        RECT 544.800 111.600 546.600 114.600 ;
        RECT 562.200 111.600 564.000 118.800 ;
        RECT 575.400 116.700 583.200 118.050 ;
        RECT 575.400 111.600 577.200 116.700 ;
        RECT 581.400 111.600 583.200 116.700 ;
        RECT 584.400 117.600 585.600 119.700 ;
        RECT 600.000 118.800 603.600 119.700 ;
        RECT 618.000 118.800 621.600 119.700 ;
        RECT 584.400 111.600 586.200 117.600 ;
        RECT 600.000 111.600 601.800 118.800 ;
        RECT 618.000 111.600 619.800 118.800 ;
        RECT 641.700 117.600 642.600 120.900 ;
        RECT 646.950 118.950 649.050 121.050 ;
        RECT 637.200 115.950 642.600 117.600 ;
        RECT 637.200 111.600 639.000 115.950 ;
        RECT 656.400 114.600 657.600 123.900 ;
        RECT 659.100 122.100 660.900 122.850 ;
        RECT 665.550 121.050 666.450 133.950 ;
        RECT 674.700 131.400 676.500 143.400 ;
        RECT 691.200 131.400 693.000 143.400 ;
        RECT 697.800 137.400 699.600 143.400 ;
        RECT 712.800 137.400 714.600 143.400 ;
        RECT 674.850 128.100 676.050 131.400 ;
        RECT 670.800 124.950 673.050 127.050 ;
        RECT 674.850 125.100 675.900 128.100 ;
        RECT 676.950 124.950 679.050 127.050 ;
        RECT 680.100 125.100 681.900 125.850 ;
        RECT 691.950 125.100 693.000 131.400 ;
        RECT 694.950 124.950 697.050 127.050 ;
        RECT 671.100 123.150 672.900 123.900 ;
        RECT 673.950 121.950 676.050 124.050 ;
        RECT 677.100 123.150 678.900 123.900 ;
        RECT 679.950 121.950 682.050 124.050 ;
        RECT 691.950 123.450 694.050 124.050 ;
        RECT 686.550 122.550 694.050 123.450 ;
        RECT 695.100 123.150 696.900 123.900 ;
        RECT 658.950 118.950 661.050 121.050 ;
        RECT 665.100 118.950 667.200 121.050 ;
        RECT 673.950 120.750 675.150 120.900 ;
        RECT 671.400 119.700 675.150 120.750 ;
        RECT 671.400 117.600 672.600 119.700 ;
        RECT 655.800 111.600 657.600 114.600 ;
        RECT 670.800 111.600 672.600 117.600 ;
        RECT 673.800 116.700 681.600 118.050 ;
        RECT 673.800 111.600 675.600 116.700 ;
        RECT 679.800 111.600 681.600 116.700 ;
        RECT 686.550 115.050 687.450 122.550 ;
        RECT 691.950 121.950 694.050 122.550 ;
        RECT 693.150 117.600 694.050 120.900 ;
        RECT 698.550 120.300 699.600 137.400 ;
        RECT 713.700 137.100 714.600 137.400 ;
        RECT 718.800 137.400 720.600 143.400 ;
        RECT 733.800 137.400 735.600 143.400 ;
        RECT 748.800 137.400 750.600 143.400 ;
        RECT 757.950 139.950 760.050 142.050 ;
        RECT 718.800 137.100 720.300 137.400 ;
        RECT 713.700 136.200 720.300 137.100 ;
        RECT 706.950 133.950 709.050 136.050 ;
        RECT 701.100 125.100 702.900 125.850 ;
        RECT 700.950 121.950 703.050 124.050 ;
        RECT 695.100 119.100 702.600 120.300 ;
        RECT 695.100 118.500 696.900 119.100 ;
        RECT 693.150 115.800 695.100 117.600 ;
        RECT 685.950 112.950 688.050 115.050 ;
        RECT 693.300 111.600 695.100 115.800 ;
        RECT 700.800 111.600 702.600 119.100 ;
        RECT 707.550 115.050 708.450 133.950 ;
        RECT 713.700 131.100 714.600 136.200 ;
        RECT 727.800 133.950 729.900 136.050 ;
        RECT 719.100 131.100 720.900 131.850 ;
        RECT 709.950 127.950 715.050 130.050 ;
        RECT 718.950 127.950 721.050 130.050 ;
        RECT 713.700 121.650 714.600 126.900 ;
        RECT 715.950 124.950 718.050 127.050 ;
        RECT 721.950 124.950 724.200 127.050 ;
        RECT 728.550 126.450 729.450 133.950 ;
        RECT 734.400 128.100 735.600 137.400 ;
        RECT 749.400 128.100 750.600 137.400 ;
        RECT 733.950 126.450 736.050 127.050 ;
        RECT 728.550 125.550 736.050 126.450 ;
        RECT 733.950 124.950 736.050 125.550 ;
        RECT 748.950 124.950 754.200 127.050 ;
        RECT 758.550 124.050 759.450 139.950 ;
        RECT 767.700 131.400 769.500 143.400 ;
        RECT 787.800 137.400 789.600 143.400 ;
        RECT 767.850 128.100 769.050 131.400 ;
        RECT 763.950 124.950 766.050 127.050 ;
        RECT 767.850 125.100 768.900 128.100 ;
        RECT 778.950 127.950 781.050 130.050 ;
        RECT 784.950 127.950 787.050 130.050 ;
        RECT 788.400 128.100 789.600 137.400 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 790.950 127.950 793.050 130.050 ;
        RECT 769.950 124.950 772.050 127.050 ;
        RECT 773.100 125.100 774.900 125.850 ;
        RECT 716.100 123.150 717.900 123.900 ;
        RECT 722.100 123.150 723.900 123.900 ;
        RECT 713.700 120.000 717.900 121.650 ;
        RECT 706.950 112.950 709.050 115.050 ;
        RECT 716.100 111.600 717.900 120.000 ;
        RECT 734.400 114.600 735.600 123.900 ;
        RECT 737.100 122.100 738.900 122.850 ;
        RECT 736.950 118.950 739.050 121.050 ;
        RECT 749.400 114.600 750.600 123.900 ;
        RECT 752.100 122.100 753.900 122.850 ;
        RECT 757.950 121.950 760.050 124.050 ;
        RECT 764.100 123.150 765.900 123.900 ;
        RECT 766.950 121.950 769.050 124.050 ;
        RECT 770.100 123.150 771.900 123.900 ;
        RECT 772.950 121.950 775.050 124.050 ;
        RECT 779.550 121.050 780.450 127.950 ;
        RECT 785.100 126.150 786.900 126.900 ;
        RECT 787.950 124.950 790.050 127.050 ;
        RECT 791.100 126.150 792.900 126.900 ;
        RECT 751.950 118.950 754.050 121.050 ;
        RECT 766.950 120.750 768.150 120.900 ;
        RECT 764.400 119.700 768.150 120.750 ;
        RECT 764.400 117.600 765.600 119.700 ;
        RECT 778.950 118.950 781.050 121.050 ;
        RECT 788.400 119.700 789.600 123.900 ;
        RECT 786.000 118.800 789.600 119.700 ;
        RECT 733.800 111.600 735.600 114.600 ;
        RECT 748.800 111.600 750.600 114.600 ;
        RECT 763.800 111.600 765.600 117.600 ;
        RECT 766.800 116.700 774.600 118.050 ;
        RECT 766.800 111.600 768.600 116.700 ;
        RECT 772.800 111.600 774.600 116.700 ;
        RECT 786.000 111.600 787.800 118.800 ;
        RECT 797.550 115.050 798.450 133.950 ;
        RECT 806.700 131.400 808.500 143.400 ;
        RECT 817.950 139.950 820.050 142.050 ;
        RECT 806.850 128.100 808.050 131.400 ;
        RECT 802.950 124.950 805.050 127.050 ;
        RECT 806.850 125.100 807.900 128.100 ;
        RECT 808.950 124.950 811.050 127.050 ;
        RECT 812.100 125.100 813.900 125.850 ;
        RECT 803.100 123.150 804.900 123.900 ;
        RECT 805.800 121.950 808.050 124.050 ;
        RECT 809.100 123.150 810.900 123.900 ;
        RECT 811.800 121.950 814.050 124.050 ;
        RECT 805.950 120.750 807.150 120.900 ;
        RECT 803.400 119.700 807.150 120.750 ;
        RECT 803.400 117.600 804.600 119.700 ;
        RECT 796.950 112.950 799.050 115.050 ;
        RECT 802.800 111.600 804.600 117.600 ;
        RECT 805.800 116.700 813.600 118.050 ;
        RECT 805.800 111.600 807.600 116.700 ;
        RECT 811.800 111.600 813.600 116.700 ;
        RECT 818.550 115.050 819.450 139.950 ;
        RECT 827.700 131.400 829.500 143.400 ;
        RECT 847.500 131.400 849.300 143.400 ;
        RECT 827.850 128.100 829.050 131.400 ;
        RECT 847.950 128.100 849.150 131.400 ;
        RECT 850.950 129.000 853.050 133.050 ;
        RECT 823.950 124.950 826.050 127.050 ;
        RECT 827.850 125.100 828.900 128.100 ;
        RECT 829.950 124.950 832.050 127.050 ;
        RECT 833.100 125.100 834.900 125.850 ;
        RECT 842.100 125.100 843.900 125.850 ;
        RECT 844.950 124.950 847.050 127.050 ;
        RECT 848.100 125.100 849.150 128.100 ;
        RECT 851.550 127.050 852.450 129.000 ;
        RECT 850.950 124.950 853.050 127.050 ;
        RECT 824.100 123.150 825.900 123.900 ;
        RECT 826.800 121.950 829.050 124.050 ;
        RECT 830.100 123.150 831.900 123.900 ;
        RECT 832.950 121.950 835.050 124.050 ;
        RECT 841.950 121.950 844.050 124.050 ;
        RECT 845.100 123.150 846.900 123.900 ;
        RECT 847.950 121.950 850.200 124.050 ;
        RECT 851.100 123.150 852.900 123.900 ;
        RECT 826.950 120.750 828.150 120.900 ;
        RECT 824.400 119.700 828.150 120.750 ;
        RECT 848.850 120.750 850.050 120.900 ;
        RECT 848.850 119.700 852.600 120.750 ;
        RECT 824.400 117.600 825.600 119.700 ;
        RECT 817.950 112.950 820.050 115.050 ;
        RECT 823.800 111.600 825.600 117.600 ;
        RECT 826.800 116.700 834.600 118.050 ;
        RECT 826.800 111.600 828.600 116.700 ;
        RECT 832.800 111.600 834.600 116.700 ;
        RECT 842.400 116.700 850.200 118.050 ;
        RECT 842.400 111.600 844.200 116.700 ;
        RECT 848.400 111.600 850.200 116.700 ;
        RECT 851.400 117.600 852.600 119.700 ;
        RECT 851.400 111.600 853.200 117.600 ;
        RECT 10.800 104.400 12.600 107.400 ;
        RECT 11.400 95.100 12.600 104.400 ;
        RECT 25.800 101.400 27.600 107.400 ;
        RECT 13.950 97.950 16.050 100.050 ;
        RECT 26.400 99.300 27.600 101.400 ;
        RECT 28.800 102.300 30.600 107.400 ;
        RECT 34.800 102.300 36.600 107.400 ;
        RECT 28.800 100.950 36.600 102.300 ;
        RECT 26.400 98.250 30.150 99.300 ;
        RECT 50.100 99.000 51.900 107.400 ;
        RECT 70.200 103.050 72.000 107.400 ;
        RECT 93.000 103.050 94.800 107.400 ;
        RECT 70.200 101.400 75.600 103.050 ;
        RECT 28.950 98.100 30.150 98.250 ;
        RECT 47.700 97.350 51.900 99.000 ;
        RECT 74.700 98.100 75.600 101.400 ;
        RECT 82.950 100.950 85.050 103.050 ;
        RECT 89.400 101.400 94.800 103.050 ;
        RECT 14.100 96.150 15.900 96.900 ;
        RECT 26.100 95.100 27.900 95.850 ;
        RECT 28.950 94.950 31.050 97.050 ;
        RECT 32.100 95.100 33.900 95.850 ;
        RECT 34.950 94.950 37.050 97.050 ;
        RECT 10.950 91.950 16.050 94.050 ;
        RECT 25.950 91.950 28.050 94.050 ;
        RECT 29.850 90.900 30.900 93.900 ;
        RECT 31.950 91.950 34.050 94.050 ;
        RECT 35.100 93.150 36.900 93.900 ;
        RECT 47.700 92.100 48.600 97.350 ;
        RECT 50.100 95.100 51.900 95.850 ;
        RECT 56.100 95.100 57.900 95.850 ;
        RECT 65.100 95.100 66.900 95.850 ;
        RECT 67.950 94.950 70.050 97.050 ;
        RECT 71.100 95.100 72.900 95.850 ;
        RECT 73.950 94.950 79.050 97.050 ;
        RECT 83.550 96.450 84.450 100.950 ;
        RECT 89.400 98.100 90.300 101.400 ;
        RECT 113.100 99.000 114.900 107.400 ;
        RECT 134.100 99.000 135.900 107.400 ;
        RECT 151.800 101.400 153.600 107.400 ;
        RECT 110.700 97.350 114.900 99.000 ;
        RECT 131.700 97.350 135.900 99.000 ;
        RECT 152.400 99.300 153.600 101.400 ;
        RECT 154.800 102.300 156.600 107.400 ;
        RECT 160.800 102.300 162.600 107.400 ;
        RECT 154.800 100.950 162.600 102.300 ;
        RECT 170.400 102.300 172.200 107.400 ;
        RECT 176.400 102.300 178.200 107.400 ;
        RECT 170.400 100.950 178.200 102.300 ;
        RECT 179.400 101.400 181.200 107.400 ;
        RECT 193.800 101.400 195.600 107.400 ;
        RECT 179.400 99.300 180.600 101.400 ;
        RECT 152.400 98.250 156.150 99.300 ;
        RECT 154.950 98.100 156.150 98.250 ;
        RECT 176.850 98.250 180.600 99.300 ;
        RECT 176.850 98.100 178.050 98.250 ;
        RECT 184.950 97.950 187.050 100.050 ;
        RECT 194.400 99.300 195.600 101.400 ;
        RECT 196.800 102.300 198.600 107.400 ;
        RECT 202.800 102.300 204.600 107.400 ;
        RECT 196.800 100.950 204.600 102.300 ;
        RECT 208.950 100.950 211.050 103.050 ;
        RECT 194.400 98.250 198.150 99.300 ;
        RECT 196.950 98.100 198.150 98.250 ;
        RECT 88.950 96.450 91.050 97.050 ;
        RECT 83.550 95.550 91.050 96.450 ;
        RECT 88.950 94.950 91.050 95.550 ;
        RECT 92.100 95.100 93.900 95.850 ;
        RECT 94.950 94.950 97.050 97.050 ;
        RECT 98.100 95.100 99.900 95.850 ;
        RECT 49.950 91.950 52.050 94.050 ;
        RECT 55.950 91.950 58.200 94.050 ;
        RECT 64.950 91.950 67.050 94.050 ;
        RECT 68.100 93.150 69.900 93.900 ;
        RECT 70.950 91.950 73.050 94.050 ;
        RECT 11.400 81.600 12.600 90.900 ;
        RECT 29.850 87.600 31.050 90.900 ;
        RECT 46.950 88.950 49.050 91.050 ;
        RECT 52.950 88.950 55.050 91.050 ;
        RECT 10.800 75.600 12.600 81.600 ;
        RECT 29.700 75.600 31.500 87.600 ;
        RECT 47.700 82.800 48.600 87.900 ;
        RECT 53.100 87.150 54.900 87.900 ;
        RECT 74.700 87.600 75.600 93.900 ;
        RECT 89.400 87.600 90.300 93.900 ;
        RECT 91.800 91.950 94.050 94.050 ;
        RECT 95.100 93.150 96.900 93.900 ;
        RECT 97.950 91.950 100.050 94.050 ;
        RECT 110.700 92.100 111.600 97.350 ;
        RECT 113.100 95.100 114.900 95.850 ;
        RECT 119.100 95.100 120.900 95.850 ;
        RECT 112.950 91.950 115.050 94.050 ;
        RECT 118.950 91.950 121.050 94.050 ;
        RECT 131.700 92.100 132.600 97.350 ;
        RECT 134.100 95.100 135.900 95.850 ;
        RECT 140.100 95.100 141.900 95.850 ;
        RECT 152.100 95.100 153.900 95.850 ;
        RECT 154.950 94.950 157.050 97.050 ;
        RECT 158.100 95.100 159.900 95.850 ;
        RECT 160.950 94.950 163.050 97.050 ;
        RECT 169.950 94.950 172.050 97.050 ;
        RECT 173.100 95.100 174.900 95.850 ;
        RECT 175.950 94.950 178.050 97.050 ;
        RECT 179.100 95.100 180.900 95.850 ;
        RECT 133.950 91.950 136.050 94.050 ;
        RECT 139.950 91.950 142.050 94.050 ;
        RECT 145.800 91.950 147.900 94.050 ;
        RECT 151.950 91.950 154.050 94.050 ;
        RECT 106.950 88.950 112.050 91.050 ;
        RECT 115.950 88.950 118.050 91.050 ;
        RECT 130.950 90.450 133.050 91.050 ;
        RECT 125.550 89.550 133.050 90.450 ;
        RECT 65.400 86.700 73.200 87.600 ;
        RECT 47.700 81.900 54.300 82.800 ;
        RECT 47.700 81.600 48.600 81.900 ;
        RECT 46.800 75.600 48.600 81.600 ;
        RECT 52.800 81.600 54.300 81.900 ;
        RECT 52.800 75.600 54.600 81.600 ;
        RECT 65.400 75.600 67.200 86.700 ;
        RECT 71.400 75.600 73.200 86.700 ;
        RECT 74.400 75.600 76.200 87.600 ;
        RECT 88.800 75.600 90.600 87.600 ;
        RECT 91.800 86.700 99.600 87.600 ;
        RECT 91.800 75.600 93.600 86.700 ;
        RECT 97.800 75.600 99.600 86.700 ;
        RECT 110.700 82.800 111.600 87.900 ;
        RECT 116.100 87.150 117.900 87.900 ;
        RECT 125.550 85.050 126.450 89.550 ;
        RECT 130.950 88.950 133.050 89.550 ;
        RECT 136.950 88.950 139.050 91.050 ;
        RECT 146.550 88.050 147.450 91.950 ;
        RECT 155.850 90.900 156.900 93.900 ;
        RECT 157.950 91.950 160.050 94.050 ;
        RECT 161.100 93.150 162.900 93.900 ;
        RECT 170.100 93.150 171.900 93.900 ;
        RECT 172.950 91.950 175.050 94.050 ;
        RECT 176.100 90.900 177.150 93.900 ;
        RECT 178.950 91.950 181.200 94.050 ;
        RECT 124.950 82.950 127.050 85.050 ;
        RECT 131.700 82.800 132.600 87.900 ;
        RECT 137.100 87.150 138.900 87.900 ;
        RECT 145.950 85.950 148.050 88.050 ;
        RECT 155.850 87.600 157.050 90.900 ;
        RECT 175.950 87.600 177.150 90.900 ;
        RECT 179.550 90.000 180.450 91.950 ;
        RECT 110.700 81.900 117.300 82.800 ;
        RECT 110.700 81.600 111.600 81.900 ;
        RECT 109.800 75.600 111.600 81.600 ;
        RECT 115.800 81.600 117.300 81.900 ;
        RECT 131.700 81.900 138.300 82.800 ;
        RECT 131.700 81.600 132.600 81.900 ;
        RECT 115.800 75.600 117.600 81.600 ;
        RECT 130.800 75.600 132.600 81.600 ;
        RECT 136.800 81.600 138.300 81.900 ;
        RECT 136.800 75.600 138.600 81.600 ;
        RECT 155.700 75.600 157.500 87.600 ;
        RECT 175.500 75.600 177.300 87.600 ;
        RECT 178.950 85.950 181.050 90.000 ;
        RECT 185.550 79.050 186.450 97.950 ;
        RECT 194.100 95.100 195.900 95.850 ;
        RECT 196.950 94.950 199.050 97.050 ;
        RECT 200.100 95.100 201.900 95.850 ;
        RECT 202.950 94.950 205.050 97.050 ;
        RECT 209.550 94.050 210.450 100.950 ;
        RECT 218.100 99.000 219.900 107.400 ;
        RECT 240.000 103.050 241.800 107.400 ;
        RECT 215.700 97.350 219.900 99.000 ;
        RECT 236.400 101.400 241.800 103.050 ;
        RECT 256.800 101.400 258.600 107.400 ;
        RECT 236.400 98.100 237.300 101.400 ;
        RECT 250.950 97.950 253.050 100.050 ;
        RECT 257.400 99.300 258.600 101.400 ;
        RECT 259.800 102.300 261.600 107.400 ;
        RECT 265.800 102.300 267.600 107.400 ;
        RECT 259.800 100.950 267.600 102.300 ;
        RECT 278.400 104.400 280.200 107.400 ;
        RECT 257.400 98.250 261.150 99.300 ;
        RECT 259.950 98.100 261.150 98.250 ;
        RECT 274.950 97.950 277.050 100.050 ;
        RECT 193.950 91.950 196.050 94.050 ;
        RECT 197.850 90.900 198.900 93.900 ;
        RECT 199.950 91.950 202.050 94.050 ;
        RECT 203.100 93.150 204.900 93.900 ;
        RECT 208.950 91.950 211.050 94.050 ;
        RECT 215.700 92.100 216.600 97.350 ;
        RECT 229.950 96.450 234.000 97.050 ;
        RECT 235.950 96.450 238.050 97.050 ;
        RECT 218.100 95.100 219.900 95.850 ;
        RECT 224.100 95.100 225.900 95.850 ;
        RECT 229.950 95.550 238.050 96.450 ;
        RECT 229.950 94.950 234.000 95.550 ;
        RECT 235.950 94.950 238.050 95.550 ;
        RECT 239.100 95.100 240.900 95.850 ;
        RECT 241.950 94.950 244.200 97.050 ;
        RECT 245.100 95.100 246.900 95.850 ;
        RECT 217.950 91.950 220.050 94.050 ;
        RECT 223.950 91.950 226.050 94.050 ;
        RECT 197.850 87.600 199.050 90.900 ;
        RECT 214.950 90.450 217.050 91.050 ;
        RECT 209.550 89.550 217.050 90.450 ;
        RECT 184.950 76.950 187.050 79.050 ;
        RECT 197.700 75.600 199.500 87.600 ;
        RECT 209.550 85.050 210.450 89.550 ;
        RECT 214.950 88.950 217.050 89.550 ;
        RECT 220.950 88.950 223.050 91.050 ;
        RECT 208.950 82.950 211.050 85.050 ;
        RECT 215.700 82.800 216.600 87.900 ;
        RECT 221.100 87.150 222.900 87.900 ;
        RECT 236.400 87.600 237.300 93.900 ;
        RECT 238.950 91.950 241.050 94.050 ;
        RECT 242.100 93.150 243.900 93.900 ;
        RECT 244.950 91.950 247.050 94.050 ;
        RECT 251.550 91.050 252.450 97.950 ;
        RECT 257.100 95.100 258.900 95.850 ;
        RECT 259.950 94.950 262.050 97.050 ;
        RECT 263.100 95.100 264.900 95.850 ;
        RECT 265.950 94.950 268.200 97.050 ;
        RECT 275.100 96.150 276.900 96.900 ;
        RECT 278.400 95.100 279.600 104.400 ;
        RECT 296.100 99.000 297.900 107.400 ;
        RECT 317.100 99.000 318.900 107.400 ;
        RECT 337.200 103.050 339.000 107.400 ;
        RECT 337.200 101.400 342.600 103.050 ;
        RECT 355.800 101.400 357.600 107.400 ;
        RECT 296.100 97.350 300.300 99.000 ;
        RECT 290.100 95.100 291.900 95.850 ;
        RECT 296.100 95.100 297.900 95.850 ;
        RECT 256.950 91.950 259.050 94.050 ;
        RECT 250.950 88.950 253.050 91.050 ;
        RECT 260.850 90.900 261.900 93.900 ;
        RECT 262.950 91.950 265.050 94.050 ;
        RECT 266.100 93.150 267.900 93.900 ;
        RECT 277.950 91.950 283.050 94.050 ;
        RECT 289.950 91.950 292.050 94.050 ;
        RECT 295.950 91.950 298.050 94.050 ;
        RECT 299.400 92.100 300.300 97.350 ;
        RECT 314.700 97.350 318.900 99.000 ;
        RECT 341.700 98.100 342.600 101.400 ;
        RECT 356.400 99.300 357.600 101.400 ;
        RECT 358.800 102.300 360.600 107.400 ;
        RECT 364.800 102.300 366.600 107.400 ;
        RECT 358.800 100.950 366.600 102.300 ;
        RECT 377.400 104.400 379.200 107.400 ;
        RECT 356.400 98.250 360.150 99.300 ;
        RECT 358.950 98.100 360.150 98.250 ;
        RECT 370.950 97.950 376.050 100.050 ;
        RECT 314.700 92.100 315.600 97.350 ;
        RECT 317.100 95.100 318.900 95.850 ;
        RECT 323.100 95.100 324.900 95.850 ;
        RECT 332.100 95.100 333.900 95.850 ;
        RECT 334.950 94.950 337.050 97.050 ;
        RECT 338.100 95.100 339.900 95.850 ;
        RECT 340.950 94.950 343.050 97.050 ;
        RECT 356.100 95.100 357.900 95.850 ;
        RECT 358.800 94.950 361.050 97.050 ;
        RECT 362.100 95.100 363.900 95.850 ;
        RECT 364.950 94.950 367.050 97.050 ;
        RECT 374.100 96.150 375.900 96.900 ;
        RECT 377.400 95.100 378.600 104.400 ;
        RECT 391.800 101.400 393.600 107.400 ;
        RECT 392.400 99.300 393.600 101.400 ;
        RECT 394.800 102.300 396.600 107.400 ;
        RECT 400.800 102.300 402.600 107.400 ;
        RECT 394.800 100.950 402.600 102.300 ;
        RECT 410.400 102.300 412.200 107.400 ;
        RECT 416.400 102.300 418.200 107.400 ;
        RECT 410.400 100.950 418.200 102.300 ;
        RECT 419.400 101.400 421.200 107.400 ;
        RECT 419.400 99.300 420.600 101.400 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 392.400 98.250 396.150 99.300 ;
        RECT 394.950 98.100 396.150 98.250 ;
        RECT 416.850 98.250 420.600 99.300 ;
        RECT 416.850 98.100 418.050 98.250 ;
        RECT 385.950 94.950 388.050 97.050 ;
        RECT 392.100 95.100 393.900 95.850 ;
        RECT 394.950 94.950 397.050 97.050 ;
        RECT 398.100 95.100 399.900 95.850 ;
        RECT 400.950 94.950 403.050 97.050 ;
        RECT 409.950 94.950 412.050 97.050 ;
        RECT 413.100 95.100 414.900 95.850 ;
        RECT 415.950 94.950 418.050 97.050 ;
        RECT 419.100 95.100 420.900 95.850 ;
        RECT 316.950 91.950 319.050 94.050 ;
        RECT 322.950 91.950 325.050 94.050 ;
        RECT 331.950 91.950 334.050 94.050 ;
        RECT 335.100 93.150 336.900 93.900 ;
        RECT 337.950 91.950 340.050 94.050 ;
        RECT 260.850 87.600 262.050 90.900 ;
        RECT 215.700 81.900 222.300 82.800 ;
        RECT 215.700 81.600 216.600 81.900 ;
        RECT 214.800 75.600 216.600 81.600 ;
        RECT 220.800 81.600 222.300 81.900 ;
        RECT 220.800 75.600 222.600 81.600 ;
        RECT 235.800 75.600 237.600 87.600 ;
        RECT 238.800 86.700 246.600 87.600 ;
        RECT 238.800 75.600 240.600 86.700 ;
        RECT 244.800 75.600 246.600 86.700 ;
        RECT 260.700 75.600 262.500 87.600 ;
        RECT 278.400 81.600 279.600 90.900 ;
        RECT 292.950 88.950 295.050 91.050 ;
        RECT 298.950 88.950 304.050 91.050 ;
        RECT 313.950 90.450 316.050 91.050 ;
        RECT 308.550 89.550 316.050 90.450 ;
        RECT 293.100 87.150 294.900 87.900 ;
        RECT 299.400 82.800 300.300 87.900 ;
        RECT 293.700 81.900 300.300 82.800 ;
        RECT 308.550 82.050 309.450 89.550 ;
        RECT 313.950 88.950 316.050 89.550 ;
        RECT 319.950 88.950 322.050 91.050 ;
        RECT 314.700 82.800 315.600 87.900 ;
        RECT 320.100 87.150 321.900 87.900 ;
        RECT 341.700 87.600 342.600 93.900 ;
        RECT 355.800 91.950 358.050 94.050 ;
        RECT 332.400 86.700 340.200 87.600 ;
        RECT 293.700 81.600 295.200 81.900 ;
        RECT 278.400 75.600 280.200 81.600 ;
        RECT 293.400 75.600 295.200 81.600 ;
        RECT 299.400 81.600 300.300 81.900 ;
        RECT 299.400 75.600 301.200 81.600 ;
        RECT 307.950 79.950 310.050 82.050 ;
        RECT 314.700 81.900 321.300 82.800 ;
        RECT 314.700 81.600 315.600 81.900 ;
        RECT 313.800 75.600 315.600 81.600 ;
        RECT 319.800 81.600 321.300 81.900 ;
        RECT 319.800 75.600 321.600 81.600 ;
        RECT 332.400 75.600 334.200 86.700 ;
        RECT 338.400 75.600 340.200 86.700 ;
        RECT 341.400 75.600 343.200 87.600 ;
        RECT 356.550 85.050 357.450 91.950 ;
        RECT 359.850 90.900 360.900 93.900 ;
        RECT 361.950 91.950 364.200 94.050 ;
        RECT 365.100 93.150 366.900 93.900 ;
        RECT 373.950 91.950 379.050 94.050 ;
        RECT 359.850 87.600 361.050 90.900 ;
        RECT 355.950 82.950 358.050 85.050 ;
        RECT 359.700 75.600 361.500 87.600 ;
        RECT 377.400 81.600 378.600 90.900 ;
        RECT 377.400 75.600 379.200 81.600 ;
        RECT 386.550 79.050 387.450 94.950 ;
        RECT 428.550 94.050 429.450 100.950 ;
        RECT 437.100 99.000 438.900 107.400 ;
        RECT 457.200 103.050 459.000 107.400 ;
        RECT 457.200 101.400 462.600 103.050 ;
        RECT 434.700 97.350 438.900 99.000 ;
        RECT 461.700 98.100 462.600 101.400 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 391.950 91.950 394.050 94.050 ;
        RECT 395.850 90.900 396.900 93.900 ;
        RECT 397.950 91.950 400.050 94.050 ;
        RECT 401.100 93.150 402.900 93.900 ;
        RECT 410.100 93.150 411.900 93.900 ;
        RECT 412.950 91.950 415.050 94.050 ;
        RECT 416.100 90.900 417.150 93.900 ;
        RECT 418.950 91.950 421.050 94.050 ;
        RECT 427.950 91.950 430.050 94.050 ;
        RECT 434.700 92.100 435.600 97.350 ;
        RECT 437.100 95.100 438.900 95.850 ;
        RECT 443.100 95.100 444.900 95.850 ;
        RECT 452.100 95.100 453.900 95.850 ;
        RECT 454.800 94.950 457.050 97.050 ;
        RECT 458.100 95.100 459.900 95.850 ;
        RECT 460.950 94.950 463.050 97.050 ;
        RECT 436.950 91.950 439.050 94.050 ;
        RECT 442.950 91.950 445.050 94.050 ;
        RECT 451.950 91.950 454.050 94.050 ;
        RECT 455.100 93.150 456.900 93.900 ;
        RECT 457.950 91.950 460.050 94.050 ;
        RECT 395.850 87.600 397.050 90.900 ;
        RECT 415.950 87.600 417.150 90.900 ;
        RECT 433.950 90.450 436.050 91.050 ;
        RECT 428.550 89.550 436.050 90.450 ;
        RECT 385.950 76.950 388.050 79.050 ;
        RECT 395.700 75.600 397.500 87.600 ;
        RECT 415.500 75.600 417.300 87.600 ;
        RECT 428.550 82.050 429.450 89.550 ;
        RECT 433.950 88.950 436.050 89.550 ;
        RECT 439.800 88.950 442.050 91.050 ;
        RECT 434.700 82.800 435.600 87.900 ;
        RECT 440.100 87.150 441.900 87.900 ;
        RECT 461.700 87.600 462.600 93.900 ;
        RECT 452.400 86.700 460.200 87.600 ;
        RECT 427.950 79.950 430.050 82.050 ;
        RECT 434.700 81.900 441.300 82.800 ;
        RECT 434.700 81.600 435.600 81.900 ;
        RECT 433.800 75.600 435.600 81.600 ;
        RECT 439.800 81.600 441.300 81.900 ;
        RECT 439.800 75.600 441.600 81.600 ;
        RECT 452.400 75.600 454.200 86.700 ;
        RECT 458.400 75.600 460.200 86.700 ;
        RECT 461.400 75.600 463.200 87.600 ;
        RECT 467.550 79.050 468.450 100.950 ;
        RECT 477.000 100.200 478.800 107.400 ;
        RECT 494.400 104.400 496.200 107.400 ;
        RECT 477.000 99.300 480.600 100.200 ;
        RECT 479.400 95.100 480.600 99.300 ;
        RECT 490.950 97.950 493.050 100.050 ;
        RECT 491.100 96.150 492.900 96.900 ;
        RECT 494.400 95.100 495.600 104.400 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 476.100 92.100 477.900 92.850 ;
        RECT 478.800 91.950 481.050 94.050 ;
        RECT 493.950 93.450 496.050 94.050 ;
        RECT 482.100 92.100 483.900 92.850 ;
        RECT 488.550 92.550 496.050 93.450 ;
        RECT 475.950 88.950 478.050 91.050 ;
        RECT 479.400 81.600 480.600 90.900 ;
        RECT 481.950 88.950 484.050 91.050 ;
        RECT 488.550 85.050 489.450 92.550 ;
        RECT 493.950 91.950 496.050 92.550 ;
        RECT 503.550 91.050 504.450 100.950 ;
        RECT 510.000 100.200 511.800 107.400 ;
        RECT 531.000 103.050 532.800 107.400 ;
        RECT 527.400 101.400 532.800 103.050 ;
        RECT 545.400 102.300 547.200 107.400 ;
        RECT 551.400 102.300 553.200 107.400 ;
        RECT 510.000 99.300 513.600 100.200 ;
        RECT 512.400 95.100 513.600 99.300 ;
        RECT 527.400 98.100 528.300 101.400 ;
        RECT 545.400 100.950 553.200 102.300 ;
        RECT 554.400 101.400 556.200 107.400 ;
        RECT 554.400 99.300 555.600 101.400 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 551.850 98.250 555.600 99.300 ;
        RECT 551.850 98.100 553.050 98.250 ;
        RECT 520.950 96.450 525.000 97.050 ;
        RECT 526.950 96.450 529.050 97.050 ;
        RECT 520.950 95.550 529.050 96.450 ;
        RECT 520.950 94.950 525.000 95.550 ;
        RECT 526.950 94.950 529.050 95.550 ;
        RECT 530.100 95.100 531.900 95.850 ;
        RECT 532.950 94.950 535.050 97.050 ;
        RECT 536.100 95.100 537.900 95.850 ;
        RECT 544.950 94.950 547.050 97.050 ;
        RECT 548.100 95.100 549.900 95.850 ;
        RECT 550.950 94.950 553.050 97.050 ;
        RECT 554.100 95.100 555.900 95.850 ;
        RECT 509.100 92.100 510.900 92.850 ;
        RECT 511.950 91.950 514.050 94.050 ;
        RECT 515.100 92.100 516.900 92.850 ;
        RECT 487.950 82.950 490.050 85.050 ;
        RECT 466.950 76.950 469.050 79.050 ;
        RECT 478.800 75.600 480.600 81.600 ;
        RECT 494.400 81.600 495.600 90.900 ;
        RECT 502.950 88.950 505.050 91.050 ;
        RECT 508.950 88.950 511.050 91.050 ;
        RECT 512.400 81.600 513.600 90.900 ;
        RECT 514.950 88.950 517.050 91.050 ;
        RECT 515.550 87.000 516.450 88.950 ;
        RECT 527.400 87.600 528.300 93.900 ;
        RECT 529.950 91.950 532.050 94.050 ;
        RECT 533.100 93.150 534.900 93.900 ;
        RECT 535.950 91.950 538.050 94.050 ;
        RECT 545.100 93.150 546.900 93.900 ;
        RECT 547.950 91.950 550.050 94.050 ;
        RECT 551.100 90.900 552.150 93.900 ;
        RECT 553.950 91.950 556.050 94.050 ;
        RECT 560.550 91.050 561.450 100.950 ;
        RECT 570.000 100.200 571.800 107.400 ;
        RECT 588.300 103.200 590.100 107.400 ;
        RECT 588.150 101.400 590.100 103.200 ;
        RECT 570.000 99.300 573.600 100.200 ;
        RECT 572.400 95.100 573.600 99.300 ;
        RECT 588.150 98.100 589.050 101.400 ;
        RECT 590.100 99.900 591.900 100.500 ;
        RECT 595.800 99.900 597.600 107.400 ;
        RECT 608.400 104.400 610.200 107.400 ;
        RECT 628.800 104.400 630.600 107.400 ;
        RECT 608.400 101.100 609.600 104.400 ;
        RECT 629.400 101.100 630.600 104.400 ;
        RECT 644.400 104.400 646.200 107.400 ;
        RECT 662.400 104.400 664.200 107.400 ;
        RECT 644.400 101.100 645.600 104.400 ;
        RECT 662.400 101.100 663.600 104.400 ;
        RECT 682.200 103.050 684.000 107.400 ;
        RECT 670.950 100.950 673.050 103.050 ;
        RECT 682.200 101.400 687.600 103.050 ;
        RECT 590.100 98.700 597.600 99.900 ;
        RECT 586.950 94.950 589.050 97.050 ;
        RECT 590.100 95.100 591.900 95.850 ;
        RECT 569.100 92.100 570.900 92.850 ;
        RECT 571.950 91.950 574.050 94.050 ;
        RECT 575.100 92.100 576.900 92.850 ;
        RECT 550.950 87.600 552.150 90.900 ;
        RECT 559.950 88.950 562.050 91.050 ;
        RECT 568.950 88.950 571.050 91.050 ;
        RECT 514.950 82.950 517.050 87.000 ;
        RECT 494.400 75.600 496.200 81.600 ;
        RECT 511.800 75.600 513.600 81.600 ;
        RECT 526.800 75.600 528.600 87.600 ;
        RECT 529.800 86.700 537.600 87.600 ;
        RECT 529.800 75.600 531.600 86.700 ;
        RECT 535.800 75.600 537.600 86.700 ;
        RECT 550.500 75.600 552.300 87.600 ;
        RECT 572.400 81.600 573.600 90.900 ;
        RECT 574.950 88.950 580.050 91.050 ;
        RECT 586.950 87.600 588.000 93.900 ;
        RECT 589.950 91.950 592.050 94.050 ;
        RECT 571.800 75.600 573.600 81.600 ;
        RECT 586.200 75.600 588.000 87.600 ;
        RECT 593.550 81.600 594.600 98.700 ;
        RECT 607.950 97.950 610.050 100.050 ;
        RECT 628.950 97.950 631.050 100.050 ;
        RECT 643.950 97.950 646.200 100.050 ;
        RECT 661.800 97.950 664.050 100.050 ;
        RECT 595.950 94.950 598.050 97.050 ;
        RECT 604.950 94.950 607.050 97.050 ;
        RECT 608.700 93.900 609.900 96.900 ;
        RECT 610.950 94.950 613.050 97.050 ;
        RECT 616.950 94.950 619.050 97.050 ;
        RECT 625.950 94.950 628.050 97.050 ;
        RECT 596.100 93.150 597.900 93.900 ;
        RECT 605.100 93.150 606.900 93.900 ;
        RECT 608.700 88.650 610.050 93.900 ;
        RECT 611.100 93.150 612.900 93.900 ;
        RECT 617.550 91.050 618.450 94.950 ;
        RECT 629.100 93.900 630.300 96.900 ;
        RECT 631.950 94.950 634.050 97.050 ;
        RECT 640.950 94.950 643.050 97.050 ;
        RECT 644.700 93.900 645.900 96.900 ;
        RECT 646.950 94.950 649.050 97.050 ;
        RECT 658.950 94.950 661.050 97.050 ;
        RECT 662.700 93.900 663.900 96.900 ;
        RECT 664.950 94.950 667.200 97.050 ;
        RECT 626.100 93.150 627.900 93.900 ;
        RECT 616.950 88.950 619.050 91.050 ;
        RECT 628.950 88.650 630.300 93.900 ;
        RECT 632.100 93.150 633.900 93.900 ;
        RECT 641.100 93.150 642.900 93.900 ;
        RECT 608.700 87.600 611.400 88.650 ;
        RECT 592.800 75.600 594.600 81.600 ;
        RECT 609.600 75.600 611.400 87.600 ;
        RECT 627.600 87.600 630.300 88.650 ;
        RECT 644.700 88.650 646.050 93.900 ;
        RECT 647.100 93.150 648.900 93.900 ;
        RECT 659.100 93.150 660.900 93.900 ;
        RECT 662.700 88.650 664.050 93.900 ;
        RECT 665.100 93.150 666.900 93.900 ;
        RECT 644.700 87.600 647.400 88.650 ;
        RECT 662.700 87.600 665.400 88.650 ;
        RECT 627.600 75.600 629.400 87.600 ;
        RECT 645.600 75.600 647.400 87.600 ;
        RECT 663.600 75.600 665.400 87.600 ;
        RECT 671.550 79.050 672.450 100.950 ;
        RECT 686.700 98.100 687.600 101.400 ;
        RECT 698.400 102.300 700.200 107.400 ;
        RECT 704.400 102.300 706.200 107.400 ;
        RECT 698.400 100.950 706.200 102.300 ;
        RECT 707.400 101.400 709.200 107.400 ;
        RECT 707.400 99.300 708.600 101.400 ;
        RECT 724.200 100.200 726.000 107.400 ;
        RECT 739.800 104.400 741.600 107.400 ;
        RECT 704.850 98.250 708.600 99.300 ;
        RECT 722.400 99.300 726.000 100.200 ;
        RECT 704.850 98.100 706.050 98.250 ;
        RECT 677.100 95.100 678.900 95.850 ;
        RECT 679.950 94.950 682.050 97.050 ;
        RECT 685.950 96.450 688.050 97.050 ;
        RECT 683.100 95.100 684.900 95.850 ;
        RECT 685.950 95.550 693.450 96.450 ;
        RECT 685.950 94.950 688.050 95.550 ;
        RECT 676.950 91.950 679.050 94.050 ;
        RECT 680.100 93.150 681.900 93.900 ;
        RECT 682.950 91.950 685.050 94.050 ;
        RECT 686.700 87.600 687.600 93.900 ;
        RECT 692.550 88.050 693.450 95.550 ;
        RECT 697.950 94.950 700.050 97.050 ;
        RECT 701.100 95.100 702.900 95.850 ;
        RECT 703.950 94.950 706.050 97.050 ;
        RECT 707.100 95.100 708.900 95.850 ;
        RECT 722.400 95.100 723.600 99.300 ;
        RECT 740.400 95.100 741.600 104.400 ;
        RECT 742.950 97.950 745.050 103.050 ;
        RECT 752.400 102.300 754.200 107.400 ;
        RECT 758.400 102.300 760.200 107.400 ;
        RECT 752.400 100.950 760.200 102.300 ;
        RECT 761.400 101.400 763.200 107.400 ;
        RECT 766.950 103.950 769.050 106.050 ;
        RECT 761.400 99.300 762.600 101.400 ;
        RECT 758.850 98.250 762.600 99.300 ;
        RECT 758.850 98.100 760.050 98.250 ;
        RECT 743.100 96.150 744.900 96.900 ;
        RECT 751.950 94.950 754.050 97.050 ;
        RECT 755.100 95.100 756.900 95.850 ;
        RECT 757.950 94.950 760.200 97.050 ;
        RECT 761.100 95.100 762.900 95.850 ;
        RECT 767.550 94.050 768.450 103.950 ;
        RECT 779.100 99.000 780.900 107.400 ;
        RECT 799.200 103.050 801.000 107.400 ;
        RECT 818.400 104.400 820.200 107.400 ;
        RECT 799.200 101.400 804.600 103.050 ;
        RECT 776.700 97.350 780.900 99.000 ;
        RECT 803.700 98.100 804.600 101.400 ;
        RECT 814.950 97.950 817.050 100.050 ;
        RECT 698.100 93.150 699.900 93.900 ;
        RECT 700.950 91.950 703.050 94.050 ;
        RECT 704.100 90.900 705.150 93.900 ;
        RECT 706.950 91.950 709.050 94.050 ;
        RECT 719.100 92.100 720.900 92.850 ;
        RECT 721.800 91.950 724.050 94.050 ;
        RECT 725.100 92.100 726.900 92.850 ;
        RECT 736.950 91.950 742.050 94.050 ;
        RECT 752.100 93.150 753.900 93.900 ;
        RECT 754.950 91.950 757.050 94.050 ;
        RECT 677.400 86.700 685.200 87.600 ;
        RECT 670.950 76.950 673.050 79.050 ;
        RECT 677.400 75.600 679.200 86.700 ;
        RECT 683.400 75.600 685.200 86.700 ;
        RECT 686.400 75.600 688.200 87.600 ;
        RECT 691.950 85.950 694.050 88.050 ;
        RECT 703.950 87.600 705.150 90.900 ;
        RECT 718.950 88.950 721.050 91.050 ;
        RECT 703.500 75.600 705.300 87.600 ;
        RECT 722.400 81.600 723.600 90.900 ;
        RECT 724.950 88.950 727.200 91.050 ;
        RECT 758.100 90.900 759.150 93.900 ;
        RECT 760.950 91.950 763.050 94.050 ;
        RECT 766.950 91.950 769.050 94.050 ;
        RECT 776.700 92.100 777.600 97.350 ;
        RECT 779.100 95.100 780.900 95.850 ;
        RECT 785.100 95.100 786.900 95.850 ;
        RECT 794.100 95.100 795.900 95.850 ;
        RECT 796.950 94.950 799.050 97.050 ;
        RECT 800.100 95.100 801.900 95.850 ;
        RECT 802.950 94.950 805.050 97.050 ;
        RECT 815.100 96.150 816.900 96.900 ;
        RECT 818.400 95.100 819.600 104.400 ;
        RECT 835.200 100.200 837.000 107.400 ;
        RECT 850.800 104.400 852.600 107.400 ;
        RECT 833.400 99.300 837.000 100.200 ;
        RECT 833.400 95.100 834.600 99.300 ;
        RECT 851.400 95.100 852.600 104.400 ;
        RECT 853.950 97.950 856.050 100.050 ;
        RECT 854.100 96.150 855.900 96.900 ;
        RECT 778.950 91.950 781.050 94.050 ;
        RECT 784.950 91.950 787.050 94.050 ;
        RECT 793.950 91.950 796.050 94.050 ;
        RECT 797.100 93.150 798.900 93.900 ;
        RECT 799.950 91.950 802.050 94.050 ;
        RECT 740.400 81.600 741.600 90.900 ;
        RECT 757.950 87.600 759.150 90.900 ;
        RECT 772.950 88.950 778.050 91.050 ;
        RECT 781.800 88.950 784.050 91.050 ;
        RECT 722.400 75.600 724.200 81.600 ;
        RECT 739.800 75.600 741.600 81.600 ;
        RECT 757.500 75.600 759.300 87.600 ;
        RECT 776.700 82.800 777.600 87.900 ;
        RECT 782.100 87.150 783.900 87.900 ;
        RECT 803.700 87.600 804.600 93.900 ;
        RECT 817.950 91.950 823.050 94.050 ;
        RECT 830.100 92.100 831.900 92.850 ;
        RECT 832.950 91.950 835.050 94.050 ;
        RECT 836.100 92.100 837.900 92.850 ;
        RECT 847.950 91.950 853.050 94.050 ;
        RECT 794.400 86.700 802.200 87.600 ;
        RECT 776.700 81.900 783.300 82.800 ;
        RECT 776.700 81.600 777.600 81.900 ;
        RECT 775.800 75.600 777.600 81.600 ;
        RECT 781.800 81.600 783.300 81.900 ;
        RECT 781.800 75.600 783.600 81.600 ;
        RECT 794.400 75.600 796.200 86.700 ;
        RECT 800.400 75.600 802.200 86.700 ;
        RECT 803.400 75.600 805.200 87.600 ;
        RECT 818.400 81.600 819.600 90.900 ;
        RECT 829.950 88.950 832.050 91.050 ;
        RECT 833.400 81.600 834.600 90.900 ;
        RECT 835.950 85.950 838.050 91.050 ;
        RECT 851.400 81.600 852.600 90.900 ;
        RECT 818.400 75.600 820.200 81.600 ;
        RECT 833.400 75.600 835.200 81.600 ;
        RECT 850.800 75.600 852.600 81.600 ;
        RECT 10.800 65.400 12.600 71.400 ;
        RECT 11.700 65.100 12.600 65.400 ;
        RECT 16.800 65.400 18.600 71.400 ;
        RECT 16.800 65.100 18.300 65.400 ;
        RECT 11.700 64.200 18.300 65.100 ;
        RECT 11.700 59.100 12.600 64.200 ;
        RECT 29.400 60.300 31.200 71.400 ;
        RECT 35.400 60.300 37.200 71.400 ;
        RECT 17.100 59.100 18.900 59.850 ;
        RECT 29.400 59.400 37.200 60.300 ;
        RECT 38.400 59.400 40.200 71.400 ;
        RECT 55.500 59.400 57.300 71.400 ;
        RECT 73.800 65.400 75.600 71.400 ;
        RECT 74.700 65.100 75.600 65.400 ;
        RECT 79.800 65.400 81.600 71.400 ;
        RECT 94.800 70.500 102.600 71.400 ;
        RECT 79.800 65.100 81.300 65.400 ;
        RECT 74.700 64.200 81.300 65.100 ;
        RECT 10.950 57.450 13.050 58.050 ;
        RECT 5.550 56.550 13.050 57.450 ;
        RECT 5.550 43.050 6.450 56.550 ;
        RECT 10.950 55.950 13.050 56.550 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 11.700 49.650 12.600 54.900 ;
        RECT 13.950 52.950 16.050 55.050 ;
        RECT 19.950 52.950 22.050 55.050 ;
        RECT 28.800 52.950 31.050 55.050 ;
        RECT 32.100 53.100 33.900 53.850 ;
        RECT 34.950 52.950 37.050 55.050 ;
        RECT 38.700 53.100 39.600 59.400 ;
        RECT 43.950 55.950 46.050 58.050 ;
        RECT 55.950 56.100 57.150 59.400 ;
        RECT 74.700 59.100 75.600 64.200 ;
        RECT 80.100 59.100 81.900 59.850 ;
        RECT 94.800 59.400 96.600 70.500 ;
        RECT 97.800 58.500 99.600 69.600 ;
        RECT 100.800 60.600 102.600 70.500 ;
        RECT 106.800 60.600 108.600 71.400 ;
        RECT 113.100 64.950 115.200 67.050 ;
        RECT 100.800 59.700 108.600 60.600 ;
        RECT 14.100 51.150 15.900 51.900 ;
        RECT 20.100 51.150 21.900 51.900 ;
        RECT 29.100 51.150 30.900 51.900 ;
        RECT 31.950 49.950 34.050 52.050 ;
        RECT 35.100 51.150 36.900 51.900 ;
        RECT 37.950 51.450 40.050 52.050 ;
        RECT 44.550 51.450 45.450 55.950 ;
        RECT 50.100 53.100 51.900 53.850 ;
        RECT 52.950 52.950 55.050 55.050 ;
        RECT 56.100 53.100 57.150 56.100 ;
        RECT 73.950 55.950 76.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 88.950 55.950 91.050 58.050 ;
        RECT 97.800 57.600 101.850 58.500 ;
        RECT 113.550 58.050 114.450 64.950 ;
        RECT 122.700 59.400 124.500 71.400 ;
        RECT 139.800 65.400 141.600 71.400 ;
        RECT 140.700 65.100 141.600 65.400 ;
        RECT 145.800 65.400 147.600 71.400 ;
        RECT 145.800 65.100 147.300 65.400 ;
        RECT 140.700 64.200 147.300 65.100 ;
        RECT 100.950 56.100 101.850 57.600 ;
        RECT 58.950 52.950 61.050 55.050 ;
        RECT 37.950 50.550 45.450 51.450 ;
        RECT 37.950 49.950 40.050 50.550 ;
        RECT 11.700 48.000 15.900 49.650 ;
        RECT 4.950 40.950 7.050 43.050 ;
        RECT 14.100 39.600 15.900 48.000 ;
        RECT 38.700 45.600 39.600 48.900 ;
        RECT 44.550 46.050 45.450 50.550 ;
        RECT 46.950 49.950 52.050 52.050 ;
        RECT 53.100 51.150 54.900 51.900 ;
        RECT 55.950 49.950 58.050 52.050 ;
        RECT 59.100 51.150 60.900 51.900 ;
        RECT 74.700 49.650 75.600 54.900 ;
        RECT 76.950 52.950 79.050 55.050 ;
        RECT 82.950 52.950 85.050 55.050 ;
        RECT 89.550 52.050 90.450 55.950 ;
        RECT 95.100 53.100 96.900 53.850 ;
        RECT 97.800 52.950 100.050 55.050 ;
        RECT 101.100 53.100 101.850 56.100 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 122.850 56.100 124.050 59.400 ;
        RECT 140.700 59.100 141.600 64.200 ;
        RECT 158.400 60.300 160.200 71.400 ;
        RECT 164.400 60.300 166.200 71.400 ;
        RECT 146.100 59.100 147.900 59.850 ;
        RECT 158.400 59.400 166.200 60.300 ;
        RECT 167.400 59.400 169.200 71.400 ;
        RECT 175.950 67.950 178.050 70.050 ;
        RECT 103.950 52.950 106.050 55.050 ;
        RECT 107.100 53.100 108.750 53.850 ;
        RECT 118.950 52.950 121.050 55.050 ;
        RECT 122.850 53.100 123.900 56.100 ;
        RECT 136.950 55.950 142.050 58.050 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 124.950 52.950 127.050 55.050 ;
        RECT 128.100 53.100 129.900 53.850 ;
        RECT 77.100 51.150 78.900 51.900 ;
        RECT 83.100 51.150 84.900 51.900 ;
        RECT 88.950 49.950 91.050 52.050 ;
        RECT 94.800 49.950 97.050 52.050 ;
        RECT 98.250 51.150 99.900 51.900 ;
        RECT 100.950 49.950 103.050 52.050 ;
        RECT 104.100 51.150 105.750 51.900 ;
        RECT 106.800 49.950 109.050 52.050 ;
        RECT 119.100 51.150 120.900 51.900 ;
        RECT 121.950 49.950 124.050 52.050 ;
        RECT 125.100 51.150 126.900 51.900 ;
        RECT 127.950 49.950 130.050 52.050 ;
        RECT 140.700 49.650 141.600 54.900 ;
        RECT 142.950 52.950 145.050 55.050 ;
        RECT 148.950 52.950 151.050 55.050 ;
        RECT 157.950 52.950 160.050 55.050 ;
        RECT 161.100 53.100 162.900 53.850 ;
        RECT 163.950 52.950 166.050 55.050 ;
        RECT 167.700 53.100 168.600 59.400 ;
        RECT 173.100 58.950 175.200 61.050 ;
        RECT 143.100 51.150 144.900 51.900 ;
        RECT 149.100 51.150 150.900 51.900 ;
        RECT 158.100 51.150 159.900 51.900 ;
        RECT 56.850 48.750 58.050 48.900 ;
        RECT 56.850 47.700 60.600 48.750 ;
        RECT 74.700 48.000 78.900 49.650 ;
        RECT 34.200 43.950 39.600 45.600 ;
        RECT 43.950 43.950 46.050 46.050 ;
        RECT 50.400 44.700 58.200 46.050 ;
        RECT 34.200 39.600 36.000 43.950 ;
        RECT 50.400 39.600 52.200 44.700 ;
        RECT 56.400 39.600 58.200 44.700 ;
        RECT 59.400 45.600 60.600 47.700 ;
        RECT 59.400 39.600 61.200 45.600 ;
        RECT 77.100 39.600 78.900 48.000 ;
        RECT 102.000 45.600 103.050 48.900 ;
        RECT 121.950 48.750 123.150 48.900 ;
        RECT 119.400 47.700 123.150 48.750 ;
        RECT 140.700 48.000 144.900 49.650 ;
        RECT 119.400 45.600 120.600 47.700 ;
        RECT 102.000 39.600 103.800 45.600 ;
        RECT 118.800 39.600 120.600 45.600 ;
        RECT 121.800 44.700 129.600 46.050 ;
        RECT 121.800 39.600 123.600 44.700 ;
        RECT 127.800 39.600 129.600 44.700 ;
        RECT 143.100 39.600 144.900 48.000 ;
        RECT 160.950 46.950 163.050 52.050 ;
        RECT 164.100 51.150 165.900 51.900 ;
        RECT 166.950 51.450 169.050 52.050 ;
        RECT 173.550 51.450 174.450 58.950 ;
        RECT 176.550 52.050 177.450 67.950 ;
        RECT 185.700 59.400 187.500 71.400 ;
        RECT 196.950 67.950 199.050 70.050 ;
        RECT 185.850 56.100 187.050 59.400 ;
        RECT 181.950 52.950 184.050 55.050 ;
        RECT 185.850 53.100 186.900 56.100 ;
        RECT 187.950 52.950 190.050 55.050 ;
        RECT 191.100 53.100 192.900 53.850 ;
        RECT 197.550 52.050 198.450 67.950 ;
        RECT 202.800 65.400 204.600 71.400 ;
        RECT 203.700 65.100 204.600 65.400 ;
        RECT 208.800 65.400 210.600 71.400 ;
        RECT 208.800 65.100 210.300 65.400 ;
        RECT 203.700 64.200 210.300 65.100 ;
        RECT 217.950 64.950 220.050 67.050 ;
        RECT 203.700 59.100 204.600 64.200 ;
        RECT 209.100 59.100 210.900 59.850 ;
        RECT 199.950 55.950 205.050 58.050 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 166.950 50.550 174.450 51.450 ;
        RECT 166.950 49.950 169.050 50.550 ;
        RECT 175.950 49.950 178.050 52.050 ;
        RECT 182.100 51.150 183.900 51.900 ;
        RECT 184.950 49.950 187.050 52.050 ;
        RECT 188.100 51.150 189.900 51.900 ;
        RECT 190.950 49.950 193.050 52.050 ;
        RECT 196.950 49.950 199.050 52.050 ;
        RECT 203.700 49.650 204.600 54.900 ;
        RECT 205.950 52.950 208.050 55.050 ;
        RECT 211.950 52.950 214.050 55.050 ;
        RECT 206.100 51.150 207.900 51.900 ;
        RECT 212.100 51.150 213.900 51.900 ;
        RECT 218.550 51.450 219.450 64.950 ;
        RECT 223.800 59.400 225.600 71.400 ;
        RECT 226.800 60.300 228.600 71.400 ;
        RECT 232.800 60.300 234.600 71.400 ;
        RECT 226.800 59.400 234.600 60.300 ;
        RECT 244.200 59.400 246.000 71.400 ;
        RECT 250.800 65.400 252.600 71.400 ;
        RECT 224.400 53.100 225.300 59.400 ;
        RECT 226.950 52.950 229.050 55.050 ;
        RECT 230.100 53.100 231.900 53.850 ;
        RECT 232.950 52.950 235.200 55.050 ;
        RECT 244.950 53.100 246.000 59.400 ;
        RECT 247.950 52.950 250.050 55.050 ;
        RECT 223.950 51.450 226.050 52.050 ;
        RECT 218.550 50.550 226.050 51.450 ;
        RECT 227.100 51.150 228.900 51.900 ;
        RECT 223.950 49.950 226.050 50.550 ;
        RECT 229.950 49.950 232.050 52.050 ;
        RECT 233.100 51.150 234.900 51.900 ;
        RECT 241.950 49.950 247.050 52.050 ;
        RECT 248.100 51.150 249.900 51.900 ;
        RECT 167.700 45.600 168.600 48.900 ;
        RECT 184.950 48.750 186.150 48.900 ;
        RECT 182.400 47.700 186.150 48.750 ;
        RECT 203.700 48.000 207.900 49.650 ;
        RECT 182.400 45.600 183.600 47.700 ;
        RECT 163.200 43.950 168.600 45.600 ;
        RECT 163.200 39.600 165.000 43.950 ;
        RECT 181.800 39.600 183.600 45.600 ;
        RECT 184.800 44.700 192.600 46.050 ;
        RECT 184.800 39.600 186.600 44.700 ;
        RECT 190.800 39.600 192.600 44.700 ;
        RECT 206.100 39.600 207.900 48.000 ;
        RECT 224.400 45.600 225.300 48.900 ;
        RECT 246.150 45.600 247.050 48.900 ;
        RECT 251.550 48.300 252.600 65.400 ;
        RECT 266.400 65.400 268.200 71.400 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 266.400 56.100 267.600 65.400 ;
        RECT 281.400 60.300 283.200 71.400 ;
        RECT 287.400 60.300 289.200 71.400 ;
        RECT 281.400 59.400 289.200 60.300 ;
        RECT 290.400 59.400 292.200 71.400 ;
        RECT 295.950 64.950 298.050 67.050 ;
        RECT 305.400 65.400 307.200 71.400 ;
        RECT 305.700 65.100 307.200 65.400 ;
        RECT 311.400 65.400 313.200 71.400 ;
        RECT 326.400 65.400 328.200 71.400 ;
        RECT 343.800 65.400 345.600 71.400 ;
        RECT 359.400 65.400 361.200 71.400 ;
        RECT 311.400 65.100 312.300 65.400 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 263.100 54.150 264.900 54.900 ;
        RECT 254.100 53.100 255.900 53.850 ;
        RECT 265.950 52.950 268.050 55.050 ;
        RECT 269.100 54.150 270.900 54.900 ;
        RECT 280.950 52.950 283.050 58.050 ;
        RECT 284.100 53.100 285.900 53.850 ;
        RECT 286.950 52.950 289.050 55.050 ;
        RECT 290.700 53.100 291.600 59.400 ;
        RECT 253.950 49.950 256.050 52.050 ;
        RECT 248.100 47.100 255.600 48.300 ;
        RECT 248.100 46.500 249.900 47.100 ;
        RECT 224.400 43.950 229.800 45.600 ;
        RECT 228.000 39.600 229.800 43.950 ;
        RECT 246.150 43.800 248.100 45.600 ;
        RECT 246.300 39.600 248.100 43.800 ;
        RECT 253.800 39.600 255.600 47.100 ;
        RECT 266.400 47.700 267.600 51.900 ;
        RECT 281.100 51.150 282.900 51.900 ;
        RECT 283.950 49.950 286.050 52.050 ;
        RECT 287.100 51.150 288.900 51.900 ;
        RECT 289.950 51.450 292.050 52.050 ;
        RECT 296.550 51.450 297.450 64.950 ;
        RECT 305.700 64.200 312.300 65.100 ;
        RECT 305.100 59.100 306.900 59.850 ;
        RECT 311.400 59.100 312.300 64.200 ;
        RECT 316.950 61.950 319.050 64.050 ;
        RECT 304.950 55.950 307.050 58.050 ;
        RECT 310.950 57.450 313.050 58.050 ;
        RECT 317.550 57.450 318.450 61.950 ;
        RECT 310.950 56.550 318.450 57.450 ;
        RECT 310.950 55.950 313.050 56.550 ;
        RECT 322.950 55.950 325.050 58.050 ;
        RECT 326.400 56.100 327.600 65.400 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 344.400 56.100 345.600 65.400 ;
        RECT 359.700 65.100 361.200 65.400 ;
        RECT 365.400 65.400 367.200 71.400 ;
        RECT 379.800 65.400 381.600 71.400 ;
        RECT 365.400 65.100 366.300 65.400 ;
        RECT 359.700 64.200 366.300 65.100 ;
        RECT 349.950 61.950 352.050 64.050 ;
        RECT 301.950 52.950 304.050 55.050 ;
        RECT 307.950 52.950 310.050 55.050 ;
        RECT 289.950 50.550 297.450 51.450 ;
        RECT 302.100 51.150 303.900 51.900 ;
        RECT 308.100 51.150 309.900 51.900 ;
        RECT 289.950 49.950 292.050 50.550 ;
        RECT 311.400 49.650 312.300 54.900 ;
        RECT 323.100 54.150 324.900 54.900 ;
        RECT 325.950 52.950 328.050 55.050 ;
        RECT 329.100 54.150 330.900 54.900 ;
        RECT 343.950 54.450 346.050 55.050 ;
        RECT 350.550 54.450 351.450 61.950 ;
        RECT 359.100 59.100 360.900 59.850 ;
        RECT 365.400 59.100 366.300 64.200 ;
        RECT 380.700 65.100 381.600 65.400 ;
        RECT 385.800 65.400 387.600 71.400 ;
        RECT 401.400 65.400 403.200 71.400 ;
        RECT 409.950 67.950 412.050 70.050 ;
        RECT 385.800 65.100 387.300 65.400 ;
        RECT 380.700 64.200 387.300 65.100 ;
        RECT 380.700 59.100 381.600 64.200 ;
        RECT 386.100 59.100 387.900 59.850 ;
        RECT 358.950 55.950 361.200 58.050 ;
        RECT 364.950 57.450 367.050 58.050 ;
        RECT 364.950 56.550 372.450 57.450 ;
        RECT 364.950 55.950 367.050 56.550 ;
        RECT 371.550 55.050 372.450 56.550 ;
        RECT 376.950 55.950 382.050 58.050 ;
        RECT 385.950 55.950 388.050 58.050 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 401.400 56.100 402.600 65.400 ;
        RECT 403.950 55.950 406.050 58.050 ;
        RECT 410.550 55.050 411.450 67.950 ;
        RECT 416.400 60.300 418.200 71.400 ;
        RECT 422.400 60.300 424.200 71.400 ;
        RECT 416.400 59.400 424.200 60.300 ;
        RECT 425.400 59.400 427.200 71.400 ;
        RECT 437.400 60.600 439.200 71.400 ;
        RECT 443.400 70.500 451.200 71.400 ;
        RECT 443.400 60.600 445.200 70.500 ;
        RECT 437.400 59.700 445.200 60.600 ;
        RECT 343.950 53.550 351.450 54.450 ;
        RECT 343.950 52.950 346.050 53.550 ;
        RECT 355.950 52.950 358.050 55.050 ;
        RECT 361.950 52.950 364.050 55.050 ;
        RECT 313.950 49.950 316.050 52.050 ;
        RECT 266.400 46.800 270.000 47.700 ;
        RECT 268.200 39.600 270.000 46.800 ;
        RECT 290.700 45.600 291.600 48.900 ;
        RECT 286.200 43.950 291.600 45.600 ;
        RECT 308.100 48.000 312.300 49.650 ;
        RECT 286.200 39.600 288.000 43.950 ;
        RECT 308.100 39.600 309.900 48.000 ;
        RECT 314.550 43.050 315.450 49.950 ;
        RECT 326.400 47.700 327.600 51.900 ;
        RECT 326.400 46.800 330.000 47.700 ;
        RECT 313.800 40.950 315.900 43.050 ;
        RECT 328.200 39.600 330.000 46.800 ;
        RECT 344.400 42.600 345.600 51.900 ;
        RECT 356.100 51.150 357.900 51.900 ;
        RECT 362.100 51.150 363.900 51.900 ;
        RECT 347.100 50.100 348.900 50.850 ;
        RECT 365.400 49.650 366.300 54.900 ;
        RECT 371.550 53.550 376.050 55.050 ;
        RECT 372.000 52.950 376.050 53.550 ;
        RECT 346.950 46.950 349.050 49.050 ;
        RECT 362.100 48.000 366.300 49.650 ;
        RECT 380.700 49.650 381.600 54.900 ;
        RECT 382.950 52.950 385.050 55.050 ;
        RECT 388.950 52.950 391.050 55.050 ;
        RECT 398.100 54.150 399.900 54.900 ;
        RECT 400.950 52.950 403.050 55.050 ;
        RECT 404.100 54.150 405.900 54.900 ;
        RECT 409.800 52.950 411.900 55.050 ;
        RECT 415.950 52.950 418.050 55.050 ;
        RECT 419.100 53.100 420.900 53.850 ;
        RECT 421.950 52.950 424.050 55.050 ;
        RECT 425.700 53.100 426.600 59.400 ;
        RECT 446.400 58.500 448.200 69.600 ;
        RECT 449.400 59.400 451.200 70.500 ;
        RECT 455.550 59.400 457.350 71.400 ;
        RECT 463.050 65.400 464.850 71.400 ;
        RECT 460.950 63.300 464.850 65.400 ;
        RECT 470.850 64.500 472.650 71.400 ;
        RECT 478.650 65.400 480.450 71.400 ;
        RECT 479.250 64.500 480.450 65.400 ;
        RECT 469.950 63.450 476.550 64.500 ;
        RECT 469.950 62.700 471.750 63.450 ;
        RECT 474.750 62.700 476.550 63.450 ;
        RECT 479.250 62.400 484.050 64.500 ;
        RECT 462.150 60.600 464.850 62.400 ;
        RECT 465.750 61.800 467.550 62.400 ;
        RECT 465.750 60.900 472.050 61.800 ;
        RECT 479.250 61.500 480.450 62.400 ;
        RECT 465.750 60.600 467.550 60.900 ;
        RECT 463.950 59.700 464.850 60.600 ;
        RECT 430.950 55.950 433.050 58.050 ;
        RECT 444.150 57.600 448.200 58.500 ;
        RECT 444.150 56.100 445.050 57.600 ;
        RECT 383.100 51.150 384.900 51.900 ;
        RECT 389.100 51.150 390.900 51.900 ;
        RECT 380.700 48.000 384.900 49.650 ;
        RECT 343.800 39.600 345.600 42.600 ;
        RECT 362.100 39.600 363.900 48.000 ;
        RECT 383.100 39.600 384.900 48.000 ;
        RECT 401.400 47.700 402.600 51.900 ;
        RECT 416.100 51.150 417.900 51.900 ;
        RECT 418.950 49.950 421.050 52.050 ;
        RECT 422.100 51.150 423.900 51.900 ;
        RECT 424.950 51.450 427.050 52.050 ;
        RECT 431.550 51.450 432.450 55.950 ;
        RECT 437.250 53.100 438.900 53.850 ;
        RECT 439.800 52.950 442.050 55.050 ;
        RECT 444.150 53.100 444.900 56.100 ;
        RECT 445.950 52.950 448.200 55.050 ;
        RECT 449.100 53.100 450.900 53.850 ;
        RECT 455.550 52.050 456.750 59.400 ;
        RECT 460.950 58.800 463.050 59.700 ;
        RECT 463.950 58.800 469.950 59.700 ;
        RECT 458.850 57.600 463.050 58.800 ;
        RECT 457.950 55.800 459.750 57.600 ;
        RECT 469.050 53.100 469.950 58.800 ;
        RECT 471.150 58.800 472.050 60.900 ;
        RECT 472.950 60.300 480.450 61.500 ;
        RECT 472.950 59.700 474.750 60.300 ;
        RECT 487.050 59.400 488.850 71.400 ;
        RECT 477.750 58.800 488.850 59.400 ;
        RECT 471.150 58.200 488.850 58.800 ;
        RECT 471.150 57.900 479.550 58.200 ;
        RECT 477.750 57.600 479.550 57.900 ;
        RECT 482.100 52.800 483.900 53.100 ;
        RECT 424.950 50.550 432.450 51.450 ;
        RECT 424.950 49.950 427.050 50.550 ;
        RECT 436.950 49.950 439.050 52.050 ;
        RECT 440.250 51.150 441.900 51.900 ;
        RECT 442.800 49.950 445.050 52.050 ;
        RECT 446.100 51.150 447.750 51.900 ;
        RECT 448.950 49.950 451.050 52.050 ;
        RECT 455.550 49.950 456.900 52.050 ;
        RECT 457.950 49.950 460.050 52.050 ;
        RECT 461.100 49.950 461.850 51.750 ;
        RECT 469.800 49.950 472.050 52.050 ;
        RECT 475.950 49.950 478.050 52.050 ;
        RECT 479.100 51.900 483.900 52.800 ;
        RECT 482.100 51.300 483.900 51.900 ;
        RECT 485.100 51.150 486.900 52.950 ;
        RECT 479.100 50.400 480.900 51.000 ;
        RECT 485.100 50.400 486.000 51.150 ;
        RECT 401.400 46.800 405.000 47.700 ;
        RECT 403.200 39.600 405.000 46.800 ;
        RECT 425.700 45.600 426.600 48.900 ;
        RECT 442.950 45.600 444.000 48.900 ;
        RECT 421.200 43.950 426.600 45.600 ;
        RECT 421.200 39.600 423.000 43.950 ;
        RECT 442.200 39.600 444.000 45.600 ;
        RECT 455.550 45.600 456.750 49.950 ;
        RECT 479.100 49.200 486.000 50.400 ;
        RECT 469.050 48.000 469.950 48.900 ;
        RECT 479.100 48.000 480.150 49.200 ;
        RECT 469.050 47.100 480.150 48.000 ;
        RECT 469.050 46.800 469.950 47.100 ;
        RECT 455.550 39.600 457.350 45.600 ;
        RECT 460.950 44.700 463.050 45.600 ;
        RECT 468.150 45.000 469.950 46.800 ;
        RECT 479.100 46.200 480.150 47.100 ;
        RECT 475.350 45.450 477.150 46.200 ;
        RECT 460.950 43.500 464.700 44.700 ;
        RECT 463.650 42.600 464.700 43.500 ;
        RECT 472.200 44.400 477.150 45.450 ;
        RECT 478.650 44.400 480.450 46.200 ;
        RECT 487.950 45.600 488.850 58.200 ;
        RECT 500.400 65.400 502.200 71.400 ;
        RECT 500.400 56.100 501.600 65.400 ;
        RECT 512.400 60.600 514.200 71.400 ;
        RECT 518.400 70.500 526.200 71.400 ;
        RECT 518.400 60.600 520.200 70.500 ;
        RECT 512.400 59.700 520.200 60.600 ;
        RECT 521.400 58.500 523.200 69.600 ;
        RECT 524.400 59.400 526.200 70.500 ;
        RECT 536.400 65.400 538.200 71.400 ;
        RECT 519.150 57.600 523.200 58.500 ;
        RECT 536.400 58.500 537.600 65.400 ;
        RECT 542.700 59.400 544.500 71.400 ;
        RECT 556.500 59.400 558.300 71.400 ;
        RECT 562.800 65.400 564.600 71.400 ;
        RECT 574.800 65.400 576.600 71.400 ;
        RECT 536.400 57.600 542.100 58.500 ;
        RECT 519.150 56.100 520.050 57.600 ;
        RECT 540.150 56.700 542.100 57.600 ;
        RECT 499.950 52.950 505.050 55.050 ;
        RECT 512.250 53.100 513.900 53.850 ;
        RECT 514.950 52.950 517.050 55.050 ;
        RECT 519.150 53.100 519.900 56.100 ;
        RECT 520.950 52.950 523.050 55.050 ;
        RECT 524.100 53.100 525.900 53.850 ;
        RECT 536.100 53.100 537.900 53.850 ;
        RECT 540.150 53.100 541.050 56.700 ;
        RECT 543.000 53.100 544.200 59.400 ;
        RECT 556.800 53.100 558.000 59.400 ;
        RECT 563.400 58.500 564.600 65.400 ;
        RECT 575.700 65.100 576.600 65.400 ;
        RECT 580.800 65.400 582.600 71.400 ;
        RECT 580.800 65.100 582.300 65.400 ;
        RECT 575.700 64.200 582.300 65.100 ;
        RECT 575.700 59.100 576.600 64.200 ;
        RECT 581.100 59.100 582.900 59.850 ;
        RECT 599.700 59.400 601.500 71.400 ;
        RECT 617.400 65.400 619.200 71.400 ;
        RECT 631.800 65.400 633.600 71.400 ;
        RECT 558.900 57.600 564.600 58.500 ;
        RECT 558.900 56.700 560.850 57.600 ;
        RECT 559.950 53.100 560.850 56.700 ;
        RECT 571.950 55.950 577.050 58.050 ;
        RECT 580.950 55.950 583.050 58.050 ;
        RECT 599.850 56.100 601.050 59.400 ;
        RECT 617.400 56.100 618.600 65.400 ;
        RECT 632.700 65.100 633.600 65.400 ;
        RECT 637.800 65.400 639.600 71.400 ;
        RECT 653.400 65.400 655.200 71.400 ;
        RECT 637.800 65.100 639.300 65.400 ;
        RECT 632.700 64.200 639.300 65.100 ;
        RECT 632.700 59.100 633.600 64.200 ;
        RECT 638.100 59.100 639.900 59.850 ;
        RECT 563.100 53.100 564.900 53.850 ;
        RECT 497.100 50.100 498.900 50.850 ;
        RECT 493.950 46.950 499.050 49.050 ;
        RECT 472.200 42.600 473.250 44.400 ;
        RECT 481.950 43.500 484.050 45.600 ;
        RECT 481.950 42.600 483.000 43.500 ;
        RECT 463.650 39.600 465.450 42.600 ;
        RECT 471.450 39.600 473.250 42.600 ;
        RECT 479.250 41.700 483.000 42.600 ;
        RECT 479.250 39.600 481.050 41.700 ;
        RECT 487.050 39.600 488.850 45.600 ;
        RECT 500.400 42.600 501.600 51.900 ;
        RECT 511.950 49.950 514.050 52.050 ;
        RECT 515.250 51.150 516.900 51.900 ;
        RECT 517.950 49.950 520.050 52.050 ;
        RECT 521.100 51.150 522.750 51.900 ;
        RECT 523.950 49.950 526.050 52.050 ;
        RECT 535.950 49.950 538.050 52.050 ;
        RECT 540.150 48.900 540.900 53.100 ;
        RECT 560.100 48.900 560.850 53.100 ;
        RECT 562.950 49.950 565.050 52.050 ;
        RECT 517.950 45.600 519.000 48.900 ;
        RECT 540.150 48.300 541.050 48.900 ;
        RECT 540.150 47.400 542.100 48.300 ;
        RECT 500.400 39.600 502.200 42.600 ;
        RECT 517.200 39.600 519.000 45.600 ;
        RECT 537.000 46.500 542.100 47.400 ;
        RECT 537.000 42.600 538.200 46.500 ;
        RECT 543.000 45.600 544.200 48.900 ;
        RECT 556.800 45.600 558.000 48.900 ;
        RECT 559.950 48.300 560.850 48.900 ;
        RECT 558.900 47.400 560.850 48.300 ;
        RECT 575.700 49.650 576.600 54.900 ;
        RECT 577.950 52.950 580.050 55.050 ;
        RECT 599.850 53.100 600.900 56.100 ;
        RECT 631.950 55.950 634.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 649.800 55.950 652.050 58.050 ;
        RECT 653.400 56.100 654.600 65.400 ;
        RECT 664.950 64.950 667.050 67.050 ;
        RECT 673.800 65.400 675.600 71.400 ;
        RECT 691.800 65.400 693.600 71.400 ;
        RECT 706.800 65.400 708.600 71.400 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 601.950 52.950 604.050 55.050 ;
        RECT 605.100 53.100 606.900 53.850 ;
        RECT 616.950 52.950 622.050 55.050 ;
        RECT 578.100 51.150 579.900 51.900 ;
        RECT 584.100 51.150 585.900 51.900 ;
        RECT 596.100 51.150 597.900 51.900 ;
        RECT 598.950 49.950 601.050 52.050 ;
        RECT 602.100 51.150 603.900 51.900 ;
        RECT 604.950 49.950 607.050 52.050 ;
        RECT 614.100 50.100 615.900 50.850 ;
        RECT 575.700 48.000 579.900 49.650 ;
        RECT 598.950 48.750 600.150 48.900 ;
        RECT 558.900 46.500 564.000 47.400 ;
        RECT 536.400 39.600 538.200 42.600 ;
        RECT 542.700 39.600 544.500 45.600 ;
        RECT 556.500 39.600 558.300 45.600 ;
        RECT 562.800 42.600 564.000 46.500 ;
        RECT 562.800 39.600 564.600 42.600 ;
        RECT 578.100 39.600 579.900 48.000 ;
        RECT 596.400 47.700 600.150 48.750 ;
        RECT 596.400 45.600 597.600 47.700 ;
        RECT 613.950 46.950 616.050 49.050 ;
        RECT 595.800 39.600 597.600 45.600 ;
        RECT 598.800 44.700 606.600 46.050 ;
        RECT 598.800 39.600 600.600 44.700 ;
        RECT 604.800 39.600 606.600 44.700 ;
        RECT 617.400 42.600 618.600 51.900 ;
        RECT 632.700 49.650 633.600 54.900 ;
        RECT 634.950 52.950 637.050 55.050 ;
        RECT 640.950 52.950 643.050 55.050 ;
        RECT 650.100 54.150 651.900 54.900 ;
        RECT 652.950 52.950 655.050 55.050 ;
        RECT 656.100 54.150 657.900 54.900 ;
        RECT 665.550 52.050 666.450 64.950 ;
        RECT 670.950 55.950 673.050 58.050 ;
        RECT 674.400 56.100 675.600 65.400 ;
        RECT 676.950 55.950 679.050 58.050 ;
        RECT 688.800 55.950 691.050 58.050 ;
        RECT 692.400 56.100 693.600 65.400 ;
        RECT 707.700 65.100 708.600 65.400 ;
        RECT 712.800 65.400 714.600 71.400 ;
        RECT 712.800 65.100 714.300 65.400 ;
        RECT 707.700 64.200 714.300 65.100 ;
        RECT 700.950 61.950 703.050 64.050 ;
        RECT 694.950 55.950 697.050 58.050 ;
        RECT 701.550 57.450 702.450 61.950 ;
        RECT 707.700 59.100 708.600 64.200 ;
        RECT 725.400 60.300 727.200 71.400 ;
        RECT 731.400 60.300 733.200 71.400 ;
        RECT 713.100 59.100 714.900 59.850 ;
        RECT 725.400 59.400 733.200 60.300 ;
        RECT 734.400 59.400 736.200 71.400 ;
        RECT 739.950 64.950 742.050 67.050 ;
        RECT 751.800 65.400 753.600 71.400 ;
        RECT 766.800 65.400 768.600 71.400 ;
        RECT 706.950 57.450 709.050 58.050 ;
        RECT 701.550 56.550 709.050 57.450 ;
        RECT 706.950 55.950 709.050 56.550 ;
        RECT 712.950 55.950 715.050 58.050 ;
        RECT 671.100 54.150 672.900 54.900 ;
        RECT 673.950 52.950 676.200 55.050 ;
        RECT 677.100 54.150 678.900 54.900 ;
        RECT 689.100 54.150 690.900 54.900 ;
        RECT 691.950 52.950 694.050 55.050 ;
        RECT 695.100 54.150 696.900 54.900 ;
        RECT 635.100 51.150 636.900 51.900 ;
        RECT 641.100 51.150 642.900 51.900 ;
        RECT 632.700 48.000 636.900 49.650 ;
        RECT 617.400 39.600 619.200 42.600 ;
        RECT 635.100 39.600 636.900 48.000 ;
        RECT 653.400 47.700 654.600 51.900 ;
        RECT 664.950 49.950 667.050 52.050 ;
        RECT 674.400 47.700 675.600 51.900 ;
        RECT 692.400 47.700 693.600 51.900 ;
        RECT 707.700 49.650 708.600 54.900 ;
        RECT 709.950 52.950 712.050 55.050 ;
        RECT 715.950 52.950 718.050 55.050 ;
        RECT 724.950 52.950 727.050 55.050 ;
        RECT 728.100 53.100 729.900 53.850 ;
        RECT 730.950 52.950 733.050 55.050 ;
        RECT 734.700 53.100 735.600 59.400 ;
        RECT 740.550 55.050 741.450 64.950 ;
        RECT 748.950 55.950 751.050 58.050 ;
        RECT 752.400 56.100 753.600 65.400 ;
        RECT 767.700 65.100 768.600 65.400 ;
        RECT 772.800 65.400 774.600 71.400 ;
        RECT 787.800 65.400 789.600 71.400 ;
        RECT 772.800 65.100 774.300 65.400 ;
        RECT 767.700 64.200 774.300 65.100 ;
        RECT 788.700 65.100 789.600 65.400 ;
        RECT 793.800 65.400 795.600 71.400 ;
        RECT 793.800 65.100 795.300 65.400 ;
        RECT 788.700 64.200 795.300 65.100 ;
        RECT 767.700 59.100 768.600 64.200 ;
        RECT 773.100 59.100 774.900 59.850 ;
        RECT 788.700 59.100 789.600 64.200 ;
        RECT 802.950 61.950 805.050 64.050 ;
        RECT 794.100 59.100 795.900 59.850 ;
        RECT 754.950 55.950 757.050 58.050 ;
        RECT 766.950 57.450 769.050 58.050 ;
        RECT 761.550 56.550 769.050 57.450 ;
        RECT 739.950 52.950 742.050 55.050 ;
        RECT 749.100 54.150 750.900 54.900 ;
        RECT 751.950 52.950 754.050 55.050 ;
        RECT 755.100 54.150 756.900 54.900 ;
        RECT 710.100 51.150 711.900 51.900 ;
        RECT 716.100 51.150 717.900 51.900 ;
        RECT 725.100 51.150 726.900 51.900 ;
        RECT 727.950 49.950 730.050 52.050 ;
        RECT 731.100 51.150 732.900 51.900 ;
        RECT 733.950 51.450 736.050 52.050 ;
        RECT 733.950 50.550 741.450 51.450 ;
        RECT 733.950 49.950 736.050 50.550 ;
        RECT 707.700 48.000 711.900 49.650 ;
        RECT 653.400 46.800 657.000 47.700 ;
        RECT 655.200 39.600 657.000 46.800 ;
        RECT 672.000 46.800 675.600 47.700 ;
        RECT 690.000 46.800 693.600 47.700 ;
        RECT 672.000 39.600 673.800 46.800 ;
        RECT 690.000 39.600 691.800 46.800 ;
        RECT 710.100 39.600 711.900 48.000 ;
        RECT 734.700 45.600 735.600 48.900 ;
        RECT 740.550 46.050 741.450 50.550 ;
        RECT 752.400 47.700 753.600 51.900 ;
        RECT 750.000 46.800 753.600 47.700 ;
        RECT 730.200 43.950 735.600 45.600 ;
        RECT 739.950 43.950 742.050 46.050 ;
        RECT 730.200 39.600 732.000 43.950 ;
        RECT 750.000 39.600 751.800 46.800 ;
        RECT 761.550 43.050 762.450 56.550 ;
        RECT 766.950 55.950 769.050 56.550 ;
        RECT 772.950 55.950 775.050 58.050 ;
        RECT 781.950 57.450 786.000 58.050 ;
        RECT 787.950 57.450 790.050 58.050 ;
        RECT 781.950 56.550 790.050 57.450 ;
        RECT 781.950 55.950 786.000 56.550 ;
        RECT 787.950 55.950 790.050 56.550 ;
        RECT 793.950 55.950 796.050 58.050 ;
        RECT 767.700 49.650 768.600 54.900 ;
        RECT 769.950 52.950 772.050 55.050 ;
        RECT 775.800 52.950 778.050 55.050 ;
        RECT 770.100 51.150 771.900 51.900 ;
        RECT 776.100 51.150 777.900 51.900 ;
        RECT 788.700 49.650 789.600 54.900 ;
        RECT 790.800 52.950 793.050 55.050 ;
        RECT 796.950 52.950 799.050 55.050 ;
        RECT 791.100 51.150 792.900 51.900 ;
        RECT 797.100 51.150 798.900 51.900 ;
        RECT 767.700 48.000 771.900 49.650 ;
        RECT 788.700 48.000 792.900 49.650 ;
        RECT 803.550 49.050 804.450 61.950 ;
        RECT 812.700 59.400 814.500 71.400 ;
        RECT 823.950 61.950 826.050 64.050 ;
        RECT 812.850 56.100 814.050 59.400 ;
        RECT 808.950 52.950 811.050 55.050 ;
        RECT 812.850 53.100 813.900 56.100 ;
        RECT 814.950 52.950 817.050 55.050 ;
        RECT 818.100 53.100 819.900 53.850 ;
        RECT 824.550 52.050 825.450 61.950 ;
        RECT 833.700 59.400 835.500 71.400 ;
        RECT 850.800 65.400 852.600 71.400 ;
        RECT 833.850 56.100 835.050 59.400 ;
        RECT 851.400 56.100 852.600 65.400 ;
        RECT 829.950 52.950 832.050 55.050 ;
        RECT 833.850 53.100 834.900 56.100 ;
        RECT 835.950 52.950 838.050 55.050 ;
        RECT 839.100 53.100 840.900 53.850 ;
        RECT 847.950 52.950 853.050 55.050 ;
        RECT 809.100 51.150 810.900 51.900 ;
        RECT 811.950 49.950 814.050 52.050 ;
        RECT 815.100 51.150 816.900 51.900 ;
        RECT 817.950 49.950 820.050 52.050 ;
        RECT 823.950 49.950 826.050 52.050 ;
        RECT 830.100 51.150 831.900 51.900 ;
        RECT 832.950 49.950 835.050 52.050 ;
        RECT 836.100 51.150 837.900 51.900 ;
        RECT 838.950 49.950 841.050 52.050 ;
        RECT 760.950 40.950 763.050 43.050 ;
        RECT 770.100 39.600 771.900 48.000 ;
        RECT 791.100 39.600 792.900 48.000 ;
        RECT 802.950 46.950 805.050 49.050 ;
        RECT 811.950 48.750 813.150 48.900 ;
        RECT 832.950 48.750 834.150 48.900 ;
        RECT 809.400 47.700 813.150 48.750 ;
        RECT 830.400 47.700 834.150 48.750 ;
        RECT 809.400 45.600 810.600 47.700 ;
        RECT 808.800 39.600 810.600 45.600 ;
        RECT 811.800 44.700 819.600 46.050 ;
        RECT 830.400 45.600 831.600 47.700 ;
        RECT 811.800 39.600 813.600 44.700 ;
        RECT 817.800 39.600 819.600 44.700 ;
        RECT 829.800 39.600 831.600 45.600 ;
        RECT 832.800 44.700 840.600 46.050 ;
        RECT 832.800 39.600 834.600 44.700 ;
        RECT 838.800 39.600 840.600 44.700 ;
        RECT 851.400 42.600 852.600 51.900 ;
        RECT 854.100 50.100 855.900 50.850 ;
        RECT 853.950 46.950 856.050 49.050 ;
        RECT 850.800 39.600 852.600 42.600 ;
        RECT 10.800 32.400 12.600 35.400 ;
        RECT 11.400 23.100 12.600 32.400 ;
        RECT 13.950 25.950 16.050 28.050 ;
        RECT 29.100 27.000 30.900 35.400 ;
        RECT 46.800 29.400 48.600 35.400 ;
        RECT 47.400 27.300 48.600 29.400 ;
        RECT 49.800 30.300 51.600 35.400 ;
        RECT 55.800 30.300 57.600 35.400 ;
        RECT 49.800 28.950 57.600 30.300 ;
        RECT 65.400 30.300 67.200 35.400 ;
        RECT 71.400 30.300 73.200 35.400 ;
        RECT 65.400 28.950 73.200 30.300 ;
        RECT 74.400 29.400 76.200 35.400 ;
        RECT 74.400 27.300 75.600 29.400 ;
        RECT 29.100 25.350 33.300 27.000 ;
        RECT 47.400 26.250 51.150 27.300 ;
        RECT 49.950 26.100 51.150 26.250 ;
        RECT 71.850 26.250 75.600 27.300 ;
        RECT 92.100 27.000 93.900 35.400 ;
        RECT 113.100 27.000 114.900 35.400 ;
        RECT 134.100 27.000 135.900 35.400 ;
        RECT 152.400 32.400 154.200 35.400 ;
        RECT 71.850 26.100 73.050 26.250 ;
        RECT 92.100 25.350 96.300 27.000 ;
        RECT 113.100 25.350 117.300 27.000 ;
        RECT 134.100 25.350 138.300 27.000 ;
        RECT 148.950 25.950 151.050 28.050 ;
        RECT 14.100 24.150 15.900 24.900 ;
        RECT 23.100 23.100 24.900 23.850 ;
        RECT 29.100 23.100 30.900 23.850 ;
        RECT 10.950 19.950 16.050 22.050 ;
        RECT 22.800 19.950 25.050 22.050 ;
        RECT 28.950 19.950 31.050 22.050 ;
        RECT 32.400 20.100 33.300 25.350 ;
        RECT 47.100 23.100 48.900 23.850 ;
        RECT 49.950 22.950 52.050 25.050 ;
        RECT 53.100 23.100 54.900 23.850 ;
        RECT 55.950 22.950 58.050 25.050 ;
        RECT 64.950 22.950 67.050 25.050 ;
        RECT 68.100 23.100 69.900 23.850 ;
        RECT 70.950 22.950 73.050 25.050 ;
        RECT 74.100 23.100 75.900 23.850 ;
        RECT 86.100 23.100 87.900 23.850 ;
        RECT 92.100 23.100 93.900 23.850 ;
        RECT 46.950 19.950 49.050 22.050 ;
        RECT 11.400 9.600 12.600 18.900 ;
        RECT 25.950 16.950 28.050 19.050 ;
        RECT 31.950 18.450 34.050 19.050 ;
        RECT 50.850 18.900 51.900 21.900 ;
        RECT 52.950 19.950 55.050 22.050 ;
        RECT 56.100 21.150 57.900 21.900 ;
        RECT 65.100 21.150 66.900 21.900 ;
        RECT 67.950 19.950 70.050 22.050 ;
        RECT 71.100 18.900 72.150 21.900 ;
        RECT 73.950 19.950 76.050 22.050 ;
        RECT 85.950 19.950 88.050 22.050 ;
        RECT 91.950 19.950 94.050 22.050 ;
        RECT 95.400 20.100 96.300 25.350 ;
        RECT 107.100 23.100 108.900 23.850 ;
        RECT 113.100 23.100 114.900 23.850 ;
        RECT 106.950 19.950 109.050 22.050 ;
        RECT 112.950 19.950 115.050 22.050 ;
        RECT 116.400 20.100 117.300 25.350 ;
        RECT 128.100 23.100 129.900 23.850 ;
        RECT 134.100 23.100 135.900 23.850 ;
        RECT 127.950 19.950 130.050 22.050 ;
        RECT 133.950 19.950 136.050 22.050 ;
        RECT 137.400 20.100 138.300 25.350 ;
        RECT 149.100 24.150 150.900 24.900 ;
        RECT 152.400 23.100 153.600 32.400 ;
        RECT 160.950 25.950 163.050 28.050 ;
        RECT 170.100 27.000 171.900 35.400 ;
        RECT 190.200 31.050 192.000 35.400 ;
        RECT 212.400 32.400 214.200 35.400 ;
        RECT 218.400 32.400 220.200 35.400 ;
        RECT 213.150 31.500 214.200 32.400 ;
        RECT 219.150 31.500 220.200 32.400 ;
        RECT 190.200 29.400 195.600 31.050 ;
        RECT 213.150 30.600 223.950 31.500 ;
        RECT 148.950 19.950 154.050 22.050 ;
        RECT 31.950 17.550 39.450 18.450 ;
        RECT 31.950 16.950 34.050 17.550 ;
        RECT 26.100 15.150 27.900 15.900 ;
        RECT 32.400 10.800 33.300 15.900 ;
        RECT 26.700 9.900 33.300 10.800 ;
        RECT 26.700 9.600 28.200 9.900 ;
        RECT 10.800 3.600 12.600 9.600 ;
        RECT 26.400 3.600 28.200 9.600 ;
        RECT 32.400 9.600 33.300 9.900 ;
        RECT 32.400 3.600 34.200 9.600 ;
        RECT 38.550 7.050 39.450 17.550 ;
        RECT 50.850 15.600 52.050 18.900 ;
        RECT 70.950 15.600 72.150 18.900 ;
        RECT 88.950 16.950 91.050 19.050 ;
        RECT 94.950 16.950 100.050 19.050 ;
        RECT 109.950 16.950 112.050 19.050 ;
        RECT 115.950 18.450 118.050 19.050 ;
        RECT 120.000 18.450 124.050 19.050 ;
        RECT 115.950 17.550 124.050 18.450 ;
        RECT 115.950 16.950 118.050 17.550 ;
        RECT 120.000 16.950 124.050 17.550 ;
        RECT 130.950 16.950 133.050 19.050 ;
        RECT 136.950 18.450 139.050 19.050 ;
        RECT 136.950 17.550 144.450 18.450 ;
        RECT 136.950 16.950 139.050 17.550 ;
        RECT 37.950 4.950 40.050 7.050 ;
        RECT 50.700 3.600 52.500 15.600 ;
        RECT 70.500 3.600 72.300 15.600 ;
        RECT 89.100 15.150 90.900 15.900 ;
        RECT 95.400 10.800 96.300 15.900 ;
        RECT 110.100 15.150 111.900 15.900 ;
        RECT 116.400 10.800 117.300 15.900 ;
        RECT 131.100 15.150 132.900 15.900 ;
        RECT 137.400 10.800 138.300 15.900 ;
        RECT 143.550 13.050 144.450 17.550 ;
        RECT 142.950 10.950 145.050 13.050 ;
        RECT 89.700 9.900 96.300 10.800 ;
        RECT 89.700 9.600 91.200 9.900 ;
        RECT 89.400 3.600 91.200 9.600 ;
        RECT 95.400 9.600 96.300 9.900 ;
        RECT 110.700 9.900 117.300 10.800 ;
        RECT 110.700 9.600 112.200 9.900 ;
        RECT 95.400 3.600 97.200 9.600 ;
        RECT 110.400 3.600 112.200 9.600 ;
        RECT 116.400 9.600 117.300 9.900 ;
        RECT 131.700 9.900 138.300 10.800 ;
        RECT 131.700 9.600 133.200 9.900 ;
        RECT 116.400 3.600 118.200 9.600 ;
        RECT 131.400 3.600 133.200 9.600 ;
        RECT 137.400 9.600 138.300 9.900 ;
        RECT 152.400 9.600 153.600 18.900 ;
        RECT 161.550 18.450 162.450 25.950 ;
        RECT 167.700 25.350 171.900 27.000 ;
        RECT 194.700 26.100 195.600 29.400 ;
        RECT 167.700 20.100 168.600 25.350 ;
        RECT 196.950 25.050 199.050 25.200 ;
        RECT 170.100 23.100 171.900 23.850 ;
        RECT 176.100 23.100 177.900 23.850 ;
        RECT 185.100 23.100 186.900 23.850 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 191.100 23.100 192.900 23.850 ;
        RECT 193.950 23.100 199.050 25.050 ;
        RECT 208.950 23.100 211.050 25.200 ;
        RECT 215.100 23.250 216.900 24.000 ;
        RECT 217.950 23.100 220.050 28.050 ;
        RECT 222.750 23.250 223.950 30.600 ;
        RECT 229.950 28.950 232.050 31.050 ;
        RECT 239.400 30.300 241.200 35.400 ;
        RECT 245.400 30.300 247.200 35.400 ;
        RECT 239.400 28.950 247.200 30.300 ;
        RECT 248.400 29.400 250.200 35.400 ;
        RECT 263.400 32.400 265.200 35.400 ;
        RECT 193.950 22.950 198.450 23.100 ;
        RECT 169.950 19.950 172.050 22.050 ;
        RECT 175.950 19.950 178.200 22.050 ;
        RECT 184.950 19.950 187.050 22.050 ;
        RECT 188.100 21.150 189.900 21.900 ;
        RECT 190.950 19.950 193.050 22.050 ;
        RECT 166.950 18.450 169.050 19.050 ;
        RECT 161.550 17.550 169.050 18.450 ;
        RECT 166.950 16.950 169.050 17.550 ;
        RECT 172.950 16.950 175.050 19.050 ;
        RECT 167.700 10.800 168.600 15.900 ;
        RECT 173.100 15.150 174.900 15.900 ;
        RECT 194.700 15.600 195.600 21.900 ;
        RECT 209.100 21.300 210.900 22.050 ;
        RECT 214.950 19.950 217.050 22.200 ;
        RECT 218.100 21.300 219.900 22.050 ;
        RECT 222.750 19.050 222.900 23.250 ;
        RECT 223.950 21.450 226.050 22.200 ;
        RECT 230.550 21.450 231.450 28.950 ;
        RECT 248.400 27.300 249.600 29.400 ;
        RECT 245.850 26.250 249.600 27.300 ;
        RECT 245.850 26.100 247.050 26.250 ;
        RECT 259.950 25.950 262.050 28.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 242.100 23.100 243.900 23.850 ;
        RECT 244.950 22.950 247.050 25.050 ;
        RECT 260.100 24.150 261.900 24.900 ;
        RECT 248.100 23.100 249.900 23.850 ;
        RECT 263.400 23.100 264.600 32.400 ;
        RECT 277.800 29.400 279.600 35.400 ;
        RECT 278.400 27.300 279.600 29.400 ;
        RECT 280.800 30.300 282.600 35.400 ;
        RECT 286.800 30.300 288.600 35.400 ;
        RECT 280.800 28.950 288.600 30.300 ;
        RECT 299.400 32.400 301.200 35.400 ;
        RECT 278.400 26.250 282.150 27.300 ;
        RECT 280.950 26.100 282.150 26.250 ;
        RECT 295.950 25.950 298.050 28.050 ;
        RECT 278.100 23.100 279.900 23.850 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 284.100 23.100 285.900 23.850 ;
        RECT 286.950 22.950 289.050 25.050 ;
        RECT 296.100 24.150 297.900 24.900 ;
        RECT 299.400 23.100 300.600 32.400 ;
        RECT 311.400 30.300 313.200 35.400 ;
        RECT 317.400 30.300 319.200 35.400 ;
        RECT 311.400 28.950 319.200 30.300 ;
        RECT 320.400 29.400 322.200 35.400 ;
        RECT 320.400 27.300 321.600 29.400 ;
        RECT 337.200 28.200 339.000 35.400 ;
        RECT 352.800 29.400 354.600 35.400 ;
        RECT 317.850 26.250 321.600 27.300 ;
        RECT 335.400 27.300 339.000 28.200 ;
        RECT 353.400 27.300 354.600 29.400 ;
        RECT 355.800 30.300 357.600 35.400 ;
        RECT 361.800 30.300 363.600 35.400 ;
        RECT 355.800 28.950 363.600 30.300 ;
        RECT 375.000 28.200 376.800 35.400 ;
        RECT 391.800 32.400 393.600 35.400 ;
        RECT 404.400 32.400 406.200 35.400 ;
        RECT 375.000 27.300 378.600 28.200 ;
        RECT 317.850 26.100 319.050 26.250 ;
        RECT 310.950 22.950 313.050 25.050 ;
        RECT 314.100 23.100 315.900 23.850 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 320.100 23.100 321.900 23.850 ;
        RECT 335.400 23.100 336.600 27.300 ;
        RECT 353.400 26.250 357.150 27.300 ;
        RECT 355.950 26.100 357.150 26.250 ;
        RECT 353.100 23.100 354.900 23.850 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 359.100 23.100 360.900 23.850 ;
        RECT 361.950 22.950 364.050 25.050 ;
        RECT 377.400 23.100 378.600 27.300 ;
        RECT 392.400 23.100 393.600 32.400 ;
        RECT 405.000 28.500 406.200 32.400 ;
        RECT 410.700 29.400 412.500 35.400 ;
        RECT 424.800 32.400 426.600 35.400 ;
        RECT 394.950 25.950 400.050 28.050 ;
        RECT 405.000 27.600 410.100 28.500 ;
        RECT 408.150 26.700 410.100 27.600 ;
        RECT 408.150 26.100 409.050 26.700 ;
        RECT 411.000 26.100 412.200 29.400 ;
        RECT 395.100 24.150 396.900 24.900 ;
        RECT 403.800 22.950 406.050 25.050 ;
        RECT 223.950 20.550 231.450 21.450 ;
        RECT 239.100 21.150 240.900 21.900 ;
        RECT 223.950 20.100 226.050 20.550 ;
        RECT 241.950 19.950 244.050 22.050 ;
        RECT 222.750 16.800 223.950 19.050 ;
        RECT 245.100 18.900 246.150 21.900 ;
        RECT 247.950 19.950 250.050 22.050 ;
        RECT 262.950 21.450 265.050 22.050 ;
        RECT 267.000 21.450 271.050 22.050 ;
        RECT 262.950 20.550 271.050 21.450 ;
        RECT 262.950 19.950 265.050 20.550 ;
        RECT 267.000 19.950 271.050 20.550 ;
        RECT 277.950 19.950 280.050 22.050 ;
        RECT 281.850 18.900 282.900 21.900 ;
        RECT 283.950 19.950 286.200 22.050 ;
        RECT 287.100 21.150 288.900 21.900 ;
        RECT 298.950 19.950 304.050 22.050 ;
        RECT 311.100 21.150 312.900 21.900 ;
        RECT 313.950 19.950 316.050 22.050 ;
        RECT 317.100 18.900 318.150 21.900 ;
        RECT 319.950 19.950 322.050 22.050 ;
        RECT 332.100 20.100 333.900 20.850 ;
        RECT 334.950 19.950 337.050 22.050 ;
        RECT 338.100 20.100 339.900 20.850 ;
        RECT 352.800 19.950 355.050 22.050 ;
        RECT 222.750 15.600 226.200 16.800 ;
        RECT 244.950 15.600 246.150 18.900 ;
        RECT 185.400 14.700 193.200 15.600 ;
        RECT 167.700 9.900 174.300 10.800 ;
        RECT 167.700 9.600 168.600 9.900 ;
        RECT 137.400 3.600 139.200 9.600 ;
        RECT 152.400 3.600 154.200 9.600 ;
        RECT 166.800 3.600 168.600 9.600 ;
        RECT 172.800 9.600 174.300 9.900 ;
        RECT 172.800 3.600 174.600 9.600 ;
        RECT 185.400 3.600 187.200 14.700 ;
        RECT 191.400 3.600 193.200 14.700 ;
        RECT 194.400 3.600 196.200 15.600 ;
        RECT 206.400 13.500 214.200 14.400 ;
        RECT 206.400 3.600 208.200 13.500 ;
        RECT 212.400 4.500 214.200 13.500 ;
        RECT 215.400 13.200 223.800 14.100 ;
        RECT 215.400 5.400 217.200 13.200 ;
        RECT 218.400 4.500 220.200 12.300 ;
        RECT 212.400 3.600 220.200 4.500 ;
        RECT 222.000 4.500 223.800 13.200 ;
        RECT 225.000 13.200 226.200 15.600 ;
        RECT 225.000 5.400 226.800 13.200 ;
        RECT 228.000 4.500 229.800 13.800 ;
        RECT 222.000 3.600 229.800 4.500 ;
        RECT 244.500 3.600 246.300 15.600 ;
        RECT 263.400 9.600 264.600 18.900 ;
        RECT 281.850 15.600 283.050 18.900 ;
        RECT 263.400 3.600 265.200 9.600 ;
        RECT 281.700 3.600 283.500 15.600 ;
        RECT 299.400 9.600 300.600 18.900 ;
        RECT 316.950 15.600 318.150 18.900 ;
        RECT 331.950 16.950 334.050 19.050 ;
        RECT 299.400 3.600 301.200 9.600 ;
        RECT 316.500 3.600 318.300 15.600 ;
        RECT 335.400 9.600 336.600 18.900 ;
        RECT 337.950 16.950 340.200 19.050 ;
        RECT 356.850 18.900 357.900 21.900 ;
        RECT 358.950 19.950 361.050 22.050 ;
        RECT 362.100 21.150 363.900 21.900 ;
        RECT 374.100 20.100 375.900 20.850 ;
        RECT 376.950 19.950 379.050 22.050 ;
        RECT 380.100 20.100 381.900 20.850 ;
        RECT 391.950 19.950 397.050 22.050 ;
        RECT 408.150 21.900 408.900 26.100 ;
        RECT 425.400 23.100 426.600 32.400 ;
        RECT 432.150 29.400 433.950 35.400 ;
        RECT 439.950 33.300 441.750 35.400 ;
        RECT 438.000 32.400 441.750 33.300 ;
        RECT 447.750 32.400 449.550 35.400 ;
        RECT 455.550 32.400 457.350 35.400 ;
        RECT 438.000 31.500 439.050 32.400 ;
        RECT 436.950 29.400 439.050 31.500 ;
        RECT 447.750 30.600 448.800 32.400 ;
        RECT 427.950 25.950 430.050 28.050 ;
        RECT 428.100 24.150 429.900 24.900 ;
        RECT 404.100 21.150 405.900 21.900 ;
        RECT 356.850 15.600 358.050 18.900 ;
        RECT 373.950 16.950 376.050 19.050 ;
        RECT 335.400 3.600 337.200 9.600 ;
        RECT 356.700 3.600 358.500 15.600 ;
        RECT 377.400 9.600 378.600 18.900 ;
        RECT 379.950 16.950 385.050 19.050 ;
        RECT 392.400 9.600 393.600 18.900 ;
        RECT 408.150 18.300 409.050 21.900 ;
        RECT 408.150 17.400 410.100 18.300 ;
        RECT 376.800 3.600 378.600 9.600 ;
        RECT 391.800 3.600 393.600 9.600 ;
        RECT 404.400 16.500 410.100 17.400 ;
        RECT 404.400 9.600 405.600 16.500 ;
        RECT 411.000 15.600 412.200 21.900 ;
        RECT 424.950 19.950 427.050 22.050 ;
        RECT 404.400 3.600 406.200 9.600 ;
        RECT 410.700 3.600 412.500 15.600 ;
        RECT 425.400 9.600 426.600 18.900 ;
        RECT 424.800 3.600 426.600 9.600 ;
        RECT 432.150 16.800 433.050 29.400 ;
        RECT 440.550 28.800 442.350 30.600 ;
        RECT 443.850 29.550 448.800 30.600 ;
        RECT 456.300 31.500 457.350 32.400 ;
        RECT 456.300 30.300 460.050 31.500 ;
        RECT 443.850 28.800 445.650 29.550 ;
        RECT 440.850 27.900 441.900 28.800 ;
        RECT 451.050 28.200 452.850 30.000 ;
        RECT 457.950 29.400 460.050 30.300 ;
        RECT 463.650 29.400 465.450 35.400 ;
        RECT 475.500 29.400 477.300 35.400 ;
        RECT 481.800 32.400 483.600 35.400 ;
        RECT 451.050 27.900 451.950 28.200 ;
        RECT 440.850 27.000 451.950 27.900 ;
        RECT 440.850 25.800 441.900 27.000 ;
        RECT 451.050 26.100 451.950 27.000 ;
        RECT 435.000 24.600 441.900 25.800 ;
        RECT 464.250 25.050 465.450 29.400 ;
        RECT 475.800 26.100 477.000 29.400 ;
        RECT 481.800 28.500 483.000 32.400 ;
        RECT 493.500 29.400 495.300 35.400 ;
        RECT 499.800 32.400 501.600 35.400 ;
        RECT 511.800 32.400 513.600 35.400 ;
        RECT 477.900 27.600 483.000 28.500 ;
        RECT 477.900 26.700 479.850 27.600 ;
        RECT 478.950 26.100 479.850 26.700 ;
        RECT 493.800 26.100 495.000 29.400 ;
        RECT 499.800 28.500 501.000 32.400 ;
        RECT 495.900 27.600 501.000 28.500 ;
        RECT 495.900 26.700 497.850 27.600 ;
        RECT 496.950 26.100 497.850 26.700 ;
        RECT 435.000 23.850 435.900 24.600 ;
        RECT 440.100 24.000 441.900 24.600 ;
        RECT 434.100 22.050 435.900 23.850 ;
        RECT 437.100 23.100 438.900 23.700 ;
        RECT 437.100 22.200 441.900 23.100 ;
        RECT 442.950 22.950 445.050 25.050 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 459.150 23.250 459.900 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 464.100 22.950 465.450 25.050 ;
        RECT 437.100 21.900 438.900 22.200 ;
        RECT 441.450 17.100 443.250 17.400 ;
        RECT 441.450 16.800 449.850 17.100 ;
        RECT 432.150 16.200 449.850 16.800 ;
        RECT 432.150 15.600 443.250 16.200 ;
        RECT 432.150 3.600 433.950 15.600 ;
        RECT 446.250 14.700 448.050 15.300 ;
        RECT 440.550 13.500 448.050 14.700 ;
        RECT 448.950 14.100 449.850 16.200 ;
        RECT 451.050 16.200 451.950 21.900 ;
        RECT 461.250 17.400 463.050 19.200 ;
        RECT 457.950 16.200 462.150 17.400 ;
        RECT 451.050 15.300 457.050 16.200 ;
        RECT 457.950 15.300 460.050 16.200 ;
        RECT 464.250 15.600 465.450 22.950 ;
        RECT 479.100 21.900 479.850 26.100 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 497.100 21.900 497.850 26.100 ;
        RECT 499.950 22.950 502.050 25.050 ;
        RECT 512.400 23.100 513.600 32.400 ;
        RECT 528.000 28.200 529.800 35.400 ;
        RECT 546.000 28.200 547.800 35.400 ;
        RECT 514.950 27.450 517.050 28.050 ;
        RECT 514.950 26.550 522.450 27.450 ;
        RECT 528.000 27.300 531.600 28.200 ;
        RECT 546.000 27.300 549.600 28.200 ;
        RECT 514.950 25.950 517.050 26.550 ;
        RECT 515.100 24.150 516.900 24.900 ;
        RECT 521.550 22.050 522.450 26.550 ;
        RECT 530.400 23.100 531.600 27.300 ;
        RECT 548.400 23.100 549.600 27.300 ;
        RECT 566.100 27.000 567.900 35.400 ;
        RECT 583.800 29.400 585.600 35.400 ;
        RECT 563.700 25.350 567.900 27.000 ;
        RECT 584.400 27.300 585.600 29.400 ;
        RECT 586.800 30.300 588.600 35.400 ;
        RECT 592.800 30.300 594.600 35.400 ;
        RECT 586.800 28.950 594.600 30.300 ;
        RECT 604.500 29.400 606.300 35.400 ;
        RECT 610.800 32.400 612.600 35.400 ;
        RECT 584.400 26.250 588.150 27.300 ;
        RECT 586.950 26.100 588.150 26.250 ;
        RECT 604.800 26.100 606.000 29.400 ;
        RECT 610.800 28.500 612.000 32.400 ;
        RECT 624.300 31.200 626.100 35.400 ;
        RECT 606.900 27.600 612.000 28.500 ;
        RECT 624.150 29.400 626.100 31.200 ;
        RECT 606.900 26.700 608.850 27.600 ;
        RECT 607.950 26.100 608.850 26.700 ;
        RECT 624.150 26.100 625.050 29.400 ;
        RECT 626.100 27.900 627.900 28.500 ;
        RECT 631.800 27.900 633.600 35.400 ;
        RECT 646.200 28.200 648.000 35.400 ;
        RECT 664.200 28.200 666.000 35.400 ;
        RECT 626.100 26.700 633.600 27.900 ;
        RECT 644.400 27.300 648.000 28.200 ;
        RECT 475.800 15.600 477.000 21.900 ;
        RECT 478.950 18.300 479.850 21.900 ;
        RECT 482.100 21.150 483.900 21.900 ;
        RECT 477.900 17.400 479.850 18.300 ;
        RECT 477.900 16.500 483.600 17.400 ;
        RECT 456.150 14.400 457.050 15.300 ;
        RECT 453.450 14.100 455.250 14.400 ;
        RECT 440.550 12.600 441.750 13.500 ;
        RECT 448.950 13.200 455.250 14.100 ;
        RECT 453.450 12.600 455.250 13.200 ;
        RECT 456.150 12.600 458.850 14.400 ;
        RECT 436.950 10.500 441.750 12.600 ;
        RECT 444.450 11.550 446.250 12.300 ;
        RECT 449.250 11.550 451.050 12.300 ;
        RECT 444.450 10.500 451.050 11.550 ;
        RECT 440.550 9.600 441.750 10.500 ;
        RECT 440.550 3.600 442.350 9.600 ;
        RECT 448.350 3.600 450.150 10.500 ;
        RECT 456.150 9.600 460.050 11.700 ;
        RECT 456.150 3.600 457.950 9.600 ;
        RECT 463.650 3.600 465.450 15.600 ;
        RECT 475.500 3.600 477.300 15.600 ;
        RECT 482.400 9.600 483.600 16.500 ;
        RECT 493.800 15.600 495.000 21.900 ;
        RECT 496.950 18.300 497.850 21.900 ;
        RECT 500.100 21.150 501.900 21.900 ;
        RECT 508.950 19.950 514.050 22.050 ;
        RECT 520.950 19.950 523.050 22.050 ;
        RECT 527.100 20.100 528.900 20.850 ;
        RECT 529.950 19.950 532.050 22.050 ;
        RECT 533.100 20.100 534.900 20.850 ;
        RECT 538.950 19.950 541.050 22.050 ;
        RECT 545.100 20.100 546.900 20.850 ;
        RECT 547.950 19.950 550.050 22.050 ;
        RECT 551.100 20.100 552.900 20.850 ;
        RECT 563.700 20.100 564.600 25.350 ;
        RECT 566.100 23.100 567.900 23.850 ;
        RECT 572.100 23.100 573.900 23.850 ;
        RECT 584.100 23.100 585.900 23.850 ;
        RECT 586.950 22.950 589.050 25.050 ;
        RECT 590.100 23.100 591.900 23.850 ;
        RECT 592.950 22.950 595.200 25.050 ;
        RECT 565.800 19.950 568.050 22.050 ;
        RECT 571.950 19.950 574.200 22.050 ;
        RECT 583.950 19.950 586.050 22.050 ;
        RECT 495.900 17.400 497.850 18.300 ;
        RECT 495.900 16.500 501.600 17.400 ;
        RECT 481.800 3.600 483.600 9.600 ;
        RECT 493.500 3.600 495.300 15.600 ;
        RECT 500.400 9.600 501.600 16.500 ;
        RECT 512.400 9.600 513.600 18.900 ;
        RECT 526.950 16.950 529.050 19.050 ;
        RECT 530.400 9.600 531.600 18.900 ;
        RECT 532.950 16.950 535.050 19.050 ;
        RECT 539.550 13.050 540.450 19.950 ;
        RECT 544.950 16.950 547.050 19.050 ;
        RECT 538.950 10.950 541.050 13.050 ;
        RECT 548.400 9.600 549.600 18.900 ;
        RECT 550.950 16.950 553.050 19.050 ;
        RECT 559.950 16.950 565.050 19.050 ;
        RECT 568.950 16.950 571.200 19.050 ;
        RECT 587.850 18.900 588.900 21.900 ;
        RECT 589.950 19.950 592.050 22.050 ;
        RECT 608.100 21.900 608.850 26.100 ;
        RECT 610.950 22.950 616.050 25.050 ;
        RECT 622.950 24.450 625.050 25.050 ;
        RECT 617.550 23.550 625.050 24.450 ;
        RECT 593.100 21.150 594.900 21.900 ;
        RECT 563.700 10.800 564.600 15.900 ;
        RECT 569.100 15.150 570.900 15.900 ;
        RECT 587.850 15.600 589.050 18.900 ;
        RECT 604.800 15.600 606.000 21.900 ;
        RECT 607.950 18.300 608.850 21.900 ;
        RECT 611.100 21.150 612.900 21.900 ;
        RECT 606.900 17.400 608.850 18.300 ;
        RECT 606.900 16.500 612.600 17.400 ;
        RECT 563.700 9.900 570.300 10.800 ;
        RECT 563.700 9.600 564.600 9.900 ;
        RECT 499.800 3.600 501.600 9.600 ;
        RECT 511.800 3.600 513.600 9.600 ;
        RECT 529.800 3.600 531.600 9.600 ;
        RECT 547.800 3.600 549.600 9.600 ;
        RECT 562.800 3.600 564.600 9.600 ;
        RECT 568.800 9.600 570.300 9.900 ;
        RECT 568.800 3.600 570.600 9.600 ;
        RECT 587.700 3.600 589.500 15.600 ;
        RECT 604.500 3.600 606.300 15.600 ;
        RECT 611.400 9.600 612.600 16.500 ;
        RECT 617.550 13.050 618.450 23.550 ;
        RECT 622.950 22.950 625.050 23.550 ;
        RECT 626.100 23.100 627.900 23.850 ;
        RECT 622.950 15.600 624.000 21.900 ;
        RECT 625.950 19.950 628.050 22.050 ;
        RECT 616.950 10.950 619.050 13.050 ;
        RECT 610.800 3.600 612.600 9.600 ;
        RECT 622.200 3.600 624.000 15.600 ;
        RECT 629.550 9.600 630.600 26.700 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 644.400 23.100 645.600 27.300 ;
        RECT 652.950 25.950 655.050 28.050 ;
        RECT 662.400 27.300 666.000 28.200 ;
        RECT 653.550 22.050 654.450 25.950 ;
        RECT 662.400 23.100 663.600 27.300 ;
        RECT 683.100 27.000 684.900 35.400 ;
        RECT 700.800 32.400 702.600 35.400 ;
        RECT 680.700 25.350 684.900 27.000 ;
        RECT 632.100 21.150 633.900 21.900 ;
        RECT 641.100 20.100 642.900 20.850 ;
        RECT 643.950 19.950 646.050 22.050 ;
        RECT 647.100 20.100 648.900 20.850 ;
        RECT 652.950 19.950 655.050 22.050 ;
        RECT 659.100 20.100 660.900 20.850 ;
        RECT 661.950 19.950 664.050 22.050 ;
        RECT 665.100 20.100 666.900 20.850 ;
        RECT 680.700 20.100 681.600 25.350 ;
        RECT 683.100 23.100 684.900 23.850 ;
        RECT 689.100 23.100 690.900 23.850 ;
        RECT 701.400 23.100 702.600 32.400 ;
        RECT 703.950 25.950 706.050 28.050 ;
        RECT 719.100 27.000 720.900 35.400 ;
        RECT 739.200 28.200 741.000 35.400 ;
        RECT 716.700 25.350 720.900 27.000 ;
        RECT 737.400 27.300 741.000 28.200 ;
        RECT 746.550 29.400 748.350 35.400 ;
        RECT 754.650 32.400 756.450 35.400 ;
        RECT 762.450 32.400 764.250 35.400 ;
        RECT 770.250 33.300 772.050 35.400 ;
        RECT 770.250 32.400 774.000 33.300 ;
        RECT 754.650 31.500 755.700 32.400 ;
        RECT 751.950 30.300 755.700 31.500 ;
        RECT 763.200 30.600 764.250 32.400 ;
        RECT 772.950 31.500 774.000 32.400 ;
        RECT 751.950 29.400 754.050 30.300 ;
        RECT 704.100 24.150 705.900 24.900 ;
        RECT 682.800 19.950 685.050 22.050 ;
        RECT 688.950 19.950 691.200 22.050 ;
        RECT 697.950 19.950 703.050 22.050 ;
        RECT 716.700 20.100 717.600 25.350 ;
        RECT 719.100 23.100 720.900 23.850 ;
        RECT 725.100 23.100 726.900 23.850 ;
        RECT 737.400 23.100 738.600 27.300 ;
        RECT 746.550 25.050 747.750 29.400 ;
        RECT 759.150 28.200 760.950 30.000 ;
        RECT 763.200 29.550 768.150 30.600 ;
        RECT 766.350 28.800 768.150 29.550 ;
        RECT 769.650 28.800 771.450 30.600 ;
        RECT 772.950 29.400 775.050 31.500 ;
        RECT 778.050 29.400 779.850 35.400 ;
        RECT 793.200 31.050 795.000 35.400 ;
        RECT 802.950 31.950 805.050 34.050 ;
        RECT 793.200 29.400 798.600 31.050 ;
        RECT 760.050 27.900 760.950 28.200 ;
        RECT 770.100 27.900 771.150 28.800 ;
        RECT 760.050 27.000 771.150 27.900 ;
        RECT 760.050 26.100 760.950 27.000 ;
        RECT 770.100 25.800 771.150 27.000 ;
        RECT 746.550 22.950 747.900 25.050 ;
        RECT 748.950 22.950 751.050 25.050 ;
        RECT 752.100 23.250 752.850 25.050 ;
        RECT 760.950 22.950 763.050 25.050 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 770.100 24.600 777.000 25.800 ;
        RECT 770.100 24.000 771.900 24.600 ;
        RECT 776.100 23.850 777.000 24.600 ;
        RECT 773.100 23.100 774.900 23.700 ;
        RECT 718.950 19.950 721.050 22.050 ;
        RECT 724.950 19.950 727.050 22.050 ;
        RECT 734.100 20.100 735.900 20.850 ;
        RECT 736.950 19.950 739.050 22.050 ;
        RECT 740.100 20.100 741.900 20.850 ;
        RECT 640.950 16.950 643.050 19.050 ;
        RECT 628.800 3.600 630.600 9.600 ;
        RECT 644.400 9.600 645.600 18.900 ;
        RECT 646.950 16.950 649.050 19.050 ;
        RECT 658.950 16.950 661.050 19.050 ;
        RECT 662.400 9.600 663.600 18.900 ;
        RECT 664.950 16.950 667.050 19.050 ;
        RECT 679.950 18.450 682.050 19.050 ;
        RECT 674.550 18.000 682.050 18.450 ;
        RECT 673.950 17.550 682.050 18.000 ;
        RECT 673.950 13.950 676.050 17.550 ;
        RECT 679.950 16.950 682.050 17.550 ;
        RECT 685.950 16.950 688.050 19.050 ;
        RECT 680.700 10.800 681.600 15.900 ;
        RECT 686.100 15.150 687.900 15.900 ;
        RECT 680.700 9.900 687.300 10.800 ;
        RECT 680.700 9.600 681.600 9.900 ;
        RECT 644.400 3.600 646.200 9.600 ;
        RECT 662.400 3.600 664.200 9.600 ;
        RECT 679.800 3.600 681.600 9.600 ;
        RECT 685.800 9.600 687.300 9.900 ;
        RECT 701.400 9.600 702.600 18.900 ;
        RECT 715.950 18.450 718.050 19.050 ;
        RECT 710.550 17.550 718.050 18.450 ;
        RECT 710.550 13.050 711.450 17.550 ;
        RECT 715.950 16.950 718.050 17.550 ;
        RECT 721.950 16.950 724.050 19.050 ;
        RECT 733.950 16.950 736.050 19.050 ;
        RECT 709.950 10.950 712.050 13.050 ;
        RECT 716.700 10.800 717.600 15.900 ;
        RECT 722.100 15.150 723.900 15.900 ;
        RECT 716.700 9.900 723.300 10.800 ;
        RECT 716.700 9.600 717.600 9.900 ;
        RECT 685.800 3.600 687.600 9.600 ;
        RECT 700.800 3.600 702.600 9.600 ;
        RECT 715.800 3.600 717.600 9.600 ;
        RECT 721.800 9.600 723.300 9.900 ;
        RECT 737.400 9.600 738.600 18.900 ;
        RECT 739.950 16.950 742.050 19.050 ;
        RECT 746.550 15.600 747.750 22.950 ;
        RECT 770.100 22.200 774.900 23.100 ;
        RECT 773.100 21.900 774.900 22.200 ;
        RECT 776.100 22.050 777.900 23.850 ;
        RECT 748.950 17.400 750.750 19.200 ;
        RECT 749.850 16.200 754.050 17.400 ;
        RECT 760.050 16.200 760.950 21.900 ;
        RECT 768.750 17.100 770.550 17.400 ;
        RECT 721.800 3.600 723.600 9.600 ;
        RECT 737.400 3.600 739.200 9.600 ;
        RECT 746.550 3.600 748.350 15.600 ;
        RECT 751.950 15.300 754.050 16.200 ;
        RECT 754.950 15.300 760.950 16.200 ;
        RECT 762.150 16.800 770.550 17.100 ;
        RECT 778.950 16.800 779.850 29.400 ;
        RECT 797.700 26.100 798.600 29.400 ;
        RECT 788.100 23.100 789.900 23.850 ;
        RECT 790.950 22.950 793.050 25.050 ;
        RECT 796.950 24.450 799.050 25.050 ;
        RECT 803.550 24.450 804.450 31.950 ;
        RECT 809.400 30.300 811.200 35.400 ;
        RECT 815.400 30.300 817.200 35.400 ;
        RECT 809.400 28.950 817.200 30.300 ;
        RECT 818.400 29.400 820.200 35.400 ;
        RECT 830.400 32.400 832.200 35.400 ;
        RECT 818.400 27.300 819.600 29.400 ;
        RECT 823.950 28.950 826.050 31.050 ;
        RECT 815.850 26.250 819.600 27.300 ;
        RECT 815.850 26.100 817.050 26.250 ;
        RECT 794.100 23.100 795.900 23.850 ;
        RECT 796.950 23.550 804.450 24.450 ;
        RECT 796.950 22.950 799.050 23.550 ;
        RECT 808.950 22.950 811.050 25.050 ;
        RECT 812.100 23.100 813.900 23.850 ;
        RECT 814.950 22.950 817.050 25.050 ;
        RECT 824.550 24.450 825.450 28.950 ;
        RECT 831.000 28.500 832.200 32.400 ;
        RECT 836.700 29.400 838.500 35.400 ;
        RECT 851.400 32.400 853.200 35.400 ;
        RECT 831.000 27.600 836.100 28.500 ;
        RECT 834.150 26.700 836.100 27.600 ;
        RECT 834.150 26.100 835.050 26.700 ;
        RECT 837.000 26.100 838.200 29.400 ;
        RECT 829.950 24.450 832.050 25.050 ;
        RECT 818.100 23.100 819.900 23.850 ;
        RECT 824.550 23.550 832.050 24.450 ;
        RECT 829.950 22.950 832.050 23.550 ;
        RECT 787.950 19.950 790.050 22.050 ;
        RECT 791.100 21.150 792.900 21.900 ;
        RECT 793.950 19.950 796.050 22.050 ;
        RECT 762.150 16.200 779.850 16.800 ;
        RECT 754.950 14.400 755.850 15.300 ;
        RECT 753.150 12.600 755.850 14.400 ;
        RECT 756.750 14.100 758.550 14.400 ;
        RECT 762.150 14.100 763.050 16.200 ;
        RECT 768.750 15.600 779.850 16.200 ;
        RECT 797.700 15.600 798.600 21.900 ;
        RECT 809.100 21.150 810.900 21.900 ;
        RECT 811.950 19.950 814.050 22.050 ;
        RECT 815.100 18.900 816.150 21.900 ;
        RECT 817.950 19.950 820.050 22.050 ;
        RECT 834.150 21.900 834.900 26.100 ;
        RECT 847.950 25.950 850.050 28.050 ;
        RECT 835.950 22.950 838.050 25.050 ;
        RECT 848.100 24.150 849.900 24.900 ;
        RECT 851.400 23.100 852.600 32.400 ;
        RECT 830.100 21.150 831.900 21.900 ;
        RECT 814.950 15.600 816.150 18.900 ;
        RECT 834.150 18.300 835.050 21.900 ;
        RECT 834.150 17.400 836.100 18.300 ;
        RECT 830.400 16.500 836.100 17.400 ;
        RECT 756.750 13.200 763.050 14.100 ;
        RECT 763.950 14.700 765.750 15.300 ;
        RECT 763.950 13.500 771.450 14.700 ;
        RECT 756.750 12.600 758.550 13.200 ;
        RECT 770.250 12.600 771.450 13.500 ;
        RECT 751.950 9.600 755.850 11.700 ;
        RECT 760.950 11.550 762.750 12.300 ;
        RECT 765.750 11.550 767.550 12.300 ;
        RECT 760.950 10.500 767.550 11.550 ;
        RECT 770.250 10.500 775.050 12.600 ;
        RECT 754.050 3.600 755.850 9.600 ;
        RECT 761.850 3.600 763.650 10.500 ;
        RECT 770.250 9.600 771.450 10.500 ;
        RECT 769.650 3.600 771.450 9.600 ;
        RECT 778.050 3.600 779.850 15.600 ;
        RECT 788.400 14.700 796.200 15.600 ;
        RECT 788.400 3.600 790.200 14.700 ;
        RECT 794.400 3.600 796.200 14.700 ;
        RECT 797.400 3.600 799.200 15.600 ;
        RECT 814.500 3.600 816.300 15.600 ;
        RECT 830.400 9.600 831.600 16.500 ;
        RECT 837.000 15.600 838.200 21.900 ;
        RECT 847.950 19.950 853.050 22.050 ;
        RECT 830.400 3.600 832.200 9.600 ;
        RECT 836.700 3.600 838.500 15.600 ;
        RECT 851.400 9.600 852.600 18.900 ;
        RECT 851.400 3.600 853.200 9.600 ;
      LAYER metal2 ;
        RECT 640.950 867.450 643.050 868.050 ;
        RECT 718.950 867.450 721.050 868.050 ;
        RECT 640.950 866.400 721.050 867.450 ;
        RECT 640.950 865.950 643.050 866.400 ;
        RECT 718.950 865.950 721.050 866.400 ;
        RECT 739.950 867.450 742.050 868.050 ;
        RECT 814.950 867.450 817.050 868.050 ;
        RECT 739.950 866.400 817.050 867.450 ;
        RECT 739.950 865.950 742.050 866.400 ;
        RECT 814.950 865.950 817.050 866.400 ;
        RECT 601.950 864.450 604.050 865.050 ;
        RECT 634.950 864.450 637.050 865.050 ;
        RECT 601.950 863.400 637.050 864.450 ;
        RECT 601.950 862.950 604.050 863.400 ;
        RECT 634.950 862.950 637.050 863.400 ;
        RECT 184.950 861.450 187.050 862.050 ;
        RECT 226.950 861.450 229.050 862.050 ;
        RECT 283.950 861.450 286.050 862.050 ;
        RECT 184.950 860.400 286.050 861.450 ;
        RECT 184.950 859.950 187.050 860.400 ;
        RECT 226.950 859.950 229.050 860.400 ;
        RECT 283.950 859.950 286.050 860.400 ;
        RECT 88.950 858.450 91.050 859.050 ;
        RECT 196.950 858.450 199.050 859.050 ;
        RECT 88.950 857.400 199.050 858.450 ;
        RECT 88.950 856.950 91.050 857.400 ;
        RECT 196.950 856.950 199.050 857.400 ;
        RECT 583.950 857.100 586.050 859.200 ;
        RECT 91.950 855.450 94.050 856.050 ;
        RECT 316.950 855.450 319.050 856.050 ;
        RECT 91.950 854.400 319.050 855.450 ;
        RECT 91.950 853.950 94.050 854.400 ;
        RECT 316.950 853.950 319.050 854.400 ;
        RECT 343.950 855.450 346.050 856.050 ;
        RECT 439.950 855.450 442.050 856.050 ;
        RECT 343.950 854.400 442.050 855.450 ;
        RECT 343.950 853.950 346.050 854.400 ;
        RECT 439.950 853.950 442.050 854.400 ;
        RECT 584.550 853.350 585.750 857.100 ;
        RECT 586.950 855.300 589.050 857.400 ;
        RECT 589.950 855.300 592.050 857.400 ;
        RECT 593.850 855.300 595.950 857.400 ;
        RECT 607.950 856.950 610.050 859.050 ;
        RECT 610.950 856.950 613.050 859.050 ;
        RECT 613.950 856.950 616.050 859.050 ;
        RECT 673.950 857.100 676.050 859.200 ;
        RECT 46.950 852.450 49.050 853.050 ;
        RECT 124.950 852.450 127.050 853.050 ;
        RECT 17.400 852.000 127.050 852.450 ;
        RECT 16.950 851.400 127.050 852.000 ;
        RECT 16.950 847.950 19.050 851.400 ;
        RECT 31.950 847.950 34.050 851.400 ;
        RECT 46.950 850.950 49.050 851.400 ;
        RECT 124.950 850.950 127.050 851.400 ;
        RECT 130.950 852.450 133.050 853.050 ;
        RECT 151.950 852.450 154.050 853.050 ;
        RECT 130.950 851.400 154.050 852.450 ;
        RECT 130.950 850.950 133.050 851.400 ;
        RECT 151.950 850.950 154.050 851.400 ;
        RECT 241.950 852.450 244.050 853.050 ;
        RECT 256.950 852.450 259.050 853.050 ;
        RECT 265.950 852.450 268.050 853.050 ;
        RECT 241.950 851.400 268.050 852.450 ;
        RECT 241.950 850.950 244.050 851.400 ;
        RECT 256.950 850.950 259.050 851.400 ;
        RECT 265.950 850.950 268.050 851.400 ;
        RECT 319.950 852.450 322.050 853.050 ;
        RECT 421.950 852.450 424.050 853.050 ;
        RECT 319.950 851.400 424.050 852.450 ;
        RECT 319.950 850.950 322.050 851.400 ;
        RECT 421.950 850.950 424.050 851.400 ;
        RECT 118.950 849.450 121.050 850.050 ;
        RECT 136.950 849.450 142.050 850.050 ;
        RECT 118.950 848.400 142.050 849.450 ;
        RECT 118.950 847.950 121.050 848.400 ;
        RECT 136.950 847.950 142.050 848.400 ;
        RECT 7.950 846.450 10.050 847.050 ;
        RECT 13.950 846.450 16.050 847.050 ;
        RECT 7.950 845.400 16.050 846.450 ;
        RECT 7.950 844.950 10.050 845.400 ;
        RECT 13.950 844.950 16.050 845.400 ;
        RECT 19.950 846.450 22.050 847.050 ;
        RECT 28.950 846.450 31.050 847.050 ;
        RECT 19.950 845.400 31.050 846.450 ;
        RECT 19.950 844.950 22.050 845.400 ;
        RECT 28.950 841.950 31.050 845.400 ;
        RECT 34.950 841.950 37.050 847.050 ;
        RECT 46.950 844.950 52.050 847.050 ;
        RECT 55.950 844.950 61.050 847.050 ;
        RECT 73.800 846.450 75.900 847.050 ;
        RECT 68.400 845.400 75.900 846.450 ;
        RECT 49.950 841.950 55.050 844.050 ;
        RECT 61.950 843.450 64.050 844.050 ;
        RECT 68.400 843.450 69.450 845.400 ;
        RECT 73.800 844.950 75.900 845.400 ;
        RECT 77.100 844.950 82.050 847.050 ;
        RECT 94.950 844.050 97.050 847.050 ;
        RECT 100.950 846.450 103.050 847.050 ;
        RECT 112.950 846.450 115.050 847.050 ;
        RECT 130.800 846.450 132.900 847.050 ;
        RECT 100.950 845.400 132.900 846.450 ;
        RECT 134.100 846.000 136.200 847.050 ;
        RECT 100.950 844.950 103.050 845.400 ;
        RECT 112.950 844.950 115.050 845.400 ;
        RECT 130.800 844.950 132.900 845.400 ;
        RECT 133.950 844.950 136.200 846.000 ;
        RECT 139.950 844.950 145.050 847.050 ;
        RECT 151.950 844.950 154.050 850.050 ;
        RECT 208.950 847.950 214.050 850.050 ;
        RECT 217.950 847.950 223.050 850.050 ;
        RECT 225.000 849.450 229.050 850.050 ;
        RECT 224.400 847.950 229.050 849.450 ;
        RECT 232.950 847.950 238.050 850.050 ;
        RECT 358.950 849.450 361.050 850.050 ;
        RECT 376.950 849.450 379.050 850.050 ;
        RECT 412.950 849.450 415.050 850.050 ;
        RECT 257.400 849.000 291.450 849.450 ;
        RECT 256.950 848.400 291.450 849.000 ;
        RECT 157.950 844.950 163.050 847.050 ;
        RECT 166.950 844.950 172.050 847.050 ;
        RECT 175.950 844.950 181.050 847.050 ;
        RECT 196.950 846.450 199.050 847.050 ;
        RECT 205.950 846.450 208.050 847.050 ;
        RECT 196.950 845.400 208.050 846.450 ;
        RECT 196.950 844.950 199.050 845.400 ;
        RECT 205.950 844.950 208.050 845.400 ;
        RECT 211.950 846.450 214.050 847.050 ;
        RECT 224.400 846.450 225.450 847.950 ;
        RECT 211.950 845.400 225.450 846.450 ;
        RECT 226.950 846.450 229.050 847.050 ;
        RECT 232.950 846.450 235.050 847.050 ;
        RECT 226.950 845.400 235.050 846.450 ;
        RECT 211.950 844.950 214.050 845.400 ;
        RECT 226.950 844.950 229.050 845.400 ;
        RECT 232.950 844.950 235.050 845.400 ;
        RECT 238.950 844.950 243.900 847.050 ;
        RECT 245.100 846.450 247.200 847.050 ;
        RECT 250.950 846.450 253.050 847.050 ;
        RECT 245.100 845.400 253.050 846.450 ;
        RECT 245.100 844.950 247.200 845.400 ;
        RECT 250.950 844.950 253.050 845.400 ;
        RECT 256.950 844.950 259.050 848.400 ;
        RECT 283.950 844.950 289.050 847.050 ;
        RECT 290.400 846.450 291.450 848.400 ;
        RECT 358.950 849.000 369.600 849.450 ;
        RECT 358.950 848.400 370.050 849.000 ;
        RECT 358.950 847.950 361.050 848.400 ;
        RECT 367.950 847.050 370.050 848.400 ;
        RECT 376.950 848.400 415.050 849.450 ;
        RECT 376.950 847.950 379.050 848.400 ;
        RECT 292.950 846.450 295.050 847.050 ;
        RECT 304.950 846.450 307.050 847.050 ;
        RECT 319.800 846.450 321.900 847.050 ;
        RECT 290.400 845.400 321.900 846.450 ;
        RECT 292.950 844.950 295.050 845.400 ;
        RECT 304.950 844.950 307.050 845.400 ;
        RECT 319.800 844.950 321.900 845.400 ;
        RECT 323.100 846.450 325.200 847.050 ;
        RECT 337.950 846.450 340.050 847.050 ;
        RECT 323.100 845.400 340.050 846.450 ;
        RECT 323.100 844.950 325.200 845.400 ;
        RECT 337.950 844.950 340.050 845.400 ;
        RECT 133.950 844.050 136.050 844.950 ;
        RECT 61.950 842.400 69.450 843.450 ;
        RECT 61.950 841.950 64.050 842.400 ;
        RECT 70.950 841.950 75.900 844.050 ;
        RECT 77.100 843.450 79.200 844.050 ;
        RECT 91.800 843.450 93.900 844.050 ;
        RECT 77.100 842.400 93.900 843.450 ;
        RECT 94.950 843.000 97.200 844.050 ;
        RECT 98.100 843.000 100.200 844.050 ;
        RECT 77.100 841.950 79.200 842.400 ;
        RECT 91.800 841.950 93.900 842.400 ;
        RECT 95.100 841.950 97.200 843.000 ;
        RECT 97.950 841.950 100.200 843.000 ;
        RECT 43.950 840.450 46.050 841.050 ;
        RECT 76.950 840.450 79.050 841.050 ;
        RECT 43.950 839.400 79.050 840.450 ;
        RECT 43.950 838.950 46.050 839.400 ;
        RECT 76.950 838.950 79.050 839.400 ;
        RECT 82.950 840.450 85.050 841.050 ;
        RECT 97.950 840.450 100.050 841.950 ;
        RECT 82.950 840.000 100.050 840.450 ;
        RECT 82.950 839.400 99.450 840.000 ;
        RECT 82.950 838.950 85.050 839.400 ;
        RECT 103.950 838.950 106.050 844.050 ;
        RECT 118.950 838.950 121.050 844.050 ;
        RECT 133.950 843.000 136.200 844.050 ;
        RECT 134.100 841.950 136.200 843.000 ;
        RECT 148.950 838.950 151.050 844.050 ;
        RECT 154.950 840.450 157.050 844.050 ;
        RECT 172.950 843.450 175.050 844.050 ;
        RECT 193.950 843.450 196.050 844.050 ;
        RECT 172.950 842.400 196.050 843.450 ;
        RECT 172.950 841.950 175.050 842.400 ;
        RECT 193.950 841.950 196.050 842.400 ;
        RECT 247.950 843.450 250.050 844.050 ;
        RECT 253.950 843.450 256.050 844.050 ;
        RECT 247.950 842.400 256.050 843.450 ;
        RECT 247.950 841.950 250.050 842.400 ;
        RECT 253.950 841.950 256.050 842.400 ;
        RECT 181.950 840.450 184.050 841.050 ;
        RECT 154.950 840.000 184.050 840.450 ;
        RECT 155.400 839.400 184.050 840.000 ;
        RECT 181.950 838.950 184.050 839.400 ;
        RECT 196.950 840.450 199.050 841.050 ;
        RECT 214.950 840.450 217.050 841.050 ;
        RECT 196.950 839.400 217.050 840.450 ;
        RECT 259.950 840.450 262.050 844.050 ;
        RECT 274.950 840.450 277.050 841.050 ;
        RECT 259.950 840.000 277.050 840.450 ;
        RECT 260.400 839.400 277.050 840.000 ;
        RECT 196.950 838.950 199.050 839.400 ;
        RECT 214.950 838.950 217.050 839.400 ;
        RECT 34.950 837.450 37.050 838.050 ;
        RECT 58.950 837.450 61.050 838.050 ;
        RECT 34.950 836.400 61.050 837.450 ;
        RECT 34.950 835.950 37.050 836.400 ;
        RECT 58.950 835.950 61.050 836.400 ;
        RECT 133.950 837.450 136.050 838.050 ;
        RECT 169.950 837.450 172.050 838.050 ;
        RECT 133.950 836.400 172.050 837.450 ;
        RECT 133.950 835.950 136.050 836.400 ;
        RECT 169.950 835.950 172.050 836.400 ;
        RECT 211.950 837.450 214.050 838.050 ;
        RECT 247.950 837.450 250.050 838.050 ;
        RECT 211.950 836.400 250.050 837.450 ;
        RECT 274.950 837.450 277.050 839.400 ;
        RECT 289.950 838.950 292.050 844.050 ;
        RECT 295.950 841.950 301.050 844.050 ;
        RECT 328.950 841.050 331.050 844.050 ;
        RECT 343.950 841.950 346.050 847.050 ;
        RECT 361.950 844.950 366.900 847.050 ;
        RECT 367.950 846.000 370.200 847.050 ;
        RECT 368.100 844.950 370.200 846.000 ;
        RECT 373.950 846.450 376.050 847.050 ;
        RECT 385.950 846.450 388.050 847.050 ;
        RECT 373.950 846.000 396.450 846.450 ;
        RECT 373.950 845.400 397.050 846.000 ;
        RECT 373.950 844.950 376.050 845.400 ;
        RECT 385.950 844.950 388.050 845.400 ;
        RECT 349.950 841.950 355.050 844.050 ;
        RECT 304.950 840.450 307.050 841.050 ;
        RECT 328.800 840.450 331.050 841.050 ;
        RECT 304.950 840.000 331.050 840.450 ;
        RECT 332.100 840.450 334.200 841.050 ;
        RECT 343.800 840.450 345.900 841.050 ;
        RECT 304.950 839.400 330.900 840.000 ;
        RECT 304.950 838.950 307.050 839.400 ;
        RECT 328.800 838.950 330.900 839.400 ;
        RECT 332.100 839.400 345.900 840.450 ;
        RECT 332.100 838.950 334.200 839.400 ;
        RECT 343.800 838.950 345.900 839.400 ;
        RECT 347.100 840.450 349.200 841.050 ;
        RECT 358.950 840.450 361.050 841.050 ;
        RECT 347.100 839.400 361.050 840.450 ;
        RECT 347.100 838.950 349.200 839.400 ;
        RECT 358.950 838.950 361.050 839.400 ;
        RECT 364.950 838.950 367.050 844.050 ;
        RECT 370.950 843.450 373.050 844.050 ;
        RECT 376.950 843.450 379.050 844.050 ;
        RECT 370.950 842.400 379.050 843.450 ;
        RECT 370.950 841.950 373.050 842.400 ;
        RECT 376.950 841.950 379.050 842.400 ;
        RECT 394.950 841.950 397.050 845.400 ;
        RECT 397.950 844.950 400.050 848.400 ;
        RECT 412.950 847.950 415.050 848.400 ;
        RECT 433.950 847.950 439.050 850.050 ;
        RECT 442.950 849.450 445.050 850.050 ;
        RECT 448.950 849.450 451.050 850.050 ;
        RECT 442.950 848.400 451.050 849.450 ;
        RECT 442.950 847.950 445.050 848.400 ;
        RECT 448.950 847.950 451.050 848.400 ;
        RECT 484.950 847.950 487.050 853.050 ;
        RECT 559.950 852.450 562.050 853.050 ;
        RECT 574.950 852.450 577.050 853.050 ;
        RECT 559.950 851.400 577.050 852.450 ;
        RECT 559.950 850.950 562.050 851.400 ;
        RECT 574.950 850.950 577.050 851.400 ;
        RECT 583.950 851.250 586.050 853.350 ;
        RECT 511.950 847.950 517.050 850.050 ;
        RECT 520.950 849.450 523.050 850.050 ;
        RECT 526.950 849.450 529.050 850.050 ;
        RECT 520.950 848.400 529.050 849.450 ;
        RECT 520.950 847.950 523.050 848.400 ;
        RECT 526.950 847.950 529.050 848.400 ;
        RECT 403.950 844.950 409.050 847.050 ;
        RECT 418.950 844.950 424.050 847.050 ;
        RECT 427.950 844.950 433.050 847.050 ;
        RECT 439.950 844.950 445.050 847.050 ;
        RECT 466.950 846.450 469.050 847.050 ;
        RECT 475.950 846.450 478.050 847.050 ;
        RECT 466.950 845.400 478.050 846.450 ;
        RECT 466.950 844.950 469.050 845.400 ;
        RECT 475.950 844.950 478.050 845.400 ;
        RECT 400.950 841.950 406.050 844.050 ;
        RECT 385.950 840.450 388.050 841.050 ;
        RECT 412.950 840.450 415.050 841.050 ;
        RECT 385.950 839.400 415.050 840.450 ;
        RECT 424.950 840.450 427.050 844.050 ;
        RECT 457.950 843.450 460.050 844.050 ;
        RECT 469.950 843.450 472.050 844.050 ;
        RECT 457.950 842.400 472.050 843.450 ;
        RECT 481.950 843.450 484.050 847.050 ;
        RECT 487.950 846.450 490.050 847.050 ;
        RECT 496.950 846.450 499.050 847.050 ;
        RECT 487.950 845.400 499.050 846.450 ;
        RECT 487.950 844.950 490.050 845.400 ;
        RECT 496.950 844.950 499.050 845.400 ;
        RECT 517.950 846.450 520.050 847.050 ;
        RECT 526.950 846.450 529.050 847.050 ;
        RECT 517.950 845.400 529.050 846.450 ;
        RECT 517.950 844.950 520.050 845.400 ;
        RECT 526.950 844.950 529.050 845.400 ;
        RECT 562.950 844.950 565.050 847.050 ;
        RECT 566.250 844.950 567.150 847.050 ;
        RECT 572.850 844.950 573.750 847.050 ;
        RECT 574.950 844.950 577.050 847.050 ;
        RECT 511.950 843.450 514.050 844.050 ;
        RECT 481.950 843.000 514.050 843.450 ;
        RECT 482.400 842.400 514.050 843.000 ;
        RECT 457.950 841.950 460.050 842.400 ;
        RECT 469.950 841.950 472.050 842.400 ;
        RECT 511.950 841.950 514.050 842.400 ;
        RECT 436.950 840.450 439.050 841.050 ;
        RECT 454.950 840.450 457.050 841.050 ;
        RECT 472.950 840.450 475.050 841.050 ;
        RECT 424.950 840.000 475.050 840.450 ;
        RECT 425.400 839.400 475.050 840.000 ;
        RECT 385.950 838.950 388.050 839.400 ;
        RECT 412.950 838.950 415.050 839.400 ;
        RECT 436.950 838.950 439.050 839.400 ;
        RECT 454.950 838.950 457.050 839.400 ;
        RECT 472.950 838.950 475.050 839.400 ;
        RECT 502.950 840.450 505.050 841.050 ;
        RECT 568.950 840.450 571.050 841.050 ;
        RECT 502.950 839.400 571.050 840.450 ;
        RECT 502.950 838.950 505.050 839.400 ;
        RECT 568.950 838.950 571.050 839.400 ;
        RECT 295.950 837.450 298.050 838.050 ;
        RECT 274.950 837.000 298.050 837.450 ;
        RECT 275.400 836.400 298.050 837.000 ;
        RECT 211.950 835.950 214.050 836.400 ;
        RECT 247.950 835.950 250.050 836.400 ;
        RECT 295.950 835.950 298.050 836.400 ;
        RECT 328.950 837.450 331.050 838.050 ;
        RECT 349.950 837.450 352.050 838.050 ;
        RECT 328.950 836.400 352.050 837.450 ;
        RECT 328.950 835.950 331.050 836.400 ;
        RECT 349.950 835.950 352.050 836.400 ;
        RECT 427.950 837.450 430.050 838.050 ;
        RECT 448.950 837.450 451.050 838.050 ;
        RECT 517.950 837.450 520.050 838.050 ;
        RECT 427.950 836.400 520.050 837.450 ;
        RECT 427.950 835.950 430.050 836.400 ;
        RECT 448.950 835.950 451.050 836.400 ;
        RECT 517.950 835.950 520.050 836.400 ;
        RECT 553.950 837.450 556.050 838.050 ;
        RECT 562.950 837.450 565.050 838.050 ;
        RECT 584.550 837.600 585.750 851.250 ;
        RECT 586.950 837.600 588.150 855.300 ;
        RECT 589.950 853.350 591.150 855.300 ;
        RECT 589.950 851.250 592.050 853.350 ;
        RECT 589.950 837.600 591.450 851.250 ;
        RECT 593.850 845.550 595.050 855.300 ;
        RECT 598.950 854.400 601.050 856.500 ;
        RECT 599.850 848.250 601.050 854.400 ;
        RECT 598.950 846.150 601.050 848.250 ;
        RECT 593.850 843.450 596.850 845.550 ;
        RECT 593.850 837.600 595.050 843.450 ;
        RECT 599.850 842.250 601.050 846.150 ;
        RECT 601.950 842.250 604.050 843.150 ;
        RECT 599.850 837.750 600.750 842.250 ;
        RECT 601.950 838.950 604.050 841.050 ;
        RECT 607.950 838.050 609.150 856.950 ;
        RECT 610.950 852.750 612.150 856.950 ;
        RECT 610.950 850.650 613.050 852.750 ;
        RECT 610.950 838.050 612.150 850.650 ;
        RECT 613.950 838.050 615.150 856.950 ;
        RECT 674.550 853.350 675.750 857.100 ;
        RECT 676.950 855.300 679.050 857.400 ;
        RECT 679.950 855.300 682.050 857.400 ;
        RECT 683.850 855.300 685.950 857.400 ;
        RECT 697.950 856.950 700.050 859.050 ;
        RECT 700.950 856.950 703.050 859.050 ;
        RECT 703.950 856.950 706.050 859.050 ;
        RECT 640.800 852.000 642.900 853.050 ;
        RECT 640.800 850.950 643.050 852.000 ;
        RECT 673.950 851.250 676.050 853.350 ;
        RECT 640.950 850.050 643.050 850.950 ;
        RECT 619.950 848.250 622.050 849.150 ;
        RECT 640.800 849.000 643.050 850.050 ;
        RECT 640.800 847.950 642.900 849.000 ;
        RECT 644.100 847.950 649.050 850.050 ;
        RECT 619.950 844.950 622.050 847.050 ;
        RECT 625.950 845.850 628.050 846.750 ;
        RECT 634.950 846.450 637.050 847.050 ;
        RECT 643.950 846.450 646.050 847.050 ;
        RECT 634.950 845.400 646.050 846.450 ;
        RECT 634.950 844.950 637.050 845.400 ;
        RECT 643.950 844.950 646.050 845.400 ;
        RECT 649.950 844.950 655.050 847.050 ;
        RECT 656.250 844.950 657.150 847.050 ;
        RECT 662.850 844.950 663.750 847.050 ;
        RECT 664.950 844.950 667.050 847.050 ;
        RECT 620.400 840.450 621.450 844.950 ;
        RECT 631.950 840.450 634.050 841.050 ;
        RECT 620.400 839.400 634.050 840.450 ;
        RECT 631.950 838.950 634.050 839.400 ;
        RECT 599.850 837.600 601.050 837.750 ;
        RECT 553.950 836.400 565.050 837.450 ;
        RECT 553.950 835.950 556.050 836.400 ;
        RECT 562.950 835.950 565.050 836.400 ;
        RECT 583.950 835.500 586.050 837.600 ;
        RECT 586.950 835.500 589.050 837.600 ;
        RECT 589.950 835.500 592.050 837.600 ;
        RECT 593.850 835.500 595.950 837.600 ;
        RECT 598.950 835.500 601.050 837.600 ;
        RECT 607.950 835.950 610.050 838.050 ;
        RECT 610.950 835.950 613.050 838.050 ;
        RECT 613.950 835.950 616.050 838.050 ;
        RECT 674.550 837.600 675.750 851.250 ;
        RECT 676.950 837.600 678.150 855.300 ;
        RECT 679.950 853.350 681.150 855.300 ;
        RECT 679.950 851.250 682.050 853.350 ;
        RECT 679.950 837.600 681.450 851.250 ;
        RECT 683.850 845.550 685.050 855.300 ;
        RECT 688.950 854.400 691.050 856.500 ;
        RECT 689.850 848.250 691.050 854.400 ;
        RECT 688.950 846.150 691.050 848.250 ;
        RECT 683.850 843.450 686.850 845.550 ;
        RECT 683.850 837.600 685.050 843.450 ;
        RECT 689.850 842.250 691.050 846.150 ;
        RECT 691.950 842.250 694.050 843.150 ;
        RECT 689.850 837.750 690.750 842.250 ;
        RECT 691.950 838.950 694.050 841.050 ;
        RECT 697.950 838.050 699.150 856.950 ;
        RECT 700.950 852.750 702.150 856.950 ;
        RECT 700.950 850.650 703.050 852.750 ;
        RECT 700.950 838.050 702.150 850.650 ;
        RECT 703.950 838.050 705.150 856.950 ;
        RECT 796.950 855.300 799.050 857.400 ;
        RECT 797.850 851.700 799.050 855.300 ;
        RECT 817.950 854.400 820.050 856.500 ;
        RECT 709.950 848.250 712.050 849.150 ;
        RECT 715.950 847.950 718.050 850.050 ;
        RECT 760.950 849.450 763.050 850.050 ;
        RECT 796.950 849.600 799.050 851.700 ;
        RECT 737.250 849.000 763.050 849.450 ;
        RECT 736.950 848.400 763.050 849.000 ;
        RECT 736.950 847.050 739.050 848.400 ;
        RECT 760.950 847.950 763.050 848.400 ;
        RECT 715.950 845.850 718.050 846.750 ;
        RECT 736.800 846.000 739.050 847.050 ;
        RECT 740.100 846.000 742.200 847.050 ;
        RECT 736.800 844.950 738.900 846.000 ;
        RECT 739.950 844.950 742.200 846.000 ;
        RECT 772.950 844.950 778.050 847.050 ;
        RECT 781.950 844.950 787.050 847.050 ;
        RECT 718.950 843.450 721.050 844.050 ;
        RECT 733.950 843.450 736.050 844.050 ;
        RECT 718.950 842.400 736.050 843.450 ;
        RECT 718.950 841.950 721.050 842.400 ;
        RECT 733.950 841.950 736.050 842.400 ;
        RECT 739.950 841.950 742.050 844.950 ;
        RECT 727.950 840.450 730.050 841.050 ;
        RECT 751.950 840.450 754.050 844.050 ;
        RECT 791.100 841.950 796.050 844.050 ;
        RECT 727.950 840.000 754.050 840.450 ;
        RECT 754.950 840.450 757.050 841.050 ;
        RECT 760.950 840.450 763.050 841.050 ;
        RECT 727.950 839.400 753.450 840.000 ;
        RECT 754.950 839.400 763.050 840.450 ;
        RECT 727.950 838.950 730.050 839.400 ;
        RECT 754.950 838.950 757.050 839.400 ;
        RECT 760.950 838.950 763.050 839.400 ;
        RECT 689.850 837.600 691.050 837.750 ;
        RECT 673.950 835.500 676.050 837.600 ;
        RECT 676.950 835.500 679.050 837.600 ;
        RECT 679.950 835.500 682.050 837.600 ;
        RECT 683.850 835.500 685.950 837.600 ;
        RECT 688.950 835.500 691.050 837.600 ;
        RECT 697.950 835.950 700.050 838.050 ;
        RECT 700.950 835.950 703.050 838.050 ;
        RECT 703.950 835.950 706.050 838.050 ;
        RECT 797.850 837.600 799.050 849.600 ;
        RECT 805.800 843.000 807.900 844.050 ;
        RECT 805.800 841.950 808.050 843.000 ;
        RECT 809.100 841.950 814.050 844.050 ;
        RECT 805.950 841.050 808.050 841.950 ;
        RECT 805.800 840.000 808.050 841.050 ;
        RECT 805.800 838.950 807.900 840.000 ;
        RECT 818.100 837.600 819.300 854.400 ;
        RECT 835.950 841.950 841.050 844.050 ;
        RECT 796.950 835.500 799.050 837.600 ;
        RECT 817.950 835.500 820.050 837.600 ;
        RECT 4.950 834.450 7.050 835.050 ;
        RECT 28.950 834.450 31.050 835.050 ;
        RECT 49.950 834.450 52.050 835.050 ;
        RECT 82.950 834.450 85.050 835.050 ;
        RECT 4.950 833.400 18.450 834.450 ;
        RECT 4.950 832.950 7.050 833.400 ;
        RECT 17.400 831.450 18.450 833.400 ;
        RECT 28.950 833.400 85.050 834.450 ;
        RECT 28.950 832.950 31.050 833.400 ;
        RECT 49.950 832.950 52.050 833.400 ;
        RECT 82.950 832.950 85.050 833.400 ;
        RECT 94.950 834.450 97.050 835.050 ;
        RECT 124.950 834.450 127.050 835.050 ;
        RECT 94.950 833.400 127.050 834.450 ;
        RECT 94.950 832.950 97.050 833.400 ;
        RECT 124.950 832.950 127.050 833.400 ;
        RECT 142.950 834.450 145.050 835.050 ;
        RECT 160.950 834.450 163.050 835.050 ;
        RECT 142.950 833.400 163.050 834.450 ;
        RECT 142.950 832.950 145.050 833.400 ;
        RECT 160.950 832.950 163.050 833.400 ;
        RECT 181.950 834.450 184.050 835.050 ;
        RECT 241.950 834.450 247.050 835.050 ;
        RECT 181.950 833.400 247.050 834.450 ;
        RECT 181.950 832.950 184.050 833.400 ;
        RECT 241.950 832.950 247.050 833.400 ;
        RECT 337.950 834.450 340.050 835.050 ;
        RECT 406.950 834.450 409.050 835.050 ;
        RECT 337.950 833.400 409.050 834.450 ;
        RECT 337.950 832.950 340.050 833.400 ;
        RECT 406.950 832.950 409.050 833.400 ;
        RECT 484.950 834.450 487.050 835.050 ;
        RECT 526.950 834.450 529.050 835.050 ;
        RECT 577.950 834.450 580.050 835.050 ;
        RECT 484.950 833.400 580.050 834.450 ;
        RECT 484.950 832.950 487.050 833.400 ;
        RECT 526.950 832.950 529.050 833.400 ;
        RECT 577.950 832.950 580.050 833.400 ;
        RECT 616.950 834.450 619.050 835.050 ;
        RECT 655.950 834.450 658.050 835.050 ;
        RECT 664.950 834.450 667.050 835.050 ;
        RECT 616.950 833.400 667.050 834.450 ;
        RECT 616.950 832.950 619.050 833.400 ;
        RECT 655.950 832.950 658.050 833.400 ;
        RECT 664.950 832.950 667.050 833.400 ;
        RECT 34.950 831.450 37.050 832.050 ;
        RECT 17.400 830.400 37.050 831.450 ;
        RECT 34.950 829.950 37.050 830.400 ;
        RECT 103.950 831.450 106.050 832.050 ;
        RECT 178.950 831.450 181.050 832.050 ;
        RECT 103.950 830.400 181.050 831.450 ;
        RECT 103.950 829.950 106.050 830.400 ;
        RECT 178.950 829.950 181.050 830.400 ;
        RECT 220.950 831.450 223.050 832.050 ;
        RECT 274.950 831.450 277.050 832.050 ;
        RECT 310.950 831.450 313.050 832.050 ;
        RECT 220.950 830.400 313.050 831.450 ;
        RECT 220.950 829.950 223.050 830.400 ;
        RECT 274.950 829.950 277.050 830.400 ;
        RECT 310.950 829.950 313.050 830.400 ;
        RECT 757.950 831.450 760.050 832.050 ;
        RECT 802.950 831.450 805.050 832.050 ;
        RECT 850.950 831.450 853.050 832.050 ;
        RECT 757.950 830.400 853.050 831.450 ;
        RECT 757.950 829.950 760.050 830.400 ;
        RECT 802.950 829.950 805.050 830.400 ;
        RECT 850.950 829.950 853.050 830.400 ;
        RECT 76.950 828.450 79.050 829.050 ;
        RECT 109.950 828.450 112.050 829.050 ;
        RECT 226.950 828.450 229.050 829.050 ;
        RECT 76.950 827.400 229.050 828.450 ;
        RECT 76.950 826.950 79.050 827.400 ;
        RECT 109.950 826.950 112.050 827.400 ;
        RECT 226.950 826.950 229.050 827.400 ;
        RECT 295.950 828.450 298.050 829.050 ;
        RECT 508.800 828.450 510.900 829.050 ;
        RECT 295.950 827.400 510.900 828.450 ;
        RECT 295.950 826.950 298.050 827.400 ;
        RECT 508.800 826.950 510.900 827.400 ;
        RECT 512.100 828.450 514.200 829.050 ;
        RECT 565.950 828.450 568.050 829.050 ;
        RECT 512.100 827.400 568.050 828.450 ;
        RECT 512.100 826.950 514.200 827.400 ;
        RECT 565.950 826.950 568.050 827.400 ;
        RECT 571.950 828.450 574.050 829.050 ;
        RECT 616.950 828.450 619.050 829.050 ;
        RECT 571.950 827.400 619.050 828.450 ;
        RECT 571.950 826.950 574.050 827.400 ;
        RECT 616.950 826.950 619.050 827.400 ;
        RECT 631.950 828.450 634.050 829.050 ;
        RECT 715.950 828.450 718.050 829.050 ;
        RECT 631.950 827.400 718.050 828.450 ;
        RECT 631.950 826.950 634.050 827.400 ;
        RECT 715.950 826.950 718.050 827.400 ;
        RECT 766.950 828.450 769.050 829.050 ;
        RECT 805.950 828.450 808.050 829.050 ;
        RECT 766.950 827.400 808.050 828.450 ;
        RECT 766.950 826.950 769.050 827.400 ;
        RECT 805.950 826.950 808.050 827.400 ;
        RECT 40.950 825.450 43.050 826.050 ;
        RECT 70.950 825.450 73.050 826.050 ;
        RECT 88.950 825.450 91.050 826.050 ;
        RECT 40.950 824.400 91.050 825.450 ;
        RECT 40.950 823.950 43.050 824.400 ;
        RECT 70.950 823.950 73.050 824.400 ;
        RECT 88.950 823.950 91.050 824.400 ;
        RECT 136.950 825.450 139.050 826.050 ;
        RECT 193.950 825.450 196.050 826.050 ;
        RECT 136.950 824.400 196.050 825.450 ;
        RECT 136.950 823.950 139.050 824.400 ;
        RECT 193.950 823.950 196.050 824.400 ;
        RECT 673.950 825.450 676.050 826.050 ;
        RECT 709.950 825.450 712.050 826.050 ;
        RECT 673.950 824.400 712.050 825.450 ;
        RECT 716.400 825.450 717.450 826.950 ;
        RECT 760.950 825.450 763.050 826.050 ;
        RECT 784.950 825.450 787.050 826.050 ;
        RECT 716.400 824.400 787.050 825.450 ;
        RECT 673.950 823.950 676.050 824.400 ;
        RECT 709.950 823.950 712.050 824.400 ;
        RECT 760.950 823.950 763.050 824.400 ;
        RECT 784.950 823.950 787.050 824.400 ;
        RECT 793.950 825.450 796.050 826.050 ;
        RECT 835.950 825.450 838.050 826.050 ;
        RECT 793.950 824.400 838.050 825.450 ;
        RECT 793.950 823.950 796.050 824.400 ;
        RECT 835.950 823.950 838.050 824.400 ;
        RECT 7.950 822.450 10.050 823.050 ;
        RECT 67.950 822.450 70.050 823.050 ;
        RECT 7.950 821.400 70.050 822.450 ;
        RECT 7.950 820.950 10.050 821.400 ;
        RECT 67.950 820.950 70.050 821.400 ;
        RECT 100.950 822.450 103.050 823.050 ;
        RECT 124.950 822.450 127.050 823.050 ;
        RECT 100.950 821.400 127.050 822.450 ;
        RECT 100.950 820.950 103.050 821.400 ;
        RECT 124.950 820.950 127.050 821.400 ;
        RECT 169.950 822.450 172.050 823.050 ;
        RECT 181.950 822.450 184.050 823.050 ;
        RECT 169.950 821.400 184.050 822.450 ;
        RECT 169.950 820.950 172.050 821.400 ;
        RECT 181.950 820.950 184.050 821.400 ;
        RECT 235.950 822.450 238.050 823.050 ;
        RECT 277.950 822.450 280.050 823.050 ;
        RECT 235.950 821.400 280.050 822.450 ;
        RECT 235.950 820.950 238.050 821.400 ;
        RECT 277.950 820.950 280.050 821.400 ;
        RECT 502.950 822.450 505.050 823.050 ;
        RECT 514.950 822.450 517.050 823.050 ;
        RECT 502.950 821.400 517.050 822.450 ;
        RECT 502.950 820.950 505.050 821.400 ;
        RECT 514.950 820.950 517.050 821.400 ;
        RECT 97.950 819.450 100.050 820.050 ;
        RECT 103.950 819.450 106.050 820.050 ;
        RECT 112.950 819.450 115.050 820.050 ;
        RECT 62.400 819.000 90.450 819.450 ;
        RECT 61.950 818.400 90.450 819.000 ;
        RECT 4.950 814.950 10.050 817.050 ;
        RECT 13.950 814.950 19.050 817.050 ;
        RECT 46.950 816.450 49.050 817.050 ;
        RECT 55.950 816.450 58.050 817.050 ;
        RECT 46.950 815.400 58.050 816.450 ;
        RECT 46.950 814.950 49.050 815.400 ;
        RECT 55.950 814.950 58.050 815.400 ;
        RECT 61.950 814.950 64.050 818.400 ;
        RECT 89.400 817.050 90.450 818.400 ;
        RECT 97.950 818.400 115.050 819.450 ;
        RECT 97.950 817.950 100.050 818.400 ;
        RECT 103.950 817.950 106.050 818.400 ;
        RECT 112.950 817.950 115.050 818.400 ;
        RECT 160.950 819.450 163.050 820.050 ;
        RECT 175.950 819.450 178.050 820.050 ;
        RECT 160.950 818.400 178.050 819.450 ;
        RECT 160.950 817.950 163.050 818.400 ;
        RECT 175.950 817.950 178.050 818.400 ;
        RECT 76.950 814.950 81.900 817.050 ;
        RECT 83.100 816.450 85.200 817.050 ;
        RECT 88.950 816.450 91.050 817.050 ;
        RECT 83.100 815.400 91.050 816.450 ;
        RECT 83.100 814.950 85.200 815.400 ;
        RECT 88.950 814.950 91.050 815.400 ;
        RECT 133.950 814.950 139.050 817.050 ;
        RECT 13.950 811.050 16.050 814.050 ;
        RECT 19.950 811.950 25.050 814.050 ;
        RECT 31.950 811.950 37.050 814.050 ;
        RECT 40.950 811.950 46.050 814.050 ;
        RECT 13.950 810.000 19.050 811.050 ;
        RECT 14.400 809.400 19.050 810.000 ;
        RECT 15.000 808.950 19.050 809.400 ;
        RECT 37.950 810.450 40.050 811.050 ;
        RECT 46.950 810.450 49.050 811.050 ;
        RECT 37.950 809.400 49.050 810.450 ;
        RECT 37.950 808.950 40.050 809.400 ;
        RECT 46.950 808.950 49.050 809.400 ;
        RECT 52.950 808.950 55.050 814.050 ;
        RECT 58.950 810.450 61.050 814.050 ;
        RECT 67.950 813.450 70.050 814.050 ;
        RECT 73.950 813.450 76.050 814.050 ;
        RECT 67.950 812.400 76.050 813.450 ;
        RECT 67.950 811.950 70.050 812.400 ;
        RECT 73.950 811.950 76.050 812.400 ;
        RECT 79.950 810.450 82.050 814.050 ;
        RECT 100.800 813.450 102.900 814.050 ;
        RECT 86.400 812.400 102.900 813.450 ;
        RECT 86.400 810.450 87.450 812.400 ;
        RECT 100.800 811.950 102.900 812.400 ;
        RECT 104.100 811.950 109.050 814.050 ;
        RECT 112.950 811.950 118.050 814.050 ;
        RECT 124.950 813.450 127.050 814.050 ;
        RECT 130.950 813.450 136.050 814.050 ;
        RECT 124.950 812.400 136.050 813.450 ;
        RECT 124.950 811.950 127.050 812.400 ;
        RECT 130.950 811.950 136.050 812.400 ;
        RECT 139.950 813.450 142.050 814.050 ;
        RECT 148.950 813.450 151.050 814.050 ;
        RECT 139.950 812.400 151.050 813.450 ;
        RECT 139.950 811.950 142.050 812.400 ;
        RECT 148.950 811.950 151.050 812.400 ;
        RECT 157.950 811.950 160.050 817.050 ;
        RECT 184.950 816.450 187.050 817.050 ;
        RECT 190.950 816.450 193.050 817.050 ;
        RECT 184.950 815.400 193.050 816.450 ;
        RECT 184.950 814.950 187.050 815.400 ;
        RECT 190.950 814.950 193.050 815.400 ;
        RECT 196.950 814.950 199.050 820.050 ;
        RECT 232.950 819.450 235.050 820.050 ;
        RECT 250.950 819.450 253.050 820.050 ;
        RECT 304.950 819.450 307.050 820.050 ;
        RECT 232.950 818.400 307.050 819.450 ;
        RECT 232.950 817.950 235.050 818.400 ;
        RECT 250.950 817.950 253.050 818.400 ;
        RECT 304.950 817.950 307.050 818.400 ;
        RECT 202.950 816.450 205.050 817.050 ;
        RECT 217.950 816.450 220.050 817.050 ;
        RECT 202.950 815.400 220.050 816.450 ;
        RECT 202.950 814.950 205.050 815.400 ;
        RECT 217.950 814.950 220.050 815.400 ;
        RECT 163.950 813.450 166.050 814.050 ;
        RECT 172.950 813.450 175.050 814.050 ;
        RECT 163.950 812.400 175.050 813.450 ;
        RECT 163.950 811.950 166.050 812.400 ;
        RECT 172.950 811.950 175.050 812.400 ;
        RECT 58.950 810.000 87.450 810.450 ;
        RECT 59.400 809.400 87.450 810.000 ;
        RECT 106.950 808.950 112.050 811.050 ;
        RECT 157.950 810.450 160.050 811.050 ;
        RECT 169.950 810.450 172.050 811.050 ;
        RECT 157.950 809.400 172.050 810.450 ;
        RECT 157.950 808.950 160.050 809.400 ;
        RECT 52.950 807.450 55.050 808.050 ;
        RECT 58.950 807.450 61.050 808.050 ;
        RECT 52.950 806.400 61.050 807.450 ;
        RECT 52.950 805.950 55.050 806.400 ;
        RECT 58.950 805.950 61.050 806.400 ;
        RECT 79.950 807.450 82.050 808.050 ;
        RECT 115.950 807.450 118.050 808.050 ;
        RECT 79.950 806.400 118.050 807.450 ;
        RECT 79.950 805.950 82.050 806.400 ;
        RECT 115.950 805.950 118.050 806.400 ;
        RECT 136.950 807.450 139.050 808.050 ;
        RECT 163.950 807.450 166.050 808.050 ;
        RECT 136.950 806.400 166.050 807.450 ;
        RECT 136.950 805.950 139.050 806.400 ;
        RECT 163.950 805.950 166.050 806.400 ;
        RECT 169.950 805.950 172.050 809.400 ;
        RECT 175.950 805.950 178.050 811.050 ;
        RECT 193.950 808.950 196.050 814.050 ;
        RECT 199.950 811.950 205.050 814.050 ;
        RECT 208.950 813.450 211.050 814.050 ;
        RECT 214.950 813.450 217.050 814.050 ;
        RECT 208.950 812.400 217.050 813.450 ;
        RECT 208.950 811.950 211.050 812.400 ;
        RECT 214.950 811.950 217.050 812.400 ;
        RECT 226.950 811.950 232.050 814.050 ;
        RECT 235.950 811.950 241.050 814.050 ;
        RECT 250.950 811.950 253.050 817.050 ;
        RECT 256.950 811.950 259.050 817.050 ;
        RECT 277.950 811.950 280.050 817.050 ;
        RECT 311.100 816.000 313.200 817.050 ;
        RECT 310.950 814.950 313.200 816.000 ;
        RECT 310.950 814.050 313.050 814.950 ;
        RECT 289.950 813.450 292.050 814.050 ;
        RECT 295.950 813.450 298.050 814.050 ;
        RECT 289.950 812.400 298.050 813.450 ;
        RECT 289.950 811.950 292.050 812.400 ;
        RECT 295.950 811.950 298.050 812.400 ;
        RECT 301.950 813.450 304.050 814.050 ;
        RECT 307.800 813.450 309.900 814.050 ;
        RECT 301.950 812.400 309.900 813.450 ;
        RECT 310.950 813.000 313.200 814.050 ;
        RECT 301.950 811.950 304.050 812.400 ;
        RECT 307.800 811.950 309.900 812.400 ;
        RECT 311.100 811.950 313.200 813.000 ;
        RECT 316.950 811.950 319.050 817.050 ;
        RECT 355.950 816.450 358.050 820.050 ;
        RECT 376.950 819.450 379.050 820.050 ;
        RECT 385.950 819.450 388.050 820.050 ;
        RECT 376.950 818.400 388.050 819.450 ;
        RECT 376.950 817.950 379.050 818.400 ;
        RECT 385.950 817.950 388.050 818.400 ;
        RECT 403.950 819.450 406.050 820.050 ;
        RECT 424.950 819.450 427.050 820.050 ;
        RECT 403.950 818.400 427.050 819.450 ;
        RECT 403.950 817.950 406.050 818.400 ;
        RECT 424.950 817.950 427.050 818.400 ;
        RECT 445.950 819.450 448.050 820.050 ;
        RECT 457.950 819.450 460.050 820.050 ;
        RECT 445.950 818.400 460.050 819.450 ;
        RECT 445.950 817.950 448.050 818.400 ;
        RECT 457.950 817.950 460.050 818.400 ;
        RECT 472.950 819.450 475.050 820.050 ;
        RECT 484.950 819.450 487.050 820.050 ;
        RECT 472.950 818.400 487.050 819.450 ;
        RECT 472.950 817.950 475.050 818.400 ;
        RECT 484.950 817.950 487.050 818.400 ;
        RECT 505.950 817.050 508.050 820.050 ;
        RECT 335.400 816.000 372.450 816.450 ;
        RECT 334.950 815.400 373.050 816.000 ;
        RECT 334.950 811.950 337.050 815.400 ;
        RECT 355.950 811.950 360.900 814.050 ;
        RECT 362.100 811.950 367.050 814.050 ;
        RECT 370.950 811.950 373.050 815.400 ;
        RECT 469.950 814.950 472.050 817.050 ;
        RECT 475.950 816.450 478.050 817.050 ;
        RECT 502.800 816.450 504.900 817.050 ;
        RECT 475.950 816.000 504.900 816.450 ;
        RECT 505.950 816.000 508.200 817.050 ;
        RECT 475.950 815.400 505.050 816.000 ;
        RECT 475.950 814.950 478.050 815.400 ;
        RECT 502.800 814.950 505.050 815.400 ;
        RECT 506.100 814.950 508.200 816.000 ;
        RECT 511.950 814.950 514.050 820.050 ;
        RECT 580.950 819.450 583.050 820.050 ;
        RECT 604.950 819.450 607.050 820.050 ;
        RECT 634.950 819.450 637.050 820.050 ;
        RECT 580.950 818.400 637.050 819.450 ;
        RECT 580.950 817.950 583.050 818.400 ;
        RECT 604.950 817.950 607.050 818.400 ;
        RECT 634.950 817.950 637.050 818.400 ;
        RECT 682.950 819.450 685.050 820.050 ;
        RECT 694.950 819.450 697.050 820.050 ;
        RECT 751.950 819.450 754.050 820.050 ;
        RECT 757.950 819.450 760.050 820.050 ;
        RECT 682.950 819.000 693.450 819.450 ;
        RECT 694.950 819.000 714.600 819.450 ;
        RECT 682.950 818.400 694.050 819.000 ;
        RECT 682.950 817.950 685.050 818.400 ;
        RECT 535.950 816.450 538.050 817.050 ;
        RECT 544.950 816.450 547.050 817.050 ;
        RECT 535.950 815.400 547.050 816.450 ;
        RECT 535.950 814.950 538.050 815.400 ;
        RECT 544.950 814.950 547.050 815.400 ;
        RECT 550.950 816.450 553.050 817.050 ;
        RECT 568.800 816.450 570.900 817.050 ;
        RECT 550.950 815.400 570.900 816.450 ;
        RECT 550.950 814.950 553.050 815.400 ;
        RECT 568.800 814.950 570.900 815.400 ;
        RECT 572.100 816.450 574.200 817.050 ;
        RECT 586.950 816.450 589.050 817.050 ;
        RECT 595.950 816.450 598.050 817.050 ;
        RECT 572.100 815.400 598.050 816.450 ;
        RECT 635.100 816.000 637.200 817.050 ;
        RECT 572.100 814.950 574.200 815.400 ;
        RECT 586.950 814.950 589.050 815.400 ;
        RECT 595.950 814.950 598.050 815.400 ;
        RECT 634.950 814.950 637.200 816.000 ;
        RECT 671.100 816.450 673.200 817.050 ;
        RECT 685.950 816.450 688.050 817.050 ;
        RECT 671.100 815.400 688.050 816.450 ;
        RECT 671.100 814.950 673.200 815.400 ;
        RECT 685.950 814.950 688.050 815.400 ;
        RECT 691.950 814.950 694.050 818.400 ;
        RECT 694.950 818.400 715.050 819.000 ;
        RECT 694.950 817.950 697.050 818.400 ;
        RECT 712.950 817.050 715.050 818.400 ;
        RECT 751.950 818.400 760.050 819.450 ;
        RECT 751.950 817.950 754.050 818.400 ;
        RECT 757.950 817.950 760.050 818.400 ;
        RECT 769.950 817.950 772.050 823.050 ;
        RECT 787.950 822.450 790.050 823.050 ;
        RECT 811.950 822.450 814.050 823.050 ;
        RECT 787.950 821.400 814.050 822.450 ;
        RECT 787.950 820.950 790.050 821.400 ;
        RECT 811.950 820.950 814.050 821.400 ;
        RECT 781.950 817.950 786.900 820.050 ;
        RECT 788.100 819.000 790.200 820.050 ;
        RECT 787.950 817.950 790.200 819.000 ;
        RECT 706.950 814.950 711.900 817.050 ;
        RECT 712.950 816.000 715.200 817.050 ;
        RECT 727.950 816.450 730.050 817.050 ;
        RECT 716.400 816.000 730.050 816.450 ;
        RECT 713.100 814.950 715.200 816.000 ;
        RECT 715.950 815.400 730.050 816.000 ;
        RECT 391.950 813.450 394.050 814.050 ;
        RECT 406.950 813.450 409.050 814.050 ;
        RECT 391.950 812.400 409.050 813.450 ;
        RECT 391.950 811.950 394.050 812.400 ;
        RECT 406.950 811.950 409.050 812.400 ;
        RECT 412.950 811.950 418.050 814.050 ;
        RECT 424.950 811.950 430.050 814.050 ;
        RECT 203.400 810.450 204.450 811.950 ;
        RECT 433.950 811.050 436.050 814.050 ;
        RECT 448.950 813.450 451.050 814.050 ;
        RECT 466.950 813.450 469.050 814.050 ;
        RECT 448.950 812.400 469.050 813.450 ;
        RECT 448.950 811.950 451.050 812.400 ;
        RECT 466.950 811.950 469.050 812.400 ;
        RECT 211.950 810.450 214.050 811.050 ;
        RECT 203.400 809.400 214.050 810.450 ;
        RECT 211.950 808.950 214.050 809.400 ;
        RECT 217.950 810.450 220.050 811.050 ;
        RECT 223.950 810.450 226.050 811.050 ;
        RECT 217.950 809.400 226.050 810.450 ;
        RECT 217.950 808.950 220.050 809.400 ;
        RECT 223.950 808.950 226.050 809.400 ;
        RECT 184.950 807.450 187.050 808.050 ;
        RECT 232.950 807.450 235.050 811.050 ;
        RECT 241.950 810.450 244.050 811.050 ;
        RECT 253.950 810.450 256.050 811.050 ;
        RECT 241.950 809.400 256.050 810.450 ;
        RECT 241.950 808.950 244.050 809.400 ;
        RECT 253.950 808.950 256.050 809.400 ;
        RECT 184.950 807.000 235.050 807.450 ;
        RECT 184.950 806.400 234.450 807.000 ;
        RECT 184.950 805.950 187.050 806.400 ;
        RECT 274.950 805.950 277.050 811.050 ;
        RECT 280.950 810.450 283.050 811.050 ;
        RECT 289.950 810.450 292.050 811.050 ;
        RECT 280.950 809.400 292.050 810.450 ;
        RECT 280.950 808.950 283.050 809.400 ;
        RECT 289.950 808.950 292.050 809.400 ;
        RECT 295.950 808.950 301.050 811.050 ;
        RECT 313.950 810.450 316.050 811.050 ;
        RECT 302.400 809.400 316.050 810.450 ;
        RECT 280.950 807.450 283.050 808.050 ;
        RECT 302.400 807.450 303.450 809.400 ;
        RECT 313.950 808.950 316.050 809.400 ;
        RECT 322.950 808.950 327.900 811.050 ;
        RECT 329.100 808.950 334.050 811.050 ;
        RECT 337.950 807.450 340.050 811.050 ;
        RECT 367.950 810.450 370.050 811.050 ;
        RECT 400.950 810.450 403.050 811.050 ;
        RECT 367.950 809.400 403.050 810.450 ;
        RECT 367.950 808.950 370.050 809.400 ;
        RECT 400.950 808.950 403.050 809.400 ;
        RECT 406.950 808.950 412.050 811.050 ;
        RECT 418.950 808.950 424.050 811.050 ;
        RECT 430.800 810.000 432.900 811.050 ;
        RECT 433.950 810.000 436.200 811.050 ;
        RECT 430.800 808.950 433.050 810.000 ;
        RECT 434.100 808.950 436.200 810.000 ;
        RECT 280.950 807.000 340.050 807.450 ;
        RECT 430.950 807.450 433.050 808.950 ;
        RECT 445.950 807.450 448.050 811.050 ;
        RECT 430.950 807.000 448.050 807.450 ;
        RECT 451.950 807.450 454.050 811.050 ;
        RECT 470.400 810.450 471.450 814.950 ;
        RECT 475.950 813.450 478.050 814.050 ;
        RECT 484.950 813.450 487.050 814.050 ;
        RECT 475.950 812.400 487.050 813.450 ;
        RECT 475.950 811.950 478.050 812.400 ;
        RECT 484.950 811.950 487.050 812.400 ;
        RECT 502.950 811.950 505.050 814.950 ;
        RECT 634.950 814.050 637.050 814.950 ;
        RECT 508.950 813.450 511.050 814.050 ;
        RECT 526.950 813.450 529.050 814.050 ;
        RECT 506.400 812.400 529.050 813.450 ;
        RECT 478.950 810.450 483.900 811.050 ;
        RECT 470.400 809.400 483.900 810.450 ;
        RECT 478.950 808.950 483.900 809.400 ;
        RECT 485.100 810.450 490.050 811.050 ;
        RECT 506.400 810.450 507.450 812.400 ;
        RECT 508.950 811.950 511.050 812.400 ;
        RECT 526.950 811.950 529.050 812.400 ;
        RECT 532.950 813.450 535.050 814.050 ;
        RECT 541.800 813.450 543.900 814.050 ;
        RECT 532.950 812.400 543.900 813.450 ;
        RECT 532.950 811.950 535.050 812.400 ;
        RECT 541.800 811.950 543.900 812.400 ;
        RECT 545.100 811.950 550.050 814.050 ;
        RECT 565.800 813.000 567.900 814.050 ;
        RECT 565.800 811.950 568.050 813.000 ;
        RECT 565.950 811.050 568.050 811.950 ;
        RECT 571.950 811.050 574.050 811.200 ;
        RECT 485.100 809.400 507.450 810.450 ;
        RECT 514.950 810.450 517.050 811.050 ;
        RECT 523.950 810.450 526.050 811.050 ;
        RECT 514.950 809.400 526.050 810.450 ;
        RECT 485.100 808.950 490.050 809.400 ;
        RECT 514.950 808.950 517.050 809.400 ;
        RECT 523.950 808.950 526.050 809.400 ;
        RECT 529.950 810.450 532.050 811.050 ;
        RECT 535.950 810.450 538.050 811.050 ;
        RECT 529.950 809.400 538.050 810.450 ;
        RECT 529.950 808.950 532.050 809.400 ;
        RECT 535.950 808.950 538.050 809.400 ;
        RECT 562.800 810.000 564.900 811.050 ;
        RECT 565.800 810.000 568.050 811.050 ;
        RECT 562.800 808.950 565.050 810.000 ;
        RECT 565.800 808.950 567.900 810.000 ;
        RECT 569.100 809.100 574.050 811.050 ;
        RECT 569.100 808.950 573.000 809.100 ;
        RECT 583.950 808.950 586.050 814.050 ;
        RECT 589.950 808.950 592.050 814.050 ;
        RECT 595.950 813.450 598.050 814.050 ;
        RECT 601.950 813.450 604.050 814.050 ;
        RECT 595.950 812.400 604.050 813.450 ;
        RECT 595.950 811.950 598.050 812.400 ;
        RECT 601.950 811.950 604.050 812.400 ;
        RECT 619.950 813.450 622.050 814.050 ;
        RECT 628.950 813.450 633.900 814.050 ;
        RECT 619.950 812.400 633.900 813.450 ;
        RECT 634.950 813.000 637.200 814.050 ;
        RECT 619.950 811.950 622.050 812.400 ;
        RECT 628.950 811.950 633.900 812.400 ;
        RECT 635.100 811.950 637.200 813.000 ;
        RECT 562.950 808.050 565.050 808.950 ;
        RECT 457.950 807.450 460.050 808.050 ;
        RECT 475.950 807.450 478.050 808.050 ;
        RECT 451.950 807.000 478.050 807.450 ;
        RECT 280.950 806.400 339.450 807.000 ;
        RECT 431.250 806.400 448.050 807.000 ;
        RECT 452.400 806.400 478.050 807.000 ;
        RECT 280.950 805.950 283.050 806.400 ;
        RECT 445.950 805.950 448.050 806.400 ;
        RECT 457.950 805.950 460.050 806.400 ;
        RECT 475.950 805.950 478.050 806.400 ;
        RECT 562.800 807.000 565.050 808.050 ;
        RECT 571.950 807.450 574.050 807.900 ;
        RECT 583.950 807.450 586.050 808.050 ;
        RECT 562.800 805.950 564.900 807.000 ;
        RECT 571.950 806.400 586.050 807.450 ;
        RECT 571.950 805.800 574.050 806.400 ;
        RECT 583.950 805.950 586.050 806.400 ;
        RECT 595.950 807.450 598.050 808.050 ;
        RECT 604.950 807.450 607.050 808.050 ;
        RECT 595.950 806.400 607.050 807.450 ;
        RECT 631.950 807.450 634.050 811.050 ;
        RECT 673.950 808.950 676.050 814.050 ;
        RECT 688.950 811.950 693.900 814.050 ;
        RECT 695.100 813.450 697.200 814.050 ;
        RECT 700.950 813.450 703.050 814.050 ;
        RECT 695.100 812.400 703.050 813.450 ;
        RECT 695.100 811.950 697.200 812.400 ;
        RECT 700.950 811.950 703.050 812.400 ;
        RECT 709.950 810.450 712.050 814.050 ;
        RECT 715.950 811.950 718.050 815.400 ;
        RECT 727.950 814.950 730.050 815.400 ;
        RECT 730.950 814.050 733.050 814.200 ;
        RECT 730.950 812.100 736.050 814.050 ;
        RECT 732.000 811.950 736.050 812.100 ;
        RECT 739.950 811.950 742.050 817.050 ;
        RECT 754.950 813.450 757.050 817.050 ;
        RECT 772.950 814.950 778.050 817.050 ;
        RECT 787.950 814.950 790.050 817.950 ;
        RECT 802.950 814.950 808.050 817.050 ;
        RECT 811.950 814.950 814.050 820.050 ;
        RECT 817.950 816.450 820.050 817.050 ;
        RECT 823.950 816.450 826.050 817.050 ;
        RECT 817.950 815.400 826.050 816.450 ;
        RECT 817.950 814.950 820.050 815.400 ;
        RECT 823.950 814.950 826.050 815.400 ;
        RECT 773.400 813.450 774.450 814.950 ;
        RECT 832.950 814.050 835.050 817.050 ;
        RECT 838.950 814.950 841.050 820.050 ;
        RECT 844.950 814.050 847.050 817.050 ;
        RECT 754.950 812.400 774.450 813.450 ;
        RECT 787.950 813.450 790.050 814.050 ;
        RECT 793.950 813.450 796.050 814.050 ;
        RECT 787.950 812.400 796.050 813.450 ;
        RECT 754.950 811.950 757.050 812.400 ;
        RECT 787.950 811.950 790.050 812.400 ;
        RECT 793.950 811.950 796.050 812.400 ;
        RECT 808.950 811.050 811.050 814.050 ;
        RECT 814.950 811.950 817.050 814.050 ;
        RECT 832.800 813.000 835.050 814.050 ;
        RECT 836.100 813.000 838.200 814.050 ;
        RECT 832.800 811.950 834.900 813.000 ;
        RECT 835.950 811.950 838.200 813.000 ;
        RECT 841.800 813.000 843.900 814.050 ;
        RECT 844.950 813.000 847.200 814.050 ;
        RECT 841.800 811.950 844.050 813.000 ;
        RECT 845.100 811.950 847.200 813.000 ;
        RECT 730.950 810.450 733.050 810.900 ;
        RECT 709.950 810.000 733.050 810.450 ;
        RECT 808.950 810.000 814.050 811.050 ;
        RECT 710.400 809.400 733.050 810.000 ;
        RECT 809.400 809.400 814.050 810.000 ;
        RECT 730.950 808.800 733.050 809.400 ;
        RECT 810.000 808.950 814.050 809.400 ;
        RECT 815.400 810.450 816.450 811.950 ;
        RECT 835.950 810.450 838.050 811.950 ;
        RECT 815.400 810.000 838.050 810.450 ;
        RECT 841.950 810.450 844.050 811.950 ;
        RECT 850.950 810.450 853.050 811.050 ;
        RECT 841.950 810.000 853.050 810.450 ;
        RECT 815.400 809.400 837.600 810.000 ;
        RECT 842.250 809.400 853.050 810.000 ;
        RECT 646.950 807.450 649.050 808.050 ;
        RECT 697.950 807.450 700.050 808.050 ;
        RECT 631.950 807.000 700.050 807.450 ;
        RECT 632.400 806.400 700.050 807.000 ;
        RECT 595.950 805.950 598.050 806.400 ;
        RECT 604.950 805.950 607.050 806.400 ;
        RECT 646.950 805.950 649.050 806.400 ;
        RECT 697.950 805.950 700.050 806.400 ;
        RECT 709.950 807.450 712.050 808.050 ;
        RECT 754.950 807.450 757.050 808.050 ;
        RECT 709.950 806.400 757.050 807.450 ;
        RECT 709.950 805.950 712.050 806.400 ;
        RECT 754.950 805.950 757.050 806.400 ;
        RECT 769.950 807.450 772.050 808.050 ;
        RECT 815.400 807.450 816.450 809.400 ;
        RECT 850.950 808.950 853.050 809.400 ;
        RECT 769.950 806.400 816.450 807.450 ;
        RECT 769.950 805.950 772.050 806.400 ;
        RECT 25.950 804.450 28.050 805.050 ;
        RECT 61.950 804.450 64.050 805.050 ;
        RECT 25.950 803.400 64.050 804.450 ;
        RECT 25.950 802.950 28.050 803.400 ;
        RECT 61.950 802.950 64.050 803.400 ;
        RECT 175.950 804.450 178.050 805.050 ;
        RECT 232.950 804.450 235.050 805.050 ;
        RECT 175.950 803.400 235.050 804.450 ;
        RECT 175.950 802.950 178.050 803.400 ;
        RECT 232.950 802.950 235.050 803.400 ;
        RECT 265.950 804.450 268.050 805.050 ;
        RECT 298.950 804.450 301.050 805.050 ;
        RECT 331.950 804.450 334.050 805.050 ;
        RECT 265.950 803.400 334.050 804.450 ;
        RECT 265.950 802.950 268.050 803.400 ;
        RECT 298.950 802.950 301.050 803.400 ;
        RECT 331.950 802.950 334.050 803.400 ;
        RECT 379.950 804.450 382.050 805.050 ;
        RECT 460.950 804.450 463.050 805.050 ;
        RECT 379.950 803.400 463.050 804.450 ;
        RECT 379.950 802.950 382.050 803.400 ;
        RECT 460.950 802.950 463.050 803.400 ;
        RECT 526.950 804.450 529.050 805.050 ;
        RECT 547.950 804.450 550.050 805.050 ;
        RECT 526.950 803.400 550.050 804.450 ;
        RECT 526.950 802.950 529.050 803.400 ;
        RECT 547.950 802.950 550.050 803.400 ;
        RECT 595.950 804.450 598.050 805.050 ;
        RECT 700.950 804.450 706.050 805.050 ;
        RECT 595.950 803.400 706.050 804.450 ;
        RECT 595.950 802.950 598.050 803.400 ;
        RECT 700.950 802.950 706.050 803.400 ;
        RECT 727.950 804.450 730.050 805.050 ;
        RECT 781.950 804.450 784.050 805.050 ;
        RECT 727.950 803.400 784.050 804.450 ;
        RECT 727.950 802.950 730.050 803.400 ;
        RECT 781.950 802.950 784.050 803.400 ;
        RECT 121.950 801.450 124.050 802.050 ;
        RECT 166.950 801.450 169.050 802.050 ;
        RECT 184.950 801.450 187.050 802.050 ;
        RECT 208.950 801.450 211.050 802.050 ;
        RECT 121.950 800.400 187.050 801.450 ;
        RECT 121.950 799.950 124.050 800.400 ;
        RECT 166.950 799.950 169.050 800.400 ;
        RECT 184.950 799.950 187.050 800.400 ;
        RECT 188.400 800.400 211.050 801.450 ;
        RECT 130.950 798.450 133.050 799.050 ;
        RECT 148.950 798.450 151.050 799.050 ;
        RECT 188.400 798.450 189.450 800.400 ;
        RECT 208.950 799.950 211.050 800.400 ;
        RECT 214.950 801.450 217.050 802.050 ;
        RECT 307.950 801.450 310.050 802.050 ;
        RECT 214.950 800.400 310.050 801.450 ;
        RECT 214.950 799.950 217.050 800.400 ;
        RECT 307.950 799.950 310.050 800.400 ;
        RECT 469.950 801.450 472.050 802.050 ;
        RECT 532.950 801.450 535.050 802.050 ;
        RECT 469.950 800.400 535.050 801.450 ;
        RECT 469.950 799.950 472.050 800.400 ;
        RECT 532.950 799.950 535.050 800.400 ;
        RECT 643.950 801.450 646.050 802.050 ;
        RECT 733.950 801.450 736.050 802.050 ;
        RECT 643.950 800.400 736.050 801.450 ;
        RECT 643.950 799.950 646.050 800.400 ;
        RECT 733.950 799.950 736.050 800.400 ;
        RECT 739.950 801.450 742.050 802.050 ;
        RECT 838.950 801.450 841.050 802.050 ;
        RECT 739.950 800.400 841.050 801.450 ;
        RECT 739.950 799.950 742.050 800.400 ;
        RECT 838.950 799.950 841.050 800.400 ;
        RECT 130.950 797.400 189.450 798.450 ;
        RECT 193.950 798.450 196.050 799.050 ;
        RECT 205.950 798.450 208.050 799.050 ;
        RECT 193.950 797.400 208.050 798.450 ;
        RECT 130.950 796.950 133.050 797.400 ;
        RECT 148.950 796.950 151.050 797.400 ;
        RECT 193.950 796.950 196.050 797.400 ;
        RECT 205.950 796.950 208.050 797.400 ;
        RECT 244.950 798.450 247.050 799.050 ;
        RECT 292.950 798.450 295.050 799.050 ;
        RECT 244.950 797.400 295.050 798.450 ;
        RECT 244.950 796.950 247.050 797.400 ;
        RECT 292.950 796.950 295.050 797.400 ;
        RECT 433.950 798.450 436.050 799.050 ;
        RECT 457.950 798.450 460.050 799.050 ;
        RECT 433.950 797.400 460.050 798.450 ;
        RECT 433.950 796.950 436.050 797.400 ;
        RECT 457.950 796.950 460.050 797.400 ;
        RECT 478.950 798.450 481.050 799.050 ;
        RECT 511.950 798.450 514.050 799.050 ;
        RECT 574.800 798.450 576.900 799.050 ;
        RECT 478.950 797.400 576.900 798.450 ;
        RECT 478.950 796.950 481.050 797.400 ;
        RECT 511.950 796.950 514.050 797.400 ;
        RECT 574.800 796.950 576.900 797.400 ;
        RECT 578.100 798.450 580.200 799.050 ;
        RECT 622.950 798.450 625.050 799.050 ;
        RECT 578.100 797.400 625.050 798.450 ;
        RECT 578.100 796.950 580.200 797.400 ;
        RECT 622.950 796.950 625.050 797.400 ;
        RECT 682.950 798.450 685.050 799.050 ;
        RECT 727.950 798.450 730.050 799.050 ;
        RECT 682.950 797.400 730.050 798.450 ;
        RECT 682.950 796.950 685.050 797.400 ;
        RECT 727.950 796.950 730.050 797.400 ;
        RECT 760.950 796.950 766.050 799.050 ;
        RECT 814.950 798.450 817.050 799.050 ;
        RECT 832.950 798.450 835.050 799.050 ;
        RECT 814.950 797.400 835.050 798.450 ;
        RECT 814.950 796.950 817.050 797.400 ;
        RECT 832.950 796.950 835.050 797.400 ;
        RECT 112.950 795.450 115.050 796.050 ;
        RECT 133.950 795.450 136.050 796.050 ;
        RECT 112.950 794.400 136.050 795.450 ;
        RECT 112.950 793.950 115.050 794.400 ;
        RECT 133.950 793.950 136.050 794.400 ;
        RECT 181.950 795.450 184.050 796.050 ;
        RECT 238.950 795.450 241.050 796.050 ;
        RECT 181.950 794.400 241.050 795.450 ;
        RECT 181.950 793.950 184.050 794.400 ;
        RECT 238.950 793.950 241.050 794.400 ;
        RECT 583.950 795.450 586.050 796.050 ;
        RECT 595.950 795.450 598.050 796.050 ;
        RECT 583.950 794.400 598.050 795.450 ;
        RECT 583.950 793.950 586.050 794.400 ;
        RECT 595.950 793.950 598.050 794.400 ;
        RECT 631.950 795.450 634.050 796.050 ;
        RECT 688.800 795.450 690.900 796.050 ;
        RECT 631.950 794.400 690.900 795.450 ;
        RECT 631.950 793.950 634.050 794.400 ;
        RECT 688.800 793.950 690.900 794.400 ;
        RECT 692.100 795.450 694.200 796.050 ;
        RECT 730.950 795.450 733.050 796.050 ;
        RECT 692.100 794.400 733.050 795.450 ;
        RECT 692.100 793.950 694.200 794.400 ;
        RECT 730.950 793.950 733.050 794.400 ;
        RECT 223.950 792.450 226.050 793.050 ;
        RECT 262.950 792.450 265.050 793.050 ;
        RECT 223.950 791.400 265.050 792.450 ;
        RECT 223.950 790.950 226.050 791.400 ;
        RECT 262.950 790.950 265.050 791.400 ;
        RECT 406.950 792.450 409.050 793.050 ;
        RECT 454.950 792.450 457.050 793.050 ;
        RECT 406.950 791.400 457.050 792.450 ;
        RECT 406.950 790.950 409.050 791.400 ;
        RECT 454.950 790.950 457.050 791.400 ;
        RECT 535.950 792.450 538.050 793.050 ;
        RECT 580.950 792.450 583.050 793.050 ;
        RECT 535.950 791.400 583.050 792.450 ;
        RECT 535.950 790.950 538.050 791.400 ;
        RECT 580.950 790.950 583.050 791.400 ;
        RECT 655.950 792.450 658.050 793.050 ;
        RECT 709.950 792.450 712.050 793.050 ;
        RECT 814.950 792.450 817.050 793.050 ;
        RECT 655.950 791.400 817.050 792.450 ;
        RECT 655.950 790.950 658.050 791.400 ;
        RECT 709.950 790.950 712.050 791.400 ;
        RECT 814.950 790.950 817.050 791.400 ;
        RECT 16.950 789.450 19.050 790.050 ;
        RECT 22.950 789.450 25.050 790.050 ;
        RECT 16.950 788.400 25.050 789.450 ;
        RECT 16.950 787.950 19.050 788.400 ;
        RECT 22.950 787.950 25.050 788.400 ;
        RECT 142.950 789.450 145.050 790.050 ;
        RECT 184.950 789.450 187.050 790.050 ;
        RECT 265.950 789.450 268.050 790.050 ;
        RECT 142.950 788.400 268.050 789.450 ;
        RECT 142.950 787.950 145.050 788.400 ;
        RECT 184.950 787.950 187.050 788.400 ;
        RECT 265.950 787.950 268.050 788.400 ;
        RECT 349.950 789.450 352.050 790.050 ;
        RECT 478.950 789.450 481.050 790.050 ;
        RECT 349.950 788.400 481.050 789.450 ;
        RECT 349.950 787.950 352.050 788.400 ;
        RECT 478.950 787.950 481.050 788.400 ;
        RECT 577.950 789.450 580.050 790.050 ;
        RECT 661.950 789.450 664.050 790.050 ;
        RECT 577.950 788.400 664.050 789.450 ;
        RECT 577.950 787.950 580.050 788.400 ;
        RECT 661.950 787.950 664.050 788.400 ;
        RECT 13.950 786.450 16.050 787.050 ;
        RECT 40.950 786.450 43.050 787.050 ;
        RECT 13.950 785.400 43.050 786.450 ;
        RECT 13.950 784.950 16.050 785.400 ;
        RECT 40.950 784.950 43.050 785.400 ;
        RECT 169.950 786.450 172.050 787.050 ;
        RECT 193.950 786.450 196.050 787.050 ;
        RECT 214.950 786.450 217.050 787.050 ;
        RECT 289.950 786.450 292.050 787.050 ;
        RECT 169.950 785.400 292.050 786.450 ;
        RECT 169.950 784.950 172.050 785.400 ;
        RECT 193.950 784.950 196.050 785.400 ;
        RECT 214.950 784.950 217.050 785.400 ;
        RECT 289.950 784.950 292.050 785.400 ;
        RECT 316.950 786.450 319.050 787.050 ;
        RECT 355.950 786.450 358.050 787.050 ;
        RECT 448.950 786.450 451.050 787.050 ;
        RECT 316.950 785.400 342.450 786.450 ;
        RECT 316.950 784.950 319.050 785.400 ;
        RECT 341.400 784.050 342.450 785.400 ;
        RECT 355.950 785.400 451.050 786.450 ;
        RECT 355.950 784.950 358.050 785.400 ;
        RECT 448.950 784.950 451.050 785.400 ;
        RECT 562.950 786.450 565.050 787.050 ;
        RECT 589.950 786.450 592.050 787.200 ;
        RECT 640.800 786.450 642.900 787.050 ;
        RECT 562.950 785.400 642.900 786.450 ;
        RECT 562.950 784.950 565.050 785.400 ;
        RECT 589.950 785.100 592.050 785.400 ;
        RECT 640.800 784.950 642.900 785.400 ;
        RECT 644.100 786.450 646.200 787.050 ;
        RECT 673.950 786.450 676.050 787.050 ;
        RECT 644.100 785.400 676.050 786.450 ;
        RECT 644.100 784.950 646.200 785.400 ;
        RECT 673.950 784.950 676.050 785.400 ;
        RECT 775.950 784.950 778.050 787.050 ;
        RECT 778.950 784.950 781.050 787.050 ;
        RECT 781.950 784.950 784.050 787.050 ;
        RECT 19.950 783.450 22.050 784.050 ;
        RECT 49.950 783.450 52.050 784.050 ;
        RECT 70.950 783.450 73.050 784.050 ;
        RECT 19.950 782.400 73.050 783.450 ;
        RECT 19.950 781.950 22.050 782.400 ;
        RECT 49.950 781.950 52.050 782.400 ;
        RECT 70.950 781.950 73.050 782.400 ;
        RECT 199.950 783.450 202.050 784.050 ;
        RECT 253.950 783.450 256.050 784.050 ;
        RECT 331.950 783.450 334.050 784.050 ;
        RECT 199.950 782.400 334.050 783.450 ;
        RECT 199.950 781.950 202.050 782.400 ;
        RECT 253.950 781.950 256.050 782.400 ;
        RECT 331.950 781.950 334.050 782.400 ;
        RECT 340.950 783.450 343.050 784.050 ;
        RECT 352.950 783.450 355.050 784.050 ;
        RECT 340.950 782.400 355.050 783.450 ;
        RECT 340.950 781.950 343.050 782.400 ;
        RECT 352.950 781.950 355.050 782.400 ;
        RECT 400.950 783.450 403.050 784.050 ;
        RECT 430.950 783.450 433.050 784.050 ;
        RECT 400.950 782.400 433.050 783.450 ;
        RECT 400.950 781.950 403.050 782.400 ;
        RECT 430.950 781.950 433.050 782.400 ;
        RECT 505.950 783.450 508.050 784.050 ;
        RECT 517.950 783.450 520.050 784.050 ;
        RECT 505.950 782.400 520.050 783.450 ;
        RECT 505.950 781.950 508.050 782.400 ;
        RECT 517.950 781.950 520.050 782.400 ;
        RECT 553.950 783.450 556.050 784.050 ;
        RECT 589.950 783.450 592.050 783.900 ;
        RECT 553.950 782.400 592.050 783.450 ;
        RECT 553.950 781.950 556.050 782.400 ;
        RECT 589.950 781.800 592.050 782.400 ;
        RECT 40.950 780.450 43.050 781.050 ;
        RECT 115.950 780.450 118.050 781.050 ;
        RECT 145.950 780.450 148.050 781.050 ;
        RECT 40.950 780.000 69.450 780.450 ;
        RECT 40.950 779.400 70.050 780.000 ;
        RECT 40.950 778.950 43.050 779.400 ;
        RECT 10.950 777.450 13.050 778.050 ;
        RECT 25.950 777.450 31.050 778.050 ;
        RECT 10.950 776.400 31.050 777.450 ;
        RECT 10.950 775.950 13.050 776.400 ;
        RECT 25.950 775.950 31.050 776.400 ;
        RECT 34.950 775.950 40.050 778.050 ;
        RECT 10.950 769.950 13.050 775.050 ;
        RECT 31.950 774.450 34.050 775.050 ;
        RECT 40.950 774.450 43.050 775.050 ;
        RECT 31.950 773.400 43.050 774.450 ;
        RECT 31.950 772.950 34.050 773.400 ;
        RECT 40.950 772.950 43.050 773.400 ;
        RECT 49.950 772.950 52.050 778.050 ;
        RECT 67.950 777.450 70.050 779.400 ;
        RECT 115.950 779.400 148.050 780.450 ;
        RECT 115.950 778.950 118.050 779.400 ;
        RECT 145.950 778.950 148.050 779.400 ;
        RECT 166.950 780.450 169.050 781.050 ;
        RECT 184.950 780.450 187.050 781.050 ;
        RECT 166.950 779.400 187.050 780.450 ;
        RECT 166.950 778.950 169.050 779.400 ;
        RECT 184.950 778.950 187.050 779.400 ;
        RECT 232.950 780.450 235.050 781.050 ;
        RECT 265.950 780.450 268.050 781.050 ;
        RECT 232.950 779.400 268.050 780.450 ;
        RECT 232.950 778.950 235.050 779.400 ;
        RECT 265.950 778.950 268.050 779.400 ;
        RECT 274.950 780.450 279.000 781.050 ;
        RECT 280.950 780.450 283.050 781.050 ;
        RECT 364.950 780.450 367.050 781.050 ;
        RECT 430.950 780.450 433.050 781.050 ;
        RECT 562.950 780.450 565.050 781.050 ;
        RECT 274.950 780.000 279.300 780.450 ;
        RECT 274.950 778.950 280.050 780.000 ;
        RECT 280.950 779.400 363.450 780.450 ;
        RECT 280.950 778.950 283.050 779.400 ;
        RECT 277.950 778.050 280.050 778.950 ;
        RECT 56.400 777.000 70.050 777.450 ;
        RECT 55.950 776.400 70.050 777.000 ;
        RECT 55.950 772.950 58.050 776.400 ;
        RECT 67.950 775.950 70.050 776.400 ;
        RECT 76.950 777.450 79.050 778.050 ;
        RECT 85.950 777.450 88.050 778.050 ;
        RECT 103.950 777.450 106.050 778.050 ;
        RECT 76.950 776.400 88.050 777.450 ;
        RECT 92.400 777.000 106.050 777.450 ;
        RECT 116.100 777.000 118.200 778.050 ;
        RECT 76.950 775.950 79.050 776.400 ;
        RECT 85.950 775.950 88.050 776.400 ;
        RECT 91.950 776.400 106.050 777.000 ;
        RECT 16.950 769.950 22.050 772.050 ;
        RECT 43.950 769.950 49.050 772.050 ;
        RECT 13.950 768.450 16.050 769.050 ;
        RECT 22.950 768.450 25.050 769.050 ;
        RECT 13.950 767.400 25.050 768.450 ;
        RECT 13.950 766.950 16.050 767.400 ;
        RECT 22.950 766.950 25.050 767.400 ;
        RECT 52.950 768.450 55.050 772.050 ;
        RECT 64.950 769.950 67.050 775.050 ;
        RECT 70.950 771.450 73.050 775.050 ;
        RECT 91.950 772.950 94.050 776.400 ;
        RECT 103.950 775.950 106.050 776.400 ;
        RECT 115.950 775.950 118.200 777.000 ;
        RECT 115.950 775.050 118.050 775.950 ;
        RECT 109.950 772.950 114.900 775.050 ;
        RECT 115.950 774.000 118.200 775.050 ;
        RECT 130.800 774.450 132.900 775.050 ;
        RECT 116.100 772.950 118.200 774.000 ;
        RECT 125.400 773.400 132.900 774.450 ;
        RECT 85.950 771.450 88.050 772.050 ;
        RECT 70.950 771.000 88.050 771.450 ;
        RECT 71.400 770.400 88.050 771.000 ;
        RECT 85.950 769.950 88.050 770.400 ;
        RECT 97.950 769.950 102.900 772.050 ;
        RECT 104.100 771.450 106.200 772.050 ;
        RECT 112.950 771.450 115.050 772.050 ;
        RECT 104.100 770.400 115.050 771.450 ;
        RECT 104.100 769.950 106.200 770.400 ;
        RECT 112.950 769.950 115.050 770.400 ;
        RECT 118.950 771.450 121.050 772.050 ;
        RECT 125.400 771.450 126.450 773.400 ;
        RECT 130.800 772.950 132.900 773.400 ;
        RECT 133.800 774.000 135.900 775.050 ;
        RECT 137.100 774.450 139.200 775.050 ;
        RECT 145.950 774.450 148.050 775.050 ;
        RECT 133.800 772.950 136.050 774.000 ;
        RECT 137.100 773.400 148.050 774.450 ;
        RECT 137.100 772.950 139.200 773.400 ;
        RECT 145.950 772.950 148.050 773.400 ;
        RECT 133.950 772.050 136.050 772.950 ;
        RECT 118.950 770.400 126.450 771.450 ;
        RECT 64.950 768.450 67.050 769.050 ;
        RECT 52.950 767.400 67.050 768.450 ;
        RECT 52.950 766.950 55.050 767.400 ;
        RECT 64.950 766.950 67.050 767.400 ;
        RECT 118.950 766.950 121.050 770.400 ;
        RECT 127.950 766.950 130.050 772.050 ;
        RECT 133.800 771.000 136.050 772.050 ;
        RECT 133.800 769.950 135.900 771.000 ;
        RECT 154.950 769.950 157.050 775.050 ;
        RECT 193.950 772.950 196.050 778.050 ;
        RECT 205.950 775.950 211.050 778.050 ;
        RECT 217.950 775.950 223.050 778.050 ;
        RECT 160.950 766.950 163.050 772.050 ;
        RECT 166.950 769.950 172.050 772.050 ;
        RECT 175.800 771.000 177.900 772.050 ;
        RECT 179.100 771.450 181.200 772.050 ;
        RECT 187.950 771.450 190.050 772.050 ;
        RECT 175.800 769.950 178.050 771.000 ;
        RECT 179.100 770.400 190.050 771.450 ;
        RECT 179.100 769.950 181.200 770.400 ;
        RECT 187.950 769.950 190.050 770.400 ;
        RECT 175.950 769.050 178.050 769.950 ;
        RECT 172.800 768.450 174.900 769.050 ;
        RECT 164.400 767.400 174.900 768.450 ;
        RECT 175.950 768.000 178.200 769.050 ;
        RECT 196.950 768.450 199.050 772.050 ;
        RECT 199.950 771.450 202.050 775.050 ;
        RECT 211.950 772.950 217.050 775.050 ;
        RECT 220.950 774.450 223.050 775.050 ;
        RECT 229.950 774.450 232.050 778.050 ;
        RECT 235.950 775.050 238.050 778.050 ;
        RECT 277.800 777.000 280.050 778.050 ;
        RECT 281.100 777.000 283.200 778.050 ;
        RECT 288.000 777.450 292.050 778.050 ;
        RECT 277.800 775.950 279.900 777.000 ;
        RECT 280.950 775.950 283.200 777.000 ;
        RECT 287.400 775.950 292.050 777.450 ;
        RECT 295.950 775.950 298.050 779.400 ;
        RECT 358.950 777.450 361.050 778.050 ;
        RECT 338.400 777.000 361.050 777.450 ;
        RECT 337.950 776.400 361.050 777.000 ;
        RECT 362.400 777.450 363.450 779.400 ;
        RECT 364.950 780.000 426.450 780.450 ;
        RECT 430.950 780.000 465.450 780.450 ;
        RECT 364.950 779.400 427.050 780.000 ;
        RECT 364.950 778.950 367.050 779.400 ;
        RECT 388.950 777.450 391.050 778.050 ;
        RECT 362.400 776.400 391.050 777.450 ;
        RECT 220.950 774.000 232.050 774.450 ;
        RECT 232.800 774.000 234.900 775.050 ;
        RECT 235.950 774.000 238.200 775.050 ;
        RECT 220.950 773.400 231.450 774.000 ;
        RECT 220.950 771.450 223.050 773.400 ;
        RECT 232.800 772.950 235.050 774.000 ;
        RECT 236.100 772.950 238.200 774.000 ;
        RECT 253.950 772.950 259.050 775.050 ;
        RECT 265.950 774.450 268.050 775.050 ;
        RECT 274.950 774.450 277.050 775.050 ;
        RECT 265.950 773.400 277.050 774.450 ;
        RECT 265.950 772.950 268.050 773.400 ;
        RECT 274.950 772.950 277.050 773.400 ;
        RECT 280.950 772.950 283.050 775.950 ;
        RECT 199.950 771.000 223.050 771.450 ;
        RECT 200.400 770.400 223.050 771.000 ;
        RECT 220.950 769.950 223.050 770.400 ;
        RECT 232.950 769.950 235.050 772.950 ;
        RECT 287.400 772.050 288.450 775.950 ;
        RECT 289.950 772.950 295.050 775.050 ;
        RECT 301.950 774.450 304.050 775.050 ;
        RECT 310.950 774.450 313.050 775.050 ;
        RECT 301.950 773.400 313.050 774.450 ;
        RECT 301.950 772.950 304.050 773.400 ;
        RECT 310.950 772.950 313.050 773.400 ;
        RECT 316.950 772.950 322.050 775.050 ;
        RECT 330.000 774.450 334.050 775.050 ;
        RECT 329.400 772.950 334.050 774.450 ;
        RECT 337.950 772.950 340.050 776.400 ;
        RECT 358.950 775.950 361.050 776.400 ;
        RECT 388.950 775.950 391.050 776.400 ;
        RECT 394.950 775.950 400.050 778.050 ;
        RECT 424.950 775.950 427.050 779.400 ;
        RECT 430.950 779.400 466.050 780.000 ;
        RECT 430.950 775.950 433.050 779.400 ;
        RECT 436.950 777.450 439.050 778.050 ;
        RECT 442.800 777.450 444.900 778.050 ;
        RECT 436.950 776.400 444.900 777.450 ;
        RECT 436.950 775.950 439.050 776.400 ;
        RECT 442.800 775.950 444.900 776.400 ;
        RECT 446.100 775.950 451.050 778.050 ;
        RECT 463.950 775.950 466.050 779.400 ;
        RECT 509.400 779.400 565.050 780.450 ;
        RECT 472.950 777.450 475.050 778.050 ;
        RECT 478.950 777.450 481.050 778.050 ;
        RECT 472.950 776.400 481.050 777.450 ;
        RECT 472.950 775.950 475.050 776.400 ;
        RECT 478.950 775.950 481.050 776.400 ;
        RECT 490.950 775.950 496.050 778.050 ;
        RECT 509.400 777.450 510.450 779.400 ;
        RECT 562.950 778.950 565.050 779.400 ;
        RECT 592.950 780.450 595.050 781.050 ;
        RECT 634.800 780.450 636.900 781.050 ;
        RECT 592.950 779.400 636.900 780.450 ;
        RECT 592.950 778.950 595.050 779.400 ;
        RECT 634.800 778.950 636.900 779.400 ;
        RECT 638.100 780.450 640.200 781.050 ;
        RECT 649.950 780.450 652.050 781.050 ;
        RECT 638.100 779.400 652.050 780.450 ;
        RECT 638.100 778.950 640.200 779.400 ;
        RECT 649.950 778.950 652.050 779.400 ;
        RECT 680.400 779.400 723.450 780.450 ;
        RECT 497.400 776.400 510.450 777.450 ;
        RECT 497.400 775.050 498.450 776.400 ;
        RECT 509.400 775.050 510.450 776.400 ;
        RECT 370.950 772.950 376.050 775.050 ;
        RECT 391.950 772.950 397.050 775.050 ;
        RECT 400.950 774.450 403.050 775.050 ;
        RECT 409.950 774.450 412.050 775.050 ;
        RECT 400.950 773.400 412.050 774.450 ;
        RECT 400.950 772.950 403.050 773.400 ;
        RECT 409.950 772.950 412.050 773.400 ;
        RECT 238.950 771.450 241.050 772.050 ;
        RECT 247.950 771.450 250.050 772.050 ;
        RECT 238.950 770.400 250.050 771.450 ;
        RECT 238.950 769.950 241.050 770.400 ;
        RECT 247.950 769.950 250.050 770.400 ;
        RECT 259.950 769.950 265.050 772.050 ;
        RECT 286.950 769.950 289.050 772.050 ;
        RECT 307.950 771.450 310.050 772.050 ;
        RECT 313.950 771.450 316.050 772.050 ;
        RECT 307.950 770.400 316.050 771.450 ;
        RECT 307.950 769.950 310.050 770.400 ;
        RECT 313.950 769.950 316.050 770.400 ;
        RECT 319.950 771.450 322.050 772.050 ;
        RECT 329.400 771.450 330.450 772.950 ;
        RECT 319.950 770.400 330.450 771.450 ;
        RECT 196.950 768.000 219.450 768.450 ;
        RECT 118.950 765.450 121.050 766.050 ;
        RECT 164.400 765.450 165.450 767.400 ;
        RECT 172.800 766.950 174.900 767.400 ;
        RECT 176.100 766.950 178.200 768.000 ;
        RECT 197.400 767.400 219.450 768.000 ;
        RECT 218.400 766.050 219.450 767.400 ;
        RECT 319.950 766.950 322.050 770.400 ;
        RECT 331.950 769.950 337.050 772.050 ;
        RECT 340.950 769.950 346.050 772.050 ;
        RECT 348.000 771.450 351.900 772.050 ;
        RECT 347.400 771.000 351.900 771.450 ;
        RECT 346.950 769.950 351.900 771.000 ;
        RECT 352.800 771.000 354.900 772.050 ;
        RECT 356.100 771.450 358.200 772.050 ;
        RECT 364.950 771.450 370.050 772.050 ;
        RECT 376.950 771.450 379.050 772.050 ;
        RECT 352.800 769.950 355.050 771.000 ;
        RECT 356.100 770.400 370.050 771.450 ;
        RECT 356.100 769.950 358.200 770.400 ;
        RECT 364.950 769.950 370.050 770.400 ;
        RECT 371.400 770.400 379.050 771.450 ;
        RECT 427.950 771.450 430.050 775.050 ;
        RECT 444.000 774.450 448.050 775.050 ;
        RECT 443.400 774.000 448.050 774.450 ;
        RECT 442.950 772.950 448.050 774.000 ;
        RECT 454.950 774.450 457.050 775.050 ;
        RECT 460.950 774.450 463.050 775.050 ;
        RECT 454.950 773.400 463.050 774.450 ;
        RECT 454.950 772.950 457.050 773.400 ;
        RECT 460.950 772.950 463.050 773.400 ;
        RECT 436.950 771.450 439.050 772.050 ;
        RECT 427.950 771.000 439.050 771.450 ;
        RECT 428.400 770.400 439.050 771.000 ;
        RECT 346.950 766.950 349.050 769.950 ;
        RECT 352.950 769.050 355.050 769.950 ;
        RECT 352.800 768.000 355.050 769.050 ;
        RECT 358.950 768.450 361.050 769.050 ;
        RECT 371.400 768.450 372.450 770.400 ;
        RECT 376.950 769.950 379.050 770.400 ;
        RECT 436.950 769.950 439.050 770.400 ;
        RECT 442.950 769.950 445.050 772.950 ;
        RECT 466.950 769.950 469.050 775.050 ;
        RECT 484.950 772.950 490.050 775.050 ;
        RECT 493.950 773.400 498.450 775.050 ;
        RECT 493.950 772.950 498.000 773.400 ;
        RECT 499.950 772.950 505.050 775.050 ;
        RECT 508.950 772.950 511.050 775.050 ;
        RECT 526.950 772.950 529.050 778.050 ;
        RECT 533.400 777.000 576.450 777.450 ;
        RECT 629.100 777.000 631.200 778.050 ;
        RECT 532.950 776.400 576.450 777.000 ;
        RECT 532.950 772.950 535.050 776.400 ;
        RECT 553.950 775.050 556.050 776.400 ;
        RECT 541.950 774.450 544.050 775.050 ;
        RECT 547.950 774.450 550.050 775.050 ;
        RECT 541.950 773.400 550.050 774.450 ;
        RECT 541.950 772.950 544.050 773.400 ;
        RECT 547.950 772.950 550.050 773.400 ;
        RECT 553.800 774.000 556.050 775.050 ;
        RECT 557.100 774.450 559.200 775.050 ;
        RECT 571.950 774.450 574.050 775.050 ;
        RECT 553.800 772.950 555.900 774.000 ;
        RECT 557.100 773.400 574.050 774.450 ;
        RECT 575.400 774.450 576.450 776.400 ;
        RECT 628.950 775.950 631.200 777.000 ;
        RECT 673.950 777.450 676.050 778.050 ;
        RECT 680.400 777.450 681.450 779.400 ;
        RECT 694.950 777.450 697.050 778.050 ;
        RECT 673.950 776.400 681.450 777.450 ;
        RECT 683.250 777.000 697.050 777.450 ;
        RECT 682.950 776.400 697.050 777.000 ;
        RECT 673.950 775.950 676.050 776.400 ;
        RECT 628.950 775.050 631.050 775.950 ;
        RECT 682.950 775.050 685.050 776.400 ;
        RECT 694.950 775.950 697.050 776.400 ;
        RECT 722.400 775.050 723.450 779.400 ;
        RECT 731.400 777.000 747.450 777.450 ;
        RECT 730.950 776.400 747.450 777.000 ;
        RECT 586.950 774.450 589.050 775.050 ;
        RECT 575.400 773.400 589.050 774.450 ;
        RECT 557.100 772.950 559.200 773.400 ;
        RECT 571.950 772.950 574.050 773.400 ;
        RECT 586.950 772.950 589.050 773.400 ;
        RECT 622.950 772.950 627.900 775.050 ;
        RECT 628.950 774.000 631.200 775.050 ;
        RECT 649.800 774.450 651.900 775.050 ;
        RECT 629.100 772.950 631.200 774.000 ;
        RECT 635.400 773.400 651.900 774.450 ;
        RECT 553.800 772.050 555.900 772.200 ;
        RECT 635.400 772.050 636.450 773.400 ;
        RECT 649.800 772.950 651.900 773.400 ;
        RECT 653.100 772.950 658.050 775.050 ;
        RECT 682.800 774.000 685.050 775.050 ;
        RECT 682.800 772.950 684.900 774.000 ;
        RECT 686.100 772.950 691.050 775.050 ;
        RECT 703.950 772.950 709.050 775.050 ;
        RECT 712.950 774.450 715.050 775.050 ;
        RECT 718.950 774.450 721.050 775.050 ;
        RECT 712.950 773.400 721.050 774.450 ;
        RECT 722.400 773.400 727.050 775.050 ;
        RECT 712.950 772.950 715.050 773.400 ;
        RECT 718.950 772.950 721.050 773.400 ;
        RECT 723.000 772.950 727.050 773.400 ;
        RECT 730.950 772.950 733.050 776.400 ;
        RECT 746.400 775.050 747.450 776.400 ;
        RECT 745.950 772.950 751.050 775.050 ;
        RECT 754.950 772.950 757.050 778.050 ;
        RECT 763.950 775.950 766.050 778.050 ;
        RECT 769.950 776.250 772.050 777.150 ;
        RECT 763.950 773.850 766.050 774.750 ;
        RECT 493.950 771.450 496.050 772.050 ;
        RECT 505.800 771.450 507.900 772.050 ;
        RECT 493.950 770.400 507.900 771.450 ;
        RECT 493.950 769.950 496.050 770.400 ;
        RECT 505.800 769.950 507.900 770.400 ;
        RECT 509.100 769.950 514.050 772.050 ;
        RECT 517.950 771.450 520.050 772.050 ;
        RECT 529.950 771.450 532.050 772.050 ;
        RECT 517.950 770.400 532.050 771.450 ;
        RECT 517.950 769.950 520.050 770.400 ;
        RECT 529.950 769.950 532.050 770.400 ;
        RECT 535.950 769.950 541.050 772.050 ;
        RECT 550.950 770.100 555.900 772.050 ;
        RECT 557.100 771.450 559.200 772.050 ;
        RECT 562.950 771.450 565.050 772.050 ;
        RECT 557.100 770.400 565.050 771.450 ;
        RECT 550.950 769.950 555.000 770.100 ;
        RECT 557.100 769.950 559.200 770.400 ;
        RECT 562.950 769.950 565.050 770.400 ;
        RECT 574.950 769.950 580.050 772.050 ;
        RECT 598.950 769.950 604.050 772.050 ;
        RECT 607.950 771.450 610.050 772.050 ;
        RECT 613.950 771.450 616.050 772.050 ;
        RECT 618.000 771.450 621.900 772.050 ;
        RECT 607.950 770.400 616.050 771.450 ;
        RECT 607.950 769.950 610.050 770.400 ;
        RECT 613.950 769.950 616.050 770.400 ;
        RECT 617.400 769.950 621.900 771.450 ;
        RECT 623.100 769.950 628.050 772.050 ;
        RECT 631.950 769.950 637.050 772.050 ;
        RECT 643.950 771.450 646.050 772.050 ;
        RECT 652.950 771.450 655.050 772.050 ;
        RECT 643.950 770.400 655.050 771.450 ;
        RECT 643.950 769.950 646.050 770.400 ;
        RECT 652.950 769.950 655.050 770.400 ;
        RECT 667.950 771.450 670.050 772.050 ;
        RECT 679.950 771.450 682.050 772.050 ;
        RECT 667.950 770.400 682.050 771.450 ;
        RECT 667.950 769.950 670.050 770.400 ;
        RECT 679.950 769.950 682.050 770.400 ;
        RECT 352.800 766.950 354.900 768.000 ;
        RECT 358.950 767.400 372.450 768.450 ;
        RECT 388.950 768.450 391.050 769.050 ;
        RECT 409.950 768.450 412.050 769.050 ;
        RECT 388.950 767.400 412.050 768.450 ;
        RECT 358.950 766.950 361.050 767.400 ;
        RECT 388.950 766.950 391.050 767.400 ;
        RECT 409.950 766.950 412.050 767.400 ;
        RECT 484.950 768.450 487.050 769.050 ;
        RECT 502.950 768.450 505.050 769.050 ;
        RECT 484.950 767.400 505.050 768.450 ;
        RECT 484.950 766.950 487.050 767.400 ;
        RECT 502.950 766.950 505.050 767.400 ;
        RECT 514.950 768.450 517.050 769.050 ;
        RECT 541.950 768.450 544.050 769.050 ;
        RECT 514.950 767.400 544.050 768.450 ;
        RECT 514.950 766.950 517.050 767.400 ;
        RECT 541.950 766.950 544.050 767.400 ;
        RECT 553.950 768.450 556.050 768.900 ;
        RECT 583.950 768.450 586.050 769.050 ;
        RECT 553.950 767.400 586.050 768.450 ;
        RECT 118.950 764.400 165.450 765.450 ;
        RECT 217.950 765.450 220.050 766.050 ;
        RECT 235.950 765.450 238.050 766.050 ;
        RECT 217.950 764.400 238.050 765.450 ;
        RECT 118.950 763.950 121.050 764.400 ;
        RECT 217.950 763.950 220.050 764.400 ;
        RECT 235.950 763.950 238.050 764.400 ;
        RECT 256.950 765.450 259.050 766.050 ;
        RECT 319.950 765.450 322.050 766.050 ;
        RECT 256.950 764.400 322.050 765.450 ;
        RECT 347.400 765.450 348.450 766.950 ;
        RECT 553.950 766.800 556.050 767.400 ;
        RECT 583.950 766.950 586.050 767.400 ;
        RECT 373.950 765.450 376.050 766.050 ;
        RECT 347.400 764.400 376.050 765.450 ;
        RECT 256.950 763.950 259.050 764.400 ;
        RECT 319.950 763.950 322.050 764.400 ;
        RECT 373.950 763.950 376.050 764.400 ;
        RECT 544.950 765.450 547.050 766.050 ;
        RECT 592.950 765.450 595.050 769.050 ;
        RECT 604.950 766.950 610.050 769.050 ;
        RECT 617.400 768.450 618.450 769.950 ;
        RECT 611.400 767.400 618.450 768.450 ;
        RECT 652.950 768.450 655.050 769.050 ;
        RECT 664.950 768.450 667.050 769.050 ;
        RECT 652.950 767.400 667.050 768.450 ;
        RECT 611.400 765.450 612.450 767.400 ;
        RECT 652.950 766.950 655.050 767.400 ;
        RECT 664.950 766.950 667.050 767.400 ;
        RECT 673.950 768.450 676.050 769.050 ;
        RECT 685.950 768.450 688.050 772.050 ;
        RECT 673.950 768.000 688.050 768.450 ;
        RECT 691.950 768.450 694.050 772.050 ;
        RECT 697.950 771.450 700.050 772.050 ;
        RECT 703.950 771.450 706.050 772.050 ;
        RECT 697.950 770.400 706.050 771.450 ;
        RECT 697.950 769.950 700.050 770.400 ;
        RECT 703.950 769.950 706.050 770.400 ;
        RECT 709.950 768.450 712.050 772.050 ;
        RECT 691.950 768.000 712.050 768.450 ;
        RECT 727.950 769.050 730.050 772.050 ;
        RECT 733.950 769.950 739.050 772.050 ;
        RECT 727.950 768.450 733.050 769.050 ;
        RECT 745.950 768.450 748.050 772.050 ;
        RECT 727.950 768.000 748.050 768.450 ;
        RECT 673.950 767.400 687.450 768.000 ;
        RECT 692.400 767.400 711.450 768.000 ;
        RECT 728.400 767.400 747.450 768.000 ;
        RECT 673.950 766.950 676.050 767.400 ;
        RECT 729.000 766.950 733.050 767.400 ;
        RECT 751.950 766.950 754.050 772.050 ;
        RECT 776.850 766.050 778.050 784.950 ;
        RECT 779.850 780.750 781.050 784.950 ;
        RECT 778.950 778.650 781.050 780.750 ;
        RECT 779.850 766.050 781.050 778.650 ;
        RECT 782.850 766.050 784.050 784.950 ;
        RECT 790.950 782.400 793.050 784.500 ;
        RECT 796.050 783.300 798.150 785.400 ;
        RECT 799.950 783.300 802.050 785.400 ;
        RECT 802.950 783.300 805.050 785.400 ;
        RECT 805.950 785.100 808.050 787.200 ;
        RECT 790.950 776.250 792.150 782.400 ;
        RECT 790.950 774.150 793.050 776.250 ;
        RECT 787.950 770.250 790.050 771.150 ;
        RECT 790.950 770.250 792.150 774.150 ;
        RECT 796.950 773.550 798.150 783.300 ;
        RECT 800.850 781.350 802.050 783.300 ;
        RECT 799.950 779.250 802.050 781.350 ;
        RECT 795.150 771.450 798.150 773.550 ;
        RECT 787.950 766.950 790.050 769.050 ;
        RECT 544.950 765.000 595.050 765.450 ;
        RECT 544.950 764.400 594.450 765.000 ;
        RECT 599.400 764.400 612.450 765.450 ;
        RECT 613.950 765.450 616.050 766.050 ;
        RECT 622.950 765.450 625.050 766.050 ;
        RECT 613.950 764.400 625.050 765.450 ;
        RECT 544.950 763.950 547.050 764.400 ;
        RECT 599.400 763.050 600.450 764.400 ;
        RECT 613.950 763.950 616.050 764.400 ;
        RECT 622.950 763.950 625.050 764.400 ;
        RECT 637.950 765.450 640.050 766.050 ;
        RECT 658.950 765.450 661.050 766.050 ;
        RECT 637.950 764.400 661.050 765.450 ;
        RECT 637.950 763.950 640.050 764.400 ;
        RECT 658.950 763.950 661.050 764.400 ;
        RECT 688.950 765.450 691.050 766.050 ;
        RECT 709.950 765.450 712.050 766.050 ;
        RECT 715.950 765.450 718.050 766.050 ;
        RECT 688.950 764.400 718.050 765.450 ;
        RECT 688.950 763.950 691.050 764.400 ;
        RECT 709.950 763.950 712.050 764.400 ;
        RECT 715.950 763.950 718.050 764.400 ;
        RECT 748.950 765.450 751.050 766.050 ;
        RECT 757.950 765.450 760.050 766.050 ;
        RECT 748.950 764.400 760.050 765.450 ;
        RECT 748.950 763.950 751.050 764.400 ;
        RECT 757.950 763.950 760.050 764.400 ;
        RECT 775.950 763.950 778.050 766.050 ;
        RECT 778.950 763.950 781.050 766.050 ;
        RECT 781.950 763.950 784.050 766.050 ;
        RECT 791.250 765.750 792.150 770.250 ;
        RECT 790.950 765.600 792.150 765.750 ;
        RECT 796.950 765.600 798.150 771.450 ;
        RECT 800.550 765.600 802.050 779.250 ;
        RECT 803.850 765.600 805.050 783.300 ;
        RECT 806.250 781.350 807.450 785.100 ;
        RECT 823.950 783.450 826.050 784.050 ;
        RECT 829.950 783.450 832.050 784.050 ;
        RECT 823.950 782.400 832.050 783.450 ;
        RECT 823.950 781.950 826.050 782.400 ;
        RECT 829.950 781.950 832.050 782.400 ;
        RECT 805.950 779.250 808.050 781.350 ;
        RECT 806.250 765.600 807.450 779.250 ;
        RECT 814.950 772.950 817.050 775.050 ;
        RECT 818.250 772.950 819.150 775.050 ;
        RECT 824.850 772.950 825.750 775.050 ;
        RECT 826.950 772.950 829.050 775.050 ;
        RECT 844.950 772.950 850.050 775.050 ;
        RECT 823.950 768.450 826.050 769.050 ;
        RECT 829.950 768.450 832.050 769.050 ;
        RECT 823.950 767.400 832.050 768.450 ;
        RECT 823.950 766.950 826.050 767.400 ;
        RECT 829.950 766.950 832.050 767.400 ;
        RECT 790.950 763.500 793.050 765.600 ;
        RECT 796.050 763.500 798.150 765.600 ;
        RECT 799.950 763.500 802.050 765.600 ;
        RECT 802.950 763.500 805.050 765.600 ;
        RECT 805.950 763.500 808.050 765.600 ;
        RECT 838.950 763.950 841.050 769.050 ;
        RECT 13.950 762.450 16.050 763.050 ;
        RECT 34.950 762.450 37.050 763.050 ;
        RECT 13.950 761.400 37.050 762.450 ;
        RECT 13.950 760.950 16.050 761.400 ;
        RECT 34.950 760.950 37.050 761.400 ;
        RECT 100.950 762.450 103.050 763.050 ;
        RECT 115.950 762.450 118.050 763.050 ;
        RECT 100.950 761.400 118.050 762.450 ;
        RECT 100.950 760.950 103.050 761.400 ;
        RECT 115.950 760.950 118.050 761.400 ;
        RECT 274.950 762.450 277.050 763.050 ;
        RECT 286.950 762.450 289.050 763.050 ;
        RECT 340.950 762.450 343.050 763.050 ;
        RECT 274.950 761.400 343.050 762.450 ;
        RECT 274.950 760.950 277.050 761.400 ;
        RECT 286.950 760.950 289.050 761.400 ;
        RECT 340.950 760.950 343.050 761.400 ;
        RECT 502.950 762.450 505.050 763.050 ;
        RECT 517.950 762.450 520.050 763.050 ;
        RECT 502.950 761.400 520.050 762.450 ;
        RECT 502.950 760.950 505.050 761.400 ;
        RECT 517.950 760.950 520.050 761.400 ;
        RECT 550.950 762.450 553.050 763.050 ;
        RECT 598.800 762.450 600.900 763.050 ;
        RECT 550.950 761.400 600.900 762.450 ;
        RECT 550.950 760.950 553.050 761.400 ;
        RECT 598.800 760.950 600.900 761.400 ;
        RECT 602.100 762.450 604.200 763.050 ;
        RECT 718.950 762.450 721.050 763.200 ;
        RECT 751.950 762.450 754.050 763.050 ;
        RECT 602.100 761.400 672.450 762.450 ;
        RECT 602.100 760.950 604.200 761.400 ;
        RECT 61.950 759.450 64.050 760.050 ;
        RECT 193.950 759.450 196.050 760.050 ;
        RECT 61.950 758.400 196.050 759.450 ;
        RECT 61.950 757.950 64.050 758.400 ;
        RECT 193.950 757.950 196.050 758.400 ;
        RECT 421.950 759.450 424.050 760.050 ;
        RECT 469.950 759.450 472.050 760.050 ;
        RECT 421.950 758.400 472.050 759.450 ;
        RECT 421.950 757.950 424.050 758.400 ;
        RECT 469.950 757.950 472.050 758.400 ;
        RECT 571.950 759.450 574.050 760.050 ;
        RECT 583.950 759.450 586.050 760.050 ;
        RECT 628.950 759.450 631.050 760.050 ;
        RECT 571.950 758.400 631.050 759.450 ;
        RECT 571.950 757.950 574.050 758.400 ;
        RECT 583.950 757.950 586.050 758.400 ;
        RECT 628.950 757.950 631.050 758.400 ;
        RECT 640.950 759.450 643.050 760.050 ;
        RECT 664.950 759.450 667.050 760.050 ;
        RECT 640.950 758.400 667.050 759.450 ;
        RECT 671.400 759.450 672.450 761.400 ;
        RECT 718.950 761.400 754.050 762.450 ;
        RECT 718.950 761.100 721.050 761.400 ;
        RECT 751.950 760.950 754.050 761.400 ;
        RECT 811.950 762.450 814.050 763.050 ;
        RECT 838.950 762.450 841.050 763.050 ;
        RECT 811.950 761.400 841.050 762.450 ;
        RECT 811.950 760.950 814.050 761.400 ;
        RECT 838.950 760.950 841.050 761.400 ;
        RECT 718.950 759.450 721.050 759.900 ;
        RECT 671.400 758.400 721.050 759.450 ;
        RECT 640.950 757.950 643.050 758.400 ;
        RECT 664.950 757.950 667.050 758.400 ;
        RECT 718.950 757.800 721.050 758.400 ;
        RECT 727.950 759.450 730.050 760.050 ;
        RECT 772.950 759.450 775.050 760.050 ;
        RECT 727.950 758.400 775.050 759.450 ;
        RECT 727.950 757.950 730.050 758.400 ;
        RECT 772.950 757.950 775.050 758.400 ;
        RECT 109.950 756.450 112.050 757.050 ;
        RECT 127.950 756.450 130.050 757.050 ;
        RECT 208.950 756.450 211.050 757.050 ;
        RECT 109.950 755.400 211.050 756.450 ;
        RECT 109.950 754.950 112.050 755.400 ;
        RECT 127.950 754.950 130.050 755.400 ;
        RECT 208.950 754.950 211.050 755.400 ;
        RECT 415.950 756.450 418.050 757.050 ;
        RECT 514.950 756.450 517.050 757.050 ;
        RECT 415.950 755.400 517.050 756.450 ;
        RECT 415.950 754.950 418.050 755.400 ;
        RECT 514.950 754.950 517.050 755.400 ;
        RECT 589.950 756.450 592.050 757.050 ;
        RECT 634.950 756.450 637.050 757.050 ;
        RECT 763.950 756.450 766.050 757.050 ;
        RECT 589.950 755.400 637.050 756.450 ;
        RECT 589.950 754.950 592.050 755.400 ;
        RECT 634.950 754.950 637.050 755.400 ;
        RECT 728.400 755.400 766.050 756.450 ;
        RECT 22.950 753.450 25.050 754.050 ;
        RECT 28.950 753.450 31.050 754.050 ;
        RECT 22.950 752.400 31.050 753.450 ;
        RECT 22.950 751.950 25.050 752.400 ;
        RECT 28.950 751.950 31.050 752.400 ;
        RECT 85.950 753.450 88.050 754.050 ;
        RECT 91.950 753.450 94.050 754.050 ;
        RECT 85.950 752.400 94.050 753.450 ;
        RECT 85.950 751.950 88.050 752.400 ;
        RECT 91.950 751.950 94.050 752.400 ;
        RECT 175.950 751.950 181.050 754.050 ;
        RECT 379.950 753.450 382.050 754.050 ;
        RECT 397.950 753.450 400.050 754.050 ;
        RECT 379.950 752.400 400.050 753.450 ;
        RECT 379.950 751.950 382.050 752.400 ;
        RECT 397.950 751.950 400.050 752.400 ;
        RECT 418.950 753.450 421.050 754.050 ;
        RECT 433.950 753.450 436.050 754.050 ;
        RECT 418.950 752.400 436.050 753.450 ;
        RECT 418.950 751.950 421.050 752.400 ;
        RECT 433.950 751.950 436.050 752.400 ;
        RECT 601.950 753.450 604.050 754.050 ;
        RECT 643.950 753.450 646.050 754.050 ;
        RECT 601.950 752.400 646.050 753.450 ;
        RECT 601.950 751.950 604.050 752.400 ;
        RECT 643.950 751.950 646.050 752.400 ;
        RECT 658.950 753.450 661.050 754.050 ;
        RECT 676.950 753.450 679.050 754.050 ;
        RECT 694.950 753.450 697.050 754.050 ;
        RECT 658.950 752.400 679.050 753.450 ;
        RECT 658.950 751.950 661.050 752.400 ;
        RECT 676.950 751.950 679.050 752.400 ;
        RECT 689.400 752.400 697.050 753.450 ;
        RECT 46.950 750.450 49.050 751.050 ;
        RECT 64.950 750.450 67.050 751.050 ;
        RECT 46.950 749.400 67.050 750.450 ;
        RECT 46.950 748.950 49.050 749.400 ;
        RECT 64.950 748.950 67.050 749.400 ;
        RECT 157.950 750.450 160.050 751.050 ;
        RECT 169.950 750.450 172.050 751.050 ;
        RECT 202.950 750.450 205.050 751.050 ;
        RECT 313.950 750.450 316.050 751.050 ;
        RECT 346.950 750.450 349.050 751.050 ;
        RECT 157.950 750.000 228.450 750.450 ;
        RECT 157.950 749.400 229.050 750.000 ;
        RECT 157.950 748.950 160.050 749.400 ;
        RECT 169.950 748.950 172.050 749.400 ;
        RECT 202.950 748.950 205.050 749.400 ;
        RECT 22.950 747.450 25.050 748.050 ;
        RECT 22.950 746.400 36.600 747.450 ;
        RECT 38.400 747.000 63.450 747.450 ;
        RECT 22.950 745.950 25.050 746.400 ;
        RECT 25.950 744.450 28.050 745.050 ;
        RECT 31.950 744.450 34.050 745.050 ;
        RECT 25.950 743.400 34.050 744.450 ;
        RECT 25.950 742.950 28.050 743.400 ;
        RECT 31.950 742.950 34.050 743.400 ;
        RECT 35.550 742.050 36.600 746.400 ;
        RECT 37.950 746.400 63.450 747.000 ;
        RECT 37.950 744.450 40.050 746.400 ;
        RECT 37.950 743.400 45.450 744.450 ;
        RECT 37.950 742.950 40.050 743.400 ;
        RECT 4.950 741.450 7.050 742.050 ;
        RECT 10.950 741.450 16.050 742.050 ;
        RECT 4.950 740.400 16.050 741.450 ;
        RECT 4.950 739.950 7.050 740.400 ;
        RECT 10.950 739.950 16.050 740.400 ;
        RECT 28.950 739.950 33.900 742.050 ;
        RECT 35.100 739.950 37.200 742.050 ;
        RECT 44.400 741.450 45.450 743.400 ;
        RECT 46.950 742.950 51.900 745.050 ;
        RECT 53.100 744.450 55.200 745.050 ;
        RECT 58.950 744.450 61.050 745.050 ;
        RECT 53.100 743.400 61.050 744.450 ;
        RECT 62.400 744.450 63.450 746.400 ;
        RECT 127.950 745.950 133.050 748.050 ;
        RECT 160.950 747.450 163.050 748.050 ;
        RECT 175.950 747.450 178.050 748.050 ;
        RECT 181.950 747.450 184.050 748.050 ;
        RECT 199.950 747.450 202.050 748.050 ;
        RECT 160.950 746.400 202.050 747.450 ;
        RECT 160.950 745.950 163.050 746.400 ;
        RECT 175.950 745.950 178.050 746.400 ;
        RECT 181.950 745.950 184.050 746.400 ;
        RECT 199.950 745.950 202.050 746.400 ;
        RECT 226.950 745.950 229.050 749.400 ;
        RECT 313.950 749.400 349.050 750.450 ;
        RECT 313.950 748.950 316.050 749.400 ;
        RECT 67.950 744.450 70.050 745.050 ;
        RECT 62.400 743.400 70.050 744.450 ;
        RECT 53.100 742.950 55.200 743.400 ;
        RECT 58.950 742.950 61.050 743.400 ;
        RECT 67.950 742.950 70.050 743.400 ;
        RECT 73.950 742.950 79.050 745.050 ;
        RECT 85.950 744.450 88.050 745.050 ;
        RECT 94.950 744.450 97.050 745.050 ;
        RECT 85.950 743.400 97.050 744.450 ;
        RECT 85.950 742.950 88.050 743.400 ;
        RECT 94.950 742.950 97.050 743.400 ;
        RECT 145.950 744.450 148.050 745.050 ;
        RECT 184.950 744.450 187.050 745.050 ;
        RECT 202.950 744.450 205.050 745.050 ;
        RECT 145.950 743.400 156.450 744.450 ;
        RECT 145.950 742.950 148.050 743.400 ;
        RECT 49.950 741.450 52.050 742.050 ;
        RECT 44.400 740.400 52.050 741.450 ;
        RECT 49.950 739.950 52.050 740.400 ;
        RECT 10.950 733.950 13.050 739.050 ;
        RECT 16.950 735.450 19.050 739.050 ;
        RECT 25.950 738.450 28.050 739.050 ;
        RECT 52.950 738.450 55.050 739.050 ;
        RECT 25.950 737.400 55.050 738.450 ;
        RECT 55.950 738.450 58.050 742.050 ;
        RECT 70.950 739.950 76.050 742.050 ;
        RECT 79.950 739.950 85.050 742.050 ;
        RECT 91.950 739.950 97.050 742.050 ;
        RECT 100.950 739.050 103.050 742.050 ;
        RECT 106.950 741.450 109.050 742.050 ;
        RECT 112.950 741.450 115.050 742.050 ;
        RECT 106.950 740.400 115.050 741.450 ;
        RECT 106.950 739.950 109.050 740.400 ;
        RECT 112.950 739.950 115.050 740.400 ;
        RECT 133.950 741.450 136.050 742.050 ;
        RECT 142.800 741.450 144.900 742.050 ;
        RECT 133.950 740.400 144.900 741.450 ;
        RECT 133.950 739.950 136.050 740.400 ;
        RECT 142.800 739.950 144.900 740.400 ;
        RECT 145.800 741.000 147.900 742.050 ;
        RECT 145.800 739.950 148.050 741.000 ;
        RECT 149.100 739.950 154.050 742.050 ;
        RECT 155.400 741.450 156.450 743.400 ;
        RECT 184.950 743.400 205.050 744.450 ;
        RECT 184.950 742.950 187.050 743.400 ;
        RECT 202.950 742.950 205.050 743.400 ;
        RECT 166.950 741.450 169.050 742.050 ;
        RECT 155.400 740.400 169.050 741.450 ;
        RECT 166.950 739.950 169.050 740.400 ;
        RECT 172.950 741.450 175.050 742.050 ;
        RECT 190.950 741.450 193.050 742.050 ;
        RECT 172.950 740.400 193.050 741.450 ;
        RECT 172.950 739.950 175.050 740.400 ;
        RECT 190.950 739.950 193.050 740.400 ;
        RECT 208.950 739.950 211.050 745.050 ;
        RECT 223.950 739.950 226.050 745.050 ;
        RECT 229.950 739.950 232.050 745.050 ;
        RECT 256.950 742.950 259.050 748.050 ;
        RECT 304.950 747.450 307.050 748.050 ;
        RECT 319.950 747.450 322.050 748.050 ;
        RECT 304.950 746.400 322.050 747.450 ;
        RECT 304.950 745.950 307.050 746.400 ;
        RECT 319.950 745.950 322.050 746.400 ;
        RECT 334.950 745.950 337.050 749.400 ;
        RECT 346.950 748.950 349.050 749.400 ;
        RECT 358.950 750.450 361.050 751.050 ;
        RECT 391.950 750.450 394.050 751.050 ;
        RECT 358.950 749.400 394.050 750.450 ;
        RECT 358.950 748.950 361.050 749.400 ;
        RECT 391.950 748.950 394.050 749.400 ;
        RECT 301.950 744.450 304.050 745.050 ;
        RECT 313.950 744.450 316.050 745.050 ;
        RECT 275.400 744.000 285.450 744.450 ;
        RECT 275.400 743.400 286.050 744.000 ;
        RECT 244.950 741.450 247.050 742.050 ;
        RECT 256.950 741.450 259.050 742.050 ;
        RECT 244.950 740.400 259.050 741.450 ;
        RECT 244.950 739.950 247.050 740.400 ;
        RECT 256.950 739.950 259.050 740.400 ;
        RECT 262.950 741.450 265.050 742.050 ;
        RECT 275.400 741.450 276.450 743.400 ;
        RECT 262.950 740.400 276.450 741.450 ;
        RECT 262.950 739.950 265.050 740.400 ;
        RECT 88.950 738.450 91.050 739.050 ;
        RECT 55.950 738.000 91.050 738.450 ;
        RECT 56.400 737.400 91.050 738.000 ;
        RECT 25.950 736.950 28.050 737.400 ;
        RECT 52.950 736.950 55.050 737.400 ;
        RECT 88.950 736.950 91.050 737.400 ;
        RECT 97.800 738.000 99.900 739.050 ;
        RECT 100.950 738.000 103.200 739.050 ;
        RECT 97.800 736.950 100.050 738.000 ;
        RECT 101.100 736.950 103.200 738.000 ;
        RECT 97.950 736.050 100.050 736.950 ;
        RECT 76.950 735.450 79.050 736.050 ;
        RECT 97.800 735.450 100.050 736.050 ;
        RECT 16.950 735.000 100.050 735.450 ;
        RECT 103.950 735.450 106.050 736.050 ;
        RECT 109.950 735.450 112.050 739.050 ;
        RECT 103.950 735.000 112.050 735.450 ;
        RECT 115.950 735.450 118.050 739.050 ;
        RECT 145.950 736.950 148.050 739.950 ;
        RECT 277.950 739.050 280.050 742.050 ;
        RECT 283.950 739.950 286.050 743.400 ;
        RECT 301.950 743.400 316.050 744.450 ;
        RECT 301.950 742.950 304.050 743.400 ;
        RECT 313.950 742.950 316.050 743.400 ;
        RECT 325.950 744.450 328.050 745.050 ;
        RECT 331.800 744.450 333.900 745.050 ;
        RECT 325.950 743.400 333.900 744.450 ;
        RECT 325.950 742.950 328.050 743.400 ;
        RECT 331.800 742.950 333.900 743.400 ;
        RECT 335.100 742.950 339.900 745.050 ;
        RECT 341.100 744.450 343.200 745.050 ;
        RECT 355.800 744.450 357.900 745.050 ;
        RECT 341.100 743.400 357.900 744.450 ;
        RECT 341.100 742.950 343.200 743.400 ;
        RECT 355.800 742.950 357.900 743.400 ;
        RECT 358.800 744.000 360.900 745.050 ;
        RECT 362.100 744.450 364.200 745.050 ;
        RECT 370.950 744.450 373.050 748.050 ;
        RECT 391.950 747.450 394.050 748.050 ;
        RECT 403.950 747.450 406.050 748.050 ;
        RECT 391.950 746.400 406.050 747.450 ;
        RECT 391.950 745.950 394.050 746.400 ;
        RECT 403.950 745.950 406.050 746.400 ;
        RECT 418.950 747.450 421.050 748.050 ;
        RECT 418.950 747.000 489.600 747.450 ;
        RECT 418.950 746.400 490.050 747.000 ;
        RECT 418.950 745.950 421.050 746.400 ;
        RECT 487.950 745.050 490.050 746.400 ;
        RECT 502.950 745.950 505.050 751.050 ;
        RECT 508.950 750.450 511.050 751.050 ;
        RECT 562.950 750.450 565.050 751.050 ;
        RECT 508.950 749.400 565.050 750.450 ;
        RECT 508.950 748.950 511.050 749.400 ;
        RECT 562.950 748.950 565.050 749.400 ;
        RECT 397.800 744.450 399.900 745.050 ;
        RECT 358.800 742.950 361.050 744.000 ;
        RECT 362.100 743.400 399.900 744.450 ;
        RECT 362.100 742.950 364.200 743.400 ;
        RECT 397.800 742.950 399.900 743.400 ;
        RECT 401.100 742.950 405.900 745.050 ;
        RECT 407.100 744.450 409.200 745.050 ;
        RECT 415.950 744.450 418.050 745.050 ;
        RECT 407.100 743.400 418.050 744.450 ;
        RECT 407.100 742.950 409.200 743.400 ;
        RECT 415.950 742.950 418.050 743.400 ;
        RECT 433.950 744.450 436.050 745.050 ;
        RECT 442.800 744.450 444.900 745.050 ;
        RECT 433.950 743.400 444.900 744.450 ;
        RECT 433.950 742.950 436.050 743.400 ;
        RECT 442.800 742.950 444.900 743.400 ;
        RECT 446.100 742.950 451.050 745.050 ;
        RECT 481.950 742.950 486.900 745.050 ;
        RECT 487.950 744.000 490.200 745.050 ;
        RECT 488.100 742.950 490.200 744.000 ;
        RECT 508.950 744.450 511.050 745.050 ;
        RECT 514.950 744.450 517.050 745.050 ;
        RECT 508.950 743.400 517.050 744.450 ;
        RECT 508.950 742.950 511.050 743.400 ;
        RECT 514.950 742.950 517.050 743.400 ;
        RECT 520.950 742.950 523.050 748.050 ;
        RECT 538.950 747.450 541.050 748.050 ;
        RECT 527.400 747.000 541.050 747.450 ;
        RECT 526.950 746.400 541.050 747.000 ;
        RECT 526.950 742.950 529.050 746.400 ;
        RECT 538.950 745.950 541.050 746.400 ;
        RECT 574.950 747.450 577.050 748.050 ;
        RECT 583.950 747.450 586.050 748.050 ;
        RECT 574.950 746.400 586.050 747.450 ;
        RECT 574.950 745.950 577.050 746.400 ;
        RECT 583.950 745.950 586.050 746.400 ;
        RECT 592.950 745.950 595.050 751.050 ;
        RECT 613.950 750.450 616.050 751.050 ;
        RECT 689.400 750.450 690.450 752.400 ;
        RECT 694.950 751.950 697.050 752.400 ;
        RECT 718.950 753.450 721.050 754.050 ;
        RECT 728.400 753.450 729.450 755.400 ;
        RECT 763.950 754.950 766.050 755.400 ;
        RECT 832.950 756.450 835.050 757.050 ;
        RECT 853.950 756.450 856.050 757.050 ;
        RECT 832.950 755.400 856.050 756.450 ;
        RECT 832.950 754.950 835.050 755.400 ;
        RECT 853.950 754.950 856.050 755.400 ;
        RECT 718.950 752.400 729.450 753.450 ;
        RECT 781.950 753.450 784.050 754.050 ;
        RECT 793.950 753.450 796.050 754.050 ;
        RECT 781.950 752.400 796.050 753.450 ;
        RECT 718.950 751.950 721.050 752.400 ;
        RECT 781.950 751.950 784.050 752.400 ;
        RECT 793.950 751.950 796.050 752.400 ;
        RECT 613.950 749.400 690.450 750.450 ;
        RECT 712.950 749.400 715.050 751.500 ;
        RECT 733.950 749.400 736.050 751.500 ;
        RECT 613.950 748.950 616.050 749.400 ;
        RECT 625.800 747.450 627.900 748.050 ;
        RECT 620.550 747.000 627.900 747.450 ;
        RECT 619.950 746.400 627.900 747.000 ;
        RECT 619.950 745.050 622.050 746.400 ;
        RECT 625.800 745.950 627.900 746.400 ;
        RECT 629.100 747.450 631.200 748.050 ;
        RECT 634.950 747.450 637.050 748.050 ;
        RECT 629.100 746.400 637.050 747.450 ;
        RECT 629.100 745.950 631.200 746.400 ;
        RECT 634.950 745.950 637.050 746.400 ;
        RECT 649.950 747.450 652.050 748.050 ;
        RECT 658.800 747.450 660.900 748.050 ;
        RECT 649.950 747.000 660.900 747.450 ;
        RECT 662.100 747.450 664.200 748.050 ;
        RECT 670.950 747.450 673.050 748.050 ;
        RECT 649.950 746.400 661.050 747.000 ;
        RECT 649.950 745.950 652.050 746.400 ;
        RECT 658.800 745.950 661.050 746.400 ;
        RECT 662.100 746.400 673.050 747.450 ;
        RECT 662.100 745.950 664.200 746.400 ;
        RECT 670.950 745.950 673.050 746.400 ;
        RECT 676.800 747.000 678.900 748.050 ;
        RECT 680.100 747.450 682.200 748.050 ;
        RECT 685.950 747.450 688.050 748.050 ;
        RECT 676.800 745.950 679.050 747.000 ;
        RECT 680.100 746.400 688.050 747.450 ;
        RECT 680.100 745.950 682.200 746.400 ;
        RECT 685.950 745.950 688.050 746.400 ;
        RECT 571.950 744.450 574.050 745.050 ;
        RECT 530.400 743.400 574.050 744.450 ;
        RECT 301.950 741.450 304.050 742.050 ;
        RECT 316.950 741.450 319.050 742.050 ;
        RECT 287.400 740.400 319.050 741.450 ;
        RECT 151.950 735.450 154.050 739.050 ;
        RECT 157.950 738.450 160.050 739.050 ;
        RECT 163.950 738.450 166.050 739.050 ;
        RECT 157.950 737.400 166.050 738.450 ;
        RECT 157.950 736.950 160.050 737.400 ;
        RECT 163.950 736.950 166.050 737.400 ;
        RECT 169.950 738.450 172.050 739.050 ;
        RECT 175.950 738.450 178.050 739.050 ;
        RECT 169.950 737.400 178.050 738.450 ;
        RECT 169.950 736.950 172.050 737.400 ;
        RECT 175.950 736.950 178.050 737.400 ;
        RECT 115.950 735.000 154.050 735.450 ;
        RECT 16.950 734.400 99.900 735.000 ;
        RECT 16.950 733.950 19.050 734.400 ;
        RECT 76.950 733.950 79.050 734.400 ;
        RECT 97.800 733.950 99.900 734.400 ;
        RECT 103.950 734.400 111.450 735.000 ;
        RECT 116.400 734.400 153.450 735.000 ;
        RECT 103.950 733.950 106.050 734.400 ;
        RECT 205.950 733.950 208.050 739.050 ;
        RECT 211.950 733.950 214.050 739.050 ;
        RECT 235.950 738.450 238.050 739.050 ;
        RECT 241.950 738.450 244.050 739.050 ;
        RECT 235.950 737.400 244.050 738.450 ;
        RECT 235.950 736.950 238.050 737.400 ;
        RECT 241.950 736.950 244.050 737.400 ;
        RECT 241.950 735.450 244.050 736.050 ;
        RECT 247.950 735.450 250.050 739.050 ;
        RECT 262.950 738.450 265.050 739.050 ;
        RECT 271.950 738.450 274.050 739.050 ;
        RECT 262.950 737.400 274.050 738.450 ;
        RECT 262.950 736.950 265.050 737.400 ;
        RECT 271.950 736.950 274.050 737.400 ;
        RECT 277.800 738.000 280.050 739.050 ;
        RECT 281.100 738.450 283.200 739.050 ;
        RECT 287.400 738.450 288.450 740.400 ;
        RECT 301.950 739.950 304.050 740.400 ;
        RECT 316.950 739.950 319.050 740.400 ;
        RECT 277.800 736.950 279.900 738.000 ;
        RECT 281.100 737.400 288.450 738.450 ;
        RECT 281.100 736.950 283.200 737.400 ;
        RECT 310.950 736.950 316.050 739.050 ;
        RECT 241.950 735.000 250.050 735.450 ;
        RECT 277.950 735.450 280.050 736.050 ;
        RECT 289.950 735.450 292.050 736.050 ;
        RECT 241.950 734.400 249.450 735.000 ;
        RECT 277.950 734.400 292.050 735.450 ;
        RECT 319.950 735.450 322.050 739.050 ;
        RECT 352.950 738.450 355.050 742.050 ;
        RECT 358.950 739.950 361.050 742.950 ;
        RECT 391.950 739.950 397.050 742.050 ;
        RECT 421.950 741.450 424.050 742.050 ;
        RECT 430.950 741.450 433.050 742.050 ;
        RECT 421.950 740.400 433.050 741.450 ;
        RECT 421.950 739.950 424.050 740.400 ;
        RECT 430.950 739.950 433.050 740.400 ;
        RECT 436.950 739.950 442.050 742.050 ;
        RECT 445.950 741.450 448.050 742.050 ;
        RECT 460.950 741.450 463.050 742.050 ;
        RECT 478.950 741.450 481.050 742.050 ;
        RECT 445.950 740.400 481.050 741.450 ;
        RECT 445.950 739.950 448.050 740.400 ;
        RECT 460.950 739.950 463.050 740.400 ;
        RECT 478.950 739.950 481.050 740.400 ;
        RECT 388.950 738.450 391.050 739.050 ;
        RECT 352.950 738.000 391.050 738.450 ;
        RECT 353.400 737.400 391.050 738.000 ;
        RECT 388.950 736.950 391.050 737.400 ;
        RECT 400.950 738.450 403.050 739.050 ;
        RECT 418.950 738.450 421.050 739.050 ;
        RECT 400.950 737.400 421.050 738.450 ;
        RECT 400.950 736.950 403.050 737.400 ;
        RECT 418.950 736.950 421.050 737.400 ;
        RECT 424.950 736.950 430.050 739.050 ;
        RECT 355.950 735.450 358.050 736.050 ;
        RECT 364.950 735.450 367.050 736.050 ;
        RECT 319.950 735.000 367.050 735.450 ;
        RECT 320.400 734.400 367.050 735.000 ;
        RECT 241.950 733.950 244.050 734.400 ;
        RECT 277.950 733.950 280.050 734.400 ;
        RECT 289.950 733.950 292.050 734.400 ;
        RECT 355.950 733.950 358.050 734.400 ;
        RECT 364.950 733.950 367.050 734.400 ;
        RECT 457.950 733.950 460.050 739.050 ;
        RECT 463.950 733.950 466.050 739.050 ;
        RECT 484.950 738.450 487.050 742.050 ;
        RECT 502.950 739.950 508.050 742.050 ;
        RECT 517.950 738.450 520.050 742.050 ;
        RECT 523.950 741.450 529.050 742.050 ;
        RECT 530.400 741.450 531.450 743.400 ;
        RECT 560.400 742.050 561.450 743.400 ;
        RECT 571.950 742.950 574.050 743.400 ;
        RECT 577.950 742.950 583.050 745.050 ;
        RECT 523.950 740.400 531.450 741.450 ;
        RECT 532.950 741.450 535.050 742.050 ;
        RECT 538.950 741.450 541.050 742.050 ;
        RECT 532.950 740.400 541.050 741.450 ;
        RECT 523.950 739.950 529.050 740.400 ;
        RECT 532.950 739.950 535.050 740.400 ;
        RECT 538.950 739.950 541.050 740.400 ;
        RECT 556.950 739.950 561.450 742.050 ;
        RECT 562.950 739.950 568.050 742.050 ;
        RECT 589.950 739.950 592.050 745.050 ;
        RECT 595.950 744.450 598.050 745.050 ;
        RECT 601.950 744.450 604.050 745.050 ;
        RECT 595.950 743.400 604.050 744.450 ;
        RECT 595.950 742.950 598.050 743.400 ;
        RECT 601.950 742.950 604.050 743.400 ;
        RECT 613.950 742.950 618.900 745.050 ;
        RECT 619.950 744.000 622.200 745.050 ;
        RECT 620.100 742.950 622.200 744.000 ;
        RECT 658.950 742.950 661.050 745.950 ;
        RECT 676.950 745.050 679.050 745.950 ;
        RECT 664.950 744.450 667.050 745.050 ;
        RECT 673.800 744.450 675.900 745.050 ;
        RECT 664.950 743.400 675.900 744.450 ;
        RECT 676.950 744.000 679.200 745.050 ;
        RECT 484.950 738.000 520.050 738.450 ;
        RECT 485.400 737.400 520.050 738.000 ;
        RECT 517.950 736.950 520.050 737.400 ;
        RECT 520.950 735.450 523.050 736.050 ;
        RECT 535.950 735.450 538.050 739.050 ;
        RECT 541.950 738.450 544.050 739.050 ;
        RECT 547.950 738.450 550.050 739.050 ;
        RECT 541.950 737.400 550.050 738.450 ;
        RECT 560.400 738.450 561.450 739.950 ;
        RECT 595.950 738.450 598.050 739.050 ;
        RECT 560.400 737.400 598.050 738.450 ;
        RECT 541.950 736.950 544.050 737.400 ;
        RECT 547.950 736.950 550.050 737.400 ;
        RECT 595.950 736.950 598.050 737.400 ;
        RECT 610.950 736.950 613.050 742.050 ;
        RECT 616.950 738.450 619.050 742.050 ;
        RECT 643.950 739.950 649.050 742.050 ;
        RECT 664.950 739.950 667.050 743.400 ;
        RECT 673.800 742.950 675.900 743.400 ;
        RECT 677.100 742.950 679.200 744.000 ;
        RECT 682.950 739.950 685.050 745.050 ;
        RECT 691.950 744.450 694.050 745.050 ;
        RECT 709.950 744.450 712.050 745.050 ;
        RECT 691.950 743.400 712.050 744.450 ;
        RECT 691.950 742.950 694.050 743.400 ;
        RECT 700.950 739.950 706.050 742.050 ;
        RECT 709.950 739.950 712.050 743.400 ;
        RECT 634.950 738.450 637.050 739.050 ;
        RECT 616.950 738.000 637.050 738.450 ;
        RECT 617.400 737.400 637.050 738.000 ;
        RECT 634.950 736.950 637.050 737.400 ;
        RECT 694.950 736.950 700.050 739.050 ;
        RECT 703.950 736.950 706.050 739.050 ;
        RECT 713.850 737.400 715.050 749.400 ;
        RECT 718.950 742.950 724.050 745.050 ;
        RECT 727.950 739.950 730.050 745.050 ;
        RECT 520.950 735.000 538.050 735.450 ;
        RECT 565.950 735.450 568.050 736.050 ;
        RECT 598.950 735.450 601.050 736.050 ;
        RECT 520.950 734.400 537.450 735.000 ;
        RECT 565.950 734.400 601.050 735.450 ;
        RECT 520.950 733.950 523.050 734.400 ;
        RECT 565.950 733.950 568.050 734.400 ;
        RECT 598.950 733.950 601.050 734.400 ;
        RECT 616.950 735.450 619.050 736.050 ;
        RECT 625.950 735.450 628.050 736.050 ;
        RECT 616.950 734.400 628.050 735.450 ;
        RECT 616.950 733.950 619.050 734.400 ;
        RECT 625.950 733.950 628.050 734.400 ;
        RECT 658.950 735.450 661.050 736.050 ;
        RECT 664.950 735.450 667.050 736.050 ;
        RECT 658.950 734.400 667.050 735.450 ;
        RECT 658.950 733.950 661.050 734.400 ;
        RECT 664.950 733.950 667.050 734.400 ;
        RECT 670.950 735.450 673.050 736.050 ;
        RECT 691.950 735.450 694.050 736.050 ;
        RECT 670.950 734.400 694.050 735.450 ;
        RECT 670.950 733.950 673.050 734.400 ;
        RECT 691.950 733.950 694.050 734.400 ;
        RECT 28.950 732.450 31.050 733.050 ;
        RECT 46.950 732.450 49.050 733.050 ;
        RECT 106.950 732.450 109.050 733.050 ;
        RECT 28.950 731.400 109.050 732.450 ;
        RECT 28.950 730.950 31.050 731.400 ;
        RECT 46.950 730.950 49.050 731.400 ;
        RECT 106.950 730.950 109.050 731.400 ;
        RECT 151.950 732.450 154.050 733.050 ;
        RECT 172.950 732.450 175.050 733.050 ;
        RECT 151.950 731.400 175.050 732.450 ;
        RECT 151.950 730.950 154.050 731.400 ;
        RECT 172.950 730.950 175.050 731.400 ;
        RECT 223.950 732.450 226.050 733.050 ;
        RECT 334.950 732.450 337.050 733.050 ;
        RECT 454.950 732.450 457.050 733.050 ;
        RECT 223.950 731.400 457.050 732.450 ;
        RECT 223.950 730.950 226.050 731.400 ;
        RECT 334.950 730.950 337.050 731.400 ;
        RECT 454.950 730.950 457.050 731.400 ;
        RECT 562.950 732.450 565.050 733.050 ;
        RECT 622.950 732.450 625.050 733.050 ;
        RECT 562.950 731.400 625.050 732.450 ;
        RECT 562.950 730.950 565.050 731.400 ;
        RECT 622.950 730.950 625.050 731.400 ;
        RECT 637.950 732.450 640.050 733.050 ;
        RECT 682.950 732.450 685.050 733.050 ;
        RECT 704.400 732.450 705.450 736.950 ;
        RECT 712.950 735.300 715.050 737.400 ;
        RECT 637.950 731.400 705.450 732.450 ;
        RECT 713.850 731.700 715.050 735.300 ;
        RECT 734.100 732.600 735.300 749.400 ;
        RECT 752.400 744.000 771.450 744.450 ;
        RECT 751.950 743.400 772.050 744.000 ;
        RECT 751.950 739.950 754.050 743.400 ;
        RECT 769.950 739.950 772.050 743.400 ;
        RECT 772.950 742.950 775.050 748.050 ;
        RECT 832.950 747.450 835.050 748.050 ;
        RECT 827.400 747.000 835.050 747.450 ;
        RECT 826.950 746.400 835.050 747.000 ;
        RECT 778.950 742.050 781.050 745.050 ;
        RECT 796.950 742.950 802.050 745.050 ;
        RECT 808.950 742.950 814.050 745.050 ;
        RECT 826.950 742.950 829.050 746.400 ;
        RECT 832.950 745.950 835.050 746.400 ;
        RECT 830.400 744.000 846.450 744.450 ;
        RECT 829.950 743.400 847.050 744.000 ;
        RECT 775.800 741.000 777.900 742.050 ;
        RECT 778.950 741.450 781.200 742.050 ;
        RECT 790.950 741.450 793.050 742.050 ;
        RECT 778.950 741.000 793.050 741.450 ;
        RECT 824.100 741.000 826.200 742.050 ;
        RECT 775.800 739.950 778.050 741.000 ;
        RECT 779.100 740.400 793.050 741.000 ;
        RECT 779.100 739.950 781.200 740.400 ;
        RECT 790.950 739.950 793.050 740.400 ;
        RECT 823.950 739.950 826.200 741.000 ;
        RECT 829.950 739.950 832.050 743.400 ;
        RECT 844.950 739.950 847.050 743.400 ;
        RECT 742.950 738.450 745.050 739.050 ;
        RECT 748.950 738.450 751.050 739.050 ;
        RECT 742.950 737.400 751.050 738.450 ;
        RECT 742.950 736.950 745.050 737.400 ;
        RECT 748.950 736.950 751.050 737.400 ;
        RECT 754.950 738.450 757.050 739.050 ;
        RECT 775.950 738.450 778.050 739.950 ;
        RECT 823.950 739.050 826.050 739.950 ;
        RECT 808.950 738.450 811.050 739.050 ;
        RECT 754.950 737.400 811.050 738.450 ;
        RECT 823.950 738.000 826.200 739.050 ;
        RECT 754.950 736.950 757.050 737.400 ;
        RECT 808.950 736.950 811.050 737.400 ;
        RECT 824.100 736.950 826.200 738.000 ;
        RECT 838.950 736.950 844.050 739.050 ;
        RECT 757.950 733.050 760.050 736.050 ;
        RECT 823.950 735.450 826.050 736.050 ;
        RECT 841.950 735.450 844.050 736.050 ;
        RECT 847.950 735.450 850.050 739.050 ;
        RECT 823.950 735.000 850.050 735.450 ;
        RECT 823.950 734.400 849.450 735.000 ;
        RECT 823.950 733.950 826.050 734.400 ;
        RECT 841.950 733.950 844.050 734.400 ;
        RECT 637.950 730.950 640.050 731.400 ;
        RECT 682.950 730.950 685.050 731.400 ;
        RECT 22.950 729.450 25.050 730.050 ;
        RECT 8.400 728.400 25.050 729.450 ;
        RECT 8.400 724.050 9.450 728.400 ;
        RECT 22.950 727.950 25.050 728.400 ;
        RECT 58.950 729.450 61.050 730.050 ;
        RECT 64.950 729.450 70.050 730.050 ;
        RECT 58.950 728.400 70.050 729.450 ;
        RECT 58.950 727.950 61.050 728.400 ;
        RECT 64.950 727.950 70.050 728.400 ;
        RECT 85.950 729.450 88.050 730.050 ;
        RECT 103.950 729.450 106.050 730.050 ;
        RECT 85.950 728.400 106.050 729.450 ;
        RECT 85.950 727.950 88.050 728.400 ;
        RECT 103.950 727.950 106.050 728.400 ;
        RECT 325.950 729.450 328.050 730.050 ;
        RECT 370.950 729.450 373.050 730.050 ;
        RECT 418.950 729.450 421.050 730.050 ;
        RECT 325.950 728.400 421.050 729.450 ;
        RECT 325.950 727.950 328.050 728.400 ;
        RECT 370.950 727.950 373.050 728.400 ;
        RECT 418.950 727.950 421.050 728.400 ;
        RECT 430.950 729.450 433.050 730.050 ;
        RECT 448.950 729.450 451.050 730.050 ;
        RECT 472.950 729.450 475.050 730.050 ;
        RECT 430.950 728.400 475.050 729.450 ;
        RECT 430.950 727.950 433.050 728.400 ;
        RECT 448.950 727.950 451.050 728.400 ;
        RECT 472.950 727.950 475.050 728.400 ;
        RECT 601.950 727.950 606.900 730.050 ;
        RECT 608.100 729.450 610.200 730.050 ;
        RECT 670.950 729.450 673.050 730.050 ;
        RECT 712.950 729.600 715.050 731.700 ;
        RECT 733.950 730.500 736.050 732.600 ;
        RECT 754.950 732.000 760.050 733.050 ;
        RECT 763.950 732.450 766.050 733.050 ;
        RECT 838.950 732.450 841.050 733.050 ;
        RECT 844.950 732.450 847.050 733.050 ;
        RECT 754.950 731.400 759.450 732.000 ;
        RECT 763.950 731.400 847.050 732.450 ;
        RECT 754.950 730.950 759.000 731.400 ;
        RECT 763.950 730.950 766.050 731.400 ;
        RECT 838.950 730.950 841.050 731.400 ;
        RECT 844.950 730.950 847.050 731.400 ;
        RECT 608.100 728.400 673.050 729.450 ;
        RECT 608.100 727.950 610.200 728.400 ;
        RECT 670.950 727.950 673.050 728.400 ;
        RECT 769.950 729.450 772.050 730.050 ;
        RECT 805.950 729.450 808.050 730.200 ;
        RECT 769.950 728.400 808.050 729.450 ;
        RECT 769.950 727.950 772.050 728.400 ;
        RECT 805.950 728.100 808.050 728.400 ;
        RECT 10.950 726.450 13.050 727.050 ;
        RECT 22.950 726.450 25.050 727.050 ;
        RECT 79.950 726.450 82.050 727.050 ;
        RECT 100.950 726.450 103.050 727.050 ;
        RECT 259.950 726.450 262.050 727.050 ;
        RECT 10.950 725.400 262.050 726.450 ;
        RECT 10.950 724.950 13.050 725.400 ;
        RECT 22.950 724.950 25.050 725.400 ;
        RECT 79.950 724.950 82.050 725.400 ;
        RECT 100.950 724.950 103.050 725.400 ;
        RECT 259.950 724.950 262.050 725.400 ;
        RECT 373.950 726.450 376.050 727.050 ;
        RECT 424.950 726.450 427.050 727.050 ;
        RECT 373.950 725.400 427.050 726.450 ;
        RECT 373.950 724.950 376.050 725.400 ;
        RECT 424.950 724.950 427.050 725.400 ;
        RECT 430.950 726.450 433.050 727.050 ;
        RECT 442.950 726.450 445.050 727.050 ;
        RECT 430.950 725.400 445.050 726.450 ;
        RECT 430.950 724.950 433.050 725.400 ;
        RECT 442.950 724.950 445.050 725.400 ;
        RECT 481.950 726.450 484.050 727.050 ;
        RECT 523.950 726.450 526.050 727.050 ;
        RECT 481.950 725.400 526.050 726.450 ;
        RECT 481.950 724.950 484.050 725.400 ;
        RECT 523.950 724.950 526.050 725.400 ;
        RECT 616.950 726.450 619.050 727.050 ;
        RECT 673.950 726.450 676.050 727.050 ;
        RECT 616.950 725.400 676.050 726.450 ;
        RECT 616.950 724.950 619.050 725.400 ;
        RECT 673.950 724.950 676.050 725.400 ;
        RECT 709.950 726.450 712.050 727.050 ;
        RECT 742.950 726.450 745.050 727.050 ;
        RECT 709.950 725.400 745.050 726.450 ;
        RECT 709.950 724.950 712.050 725.400 ;
        RECT 742.950 724.950 745.050 725.400 ;
        RECT 805.950 726.450 808.050 726.900 ;
        RECT 814.950 726.450 817.050 727.050 ;
        RECT 820.950 726.450 823.050 727.050 ;
        RECT 805.950 725.400 823.050 726.450 ;
        RECT 7.950 721.950 10.050 724.050 ;
        RECT 70.950 723.450 73.050 724.050 ;
        RECT 91.950 723.450 94.050 724.050 ;
        RECT 103.950 723.450 106.050 724.050 ;
        RECT 70.950 722.400 106.050 723.450 ;
        RECT 70.950 721.950 73.050 722.400 ;
        RECT 91.950 721.950 94.050 722.400 ;
        RECT 103.950 721.950 106.050 722.400 ;
        RECT 205.950 723.450 208.050 724.050 ;
        RECT 235.950 723.450 238.050 724.050 ;
        RECT 374.400 723.450 375.450 724.950 ;
        RECT 805.950 724.800 808.050 725.400 ;
        RECT 814.950 724.950 817.050 725.400 ;
        RECT 820.950 724.950 823.050 725.400 ;
        RECT 205.950 722.400 375.450 723.450 ;
        RECT 439.950 723.450 442.050 724.050 ;
        RECT 544.950 723.450 547.050 724.050 ;
        RECT 592.950 723.450 595.050 724.050 ;
        RECT 439.950 722.400 595.050 723.450 ;
        RECT 205.950 721.950 208.050 722.400 ;
        RECT 235.950 721.950 238.050 722.400 ;
        RECT 439.950 721.950 442.050 722.400 ;
        RECT 544.950 721.950 547.050 722.400 ;
        RECT 592.950 721.950 595.050 722.400 ;
        RECT 598.950 723.450 601.050 724.050 ;
        RECT 649.950 723.450 652.050 724.050 ;
        RECT 598.950 722.400 652.050 723.450 ;
        RECT 598.950 721.950 601.050 722.400 ;
        RECT 649.950 721.950 652.050 722.400 ;
        RECT 670.950 723.450 673.050 724.050 ;
        RECT 697.950 723.450 700.050 724.050 ;
        RECT 826.950 723.450 829.050 724.050 ;
        RECT 670.950 722.400 700.050 723.450 ;
        RECT 670.950 721.950 673.050 722.400 ;
        RECT 697.950 721.950 700.050 722.400 ;
        RECT 704.400 722.400 829.050 723.450 ;
        RECT 292.950 720.450 295.050 721.050 ;
        RECT 328.950 720.450 331.050 721.050 ;
        RECT 292.950 719.400 331.050 720.450 ;
        RECT 292.950 718.950 295.050 719.400 ;
        RECT 328.950 718.950 331.050 719.400 ;
        RECT 412.950 720.450 415.050 721.050 ;
        RECT 436.950 720.450 439.050 721.050 ;
        RECT 457.950 720.450 460.050 721.050 ;
        RECT 484.950 720.450 487.050 721.050 ;
        RECT 412.950 720.000 420.600 720.450 ;
        RECT 412.950 719.400 421.050 720.000 ;
        RECT 412.950 718.950 415.050 719.400 ;
        RECT 418.950 718.050 421.050 719.400 ;
        RECT 436.950 719.400 487.050 720.450 ;
        RECT 436.950 718.950 439.050 719.400 ;
        RECT 457.950 718.950 460.050 719.400 ;
        RECT 484.950 718.950 487.050 719.400 ;
        RECT 508.950 720.450 511.050 721.050 ;
        RECT 535.950 720.450 538.050 721.050 ;
        RECT 508.950 719.400 538.050 720.450 ;
        RECT 508.950 718.950 511.050 719.400 ;
        RECT 535.950 718.950 538.050 719.400 ;
        RECT 541.950 720.450 544.050 721.050 ;
        RECT 553.950 720.450 556.050 721.050 ;
        RECT 541.950 719.400 556.050 720.450 ;
        RECT 541.950 718.950 544.050 719.400 ;
        RECT 553.950 718.950 556.050 719.400 ;
        RECT 610.950 720.450 613.050 721.050 ;
        RECT 643.950 720.450 646.050 721.050 ;
        RECT 610.950 719.400 646.050 720.450 ;
        RECT 610.950 718.950 613.050 719.400 ;
        RECT 643.950 718.950 646.050 719.400 ;
        RECT 673.950 720.450 676.050 721.050 ;
        RECT 704.400 720.450 705.450 722.400 ;
        RECT 826.950 721.950 829.050 722.400 ;
        RECT 730.950 720.450 733.050 721.050 ;
        RECT 673.950 719.400 705.450 720.450 ;
        RECT 707.400 719.400 733.050 720.450 ;
        RECT 673.950 718.950 676.050 719.400 ;
        RECT 97.950 717.450 100.050 718.050 ;
        RECT 217.950 717.450 220.050 718.050 ;
        RECT 97.950 716.400 220.050 717.450 ;
        RECT 97.950 715.950 100.050 716.400 ;
        RECT 217.950 715.950 220.050 716.400 ;
        RECT 388.950 717.450 391.050 718.050 ;
        RECT 397.950 717.450 400.050 718.050 ;
        RECT 388.950 716.400 400.050 717.450 ;
        RECT 388.950 715.950 391.050 716.400 ;
        RECT 397.950 715.950 400.050 716.400 ;
        RECT 403.950 717.450 406.050 718.050 ;
        RECT 415.800 717.450 417.900 718.050 ;
        RECT 403.950 716.400 417.900 717.450 ;
        RECT 418.950 717.000 421.200 718.050 ;
        RECT 403.950 715.950 406.050 716.400 ;
        RECT 415.800 715.950 417.900 716.400 ;
        RECT 419.100 715.950 421.200 717.000 ;
        RECT 424.950 717.450 427.050 718.050 ;
        RECT 481.950 717.450 484.050 718.050 ;
        RECT 424.950 716.400 484.050 717.450 ;
        RECT 424.950 715.950 427.050 716.400 ;
        RECT 481.950 715.950 484.050 716.400 ;
        RECT 568.950 717.450 571.050 718.050 ;
        RECT 613.950 717.450 616.050 718.050 ;
        RECT 568.950 716.400 616.050 717.450 ;
        RECT 568.950 715.950 571.050 716.400 ;
        RECT 613.950 715.950 616.050 716.400 ;
        RECT 622.950 717.450 625.050 718.050 ;
        RECT 640.950 717.450 643.050 718.050 ;
        RECT 622.950 716.400 643.050 717.450 ;
        RECT 622.950 715.950 625.050 716.400 ;
        RECT 640.950 715.950 643.050 716.400 ;
        RECT 685.950 717.450 688.050 718.050 ;
        RECT 707.400 717.450 708.450 719.400 ;
        RECT 730.950 718.950 733.050 719.400 ;
        RECT 685.950 716.400 708.450 717.450 ;
        RECT 709.950 717.450 712.050 718.050 ;
        RECT 754.950 717.450 757.050 718.050 ;
        RECT 709.950 716.400 757.050 717.450 ;
        RECT 685.950 715.950 688.050 716.400 ;
        RECT 709.950 715.950 712.050 716.400 ;
        RECT 754.950 715.950 757.050 716.400 ;
        RECT 52.950 714.450 55.050 715.050 ;
        RECT 91.950 714.450 94.050 715.050 ;
        RECT 112.950 714.450 115.050 715.050 ;
        RECT 124.950 714.450 127.050 715.050 ;
        RECT 52.950 713.400 127.050 714.450 ;
        RECT 52.950 712.950 55.050 713.400 ;
        RECT 91.950 712.950 94.050 713.400 ;
        RECT 112.950 712.950 115.050 713.400 ;
        RECT 124.950 712.950 127.050 713.400 ;
        RECT 400.950 714.450 403.050 715.050 ;
        RECT 601.950 714.450 604.050 715.050 ;
        RECT 400.950 713.400 604.050 714.450 ;
        RECT 400.950 712.950 403.050 713.400 ;
        RECT 601.950 712.950 604.050 713.400 ;
        RECT 58.950 711.450 61.050 712.050 ;
        RECT 118.950 711.450 121.050 712.050 ;
        RECT 139.950 711.450 142.050 712.050 ;
        RECT 58.950 710.400 142.050 711.450 ;
        RECT 58.950 709.950 61.050 710.400 ;
        RECT 118.950 709.950 121.050 710.400 ;
        RECT 139.950 709.950 142.050 710.400 ;
        RECT 178.950 711.450 181.050 712.050 ;
        RECT 193.950 711.450 196.050 712.050 ;
        RECT 178.950 710.400 196.050 711.450 ;
        RECT 178.950 709.950 181.050 710.400 ;
        RECT 193.950 709.950 196.050 710.400 ;
        RECT 238.950 711.450 241.050 712.050 ;
        RECT 292.950 711.450 295.050 712.050 ;
        RECT 238.950 710.400 295.050 711.450 ;
        RECT 238.950 709.950 241.050 710.400 ;
        RECT 292.950 709.950 295.050 710.400 ;
        RECT 322.950 711.450 325.050 712.050 ;
        RECT 367.950 711.450 370.050 712.050 ;
        RECT 322.950 710.400 370.050 711.450 ;
        RECT 322.950 709.950 325.050 710.400 ;
        RECT 367.950 709.950 370.050 710.400 ;
        RECT 391.950 711.450 394.050 712.050 ;
        RECT 439.950 711.450 442.050 712.050 ;
        RECT 391.950 710.400 442.050 711.450 ;
        RECT 391.950 709.950 394.050 710.400 ;
        RECT 439.950 709.950 442.050 710.400 ;
        RECT 517.950 711.450 520.050 712.050 ;
        RECT 559.950 711.450 562.050 712.050 ;
        RECT 517.950 710.400 562.050 711.450 ;
        RECT 517.950 709.950 520.050 710.400 ;
        RECT 559.950 709.950 562.050 710.400 ;
        RECT 592.950 711.450 595.050 712.050 ;
        RECT 607.950 711.450 610.050 712.050 ;
        RECT 592.950 710.400 630.450 711.450 ;
        RECT 640.950 710.400 643.050 712.500 ;
        RECT 661.950 711.300 664.050 713.400 ;
        RECT 709.950 711.300 712.050 713.400 ;
        RECT 592.950 709.950 595.050 710.400 ;
        RECT 607.950 709.950 610.050 710.400 ;
        RECT 16.950 703.950 19.050 709.050 ;
        RECT 95.100 708.000 97.200 709.050 ;
        RECT 331.950 708.450 334.050 709.050 ;
        RECT 94.950 706.950 97.200 708.000 ;
        RECT 245.400 707.400 273.450 708.450 ;
        RECT 287.400 708.000 334.050 708.450 ;
        RECT 94.950 706.050 97.050 706.950 ;
        RECT 245.400 706.050 246.450 707.400 ;
        RECT 49.950 705.450 52.050 706.050 ;
        RECT 49.950 705.000 75.450 705.450 ;
        RECT 91.800 705.000 93.900 706.050 ;
        RECT 94.950 705.450 97.200 706.050 ;
        RECT 94.950 705.000 111.450 705.450 ;
        RECT 49.950 704.400 76.050 705.000 ;
        RECT 49.950 703.950 52.050 704.400 ;
        RECT 7.950 702.450 10.050 703.050 ;
        RECT 13.950 702.450 16.050 703.050 ;
        RECT 7.950 701.400 16.050 702.450 ;
        RECT 7.950 700.950 10.050 701.400 ;
        RECT 13.950 697.950 16.050 701.400 ;
        RECT 19.950 700.950 25.050 703.050 ;
        RECT 28.800 700.950 30.900 703.050 ;
        RECT 32.100 700.950 37.050 703.050 ;
        RECT 52.950 700.950 57.900 703.050 ;
        RECT 59.100 700.950 64.050 703.050 ;
        RECT 73.950 700.950 76.050 704.400 ;
        RECT 91.800 703.950 94.050 705.000 ;
        RECT 95.100 704.400 111.450 705.000 ;
        RECT 95.100 703.950 97.200 704.400 ;
        RECT 79.950 700.950 85.050 703.050 ;
        RECT 91.950 700.950 94.050 703.950 ;
        RECT 110.400 703.050 111.450 704.400 ;
        RECT 112.950 703.950 118.050 706.050 ;
        RECT 148.950 705.450 151.050 706.050 ;
        RECT 148.950 705.000 159.450 705.450 ;
        RECT 148.950 704.400 160.050 705.000 ;
        RECT 148.950 703.950 151.050 704.400 ;
        RECT 4.950 696.450 7.050 697.050 ;
        RECT 29.250 696.450 30.300 700.950 ;
        RECT 31.950 697.950 34.050 700.050 ;
        RECT 40.950 699.450 43.050 700.050 ;
        RECT 49.950 699.450 52.050 700.050 ;
        RECT 40.950 698.400 52.050 699.450 ;
        RECT 40.950 697.950 43.050 698.400 ;
        RECT 49.950 697.950 52.050 698.400 ;
        RECT 4.950 695.400 30.300 696.450 ;
        RECT 4.950 694.950 7.050 695.400 ;
        RECT 10.950 693.450 13.050 694.050 ;
        RECT 32.400 693.450 33.450 697.950 ;
        RECT 55.950 694.950 58.050 700.050 ;
        RECT 67.950 697.950 73.050 700.050 ;
        RECT 76.950 694.950 79.050 700.050 ;
        RECT 97.950 697.950 100.050 703.050 ;
        RECT 110.400 702.450 115.050 703.050 ;
        RECT 110.400 701.400 117.450 702.450 ;
        RECT 111.000 700.950 115.050 701.400 ;
        RECT 116.400 699.450 117.450 701.400 ;
        RECT 118.950 700.950 123.900 703.050 ;
        RECT 125.100 702.450 127.200 703.050 ;
        RECT 133.950 702.450 136.050 703.050 ;
        RECT 125.100 701.400 136.050 702.450 ;
        RECT 125.100 700.950 127.200 701.400 ;
        RECT 133.950 700.950 136.050 701.400 ;
        RECT 139.950 700.950 145.050 703.050 ;
        RECT 157.950 700.950 160.050 704.400 ;
        RECT 175.950 703.950 181.050 706.050 ;
        RECT 184.950 705.450 190.050 706.050 ;
        RECT 196.950 705.450 199.050 706.050 ;
        RECT 184.950 704.400 199.050 705.450 ;
        RECT 184.950 703.950 190.050 704.400 ;
        RECT 196.950 703.950 199.050 704.400 ;
        RECT 217.950 705.450 220.050 706.050 ;
        RECT 232.950 705.450 235.050 706.050 ;
        RECT 217.950 704.400 235.050 705.450 ;
        RECT 217.950 703.950 220.050 704.400 ;
        RECT 232.950 703.950 235.050 704.400 ;
        RECT 238.800 705.000 240.900 706.050 ;
        RECT 238.800 703.950 241.050 705.000 ;
        RECT 242.100 704.400 246.450 706.050 ;
        RECT 268.950 705.450 271.050 706.050 ;
        RECT 263.400 705.000 271.050 705.450 ;
        RECT 262.950 704.400 271.050 705.000 ;
        RECT 272.400 705.450 273.450 707.400 ;
        RECT 286.950 707.400 334.050 708.000 ;
        RECT 277.950 705.450 280.050 706.050 ;
        RECT 272.400 704.400 280.050 705.450 ;
        RECT 242.100 703.950 246.000 704.400 ;
        RECT 163.950 700.950 169.050 703.050 ;
        RECT 180.000 702.900 184.050 703.050 ;
        RECT 178.950 700.950 184.050 702.900 ;
        RECT 190.950 700.950 196.050 703.050 ;
        RECT 178.950 700.800 181.050 700.950 ;
        RECT 136.800 699.450 138.900 700.050 ;
        RECT 116.400 698.400 138.900 699.450 ;
        RECT 136.800 697.950 138.900 698.400 ;
        RECT 140.100 699.450 142.200 699.900 ;
        RECT 154.950 699.450 157.050 700.050 ;
        RECT 140.100 698.400 157.050 699.450 ;
        RECT 140.100 697.800 142.200 698.400 ;
        RECT 154.950 697.950 157.050 698.400 ;
        RECT 160.950 696.450 163.050 700.050 ;
        RECT 199.950 697.950 202.050 703.050 ;
        RECT 221.400 701.400 228.450 702.450 ;
        RECT 208.950 699.450 211.050 700.050 ;
        RECT 217.950 699.450 220.050 700.050 ;
        RECT 221.400 699.450 222.450 701.400 ;
        RECT 208.950 698.400 222.450 699.450 ;
        RECT 208.950 697.950 211.050 698.400 ;
        RECT 217.950 697.950 220.050 698.400 ;
        RECT 223.950 697.050 226.050 700.050 ;
        RECT 227.400 699.450 228.450 701.400 ;
        RECT 238.950 700.950 241.050 703.950 ;
        RECT 244.950 700.950 250.050 703.050 ;
        RECT 256.950 700.050 259.050 703.050 ;
        RECT 262.950 700.950 265.050 704.400 ;
        RECT 268.950 703.950 271.050 704.400 ;
        RECT 277.950 703.950 280.050 704.400 ;
        RECT 286.950 703.950 289.050 707.400 ;
        RECT 301.950 706.050 304.050 707.400 ;
        RECT 331.950 706.950 334.050 707.400 ;
        RECT 430.950 708.450 433.050 709.050 ;
        RECT 451.950 708.450 454.050 709.050 ;
        RECT 430.950 707.400 454.050 708.450 ;
        RECT 430.950 706.950 433.050 707.400 ;
        RECT 451.950 706.950 454.050 707.400 ;
        RECT 478.950 708.450 481.050 709.050 ;
        RECT 487.950 708.450 490.050 709.050 ;
        RECT 478.950 707.400 490.050 708.450 ;
        RECT 478.950 706.950 481.050 707.400 ;
        RECT 487.950 706.950 490.050 707.400 ;
        RECT 493.950 706.050 496.050 709.050 ;
        RECT 505.950 708.450 508.050 709.050 ;
        RECT 565.950 708.450 568.050 709.050 ;
        RECT 589.950 708.450 592.050 709.050 ;
        RECT 505.950 707.400 568.050 708.450 ;
        RECT 578.400 708.000 592.050 708.450 ;
        RECT 505.950 706.950 508.050 707.400 ;
        RECT 565.950 706.950 568.050 707.400 ;
        RECT 577.950 707.400 592.050 708.000 ;
        RECT 301.800 705.000 304.050 706.050 ;
        RECT 305.100 705.000 307.200 706.050 ;
        RECT 385.950 705.450 388.050 706.050 ;
        RECT 301.800 703.950 303.900 705.000 ;
        RECT 304.950 703.950 307.200 705.000 ;
        RECT 380.400 704.400 388.050 705.450 ;
        RECT 283.950 700.950 288.900 703.050 ;
        RECT 290.100 702.450 292.200 703.050 ;
        RECT 304.950 702.450 307.050 703.950 ;
        RECT 380.400 703.050 381.450 704.400 ;
        RECT 385.950 703.950 388.050 704.400 ;
        RECT 391.950 703.050 394.050 706.050 ;
        RECT 430.950 705.450 433.050 706.050 ;
        RECT 413.400 704.400 433.050 705.450 ;
        RECT 290.100 701.400 307.050 702.450 ;
        RECT 290.100 700.950 292.200 701.400 ;
        RECT 304.950 700.950 307.050 701.400 ;
        RECT 310.950 700.050 313.050 703.050 ;
        RECT 316.950 700.950 322.050 703.050 ;
        RECT 352.950 700.050 355.050 703.050 ;
        RECT 358.950 700.950 364.050 703.050 ;
        RECT 376.950 700.950 382.050 703.050 ;
        RECT 388.800 702.000 390.900 703.050 ;
        RECT 391.950 702.000 394.200 703.050 ;
        RECT 388.800 700.950 391.050 702.000 ;
        RECT 392.100 700.950 394.200 702.000 ;
        RECT 397.950 702.450 400.050 703.050 ;
        RECT 406.950 702.450 412.050 703.050 ;
        RECT 397.950 701.400 412.050 702.450 ;
        RECT 397.950 700.950 400.050 701.400 ;
        RECT 406.950 700.950 412.050 701.400 ;
        RECT 253.800 699.450 255.900 700.050 ;
        RECT 227.400 698.400 255.900 699.450 ;
        RECT 253.800 697.950 255.900 698.400 ;
        RECT 256.800 699.000 259.050 700.050 ;
        RECT 256.800 697.950 258.900 699.000 ;
        RECT 260.100 697.950 264.900 700.050 ;
        RECT 266.100 699.450 268.200 700.050 ;
        RECT 298.800 699.450 300.900 700.050 ;
        RECT 266.100 698.400 300.900 699.450 ;
        RECT 266.100 697.950 268.200 698.400 ;
        RECT 298.800 697.950 300.900 698.400 ;
        RECT 302.100 699.450 304.200 700.050 ;
        RECT 307.800 699.450 309.900 700.050 ;
        RECT 302.100 698.400 309.900 699.450 ;
        RECT 310.950 699.000 313.200 700.050 ;
        RECT 349.800 699.450 351.900 700.050 ;
        RECT 302.100 697.950 304.200 698.400 ;
        RECT 307.800 697.950 309.900 698.400 ;
        RECT 311.100 697.950 313.200 699.000 ;
        RECT 332.400 698.400 351.900 699.450 ;
        RECT 199.950 696.450 202.050 697.050 ;
        RECT 160.950 696.000 202.050 696.450 ;
        RECT 161.400 695.400 202.050 696.000 ;
        RECT 199.950 694.950 202.050 695.400 ;
        RECT 220.800 696.000 222.900 697.050 ;
        RECT 223.950 696.450 226.200 697.050 ;
        RECT 256.950 696.450 259.050 697.050 ;
        RECT 223.950 696.000 259.050 696.450 ;
        RECT 220.800 694.950 223.050 696.000 ;
        RECT 224.100 695.400 259.050 696.000 ;
        RECT 224.100 694.950 226.200 695.400 ;
        RECT 256.950 694.950 259.050 695.400 ;
        RECT 277.950 696.450 280.050 697.050 ;
        RECT 316.950 696.450 322.050 697.050 ;
        RECT 332.400 696.450 333.450 698.400 ;
        RECT 349.800 697.950 351.900 698.400 ;
        RECT 352.800 699.000 355.050 700.050 ;
        RECT 352.800 697.950 354.900 699.000 ;
        RECT 356.100 697.950 361.050 700.050 ;
        RECT 364.950 699.450 367.050 700.050 ;
        RECT 373.950 699.450 376.050 700.050 ;
        RECT 388.950 699.450 391.050 700.950 ;
        RECT 413.400 700.050 414.450 704.400 ;
        RECT 430.950 703.950 433.050 704.400 ;
        RECT 436.950 705.450 439.050 706.050 ;
        RECT 445.950 705.450 448.050 706.050 ;
        RECT 436.950 704.400 448.050 705.450 ;
        RECT 436.950 703.950 439.050 704.400 ;
        RECT 445.950 703.950 448.050 704.400 ;
        RECT 466.950 705.450 469.050 706.050 ;
        RECT 475.950 705.450 478.050 706.050 ;
        RECT 466.950 704.400 478.050 705.450 ;
        RECT 466.950 703.950 469.050 704.400 ;
        RECT 475.950 703.950 478.050 704.400 ;
        RECT 481.950 703.950 487.050 706.050 ;
        RECT 493.800 705.000 496.050 706.050 ;
        RECT 497.100 705.450 499.200 706.050 ;
        RECT 502.950 705.450 505.050 706.050 ;
        RECT 493.800 703.950 495.900 705.000 ;
        RECT 497.100 704.400 505.050 705.450 ;
        RECT 497.100 703.950 499.200 704.400 ;
        RECT 502.950 703.950 505.050 704.400 ;
        RECT 508.950 703.950 514.050 706.050 ;
        RECT 565.950 705.450 568.050 706.050 ;
        RECT 571.950 705.450 574.050 706.050 ;
        RECT 565.950 704.400 574.050 705.450 ;
        RECT 565.950 703.950 568.050 704.400 ;
        RECT 571.950 703.950 574.050 704.400 ;
        RECT 577.950 703.950 580.050 707.400 ;
        RECT 589.950 706.950 592.050 707.400 ;
        RECT 629.400 706.050 630.450 710.400 ;
        RECT 619.950 703.950 625.050 706.050 ;
        RECT 628.950 703.950 631.050 706.050 ;
        RECT 418.950 703.050 421.050 703.200 ;
        RECT 415.950 701.100 421.050 703.050 ;
        RECT 415.950 700.950 420.000 701.100 ;
        RECT 433.950 700.950 439.050 703.050 ;
        RECT 457.950 702.450 460.050 703.050 ;
        RECT 463.950 702.450 466.050 703.050 ;
        RECT 457.950 701.400 466.050 702.450 ;
        RECT 457.950 700.950 460.050 701.400 ;
        RECT 463.950 700.950 466.050 701.400 ;
        RECT 472.950 702.450 475.050 703.050 ;
        RECT 481.950 702.450 484.050 703.050 ;
        RECT 472.950 701.400 484.050 702.450 ;
        RECT 472.950 700.950 475.050 701.400 ;
        RECT 481.950 700.950 484.050 701.400 ;
        RECT 397.950 699.450 400.050 700.050 ;
        RECT 406.950 699.450 409.050 700.050 ;
        RECT 364.950 698.400 387.450 699.450 ;
        RECT 388.950 699.000 409.050 699.450 ;
        RECT 389.400 698.400 409.050 699.000 ;
        RECT 364.950 697.950 367.050 698.400 ;
        RECT 373.950 697.950 376.050 698.400 ;
        RECT 277.950 695.400 333.450 696.450 ;
        RECT 334.950 696.450 337.050 697.050 ;
        RECT 353.400 696.450 354.450 697.950 ;
        RECT 334.950 695.400 354.450 696.450 ;
        RECT 386.400 696.450 387.450 698.400 ;
        RECT 397.950 697.950 400.050 698.400 ;
        RECT 406.950 697.950 409.050 698.400 ;
        RECT 412.800 697.950 414.900 700.050 ;
        RECT 418.950 697.950 424.050 700.050 ;
        RECT 445.950 697.950 451.050 700.050 ;
        RECT 464.400 699.450 465.450 700.950 ;
        RECT 487.950 699.450 490.050 703.050 ;
        RECT 505.950 702.450 508.050 703.050 ;
        RECT 514.950 702.450 517.050 703.050 ;
        RECT 505.950 701.400 517.050 702.450 ;
        RECT 505.950 700.950 508.050 701.400 ;
        RECT 514.950 700.950 517.050 701.400 ;
        RECT 523.950 700.950 529.050 703.050 ;
        RECT 538.950 702.450 544.050 703.050 ;
        RECT 538.950 702.000 552.450 702.450 ;
        RECT 538.950 701.400 553.050 702.000 ;
        RECT 538.950 700.950 544.050 701.400 ;
        RECT 464.400 699.000 490.050 699.450 ;
        RECT 464.400 698.400 489.450 699.000 ;
        RECT 517.950 697.950 523.050 700.050 ;
        RECT 550.950 697.950 553.050 701.400 ;
        RECT 571.950 700.950 577.050 703.050 ;
        RECT 594.000 702.450 598.050 703.050 ;
        RECT 613.950 702.450 616.050 703.050 ;
        RECT 625.950 702.450 628.050 703.050 ;
        RECT 593.550 702.000 598.050 702.450 ;
        RECT 611.400 702.000 628.050 702.450 ;
        RECT 592.950 700.950 598.050 702.000 ;
        RECT 610.950 701.400 628.050 702.000 ;
        RECT 592.950 700.050 595.050 700.950 ;
        RECT 556.950 697.950 562.050 700.050 ;
        RECT 565.950 699.450 568.050 700.050 ;
        RECT 586.800 699.450 588.900 700.050 ;
        RECT 565.950 698.400 588.900 699.450 ;
        RECT 565.950 697.950 568.050 698.400 ;
        RECT 586.800 697.950 588.900 698.400 ;
        RECT 589.800 699.000 591.900 700.050 ;
        RECT 592.950 699.000 595.200 700.050 ;
        RECT 589.800 697.950 592.050 699.000 ;
        RECT 593.100 697.950 595.200 699.000 ;
        RECT 598.950 699.450 601.050 700.050 ;
        RECT 604.950 699.450 607.050 700.050 ;
        RECT 598.950 698.400 607.050 699.450 ;
        RECT 598.950 697.950 601.050 698.400 ;
        RECT 604.950 697.950 607.050 698.400 ;
        RECT 610.950 697.950 613.050 701.400 ;
        RECT 613.950 700.950 616.050 701.400 ;
        RECT 625.950 700.950 628.050 701.400 ;
        RECT 625.950 699.450 628.050 700.050 ;
        RECT 634.950 699.450 637.050 700.050 ;
        RECT 625.950 698.400 637.050 699.450 ;
        RECT 625.950 697.950 628.050 698.400 ;
        RECT 634.950 697.950 637.050 698.400 ;
        RECT 589.950 697.050 592.050 697.950 ;
        RECT 436.950 696.450 439.050 697.050 ;
        RECT 386.400 695.400 439.050 696.450 ;
        RECT 277.950 694.950 280.050 695.400 ;
        RECT 316.950 694.950 322.050 695.400 ;
        RECT 334.950 694.950 337.050 695.400 ;
        RECT 436.950 694.950 439.050 695.400 ;
        RECT 445.950 696.450 448.050 697.050 ;
        RECT 451.950 696.450 454.050 697.050 ;
        RECT 445.950 695.400 454.050 696.450 ;
        RECT 445.950 694.950 448.050 695.400 ;
        RECT 451.950 694.950 454.050 695.400 ;
        RECT 469.950 694.950 475.050 697.050 ;
        RECT 481.950 696.450 484.050 697.050 ;
        RECT 511.950 696.450 514.050 697.050 ;
        RECT 481.950 695.400 514.050 696.450 ;
        RECT 481.950 694.950 484.050 695.400 ;
        RECT 511.950 694.950 514.050 695.400 ;
        RECT 532.950 694.950 538.050 697.050 ;
        RECT 553.950 696.450 556.050 697.050 ;
        RECT 565.950 696.450 568.050 697.050 ;
        RECT 539.400 695.400 568.050 696.450 ;
        RECT 10.950 692.400 33.450 693.450 ;
        RECT 49.950 693.450 52.050 694.050 ;
        RECT 61.950 693.450 64.050 694.050 ;
        RECT 49.950 692.400 64.050 693.450 ;
        RECT 10.950 691.950 13.050 692.400 ;
        RECT 49.950 691.950 52.050 692.400 ;
        RECT 61.950 691.950 64.050 692.400 ;
        RECT 82.950 693.450 85.050 694.050 ;
        RECT 97.950 693.450 100.050 694.050 ;
        RECT 82.950 692.400 100.050 693.450 ;
        RECT 220.950 693.450 223.050 694.950 ;
        RECT 244.950 693.450 247.050 694.050 ;
        RECT 220.950 693.000 247.050 693.450 ;
        RECT 221.400 692.400 247.050 693.000 ;
        RECT 82.950 691.950 85.050 692.400 ;
        RECT 97.950 691.950 100.050 692.400 ;
        RECT 244.950 691.950 247.050 692.400 ;
        RECT 262.950 693.450 265.050 694.050 ;
        RECT 403.950 693.450 406.050 694.050 ;
        RECT 262.950 692.400 406.050 693.450 ;
        RECT 262.950 691.950 265.050 692.400 ;
        RECT 403.950 691.950 406.050 692.400 ;
        RECT 514.950 693.450 517.050 694.050 ;
        RECT 539.400 693.450 540.450 695.400 ;
        RECT 553.950 694.950 556.050 695.400 ;
        RECT 565.950 694.950 568.050 695.400 ;
        RECT 589.800 696.000 592.050 697.050 ;
        RECT 589.800 694.950 591.900 696.000 ;
        RECT 604.950 694.950 610.050 697.050 ;
        RECT 514.950 692.400 540.450 693.450 ;
        RECT 547.950 693.450 550.050 694.050 ;
        RECT 568.950 693.450 571.050 694.050 ;
        RECT 641.700 693.600 642.900 710.400 ;
        RECT 661.950 707.700 663.150 711.300 ;
        RECT 710.850 707.700 712.050 711.300 ;
        RECT 730.950 710.400 733.050 712.500 ;
        RECT 817.950 710.400 820.050 712.500 ;
        RECT 838.950 711.300 841.050 713.400 ;
        RECT 661.950 705.600 664.050 707.700 ;
        RECT 646.950 697.950 649.050 703.050 ;
        RECT 652.950 694.950 655.050 700.050 ;
        RECT 661.950 693.600 663.150 705.600 ;
        RECT 673.950 703.950 679.050 706.050 ;
        RECT 682.950 703.950 688.050 706.050 ;
        RECT 709.950 705.600 712.050 707.700 ;
        RECT 679.950 700.950 685.050 703.050 ;
        RECT 694.950 700.950 700.050 703.050 ;
        RECT 664.950 697.950 670.050 700.050 ;
        RECT 703.950 697.950 709.050 700.050 ;
        RECT 547.950 692.400 571.050 693.450 ;
        RECT 514.950 691.950 517.050 692.400 ;
        RECT 547.950 691.950 550.050 692.400 ;
        RECT 568.950 691.950 571.050 692.400 ;
        RECT 640.950 691.500 643.050 693.600 ;
        RECT 661.950 691.500 664.050 693.600 ;
        RECT 673.950 693.450 676.050 694.050 ;
        RECT 703.950 693.450 706.050 694.050 ;
        RECT 710.850 693.600 712.050 705.600 ;
        RECT 718.950 694.950 721.050 700.050 ;
        RECT 724.950 697.950 727.050 703.050 ;
        RECT 731.100 693.600 732.300 710.400 ;
        RECT 742.950 703.950 748.050 706.050 ;
        RECT 751.950 705.450 754.050 706.050 ;
        RECT 760.950 705.450 763.050 706.050 ;
        RECT 751.950 704.400 771.450 705.450 ;
        RECT 751.950 703.950 754.050 704.400 ;
        RECT 760.950 703.950 763.050 704.400 ;
        RECT 748.950 702.450 751.050 703.050 ;
        RECT 766.950 702.450 769.050 703.050 ;
        RECT 748.950 701.400 769.050 702.450 ;
        RECT 770.400 702.450 771.450 704.400 ;
        RECT 772.950 702.450 775.050 703.050 ;
        RECT 770.400 701.400 783.450 702.450 ;
        RECT 748.950 700.950 751.050 701.400 ;
        RECT 766.950 700.950 769.050 701.400 ;
        RECT 772.950 700.950 775.050 701.400 ;
        RECT 782.400 700.050 783.450 701.400 ;
        RECT 805.950 700.950 811.050 703.050 ;
        RECT 733.950 699.450 736.050 700.050 ;
        RECT 769.950 699.450 772.050 700.050 ;
        RECT 733.950 698.400 772.050 699.450 ;
        RECT 733.950 697.950 736.050 698.400 ;
        RECT 769.950 697.950 772.050 698.400 ;
        RECT 775.950 697.950 781.050 700.050 ;
        RECT 782.400 698.400 787.050 700.050 ;
        RECT 783.000 697.950 787.050 698.400 ;
        RECT 790.950 697.950 796.050 700.050 ;
        RECT 763.950 696.450 766.050 697.050 ;
        RECT 787.950 696.450 790.050 697.050 ;
        RECT 763.950 695.400 790.050 696.450 ;
        RECT 763.950 694.950 766.050 695.400 ;
        RECT 787.950 694.950 790.050 695.400 ;
        RECT 673.950 692.400 706.050 693.450 ;
        RECT 673.950 691.950 676.050 692.400 ;
        RECT 703.950 691.950 706.050 692.400 ;
        RECT 709.950 691.500 712.050 693.600 ;
        RECT 730.950 691.500 733.050 693.600 ;
        RECT 775.950 693.450 778.050 694.050 ;
        RECT 796.950 693.450 799.050 694.050 ;
        RECT 818.700 693.600 819.900 710.400 ;
        RECT 838.950 707.700 840.150 711.300 ;
        RECT 838.950 705.600 841.050 707.700 ;
        RECT 832.950 702.450 835.050 703.050 ;
        RECT 824.250 702.000 835.050 702.450 ;
        RECT 823.950 701.400 835.050 702.000 ;
        RECT 823.950 700.050 826.050 701.400 ;
        RECT 832.950 700.950 835.050 701.400 ;
        RECT 823.800 699.000 826.050 700.050 ;
        RECT 823.800 697.950 825.900 699.000 ;
        RECT 827.100 697.950 832.050 700.050 ;
        RECT 838.950 693.600 840.150 705.600 ;
        RECT 841.950 697.950 847.050 700.050 ;
        RECT 775.950 692.400 799.050 693.450 ;
        RECT 775.950 691.950 778.050 692.400 ;
        RECT 796.950 691.950 799.050 692.400 ;
        RECT 817.950 691.500 820.050 693.600 ;
        RECT 838.950 691.500 841.050 693.600 ;
        RECT 91.950 690.450 94.050 691.050 ;
        RECT 106.950 690.450 109.050 691.050 ;
        RECT 112.950 690.450 115.050 691.050 ;
        RECT 91.950 689.400 115.050 690.450 ;
        RECT 91.950 688.950 94.050 689.400 ;
        RECT 106.950 688.950 109.050 689.400 ;
        RECT 112.950 688.950 115.050 689.400 ;
        RECT 127.950 690.450 130.050 691.050 ;
        RECT 145.950 690.450 148.050 691.050 ;
        RECT 163.950 690.450 166.050 691.050 ;
        RECT 184.950 690.450 187.050 691.050 ;
        RECT 127.950 689.400 187.050 690.450 ;
        RECT 127.950 688.950 130.050 689.400 ;
        RECT 145.950 688.950 148.050 689.400 ;
        RECT 163.950 688.950 166.050 689.400 ;
        RECT 184.950 688.950 187.050 689.400 ;
        RECT 208.950 690.450 211.050 691.050 ;
        RECT 247.950 690.450 250.050 691.050 ;
        RECT 208.950 689.400 250.050 690.450 ;
        RECT 208.950 688.950 211.050 689.400 ;
        RECT 247.950 688.950 250.050 689.400 ;
        RECT 283.950 690.450 286.050 691.050 ;
        RECT 310.950 690.450 313.050 691.050 ;
        RECT 361.950 690.450 364.050 691.050 ;
        RECT 283.950 689.400 364.050 690.450 ;
        RECT 283.950 688.950 286.050 689.400 ;
        RECT 310.950 688.950 313.050 689.400 ;
        RECT 361.950 688.950 364.050 689.400 ;
        RECT 430.950 690.450 433.050 691.050 ;
        RECT 439.950 690.450 442.050 691.050 ;
        RECT 430.950 689.400 442.050 690.450 ;
        RECT 430.950 688.950 433.050 689.400 ;
        RECT 439.950 688.950 442.050 689.400 ;
        RECT 583.950 690.450 586.050 691.050 ;
        RECT 598.950 690.450 601.050 691.050 ;
        RECT 583.950 689.400 601.050 690.450 ;
        RECT 583.950 688.950 586.050 689.400 ;
        RECT 598.950 688.950 601.050 689.400 ;
        RECT 679.950 690.450 682.050 691.050 ;
        RECT 715.950 690.450 718.050 691.050 ;
        RECT 724.950 690.450 727.050 691.050 ;
        RECT 679.950 689.400 693.450 690.450 ;
        RECT 679.950 688.950 682.050 689.400 ;
        RECT 241.950 687.450 244.050 688.050 ;
        RECT 253.950 687.450 256.050 688.050 ;
        RECT 241.950 686.400 256.050 687.450 ;
        RECT 241.950 685.950 244.050 686.400 ;
        RECT 253.950 685.950 256.050 686.400 ;
        RECT 343.950 687.450 346.050 688.050 ;
        RECT 505.950 687.450 508.050 688.050 ;
        RECT 343.950 686.400 508.050 687.450 ;
        RECT 343.950 685.950 346.050 686.400 ;
        RECT 505.950 685.950 508.050 686.400 ;
        RECT 652.950 687.450 655.050 688.050 ;
        RECT 688.950 687.450 691.050 688.050 ;
        RECT 652.950 686.400 691.050 687.450 ;
        RECT 692.400 687.450 693.450 689.400 ;
        RECT 715.950 689.400 727.050 690.450 ;
        RECT 715.950 688.950 718.050 689.400 ;
        RECT 724.950 688.950 727.050 689.400 ;
        RECT 799.950 690.450 802.050 691.050 ;
        RECT 799.950 689.400 813.450 690.450 ;
        RECT 799.950 688.950 802.050 689.400 ;
        RECT 775.950 687.450 778.050 688.050 ;
        RECT 692.400 686.400 778.050 687.450 ;
        RECT 812.400 687.450 813.450 689.400 ;
        RECT 826.950 687.450 829.050 688.050 ;
        RECT 812.400 686.400 829.050 687.450 ;
        RECT 652.950 685.950 655.050 686.400 ;
        RECT 688.950 685.950 691.050 686.400 ;
        RECT 775.950 685.950 778.050 686.400 ;
        RECT 826.950 685.950 829.050 686.400 ;
        RECT 76.950 684.450 79.050 685.050 ;
        RECT 148.950 684.450 151.050 685.050 ;
        RECT 76.950 683.400 151.050 684.450 ;
        RECT 76.950 682.950 79.050 683.400 ;
        RECT 148.950 682.950 151.050 683.400 ;
        RECT 244.950 684.450 247.050 685.050 ;
        RECT 262.950 684.450 265.050 685.050 ;
        RECT 244.950 683.400 265.050 684.450 ;
        RECT 244.950 682.950 247.050 683.400 ;
        RECT 262.950 682.950 265.050 683.400 ;
        RECT 352.950 684.450 355.050 685.050 ;
        RECT 412.950 684.450 415.050 685.050 ;
        RECT 352.950 683.400 415.050 684.450 ;
        RECT 352.950 682.950 355.050 683.400 ;
        RECT 412.950 682.950 415.050 683.400 ;
        RECT 445.950 684.450 448.050 685.050 ;
        RECT 496.950 684.450 499.050 685.050 ;
        RECT 535.950 684.450 538.050 685.050 ;
        RECT 445.950 683.400 538.050 684.450 ;
        RECT 445.950 682.950 448.050 683.400 ;
        RECT 496.950 682.950 499.050 683.400 ;
        RECT 535.950 682.950 538.050 683.400 ;
        RECT 604.950 684.450 607.050 685.050 ;
        RECT 679.950 684.450 682.050 685.200 ;
        RECT 604.950 683.400 682.050 684.450 ;
        RECT 604.950 682.950 607.050 683.400 ;
        RECT 679.950 683.100 682.050 683.400 ;
        RECT 700.950 684.450 703.050 685.050 ;
        RECT 709.950 684.450 712.050 685.050 ;
        RECT 700.950 683.400 712.050 684.450 ;
        RECT 700.950 682.950 703.050 683.400 ;
        RECT 709.950 682.950 712.050 683.400 ;
        RECT 718.950 684.450 721.050 685.050 ;
        RECT 766.950 684.450 769.050 685.050 ;
        RECT 799.950 684.450 802.050 685.050 ;
        RECT 718.950 683.400 802.050 684.450 ;
        RECT 718.950 682.950 721.050 683.400 ;
        RECT 766.950 682.950 769.050 683.400 ;
        RECT 799.950 682.950 802.050 683.400 ;
        RECT 805.950 684.450 808.050 685.050 ;
        RECT 832.950 684.450 835.050 685.050 ;
        RECT 805.950 683.400 835.050 684.450 ;
        RECT 805.950 682.950 808.050 683.400 ;
        RECT 832.950 682.950 835.050 683.400 ;
        RECT 13.950 681.450 16.050 682.050 ;
        RECT 25.950 681.450 28.050 682.050 ;
        RECT 13.950 680.400 28.050 681.450 ;
        RECT 13.950 679.950 16.050 680.400 ;
        RECT 25.950 679.950 28.050 680.400 ;
        RECT 106.950 681.450 109.050 682.050 ;
        RECT 139.950 681.450 142.050 682.050 ;
        RECT 106.950 680.400 142.050 681.450 ;
        RECT 106.950 679.950 109.050 680.400 ;
        RECT 139.950 679.950 142.050 680.400 ;
        RECT 160.950 681.450 163.050 682.050 ;
        RECT 199.950 681.450 202.050 682.050 ;
        RECT 160.950 680.400 202.050 681.450 ;
        RECT 160.950 679.950 163.050 680.400 ;
        RECT 199.950 679.950 202.050 680.400 ;
        RECT 229.950 681.450 232.050 682.050 ;
        RECT 259.950 681.450 262.050 682.050 ;
        RECT 229.950 680.400 262.050 681.450 ;
        RECT 229.950 679.950 232.050 680.400 ;
        RECT 259.950 679.950 262.050 680.400 ;
        RECT 286.950 681.450 289.050 682.050 ;
        RECT 322.950 681.450 325.050 682.050 ;
        RECT 286.950 680.400 325.050 681.450 ;
        RECT 286.950 679.950 289.050 680.400 ;
        RECT 322.950 679.950 325.050 680.400 ;
        RECT 349.950 681.450 352.050 682.050 ;
        RECT 364.950 681.450 367.050 682.050 ;
        RECT 349.950 680.400 367.050 681.450 ;
        RECT 349.950 679.950 352.050 680.400 ;
        RECT 364.950 679.950 367.050 680.400 ;
        RECT 436.950 681.450 439.050 682.050 ;
        RECT 536.400 681.450 537.450 682.950 ;
        RECT 619.950 681.450 622.050 682.050 ;
        RECT 679.950 681.450 682.050 681.900 ;
        RECT 436.950 680.400 534.450 681.450 ;
        RECT 536.400 680.400 682.050 681.450 ;
        RECT 436.950 679.950 439.050 680.400 ;
        RECT 34.950 678.450 37.050 679.050 ;
        RECT 55.950 678.450 58.050 679.050 ;
        RECT 88.950 678.450 91.050 679.050 ;
        RECT 34.950 677.400 42.450 678.450 ;
        RECT 34.950 676.950 37.050 677.400 ;
        RECT 10.950 670.950 16.050 673.050 ;
        RECT 19.950 670.950 22.050 676.050 ;
        RECT 41.400 675.450 42.450 677.400 ;
        RECT 55.950 677.400 91.050 678.450 ;
        RECT 55.950 676.950 58.050 677.400 ;
        RECT 88.950 676.950 91.050 677.400 ;
        RECT 148.950 678.450 151.050 679.050 ;
        RECT 169.950 678.450 172.050 679.050 ;
        RECT 148.950 677.400 172.050 678.450 ;
        RECT 148.950 676.950 151.050 677.400 ;
        RECT 169.950 676.950 172.050 677.400 ;
        RECT 307.950 678.450 310.050 679.050 ;
        RECT 391.950 678.450 394.050 679.050 ;
        RECT 307.950 677.400 394.050 678.450 ;
        RECT 307.950 676.950 310.050 677.400 ;
        RECT 391.950 676.950 394.050 677.400 ;
        RECT 403.950 678.450 406.050 679.050 ;
        RECT 409.950 678.450 412.050 679.050 ;
        RECT 445.950 678.450 448.050 679.050 ;
        RECT 403.950 677.400 448.050 678.450 ;
        RECT 403.950 676.950 406.050 677.400 ;
        RECT 409.950 676.950 412.050 677.400 ;
        RECT 445.950 676.950 448.050 677.400 ;
        RECT 460.950 678.450 463.050 679.050 ;
        RECT 469.950 678.450 472.050 679.050 ;
        RECT 460.950 677.400 472.050 678.450 ;
        RECT 460.950 676.950 463.050 677.400 ;
        RECT 469.950 676.950 472.050 677.400 ;
        RECT 502.950 678.450 505.050 679.050 ;
        RECT 533.400 678.450 534.450 680.400 ;
        RECT 619.950 679.950 622.050 680.400 ;
        RECT 679.950 679.800 682.050 680.400 ;
        RECT 703.950 681.450 706.050 682.050 ;
        RECT 712.950 681.450 715.050 682.050 ;
        RECT 703.950 680.400 715.050 681.450 ;
        RECT 703.950 679.950 706.050 680.400 ;
        RECT 712.950 679.950 715.050 680.400 ;
        RECT 550.950 678.450 553.050 679.050 ;
        RECT 502.950 678.000 528.450 678.450 ;
        RECT 502.950 677.400 529.050 678.000 ;
        RECT 533.400 677.400 553.050 678.450 ;
        RECT 502.950 676.950 505.050 677.400 ;
        RECT 55.950 675.450 58.050 676.050 ;
        RECT 41.400 674.400 58.050 675.450 ;
        RECT 55.950 673.950 58.050 674.400 ;
        RECT 97.950 675.450 100.050 676.050 ;
        RECT 127.950 675.450 130.050 676.050 ;
        RECT 160.950 675.450 163.050 676.050 ;
        RECT 97.950 674.400 163.050 675.450 ;
        RECT 97.950 673.950 100.050 674.400 ;
        RECT 127.950 673.950 130.050 674.400 ;
        RECT 160.950 673.950 163.050 674.400 ;
        RECT 181.950 675.450 184.050 676.050 ;
        RECT 190.950 675.450 193.050 676.050 ;
        RECT 181.950 674.400 193.050 675.450 ;
        RECT 181.950 673.950 184.050 674.400 ;
        RECT 190.950 673.950 193.050 674.400 ;
        RECT 223.950 675.450 226.050 676.050 ;
        RECT 232.950 675.450 235.050 676.050 ;
        RECT 223.950 674.400 235.050 675.450 ;
        RECT 223.950 673.950 226.050 674.400 ;
        RECT 232.950 673.950 235.050 674.400 ;
        RECT 247.950 675.450 250.050 676.050 ;
        RECT 364.950 675.450 367.050 676.050 ;
        RECT 247.950 674.400 367.050 675.450 ;
        RECT 247.950 673.950 250.050 674.400 ;
        RECT 364.950 673.950 367.050 674.400 ;
        RECT 436.800 675.000 438.900 676.050 ;
        RECT 440.100 675.450 442.200 676.050 ;
        RECT 448.950 675.450 451.050 676.050 ;
        RECT 454.950 675.450 457.050 676.050 ;
        RECT 499.950 675.450 502.050 676.050 ;
        RECT 436.800 673.950 439.050 675.000 ;
        RECT 440.100 674.400 451.050 675.450 ;
        RECT 440.100 673.950 442.200 674.400 ;
        RECT 448.950 673.950 451.050 674.400 ;
        RECT 452.400 674.400 502.050 675.450 ;
        RECT 40.950 673.050 43.050 673.200 ;
        RECT 37.950 671.100 43.050 673.050 ;
        RECT 37.950 670.950 42.000 671.100 ;
        RECT 4.950 669.450 7.050 670.050 ;
        RECT 10.950 669.450 13.050 670.050 ;
        RECT 4.950 668.400 13.050 669.450 ;
        RECT 4.950 667.950 7.050 668.400 ;
        RECT 10.950 667.950 13.050 668.400 ;
        RECT 16.950 669.450 19.050 670.050 ;
        RECT 31.800 669.450 33.900 670.050 ;
        RECT 16.950 668.400 33.900 669.450 ;
        RECT 35.100 669.000 37.200 670.050 ;
        RECT 16.950 667.950 19.050 668.400 ;
        RECT 31.800 667.950 33.900 668.400 ;
        RECT 34.950 667.950 37.200 669.000 ;
        RECT 40.950 667.950 46.050 670.050 ;
        RECT 52.950 667.950 55.050 673.050 ;
        RECT 58.950 667.950 61.050 673.050 ;
        RECT 73.950 667.950 76.050 673.050 ;
        RECT 91.950 667.950 94.050 673.050 ;
        RECT 97.950 667.950 100.050 673.050 ;
        RECT 106.950 667.950 109.050 673.050 ;
        RECT 112.950 667.950 115.050 673.050 ;
        RECT 133.950 669.450 136.050 670.050 ;
        RECT 139.950 669.450 145.050 670.050 ;
        RECT 133.950 668.400 145.050 669.450 ;
        RECT 133.950 667.950 136.050 668.400 ;
        RECT 139.950 667.950 145.050 668.400 ;
        RECT 148.950 667.950 151.050 673.050 ;
        RECT 160.950 667.950 166.050 670.050 ;
        RECT 169.950 667.950 172.050 673.050 ;
        RECT 181.950 667.950 187.050 670.050 ;
        RECT 190.950 667.950 193.050 673.050 ;
        RECT 199.950 672.450 202.050 673.050 ;
        RECT 217.950 672.450 220.050 673.050 ;
        RECT 199.950 671.400 220.050 672.450 ;
        RECT 199.950 670.950 202.050 671.400 ;
        RECT 217.950 670.950 220.050 671.400 ;
        RECT 259.950 670.950 265.050 673.050 ;
        RECT 268.950 670.950 274.050 673.050 ;
        RECT 277.800 672.000 279.900 673.050 ;
        RECT 281.100 672.450 283.200 673.050 ;
        RECT 316.950 672.450 319.050 673.050 ;
        RECT 277.800 670.950 280.050 672.000 ;
        RECT 281.100 671.400 300.450 672.450 ;
        RECT 305.400 672.000 319.050 672.450 ;
        RECT 281.100 670.950 283.200 671.400 ;
        RECT 208.950 669.450 211.050 670.050 ;
        RECT 220.800 669.450 222.900 670.050 ;
        RECT 208.950 668.400 222.900 669.450 ;
        RECT 224.100 669.000 226.200 670.050 ;
        RECT 208.950 667.950 211.050 668.400 ;
        RECT 220.800 667.950 222.900 668.400 ;
        RECT 223.950 667.950 226.200 669.000 ;
        RECT 241.950 667.950 246.900 670.050 ;
        RECT 248.100 669.000 250.200 670.050 ;
        RECT 247.950 667.950 250.200 669.000 ;
        RECT 253.950 667.950 259.050 670.050 ;
        RECT 277.950 667.950 280.050 670.950 ;
        RECT 299.400 670.050 300.450 671.400 ;
        RECT 304.950 671.400 319.050 672.000 ;
        RECT 283.950 667.950 289.050 670.050 ;
        RECT 34.950 667.050 37.050 667.950 ;
        RECT 19.950 666.450 22.050 667.050 ;
        RECT 34.950 666.450 37.200 667.050 ;
        RECT 19.950 665.400 37.200 666.450 ;
        RECT 19.950 664.950 22.050 665.400 ;
        RECT 35.100 664.950 37.200 665.400 ;
        RECT 52.950 666.450 55.050 667.050 ;
        RECT 64.950 666.450 67.050 667.050 ;
        RECT 70.950 666.450 73.050 667.050 ;
        RECT 52.950 665.400 73.050 666.450 ;
        RECT 52.950 664.950 55.050 665.400 ;
        RECT 64.950 664.950 67.050 665.400 ;
        RECT 70.950 664.950 73.050 665.400 ;
        RECT 76.950 664.050 79.050 667.050 ;
        RECT 88.950 666.450 91.050 667.050 ;
        RECT 94.950 666.450 97.050 667.050 ;
        RECT 109.950 666.450 112.050 667.050 ;
        RECT 88.950 665.400 112.050 666.450 ;
        RECT 88.950 664.950 91.050 665.400 ;
        RECT 94.950 664.950 97.050 665.400 ;
        RECT 109.950 664.950 112.050 665.400 ;
        RECT 145.950 666.450 151.050 667.050 ;
        RECT 166.950 666.450 169.050 667.050 ;
        RECT 145.950 665.400 169.050 666.450 ;
        RECT 145.950 664.950 151.050 665.400 ;
        RECT 166.950 664.950 169.050 665.400 ;
        RECT 172.950 666.450 178.050 667.050 ;
        RECT 187.950 666.450 190.050 667.050 ;
        RECT 172.950 665.400 190.050 666.450 ;
        RECT 172.950 664.950 178.050 665.400 ;
        RECT 187.950 664.950 190.050 665.400 ;
        RECT 205.950 664.950 210.900 667.050 ;
        RECT 212.100 666.450 214.200 667.050 ;
        RECT 217.950 666.450 220.050 667.050 ;
        RECT 223.950 666.450 226.050 667.950 ;
        RECT 212.100 666.000 226.050 666.450 ;
        RECT 212.100 665.400 225.450 666.000 ;
        RECT 212.100 664.950 214.200 665.400 ;
        RECT 217.950 664.950 220.050 665.400 ;
        RECT 37.950 663.450 40.050 664.050 ;
        RECT 73.800 663.450 75.900 664.050 ;
        RECT 37.950 662.400 75.900 663.450 ;
        RECT 76.950 663.000 79.200 664.050 ;
        RECT 37.950 661.950 40.050 662.400 ;
        RECT 73.800 661.950 75.900 662.400 ;
        RECT 77.100 661.950 79.200 663.000 ;
        RECT 94.950 663.450 97.050 664.050 ;
        RECT 103.950 663.450 106.050 664.050 ;
        RECT 94.950 662.400 106.050 663.450 ;
        RECT 94.950 661.950 97.050 662.400 ;
        RECT 103.950 661.950 106.050 662.400 ;
        RECT 217.950 663.450 220.050 664.050 ;
        RECT 241.950 663.450 244.050 667.050 ;
        RECT 247.950 664.950 250.050 667.950 ;
        RECT 298.950 667.050 301.050 670.050 ;
        RECT 304.950 667.950 307.050 671.400 ;
        RECT 316.950 667.950 319.050 671.400 ;
        RECT 322.950 672.450 325.050 673.050 ;
        RECT 337.950 672.450 340.050 673.050 ;
        RECT 322.950 671.400 340.050 672.450 ;
        RECT 322.950 670.950 325.050 671.400 ;
        RECT 337.950 670.950 340.050 671.400 ;
        RECT 343.950 670.950 349.050 673.050 ;
        RECT 376.950 672.450 379.050 673.200 ;
        RECT 382.950 672.450 385.050 673.050 ;
        RECT 388.950 672.450 391.050 673.050 ;
        RECT 376.950 671.400 391.050 672.450 ;
        RECT 376.950 671.100 379.050 671.400 ;
        RECT 382.950 670.950 385.050 671.400 ;
        RECT 388.950 670.950 391.050 671.400 ;
        RECT 394.950 670.050 397.050 673.050 ;
        RECT 400.950 670.950 405.900 673.050 ;
        RECT 407.100 670.950 412.050 673.050 ;
        RECT 436.950 670.950 439.050 673.950 ;
        RECT 442.950 672.450 445.050 673.050 ;
        RECT 452.400 672.450 453.450 674.400 ;
        RECT 454.950 673.950 457.050 674.400 ;
        RECT 499.950 673.950 502.050 674.400 ;
        RECT 526.950 675.450 529.050 677.400 ;
        RECT 550.950 676.950 553.050 677.400 ;
        RECT 592.950 678.450 595.050 679.050 ;
        RECT 637.950 678.450 640.050 679.050 ;
        RECT 664.950 678.450 667.050 679.050 ;
        RECT 592.950 677.400 640.050 678.450 ;
        RECT 592.950 676.950 595.050 677.400 ;
        RECT 637.950 676.950 640.050 677.400 ;
        RECT 644.400 677.400 667.050 678.450 ;
        RECT 697.950 677.400 700.050 679.500 ;
        RECT 718.950 677.400 721.050 679.500 ;
        RECT 724.950 678.450 727.050 679.050 ;
        RECT 745.950 678.450 748.050 679.050 ;
        RECT 724.950 677.400 748.050 678.450 ;
        RECT 547.950 675.450 550.050 676.050 ;
        RECT 526.950 674.400 550.050 675.450 ;
        RECT 526.950 673.950 529.050 674.400 ;
        RECT 547.950 673.950 550.050 674.400 ;
        RECT 595.950 675.450 598.050 676.050 ;
        RECT 625.950 675.450 628.050 676.050 ;
        RECT 595.950 674.400 628.050 675.450 ;
        RECT 595.950 673.950 598.050 674.400 ;
        RECT 625.950 673.950 628.050 674.400 ;
        RECT 631.950 675.450 634.050 676.050 ;
        RECT 644.400 675.450 645.450 677.400 ;
        RECT 664.950 676.950 667.050 677.400 ;
        RECT 631.950 674.400 645.450 675.450 ;
        RECT 647.100 675.000 649.200 676.050 ;
        RECT 631.950 673.950 634.050 674.400 ;
        RECT 646.950 673.950 649.200 675.000 ;
        RECT 646.950 673.050 649.050 673.950 ;
        RECT 442.950 671.400 453.450 672.450 ;
        RECT 442.950 670.950 445.050 671.400 ;
        RECT 454.950 670.950 460.050 673.050 ;
        RECT 463.950 672.450 466.050 673.050 ;
        RECT 481.800 672.450 483.900 673.050 ;
        RECT 463.950 671.400 483.900 672.450 ;
        RECT 463.950 670.950 466.050 671.400 ;
        RECT 481.800 670.950 483.900 671.400 ;
        RECT 485.100 670.950 490.050 673.050 ;
        RECT 496.950 672.450 499.050 673.050 ;
        RECT 505.950 672.450 508.050 673.050 ;
        RECT 496.950 671.400 508.050 672.450 ;
        RECT 496.950 670.950 499.050 671.400 ;
        RECT 505.950 670.950 508.050 671.400 ;
        RECT 511.950 672.450 514.050 673.050 ;
        RECT 529.950 672.450 532.050 673.050 ;
        RECT 547.950 672.450 552.900 673.050 ;
        RECT 511.950 671.400 552.900 672.450 ;
        RECT 511.950 670.950 514.050 671.400 ;
        RECT 529.950 670.950 532.050 671.400 ;
        RECT 547.950 670.950 552.900 671.400 ;
        RECT 554.100 670.950 559.050 673.050 ;
        RECT 583.950 672.450 586.050 673.050 ;
        RECT 575.400 672.000 586.050 672.450 ;
        RECT 574.950 671.400 586.050 672.000 ;
        RECT 334.800 669.000 336.900 670.050 ;
        RECT 334.800 667.950 337.050 669.000 ;
        RECT 338.100 667.950 343.050 670.050 ;
        RECT 358.950 667.950 364.050 670.050 ;
        RECT 376.950 667.950 382.050 670.050 ;
        RECT 394.800 669.000 397.050 670.050 ;
        RECT 398.100 669.000 400.200 670.050 ;
        RECT 394.800 667.950 396.900 669.000 ;
        RECT 397.950 667.950 400.200 669.000 ;
        RECT 334.950 667.050 337.050 667.950 ;
        RECT 289.950 664.950 295.050 667.050 ;
        RECT 298.800 666.000 301.050 667.050 ;
        RECT 302.100 666.000 304.200 667.050 ;
        RECT 298.800 664.950 300.900 666.000 ;
        RECT 301.950 664.950 304.200 666.000 ;
        RECT 217.950 663.000 244.050 663.450 ;
        RECT 289.950 663.450 292.050 664.050 ;
        RECT 301.950 663.450 304.050 664.950 ;
        RECT 313.950 663.450 316.050 667.050 ;
        RECT 319.950 664.950 322.050 667.050 ;
        RECT 334.800 666.000 337.050 667.050 ;
        RECT 334.800 664.950 336.900 666.000 ;
        RECT 289.950 663.000 304.050 663.450 ;
        RECT 305.400 663.000 316.050 663.450 ;
        RECT 217.950 662.400 243.450 663.000 ;
        RECT 289.950 662.400 303.600 663.000 ;
        RECT 305.400 662.400 315.450 663.000 ;
        RECT 217.950 661.950 220.050 662.400 ;
        RECT 289.950 661.950 292.050 662.400 ;
        RECT 121.950 660.450 124.050 661.050 ;
        RECT 160.950 660.450 163.050 661.050 ;
        RECT 121.950 659.400 163.050 660.450 ;
        RECT 121.950 658.950 124.050 659.400 ;
        RECT 160.950 658.950 163.050 659.400 ;
        RECT 286.950 660.450 289.050 661.050 ;
        RECT 305.400 660.450 306.450 662.400 ;
        RECT 286.950 659.400 306.450 660.450 ;
        RECT 307.950 660.450 310.050 661.050 ;
        RECT 320.400 660.450 321.450 664.950 ;
        RECT 355.950 661.950 358.050 667.050 ;
        RECT 361.950 666.450 364.050 667.050 ;
        RECT 367.950 666.450 370.050 667.050 ;
        RECT 361.950 665.400 370.050 666.450 ;
        RECT 380.400 666.450 381.450 667.950 ;
        RECT 397.950 666.450 400.050 667.950 ;
        RECT 380.400 666.000 400.050 666.450 ;
        RECT 380.400 665.400 399.600 666.000 ;
        RECT 361.950 664.950 364.050 665.400 ;
        RECT 367.950 664.950 370.050 665.400 ;
        RECT 403.950 664.950 406.050 670.050 ;
        RECT 415.950 667.950 421.050 670.050 ;
        RECT 472.800 669.000 474.900 670.050 ;
        RECT 472.800 667.950 475.050 669.000 ;
        RECT 476.100 667.950 481.050 670.050 ;
        RECT 484.950 669.450 487.050 670.050 ;
        RECT 490.950 669.450 493.050 670.050 ;
        RECT 484.950 668.400 493.050 669.450 ;
        RECT 484.950 667.950 487.050 668.400 ;
        RECT 490.950 667.950 493.050 668.400 ;
        RECT 499.950 669.450 502.050 670.050 ;
        RECT 508.950 669.450 511.050 670.050 ;
        RECT 499.950 668.400 511.050 669.450 ;
        RECT 499.950 667.950 502.050 668.400 ;
        RECT 409.950 666.450 412.050 667.050 ;
        RECT 415.950 666.450 418.050 667.050 ;
        RECT 409.950 665.400 418.050 666.450 ;
        RECT 409.950 664.950 412.050 665.400 ;
        RECT 415.950 664.950 418.050 665.400 ;
        RECT 421.950 664.950 427.050 667.050 ;
        RECT 472.950 664.950 475.050 667.950 ;
        RECT 478.950 666.450 481.050 667.050 ;
        RECT 484.950 666.450 487.050 667.050 ;
        RECT 478.950 665.400 487.050 666.450 ;
        RECT 508.950 666.450 511.050 668.400 ;
        RECT 514.950 667.950 520.050 670.050 ;
        RECT 532.950 667.950 538.050 670.050 ;
        RECT 547.950 667.950 553.050 670.050 ;
        RECT 556.950 669.450 559.050 670.050 ;
        RECT 568.950 669.450 571.050 670.050 ;
        RECT 556.950 668.400 571.050 669.450 ;
        RECT 556.950 667.950 559.050 668.400 ;
        RECT 568.950 667.950 571.050 668.400 ;
        RECT 574.950 667.950 577.050 671.400 ;
        RECT 583.950 670.950 586.050 671.400 ;
        RECT 589.950 670.950 594.900 673.050 ;
        RECT 596.100 672.450 598.200 673.050 ;
        RECT 604.950 672.450 610.050 673.050 ;
        RECT 596.100 671.400 610.050 672.450 ;
        RECT 596.100 670.950 598.200 671.400 ;
        RECT 604.950 670.950 610.050 671.400 ;
        RECT 616.950 672.450 619.050 673.050 ;
        RECT 643.800 672.450 645.900 673.050 ;
        RECT 616.950 671.400 645.900 672.450 ;
        RECT 646.950 672.000 649.200 673.050 ;
        RECT 616.950 670.950 619.050 671.400 ;
        RECT 643.800 670.950 645.900 671.400 ;
        RECT 647.100 670.950 649.200 672.000 ;
        RECT 652.950 672.450 655.050 673.050 ;
        RECT 691.800 672.450 693.900 673.050 ;
        RECT 652.950 671.400 693.900 672.450 ;
        RECT 695.100 672.000 697.200 673.050 ;
        RECT 652.950 670.950 655.050 671.400 ;
        RECT 691.800 670.950 693.900 671.400 ;
        RECT 694.950 670.950 697.200 672.000 ;
        RECT 628.950 669.450 631.050 670.050 ;
        RECT 643.800 669.450 645.900 670.050 ;
        RECT 628.950 668.400 645.900 669.450 ;
        RECT 628.950 667.950 631.050 668.400 ;
        RECT 643.800 667.950 645.900 668.400 ;
        RECT 647.100 667.950 652.050 670.050 ;
        RECT 685.950 667.950 691.050 670.050 ;
        RECT 694.950 669.450 697.050 670.950 ;
        RECT 692.400 668.400 697.050 669.450 ;
        RECT 526.950 666.450 529.050 667.050 ;
        RECT 508.950 666.000 529.050 666.450 ;
        RECT 509.400 665.400 529.050 666.000 ;
        RECT 478.950 664.950 481.050 665.400 ;
        RECT 484.950 664.950 487.050 665.400 ;
        RECT 526.950 664.950 529.050 665.400 ;
        RECT 571.950 664.950 576.900 667.050 ;
        RECT 578.100 666.000 580.200 667.050 ;
        RECT 577.950 664.950 580.200 666.000 ;
        RECT 616.950 666.450 619.050 667.050 ;
        RECT 625.950 666.450 628.050 667.050 ;
        RECT 616.950 665.400 628.050 666.450 ;
        RECT 616.950 664.950 619.050 665.400 ;
        RECT 625.950 664.950 628.050 665.400 ;
        RECT 382.950 663.450 385.050 664.050 ;
        RECT 388.950 663.450 391.050 664.050 ;
        RECT 382.950 662.400 391.050 663.450 ;
        RECT 382.950 661.950 385.050 662.400 ;
        RECT 388.950 661.950 391.050 662.400 ;
        RECT 394.950 663.450 397.050 664.050 ;
        RECT 410.400 663.450 411.450 664.950 ;
        RECT 484.950 663.450 487.050 664.050 ;
        RECT 577.950 663.450 580.050 664.950 ;
        RECT 589.950 663.450 592.050 664.050 ;
        RECT 394.950 662.400 592.050 663.450 ;
        RECT 394.950 661.950 397.050 662.400 ;
        RECT 484.950 661.950 487.050 662.400 ;
        RECT 589.950 661.950 592.050 662.400 ;
        RECT 598.950 663.450 601.050 664.050 ;
        RECT 631.950 663.450 634.050 667.050 ;
        RECT 679.950 666.450 682.050 667.050 ;
        RECT 692.400 666.450 693.450 668.400 ;
        RECT 694.950 667.950 697.050 668.400 ;
        RECT 679.950 665.400 693.450 666.450 ;
        RECT 698.850 665.400 700.050 677.400 ;
        RECT 703.950 670.950 708.900 673.050 ;
        RECT 710.100 670.950 715.050 673.050 ;
        RECT 679.950 664.950 682.050 665.400 ;
        RECT 598.950 663.000 634.050 663.450 ;
        RECT 664.950 663.450 667.050 664.050 ;
        RECT 688.950 663.450 691.050 664.050 ;
        RECT 598.950 662.400 633.450 663.000 ;
        RECT 664.950 662.400 691.050 663.450 ;
        RECT 697.950 663.300 700.050 665.400 ;
        RECT 706.950 666.450 709.050 667.050 ;
        RECT 712.950 666.450 715.050 667.050 ;
        RECT 706.950 665.400 715.050 666.450 ;
        RECT 706.950 664.950 709.050 665.400 ;
        RECT 712.950 664.950 715.050 665.400 ;
        RECT 598.950 661.950 601.050 662.400 ;
        RECT 664.950 661.950 667.050 662.400 ;
        RECT 688.950 661.950 691.050 662.400 ;
        RECT 307.950 659.400 321.450 660.450 ;
        RECT 334.950 660.450 337.050 661.200 ;
        RECT 361.950 660.450 364.050 661.050 ;
        RECT 334.950 659.400 364.050 660.450 ;
        RECT 286.950 658.950 289.050 659.400 ;
        RECT 307.950 658.950 310.050 659.400 ;
        RECT 334.950 659.100 337.050 659.400 ;
        RECT 361.950 658.950 364.050 659.400 ;
        RECT 403.950 660.450 406.050 661.050 ;
        RECT 424.950 660.450 427.050 661.050 ;
        RECT 403.950 659.400 427.050 660.450 ;
        RECT 403.950 658.950 406.050 659.400 ;
        RECT 424.950 658.950 427.050 659.400 ;
        RECT 472.950 660.450 475.050 661.050 ;
        RECT 490.950 660.450 493.050 661.050 ;
        RECT 472.950 659.400 493.050 660.450 ;
        RECT 472.950 658.950 475.050 659.400 ;
        RECT 490.950 658.950 493.050 659.400 ;
        RECT 511.950 660.450 514.050 661.050 ;
        RECT 574.950 660.450 577.050 661.050 ;
        RECT 511.950 659.400 577.050 660.450 ;
        RECT 698.850 659.700 700.050 663.300 ;
        RECT 719.100 660.600 720.300 677.400 ;
        RECT 724.950 676.950 727.050 677.400 ;
        RECT 745.950 676.950 748.050 677.400 ;
        RECT 757.950 678.450 760.050 679.050 ;
        RECT 781.950 678.450 784.050 679.050 ;
        RECT 757.950 677.400 784.050 678.450 ;
        RECT 790.950 677.400 793.050 679.500 ;
        RECT 811.950 677.400 814.050 679.500 ;
        RECT 757.950 676.950 760.050 677.400 ;
        RECT 781.950 676.950 784.050 677.400 ;
        RECT 772.950 675.450 775.050 676.050 ;
        RECT 746.400 675.000 775.050 675.450 ;
        RECT 745.950 674.400 775.050 675.000 ;
        RECT 730.950 672.450 733.050 673.050 ;
        RECT 739.950 672.450 742.050 673.050 ;
        RECT 730.950 671.400 742.050 672.450 ;
        RECT 730.950 670.950 733.050 671.400 ;
        RECT 739.950 670.950 742.050 671.400 ;
        RECT 745.950 670.950 748.050 674.400 ;
        RECT 772.950 673.950 775.050 674.400 ;
        RECT 749.400 671.400 762.450 672.450 ;
        RECT 736.950 664.950 739.050 670.050 ;
        RECT 742.950 669.450 745.050 670.050 ;
        RECT 749.400 669.450 750.450 671.400 ;
        RECT 761.400 670.050 762.450 671.400 ;
        RECT 772.950 670.950 777.900 673.050 ;
        RECT 779.100 670.950 784.050 673.050 ;
        RECT 742.950 668.400 750.450 669.450 ;
        RECT 742.950 667.950 745.050 668.400 ;
        RECT 754.950 667.950 759.900 670.050 ;
        RECT 761.100 669.000 763.200 670.050 ;
        RECT 760.950 667.950 763.200 669.000 ;
        RECT 787.950 667.950 790.050 673.050 ;
        RECT 751.950 664.950 757.050 667.050 ;
        RECT 760.950 664.950 763.050 667.950 ;
        RECT 791.850 665.400 793.050 677.400 ;
        RECT 796.950 670.950 802.050 673.050 ;
        RECT 805.950 667.950 808.050 673.050 ;
        RECT 736.950 663.450 739.050 664.050 ;
        RECT 754.950 663.450 757.050 664.050 ;
        RECT 736.950 662.400 757.050 663.450 ;
        RECT 790.950 663.300 793.050 665.400 ;
        RECT 736.950 661.950 739.050 662.400 ;
        RECT 754.950 661.950 757.050 662.400 ;
        RECT 511.950 658.950 514.050 659.400 ;
        RECT 574.950 658.950 577.050 659.400 ;
        RECT 301.950 657.450 304.050 658.050 ;
        RECT 334.950 657.450 337.050 657.900 ;
        RECT 301.950 656.400 337.050 657.450 ;
        RECT 301.950 655.950 304.050 656.400 ;
        RECT 334.950 655.800 337.050 656.400 ;
        RECT 343.950 657.450 346.050 658.050 ;
        RECT 349.950 657.450 352.050 658.050 ;
        RECT 343.950 656.400 352.050 657.450 ;
        RECT 343.950 655.950 346.050 656.400 ;
        RECT 349.950 655.950 352.050 656.400 ;
        RECT 376.950 657.450 379.050 658.050 ;
        RECT 463.950 657.450 466.050 658.050 ;
        RECT 376.950 656.400 466.050 657.450 ;
        RECT 376.950 655.950 379.050 656.400 ;
        RECT 463.950 655.950 466.050 656.400 ;
        RECT 649.950 657.450 652.050 658.050 ;
        RECT 658.950 657.450 661.050 658.050 ;
        RECT 697.950 657.600 700.050 659.700 ;
        RECT 718.950 658.500 721.050 660.600 ;
        RECT 791.850 659.700 793.050 663.300 ;
        RECT 812.100 660.600 813.300 677.400 ;
        RECT 820.950 672.450 823.050 673.050 ;
        RECT 826.950 672.450 829.050 673.050 ;
        RECT 820.950 671.400 829.050 672.450 ;
        RECT 820.950 670.950 823.050 671.400 ;
        RECT 826.950 670.950 829.050 671.400 ;
        RECT 832.950 670.950 838.050 673.050 ;
        RECT 817.950 669.450 820.050 670.050 ;
        RECT 829.950 669.450 832.050 670.050 ;
        RECT 817.950 668.400 832.050 669.450 ;
        RECT 817.950 667.950 820.050 668.400 ;
        RECT 829.950 667.950 832.050 668.400 ;
        RECT 820.950 666.450 823.050 667.050 ;
        RECT 835.950 666.450 838.050 670.050 ;
        RECT 820.950 666.000 838.050 666.450 ;
        RECT 820.950 665.400 837.450 666.000 ;
        RECT 820.950 664.950 823.050 665.400 ;
        RECT 814.950 663.450 817.050 664.050 ;
        RECT 841.950 663.450 844.050 664.050 ;
        RECT 814.950 662.400 844.050 663.450 ;
        RECT 814.950 661.950 817.050 662.400 ;
        RECT 841.950 661.950 844.050 662.400 ;
        RECT 790.950 657.600 793.050 659.700 ;
        RECT 811.950 658.500 814.050 660.600 ;
        RECT 649.950 656.400 661.050 657.450 ;
        RECT 649.950 655.950 652.050 656.400 ;
        RECT 658.950 655.950 661.050 656.400 ;
        RECT 82.950 654.450 85.050 655.050 ;
        RECT 145.950 654.450 148.050 655.050 ;
        RECT 82.950 653.400 148.050 654.450 ;
        RECT 82.950 652.950 85.050 653.400 ;
        RECT 145.950 652.950 148.050 653.400 ;
        RECT 157.950 654.450 160.050 655.050 ;
        RECT 169.950 654.450 172.050 655.050 ;
        RECT 157.950 653.400 172.050 654.450 ;
        RECT 157.950 652.950 160.050 653.400 ;
        RECT 169.950 652.950 172.050 653.400 ;
        RECT 286.950 654.450 289.050 655.050 ;
        RECT 394.950 654.450 397.050 655.050 ;
        RECT 400.950 654.450 403.050 655.050 ;
        RECT 430.950 654.450 433.050 655.050 ;
        RECT 286.950 653.400 433.050 654.450 ;
        RECT 286.950 652.950 289.050 653.400 ;
        RECT 394.950 652.950 397.050 653.400 ;
        RECT 400.950 652.950 403.050 653.400 ;
        RECT 430.950 652.950 433.050 653.400 ;
        RECT 547.950 654.450 550.050 655.050 ;
        RECT 568.950 654.450 571.050 655.050 ;
        RECT 673.950 654.450 676.050 655.050 ;
        RECT 547.950 653.400 571.050 654.450 ;
        RECT 547.950 652.950 550.050 653.400 ;
        RECT 568.950 652.950 571.050 653.400 ;
        RECT 599.400 653.400 676.050 654.450 ;
        RECT 289.950 651.450 292.050 652.050 ;
        RECT 337.950 651.450 340.050 652.050 ;
        RECT 289.950 650.400 340.050 651.450 ;
        RECT 289.950 649.950 292.050 650.400 ;
        RECT 337.950 649.950 340.050 650.400 ;
        RECT 361.950 651.450 364.050 652.050 ;
        RECT 457.950 651.450 460.050 652.050 ;
        RECT 599.400 651.450 600.450 653.400 ;
        RECT 673.950 652.950 676.050 653.400 ;
        RECT 685.950 654.450 688.050 655.050 ;
        RECT 703.950 654.450 706.050 655.050 ;
        RECT 718.950 654.450 721.050 655.050 ;
        RECT 685.950 653.400 721.050 654.450 ;
        RECT 685.950 652.950 688.050 653.400 ;
        RECT 703.950 652.950 706.050 653.400 ;
        RECT 718.950 652.950 721.050 653.400 ;
        RECT 361.950 650.400 460.050 651.450 ;
        RECT 361.950 649.950 364.050 650.400 ;
        RECT 457.950 649.950 460.050 650.400 ;
        RECT 548.400 650.400 600.450 651.450 ;
        RECT 601.950 651.450 604.050 652.050 ;
        RECT 700.950 651.450 703.050 652.050 ;
        RECT 751.950 651.450 754.050 652.050 ;
        RECT 760.950 651.450 763.050 652.050 ;
        RECT 601.950 650.400 703.050 651.450 ;
        RECT 70.950 648.450 73.050 649.050 ;
        RECT 109.950 648.450 112.050 649.050 ;
        RECT 70.950 647.400 112.050 648.450 ;
        RECT 70.950 646.950 73.050 647.400 ;
        RECT 109.950 646.950 112.050 647.400 ;
        RECT 235.950 648.450 238.050 649.050 ;
        RECT 376.950 648.450 379.050 649.050 ;
        RECT 235.950 647.400 379.050 648.450 ;
        RECT 235.950 646.950 238.050 647.400 ;
        RECT 376.950 646.950 379.050 647.400 ;
        RECT 442.950 648.450 445.050 649.050 ;
        RECT 548.400 648.450 549.450 650.400 ;
        RECT 601.950 649.950 604.050 650.400 ;
        RECT 700.950 649.950 703.050 650.400 ;
        RECT 707.400 650.400 763.050 651.450 ;
        RECT 442.950 647.400 549.450 648.450 ;
        RECT 550.950 648.450 553.050 649.050 ;
        RECT 562.950 648.450 565.050 649.050 ;
        RECT 550.950 647.400 565.050 648.450 ;
        RECT 442.950 646.950 445.050 647.400 ;
        RECT 550.950 646.950 553.050 647.400 ;
        RECT 562.950 646.950 565.050 647.400 ;
        RECT 655.950 648.450 658.050 649.050 ;
        RECT 682.950 648.450 685.050 649.050 ;
        RECT 655.950 647.400 685.050 648.450 ;
        RECT 655.950 646.950 658.050 647.400 ;
        RECT 682.950 646.950 685.050 647.400 ;
        RECT 694.950 648.450 697.050 649.050 ;
        RECT 707.400 648.450 708.450 650.400 ;
        RECT 751.950 649.950 754.050 650.400 ;
        RECT 760.950 649.950 763.050 650.400 ;
        RECT 694.950 647.400 708.450 648.450 ;
        RECT 709.950 648.450 712.050 649.050 ;
        RECT 730.950 648.450 733.050 649.050 ;
        RECT 709.950 647.400 733.050 648.450 ;
        RECT 694.950 646.950 697.050 647.400 ;
        RECT 709.950 646.950 712.050 647.400 ;
        RECT 730.950 646.950 733.050 647.400 ;
        RECT 754.950 648.450 757.050 649.050 ;
        RECT 790.950 648.450 793.050 649.050 ;
        RECT 754.950 647.400 793.050 648.450 ;
        RECT 754.950 646.950 757.050 647.400 ;
        RECT 790.950 646.950 793.050 647.400 ;
        RECT 40.950 645.450 43.050 646.050 ;
        RECT 85.950 645.450 88.050 646.050 ;
        RECT 166.950 645.450 169.050 646.050 ;
        RECT 40.950 644.400 169.050 645.450 ;
        RECT 40.950 643.950 43.050 644.400 ;
        RECT 85.950 643.950 88.050 644.400 ;
        RECT 166.950 643.950 169.050 644.400 ;
        RECT 253.950 645.450 256.050 646.050 ;
        RECT 310.950 645.450 313.050 646.050 ;
        RECT 253.950 644.400 313.050 645.450 ;
        RECT 253.950 643.950 256.050 644.400 ;
        RECT 310.950 643.950 313.050 644.400 ;
        RECT 355.950 645.450 360.000 646.050 ;
        RECT 403.950 645.450 406.050 646.050 ;
        RECT 409.950 645.450 412.050 646.050 ;
        RECT 355.950 643.950 360.450 645.450 ;
        RECT 403.950 644.400 412.050 645.450 ;
        RECT 403.950 643.950 406.050 644.400 ;
        RECT 409.950 643.950 412.050 644.400 ;
        RECT 457.950 645.450 460.050 646.050 ;
        RECT 787.950 645.450 790.050 646.050 ;
        RECT 838.950 645.450 841.050 646.050 ;
        RECT 457.950 644.400 841.050 645.450 ;
        RECT 457.950 643.950 460.050 644.400 ;
        RECT 787.950 643.950 790.050 644.400 ;
        RECT 838.950 643.950 841.050 644.400 ;
        RECT 359.400 643.050 360.450 643.950 ;
        RECT 58.950 642.450 61.050 643.050 ;
        RECT 76.950 642.450 79.050 643.050 ;
        RECT 91.950 642.450 94.050 643.050 ;
        RECT 229.950 642.450 232.050 643.050 ;
        RECT 58.950 641.400 232.050 642.450 ;
        RECT 58.950 640.950 61.050 641.400 ;
        RECT 76.950 640.950 79.050 641.400 ;
        RECT 91.950 640.950 94.050 641.400 ;
        RECT 229.950 640.950 232.050 641.400 ;
        RECT 358.950 642.450 361.050 643.050 ;
        RECT 463.950 642.450 466.050 643.050 ;
        RECT 358.950 641.400 466.050 642.450 ;
        RECT 358.950 640.950 361.050 641.400 ;
        RECT 463.950 640.950 466.050 641.400 ;
        RECT 484.950 642.450 487.050 643.050 ;
        RECT 511.950 642.450 514.050 643.050 ;
        RECT 484.950 641.400 514.050 642.450 ;
        RECT 484.950 640.950 487.050 641.400 ;
        RECT 511.950 640.950 514.050 641.400 ;
        RECT 523.950 642.450 526.050 643.050 ;
        RECT 607.950 642.450 610.050 643.050 ;
        RECT 523.950 641.400 610.050 642.450 ;
        RECT 523.950 640.950 526.050 641.400 ;
        RECT 607.950 640.950 610.050 641.400 ;
        RECT 37.950 639.450 40.050 640.050 ;
        RECT 127.950 639.450 130.050 640.050 ;
        RECT 37.950 638.400 130.050 639.450 ;
        RECT 37.950 637.950 40.050 638.400 ;
        RECT 127.950 637.950 130.050 638.400 ;
        RECT 241.950 639.450 244.050 640.050 ;
        RECT 262.950 639.450 265.050 640.050 ;
        RECT 241.950 638.400 265.050 639.450 ;
        RECT 241.950 637.950 244.050 638.400 ;
        RECT 262.950 637.950 265.050 638.400 ;
        RECT 274.950 639.450 277.050 640.050 ;
        RECT 322.950 639.450 325.050 640.050 ;
        RECT 355.950 639.450 358.050 640.050 ;
        RECT 274.950 638.400 358.050 639.450 ;
        RECT 274.950 637.950 277.050 638.400 ;
        RECT 322.950 637.950 325.050 638.400 ;
        RECT 355.950 637.950 358.050 638.400 ;
        RECT 424.950 639.450 427.050 640.050 ;
        RECT 472.950 639.450 475.050 640.050 ;
        RECT 625.950 639.450 628.050 640.050 ;
        RECT 424.950 638.400 628.050 639.450 ;
        RECT 670.950 639.300 673.050 641.400 ;
        RECT 424.950 637.950 427.050 638.400 ;
        RECT 472.950 637.950 475.050 638.400 ;
        RECT 625.950 637.950 628.050 638.400 ;
        RECT 13.950 636.450 16.050 637.050 ;
        RECT 37.950 636.450 40.050 637.050 ;
        RECT 13.950 635.400 40.050 636.450 ;
        RECT 13.950 634.950 16.050 635.400 ;
        RECT 13.950 628.950 16.050 634.050 ;
        RECT 25.950 631.950 31.050 634.050 ;
        RECT 37.950 631.950 40.050 635.400 ;
        RECT 52.950 631.950 55.050 637.050 ;
        RECT 70.950 636.450 73.050 637.050 ;
        RECT 94.950 636.450 97.050 637.050 ;
        RECT 100.950 636.450 103.050 637.050 ;
        RECT 205.950 636.450 208.050 637.050 ;
        RECT 70.950 636.000 78.450 636.450 ;
        RECT 70.950 635.400 79.050 636.000 ;
        RECT 70.950 634.950 73.050 635.400 ;
        RECT 58.950 631.050 61.050 634.050 ;
        RECT 64.950 631.950 70.050 634.050 ;
        RECT 76.950 631.950 79.050 635.400 ;
        RECT 94.950 635.400 103.050 636.450 ;
        RECT 134.400 636.000 147.450 636.450 ;
        RECT 182.250 636.000 208.050 636.450 ;
        RECT 94.950 634.950 97.050 635.400 ;
        RECT 100.950 634.950 103.050 635.400 ;
        RECT 133.950 635.400 147.450 636.000 ;
        RECT 133.950 633.450 136.050 635.400 ;
        RECT 122.400 633.000 136.050 633.450 ;
        RECT 121.950 632.400 136.050 633.000 ;
        RECT 19.950 628.950 25.050 631.050 ;
        RECT 34.950 630.450 39.000 631.050 ;
        RECT 34.950 628.950 39.450 630.450 ;
        RECT 40.950 628.950 46.050 631.050 ;
        RECT 55.800 630.450 57.900 631.050 ;
        RECT 47.400 629.400 57.900 630.450 ;
        RECT 58.950 630.000 61.200 631.050 ;
        RECT 10.950 627.450 13.050 628.050 ;
        RECT 31.950 627.450 34.050 628.050 ;
        RECT 10.950 626.400 34.050 627.450 ;
        RECT 10.950 625.950 13.050 626.400 ;
        RECT 31.950 625.950 34.050 626.400 ;
        RECT 38.400 627.450 39.450 628.950 ;
        RECT 47.400 627.450 48.450 629.400 ;
        RECT 55.800 628.950 57.900 629.400 ;
        RECT 59.100 628.950 61.200 630.000 ;
        RECT 38.400 626.400 48.450 627.450 ;
        RECT 73.950 627.450 76.050 631.050 ;
        RECT 79.950 630.450 82.050 631.050 ;
        RECT 91.950 630.450 96.900 631.050 ;
        RECT 79.950 629.400 96.900 630.450 ;
        RECT 79.950 628.950 82.050 629.400 ;
        RECT 91.950 628.950 96.900 629.400 ;
        RECT 98.100 630.450 100.200 631.050 ;
        RECT 106.950 630.450 109.050 631.050 ;
        RECT 98.100 629.400 109.050 630.450 ;
        RECT 98.100 628.950 100.200 629.400 ;
        RECT 106.950 628.950 109.050 629.400 ;
        RECT 115.950 628.050 118.050 631.050 ;
        RECT 121.950 628.950 124.050 632.400 ;
        RECT 133.950 631.950 136.050 632.400 ;
        RECT 139.950 631.050 142.050 634.050 ;
        RECT 146.400 633.450 147.450 635.400 ;
        RECT 181.950 635.400 208.050 636.000 ;
        RECT 181.950 634.050 184.050 635.400 ;
        RECT 205.950 634.950 208.050 635.400 ;
        RECT 172.950 633.450 175.050 634.050 ;
        RECT 146.400 632.400 175.050 633.450 ;
        RECT 127.950 630.450 130.050 631.050 ;
        RECT 136.800 630.450 138.900 631.050 ;
        RECT 127.950 629.400 138.900 630.450 ;
        RECT 139.950 630.000 142.200 631.050 ;
        RECT 127.950 628.950 130.050 629.400 ;
        RECT 136.800 628.950 138.900 629.400 ;
        RECT 140.100 628.950 142.200 630.000 ;
        RECT 157.950 628.950 160.050 632.400 ;
        RECT 172.950 631.950 175.050 632.400 ;
        RECT 181.800 633.000 184.050 634.050 ;
        RECT 185.100 633.450 187.200 634.050 ;
        RECT 244.950 633.450 247.050 634.050 ;
        RECT 181.800 631.950 183.900 633.000 ;
        RECT 185.100 632.400 247.050 633.450 ;
        RECT 185.100 631.950 187.200 632.400 ;
        RECT 244.950 631.950 247.050 632.400 ;
        RECT 253.950 633.450 256.050 634.050 ;
        RECT 259.950 633.450 262.050 634.050 ;
        RECT 253.950 632.400 262.050 633.450 ;
        RECT 253.950 631.950 256.050 632.400 ;
        RECT 259.950 631.950 262.050 632.400 ;
        RECT 265.950 631.950 270.900 634.050 ;
        RECT 272.100 631.950 277.050 634.050 ;
        RECT 304.950 631.950 307.050 637.050 ;
        RECT 334.950 636.450 337.050 637.050 ;
        RECT 361.950 636.450 364.050 637.050 ;
        RECT 334.950 635.400 364.050 636.450 ;
        RECT 334.950 634.950 337.050 635.400 ;
        RECT 361.950 634.950 364.050 635.400 ;
        RECT 382.950 636.450 385.050 637.050 ;
        RECT 451.950 636.450 454.050 637.050 ;
        RECT 499.950 636.450 502.050 637.050 ;
        RECT 382.950 635.400 423.450 636.450 ;
        RECT 382.950 634.950 385.050 635.400 ;
        RECT 310.950 631.050 313.050 634.050 ;
        RECT 316.950 633.450 319.050 634.050 ;
        RECT 316.950 632.400 345.450 633.450 ;
        RECT 347.100 633.000 349.200 634.050 ;
        RECT 395.100 633.000 397.200 634.050 ;
        RECT 316.950 631.950 319.050 632.400 ;
        RECT 344.400 631.050 345.450 632.400 ;
        RECT 346.950 631.950 349.200 633.000 ;
        RECT 394.950 631.950 397.200 633.000 ;
        RECT 346.950 631.050 349.050 631.950 ;
        RECT 394.950 631.050 397.050 631.950 ;
        RECT 175.950 628.950 181.050 631.050 ;
        RECT 184.950 630.450 187.050 631.050 ;
        RECT 193.950 630.450 196.050 631.050 ;
        RECT 184.950 629.400 196.050 630.450 ;
        RECT 184.950 628.950 187.050 629.400 ;
        RECT 193.950 628.950 196.050 629.400 ;
        RECT 202.950 630.450 205.050 631.050 ;
        RECT 202.950 629.400 219.450 630.450 ;
        RECT 202.950 628.950 205.050 629.400 ;
        RECT 85.950 627.450 88.050 628.050 ;
        RECT 73.950 627.000 88.050 627.450 ;
        RECT 74.400 626.400 88.050 627.000 ;
        RECT 16.800 624.000 18.900 625.050 ;
        RECT 20.100 624.450 22.200 625.050 ;
        RECT 38.400 624.450 39.450 626.400 ;
        RECT 85.950 625.950 88.050 626.400 ;
        RECT 94.950 625.950 99.900 628.050 ;
        RECT 101.100 625.950 106.050 628.050 ;
        RECT 109.950 625.950 114.900 628.050 ;
        RECT 115.800 627.000 118.050 628.050 ;
        RECT 115.800 625.950 117.900 627.000 ;
        RECT 119.100 625.950 123.900 628.050 ;
        RECT 125.100 627.450 127.200 628.050 ;
        RECT 139.950 627.450 142.050 628.050 ;
        RECT 151.950 627.450 154.050 628.050 ;
        RECT 184.950 627.450 187.050 628.050 ;
        RECT 125.100 626.400 187.050 627.450 ;
        RECT 218.400 627.450 219.450 629.400 ;
        RECT 223.950 628.950 229.050 631.050 ;
        RECT 232.950 628.950 238.050 631.050 ;
        RECT 250.950 628.950 255.900 631.050 ;
        RECT 257.100 630.000 259.200 631.050 ;
        RECT 256.950 628.950 259.200 630.000 ;
        RECT 265.950 628.950 270.900 631.050 ;
        RECT 272.100 630.450 274.200 631.050 ;
        RECT 283.950 630.450 288.900 631.050 ;
        RECT 272.100 629.400 288.900 630.450 ;
        RECT 272.100 628.950 274.200 629.400 ;
        RECT 283.950 628.950 288.900 629.400 ;
        RECT 290.100 628.950 295.050 631.050 ;
        RECT 298.950 630.450 301.050 631.050 ;
        RECT 307.800 630.450 309.900 631.050 ;
        RECT 298.950 629.400 309.900 630.450 ;
        RECT 310.950 630.000 313.200 631.050 ;
        RECT 298.950 628.950 301.050 629.400 ;
        RECT 307.800 628.950 309.900 629.400 ;
        RECT 311.100 628.950 313.200 630.000 ;
        RECT 322.950 628.950 328.050 631.050 ;
        RECT 331.950 628.950 337.050 631.050 ;
        RECT 343.800 630.000 345.900 631.050 ;
        RECT 346.950 630.000 349.200 631.050 ;
        RECT 343.800 628.950 346.050 630.000 ;
        RECT 347.100 628.950 349.200 630.000 ;
        RECT 352.950 630.450 355.050 631.050 ;
        RECT 358.950 630.450 361.050 631.050 ;
        RECT 352.950 629.400 361.050 630.450 ;
        RECT 352.950 628.950 355.050 629.400 ;
        RECT 358.950 628.950 361.050 629.400 ;
        RECT 370.950 630.450 373.050 631.050 ;
        RECT 385.950 630.450 391.050 631.050 ;
        RECT 370.950 629.400 391.050 630.450 ;
        RECT 394.950 630.000 397.200 631.050 ;
        RECT 370.950 628.950 373.050 629.400 ;
        RECT 385.950 628.950 391.050 629.400 ;
        RECT 395.100 628.950 397.200 630.000 ;
        RECT 406.950 630.450 409.050 631.050 ;
        RECT 412.950 630.450 415.050 631.050 ;
        RECT 406.950 629.400 415.050 630.450 ;
        RECT 406.950 628.950 409.050 629.400 ;
        RECT 412.950 628.950 415.050 629.400 ;
        RECT 229.950 627.450 232.050 628.050 ;
        RECT 218.400 626.400 232.050 627.450 ;
        RECT 125.100 625.950 127.200 626.400 ;
        RECT 139.950 625.950 142.050 626.400 ;
        RECT 151.950 625.950 154.050 626.400 ;
        RECT 184.950 625.950 187.050 626.400 ;
        RECT 229.950 625.950 232.050 626.400 ;
        RECT 235.950 627.450 241.050 628.050 ;
        RECT 256.950 627.450 259.050 628.950 ;
        RECT 235.950 627.000 259.050 627.450 ;
        RECT 259.950 627.450 262.050 628.050 ;
        RECT 289.950 627.450 292.050 628.050 ;
        RECT 235.950 626.400 258.600 627.000 ;
        RECT 259.950 626.400 292.050 627.450 ;
        RECT 235.950 625.950 241.050 626.400 ;
        RECT 259.950 625.950 262.050 626.400 ;
        RECT 289.950 625.950 292.050 626.400 ;
        RECT 295.950 627.450 298.050 628.050 ;
        RECT 316.800 627.450 318.900 628.050 ;
        RECT 295.950 626.400 318.900 627.450 ;
        RECT 295.950 625.950 298.050 626.400 ;
        RECT 316.800 625.950 318.900 626.400 ;
        RECT 320.100 627.450 322.200 628.050 ;
        RECT 328.950 627.450 331.050 628.050 ;
        RECT 320.100 626.400 331.050 627.450 ;
        RECT 320.100 625.950 322.200 626.400 ;
        RECT 328.950 625.950 331.050 626.400 ;
        RECT 334.950 625.950 340.050 628.050 ;
        RECT 343.950 625.950 346.050 628.950 ;
        RECT 418.950 628.050 421.050 631.050 ;
        RECT 422.400 630.450 423.450 635.400 ;
        RECT 451.950 635.400 502.050 636.450 ;
        RECT 451.950 634.950 454.050 635.400 ;
        RECT 470.400 634.050 471.450 635.400 ;
        RECT 499.950 634.950 502.050 635.400 ;
        RECT 514.950 636.450 517.050 637.050 ;
        RECT 538.950 636.450 541.050 637.050 ;
        RECT 514.950 635.400 541.050 636.450 ;
        RECT 514.950 634.950 517.050 635.400 ;
        RECT 538.950 634.950 541.050 635.400 ;
        RECT 439.950 633.450 442.050 634.050 ;
        RECT 451.950 633.450 454.050 634.050 ;
        RECT 439.950 632.400 454.050 633.450 ;
        RECT 439.950 631.950 442.050 632.400 ;
        RECT 451.950 631.950 454.050 632.400 ;
        RECT 457.950 633.450 460.050 634.050 ;
        RECT 469.950 633.450 472.050 634.050 ;
        RECT 457.950 632.400 472.050 633.450 ;
        RECT 457.950 631.950 460.050 632.400 ;
        RECT 469.950 631.950 472.050 632.400 ;
        RECT 478.950 633.450 481.050 634.050 ;
        RECT 478.950 633.000 498.600 633.450 ;
        RECT 478.950 632.400 499.050 633.000 ;
        RECT 478.950 631.950 481.050 632.400 ;
        RECT 496.950 631.050 499.050 632.400 ;
        RECT 442.950 630.450 445.050 631.050 ;
        RECT 422.400 630.000 445.050 630.450 ;
        RECT 16.800 622.950 19.050 624.000 ;
        RECT 20.100 623.400 39.450 624.450 ;
        RECT 20.100 622.950 22.200 623.400 ;
        RECT 199.950 622.950 205.050 625.050 ;
        RECT 214.950 624.450 217.050 625.050 ;
        RECT 235.950 624.450 238.050 625.050 ;
        RECT 214.950 623.400 238.050 624.450 ;
        RECT 214.950 622.950 217.050 623.400 ;
        RECT 235.950 622.950 238.050 623.400 ;
        RECT 241.950 624.450 244.050 625.200 ;
        RECT 271.950 624.450 274.050 625.050 ;
        RECT 241.950 623.400 274.050 624.450 ;
        RECT 338.400 624.450 339.450 625.950 ;
        RECT 346.950 624.450 349.050 625.050 ;
        RECT 338.400 623.400 349.050 624.450 ;
        RECT 349.950 624.450 352.050 628.050 ;
        RECT 355.950 627.450 358.050 628.050 ;
        RECT 364.950 627.450 367.050 628.050 ;
        RECT 355.950 626.400 367.050 627.450 ;
        RECT 355.950 625.950 358.050 626.400 ;
        RECT 364.950 625.950 367.050 626.400 ;
        RECT 376.950 627.450 379.050 628.050 ;
        RECT 382.950 627.450 388.050 628.050 ;
        RECT 390.000 627.450 394.050 628.050 ;
        RECT 376.950 626.400 388.050 627.450 ;
        RECT 376.950 625.950 379.050 626.400 ;
        RECT 382.950 625.950 388.050 626.400 ;
        RECT 389.400 625.950 394.050 627.450 ;
        RECT 397.950 625.950 402.900 628.050 ;
        RECT 404.100 627.450 406.200 628.050 ;
        RECT 409.800 627.450 411.900 628.050 ;
        RECT 404.100 626.400 411.900 627.450 ;
        RECT 404.100 625.950 406.200 626.400 ;
        RECT 409.800 625.950 411.900 626.400 ;
        RECT 413.100 625.950 417.900 628.050 ;
        RECT 418.800 627.000 421.050 628.050 ;
        RECT 421.950 629.400 445.050 630.000 ;
        RECT 421.950 628.050 424.050 629.400 ;
        RECT 442.950 628.950 445.050 629.400 ;
        RECT 448.950 630.450 451.050 631.050 ;
        RECT 454.950 630.450 457.050 631.050 ;
        RECT 448.950 629.400 457.050 630.450 ;
        RECT 448.950 628.950 451.050 629.400 ;
        RECT 454.950 628.950 457.050 629.400 ;
        RECT 472.950 628.950 478.050 631.050 ;
        RECT 487.950 628.950 492.900 631.050 ;
        RECT 494.100 630.000 496.200 631.050 ;
        RECT 496.950 630.000 499.200 631.050 ;
        RECT 493.950 628.950 496.200 630.000 ;
        RECT 497.100 628.950 499.200 630.000 ;
        RECT 511.950 628.950 514.050 634.050 ;
        RECT 535.950 633.450 538.050 634.200 ;
        RECT 547.950 633.450 550.050 634.050 ;
        RECT 535.950 632.400 550.050 633.450 ;
        RECT 535.950 632.100 538.050 632.400 ;
        RECT 547.950 631.950 550.050 632.400 ;
        RECT 517.950 630.450 520.050 631.050 ;
        RECT 529.950 630.450 532.050 631.050 ;
        RECT 517.950 629.400 532.050 630.450 ;
        RECT 517.950 628.950 520.050 629.400 ;
        RECT 529.950 628.950 532.050 629.400 ;
        RECT 535.950 630.450 538.050 630.900 ;
        RECT 550.950 630.450 553.050 631.050 ;
        RECT 535.950 629.400 553.050 630.450 ;
        RECT 553.950 630.450 556.050 634.050 ;
        RECT 562.950 631.950 565.050 637.050 ;
        RECT 568.950 631.950 574.050 634.050 ;
        RECT 577.950 633.450 580.050 634.050 ;
        RECT 583.950 633.450 586.050 634.050 ;
        RECT 577.950 632.400 586.050 633.450 ;
        RECT 577.950 631.950 580.050 632.400 ;
        RECT 583.950 631.950 586.050 632.400 ;
        RECT 589.950 633.450 595.050 634.050 ;
        RECT 616.950 633.450 619.050 634.050 ;
        RECT 589.950 632.400 619.050 633.450 ;
        RECT 589.950 631.950 595.050 632.400 ;
        RECT 616.950 631.950 619.050 632.400 ;
        RECT 625.950 633.450 628.050 634.050 ;
        RECT 631.950 633.450 634.050 634.050 ;
        RECT 625.950 632.400 634.050 633.450 ;
        RECT 625.950 631.950 628.050 632.400 ;
        RECT 631.950 631.950 634.050 632.400 ;
        RECT 637.950 631.950 640.050 637.050 ;
        RECT 671.850 635.700 673.050 639.300 ;
        RECT 691.950 638.400 694.050 640.500 ;
        RECT 724.950 638.400 727.050 640.500 ;
        RECT 745.950 639.300 748.050 641.400 ;
        RECT 781.950 639.450 784.050 640.050 ;
        RECT 805.950 639.450 808.050 640.050 ;
        RECT 643.950 633.450 646.050 634.050 ;
        RECT 670.950 633.600 673.050 635.700 ;
        RECT 643.950 633.000 660.300 633.450 ;
        RECT 643.950 632.400 661.050 633.000 ;
        RECT 643.950 631.950 646.050 632.400 ;
        RECT 658.950 631.050 661.050 632.400 ;
        RECT 565.950 630.450 568.050 631.050 ;
        RECT 553.950 630.000 568.050 630.450 ;
        RECT 554.400 629.400 568.050 630.000 ;
        RECT 493.950 628.050 496.050 628.950 ;
        RECT 535.950 628.800 538.050 629.400 ;
        RECT 550.950 628.950 553.050 629.400 ;
        RECT 565.950 628.950 568.050 629.400 ;
        RECT 421.950 627.000 424.200 628.050 ;
        RECT 418.800 625.950 420.900 627.000 ;
        RECT 422.100 625.950 424.200 627.000 ;
        RECT 478.950 627.450 481.050 628.050 ;
        RECT 484.950 627.450 487.050 628.050 ;
        RECT 478.950 626.400 487.050 627.450 ;
        RECT 493.950 627.000 496.200 628.050 ;
        RECT 478.950 625.950 481.050 626.400 ;
        RECT 484.950 625.950 487.050 626.400 ;
        RECT 494.100 625.950 496.200 627.000 ;
        RECT 361.950 624.450 364.050 625.050 ;
        RECT 349.950 624.000 364.050 624.450 ;
        RECT 350.400 623.400 364.050 624.000 ;
        RECT 241.950 623.100 244.050 623.400 ;
        RECT 271.950 622.950 274.050 623.400 ;
        RECT 346.950 622.950 349.050 623.400 ;
        RECT 361.950 622.950 364.050 623.400 ;
        RECT 376.950 624.450 379.050 625.050 ;
        RECT 389.400 624.450 390.450 625.950 ;
        RECT 376.950 623.400 390.450 624.450 ;
        RECT 391.950 624.450 394.050 625.050 ;
        RECT 406.950 624.450 409.050 625.050 ;
        RECT 391.950 623.400 409.050 624.450 ;
        RECT 376.950 622.950 379.050 623.400 ;
        RECT 391.950 622.950 394.050 623.400 ;
        RECT 406.950 622.950 409.050 623.400 ;
        RECT 430.950 622.950 436.050 625.050 ;
        RECT 457.950 624.450 460.050 625.050 ;
        RECT 484.950 624.450 487.050 625.050 ;
        RECT 457.950 623.400 487.050 624.450 ;
        RECT 457.950 622.950 460.050 623.400 ;
        RECT 484.950 622.950 487.050 623.400 ;
        RECT 499.950 622.950 502.050 628.050 ;
        RECT 505.950 625.950 510.900 628.050 ;
        RECT 512.100 625.950 517.050 628.050 ;
        RECT 523.950 624.450 526.050 625.050 ;
        RECT 535.950 624.450 538.050 628.050 ;
        RECT 586.950 625.950 589.050 631.050 ;
        RECT 598.950 628.950 604.050 631.050 ;
        RECT 613.950 625.950 619.050 628.050 ;
        RECT 634.950 627.450 637.050 631.050 ;
        RECT 652.800 630.000 654.900 631.050 ;
        RECT 655.800 630.000 657.900 631.050 ;
        RECT 658.800 630.000 661.050 631.050 ;
        RECT 662.100 630.000 664.200 631.050 ;
        RECT 652.800 628.950 655.050 630.000 ;
        RECT 655.800 628.950 658.050 630.000 ;
        RECT 658.800 628.950 660.900 630.000 ;
        RECT 661.950 628.950 664.200 630.000 ;
        RECT 652.950 627.450 655.050 628.950 ;
        RECT 634.950 627.000 655.050 627.450 ;
        RECT 635.400 626.400 654.300 627.000 ;
        RECT 655.950 625.950 658.050 628.950 ;
        RECT 661.950 625.950 664.050 628.950 ;
        RECT 541.950 624.450 544.050 625.050 ;
        RECT 523.950 623.400 544.050 624.450 ;
        RECT 523.950 622.950 526.050 623.400 ;
        RECT 535.950 622.950 538.050 623.400 ;
        RECT 541.950 622.950 544.050 623.400 ;
        RECT 586.950 624.450 589.050 625.050 ;
        RECT 598.950 624.450 601.050 625.050 ;
        RECT 586.950 623.400 601.050 624.450 ;
        RECT 617.400 624.450 618.450 625.950 ;
        RECT 667.950 624.450 670.050 628.050 ;
        RECT 617.400 624.000 670.050 624.450 ;
        RECT 617.400 623.400 669.450 624.000 ;
        RECT 586.950 622.950 589.050 623.400 ;
        RECT 598.950 622.950 601.050 623.400 ;
        RECT 16.950 621.450 19.050 622.950 ;
        RECT 40.950 621.450 43.050 622.050 ;
        RECT 16.950 621.000 43.050 621.450 ;
        RECT 17.250 620.400 43.050 621.000 ;
        RECT 40.950 619.950 43.050 620.400 ;
        RECT 79.950 618.450 82.050 622.050 ;
        RECT 94.950 621.450 97.050 622.050 ;
        RECT 115.950 621.450 118.050 622.050 ;
        RECT 130.950 621.450 133.050 622.050 ;
        RECT 243.000 621.900 247.050 622.050 ;
        RECT 94.950 620.400 133.050 621.450 ;
        RECT 94.950 619.950 97.050 620.400 ;
        RECT 115.950 619.950 118.050 620.400 ;
        RECT 130.950 619.950 133.050 620.400 ;
        RECT 241.950 619.950 247.050 621.900 ;
        RECT 250.950 621.450 253.050 622.050 ;
        RECT 319.950 621.450 322.050 622.050 ;
        RECT 250.950 620.400 322.050 621.450 ;
        RECT 250.950 619.950 253.050 620.400 ;
        RECT 319.950 619.950 322.050 620.400 ;
        RECT 352.950 621.450 355.050 622.050 ;
        RECT 373.950 621.450 376.050 622.050 ;
        RECT 352.950 620.400 376.050 621.450 ;
        RECT 352.950 619.950 355.050 620.400 ;
        RECT 373.950 619.950 376.050 620.400 ;
        RECT 382.950 621.450 385.050 622.050 ;
        RECT 403.950 621.450 406.050 622.050 ;
        RECT 382.950 620.400 406.050 621.450 ;
        RECT 382.950 619.950 385.050 620.400 ;
        RECT 403.950 619.950 406.050 620.400 ;
        RECT 493.950 621.450 496.050 622.050 ;
        RECT 505.950 621.450 508.050 622.050 ;
        RECT 493.950 620.400 508.050 621.450 ;
        RECT 493.950 619.950 496.050 620.400 ;
        RECT 505.950 619.950 508.050 620.400 ;
        RECT 580.950 621.450 583.050 622.050 ;
        RECT 601.950 621.450 604.050 622.050 ;
        RECT 580.950 620.400 604.050 621.450 ;
        RECT 580.950 619.950 583.050 620.400 ;
        RECT 601.950 619.950 604.050 620.400 ;
        RECT 607.950 621.450 610.050 622.050 ;
        RECT 613.950 621.450 616.050 622.050 ;
        RECT 607.950 620.400 616.050 621.450 ;
        RECT 607.950 619.950 610.050 620.400 ;
        RECT 613.950 619.950 616.050 620.400 ;
        RECT 661.950 619.950 664.050 622.050 ;
        RECT 671.850 621.600 673.050 633.600 ;
        RECT 682.950 628.950 688.050 631.050 ;
        RECT 676.950 625.950 682.050 628.050 ;
        RECT 692.100 621.600 693.300 638.400 ;
        RECT 694.950 636.450 697.050 637.050 ;
        RECT 718.950 636.450 721.050 637.050 ;
        RECT 694.950 635.400 721.050 636.450 ;
        RECT 694.950 634.950 697.050 635.400 ;
        RECT 718.950 634.950 721.050 635.400 ;
        RECT 700.950 627.450 703.050 628.050 ;
        RECT 706.800 627.450 708.900 628.050 ;
        RECT 700.950 626.400 708.900 627.450 ;
        RECT 700.950 625.950 703.050 626.400 ;
        RECT 706.800 625.950 708.900 626.400 ;
        RECT 710.100 627.450 712.200 628.050 ;
        RECT 715.950 627.450 718.050 628.050 ;
        RECT 710.100 626.400 718.050 627.450 ;
        RECT 710.100 625.950 712.200 626.400 ;
        RECT 715.950 625.950 718.050 626.400 ;
        RECT 725.700 621.600 726.900 638.400 ;
        RECT 745.950 635.700 747.150 639.300 ;
        RECT 781.950 638.400 808.050 639.450 ;
        RECT 781.950 637.950 784.050 638.400 ;
        RECT 805.950 637.950 808.050 638.400 ;
        RECT 769.950 636.450 772.050 637.050 ;
        RECT 787.950 636.450 790.050 637.050 ;
        RECT 745.950 633.600 748.050 635.700 ;
        RECT 769.950 635.400 790.050 636.450 ;
        RECT 769.950 634.950 772.050 635.400 ;
        RECT 787.950 634.950 790.050 635.400 ;
        RECT 730.950 622.950 733.050 628.050 ;
        RECT 736.950 622.950 739.050 628.050 ;
        RECT 745.950 621.600 747.150 633.600 ;
        RECT 781.950 628.950 784.050 634.050 ;
        RECT 793.950 633.450 796.050 634.050 ;
        RECT 799.950 633.450 802.050 634.050 ;
        RECT 793.950 632.400 802.050 633.450 ;
        RECT 793.950 631.950 796.050 632.400 ;
        RECT 799.950 631.950 802.050 632.400 ;
        RECT 805.950 633.450 808.050 637.050 ;
        RECT 817.950 633.450 823.050 634.050 ;
        RECT 805.950 632.400 823.050 633.450 ;
        RECT 805.950 631.950 808.050 632.400 ;
        RECT 817.950 631.950 823.050 632.400 ;
        RECT 826.950 631.050 829.050 634.050 ;
        RECT 787.950 630.450 790.050 631.050 ;
        RECT 802.950 630.450 805.050 631.050 ;
        RECT 787.950 629.400 805.050 630.450 ;
        RECT 787.950 628.950 790.050 629.400 ;
        RECT 802.950 628.950 805.050 629.400 ;
        RECT 820.950 628.950 825.900 631.050 ;
        RECT 826.950 630.000 829.200 631.050 ;
        RECT 827.100 628.950 829.200 630.000 ;
        RECT 832.950 630.450 835.050 631.050 ;
        RECT 838.950 630.450 841.050 631.050 ;
        RECT 832.950 629.400 841.050 630.450 ;
        RECT 832.950 628.950 835.050 629.400 ;
        RECT 838.950 628.950 841.050 629.400 ;
        RECT 844.950 628.950 850.050 631.050 ;
        RECT 748.950 625.950 753.900 628.050 ;
        RECT 755.100 627.450 757.200 628.050 ;
        RECT 760.950 627.450 763.050 628.050 ;
        RECT 755.100 626.400 763.050 627.450 ;
        RECT 755.100 625.950 757.200 626.400 ;
        RECT 760.950 625.950 763.050 626.400 ;
        RECT 769.950 625.950 774.900 628.050 ;
        RECT 776.100 625.950 781.050 628.050 ;
        RECT 784.950 622.950 787.050 628.050 ;
        RECT 814.950 624.450 817.050 625.050 ;
        RECT 823.950 624.450 826.050 625.050 ;
        RECT 814.950 623.400 826.050 624.450 ;
        RECT 814.950 622.950 817.050 623.400 ;
        RECT 823.950 622.950 826.050 623.400 ;
        RECT 835.950 622.950 838.050 628.050 ;
        RECT 841.950 625.050 844.050 628.050 ;
        RECT 841.950 624.000 847.050 625.050 ;
        RECT 842.400 623.400 847.050 624.000 ;
        RECT 843.000 622.950 847.050 623.400 ;
        RECT 241.950 619.800 244.050 619.950 ;
        RECT 85.950 618.450 88.050 619.050 ;
        RECT 79.950 618.000 88.050 618.450 ;
        RECT 80.400 617.400 88.050 618.000 ;
        RECT 85.950 616.950 88.050 617.400 ;
        RECT 106.950 616.950 112.050 619.050 ;
        RECT 175.950 618.450 178.050 619.050 ;
        RECT 226.950 618.450 229.050 619.050 ;
        RECT 265.950 618.450 268.050 619.050 ;
        RECT 175.950 617.400 268.050 618.450 ;
        RECT 175.950 616.950 178.050 617.400 ;
        RECT 226.950 616.950 229.050 617.400 ;
        RECT 265.950 616.950 268.050 617.400 ;
        RECT 319.950 618.450 322.050 619.050 ;
        RECT 334.950 618.450 337.050 619.050 ;
        RECT 370.950 618.450 373.050 619.050 ;
        RECT 442.950 618.450 445.050 619.050 ;
        RECT 319.950 617.400 445.050 618.450 ;
        RECT 319.950 616.950 322.050 617.400 ;
        RECT 334.950 616.950 337.050 617.400 ;
        RECT 370.950 616.950 373.050 617.400 ;
        RECT 442.950 616.950 445.050 617.400 ;
        RECT 649.950 618.450 652.050 619.050 ;
        RECT 658.950 618.450 661.050 619.050 ;
        RECT 649.950 617.400 661.050 618.450 ;
        RECT 649.950 616.950 652.050 617.400 ;
        RECT 658.950 616.950 661.050 617.400 ;
        RECT 40.950 615.450 43.050 616.050 ;
        RECT 88.950 615.450 91.050 616.050 ;
        RECT 40.950 614.400 91.050 615.450 ;
        RECT 40.950 613.950 43.050 614.400 ;
        RECT 88.950 613.950 91.050 614.400 ;
        RECT 202.950 615.450 205.050 616.050 ;
        RECT 238.950 615.450 241.050 616.050 ;
        RECT 298.950 615.450 301.050 616.050 ;
        RECT 202.950 614.400 301.050 615.450 ;
        RECT 202.950 613.950 205.050 614.400 ;
        RECT 238.950 613.950 241.050 614.400 ;
        RECT 298.950 613.950 301.050 614.400 ;
        RECT 310.950 615.450 313.050 616.050 ;
        RECT 316.950 615.450 319.050 616.050 ;
        RECT 310.950 614.400 319.050 615.450 ;
        RECT 310.950 613.950 313.050 614.400 ;
        RECT 316.950 613.950 319.050 614.400 ;
        RECT 379.950 615.450 382.050 616.050 ;
        RECT 388.950 615.450 391.050 616.050 ;
        RECT 379.950 614.400 391.050 615.450 ;
        RECT 379.950 613.950 382.050 614.400 ;
        RECT 388.950 613.950 391.050 614.400 ;
        RECT 484.950 615.450 487.050 616.050 ;
        RECT 511.950 615.450 514.050 616.050 ;
        RECT 484.950 614.400 514.050 615.450 ;
        RECT 484.950 613.950 487.050 614.400 ;
        RECT 511.950 613.950 514.050 614.400 ;
        RECT 583.950 615.450 586.050 616.050 ;
        RECT 610.950 615.450 613.050 616.050 ;
        RECT 583.950 614.400 613.050 615.450 ;
        RECT 583.950 613.950 586.050 614.400 ;
        RECT 610.950 613.950 613.050 614.400 ;
        RECT 622.950 615.450 625.050 616.050 ;
        RECT 628.950 615.450 631.050 615.900 ;
        RECT 622.950 614.400 631.050 615.450 ;
        RECT 662.400 615.450 663.450 619.950 ;
        RECT 670.950 619.500 673.050 621.600 ;
        RECT 691.950 619.500 694.050 621.600 ;
        RECT 724.950 619.500 727.050 621.600 ;
        RECT 745.950 619.500 748.050 621.600 ;
        RECT 817.950 618.450 820.050 619.050 ;
        RECT 841.950 618.450 844.050 619.050 ;
        RECT 817.950 617.400 844.050 618.450 ;
        RECT 817.950 616.950 820.050 617.400 ;
        RECT 841.950 616.950 844.050 617.400 ;
        RECT 727.950 615.450 730.050 616.050 ;
        RECT 662.400 614.400 730.050 615.450 ;
        RECT 622.950 613.950 625.050 614.400 ;
        RECT 628.950 613.800 631.050 614.400 ;
        RECT 727.950 613.950 730.050 614.400 ;
        RECT 49.950 612.450 52.050 613.050 ;
        RECT 79.950 612.450 82.050 613.050 ;
        RECT 49.950 611.400 82.050 612.450 ;
        RECT 49.950 610.950 52.050 611.400 ;
        RECT 79.950 610.950 82.050 611.400 ;
        RECT 307.950 612.450 310.050 613.050 ;
        RECT 343.950 612.450 346.050 613.050 ;
        RECT 307.950 611.400 346.050 612.450 ;
        RECT 307.950 610.950 310.050 611.400 ;
        RECT 343.950 610.950 346.050 611.400 ;
        RECT 364.950 612.450 367.050 613.050 ;
        RECT 391.950 612.450 394.050 613.050 ;
        RECT 364.950 611.400 394.050 612.450 ;
        RECT 364.950 610.950 367.050 611.400 ;
        RECT 391.950 610.950 394.050 611.400 ;
        RECT 445.950 612.450 448.050 613.050 ;
        RECT 478.950 612.450 481.050 613.050 ;
        RECT 556.950 612.450 559.050 613.050 ;
        RECT 445.950 611.400 559.050 612.450 ;
        RECT 445.950 610.950 448.050 611.400 ;
        RECT 478.950 610.950 481.050 611.400 ;
        RECT 556.950 610.950 559.050 611.400 ;
        RECT 709.950 612.450 712.050 613.050 ;
        RECT 754.950 612.450 757.050 613.050 ;
        RECT 709.950 611.400 757.050 612.450 ;
        RECT 709.950 610.950 712.050 611.400 ;
        RECT 754.950 610.950 757.050 611.400 ;
        RECT 16.950 609.450 19.050 610.050 ;
        RECT 52.950 609.450 55.050 610.050 ;
        RECT 67.950 609.450 70.050 610.050 ;
        RECT 16.950 608.400 70.050 609.450 ;
        RECT 16.950 607.950 19.050 608.400 ;
        RECT 52.950 607.950 55.050 608.400 ;
        RECT 67.950 607.950 70.050 608.400 ;
        RECT 103.950 609.450 106.050 610.050 ;
        RECT 127.950 609.450 130.050 610.050 ;
        RECT 103.950 608.400 130.050 609.450 ;
        RECT 103.950 607.950 106.050 608.400 ;
        RECT 127.950 607.950 130.050 608.400 ;
        RECT 196.950 609.450 199.050 610.050 ;
        RECT 295.950 609.450 298.050 610.050 ;
        RECT 196.950 608.400 298.050 609.450 ;
        RECT 196.950 607.950 199.050 608.400 ;
        RECT 295.950 607.950 298.050 608.400 ;
        RECT 313.950 609.450 316.050 610.050 ;
        RECT 337.950 609.450 340.050 610.050 ;
        RECT 397.950 609.450 400.050 610.050 ;
        RECT 418.950 609.450 421.050 610.050 ;
        RECT 313.950 608.400 421.050 609.450 ;
        RECT 313.950 607.950 316.050 608.400 ;
        RECT 337.950 607.950 340.050 608.400 ;
        RECT 397.950 607.950 400.050 608.400 ;
        RECT 418.950 607.950 421.050 608.400 ;
        RECT 499.950 609.450 502.050 610.050 ;
        RECT 511.950 609.450 514.050 610.050 ;
        RECT 499.950 608.400 514.050 609.450 ;
        RECT 499.950 607.950 502.050 608.400 ;
        RECT 511.950 607.950 514.050 608.400 ;
        RECT 643.950 609.450 646.050 610.050 ;
        RECT 679.950 609.450 682.050 610.050 ;
        RECT 712.950 609.450 715.050 610.050 ;
        RECT 736.950 609.450 739.050 610.050 ;
        RECT 643.950 608.400 739.050 609.450 ;
        RECT 643.950 607.950 646.050 608.400 ;
        RECT 679.950 607.950 682.050 608.400 ;
        RECT 712.950 607.950 715.050 608.400 ;
        RECT 736.950 607.950 739.050 608.400 ;
        RECT 745.950 609.450 748.050 610.050 ;
        RECT 772.950 609.450 775.050 610.050 ;
        RECT 745.950 608.400 775.050 609.450 ;
        RECT 745.950 607.950 748.050 608.400 ;
        RECT 772.950 607.950 775.050 608.400 ;
        RECT 781.950 609.450 784.050 610.050 ;
        RECT 844.800 609.450 846.900 610.050 ;
        RECT 781.950 608.400 846.900 609.450 ;
        RECT 781.950 607.950 784.050 608.400 ;
        RECT 844.800 607.950 846.900 608.400 ;
        RECT 848.100 607.950 853.050 610.050 ;
        RECT 244.950 607.050 247.050 607.200 ;
        RECT 25.950 606.450 28.050 607.050 ;
        RECT 49.950 606.450 52.050 607.050 ;
        RECT 25.950 605.400 52.050 606.450 ;
        RECT 25.950 604.950 28.050 605.400 ;
        RECT 49.950 604.950 52.050 605.400 ;
        RECT 58.950 606.450 61.050 607.050 ;
        RECT 103.950 606.450 106.050 607.050 ;
        RECT 58.950 605.400 106.050 606.450 ;
        RECT 58.950 604.950 61.050 605.400 ;
        RECT 103.950 604.950 106.050 605.400 ;
        RECT 109.950 606.450 114.000 607.050 ;
        RECT 109.950 606.000 114.450 606.450 ;
        RECT 109.950 604.950 115.050 606.000 ;
        RECT 241.950 605.100 247.050 607.050 ;
        RECT 310.950 606.450 313.050 607.050 ;
        RECT 331.950 606.450 334.050 607.050 ;
        RECT 373.950 606.450 376.050 607.050 ;
        RECT 490.950 606.450 493.050 607.050 ;
        RECT 310.950 605.400 330.450 606.450 ;
        RECT 241.950 604.950 246.000 605.100 ;
        RECT 310.950 604.950 313.050 605.400 ;
        RECT 16.950 603.450 19.050 604.050 ;
        RECT 16.950 603.000 33.600 603.450 ;
        RECT 16.950 602.400 34.050 603.000 ;
        RECT 16.950 601.950 19.050 602.400 ;
        RECT 31.950 601.050 34.050 602.400 ;
        RECT 112.950 601.950 115.050 604.950 ;
        RECT 169.950 603.450 172.050 604.050 ;
        RECT 184.950 603.450 187.050 604.050 ;
        RECT 169.950 602.400 187.050 603.450 ;
        RECT 169.950 601.950 172.050 602.400 ;
        RECT 184.950 601.950 187.050 602.400 ;
        RECT 205.950 603.450 208.050 604.050 ;
        RECT 246.000 603.900 250.050 604.050 ;
        RECT 205.950 603.000 228.300 603.450 ;
        RECT 205.950 602.400 229.050 603.000 ;
        RECT 205.950 601.950 208.050 602.400 ;
        RECT 226.950 601.050 229.050 602.400 ;
        RECT 244.950 601.950 250.050 603.900 ;
        RECT 244.950 601.800 247.050 601.950 ;
        RECT 28.800 600.450 30.900 601.050 ;
        RECT 14.400 600.000 30.900 600.450 ;
        RECT 31.950 600.000 34.200 601.050 ;
        RECT 13.950 599.400 30.900 600.000 ;
        RECT 13.950 595.950 16.050 599.400 ;
        RECT 28.800 598.950 30.900 599.400 ;
        RECT 32.100 598.950 34.200 600.000 ;
        RECT 40.950 600.450 43.050 601.050 ;
        RECT 40.950 599.400 69.450 600.450 ;
        RECT 40.950 598.950 43.050 599.400 ;
        RECT 19.950 597.450 22.050 598.050 ;
        RECT 25.950 597.450 31.050 598.050 ;
        RECT 19.950 596.400 31.050 597.450 ;
        RECT 19.950 595.950 22.050 596.400 ;
        RECT 25.950 595.950 31.050 596.400 ;
        RECT 34.950 595.950 37.050 598.050 ;
        RECT 46.950 595.950 52.050 598.050 ;
        RECT 55.950 597.450 60.000 598.050 ;
        RECT 68.400 597.450 69.450 599.400 ;
        RECT 70.950 598.950 75.900 601.050 ;
        RECT 77.100 598.950 82.050 601.050 ;
        RECT 88.950 600.450 91.050 601.050 ;
        RECT 103.950 600.450 106.050 601.050 ;
        RECT 109.950 600.450 112.050 601.050 ;
        RECT 88.950 600.000 96.450 600.450 ;
        RECT 88.950 599.400 97.050 600.000 ;
        RECT 88.950 598.950 91.050 599.400 ;
        RECT 94.950 598.050 97.050 599.400 ;
        RECT 103.950 599.400 112.050 600.450 ;
        RECT 103.950 598.950 106.050 599.400 ;
        RECT 109.950 598.950 112.050 599.400 ;
        RECT 73.950 597.450 76.050 598.050 ;
        RECT 55.950 595.950 60.450 597.450 ;
        RECT 68.400 596.400 76.050 597.450 ;
        RECT 73.950 595.950 76.050 596.400 ;
        RECT 7.950 592.950 13.050 595.050 ;
        RECT 16.950 589.950 19.050 595.050 ;
        RECT 22.950 591.450 25.050 592.050 ;
        RECT 35.400 591.450 36.450 595.950 ;
        RECT 52.950 592.950 58.050 595.050 ;
        RECT 59.400 591.450 60.450 595.950 ;
        RECT 61.950 594.450 66.000 595.050 ;
        RECT 61.950 592.950 66.450 594.450 ;
        RECT 79.950 592.950 82.050 598.050 ;
        RECT 91.800 597.000 93.900 598.050 ;
        RECT 94.950 597.000 97.200 598.050 ;
        RECT 115.950 597.450 118.050 601.050 ;
        RECT 91.800 595.950 94.050 597.000 ;
        RECT 95.100 595.950 97.200 597.000 ;
        RECT 104.400 597.000 118.050 597.450 ;
        RECT 104.400 596.400 117.450 597.000 ;
        RECT 91.950 592.950 94.050 595.950 ;
        RECT 104.400 595.050 105.450 596.400 ;
        RECT 130.950 595.950 133.050 601.050 ;
        RECT 160.950 600.450 163.050 601.050 ;
        RECT 187.950 600.450 190.050 601.050 ;
        RECT 160.950 599.400 190.050 600.450 ;
        RECT 160.950 598.950 163.050 599.400 ;
        RECT 187.950 598.950 190.050 599.400 ;
        RECT 196.950 600.450 199.050 601.050 ;
        RECT 202.950 600.450 205.050 601.050 ;
        RECT 196.950 599.400 205.050 600.450 ;
        RECT 196.950 598.950 199.050 599.400 ;
        RECT 202.950 598.950 205.050 599.400 ;
        RECT 211.950 598.950 217.050 601.050 ;
        RECT 226.800 600.000 229.050 601.050 ;
        RECT 226.800 598.950 228.900 600.000 ;
        RECT 230.100 598.950 234.900 601.050 ;
        RECT 236.100 600.450 238.200 601.050 ;
        RECT 236.100 599.400 252.450 600.450 ;
        RECT 236.100 598.950 238.200 599.400 ;
        RECT 136.950 597.450 139.050 598.050 ;
        RECT 151.950 597.450 154.050 598.050 ;
        RECT 136.950 596.400 154.050 597.450 ;
        RECT 161.400 597.450 162.450 598.950 ;
        RECT 161.400 596.400 165.450 597.450 ;
        RECT 136.950 595.950 139.050 596.400 ;
        RECT 151.950 595.950 154.050 596.400 ;
        RECT 97.950 594.450 100.050 595.050 ;
        RECT 103.950 594.450 106.050 595.050 ;
        RECT 97.950 593.400 106.050 594.450 ;
        RECT 97.950 592.950 100.050 593.400 ;
        RECT 103.950 592.950 106.050 593.400 ;
        RECT 127.950 594.900 132.000 595.050 ;
        RECT 127.950 592.950 132.900 594.900 ;
        RECT 134.100 594.000 136.200 595.050 ;
        RECT 22.950 590.400 60.450 591.450 ;
        RECT 65.400 591.450 66.450 592.950 ;
        RECT 79.950 591.450 82.050 592.050 ;
        RECT 65.400 590.400 82.050 591.450 ;
        RECT 104.400 591.450 105.450 592.950 ;
        RECT 130.800 592.800 132.900 592.950 ;
        RECT 133.950 592.950 136.200 594.000 ;
        RECT 133.950 591.450 136.050 592.950 ;
        RECT 104.400 591.000 136.050 591.450 ;
        RECT 104.400 590.400 135.600 591.000 ;
        RECT 22.950 589.950 25.050 590.400 ;
        RECT 79.950 589.950 82.050 590.400 ;
        RECT 148.950 589.950 151.050 595.050 ;
        RECT 154.950 589.950 157.050 595.050 ;
        RECT 164.400 594.450 165.450 596.400 ;
        RECT 166.950 595.950 171.900 598.050 ;
        RECT 173.100 597.450 178.050 598.050 ;
        RECT 184.950 597.450 187.050 598.050 ;
        RECT 173.100 596.400 187.050 597.450 ;
        RECT 173.100 595.950 178.050 596.400 ;
        RECT 184.950 595.950 187.050 596.400 ;
        RECT 172.950 594.450 175.050 595.050 ;
        RECT 164.400 593.400 175.050 594.450 ;
        RECT 172.950 592.950 175.050 593.400 ;
        RECT 190.950 592.950 193.050 598.050 ;
        RECT 211.950 592.950 214.050 598.050 ;
        RECT 215.400 594.450 216.450 598.950 ;
        RECT 217.950 595.950 223.050 598.050 ;
        RECT 229.950 595.950 234.900 598.050 ;
        RECT 236.100 597.450 238.200 598.050 ;
        RECT 247.950 597.450 250.050 598.050 ;
        RECT 236.100 596.400 250.050 597.450 ;
        RECT 251.400 597.450 252.450 599.400 ;
        RECT 280.950 598.950 286.050 601.050 ;
        RECT 292.950 600.450 295.050 601.050 ;
        RECT 313.950 600.450 316.050 601.050 ;
        RECT 319.950 600.450 322.050 601.050 ;
        RECT 292.950 599.400 322.050 600.450 ;
        RECT 292.950 598.950 295.050 599.400 ;
        RECT 265.950 597.450 268.050 598.050 ;
        RECT 251.400 596.400 268.050 597.450 ;
        RECT 236.100 595.950 238.200 596.400 ;
        RECT 247.950 595.950 250.050 596.400 ;
        RECT 265.950 595.950 268.050 596.400 ;
        RECT 229.950 594.450 232.050 595.050 ;
        RECT 215.400 593.400 232.050 594.450 ;
        RECT 229.950 592.950 232.050 593.400 ;
        RECT 238.950 594.450 244.050 595.050 ;
        RECT 262.800 594.450 264.900 595.050 ;
        RECT 238.950 593.400 264.900 594.450 ;
        RECT 238.950 592.950 244.050 593.400 ;
        RECT 262.800 592.950 264.900 593.400 ;
        RECT 266.100 592.950 271.050 595.050 ;
        RECT 286.950 594.450 289.050 598.050 ;
        RECT 301.950 595.950 304.050 599.400 ;
        RECT 313.950 598.950 316.050 599.400 ;
        RECT 319.950 598.950 322.050 599.400 ;
        RECT 325.950 598.950 328.050 604.050 ;
        RECT 329.400 603.450 330.450 605.400 ;
        RECT 331.950 605.400 376.050 606.450 ;
        RECT 331.950 604.950 334.050 605.400 ;
        RECT 373.950 604.950 376.050 605.400 ;
        RECT 449.400 605.400 493.050 606.450 ;
        RECT 449.400 604.050 450.450 605.400 ;
        RECT 490.950 604.950 493.050 605.400 ;
        RECT 673.950 606.450 676.050 607.050 ;
        RECT 682.950 606.450 685.050 607.050 ;
        RECT 673.950 605.400 685.050 606.450 ;
        RECT 673.950 604.950 676.050 605.400 ;
        RECT 682.950 604.950 685.050 605.400 ;
        RECT 691.950 606.450 694.050 607.050 ;
        RECT 709.950 606.450 712.050 607.050 ;
        RECT 691.950 605.400 712.050 606.450 ;
        RECT 691.950 604.950 694.050 605.400 ;
        RECT 709.950 604.950 712.050 605.400 ;
        RECT 718.950 606.450 721.050 607.050 ;
        RECT 760.950 606.450 763.050 607.050 ;
        RECT 718.950 605.400 763.050 606.450 ;
        RECT 718.950 604.950 721.050 605.400 ;
        RECT 760.950 604.950 763.050 605.400 ;
        RECT 337.950 603.450 340.050 604.050 ;
        RECT 370.950 603.450 373.050 604.050 ;
        RECT 329.400 602.400 373.050 603.450 ;
        RECT 337.950 601.950 340.050 602.400 ;
        RECT 370.950 601.950 373.050 602.400 ;
        RECT 424.950 603.450 427.050 604.050 ;
        RECT 424.950 602.400 441.450 603.450 ;
        RECT 424.950 601.950 427.050 602.400 ;
        RECT 316.950 597.450 319.050 598.050 ;
        RECT 322.950 597.450 325.050 598.050 ;
        RECT 316.950 596.400 325.050 597.450 ;
        RECT 316.950 595.950 319.050 596.400 ;
        RECT 322.950 595.950 325.050 596.400 ;
        RECT 328.950 594.450 331.050 598.050 ;
        RECT 331.950 597.450 334.050 601.050 ;
        RECT 349.950 600.450 352.050 601.050 ;
        RECT 358.950 600.450 364.050 601.050 ;
        RECT 376.950 600.450 382.050 601.050 ;
        RECT 349.950 599.400 364.050 600.450 ;
        RECT 349.950 598.950 352.050 599.400 ;
        RECT 358.950 598.950 364.050 599.400 ;
        RECT 365.400 599.400 382.050 600.450 ;
        RECT 365.400 597.450 366.450 599.400 ;
        RECT 376.950 598.950 382.050 599.400 ;
        RECT 331.950 597.000 366.450 597.450 ;
        RECT 332.400 596.400 366.450 597.000 ;
        RECT 385.950 595.950 388.050 601.050 ;
        RECT 418.950 598.950 424.050 601.050 ;
        RECT 440.400 600.450 441.450 602.400 ;
        RECT 445.950 601.950 451.050 604.050 ;
        RECT 442.950 600.450 448.050 601.050 ;
        RECT 440.400 599.400 448.050 600.450 ;
        RECT 442.950 598.950 448.050 599.400 ;
        RECT 457.950 598.950 460.050 604.050 ;
        RECT 502.950 601.950 508.050 604.050 ;
        RECT 463.950 598.050 466.050 601.050 ;
        RECT 400.950 597.450 403.050 598.050 ;
        RECT 409.950 597.450 412.050 598.050 ;
        RECT 400.950 596.400 412.050 597.450 ;
        RECT 400.950 595.950 403.050 596.400 ;
        RECT 409.950 595.950 412.050 596.400 ;
        RECT 415.950 597.450 418.050 598.050 ;
        RECT 430.950 597.450 433.050 598.050 ;
        RECT 415.950 596.400 433.050 597.450 ;
        RECT 415.950 595.950 418.050 596.400 ;
        RECT 430.950 595.950 433.050 596.400 ;
        RECT 436.950 597.450 439.050 598.050 ;
        RECT 460.800 597.450 462.900 598.050 ;
        RECT 436.950 596.400 462.900 597.450 ;
        RECT 436.950 595.950 439.050 596.400 ;
        RECT 460.800 595.950 462.900 596.400 ;
        RECT 463.800 597.000 466.050 598.050 ;
        RECT 467.100 597.000 469.200 598.050 ;
        RECT 463.800 595.950 465.900 597.000 ;
        RECT 466.950 595.950 469.200 597.000 ;
        RECT 481.950 595.950 484.050 601.050 ;
        RECT 535.950 598.950 538.050 604.050 ;
        RECT 550.950 603.450 553.050 604.050 ;
        RECT 550.950 602.400 558.450 603.450 ;
        RECT 550.950 601.950 553.050 602.400 ;
        RECT 557.400 601.050 558.450 602.400 ;
        RECT 574.950 601.950 580.050 604.050 ;
        RECT 544.950 600.450 549.000 601.050 ;
        RECT 544.950 598.950 549.450 600.450 ;
        RECT 550.950 598.950 556.050 601.050 ;
        RECT 557.400 599.400 562.050 601.050 ;
        RECT 558.000 598.950 562.050 599.400 ;
        RECT 286.950 594.000 331.050 594.450 ;
        RECT 331.950 594.450 334.050 595.050 ;
        RECT 343.950 594.450 346.050 595.050 ;
        RECT 286.950 593.400 330.450 594.000 ;
        RECT 331.950 593.400 346.050 594.450 ;
        RECT 286.950 592.950 289.050 593.400 ;
        RECT 331.950 592.950 334.050 593.400 ;
        RECT 343.950 592.950 346.050 593.400 ;
        RECT 373.950 594.450 376.050 595.050 ;
        RECT 397.800 594.450 399.900 595.050 ;
        RECT 373.950 593.400 399.900 594.450 ;
        RECT 373.950 592.950 376.050 593.400 ;
        RECT 397.800 592.950 399.900 593.400 ;
        RECT 401.100 592.950 406.050 595.050 ;
        RECT 421.950 594.450 424.050 595.050 ;
        RECT 451.950 594.450 454.050 595.050 ;
        RECT 421.950 593.400 454.050 594.450 ;
        RECT 421.950 592.950 424.050 593.400 ;
        RECT 451.950 592.950 454.050 593.400 ;
        RECT 460.950 594.450 463.050 595.050 ;
        RECT 466.950 594.450 469.050 595.950 ;
        RECT 487.950 595.050 490.050 598.050 ;
        RECT 502.950 597.450 505.050 598.050 ;
        RECT 502.950 596.400 516.450 597.450 ;
        RECT 502.950 595.950 505.050 596.400 ;
        RECT 460.950 594.000 469.050 594.450 ;
        RECT 460.950 593.400 468.600 594.000 ;
        RECT 460.950 592.950 463.050 593.400 ;
        RECT 475.950 592.950 481.050 595.050 ;
        RECT 484.800 594.000 486.900 595.050 ;
        RECT 487.950 594.000 490.200 595.050 ;
        RECT 511.950 594.450 514.050 595.050 ;
        RECT 484.800 592.950 487.050 594.000 ;
        RECT 488.100 592.950 490.200 594.000 ;
        RECT 491.400 593.400 514.050 594.450 ;
        RECT 515.400 594.450 516.450 596.400 ;
        RECT 517.950 595.950 522.900 598.050 ;
        RECT 524.100 595.950 529.050 598.050 ;
        RECT 520.950 594.450 523.050 595.050 ;
        RECT 515.400 593.400 531.450 594.450 ;
        RECT 212.400 591.450 213.450 592.950 ;
        RECT 247.950 591.450 250.050 592.050 ;
        RECT 212.400 590.400 250.050 591.450 ;
        RECT 247.950 589.950 250.050 590.400 ;
        RECT 268.950 591.450 271.050 592.050 ;
        RECT 286.950 591.450 289.050 592.050 ;
        RECT 268.950 590.400 289.050 591.450 ;
        RECT 268.950 589.950 271.050 590.400 ;
        RECT 286.950 589.950 289.050 590.400 ;
        RECT 28.950 588.450 31.050 589.050 ;
        RECT 40.950 588.450 43.050 589.050 ;
        RECT 28.950 587.400 43.050 588.450 ;
        RECT 28.950 586.950 31.050 587.400 ;
        RECT 40.950 586.950 43.050 587.400 ;
        RECT 103.950 588.450 106.050 589.050 ;
        RECT 127.950 588.450 130.050 589.050 ;
        RECT 202.950 588.450 205.050 589.050 ;
        RECT 103.950 587.400 205.050 588.450 ;
        RECT 103.950 586.950 106.050 587.400 ;
        RECT 127.950 586.950 130.050 587.400 ;
        RECT 202.950 586.950 205.050 587.400 ;
        RECT 298.950 588.450 301.050 589.050 ;
        RECT 316.950 588.450 319.050 589.050 ;
        RECT 298.950 587.400 319.050 588.450 ;
        RECT 298.950 586.950 301.050 587.400 ;
        RECT 316.950 586.950 319.050 587.400 ;
        RECT 370.950 586.950 373.050 592.050 ;
        RECT 484.950 591.450 487.050 592.950 ;
        RECT 491.400 591.450 492.450 593.400 ;
        RECT 511.950 592.950 514.050 593.400 ;
        RECT 520.950 592.950 523.050 593.400 ;
        RECT 484.950 591.000 492.450 591.450 ;
        RECT 485.250 590.400 492.450 591.000 ;
        RECT 530.400 591.450 531.450 593.400 ;
        RECT 532.950 592.950 535.050 598.050 ;
        RECT 538.950 595.950 544.050 598.050 ;
        RECT 548.400 597.450 549.450 598.950 ;
        RECT 556.950 597.450 559.050 598.050 ;
        RECT 548.400 596.400 559.050 597.450 ;
        RECT 556.950 595.950 559.050 596.400 ;
        RECT 562.950 592.950 565.050 598.050 ;
        RECT 574.950 597.450 577.050 601.050 ;
        RECT 580.950 598.950 586.050 601.050 ;
        RECT 588.000 600.450 592.050 601.050 ;
        RECT 595.800 600.450 597.900 601.050 ;
        RECT 587.400 599.400 597.900 600.450 ;
        RECT 587.400 598.950 592.050 599.400 ;
        RECT 595.800 598.950 597.900 599.400 ;
        RECT 599.100 600.450 601.200 601.050 ;
        RECT 625.950 600.450 628.050 601.050 ;
        RECT 599.100 599.400 628.050 600.450 ;
        RECT 656.400 600.000 672.450 600.450 ;
        RECT 599.100 598.950 601.200 599.400 ;
        RECT 625.950 598.950 628.050 599.400 ;
        RECT 655.950 599.400 673.050 600.000 ;
        RECT 587.400 597.450 588.450 598.950 ;
        RECT 595.950 597.450 598.050 598.050 ;
        RECT 574.950 597.000 588.450 597.450 ;
        RECT 575.400 596.400 588.450 597.000 ;
        RECT 590.400 596.400 598.050 597.450 ;
        RECT 583.950 594.450 586.050 595.200 ;
        RECT 590.400 594.450 591.450 596.400 ;
        RECT 595.950 595.950 598.050 596.400 ;
        RECT 655.950 595.950 658.050 599.400 ;
        RECT 670.950 595.950 673.050 599.400 ;
        RECT 673.950 598.950 676.050 604.050 ;
        RECT 727.950 603.450 730.050 604.050 ;
        RECT 805.950 603.450 808.050 604.050 ;
        RECT 680.400 603.000 717.450 603.450 ;
        RECT 679.950 602.400 717.450 603.000 ;
        RECT 679.950 598.950 682.050 602.400 ;
        RECT 716.400 601.050 717.450 602.400 ;
        RECT 727.950 602.400 808.050 603.450 ;
        RECT 727.950 601.050 730.050 602.400 ;
        RECT 805.950 601.950 808.050 602.400 ;
        RECT 826.950 603.450 829.050 604.050 ;
        RECT 826.950 602.400 843.450 603.450 ;
        RECT 826.950 601.950 829.050 602.400 ;
        RECT 842.400 601.050 843.450 602.400 ;
        RECT 706.950 600.450 709.050 601.050 ;
        RECT 712.950 600.450 715.050 601.050 ;
        RECT 706.950 599.400 715.050 600.450 ;
        RECT 716.400 599.400 724.050 601.050 ;
        RECT 706.950 598.950 709.050 599.400 ;
        RECT 712.950 598.950 715.050 599.400 ;
        RECT 717.000 598.950 724.050 599.400 ;
        RECT 727.800 600.000 730.050 601.050 ;
        RECT 727.800 598.950 729.900 600.000 ;
        RECT 731.100 598.950 736.050 601.050 ;
        RECT 769.800 600.000 771.900 601.050 ;
        RECT 773.100 600.450 775.200 601.050 ;
        RECT 778.950 600.450 781.050 601.050 ;
        RECT 769.800 598.950 772.050 600.000 ;
        RECT 773.100 599.400 781.050 600.450 ;
        RECT 773.100 598.950 775.200 599.400 ;
        RECT 778.950 598.950 781.050 599.400 ;
        RECT 583.950 593.400 591.450 594.450 ;
        RECT 643.950 594.450 646.050 595.050 ;
        RECT 652.950 594.450 655.050 595.050 ;
        RECT 643.950 593.400 655.050 594.450 ;
        RECT 583.950 593.100 586.050 593.400 ;
        RECT 643.950 592.950 646.050 593.400 ;
        RECT 652.950 592.950 655.050 593.400 ;
        RECT 658.950 594.450 661.050 595.050 ;
        RECT 667.950 594.450 670.050 595.050 ;
        RECT 658.950 593.400 670.050 594.450 ;
        RECT 658.950 592.950 661.050 593.400 ;
        RECT 667.950 592.950 670.050 593.400 ;
        RECT 676.950 592.950 679.050 598.050 ;
        RECT 691.950 597.450 694.050 598.050 ;
        RECT 709.950 597.450 712.050 598.050 ;
        RECT 691.950 596.400 712.050 597.450 ;
        RECT 691.950 595.950 694.050 596.400 ;
        RECT 709.950 595.950 712.050 596.400 ;
        RECT 715.950 597.450 718.050 598.050 ;
        RECT 724.950 597.450 727.050 598.050 ;
        RECT 730.950 597.450 733.050 598.050 ;
        RECT 715.950 596.400 733.050 597.450 ;
        RECT 715.950 595.950 718.050 596.400 ;
        RECT 724.950 595.950 727.050 596.400 ;
        RECT 730.950 595.950 733.050 596.400 ;
        RECT 736.950 597.450 739.050 598.050 ;
        RECT 751.950 597.450 754.050 598.050 ;
        RECT 736.950 596.400 754.050 597.450 ;
        RECT 736.950 595.950 739.050 596.400 ;
        RECT 751.950 595.950 754.050 596.400 ;
        RECT 769.950 595.950 772.050 598.950 ;
        RECT 775.950 597.450 778.050 598.050 ;
        RECT 790.950 597.450 793.050 598.050 ;
        RECT 775.950 596.400 793.050 597.450 ;
        RECT 775.950 595.950 778.050 596.400 ;
        RECT 790.950 595.950 793.050 596.400 ;
        RECT 805.950 595.950 810.900 598.050 ;
        RECT 838.950 595.950 841.050 601.050 ;
        RECT 842.400 599.400 850.050 601.050 ;
        RECT 843.000 598.950 850.050 599.400 ;
        RECT 688.800 594.000 690.900 595.050 ;
        RECT 692.100 594.450 697.050 595.050 ;
        RECT 700.950 594.450 703.050 595.050 ;
        RECT 688.800 592.950 691.050 594.000 ;
        RECT 692.100 593.400 703.050 594.450 ;
        RECT 692.100 592.950 697.050 593.400 ;
        RECT 700.950 592.950 703.050 593.400 ;
        RECT 739.950 594.450 742.050 595.050 ;
        RECT 748.950 594.450 753.900 595.050 ;
        RECT 739.950 593.400 753.900 594.450 ;
        RECT 739.950 592.950 742.050 593.400 ;
        RECT 748.950 592.950 753.900 593.400 ;
        RECT 755.100 594.450 757.200 595.050 ;
        RECT 769.950 594.450 772.050 595.050 ;
        RECT 755.100 593.400 772.050 594.450 ;
        RECT 755.100 592.950 757.200 593.400 ;
        RECT 769.950 592.950 772.050 593.400 ;
        RECT 784.950 592.950 790.050 595.050 ;
        RECT 535.950 591.450 538.050 592.050 ;
        RECT 530.400 590.400 538.050 591.450 ;
        RECT 535.950 589.950 538.050 590.400 ;
        RECT 583.950 591.450 586.050 591.900 ;
        RECT 592.950 591.450 595.050 592.050 ;
        RECT 583.950 590.400 595.050 591.450 ;
        RECT 583.950 589.800 586.050 590.400 ;
        RECT 592.950 589.950 595.050 590.400 ;
        RECT 670.950 591.450 673.050 592.050 ;
        RECT 688.950 591.450 691.050 592.950 ;
        RECT 670.950 591.000 691.050 591.450 ;
        RECT 706.950 591.450 709.050 592.050 ;
        RECT 770.400 591.450 771.450 592.950 ;
        RECT 793.950 591.450 796.050 595.050 ;
        RECT 850.950 592.950 853.050 598.050 ;
        RECT 670.950 590.400 690.300 591.000 ;
        RECT 706.950 590.400 768.450 591.450 ;
        RECT 770.400 591.000 796.050 591.450 ;
        RECT 770.400 590.400 795.450 591.000 ;
        RECT 670.950 589.950 673.050 590.400 ;
        RECT 706.950 589.950 709.050 590.400 ;
        RECT 457.950 588.450 460.050 589.050 ;
        RECT 601.950 588.450 604.050 589.050 ;
        RECT 634.950 588.450 637.050 589.050 ;
        RECT 457.950 587.400 637.050 588.450 ;
        RECT 457.950 586.950 460.050 587.400 ;
        RECT 601.950 586.950 604.050 587.400 ;
        RECT 634.950 586.950 637.050 587.400 ;
        RECT 652.950 588.450 655.050 589.050 ;
        RECT 676.950 588.450 679.050 589.050 ;
        RECT 652.950 587.400 679.050 588.450 ;
        RECT 652.950 586.950 655.050 587.400 ;
        RECT 676.950 586.950 679.050 587.400 ;
        RECT 724.950 588.450 727.050 589.050 ;
        RECT 754.950 588.450 757.050 589.050 ;
        RECT 724.950 587.400 757.050 588.450 ;
        RECT 767.400 588.450 768.450 590.400 ;
        RECT 787.950 588.450 790.050 589.050 ;
        RECT 767.400 587.400 790.050 588.450 ;
        RECT 724.950 586.950 727.050 587.400 ;
        RECT 754.950 586.950 757.050 587.400 ;
        RECT 787.950 586.950 790.050 587.400 ;
        RECT 70.950 585.450 73.050 586.050 ;
        RECT 136.950 585.450 139.050 586.050 ;
        RECT 70.950 584.400 139.050 585.450 ;
        RECT 70.950 583.950 73.050 584.400 ;
        RECT 136.950 583.950 139.050 584.400 ;
        RECT 160.950 585.450 163.050 586.050 ;
        RECT 208.950 585.450 211.050 586.050 ;
        RECT 160.950 584.400 211.050 585.450 ;
        RECT 160.950 583.950 163.050 584.400 ;
        RECT 208.950 583.950 211.050 584.400 ;
        RECT 226.950 585.450 229.050 586.050 ;
        RECT 313.950 585.450 316.050 586.050 ;
        RECT 226.950 584.400 316.050 585.450 ;
        RECT 226.950 583.950 229.050 584.400 ;
        RECT 313.950 583.950 316.050 584.400 ;
        RECT 367.950 585.450 370.050 586.050 ;
        RECT 403.950 585.450 406.050 586.050 ;
        RECT 367.950 584.400 406.050 585.450 ;
        RECT 367.950 583.950 370.050 584.400 ;
        RECT 403.950 583.950 406.050 584.400 ;
        RECT 430.950 585.450 433.050 586.050 ;
        RECT 586.800 585.450 588.900 586.050 ;
        RECT 430.950 584.400 588.900 585.450 ;
        RECT 430.950 583.950 433.050 584.400 ;
        RECT 586.800 583.950 588.900 584.400 ;
        RECT 590.100 585.450 592.200 586.050 ;
        RECT 655.950 585.450 658.050 586.050 ;
        RECT 706.800 585.450 708.900 586.050 ;
        RECT 590.100 584.400 708.900 585.450 ;
        RECT 590.100 583.950 592.200 584.400 ;
        RECT 655.950 583.950 658.050 584.400 ;
        RECT 706.800 583.950 708.900 584.400 ;
        RECT 710.100 585.450 712.200 586.050 ;
        RECT 727.950 585.450 730.050 586.050 ;
        RECT 710.100 584.400 730.050 585.450 ;
        RECT 710.100 583.950 712.200 584.400 ;
        RECT 727.950 583.950 730.050 584.400 ;
        RECT 100.950 582.450 103.050 583.050 ;
        RECT 166.950 582.450 169.050 583.050 ;
        RECT 190.950 582.450 193.050 583.050 ;
        RECT 100.950 581.400 193.050 582.450 ;
        RECT 100.950 580.950 103.050 581.400 ;
        RECT 166.950 580.950 169.050 581.400 ;
        RECT 190.950 580.950 193.050 581.400 ;
        RECT 199.950 582.450 202.050 583.050 ;
        RECT 217.950 582.450 220.050 583.050 ;
        RECT 199.950 581.400 220.050 582.450 ;
        RECT 199.950 580.950 202.050 581.400 ;
        RECT 217.950 580.950 220.050 581.400 ;
        RECT 265.950 582.450 268.050 583.050 ;
        RECT 271.950 582.450 274.050 583.050 ;
        RECT 457.950 582.450 460.050 583.050 ;
        RECT 265.950 581.400 274.050 582.450 ;
        RECT 265.950 580.950 268.050 581.400 ;
        RECT 271.950 580.950 274.050 581.400 ;
        RECT 275.400 581.400 460.050 582.450 ;
        RECT 16.950 579.450 19.050 580.050 ;
        RECT 275.400 579.450 276.450 581.400 ;
        RECT 457.950 580.950 460.050 581.400 ;
        RECT 577.950 582.450 580.050 583.050 ;
        RECT 595.950 582.450 598.050 583.050 ;
        RECT 577.950 581.400 598.050 582.450 ;
        RECT 577.950 580.950 580.050 581.400 ;
        RECT 595.950 580.950 598.050 581.400 ;
        RECT 640.950 582.450 643.050 583.050 ;
        RECT 670.800 582.450 672.900 583.050 ;
        RECT 640.950 581.400 672.900 582.450 ;
        RECT 640.950 580.950 643.050 581.400 ;
        RECT 670.800 580.950 672.900 581.400 ;
        RECT 674.100 582.450 676.200 583.050 ;
        RECT 781.950 582.450 784.050 583.050 ;
        RECT 674.100 581.400 784.050 582.450 ;
        RECT 674.100 580.950 676.200 581.400 ;
        RECT 781.950 580.950 784.050 581.400 ;
        RECT 820.950 582.450 823.050 583.050 ;
        RECT 832.950 582.450 835.050 583.050 ;
        RECT 820.950 581.400 835.050 582.450 ;
        RECT 820.950 580.950 823.050 581.400 ;
        RECT 832.950 580.950 835.050 581.400 ;
        RECT 16.950 578.400 276.450 579.450 ;
        RECT 334.950 579.450 337.050 580.050 ;
        RECT 454.950 579.450 457.050 580.050 ;
        RECT 334.950 578.400 457.050 579.450 ;
        RECT 16.950 577.950 19.050 578.400 ;
        RECT 334.950 577.950 337.050 578.400 ;
        RECT 454.950 577.950 457.050 578.400 ;
        RECT 478.950 579.450 481.050 580.050 ;
        RECT 505.950 579.450 508.050 580.050 ;
        RECT 478.950 578.400 508.050 579.450 ;
        RECT 478.950 577.950 481.050 578.400 ;
        RECT 505.950 577.950 508.050 578.400 ;
        RECT 517.950 579.450 520.050 580.050 ;
        RECT 532.950 579.450 535.050 580.050 ;
        RECT 541.950 579.450 544.050 580.050 ;
        RECT 517.950 578.400 544.050 579.450 ;
        RECT 517.950 577.950 520.050 578.400 ;
        RECT 532.950 577.950 535.050 578.400 ;
        RECT 541.950 577.950 544.050 578.400 ;
        RECT 562.950 579.450 565.050 580.050 ;
        RECT 598.950 579.450 601.050 580.050 ;
        RECT 562.950 578.400 601.050 579.450 ;
        RECT 562.950 577.950 565.050 578.400 ;
        RECT 598.950 577.950 601.050 578.400 ;
        RECT 613.950 579.450 616.050 580.050 ;
        RECT 763.950 579.450 766.050 580.050 ;
        RECT 793.950 579.450 796.050 580.050 ;
        RECT 613.950 578.400 796.050 579.450 ;
        RECT 613.950 577.950 616.050 578.400 ;
        RECT 763.950 577.950 766.050 578.400 ;
        RECT 793.950 577.950 796.050 578.400 ;
        RECT 238.950 576.450 241.050 577.050 ;
        RECT 244.950 576.450 247.050 577.050 ;
        RECT 238.950 575.400 247.050 576.450 ;
        RECT 238.950 574.950 241.050 575.400 ;
        RECT 244.950 574.950 247.050 575.400 ;
        RECT 259.950 576.450 262.050 577.050 ;
        RECT 292.950 576.450 295.050 577.050 ;
        RECT 259.950 575.400 295.050 576.450 ;
        RECT 259.950 574.950 262.050 575.400 ;
        RECT 292.950 574.950 295.050 575.400 ;
        RECT 322.950 576.450 325.050 577.050 ;
        RECT 379.950 576.450 382.050 577.050 ;
        RECT 322.950 575.400 382.050 576.450 ;
        RECT 322.950 574.950 325.050 575.400 ;
        RECT 379.950 574.950 382.050 575.400 ;
        RECT 385.950 576.450 388.050 577.050 ;
        RECT 439.950 576.450 442.050 577.050 ;
        RECT 466.950 576.450 469.050 577.050 ;
        RECT 385.950 575.400 469.050 576.450 ;
        RECT 385.950 574.950 388.050 575.400 ;
        RECT 439.950 574.950 442.050 575.400 ;
        RECT 466.950 574.950 469.050 575.400 ;
        RECT 28.950 573.450 31.050 574.050 ;
        RECT 70.950 573.450 73.050 574.050 ;
        RECT 28.950 572.400 73.050 573.450 ;
        RECT 28.950 571.950 31.050 572.400 ;
        RECT 70.950 571.950 73.050 572.400 ;
        RECT 232.950 573.450 235.050 574.050 ;
        RECT 262.950 573.450 265.050 574.050 ;
        RECT 298.800 573.450 300.900 574.050 ;
        RECT 232.950 572.400 300.900 573.450 ;
        RECT 232.950 571.950 235.050 572.400 ;
        RECT 262.950 571.950 265.050 572.400 ;
        RECT 298.800 571.950 300.900 572.400 ;
        RECT 302.100 573.450 304.200 574.050 ;
        RECT 337.950 573.450 340.050 574.050 ;
        RECT 302.100 572.400 340.050 573.450 ;
        RECT 302.100 571.950 304.200 572.400 ;
        RECT 337.950 571.950 340.050 572.400 ;
        RECT 409.950 573.450 412.050 574.050 ;
        RECT 469.950 573.450 472.050 574.050 ;
        RECT 409.950 572.400 472.050 573.450 ;
        RECT 487.950 573.450 490.050 577.050 ;
        RECT 619.950 576.450 622.050 577.050 ;
        RECT 676.950 576.450 679.050 577.050 ;
        RECT 619.950 575.400 679.050 576.450 ;
        RECT 619.950 574.950 622.050 575.400 ;
        RECT 676.950 574.950 679.050 575.400 ;
        RECT 691.950 576.450 694.050 577.050 ;
        RECT 745.950 576.450 748.050 577.050 ;
        RECT 691.950 575.400 748.050 576.450 ;
        RECT 691.950 574.950 694.050 575.400 ;
        RECT 745.950 574.950 748.050 575.400 ;
        RECT 778.950 576.450 781.050 577.050 ;
        RECT 814.950 576.450 817.050 577.050 ;
        RECT 778.950 575.400 817.050 576.450 ;
        RECT 778.950 574.950 781.050 575.400 ;
        RECT 814.950 574.950 817.050 575.400 ;
        RECT 562.950 573.450 565.050 574.050 ;
        RECT 487.950 573.000 565.050 573.450 ;
        RECT 488.400 572.400 565.050 573.000 ;
        RECT 409.950 571.950 412.050 572.400 ;
        RECT 469.950 571.950 472.050 572.400 ;
        RECT 562.950 571.950 565.050 572.400 ;
        RECT 613.950 573.450 616.050 574.050 ;
        RECT 706.950 573.450 709.050 574.050 ;
        RECT 613.950 572.400 709.050 573.450 ;
        RECT 613.950 571.950 616.050 572.400 ;
        RECT 706.950 571.950 709.050 572.400 ;
        RECT 721.950 573.450 724.050 574.050 ;
        RECT 781.950 573.450 784.050 574.050 ;
        RECT 721.950 572.400 784.050 573.450 ;
        RECT 721.950 571.950 724.050 572.400 ;
        RECT 781.950 571.950 784.050 572.400 ;
        RECT 787.950 573.450 790.050 574.050 ;
        RECT 796.950 573.450 799.050 574.050 ;
        RECT 787.950 572.400 799.050 573.450 ;
        RECT 787.950 571.950 790.050 572.400 ;
        RECT 796.950 571.950 799.050 572.400 ;
        RECT 34.950 570.450 37.050 571.050 ;
        RECT 52.950 570.450 55.050 571.050 ;
        RECT 34.950 569.400 55.050 570.450 ;
        RECT 34.950 568.950 37.050 569.400 ;
        RECT 52.950 568.950 55.050 569.400 ;
        RECT 145.950 570.450 148.050 571.050 ;
        RECT 187.950 570.450 190.050 571.050 ;
        RECT 145.950 569.400 190.050 570.450 ;
        RECT 145.950 568.950 148.050 569.400 ;
        RECT 187.950 568.950 190.050 569.400 ;
        RECT 247.950 570.450 250.050 571.050 ;
        RECT 364.950 570.450 367.050 571.050 ;
        RECT 247.950 569.400 367.050 570.450 ;
        RECT 247.950 568.950 250.050 569.400 ;
        RECT 364.950 568.950 367.050 569.400 ;
        RECT 376.950 570.450 379.050 571.050 ;
        RECT 448.950 570.450 451.050 571.050 ;
        RECT 376.950 569.400 451.050 570.450 ;
        RECT 376.950 568.950 379.050 569.400 ;
        RECT 448.950 568.950 451.050 569.400 ;
        RECT 460.950 568.050 463.050 571.050 ;
        RECT 466.950 570.450 469.050 571.050 ;
        RECT 619.950 570.450 622.050 571.050 ;
        RECT 466.950 569.400 622.050 570.450 ;
        RECT 466.950 568.950 469.050 569.400 ;
        RECT 619.950 568.950 622.050 569.400 ;
        RECT 79.950 567.450 82.050 568.050 ;
        RECT 127.950 567.450 130.050 568.050 ;
        RECT 79.950 566.400 130.050 567.450 ;
        RECT 79.950 565.950 82.050 566.400 ;
        RECT 127.950 565.950 130.050 566.400 ;
        RECT 154.950 567.450 157.050 568.050 ;
        RECT 172.950 567.450 175.050 568.050 ;
        RECT 238.950 567.450 241.050 568.050 ;
        RECT 154.950 566.400 241.050 567.450 ;
        RECT 154.950 565.950 157.050 566.400 ;
        RECT 172.950 565.950 175.050 566.400 ;
        RECT 238.950 565.950 241.050 566.400 ;
        RECT 277.950 567.450 280.050 568.050 ;
        RECT 295.950 567.450 298.050 568.050 ;
        RECT 310.800 567.450 312.900 568.050 ;
        RECT 277.950 566.400 312.900 567.450 ;
        RECT 277.950 565.950 280.050 566.400 ;
        RECT 295.950 565.950 298.050 566.400 ;
        RECT 310.800 565.950 312.900 566.400 ;
        RECT 314.100 565.950 319.050 568.050 ;
        RECT 397.950 567.450 400.050 568.050 ;
        RECT 427.950 567.450 430.050 568.050 ;
        RECT 442.950 567.450 445.050 568.050 ;
        RECT 451.950 567.450 454.050 568.050 ;
        RECT 397.950 566.400 454.050 567.450 ;
        RECT 397.950 565.950 400.050 566.400 ;
        RECT 427.950 565.950 430.050 566.400 ;
        RECT 442.950 565.950 445.050 566.400 ;
        RECT 451.950 565.950 454.050 566.400 ;
        RECT 457.950 567.000 463.050 568.050 ;
        RECT 463.950 567.450 466.050 568.050 ;
        RECT 487.950 567.450 490.050 568.050 ;
        RECT 457.950 566.400 462.450 567.000 ;
        RECT 463.950 566.400 490.050 567.450 ;
        RECT 457.950 565.950 462.000 566.400 ;
        RECT 463.950 565.950 466.050 566.400 ;
        RECT 487.950 565.950 490.050 566.400 ;
        RECT 511.950 567.450 514.050 568.050 ;
        RECT 547.950 567.450 550.050 568.050 ;
        RECT 511.950 566.400 550.050 567.450 ;
        RECT 637.950 567.300 640.050 569.400 ;
        RECT 511.950 565.950 514.050 566.400 ;
        RECT 547.950 565.950 550.050 566.400 ;
        RECT 43.950 564.450 46.050 565.050 ;
        RECT 148.950 564.450 151.050 565.050 ;
        RECT 157.950 564.450 160.050 565.050 ;
        RECT 199.950 564.450 202.050 565.050 ;
        RECT 259.950 564.450 262.050 565.050 ;
        RECT 43.950 563.400 72.450 564.450 ;
        RECT 43.950 562.950 46.050 563.400 ;
        RECT 71.400 562.050 72.450 563.400 ;
        RECT 148.950 563.400 180.450 564.450 ;
        RECT 148.950 562.950 151.050 563.400 ;
        RECT 157.950 562.950 160.050 563.400 ;
        RECT 179.400 562.050 180.450 563.400 ;
        RECT 199.950 563.400 262.050 564.450 ;
        RECT 199.950 562.950 202.050 563.400 ;
        RECT 259.950 562.950 262.050 563.400 ;
        RECT 265.950 564.450 268.050 565.050 ;
        RECT 301.950 564.450 304.050 565.050 ;
        RECT 265.950 563.400 304.050 564.450 ;
        RECT 265.950 562.950 268.050 563.400 ;
        RECT 301.950 562.950 304.050 563.400 ;
        RECT 442.950 564.450 445.050 565.050 ;
        RECT 502.950 564.450 505.050 565.050 ;
        RECT 442.950 563.400 505.050 564.450 ;
        RECT 442.950 562.950 445.050 563.400 ;
        RECT 502.950 562.950 505.050 563.400 ;
        RECT 532.950 564.450 537.000 565.050 ;
        RECT 568.950 564.450 571.050 565.050 ;
        RECT 532.950 564.000 537.450 564.450 ;
        RECT 532.950 562.950 538.050 564.000 ;
        RECT 406.950 562.050 409.050 562.200 ;
        RECT 1.950 558.450 4.050 559.050 ;
        RECT 22.950 558.450 25.050 559.050 ;
        RECT 28.950 558.450 31.050 559.050 ;
        RECT 1.950 557.400 31.050 558.450 ;
        RECT 1.950 556.950 4.050 557.400 ;
        RECT 22.950 556.950 25.050 557.400 ;
        RECT 28.950 556.950 31.050 557.400 ;
        RECT 34.950 556.950 37.050 562.050 ;
        RECT 70.950 561.450 73.050 562.050 ;
        RECT 121.950 561.450 124.050 562.050 ;
        RECT 70.950 560.400 124.050 561.450 ;
        RECT 70.950 559.950 73.050 560.400 ;
        RECT 121.950 559.950 124.050 560.400 ;
        RECT 127.950 561.450 133.050 562.050 ;
        RECT 145.950 561.450 148.050 562.050 ;
        RECT 172.950 561.450 175.050 562.050 ;
        RECT 127.950 560.400 148.050 561.450 ;
        RECT 155.550 561.000 175.050 561.450 ;
        RECT 127.950 559.950 133.050 560.400 ;
        RECT 145.950 559.950 148.050 560.400 ;
        RECT 154.950 560.400 175.050 561.000 ;
        RECT 151.800 559.050 153.900 559.200 ;
        RECT 40.950 558.450 43.050 559.050 ;
        RECT 49.800 558.450 51.900 559.050 ;
        RECT 40.950 558.000 51.900 558.450 ;
        RECT 53.100 558.450 58.050 559.050 ;
        RECT 76.950 558.450 79.050 559.050 ;
        RECT 40.950 557.400 52.050 558.000 ;
        RECT 40.950 556.950 43.050 557.400 ;
        RECT 49.800 556.950 52.050 557.400 ;
        RECT 53.100 557.400 79.050 558.450 ;
        RECT 53.100 556.950 58.050 557.400 ;
        RECT 76.950 556.950 79.050 557.400 ;
        RECT 88.950 558.450 91.050 559.050 ;
        RECT 106.950 558.450 109.050 559.050 ;
        RECT 88.950 557.400 109.050 558.450 ;
        RECT 88.950 556.950 91.050 557.400 ;
        RECT 106.950 556.950 109.050 557.400 ;
        RECT 112.950 558.450 115.050 559.050 ;
        RECT 127.950 558.450 132.900 559.050 ;
        RECT 112.950 557.400 132.900 558.450 ;
        RECT 134.100 558.000 136.200 559.050 ;
        RECT 112.950 556.950 115.050 557.400 ;
        RECT 127.950 556.950 132.900 557.400 ;
        RECT 133.950 556.950 136.200 558.000 ;
        RECT 145.800 558.000 147.900 559.050 ;
        RECT 145.800 556.950 148.050 558.000 ;
        RECT 149.100 557.100 153.900 559.050 ;
        RECT 154.950 559.050 157.050 560.400 ;
        RECT 154.950 558.000 157.200 559.050 ;
        RECT 149.100 556.950 153.000 557.100 ;
        RECT 155.100 556.950 157.200 558.000 ;
        RECT 172.950 556.950 175.050 560.400 ;
        RECT 178.950 561.450 181.050 562.050 ;
        RECT 187.950 561.450 190.050 562.050 ;
        RECT 178.950 560.400 190.050 561.450 ;
        RECT 178.950 559.950 181.050 560.400 ;
        RECT 187.950 559.950 190.050 560.400 ;
        RECT 196.950 561.450 199.050 562.050 ;
        RECT 226.950 561.450 229.050 562.050 ;
        RECT 196.950 560.400 229.050 561.450 ;
        RECT 196.950 559.950 199.050 560.400 ;
        RECT 49.950 556.050 52.050 556.950 ;
        RECT 16.950 553.950 22.050 556.050 ;
        RECT 25.950 555.450 28.050 556.050 ;
        RECT 31.950 555.450 34.050 556.050 ;
        RECT 25.950 554.400 34.050 555.450 ;
        RECT 25.950 553.950 28.050 554.400 ;
        RECT 31.950 553.950 34.050 554.400 ;
        RECT 37.950 555.450 40.050 556.050 ;
        RECT 43.800 555.450 45.900 556.050 ;
        RECT 37.950 554.400 45.900 555.450 ;
        RECT 37.950 553.950 40.050 554.400 ;
        RECT 43.800 553.950 45.900 554.400 ;
        RECT 47.100 555.000 52.050 556.050 ;
        RECT 47.100 554.400 51.300 555.000 ;
        RECT 47.100 553.950 51.000 554.400 ;
        RECT 52.950 553.950 57.900 556.050 ;
        RECT 59.100 555.450 61.200 556.050 ;
        RECT 72.000 555.900 75.000 556.050 ;
        RECT 70.950 555.450 76.050 555.900 ;
        RECT 59.100 554.400 76.050 555.450 ;
        RECT 59.100 553.950 61.200 554.400 ;
        RECT 70.950 553.950 76.050 554.400 ;
        RECT 85.950 555.450 88.050 556.050 ;
        RECT 100.950 555.450 103.050 556.050 ;
        RECT 85.950 554.400 103.050 555.450 ;
        RECT 85.950 553.950 88.050 554.400 ;
        RECT 100.950 553.950 103.050 554.400 ;
        RECT 109.950 555.450 112.050 556.050 ;
        RECT 133.950 555.450 136.050 556.950 ;
        RECT 109.950 555.000 136.050 555.450 ;
        RECT 109.950 554.400 135.600 555.000 ;
        RECT 70.950 553.800 73.050 553.950 ;
        RECT 73.950 553.800 76.050 553.950 ;
        RECT 76.950 550.950 82.050 553.050 ;
        RECT 109.950 552.450 112.050 554.400 ;
        RECT 145.950 553.950 148.050 556.950 ;
        RECT 152.100 555.000 154.200 556.050 ;
        RECT 151.950 553.950 154.200 555.000 ;
        RECT 157.950 553.950 163.050 556.050 ;
        RECT 178.950 553.950 181.050 559.050 ;
        RECT 193.950 553.950 196.050 559.050 ;
        RECT 199.950 558.450 202.050 559.050 ;
        RECT 208.950 558.450 211.050 559.050 ;
        RECT 199.950 557.400 211.050 558.450 ;
        RECT 199.950 556.950 202.050 557.400 ;
        RECT 208.950 556.950 211.050 557.400 ;
        RECT 226.950 556.950 229.050 560.400 ;
        RECT 232.950 556.950 238.050 559.050 ;
        RECT 247.950 556.950 250.050 562.050 ;
        RECT 283.950 561.450 286.050 562.050 ;
        RECT 304.950 561.450 309.900 562.050 ;
        RECT 283.950 560.400 309.900 561.450 ;
        RECT 283.950 559.950 286.050 560.400 ;
        RECT 304.950 559.950 309.900 560.400 ;
        RECT 311.100 561.450 313.200 562.050 ;
        RECT 316.950 561.450 319.050 562.050 ;
        RECT 311.100 560.400 319.050 561.450 ;
        RECT 311.100 559.950 313.200 560.400 ;
        RECT 316.950 559.950 319.050 560.400 ;
        RECT 328.950 561.450 331.050 562.050 ;
        RECT 337.950 561.450 340.050 562.050 ;
        RECT 328.950 560.400 340.050 561.450 ;
        RECT 328.950 559.950 331.050 560.400 ;
        RECT 337.950 559.950 340.050 560.400 ;
        RECT 352.950 561.450 355.050 562.050 ;
        RECT 358.950 561.450 364.050 562.050 ;
        RECT 352.950 560.400 364.050 561.450 ;
        RECT 352.950 559.950 355.050 560.400 ;
        RECT 358.950 559.950 364.050 560.400 ;
        RECT 367.950 561.450 370.050 562.050 ;
        RECT 376.950 561.450 379.050 562.050 ;
        RECT 367.950 560.400 379.050 561.450 ;
        RECT 367.950 559.950 370.050 560.400 ;
        RECT 376.950 559.950 379.050 560.400 ;
        RECT 391.950 561.450 394.050 562.050 ;
        RECT 397.950 561.450 400.050 562.050 ;
        RECT 391.950 560.400 400.050 561.450 ;
        RECT 391.950 559.950 394.050 560.400 ;
        RECT 397.950 559.950 400.050 560.400 ;
        RECT 403.950 560.100 409.050 562.050 ;
        RECT 403.950 559.950 408.000 560.100 ;
        RECT 433.950 559.950 439.050 562.050 ;
        RECT 448.950 561.450 451.050 562.050 ;
        RECT 469.950 561.450 472.050 562.050 ;
        RECT 448.950 560.400 465.450 561.450 ;
        RECT 448.950 559.950 451.050 560.400 ;
        RECT 253.950 558.450 256.050 559.050 ;
        RECT 265.950 558.450 268.050 559.050 ;
        RECT 284.400 558.450 285.450 559.950 ;
        RECT 253.950 557.400 268.050 558.450 ;
        RECT 275.400 558.000 285.450 558.450 ;
        RECT 253.950 556.950 256.050 557.400 ;
        RECT 265.950 556.950 268.050 557.400 ;
        RECT 274.950 557.400 285.450 558.000 ;
        RECT 217.950 555.450 220.050 556.050 ;
        RECT 229.950 555.450 232.050 556.050 ;
        RECT 235.950 555.450 238.050 556.050 ;
        RECT 247.800 555.450 249.900 556.050 ;
        RECT 217.950 554.400 232.050 555.450 ;
        RECT 217.950 553.950 220.050 554.400 ;
        RECT 229.950 553.950 232.050 554.400 ;
        RECT 233.400 554.400 249.900 555.450 ;
        RECT 251.100 555.000 253.200 556.050 ;
        RECT 151.950 553.050 154.050 553.950 ;
        RECT 148.800 552.450 150.900 553.050 ;
        RECT 109.950 551.400 150.900 552.450 ;
        RECT 151.950 552.000 154.200 553.050 ;
        RECT 109.950 550.950 112.050 551.400 ;
        RECT 148.800 550.950 150.900 551.400 ;
        RECT 152.100 550.950 154.200 552.000 ;
        RECT 214.950 552.450 217.050 553.050 ;
        RECT 233.400 552.450 234.450 554.400 ;
        RECT 235.950 553.950 238.050 554.400 ;
        RECT 247.800 553.950 249.900 554.400 ;
        RECT 250.950 553.950 253.200 555.000 ;
        RECT 256.950 555.450 259.050 556.050 ;
        RECT 262.950 555.450 265.050 556.050 ;
        RECT 256.950 554.400 265.050 555.450 ;
        RECT 256.950 553.950 259.050 554.400 ;
        RECT 262.950 553.950 265.050 554.400 ;
        RECT 274.950 553.950 277.050 557.400 ;
        RECT 304.950 556.950 310.050 559.050 ;
        RECT 283.950 553.950 289.050 556.050 ;
        RECT 292.950 553.950 298.050 556.050 ;
        RECT 316.950 555.450 319.050 556.050 ;
        RECT 322.950 555.450 325.050 556.050 ;
        RECT 316.950 554.400 325.050 555.450 ;
        RECT 316.950 553.950 319.050 554.400 ;
        RECT 322.950 553.950 325.050 554.400 ;
        RECT 328.950 553.950 331.050 559.050 ;
        RECT 361.950 556.950 367.050 559.050 ;
        RECT 379.950 558.450 382.050 559.050 ;
        RECT 368.400 557.400 382.050 558.450 ;
        RECT 334.950 555.450 337.050 556.050 ;
        RECT 346.950 555.450 349.050 556.050 ;
        RECT 334.950 554.400 349.050 555.450 ;
        RECT 334.950 553.950 337.050 554.400 ;
        RECT 346.950 553.950 349.050 554.400 ;
        RECT 352.950 555.450 355.050 556.050 ;
        RECT 368.400 555.450 369.450 557.400 ;
        RECT 379.950 556.950 382.050 557.400 ;
        RECT 400.950 558.450 403.050 559.050 ;
        RECT 406.950 558.450 409.050 558.900 ;
        RECT 418.950 558.450 423.900 559.050 ;
        RECT 400.950 557.400 409.050 558.450 ;
        RECT 400.950 556.950 403.050 557.400 ;
        RECT 406.950 556.800 409.050 557.400 ;
        RECT 410.400 557.400 423.900 558.450 ;
        RECT 352.950 554.400 369.450 555.450 ;
        RECT 397.950 555.450 400.050 556.050 ;
        RECT 410.400 555.450 411.450 557.400 ;
        RECT 418.950 556.950 423.900 557.400 ;
        RECT 425.100 556.950 430.050 559.050 ;
        RECT 439.950 556.950 445.050 559.050 ;
        RECT 454.800 558.450 456.900 559.050 ;
        RECT 446.400 557.400 456.900 558.450 ;
        RECT 397.950 554.400 411.450 555.450 ;
        RECT 352.950 553.950 355.050 554.400 ;
        RECT 397.950 553.950 400.050 554.400 ;
        RECT 412.950 553.950 418.050 556.050 ;
        RECT 214.950 551.400 234.450 552.450 ;
        RECT 238.950 552.450 241.050 553.050 ;
        RECT 250.950 552.450 253.050 553.950 ;
        RECT 238.950 552.000 253.050 552.450 ;
        RECT 265.950 552.450 268.050 553.050 ;
        RECT 271.950 552.450 274.050 553.050 ;
        RECT 238.950 551.400 252.450 552.000 ;
        RECT 265.950 551.400 274.050 552.450 ;
        RECT 214.950 550.950 217.050 551.400 ;
        RECT 238.950 550.950 241.050 551.400 ;
        RECT 265.950 550.950 268.050 551.400 ;
        RECT 271.950 550.950 274.050 551.400 ;
        RECT 55.950 549.450 58.050 550.050 ;
        RECT 109.950 549.450 112.050 550.050 ;
        RECT 55.950 548.400 112.050 549.450 ;
        RECT 55.950 547.950 58.050 548.400 ;
        RECT 109.950 547.950 112.050 548.400 ;
        RECT 130.950 549.450 133.050 550.050 ;
        RECT 163.950 549.450 166.050 550.050 ;
        RECT 130.950 548.400 166.050 549.450 ;
        RECT 130.950 547.950 133.050 548.400 ;
        RECT 163.950 547.950 166.050 548.400 ;
        RECT 193.950 549.450 196.050 550.050 ;
        RECT 262.950 549.450 265.050 550.050 ;
        RECT 193.950 548.400 265.050 549.450 ;
        RECT 193.950 547.950 196.050 548.400 ;
        RECT 262.950 547.950 265.050 548.400 ;
        RECT 277.950 547.950 280.050 553.050 ;
        RECT 289.950 549.450 292.050 553.050 ;
        RECT 304.950 552.450 307.050 553.050 ;
        RECT 316.950 552.450 319.050 553.050 ;
        RECT 304.950 551.400 319.050 552.450 ;
        RECT 304.950 550.950 307.050 551.400 ;
        RECT 316.950 550.950 319.050 551.400 ;
        RECT 328.950 552.450 331.050 553.050 ;
        RECT 349.950 552.450 352.050 553.050 ;
        RECT 328.950 551.400 352.050 552.450 ;
        RECT 328.950 550.950 331.050 551.400 ;
        RECT 349.950 550.950 352.050 551.400 ;
        RECT 358.950 552.450 361.050 553.050 ;
        RECT 370.950 552.450 373.050 553.050 ;
        RECT 358.950 551.400 373.050 552.450 ;
        RECT 358.950 550.950 361.050 551.400 ;
        RECT 370.950 550.950 373.050 551.400 ;
        RECT 379.950 552.450 382.050 553.050 ;
        RECT 388.950 552.450 391.050 553.050 ;
        RECT 379.950 551.400 391.050 552.450 ;
        RECT 379.950 550.950 382.050 551.400 ;
        RECT 388.950 550.950 391.050 551.400 ;
        RECT 406.950 552.450 409.050 553.050 ;
        RECT 421.950 552.450 424.050 556.050 ;
        RECT 446.400 555.450 447.450 557.400 ;
        RECT 454.800 556.950 456.900 557.400 ;
        RECT 457.800 558.000 459.900 559.050 ;
        RECT 461.100 558.000 463.200 559.050 ;
        RECT 457.800 556.950 460.050 558.000 ;
        RECT 457.950 556.050 460.050 556.950 ;
        RECT 437.400 554.400 447.450 555.450 ;
        RECT 437.400 553.050 438.450 554.400 ;
        RECT 448.950 553.950 454.050 556.050 ;
        RECT 457.800 555.000 460.050 556.050 ;
        RECT 460.950 556.950 463.200 558.000 ;
        RECT 464.400 558.450 465.450 560.400 ;
        RECT 469.950 561.000 498.450 561.450 ;
        RECT 469.950 560.400 499.050 561.000 ;
        RECT 469.950 559.950 472.050 560.400 ;
        RECT 469.950 558.450 472.050 559.050 ;
        RECT 464.400 557.400 472.050 558.450 ;
        RECT 469.950 556.950 472.050 557.400 ;
        RECT 496.950 556.950 499.050 560.400 ;
        RECT 502.950 556.950 505.050 562.050 ;
        RECT 511.950 561.450 514.050 562.050 ;
        RECT 511.950 561.000 534.450 561.450 ;
        RECT 511.950 560.400 535.050 561.000 ;
        RECT 511.950 559.950 514.050 560.400 ;
        RECT 532.950 556.950 535.050 560.400 ;
        RECT 535.950 559.950 538.050 562.950 ;
        RECT 554.400 563.400 571.050 564.450 ;
        RECT 638.850 563.700 640.050 567.300 ;
        RECT 658.950 566.400 661.050 568.500 ;
        RECT 673.950 567.300 676.050 569.400 ;
        RECT 541.950 562.050 544.050 562.200 ;
        RECT 541.950 561.450 547.050 562.050 ;
        RECT 554.400 561.450 555.450 563.400 ;
        RECT 568.950 562.950 571.050 563.400 ;
        RECT 541.950 560.400 555.450 561.450 ;
        RECT 541.950 560.100 547.050 560.400 ;
        RECT 543.000 559.950 547.050 560.100 ;
        RECT 556.950 559.950 562.050 562.050 ;
        RECT 577.950 559.050 580.050 562.050 ;
        RECT 586.950 559.950 592.050 562.050 ;
        RECT 538.950 558.900 543.000 559.050 ;
        RECT 538.950 556.950 544.050 558.900 ;
        RECT 547.950 558.450 550.050 559.050 ;
        RECT 553.950 558.450 556.050 559.050 ;
        RECT 547.950 557.400 556.050 558.450 ;
        RECT 547.950 556.950 550.050 557.400 ;
        RECT 553.950 556.950 556.050 557.400 ;
        RECT 559.950 556.950 565.050 559.050 ;
        RECT 568.950 558.450 571.050 559.050 ;
        RECT 574.800 558.450 576.900 559.050 ;
        RECT 568.950 557.400 576.900 558.450 ;
        RECT 568.950 556.950 571.050 557.400 ;
        RECT 574.800 556.950 576.900 557.400 ;
        RECT 577.800 558.000 580.050 559.050 ;
        RECT 581.100 558.000 583.200 559.050 ;
        RECT 577.800 556.950 579.900 558.000 ;
        RECT 580.950 556.950 583.200 558.000 ;
        RECT 598.950 556.950 604.050 559.050 ;
        RECT 616.950 556.950 622.050 559.050 ;
        RECT 625.950 556.950 628.050 562.050 ;
        RECT 637.950 561.600 640.050 563.700 ;
        RECT 460.950 556.050 463.050 556.950 ;
        RECT 541.950 556.800 544.050 556.950 ;
        RECT 460.950 555.000 463.200 556.050 ;
        RECT 464.100 555.000 466.200 556.050 ;
        RECT 457.800 553.950 459.900 555.000 ;
        RECT 461.100 553.950 463.200 555.000 ;
        RECT 463.950 553.950 466.200 555.000 ;
        RECT 469.950 555.450 472.050 556.050 ;
        RECT 475.800 555.450 477.900 556.050 ;
        RECT 469.950 554.400 477.900 555.450 ;
        RECT 469.950 553.950 472.050 554.400 ;
        RECT 475.800 553.950 477.900 554.400 ;
        RECT 479.100 555.450 484.050 556.050 ;
        RECT 493.950 555.450 496.050 556.050 ;
        RECT 479.100 554.400 496.050 555.450 ;
        RECT 479.100 553.950 484.050 554.400 ;
        RECT 493.950 553.950 496.050 554.400 ;
        RECT 499.950 555.450 502.050 556.050 ;
        RECT 511.950 555.450 514.050 556.050 ;
        RECT 499.950 554.400 514.050 555.450 ;
        RECT 499.950 553.950 502.050 554.400 ;
        RECT 511.950 553.950 514.050 554.400 ;
        RECT 436.950 552.450 439.050 553.050 ;
        RECT 406.950 551.400 439.050 552.450 ;
        RECT 406.950 550.950 409.050 551.400 ;
        RECT 436.950 550.950 439.050 551.400 ;
        RECT 463.950 552.450 466.050 553.950 ;
        RECT 478.950 552.450 481.050 553.050 ;
        RECT 463.950 551.400 481.050 552.450 ;
        RECT 463.950 550.950 466.050 551.400 ;
        RECT 478.950 550.950 481.050 551.400 ;
        RECT 490.950 552.450 493.050 553.050 ;
        RECT 517.950 552.450 520.050 556.050 ;
        RECT 523.950 555.450 526.050 556.050 ;
        RECT 556.950 555.450 559.050 556.050 ;
        RECT 523.950 554.400 559.050 555.450 ;
        RECT 523.950 553.950 526.050 554.400 ;
        RECT 556.950 553.950 559.050 554.400 ;
        RECT 568.950 555.450 571.050 556.050 ;
        RECT 580.950 555.450 583.050 556.950 ;
        RECT 568.950 555.000 583.050 555.450 ;
        RECT 586.950 555.450 589.050 556.050 ;
        RECT 595.950 555.450 598.050 556.050 ;
        RECT 568.950 554.400 582.600 555.000 ;
        RECT 586.950 554.400 598.050 555.450 ;
        RECT 568.950 553.950 571.050 554.400 ;
        RECT 586.950 553.950 589.050 554.400 ;
        RECT 595.950 553.950 598.050 554.400 ;
        RECT 604.950 553.950 610.050 556.050 ;
        RECT 490.950 552.000 520.050 552.450 ;
        RECT 520.950 552.450 523.050 553.050 ;
        RECT 532.950 552.450 535.050 553.050 ;
        RECT 616.950 552.450 619.050 556.050 ;
        RECT 490.950 551.400 519.450 552.000 ;
        RECT 520.950 551.400 535.050 552.450 ;
        RECT 490.950 550.950 493.050 551.400 ;
        RECT 520.950 550.950 523.050 551.400 ;
        RECT 532.950 550.950 535.050 551.400 ;
        RECT 575.400 551.400 621.450 552.450 ;
        RECT 298.950 549.450 301.050 550.050 ;
        RECT 289.950 549.000 301.050 549.450 ;
        RECT 290.400 548.400 301.050 549.000 ;
        RECT 298.950 547.950 301.050 548.400 ;
        RECT 307.950 549.450 310.050 550.050 ;
        RECT 329.400 549.450 330.450 550.950 ;
        RECT 307.950 548.400 330.450 549.450 ;
        RECT 334.950 549.450 337.050 550.050 ;
        RECT 355.950 549.450 358.050 550.050 ;
        RECT 409.950 549.450 412.050 550.050 ;
        RECT 334.950 548.400 358.050 549.450 ;
        RECT 307.950 547.950 310.050 548.400 ;
        RECT 334.950 547.950 337.050 548.400 ;
        RECT 355.950 547.950 358.050 548.400 ;
        RECT 389.400 548.400 412.050 549.450 ;
        RECT 46.950 546.450 49.050 547.050 ;
        RECT 79.950 546.450 82.050 547.050 ;
        RECT 118.950 546.450 121.050 547.050 ;
        RECT 46.950 545.400 82.050 546.450 ;
        RECT 46.950 544.950 49.050 545.400 ;
        RECT 79.950 544.950 82.050 545.400 ;
        RECT 86.400 545.400 121.050 546.450 ;
        RECT 73.950 543.450 76.050 544.050 ;
        RECT 86.400 543.450 87.450 545.400 ;
        RECT 118.950 544.950 121.050 545.400 ;
        RECT 208.950 546.450 211.050 547.050 ;
        RECT 286.950 546.450 289.050 547.050 ;
        RECT 208.950 545.400 289.050 546.450 ;
        RECT 208.950 544.950 211.050 545.400 ;
        RECT 286.950 544.950 289.050 545.400 ;
        RECT 313.950 546.450 316.050 547.050 ;
        RECT 389.400 546.450 390.450 548.400 ;
        RECT 409.950 547.950 412.050 548.400 ;
        RECT 421.950 549.450 424.050 550.050 ;
        RECT 460.950 549.450 463.050 550.050 ;
        RECT 421.950 548.400 463.050 549.450 ;
        RECT 421.950 547.950 424.050 548.400 ;
        RECT 460.950 547.950 463.050 548.400 ;
        RECT 520.950 549.450 523.050 550.050 ;
        RECT 575.400 549.450 576.450 551.400 ;
        RECT 520.950 548.400 576.450 549.450 ;
        RECT 577.950 549.450 580.050 550.050 ;
        RECT 604.950 549.450 607.050 550.050 ;
        RECT 577.950 548.400 607.050 549.450 ;
        RECT 620.400 549.450 621.450 551.400 ;
        RECT 622.950 550.950 625.050 556.050 ;
        RECT 631.950 553.950 637.050 556.050 ;
        RECT 628.950 549.450 631.050 550.050 ;
        RECT 638.850 549.600 640.050 561.600 ;
        RECT 643.950 553.950 649.050 556.050 ;
        RECT 652.950 550.950 655.050 556.050 ;
        RECT 659.100 549.600 660.300 566.400 ;
        RECT 674.850 563.700 676.050 567.300 ;
        RECT 694.950 566.400 697.050 568.500 ;
        RECT 709.950 567.300 712.050 569.400 ;
        RECT 673.950 561.600 676.050 563.700 ;
        RECT 667.950 553.950 673.050 556.050 ;
        RECT 674.850 549.600 676.050 561.600 ;
        RECT 685.950 556.950 691.050 559.050 ;
        RECT 679.950 553.950 685.050 556.050 ;
        RECT 695.100 549.600 696.300 566.400 ;
        RECT 710.850 563.700 712.050 567.300 ;
        RECT 730.950 566.400 733.050 568.500 ;
        RECT 763.950 567.450 766.050 568.050 ;
        RECT 778.950 567.450 781.050 568.050 ;
        RECT 763.950 566.400 781.050 567.450 ;
        RECT 799.950 567.300 802.050 569.400 ;
        RECT 709.950 561.600 712.050 563.700 ;
        RECT 703.950 553.950 709.050 556.050 ;
        RECT 710.850 549.600 712.050 561.600 ;
        RECT 715.950 553.950 720.900 556.050 ;
        RECT 722.100 553.950 727.050 556.050 ;
        RECT 731.100 549.600 732.300 566.400 ;
        RECT 763.950 565.950 766.050 566.400 ;
        RECT 778.950 565.950 781.050 566.400 ;
        RECT 745.950 564.450 748.050 565.050 ;
        RECT 745.950 564.000 774.450 564.450 ;
        RECT 745.950 563.400 775.050 564.000 ;
        RECT 800.850 563.700 802.050 567.300 ;
        RECT 820.950 566.400 823.050 568.500 ;
        RECT 745.950 562.950 748.050 563.400 ;
        RECT 763.950 559.950 769.050 562.050 ;
        RECT 772.950 559.950 775.050 563.400 ;
        RECT 799.950 561.600 802.050 563.700 ;
        RECT 745.950 559.050 748.050 559.200 ;
        RECT 745.950 557.100 751.050 559.050 ;
        RECT 747.000 556.950 751.050 557.100 ;
        RECT 754.950 558.450 757.050 559.050 ;
        RECT 769.950 558.450 772.050 559.050 ;
        RECT 754.950 557.400 772.050 558.450 ;
        RECT 754.950 556.950 757.050 557.400 ;
        RECT 769.950 556.950 772.050 557.400 ;
        RECT 781.950 558.450 784.050 559.050 ;
        RECT 787.950 558.450 790.050 559.050 ;
        RECT 781.950 557.400 790.050 558.450 ;
        RECT 781.950 556.950 784.050 557.400 ;
        RECT 787.950 556.950 790.050 557.400 ;
        RECT 742.950 553.950 747.900 556.050 ;
        RECT 749.100 553.950 754.050 556.050 ;
        RECT 793.950 553.950 799.050 556.050 ;
        RECT 733.950 552.450 736.050 553.050 ;
        RECT 763.950 552.450 766.050 553.050 ;
        RECT 733.950 551.400 766.050 552.450 ;
        RECT 733.950 550.950 736.050 551.400 ;
        RECT 763.950 550.950 766.050 551.400 ;
        RECT 620.400 548.400 631.050 549.450 ;
        RECT 520.950 547.950 523.050 548.400 ;
        RECT 577.950 547.950 580.050 548.400 ;
        RECT 604.950 547.950 607.050 548.400 ;
        RECT 628.950 547.950 631.050 548.400 ;
        RECT 637.950 547.500 640.050 549.600 ;
        RECT 658.950 547.500 661.050 549.600 ;
        RECT 673.950 547.500 676.050 549.600 ;
        RECT 694.950 547.500 697.050 549.600 ;
        RECT 709.950 547.500 712.050 549.600 ;
        RECT 730.950 547.500 733.050 549.600 ;
        RECT 754.950 549.450 757.050 550.050 ;
        RECT 766.950 549.450 769.050 550.050 ;
        RECT 754.950 548.400 769.050 549.450 ;
        RECT 754.950 547.950 757.050 548.400 ;
        RECT 766.950 547.950 769.050 548.400 ;
        RECT 784.950 547.950 787.050 553.050 ;
        RECT 800.850 549.600 802.050 561.600 ;
        RECT 805.950 553.950 810.900 556.050 ;
        RECT 812.100 553.950 817.050 556.050 ;
        RECT 821.100 549.600 822.300 566.400 ;
        RECT 841.950 558.450 844.050 559.050 ;
        RECT 853.950 558.450 856.050 559.050 ;
        RECT 841.950 557.400 856.050 558.450 ;
        RECT 841.950 556.950 844.050 557.400 ;
        RECT 853.950 556.950 856.050 557.400 ;
        RECT 823.950 552.450 826.050 553.050 ;
        RECT 835.950 552.450 838.050 553.050 ;
        RECT 850.950 552.450 853.050 553.050 ;
        RECT 823.950 551.400 853.050 552.450 ;
        RECT 823.950 550.950 826.050 551.400 ;
        RECT 835.950 550.950 838.050 551.400 ;
        RECT 850.950 550.950 853.050 551.400 ;
        RECT 799.950 547.500 802.050 549.600 ;
        RECT 820.950 547.500 823.050 549.600 ;
        RECT 313.950 545.400 390.450 546.450 ;
        RECT 391.950 546.450 394.050 547.050 ;
        RECT 439.950 546.450 442.050 547.050 ;
        RECT 391.950 545.400 442.050 546.450 ;
        RECT 313.950 544.950 316.050 545.400 ;
        RECT 391.950 544.950 394.050 545.400 ;
        RECT 439.950 544.950 442.050 545.400 ;
        RECT 469.950 546.450 472.050 547.050 ;
        RECT 571.950 546.450 574.050 547.050 ;
        RECT 619.950 546.450 622.050 547.050 ;
        RECT 469.950 545.400 564.450 546.450 ;
        RECT 469.950 544.950 472.050 545.400 ;
        RECT 73.950 542.400 87.450 543.450 ;
        RECT 193.950 543.450 196.050 544.050 ;
        RECT 202.950 543.450 205.050 544.050 ;
        RECT 193.950 542.400 205.050 543.450 ;
        RECT 73.950 541.950 76.050 542.400 ;
        RECT 193.950 541.950 196.050 542.400 ;
        RECT 202.950 541.950 205.050 542.400 ;
        RECT 214.950 543.450 217.050 544.050 ;
        RECT 220.950 543.450 223.050 544.050 ;
        RECT 214.950 542.400 223.050 543.450 ;
        RECT 287.400 543.450 288.450 544.950 ;
        RECT 349.950 543.450 352.050 544.050 ;
        RECT 481.950 543.450 484.050 544.050 ;
        RECT 287.400 542.400 352.050 543.450 ;
        RECT 214.950 541.950 217.050 542.400 ;
        RECT 220.950 541.950 223.050 542.400 ;
        RECT 349.950 541.950 352.050 542.400 ;
        RECT 383.400 542.400 484.050 543.450 ;
        RECT 563.400 543.450 564.450 545.400 ;
        RECT 571.950 545.400 622.050 546.450 ;
        RECT 571.950 544.950 574.050 545.400 ;
        RECT 619.950 544.950 622.050 545.400 ;
        RECT 715.950 546.450 718.050 547.050 ;
        RECT 724.950 546.450 727.050 547.050 ;
        RECT 715.950 545.400 727.050 546.450 ;
        RECT 715.950 544.950 718.050 545.400 ;
        RECT 724.950 544.950 727.050 545.400 ;
        RECT 736.950 546.450 739.050 547.050 ;
        RECT 736.950 545.400 777.450 546.450 ;
        RECT 736.950 544.950 739.050 545.400 ;
        RECT 574.950 543.450 577.050 544.050 ;
        RECT 563.400 542.400 577.050 543.450 ;
        RECT 383.400 541.050 384.450 542.400 ;
        RECT 481.950 541.950 484.050 542.400 ;
        RECT 574.950 541.950 577.050 542.400 ;
        RECT 622.950 543.450 625.050 544.050 ;
        RECT 652.950 543.450 655.050 544.050 ;
        RECT 622.950 542.400 655.050 543.450 ;
        RECT 622.950 541.950 625.050 542.400 ;
        RECT 652.950 541.950 655.050 542.400 ;
        RECT 664.950 543.450 667.050 544.050 ;
        RECT 706.950 543.450 709.050 544.050 ;
        RECT 712.950 543.450 715.050 544.050 ;
        RECT 664.950 542.400 715.050 543.450 ;
        RECT 664.950 541.950 667.050 542.400 ;
        RECT 706.950 541.950 709.050 542.400 ;
        RECT 712.950 541.950 715.050 542.400 ;
        RECT 718.950 543.450 721.050 544.050 ;
        RECT 739.950 543.450 742.050 544.050 ;
        RECT 718.950 542.400 742.050 543.450 ;
        RECT 776.400 543.450 777.450 545.400 ;
        RECT 805.950 543.450 808.050 544.050 ;
        RECT 776.400 542.400 808.050 543.450 ;
        RECT 718.950 541.950 721.050 542.400 ;
        RECT 739.950 541.950 742.050 542.400 ;
        RECT 805.950 541.950 808.050 542.400 ;
        RECT 205.950 540.450 208.050 541.050 ;
        RECT 217.950 540.450 220.050 541.050 ;
        RECT 205.950 539.400 220.050 540.450 ;
        RECT 205.950 538.950 208.050 539.400 ;
        RECT 217.950 538.950 220.050 539.400 ;
        RECT 232.950 540.450 235.050 541.050 ;
        RECT 274.950 540.450 277.050 541.050 ;
        RECT 382.950 540.450 385.050 541.050 ;
        RECT 232.950 539.400 273.450 540.450 ;
        RECT 232.950 538.950 235.050 539.400 ;
        RECT 10.950 537.450 13.050 538.050 ;
        RECT 34.950 537.450 37.050 538.050 ;
        RECT 10.950 536.400 37.050 537.450 ;
        RECT 10.950 535.950 13.050 536.400 ;
        RECT 34.950 535.950 37.050 536.400 ;
        RECT 211.950 537.450 214.050 538.050 ;
        RECT 259.950 537.450 262.050 538.050 ;
        RECT 211.950 536.400 262.050 537.450 ;
        RECT 272.400 537.450 273.450 539.400 ;
        RECT 274.950 539.400 385.050 540.450 ;
        RECT 274.950 538.950 277.050 539.400 ;
        RECT 382.950 538.950 385.050 539.400 ;
        RECT 457.950 540.450 460.050 541.050 ;
        RECT 478.950 540.450 481.050 541.050 ;
        RECT 457.950 539.400 481.050 540.450 ;
        RECT 457.950 538.950 460.050 539.400 ;
        RECT 478.950 538.950 481.050 539.400 ;
        RECT 502.950 540.450 505.050 541.050 ;
        RECT 559.950 540.450 562.050 541.050 ;
        RECT 502.950 539.400 562.050 540.450 ;
        RECT 502.950 538.950 505.050 539.400 ;
        RECT 559.950 538.950 562.050 539.400 ;
        RECT 586.950 540.450 589.050 541.050 ;
        RECT 670.950 540.450 673.050 541.050 ;
        RECT 586.950 539.400 673.050 540.450 ;
        RECT 586.950 538.950 589.050 539.400 ;
        RECT 670.950 538.950 673.050 539.400 ;
        RECT 721.950 540.450 724.050 541.050 ;
        RECT 748.950 540.450 751.050 541.050 ;
        RECT 721.950 539.400 751.050 540.450 ;
        RECT 721.950 538.950 724.050 539.400 ;
        RECT 748.950 538.950 751.050 539.400 ;
        RECT 757.950 540.450 760.050 541.050 ;
        RECT 781.950 540.450 784.050 541.050 ;
        RECT 757.950 539.400 784.050 540.450 ;
        RECT 757.950 538.950 760.050 539.400 ;
        RECT 781.950 538.950 784.050 539.400 ;
        RECT 301.950 537.450 304.050 538.050 ;
        RECT 361.950 537.450 364.050 538.050 ;
        RECT 272.400 536.400 364.050 537.450 ;
        RECT 211.950 535.950 214.050 536.400 ;
        RECT 259.950 535.950 262.050 536.400 ;
        RECT 301.950 535.950 304.050 536.400 ;
        RECT 361.950 535.950 364.050 536.400 ;
        RECT 415.950 537.450 418.050 538.050 ;
        RECT 427.950 537.450 430.050 538.050 ;
        RECT 415.950 536.400 430.050 537.450 ;
        RECT 415.950 535.950 418.050 536.400 ;
        RECT 427.950 535.950 430.050 536.400 ;
        RECT 436.950 537.450 439.050 538.050 ;
        RECT 493.950 537.450 496.050 538.050 ;
        RECT 541.950 537.450 544.050 538.050 ;
        RECT 436.950 536.400 544.050 537.450 ;
        RECT 436.950 535.950 439.050 536.400 ;
        RECT 493.950 535.950 496.050 536.400 ;
        RECT 541.950 535.950 544.050 536.400 ;
        RECT 550.950 537.450 553.050 538.050 ;
        RECT 562.950 537.450 565.050 538.050 ;
        RECT 550.950 536.400 565.050 537.450 ;
        RECT 550.950 535.950 553.050 536.400 ;
        RECT 562.950 535.950 565.050 536.400 ;
        RECT 625.950 537.450 628.050 538.050 ;
        RECT 646.950 537.450 649.050 538.050 ;
        RECT 682.950 537.450 685.050 538.050 ;
        RECT 625.950 536.400 685.050 537.450 ;
        RECT 625.950 535.950 628.050 536.400 ;
        RECT 646.950 535.950 649.050 536.400 ;
        RECT 682.950 535.950 685.050 536.400 ;
        RECT 760.950 537.450 763.050 538.050 ;
        RECT 760.950 536.400 774.450 537.450 ;
        RECT 760.950 535.950 763.050 536.400 ;
        RECT 64.950 534.450 67.050 535.050 ;
        RECT 106.950 534.450 109.050 535.050 ;
        RECT 118.950 534.450 121.050 535.050 ;
        RECT 193.950 534.450 196.050 535.050 ;
        RECT 232.950 534.450 235.050 535.050 ;
        RECT 64.950 534.000 162.450 534.450 ;
        RECT 64.950 533.400 163.050 534.000 ;
        RECT 64.950 532.950 67.050 533.400 ;
        RECT 106.950 532.950 109.050 533.400 ;
        RECT 118.950 532.950 121.050 533.400 ;
        RECT 25.950 531.450 28.050 532.050 ;
        RECT 17.250 531.000 28.050 531.450 ;
        RECT 16.950 530.400 28.050 531.000 ;
        RECT 16.950 529.050 19.050 530.400 ;
        RECT 25.950 529.950 28.050 530.400 ;
        RECT 7.950 526.950 12.900 529.050 ;
        RECT 14.100 528.000 19.050 529.050 ;
        RECT 20.100 528.450 22.200 529.050 ;
        RECT 28.950 528.450 31.050 529.050 ;
        RECT 14.100 526.950 18.900 528.000 ;
        RECT 20.100 527.400 31.050 528.450 ;
        RECT 20.100 526.950 22.200 527.400 ;
        RECT 13.950 523.950 18.900 526.050 ;
        RECT 20.100 525.000 22.200 526.050 ;
        RECT 19.950 523.950 22.200 525.000 ;
        RECT 28.950 523.950 31.050 527.400 ;
        RECT 34.950 523.950 37.050 529.050 ;
        RECT 49.950 528.450 52.050 529.050 ;
        RECT 49.950 528.000 72.450 528.450 ;
        RECT 49.950 527.400 73.050 528.000 ;
        RECT 49.950 526.950 52.050 527.400 ;
        RECT 19.950 522.450 22.050 523.950 ;
        RECT 49.950 523.050 52.050 526.050 ;
        RECT 55.950 523.050 58.050 526.050 ;
        RECT 70.950 523.950 73.050 527.400 ;
        RECT 73.950 526.950 76.050 532.050 ;
        RECT 160.950 531.450 163.050 533.400 ;
        RECT 193.950 533.400 235.050 534.450 ;
        RECT 193.950 532.950 196.050 533.400 ;
        RECT 232.950 532.950 235.050 533.400 ;
        RECT 241.950 534.450 244.050 535.050 ;
        RECT 271.950 534.450 274.050 535.050 ;
        RECT 241.950 533.400 274.050 534.450 ;
        RECT 241.950 532.950 244.050 533.400 ;
        RECT 271.950 532.950 274.050 533.400 ;
        RECT 343.950 534.450 346.050 535.050 ;
        RECT 373.950 534.450 376.050 535.050 ;
        RECT 466.950 534.450 469.050 535.050 ;
        RECT 487.950 534.450 490.050 535.050 ;
        RECT 343.950 533.400 376.050 534.450 ;
        RECT 407.400 534.000 469.050 534.450 ;
        RECT 343.950 532.950 346.050 533.400 ;
        RECT 373.950 532.950 376.050 533.400 ;
        RECT 406.950 533.400 469.050 534.000 ;
        RECT 160.950 530.400 168.450 531.450 ;
        RECT 160.950 529.950 163.050 530.400 ;
        RECT 167.400 529.050 168.450 530.400 ;
        RECT 82.950 528.450 85.050 529.050 ;
        RECT 82.950 527.400 90.450 528.450 ;
        RECT 82.950 526.950 85.050 527.400 ;
        RECT 28.800 522.450 30.900 523.050 ;
        RECT 19.950 522.000 30.900 522.450 ;
        RECT 32.100 522.000 34.200 523.050 ;
        RECT 20.550 521.400 30.900 522.000 ;
        RECT 28.800 520.950 30.900 521.400 ;
        RECT 31.950 520.950 34.200 522.000 ;
        RECT 40.950 522.450 43.050 523.050 ;
        RECT 49.800 522.450 52.050 523.050 ;
        RECT 40.950 522.000 52.050 522.450 ;
        RECT 52.800 522.000 54.900 523.050 ;
        RECT 55.950 522.450 58.200 523.050 ;
        RECT 76.950 522.450 79.050 526.050 ;
        RECT 89.400 525.450 90.450 527.400 ;
        RECT 91.950 526.950 96.900 529.050 ;
        RECT 98.100 526.950 103.050 529.050 ;
        RECT 94.950 525.450 97.050 526.050 ;
        RECT 89.400 524.400 97.050 525.450 ;
        RECT 94.950 523.950 97.050 524.400 ;
        RECT 55.950 522.000 79.050 522.450 ;
        RECT 100.950 522.450 103.050 526.050 ;
        RECT 112.950 523.950 115.050 529.050 ;
        RECT 118.950 523.950 121.050 529.050 ;
        RECT 136.950 526.950 142.050 529.050 ;
        RECT 167.400 527.400 172.050 529.050 ;
        RECT 168.000 526.950 172.050 527.400 ;
        RECT 175.950 526.950 178.050 532.050 ;
        RECT 181.950 528.450 184.050 529.050 ;
        RECT 187.950 528.450 190.050 529.050 ;
        RECT 181.950 527.400 190.050 528.450 ;
        RECT 181.950 526.950 184.050 527.400 ;
        RECT 187.950 526.950 190.050 527.400 ;
        RECT 205.950 528.450 208.050 529.050 ;
        RECT 229.950 528.450 234.900 529.050 ;
        RECT 205.950 527.400 234.900 528.450 ;
        RECT 205.950 526.950 208.050 527.400 ;
        RECT 229.950 526.950 234.900 527.400 ;
        RECT 236.100 528.450 238.200 529.050 ;
        RECT 244.950 528.450 247.050 529.050 ;
        RECT 253.950 528.450 256.050 529.050 ;
        RECT 236.100 527.400 256.050 528.450 ;
        RECT 236.100 526.950 238.200 527.400 ;
        RECT 244.950 526.950 247.050 527.400 ;
        RECT 253.950 526.950 256.050 527.400 ;
        RECT 259.950 526.950 262.050 532.050 ;
        RECT 280.950 531.450 283.050 532.050 ;
        RECT 280.950 530.400 294.450 531.450 ;
        RECT 280.950 529.950 283.050 530.400 ;
        RECT 293.400 529.050 294.450 530.400 ;
        RECT 295.950 529.950 300.900 532.050 ;
        RECT 302.100 531.000 304.200 532.050 ;
        RECT 334.950 531.450 340.050 532.050 ;
        RECT 301.950 529.950 304.200 531.000 ;
        RECT 323.400 530.400 340.050 531.450 ;
        RECT 265.950 526.950 271.050 529.050 ;
        RECT 293.400 527.400 298.050 529.050 ;
        RECT 294.000 526.950 298.050 527.400 ;
        RECT 301.950 526.950 304.050 529.950 ;
        RECT 316.950 526.950 322.050 529.050 ;
        RECT 323.400 526.050 324.450 530.400 ;
        RECT 334.950 529.950 340.050 530.400 ;
        RECT 349.950 531.450 352.050 532.050 ;
        RECT 388.950 531.450 391.050 532.050 ;
        RECT 397.950 531.450 400.050 532.050 ;
        RECT 349.950 531.000 372.450 531.450 ;
        RECT 349.950 530.400 373.050 531.000 ;
        RECT 349.950 529.950 352.050 530.400 ;
        RECT 106.950 522.450 109.050 523.050 ;
        RECT 100.950 522.000 109.050 522.450 ;
        RECT 40.950 521.400 51.900 522.000 ;
        RECT 40.950 520.950 43.050 521.400 ;
        RECT 49.800 520.950 51.900 521.400 ;
        RECT 52.800 520.950 55.050 522.000 ;
        RECT 56.100 521.400 78.450 522.000 ;
        RECT 101.400 521.400 109.050 522.000 ;
        RECT 56.100 520.950 58.200 521.400 ;
        RECT 106.950 520.950 109.050 521.400 ;
        RECT 13.950 519.450 16.050 520.050 ;
        RECT 31.950 519.450 34.050 520.950 ;
        RECT 13.950 519.000 34.050 519.450 ;
        RECT 52.950 519.450 55.050 520.950 ;
        RECT 73.950 519.450 76.050 520.050 ;
        RECT 52.950 519.000 76.050 519.450 ;
        RECT 13.950 518.400 33.600 519.000 ;
        RECT 53.250 518.400 76.050 519.000 ;
        RECT 13.950 517.950 16.050 518.400 ;
        RECT 73.950 517.950 76.050 518.400 ;
        RECT 115.950 517.950 118.050 523.050 ;
        RECT 124.950 522.450 127.050 523.050 ;
        RECT 124.950 521.400 132.450 522.450 ;
        RECT 124.950 520.950 127.050 521.400 ;
        RECT 131.400 519.450 132.450 521.400 ;
        RECT 133.950 520.950 136.050 526.050 ;
        RECT 139.950 525.450 142.050 526.050 ;
        RECT 154.950 525.450 157.050 526.050 ;
        RECT 139.950 524.400 157.050 525.450 ;
        RECT 139.950 523.950 142.050 524.400 ;
        RECT 154.950 523.950 157.050 524.400 ;
        RECT 172.950 523.950 175.050 526.050 ;
        RECT 178.950 525.450 181.050 526.050 ;
        RECT 184.950 525.450 187.050 526.050 ;
        RECT 193.950 525.450 196.050 526.050 ;
        RECT 178.950 524.400 196.050 525.450 ;
        RECT 178.950 523.950 181.050 524.400 ;
        RECT 184.950 523.950 187.050 524.400 ;
        RECT 193.950 523.950 196.050 524.400 ;
        RECT 199.950 523.950 205.050 526.050 ;
        RECT 217.950 523.950 223.050 526.050 ;
        RECT 241.950 525.450 244.050 526.050 ;
        RECT 247.950 525.450 250.050 526.050 ;
        RECT 256.950 525.450 259.050 526.050 ;
        RECT 241.950 524.400 259.050 525.450 ;
        RECT 241.950 523.950 244.050 524.400 ;
        RECT 247.950 523.950 250.050 524.400 ;
        RECT 256.950 523.950 259.050 524.400 ;
        RECT 173.400 520.050 174.450 523.950 ;
        RECT 190.950 522.450 193.050 523.050 ;
        RECT 196.950 522.450 199.050 523.050 ;
        RECT 190.950 521.400 199.050 522.450 ;
        RECT 190.950 520.950 193.050 521.400 ;
        RECT 196.950 520.950 199.050 521.400 ;
        RECT 205.950 522.450 208.050 523.050 ;
        RECT 214.800 522.450 216.900 523.050 ;
        RECT 205.950 521.400 216.900 522.450 ;
        RECT 218.100 522.000 220.200 523.050 ;
        RECT 205.950 520.950 208.050 521.400 ;
        RECT 214.800 520.950 216.900 521.400 ;
        RECT 217.950 520.950 220.200 522.000 ;
        RECT 223.950 522.450 226.050 523.050 ;
        RECT 229.950 522.450 232.050 523.050 ;
        RECT 238.950 522.450 241.050 523.050 ;
        RECT 262.950 522.450 265.050 526.050 ;
        RECT 283.950 525.450 286.050 526.050 ;
        RECT 310.950 525.450 313.050 526.050 ;
        RECT 283.950 524.400 313.050 525.450 ;
        RECT 283.950 523.950 286.050 524.400 ;
        RECT 310.950 523.950 313.050 524.400 ;
        RECT 223.950 521.400 232.050 522.450 ;
        RECT 223.950 520.950 226.050 521.400 ;
        RECT 229.950 520.950 232.050 521.400 ;
        RECT 233.400 521.400 276.450 522.450 ;
        RECT 173.400 519.450 178.050 520.050 ;
        RECT 131.400 518.400 178.050 519.450 ;
        RECT 217.950 519.450 220.050 520.950 ;
        RECT 233.400 519.450 234.450 521.400 ;
        RECT 238.950 520.950 241.050 521.400 ;
        RECT 217.950 519.000 234.450 519.450 ;
        RECT 218.550 518.400 234.450 519.000 ;
        RECT 275.400 519.450 276.450 521.400 ;
        RECT 277.950 520.950 283.050 523.050 ;
        RECT 286.950 520.950 292.050 523.050 ;
        RECT 316.950 520.950 319.050 526.050 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 325.950 525.450 328.050 529.050 ;
        RECT 340.950 528.450 343.050 529.050 ;
        RECT 352.950 528.450 355.050 529.200 ;
        RECT 340.950 527.400 355.050 528.450 ;
        RECT 340.950 526.950 343.050 527.400 ;
        RECT 352.950 527.100 355.050 527.400 ;
        RECT 370.950 526.950 373.050 530.400 ;
        RECT 388.950 530.400 400.050 531.450 ;
        RECT 379.950 528.450 382.050 529.050 ;
        RECT 388.950 528.450 391.050 530.400 ;
        RECT 397.950 529.950 400.050 530.400 ;
        RECT 406.950 529.950 409.050 533.400 ;
        RECT 466.950 532.950 469.050 533.400 ;
        RECT 482.400 533.400 490.050 534.450 ;
        RECT 439.950 532.050 442.050 532.200 ;
        RECT 439.950 530.100 445.050 532.050 ;
        RECT 441.000 529.950 445.050 530.100 ;
        RECT 472.950 531.450 475.050 532.050 ;
        RECT 482.400 531.450 483.450 533.400 ;
        RECT 487.950 532.950 490.050 533.400 ;
        RECT 574.950 534.450 577.050 535.050 ;
        RECT 664.950 534.450 667.050 535.050 ;
        RECT 574.950 533.400 667.050 534.450 ;
        RECT 727.950 533.400 730.050 535.500 ;
        RECT 748.950 533.400 751.050 535.500 ;
        RECT 773.400 534.450 774.450 536.400 ;
        RECT 856.950 534.450 859.050 535.050 ;
        RECT 773.400 533.400 859.050 534.450 ;
        RECT 574.950 532.950 577.050 533.400 ;
        RECT 664.950 532.950 667.050 533.400 ;
        RECT 472.950 531.000 483.450 531.450 ;
        RECT 484.950 531.450 487.050 532.050 ;
        RECT 490.950 531.450 493.050 532.050 ;
        RECT 499.950 531.450 502.050 532.050 ;
        RECT 472.950 530.400 484.050 531.000 ;
        RECT 472.950 529.950 475.050 530.400 ;
        RECT 481.950 529.050 484.050 530.400 ;
        RECT 484.950 530.400 502.050 531.450 ;
        RECT 484.950 529.950 487.050 530.400 ;
        RECT 490.950 529.950 493.050 530.400 ;
        RECT 499.950 529.950 502.050 530.400 ;
        RECT 511.950 531.450 514.050 532.050 ;
        RECT 523.950 531.450 526.050 532.050 ;
        RECT 511.950 530.400 526.050 531.450 ;
        RECT 511.950 529.950 514.050 530.400 ;
        RECT 379.950 528.000 391.050 528.450 ;
        RECT 391.950 528.450 394.050 529.050 ;
        RECT 403.800 528.450 405.900 529.050 ;
        RECT 379.950 527.400 390.450 528.000 ;
        RECT 391.950 527.400 405.900 528.450 ;
        RECT 379.950 526.950 382.050 527.400 ;
        RECT 391.950 526.950 394.050 527.400 ;
        RECT 403.800 526.950 405.900 527.400 ;
        RECT 407.100 526.950 412.050 529.050 ;
        RECT 415.950 528.450 418.050 529.050 ;
        RECT 421.950 528.450 424.050 529.050 ;
        RECT 415.950 527.400 424.050 528.450 ;
        RECT 415.950 526.950 418.050 527.400 ;
        RECT 421.950 526.950 424.050 527.400 ;
        RECT 427.950 528.450 430.050 529.050 ;
        RECT 436.800 528.450 438.900 529.050 ;
        RECT 427.950 527.400 438.900 528.450 ;
        RECT 427.950 526.950 430.050 527.400 ;
        RECT 436.800 526.950 438.900 527.400 ;
        RECT 440.100 528.450 442.200 528.900 ;
        RECT 440.100 528.000 459.600 528.450 ;
        RECT 478.800 528.000 480.900 529.050 ;
        RECT 481.800 528.000 484.050 529.050 ;
        RECT 485.100 528.000 487.200 529.050 ;
        RECT 440.100 527.400 460.050 528.000 ;
        RECT 440.100 526.800 442.200 527.400 ;
        RECT 457.950 526.050 460.050 527.400 ;
        RECT 478.800 526.950 481.050 528.000 ;
        RECT 481.800 526.950 483.900 528.000 ;
        RECT 484.950 526.950 487.200 528.000 ;
        RECT 490.950 528.450 493.050 529.050 ;
        RECT 502.950 528.450 505.050 529.050 ;
        RECT 490.950 527.400 505.050 528.450 ;
        RECT 490.950 526.950 493.050 527.400 ;
        RECT 502.950 526.950 505.050 527.400 ;
        RECT 517.950 526.950 520.050 530.400 ;
        RECT 523.950 529.950 526.050 530.400 ;
        RECT 544.950 531.450 547.050 532.050 ;
        RECT 616.950 531.450 619.050 532.050 ;
        RECT 640.950 531.450 643.050 532.050 ;
        RECT 544.950 530.400 561.450 531.450 ;
        RECT 544.950 529.950 547.050 530.400 ;
        RECT 560.400 529.050 561.450 530.400 ;
        RECT 616.950 530.400 643.050 531.450 ;
        RECT 616.950 529.950 619.050 530.400 ;
        RECT 640.950 529.950 643.050 530.400 ;
        RECT 709.950 531.450 712.050 532.050 ;
        RECT 709.950 530.400 723.450 531.450 ;
        RECT 709.950 529.950 712.050 530.400 ;
        RECT 722.400 529.050 723.450 530.400 ;
        RECT 526.950 528.450 529.050 529.050 ;
        RECT 556.950 528.450 559.050 529.050 ;
        RECT 526.950 527.400 559.050 528.450 ;
        RECT 560.400 527.400 565.050 529.050 ;
        RECT 526.950 526.950 529.050 527.400 ;
        RECT 556.950 526.950 559.050 527.400 ;
        RECT 561.000 526.950 565.050 527.400 ;
        RECT 637.950 528.450 640.050 529.050 ;
        RECT 637.950 527.400 645.450 528.450 ;
        RECT 637.950 526.950 640.050 527.400 ;
        RECT 352.950 525.450 355.050 526.050 ;
        RECT 325.950 525.000 355.050 525.450 ;
        RECT 326.400 524.400 355.050 525.000 ;
        RECT 352.950 523.800 355.050 524.400 ;
        RECT 364.950 523.950 370.050 526.050 ;
        RECT 331.950 522.450 334.050 523.050 ;
        RECT 337.950 522.450 340.050 523.050 ;
        RECT 349.950 522.450 352.050 523.050 ;
        RECT 331.950 521.400 352.050 522.450 ;
        RECT 331.950 520.950 334.050 521.400 ;
        RECT 337.950 520.950 340.050 521.400 ;
        RECT 349.950 520.950 352.050 521.400 ;
        RECT 322.950 519.450 325.050 520.050 ;
        RECT 275.400 518.400 325.050 519.450 ;
        RECT 355.950 519.450 358.050 523.050 ;
        RECT 361.950 522.450 364.050 523.050 ;
        RECT 373.950 522.450 376.050 526.050 ;
        RECT 394.950 525.450 397.050 526.050 ;
        RECT 400.950 525.450 403.050 526.050 ;
        RECT 394.950 524.400 403.050 525.450 ;
        RECT 394.950 523.950 397.050 524.400 ;
        RECT 400.950 523.950 403.050 524.400 ;
        RECT 421.950 523.950 427.050 526.050 ;
        RECT 430.950 523.950 436.050 526.050 ;
        RECT 448.950 525.450 451.050 526.050 ;
        RECT 454.800 525.450 456.900 526.050 ;
        RECT 448.950 524.400 456.900 525.450 ;
        RECT 457.950 525.000 460.200 526.050 ;
        RECT 448.950 523.950 451.050 524.400 ;
        RECT 454.800 523.950 456.900 524.400 ;
        RECT 458.100 523.950 460.200 525.000 ;
        RECT 463.950 523.950 469.050 526.050 ;
        RECT 478.950 523.950 481.050 526.950 ;
        RECT 484.950 523.950 487.050 526.950 ;
        RECT 493.950 525.450 496.050 526.050 ;
        RECT 514.950 525.450 517.050 526.050 ;
        RECT 493.950 524.400 517.050 525.450 ;
        RECT 493.950 523.950 496.050 524.400 ;
        RECT 514.950 523.950 517.050 524.400 ;
        RECT 520.950 525.450 523.050 526.050 ;
        RECT 535.800 525.450 537.900 526.050 ;
        RECT 520.950 524.400 537.900 525.450 ;
        RECT 361.950 522.000 376.050 522.450 ;
        RECT 361.950 521.400 375.450 522.000 ;
        RECT 361.950 520.950 364.050 521.400 ;
        RECT 460.950 520.950 466.050 523.050 ;
        RECT 508.950 522.450 511.050 523.050 ;
        RECT 520.950 522.450 523.050 524.400 ;
        RECT 535.800 523.950 537.900 524.400 ;
        RECT 539.100 523.950 544.050 526.050 ;
        RECT 556.950 523.950 561.900 526.050 ;
        RECT 574.950 523.950 580.050 526.050 ;
        RECT 605.100 525.450 607.200 526.050 ;
        RECT 619.950 525.450 622.050 526.050 ;
        RECT 625.950 525.450 628.050 526.050 ;
        RECT 605.100 524.400 628.050 525.450 ;
        RECT 644.400 525.450 645.450 527.400 ;
        RECT 646.950 526.950 652.050 529.050 ;
        RECT 655.950 528.450 658.050 529.050 ;
        RECT 664.950 528.450 667.050 529.050 ;
        RECT 655.950 527.400 667.050 528.450 ;
        RECT 655.950 526.950 658.050 527.400 ;
        RECT 664.950 526.950 667.050 527.400 ;
        RECT 679.950 528.450 682.050 529.050 ;
        RECT 685.950 528.450 688.050 529.050 ;
        RECT 679.950 527.400 688.050 528.450 ;
        RECT 679.950 526.950 682.050 527.400 ;
        RECT 685.950 526.950 688.050 527.400 ;
        RECT 694.950 528.450 697.050 529.050 ;
        RECT 718.950 528.450 721.050 529.050 ;
        RECT 694.950 527.400 721.050 528.450 ;
        RECT 722.400 527.400 727.050 529.050 ;
        RECT 694.950 526.950 697.050 527.400 ;
        RECT 718.950 526.950 721.050 527.400 ;
        RECT 723.000 526.950 727.050 527.400 ;
        RECT 652.950 525.450 655.050 526.050 ;
        RECT 644.400 524.400 655.050 525.450 ;
        RECT 605.100 523.950 607.200 524.400 ;
        RECT 619.950 523.950 622.050 524.400 ;
        RECT 625.950 523.950 628.050 524.400 ;
        RECT 652.950 523.950 655.050 524.400 ;
        RECT 658.950 525.450 661.050 526.050 ;
        RECT 673.950 525.450 676.050 526.050 ;
        RECT 658.950 524.400 676.050 525.450 ;
        RECT 658.950 523.950 661.050 524.400 ;
        RECT 673.950 523.950 676.050 524.400 ;
        RECT 688.950 523.950 694.050 526.050 ;
        RECT 697.950 525.450 700.050 526.050 ;
        RECT 712.950 525.450 715.050 526.050 ;
        RECT 697.950 524.400 715.050 525.450 ;
        RECT 697.950 523.950 700.050 524.400 ;
        RECT 712.950 523.950 715.050 524.400 ;
        RECT 508.950 522.000 523.050 522.450 ;
        RECT 523.950 522.450 526.050 523.050 ;
        RECT 538.950 522.450 541.050 523.050 ;
        RECT 508.950 521.400 522.450 522.000 ;
        RECT 523.950 521.400 541.050 522.450 ;
        RECT 508.950 520.950 511.050 521.400 ;
        RECT 523.950 520.950 526.050 521.400 ;
        RECT 538.950 520.950 541.050 521.400 ;
        RECT 580.950 522.450 583.050 523.200 ;
        RECT 622.950 522.450 625.050 523.050 ;
        RECT 580.950 521.400 625.050 522.450 ;
        RECT 580.950 521.100 583.050 521.400 ;
        RECT 622.950 520.950 625.050 521.400 ;
        RECT 667.950 520.950 673.050 523.050 ;
        RECT 373.950 519.450 376.050 520.050 ;
        RECT 388.950 519.450 391.050 520.050 ;
        RECT 355.950 519.000 391.050 519.450 ;
        RECT 174.000 517.950 178.050 518.400 ;
        RECT 226.950 517.050 229.050 518.400 ;
        RECT 322.950 517.950 325.050 518.400 ;
        RECT 356.400 518.400 391.050 519.000 ;
        RECT 43.950 516.450 46.050 517.050 ;
        RECT 55.950 516.450 58.050 517.050 ;
        RECT 43.950 515.400 58.050 516.450 ;
        RECT 43.950 514.950 46.050 515.400 ;
        RECT 55.950 514.950 58.050 515.400 ;
        RECT 112.950 516.450 115.050 517.050 ;
        RECT 133.950 516.450 136.050 517.050 ;
        RECT 112.950 515.400 136.050 516.450 ;
        RECT 112.950 514.950 115.050 515.400 ;
        RECT 133.950 514.950 136.050 515.400 ;
        RECT 148.950 516.450 151.050 517.050 ;
        RECT 202.950 516.450 205.050 517.050 ;
        RECT 148.950 515.400 205.050 516.450 ;
        RECT 148.950 514.950 151.050 515.400 ;
        RECT 202.950 514.950 205.050 515.400 ;
        RECT 226.800 516.000 229.050 517.050 ;
        RECT 230.100 516.450 232.200 517.050 ;
        RECT 235.950 516.450 238.050 517.050 ;
        RECT 226.800 514.950 228.900 516.000 ;
        RECT 230.100 515.400 238.050 516.450 ;
        RECT 230.100 514.950 232.200 515.400 ;
        RECT 235.950 514.950 238.050 515.400 ;
        RECT 283.950 516.450 286.050 517.050 ;
        RECT 298.950 516.450 301.050 517.050 ;
        RECT 283.950 515.400 301.050 516.450 ;
        RECT 283.950 514.950 286.050 515.400 ;
        RECT 298.950 514.950 301.050 515.400 ;
        RECT 304.950 516.450 307.050 517.050 ;
        RECT 337.950 516.450 340.050 517.050 ;
        RECT 304.950 515.400 340.050 516.450 ;
        RECT 304.950 514.950 307.050 515.400 ;
        RECT 337.950 514.950 340.050 515.400 ;
        RECT 343.950 516.450 346.050 517.050 ;
        RECT 356.400 516.450 357.450 518.400 ;
        RECT 373.950 517.950 376.050 518.400 ;
        RECT 388.950 517.950 391.050 518.400 ;
        RECT 550.950 519.450 553.050 520.050 ;
        RECT 580.950 519.450 583.050 519.900 ;
        RECT 550.950 518.400 583.050 519.450 ;
        RECT 550.950 517.950 553.050 518.400 ;
        RECT 580.950 517.800 583.050 518.400 ;
        RECT 637.950 519.450 640.050 520.050 ;
        RECT 676.950 519.450 679.050 523.050 ;
        RECT 706.950 520.950 712.050 523.050 ;
        RECT 637.950 519.000 679.050 519.450 ;
        RECT 691.950 519.450 694.050 520.050 ;
        RECT 715.950 519.450 718.050 523.050 ;
        RECT 728.850 521.400 730.050 533.400 ;
        RECT 739.950 531.450 744.000 532.050 ;
        RECT 739.950 531.000 744.450 531.450 ;
        RECT 739.950 529.950 745.050 531.000 ;
        RECT 733.950 526.950 739.050 529.050 ;
        RECT 742.950 526.950 745.050 529.950 ;
        RECT 691.950 519.000 718.050 519.450 ;
        RECT 727.950 519.300 730.050 521.400 ;
        RECT 637.950 518.400 678.450 519.000 ;
        RECT 691.950 518.400 717.450 519.000 ;
        RECT 637.950 517.950 640.050 518.400 ;
        RECT 691.950 517.950 694.050 518.400 ;
        RECT 343.950 515.400 357.450 516.450 ;
        RECT 415.950 516.450 418.050 517.050 ;
        RECT 424.950 516.450 427.050 517.050 ;
        RECT 415.950 515.400 427.050 516.450 ;
        RECT 343.950 514.950 346.050 515.400 ;
        RECT 415.950 514.950 418.050 515.400 ;
        RECT 424.950 514.950 427.050 515.400 ;
        RECT 514.950 516.450 517.050 517.050 ;
        RECT 583.950 516.450 586.050 517.050 ;
        RECT 514.950 515.400 586.050 516.450 ;
        RECT 514.950 514.950 517.050 515.400 ;
        RECT 583.950 514.950 586.050 515.400 ;
        RECT 592.950 516.450 595.050 517.050 ;
        RECT 664.950 516.450 667.050 517.050 ;
        RECT 592.950 515.400 667.050 516.450 ;
        RECT 592.950 514.950 595.050 515.400 ;
        RECT 664.950 514.950 667.050 515.400 ;
        RECT 670.950 516.450 673.050 517.200 ;
        RECT 685.950 516.450 688.050 517.050 ;
        RECT 670.950 515.400 688.050 516.450 ;
        RECT 728.850 515.700 730.050 519.300 ;
        RECT 749.100 516.600 750.300 533.400 ;
        RECT 856.950 532.950 859.050 533.400 ;
        RECT 757.950 531.450 760.050 532.050 ;
        RECT 784.950 531.450 787.050 532.050 ;
        RECT 805.950 531.450 808.050 532.050 ;
        RECT 757.950 530.400 808.050 531.450 ;
        RECT 757.950 529.950 760.050 530.400 ;
        RECT 766.950 526.950 769.050 530.400 ;
        RECT 784.950 529.950 787.050 530.400 ;
        RECT 805.950 529.950 808.050 530.400 ;
        RECT 778.950 528.450 781.050 529.050 ;
        RECT 784.800 528.450 786.900 529.050 ;
        RECT 778.950 527.400 786.900 528.450 ;
        RECT 778.950 526.950 781.050 527.400 ;
        RECT 784.800 526.950 786.900 527.400 ;
        RECT 788.100 526.950 793.050 529.050 ;
        RECT 754.950 525.450 757.050 526.050 ;
        RECT 763.950 525.450 766.050 526.050 ;
        RECT 754.950 524.400 766.050 525.450 ;
        RECT 754.950 523.950 757.050 524.400 ;
        RECT 763.950 523.950 766.050 524.400 ;
        RECT 769.950 522.450 772.050 526.050 ;
        RECT 784.950 523.950 790.050 526.050 ;
        RECT 787.950 522.450 790.050 523.050 ;
        RECT 769.950 522.000 790.050 522.450 ;
        RECT 793.950 522.450 796.050 526.050 ;
        RECT 811.950 525.450 814.050 526.050 ;
        RECT 820.950 525.450 823.050 529.050 ;
        RECT 826.950 526.950 829.050 532.050 ;
        RECT 811.950 525.000 823.050 525.450 ;
        RECT 811.950 524.400 822.450 525.000 ;
        RECT 811.950 523.950 814.050 524.400 ;
        RECT 823.950 523.050 826.050 526.050 ;
        RECT 844.950 525.450 847.050 526.050 ;
        RECT 853.950 525.450 856.050 526.050 ;
        RECT 844.950 524.400 856.050 525.450 ;
        RECT 844.950 523.950 847.050 524.400 ;
        RECT 853.950 523.950 856.050 524.400 ;
        RECT 805.950 522.450 808.050 523.050 ;
        RECT 820.950 522.450 826.050 523.050 ;
        RECT 793.950 522.000 826.050 522.450 ;
        RECT 770.400 521.400 790.050 522.000 ;
        RECT 794.400 521.400 825.450 522.000 ;
        RECT 787.950 520.950 790.050 521.400 ;
        RECT 805.950 520.950 808.050 521.400 ;
        RECT 820.950 520.950 825.000 521.400 ;
        RECT 670.950 515.100 673.050 515.400 ;
        RECT 685.950 514.950 688.050 515.400 ;
        RECT 253.950 513.450 256.050 514.050 ;
        RECT 331.800 513.450 333.900 514.050 ;
        RECT 253.950 512.400 333.900 513.450 ;
        RECT 253.950 511.950 256.050 512.400 ;
        RECT 331.800 511.950 333.900 512.400 ;
        RECT 335.100 513.450 337.200 514.050 ;
        RECT 343.950 513.450 346.050 514.050 ;
        RECT 335.100 512.400 346.050 513.450 ;
        RECT 335.100 511.950 337.200 512.400 ;
        RECT 343.950 511.950 346.050 512.400 ;
        RECT 472.950 513.450 475.050 514.050 ;
        RECT 484.950 513.450 487.050 514.050 ;
        RECT 472.950 512.400 487.050 513.450 ;
        RECT 472.950 511.950 475.050 512.400 ;
        RECT 484.950 511.950 487.050 512.400 ;
        RECT 670.950 513.450 673.050 513.900 ;
        RECT 727.950 513.600 730.050 515.700 ;
        RECT 748.950 514.500 751.050 516.600 ;
        RECT 760.950 516.450 763.050 517.050 ;
        RECT 793.950 516.450 796.050 517.050 ;
        RECT 760.950 515.400 796.050 516.450 ;
        RECT 760.950 514.950 763.050 515.400 ;
        RECT 793.950 514.950 796.050 515.400 ;
        RECT 832.950 513.450 835.050 514.050 ;
        RECT 844.950 513.450 847.050 514.050 ;
        RECT 670.950 512.400 714.450 513.450 ;
        RECT 670.950 511.800 673.050 512.400 ;
        RECT 28.950 510.450 31.050 511.050 ;
        RECT 151.950 510.450 154.050 511.050 ;
        RECT 28.950 509.400 154.050 510.450 ;
        RECT 28.950 508.950 31.050 509.400 ;
        RECT 151.950 508.950 154.050 509.400 ;
        RECT 220.950 510.450 223.050 511.050 ;
        RECT 343.950 510.450 346.050 511.050 ;
        RECT 220.950 509.400 346.050 510.450 ;
        RECT 220.950 508.950 223.050 509.400 ;
        RECT 343.950 508.950 346.050 509.400 ;
        RECT 460.950 510.450 463.050 511.050 ;
        RECT 550.950 510.450 553.050 511.050 ;
        RECT 583.950 510.450 586.050 511.050 ;
        RECT 604.950 510.450 607.050 511.050 ;
        RECT 460.950 509.400 607.050 510.450 ;
        RECT 460.950 508.950 463.050 509.400 ;
        RECT 550.950 508.950 553.050 509.400 ;
        RECT 583.950 508.950 586.050 509.400 ;
        RECT 604.950 508.950 607.050 509.400 ;
        RECT 619.950 510.450 622.050 511.050 ;
        RECT 709.950 510.450 712.050 511.050 ;
        RECT 619.950 509.400 712.050 510.450 ;
        RECT 713.400 510.450 714.450 512.400 ;
        RECT 832.950 512.400 847.050 513.450 ;
        RECT 832.950 511.950 835.050 512.400 ;
        RECT 844.950 511.950 847.050 512.400 ;
        RECT 745.950 510.450 748.050 511.050 ;
        RECT 713.400 509.400 748.050 510.450 ;
        RECT 619.950 508.950 622.050 509.400 ;
        RECT 709.950 508.950 712.050 509.400 ;
        RECT 745.950 508.950 748.050 509.400 ;
        RECT 778.950 510.450 781.050 511.050 ;
        RECT 793.950 510.450 796.050 511.050 ;
        RECT 778.950 509.400 796.050 510.450 ;
        RECT 778.950 508.950 781.050 509.400 ;
        RECT 793.950 508.950 796.050 509.400 ;
        RECT 841.950 510.450 844.050 511.050 ;
        RECT 853.950 510.450 856.050 511.050 ;
        RECT 841.950 509.400 856.050 510.450 ;
        RECT 841.950 508.950 844.050 509.400 ;
        RECT 853.950 508.950 856.050 509.400 ;
        RECT 214.950 507.450 217.050 508.050 ;
        RECT 277.950 507.450 280.050 508.050 ;
        RECT 214.950 506.400 280.050 507.450 ;
        RECT 214.950 505.950 217.050 506.400 ;
        RECT 277.950 505.950 280.050 506.400 ;
        RECT 295.950 507.450 298.050 508.050 ;
        RECT 337.950 507.450 340.050 508.050 ;
        RECT 295.950 506.400 340.050 507.450 ;
        RECT 295.950 505.950 298.050 506.400 ;
        RECT 337.950 505.950 340.050 506.400 ;
        RECT 376.950 507.450 379.050 508.050 ;
        RECT 406.950 507.450 409.050 508.050 ;
        RECT 376.950 506.400 409.050 507.450 ;
        RECT 376.950 505.950 379.050 506.400 ;
        RECT 406.950 505.950 409.050 506.400 ;
        RECT 511.950 507.450 514.050 508.050 ;
        RECT 598.950 507.450 601.050 508.050 ;
        RECT 616.950 507.450 619.050 508.050 ;
        RECT 511.950 506.400 601.050 507.450 ;
        RECT 511.950 505.950 514.050 506.400 ;
        RECT 598.950 505.950 601.050 506.400 ;
        RECT 605.400 506.400 619.050 507.450 ;
        RECT 16.950 504.450 19.050 505.050 ;
        RECT 115.950 504.450 118.050 505.050 ;
        RECT 124.950 504.450 127.050 505.050 ;
        RECT 136.950 504.450 139.050 505.050 ;
        RECT 16.950 503.400 139.050 504.450 ;
        RECT 16.950 502.950 19.050 503.400 ;
        RECT 115.950 502.950 118.050 503.400 ;
        RECT 124.950 502.950 127.050 503.400 ;
        RECT 136.950 502.950 139.050 503.400 ;
        RECT 172.950 504.450 175.050 505.050 ;
        RECT 280.950 504.450 283.050 505.050 ;
        RECT 172.950 503.400 283.050 504.450 ;
        RECT 172.950 502.950 175.050 503.400 ;
        RECT 280.950 502.950 283.050 503.400 ;
        RECT 298.950 504.450 301.050 505.050 ;
        RECT 445.950 504.450 448.050 505.050 ;
        RECT 298.950 503.400 448.050 504.450 ;
        RECT 298.950 502.950 301.050 503.400 ;
        RECT 445.950 502.950 448.050 503.400 ;
        RECT 472.950 504.450 475.050 505.050 ;
        RECT 505.950 504.450 508.050 505.200 ;
        RECT 472.950 503.400 508.050 504.450 ;
        RECT 472.950 502.950 475.050 503.400 ;
        RECT 505.950 503.100 508.050 503.400 ;
        RECT 577.950 504.450 580.050 505.050 ;
        RECT 605.400 504.450 606.450 506.400 ;
        RECT 616.950 505.950 619.050 506.400 ;
        RECT 685.950 507.450 688.050 508.050 ;
        RECT 754.950 507.450 757.050 508.050 ;
        RECT 778.950 507.450 781.050 508.050 ;
        RECT 685.950 506.400 781.050 507.450 ;
        RECT 685.950 505.950 688.050 506.400 ;
        RECT 754.950 505.950 757.050 506.400 ;
        RECT 778.950 505.950 781.050 506.400 ;
        RECT 634.950 504.450 637.050 505.050 ;
        RECT 577.950 503.400 606.450 504.450 ;
        RECT 608.400 503.400 637.050 504.450 ;
        RECT 577.950 502.950 580.050 503.400 ;
        RECT 199.950 501.450 202.050 502.050 ;
        RECT 232.950 501.450 235.050 502.050 ;
        RECT 199.950 500.400 235.050 501.450 ;
        RECT 199.950 499.950 202.050 500.400 ;
        RECT 232.950 499.950 235.050 500.400 ;
        RECT 259.950 501.450 262.050 502.050 ;
        RECT 313.950 501.450 319.050 502.050 ;
        RECT 259.950 500.400 319.050 501.450 ;
        RECT 259.950 499.950 262.050 500.400 ;
        RECT 313.950 499.950 319.050 500.400 ;
        RECT 343.950 501.450 346.050 502.050 ;
        RECT 406.950 501.450 409.050 502.050 ;
        RECT 343.950 500.400 409.050 501.450 ;
        RECT 343.950 499.950 346.050 500.400 ;
        RECT 406.950 499.950 409.050 500.400 ;
        RECT 415.950 501.450 418.050 502.050 ;
        RECT 439.950 501.450 442.050 502.050 ;
        RECT 415.950 500.400 442.050 501.450 ;
        RECT 415.950 499.950 418.050 500.400 ;
        RECT 439.950 499.950 442.050 500.400 ;
        RECT 505.950 501.450 508.050 501.900 ;
        RECT 517.950 501.450 520.050 502.050 ;
        RECT 505.950 500.400 520.050 501.450 ;
        RECT 67.950 498.450 70.050 499.050 ;
        RECT 106.950 498.450 109.050 499.050 ;
        RECT 127.950 498.450 130.050 499.050 ;
        RECT 67.950 497.400 105.450 498.450 ;
        RECT 67.950 496.950 70.050 497.400 ;
        RECT 70.950 495.450 73.050 496.050 ;
        RECT 79.950 495.450 82.050 496.050 ;
        RECT 70.950 494.400 82.050 495.450 ;
        RECT 104.400 495.450 105.450 497.400 ;
        RECT 106.950 497.400 130.050 498.450 ;
        RECT 106.950 496.950 109.050 497.400 ;
        RECT 127.950 496.950 130.050 497.400 ;
        RECT 184.950 498.450 187.050 499.050 ;
        RECT 295.950 498.450 298.050 499.050 ;
        RECT 367.950 498.450 370.050 499.050 ;
        RECT 184.950 497.400 294.450 498.450 ;
        RECT 184.950 496.950 187.050 497.400 ;
        RECT 169.950 495.450 172.050 496.050 ;
        RECT 104.400 494.400 172.050 495.450 ;
        RECT 70.950 493.950 73.050 494.400 ;
        RECT 79.950 493.950 82.050 494.400 ;
        RECT 169.950 493.950 172.050 494.400 ;
        RECT 220.950 495.450 223.050 496.050 ;
        RECT 241.950 495.450 244.050 496.050 ;
        RECT 259.950 495.450 262.050 496.050 ;
        RECT 220.950 494.400 244.050 495.450 ;
        RECT 220.950 493.950 223.050 494.400 ;
        RECT 241.950 493.950 244.050 494.400 ;
        RECT 251.400 494.400 262.050 495.450 ;
        RECT 293.400 495.450 294.450 497.400 ;
        RECT 295.950 497.400 370.050 498.450 ;
        RECT 407.400 498.450 408.450 499.950 ;
        RECT 505.950 499.800 508.050 500.400 ;
        RECT 517.950 499.950 520.050 500.400 ;
        RECT 556.950 501.450 559.050 502.050 ;
        RECT 608.400 501.450 609.450 503.400 ;
        RECT 634.950 502.950 637.050 503.400 ;
        RECT 655.950 504.450 658.050 505.050 ;
        RECT 691.950 504.450 694.050 505.050 ;
        RECT 655.950 503.400 694.050 504.450 ;
        RECT 655.950 502.950 658.050 503.400 ;
        RECT 691.950 502.950 694.050 503.400 ;
        RECT 712.950 504.450 715.050 505.050 ;
        RECT 730.950 504.450 733.050 505.050 ;
        RECT 712.950 503.400 733.050 504.450 ;
        RECT 712.950 502.950 715.050 503.400 ;
        RECT 730.950 502.950 733.050 503.400 ;
        RECT 739.950 504.450 742.050 505.050 ;
        RECT 829.950 504.450 832.050 505.050 ;
        RECT 739.950 503.400 832.050 504.450 ;
        RECT 739.950 502.950 742.050 503.400 ;
        RECT 829.950 502.950 832.050 503.400 ;
        RECT 556.950 500.400 609.450 501.450 ;
        RECT 610.950 501.450 613.050 502.050 ;
        RECT 772.950 501.450 775.050 502.050 ;
        RECT 610.950 500.400 775.050 501.450 ;
        RECT 556.950 499.950 559.050 500.400 ;
        RECT 610.950 499.950 613.050 500.400 ;
        RECT 772.950 499.950 775.050 500.400 ;
        RECT 421.950 498.450 424.050 499.050 ;
        RECT 407.400 497.400 424.050 498.450 ;
        RECT 604.950 498.450 607.050 499.050 ;
        RECT 658.800 498.450 660.900 499.050 ;
        RECT 604.950 497.400 660.900 498.450 ;
        RECT 295.950 496.950 298.050 497.400 ;
        RECT 367.950 496.950 370.050 497.400 ;
        RECT 421.950 496.950 424.050 497.400 ;
        RECT 328.950 495.450 331.050 496.050 ;
        RECT 364.950 495.450 367.050 496.050 ;
        RECT 293.400 494.400 367.050 495.450 ;
        RECT 10.950 492.450 13.050 493.050 ;
        RECT 34.950 492.450 37.050 493.050 ;
        RECT 73.950 492.450 76.050 493.050 ;
        RECT 10.950 491.400 37.050 492.450 ;
        RECT 10.950 490.950 13.050 491.400 ;
        RECT 17.400 487.050 18.450 491.400 ;
        RECT 34.950 490.950 37.050 491.400 ;
        RECT 59.400 491.400 76.050 492.450 ;
        RECT 49.800 489.000 51.900 490.050 ;
        RECT 53.100 489.450 55.200 490.050 ;
        RECT 59.400 489.450 60.450 491.400 ;
        RECT 73.950 490.950 76.050 491.400 ;
        RECT 49.800 487.950 52.050 489.000 ;
        RECT 53.100 488.400 60.450 489.450 ;
        RECT 61.950 489.450 64.050 490.050 ;
        RECT 61.950 488.400 75.450 489.450 ;
        RECT 53.100 487.950 55.200 488.400 ;
        RECT 61.950 487.950 64.050 488.400 ;
        RECT 7.950 484.950 13.050 487.050 ;
        RECT 16.950 484.950 19.050 487.050 ;
        RECT 28.800 486.000 30.900 487.050 ;
        RECT 28.800 484.950 31.050 486.000 ;
        RECT 32.100 484.950 36.900 487.050 ;
        RECT 38.100 486.450 40.200 487.050 ;
        RECT 43.950 486.450 46.050 487.050 ;
        RECT 38.100 485.400 46.050 486.450 ;
        RECT 38.100 484.950 40.200 485.400 ;
        RECT 43.950 484.950 46.050 485.400 ;
        RECT 49.950 484.950 52.050 487.950 ;
        RECT 74.400 487.050 75.450 488.400 ;
        RECT 79.950 487.950 82.050 493.050 ;
        RECT 106.950 492.450 109.050 493.050 ;
        RECT 151.950 492.450 154.050 493.050 ;
        RECT 106.950 491.400 154.050 492.450 ;
        RECT 106.950 490.950 109.050 491.400 ;
        RECT 151.950 490.950 154.050 491.400 ;
        RECT 196.950 492.450 201.000 493.050 ;
        RECT 196.950 490.950 201.450 492.450 ;
        RECT 175.950 490.050 178.050 490.200 ;
        RECT 13.950 481.950 18.900 484.050 ;
        RECT 20.100 483.450 22.200 484.050 ;
        RECT 28.950 483.450 31.050 484.950 ;
        RECT 20.100 482.400 31.050 483.450 ;
        RECT 20.100 481.950 22.200 482.400 ;
        RECT 28.950 481.950 31.050 482.400 ;
        RECT 34.950 483.450 37.050 484.050 ;
        RECT 34.950 482.400 54.450 483.450 ;
        RECT 34.950 481.950 37.050 482.400 ;
        RECT 53.400 480.450 54.450 482.400 ;
        RECT 55.950 481.950 58.050 487.050 ;
        RECT 74.400 485.400 79.050 487.050 ;
        RECT 75.000 484.950 79.050 485.400 ;
        RECT 82.800 486.000 84.900 487.050 ;
        RECT 86.100 486.450 88.200 487.050 ;
        RECT 91.800 486.450 93.900 487.050 ;
        RECT 82.800 484.950 85.050 486.000 ;
        RECT 86.100 485.400 93.900 486.450 ;
        RECT 86.100 484.950 88.200 485.400 ;
        RECT 91.800 484.950 93.900 485.400 ;
        RECT 95.100 486.450 100.050 487.050 ;
        RECT 112.950 486.450 115.050 487.050 ;
        RECT 95.100 485.400 115.050 486.450 ;
        RECT 95.100 484.950 100.050 485.400 ;
        RECT 112.950 484.950 115.050 485.400 ;
        RECT 124.950 484.950 130.050 487.050 ;
        RECT 133.950 484.950 136.050 490.050 ;
        RECT 151.950 484.950 154.050 490.050 ;
        RECT 169.800 489.000 171.900 490.050 ;
        RECT 169.800 487.950 172.050 489.000 ;
        RECT 173.100 488.100 178.050 490.050 ;
        RECT 173.100 487.950 177.000 488.100 ;
        RECT 157.950 486.450 160.050 487.050 ;
        RECT 163.950 486.450 166.050 487.050 ;
        RECT 157.950 485.400 166.050 486.450 ;
        RECT 157.950 484.950 160.050 485.400 ;
        RECT 163.950 484.950 166.050 485.400 ;
        RECT 169.950 484.950 172.050 487.950 ;
        RECT 200.400 487.050 201.450 490.950 ;
        RECT 208.950 489.450 211.050 490.050 ;
        RECT 244.950 489.450 247.050 490.050 ;
        RECT 208.950 488.400 247.050 489.450 ;
        RECT 208.950 487.950 211.050 488.400 ;
        RECT 244.950 487.950 247.050 488.400 ;
        RECT 251.400 487.050 252.450 494.400 ;
        RECT 259.950 493.950 262.050 494.400 ;
        RECT 328.950 493.950 331.050 494.400 ;
        RECT 364.950 493.950 367.050 494.400 ;
        RECT 409.950 495.450 412.050 496.050 ;
        RECT 424.950 495.450 427.050 496.050 ;
        RECT 409.950 494.400 427.050 495.450 ;
        RECT 541.950 495.300 544.050 497.400 ;
        RECT 409.950 493.950 412.050 494.400 ;
        RECT 424.950 493.950 427.050 494.400 ;
        RECT 253.800 492.000 255.900 493.050 ;
        RECT 257.100 492.450 259.200 493.050 ;
        RECT 268.950 492.450 271.050 493.050 ;
        RECT 253.800 490.950 256.050 492.000 ;
        RECT 257.100 491.400 271.050 492.450 ;
        RECT 257.100 490.950 259.200 491.400 ;
        RECT 268.950 490.950 271.050 491.400 ;
        RECT 253.950 487.950 256.050 490.950 ;
        RECT 259.950 489.450 262.050 490.050 ;
        RECT 265.950 489.450 268.050 490.050 ;
        RECT 259.950 488.400 268.050 489.450 ;
        RECT 259.950 487.950 262.050 488.400 ;
        RECT 265.950 487.950 268.050 488.400 ;
        RECT 283.950 487.950 289.050 490.050 ;
        RECT 292.950 489.450 298.050 490.050 ;
        RECT 301.950 489.450 304.050 490.050 ;
        RECT 292.950 488.400 304.050 489.450 ;
        RECT 292.950 487.950 298.050 488.400 ;
        RECT 301.950 487.950 304.050 488.400 ;
        RECT 307.950 487.950 313.050 490.050 ;
        RECT 316.950 489.450 319.050 490.050 ;
        RECT 322.950 489.450 325.050 490.050 ;
        RECT 316.950 488.400 325.050 489.450 ;
        RECT 316.950 487.950 319.050 488.400 ;
        RECT 322.950 487.950 325.050 488.400 ;
        RECT 328.950 487.950 331.050 493.050 ;
        RECT 340.950 492.450 343.050 493.050 ;
        RECT 394.950 492.450 397.050 493.050 ;
        RECT 418.950 492.450 421.050 493.050 ;
        RECT 448.950 492.450 451.050 493.050 ;
        RECT 340.950 492.000 360.450 492.450 ;
        RECT 340.950 491.400 361.050 492.000 ;
        RECT 340.950 490.950 343.050 491.400 ;
        RECT 337.950 487.950 342.900 490.050 ;
        RECT 343.800 489.000 345.900 490.050 ;
        RECT 347.100 489.450 351.000 490.050 ;
        RECT 343.800 487.950 346.050 489.000 ;
        RECT 347.100 487.950 351.450 489.450 ;
        RECT 358.950 487.950 361.050 491.400 ;
        RECT 394.950 491.400 451.050 492.450 ;
        RECT 394.950 490.950 397.050 491.400 ;
        RECT 418.950 490.950 421.050 491.400 ;
        RECT 448.950 490.950 451.050 491.400 ;
        RECT 454.950 492.450 457.050 493.050 ;
        RECT 535.950 492.450 538.050 493.050 ;
        RECT 454.950 491.400 538.050 492.450 ;
        RECT 542.850 491.700 544.050 495.300 ;
        RECT 562.950 494.400 565.050 496.500 ;
        RECT 577.950 495.300 580.050 497.400 ;
        RECT 604.950 496.950 607.050 497.400 ;
        RECT 658.800 496.950 660.900 497.400 ;
        RECT 688.950 498.450 691.050 499.050 ;
        RECT 739.950 498.450 742.050 499.050 ;
        RECT 688.950 497.400 742.050 498.450 ;
        RECT 688.950 496.950 691.050 497.400 ;
        RECT 739.950 496.950 742.050 497.400 ;
        RECT 781.950 498.450 784.050 499.050 ;
        RECT 787.950 498.450 790.050 499.050 ;
        RECT 781.950 497.400 790.050 498.450 ;
        RECT 781.950 496.950 784.050 497.400 ;
        RECT 787.950 496.950 790.050 497.400 ;
        RECT 454.950 490.950 457.050 491.400 ;
        RECT 535.950 490.950 538.050 491.400 ;
        RECT 367.950 489.450 370.050 490.050 ;
        RECT 367.950 489.000 378.450 489.450 ;
        RECT 367.950 488.400 379.050 489.000 ;
        RECT 367.950 487.950 370.050 488.400 ;
        RECT 343.950 487.050 346.050 487.950 ;
        RECT 350.400 487.050 351.450 487.950 ;
        RECT 175.950 484.950 181.050 487.050 ;
        RECT 190.950 484.950 196.050 487.050 ;
        RECT 199.950 484.950 202.050 487.050 ;
        RECT 211.950 486.450 214.050 487.050 ;
        RECT 206.400 485.400 214.050 486.450 ;
        RECT 82.950 483.450 85.050 484.950 ;
        RECT 206.400 484.050 207.450 485.400 ;
        RECT 211.950 484.950 214.050 485.400 ;
        RECT 250.950 484.950 253.050 487.050 ;
        RECT 256.950 486.450 259.050 487.050 ;
        RECT 265.950 486.450 268.050 487.050 ;
        RECT 256.950 485.400 268.050 486.450 ;
        RECT 256.950 484.950 259.050 485.400 ;
        RECT 265.950 484.950 268.050 485.400 ;
        RECT 286.950 484.950 292.050 487.050 ;
        RECT 304.950 486.450 307.050 487.050 ;
        RECT 316.950 486.450 319.050 487.050 ;
        RECT 304.950 485.400 319.050 486.450 ;
        RECT 304.950 484.950 307.050 485.400 ;
        RECT 316.950 484.950 319.050 485.400 ;
        RECT 91.800 483.450 93.900 484.050 ;
        RECT 82.950 483.000 93.900 483.450 ;
        RECT 95.100 483.000 97.200 484.050 ;
        RECT 83.250 482.400 93.900 483.000 ;
        RECT 91.800 481.950 93.900 482.400 ;
        RECT 94.950 481.950 97.200 483.000 ;
        RECT 124.950 483.450 127.050 484.050 ;
        RECT 130.950 483.450 133.050 484.050 ;
        RECT 124.950 482.400 133.050 483.450 ;
        RECT 124.950 481.950 127.050 482.400 ;
        RECT 130.950 481.950 133.050 482.400 ;
        RECT 139.950 483.450 142.050 484.050 ;
        RECT 148.950 483.450 151.050 484.050 ;
        RECT 139.950 482.400 151.050 483.450 ;
        RECT 139.950 481.950 142.050 482.400 ;
        RECT 148.950 481.950 151.050 482.400 ;
        RECT 154.800 483.000 156.900 484.050 ;
        RECT 158.100 483.450 160.200 484.050 ;
        RECT 196.950 483.450 199.050 484.050 ;
        RECT 154.800 481.950 157.050 483.000 ;
        RECT 158.100 482.400 199.050 483.450 ;
        RECT 158.100 481.950 160.200 482.400 ;
        RECT 196.950 481.950 199.050 482.400 ;
        RECT 202.950 482.400 207.450 484.050 ;
        RECT 226.950 483.450 229.050 484.050 ;
        RECT 235.800 483.450 237.900 484.050 ;
        RECT 218.400 483.000 237.900 483.450 ;
        RECT 217.950 482.400 237.900 483.000 ;
        RECT 202.950 481.950 207.000 482.400 ;
        RECT 70.950 480.450 73.050 481.050 ;
        RECT 94.950 480.450 97.050 481.950 ;
        RECT 53.400 480.000 97.050 480.450 ;
        RECT 118.950 480.450 121.050 481.050 ;
        RECT 127.950 480.450 130.050 481.050 ;
        RECT 133.950 480.450 136.050 481.050 ;
        RECT 53.400 479.400 96.600 480.000 ;
        RECT 118.950 479.400 136.050 480.450 ;
        RECT 154.950 480.450 157.050 481.950 ;
        RECT 187.950 480.450 190.050 481.050 ;
        RECT 154.950 480.000 190.050 480.450 ;
        RECT 155.400 479.400 190.050 480.000 ;
        RECT 70.950 478.950 73.050 479.400 ;
        RECT 118.950 478.950 121.050 479.400 ;
        RECT 127.950 478.950 130.050 479.400 ;
        RECT 133.950 478.950 136.050 479.400 ;
        RECT 187.950 478.950 190.050 479.400 ;
        RECT 193.950 480.450 196.050 481.050 ;
        RECT 202.950 480.450 205.050 481.050 ;
        RECT 193.950 479.400 205.050 480.450 ;
        RECT 193.950 478.950 196.050 479.400 ;
        RECT 202.950 478.950 205.050 479.400 ;
        RECT 217.950 478.950 220.050 482.400 ;
        RECT 226.950 481.950 229.050 482.400 ;
        RECT 235.800 481.950 237.900 482.400 ;
        RECT 239.100 483.450 241.200 484.050 ;
        RECT 247.950 483.450 250.050 484.050 ;
        RECT 239.100 482.400 250.050 483.450 ;
        RECT 239.100 481.950 241.200 482.400 ;
        RECT 247.950 481.950 250.050 482.400 ;
        RECT 280.950 483.450 283.050 484.050 ;
        RECT 295.950 483.450 298.050 484.050 ;
        RECT 280.950 482.400 298.050 483.450 ;
        RECT 280.950 481.950 283.050 482.400 ;
        RECT 295.950 481.950 298.050 482.400 ;
        RECT 325.950 481.950 328.050 487.050 ;
        RECT 343.800 486.000 346.050 487.050 ;
        RECT 349.950 486.450 352.050 487.050 ;
        RECT 355.950 486.450 358.050 487.050 ;
        RECT 343.800 484.950 345.900 486.000 ;
        RECT 349.950 485.400 358.050 486.450 ;
        RECT 349.950 484.950 352.050 485.400 ;
        RECT 355.950 484.950 358.050 485.400 ;
        RECT 361.950 481.950 364.050 487.050 ;
        RECT 376.950 484.950 379.050 488.400 ;
        RECT 382.950 484.950 388.050 487.050 ;
        RECT 397.950 484.950 403.050 487.050 ;
        RECT 406.950 484.950 409.050 490.050 ;
        RECT 436.950 486.450 439.050 487.050 ;
        RECT 428.400 486.000 439.050 486.450 ;
        RECT 427.950 485.400 439.050 486.000 ;
        RECT 166.950 477.450 169.050 478.050 ;
        RECT 190.950 477.450 193.050 478.050 ;
        RECT 166.950 476.400 193.050 477.450 ;
        RECT 271.950 477.450 274.050 481.050 ;
        RECT 322.950 480.450 325.050 481.050 ;
        RECT 355.950 480.450 358.050 481.050 ;
        RECT 322.950 479.400 358.050 480.450 ;
        RECT 379.950 480.450 382.050 484.050 ;
        RECT 394.950 483.450 397.050 484.050 ;
        RECT 403.950 483.450 406.050 484.050 ;
        RECT 394.950 482.400 406.050 483.450 ;
        RECT 394.950 481.950 397.050 482.400 ;
        RECT 403.950 481.950 406.050 482.400 ;
        RECT 397.950 480.450 400.050 481.050 ;
        RECT 379.950 480.000 400.050 480.450 ;
        RECT 380.400 479.400 400.050 480.000 ;
        RECT 322.950 478.950 325.050 479.400 ;
        RECT 355.950 478.950 358.050 479.400 ;
        RECT 397.950 478.950 400.050 479.400 ;
        RECT 409.950 478.950 412.050 484.050 ;
        RECT 418.950 481.950 424.050 484.050 ;
        RECT 427.950 483.450 430.050 485.400 ;
        RECT 436.950 484.950 439.050 485.400 ;
        RECT 448.950 484.950 454.050 487.050 ;
        RECT 457.950 486.450 460.050 490.050 ;
        RECT 463.950 489.450 466.050 490.050 ;
        RECT 481.950 489.450 487.050 490.050 ;
        RECT 541.950 489.600 544.050 491.700 ;
        RECT 463.950 488.400 487.050 489.450 ;
        RECT 463.950 487.950 466.050 488.400 ;
        RECT 481.950 487.950 487.050 488.400 ;
        RECT 487.950 486.450 490.050 487.050 ;
        RECT 493.950 486.450 496.050 487.050 ;
        RECT 457.950 485.400 477.450 486.450 ;
        RECT 457.950 484.950 460.050 485.400 ;
        RECT 454.950 483.450 457.050 484.050 ;
        RECT 427.950 482.400 457.050 483.450 ;
        RECT 427.950 481.950 430.050 482.400 ;
        RECT 454.950 481.950 457.050 482.400 ;
        RECT 463.950 483.450 466.050 484.050 ;
        RECT 469.950 483.450 472.050 484.050 ;
        RECT 476.400 483.900 477.450 485.400 ;
        RECT 487.950 485.400 496.050 486.450 ;
        RECT 487.950 484.950 490.050 485.400 ;
        RECT 493.950 484.950 496.050 485.400 ;
        RECT 511.950 484.950 517.050 487.050 ;
        RECT 520.950 484.950 526.050 487.050 ;
        RECT 463.950 482.400 472.050 483.450 ;
        RECT 463.950 481.950 466.050 482.400 ;
        RECT 469.950 481.950 472.050 482.400 ;
        RECT 475.950 481.800 478.050 483.900 ;
        RECT 514.950 481.950 520.050 484.050 ;
        RECT 526.950 483.450 529.050 484.050 ;
        RECT 521.400 482.400 529.050 483.450 ;
        RECT 415.950 480.450 418.050 481.050 ;
        RECT 424.950 480.450 427.050 481.050 ;
        RECT 415.950 479.400 427.050 480.450 ;
        RECT 415.950 478.950 418.050 479.400 ;
        RECT 424.950 478.950 427.050 479.400 ;
        RECT 433.950 480.450 436.050 481.050 ;
        RECT 442.950 480.450 445.050 481.050 ;
        RECT 433.950 479.400 445.050 480.450 ;
        RECT 433.950 478.950 436.050 479.400 ;
        RECT 442.950 478.950 445.050 479.400 ;
        RECT 274.950 477.450 277.050 478.050 ;
        RECT 352.950 477.450 355.050 478.050 ;
        RECT 271.950 477.000 355.050 477.450 ;
        RECT 272.400 476.400 355.050 477.000 ;
        RECT 166.950 475.950 169.050 476.400 ;
        RECT 190.950 475.950 193.050 476.400 ;
        RECT 274.950 475.950 277.050 476.400 ;
        RECT 352.950 475.950 355.050 476.400 ;
        RECT 361.950 477.450 364.050 478.050 ;
        RECT 415.950 477.450 421.050 478.050 ;
        RECT 361.950 476.400 421.050 477.450 ;
        RECT 361.950 475.950 364.050 476.400 ;
        RECT 415.950 475.950 421.050 476.400 ;
        RECT 484.950 475.950 487.050 481.050 ;
        RECT 511.950 480.450 514.050 481.050 ;
        RECT 517.950 480.450 520.050 481.050 ;
        RECT 521.400 480.450 522.450 482.400 ;
        RECT 526.950 481.950 529.050 482.400 ;
        RECT 535.950 481.950 541.050 484.050 ;
        RECT 511.950 479.400 522.450 480.450 ;
        RECT 511.950 478.950 514.050 479.400 ;
        RECT 517.950 478.950 520.050 479.400 ;
        RECT 505.950 477.450 508.050 478.050 ;
        RECT 511.950 477.450 514.050 478.050 ;
        RECT 542.850 477.600 544.050 489.600 ;
        RECT 557.100 486.000 559.200 487.050 ;
        RECT 556.950 484.950 559.200 486.000 ;
        RECT 556.950 484.050 559.050 484.950 ;
        RECT 550.950 481.950 555.900 484.050 ;
        RECT 556.950 483.000 559.200 484.050 ;
        RECT 557.100 481.950 559.200 483.000 ;
        RECT 563.100 477.600 564.300 494.400 ;
        RECT 578.850 491.700 580.050 495.300 ;
        RECT 598.950 494.400 601.050 496.500 ;
        RECT 613.950 495.450 616.050 496.050 ;
        RECT 637.950 495.450 640.050 496.050 ;
        RECT 613.950 494.400 640.050 495.450 ;
        RECT 577.950 489.600 580.050 491.700 ;
        RECT 565.950 483.450 568.050 484.050 ;
        RECT 574.950 483.450 577.050 484.050 ;
        RECT 565.950 482.400 577.050 483.450 ;
        RECT 565.950 481.950 568.050 482.400 ;
        RECT 574.950 481.950 577.050 482.400 ;
        RECT 578.850 477.600 580.050 489.600 ;
        RECT 583.950 481.950 589.050 484.050 ;
        RECT 592.950 481.950 595.050 487.050 ;
        RECT 599.100 477.600 600.300 494.400 ;
        RECT 613.950 493.950 616.050 494.400 ;
        RECT 637.950 493.950 640.050 494.400 ;
        RECT 649.950 495.450 652.050 496.050 ;
        RECT 655.950 495.450 658.050 496.050 ;
        RECT 679.950 495.450 682.050 496.050 ;
        RECT 649.950 494.400 682.050 495.450 ;
        RECT 649.950 493.950 652.050 494.400 ;
        RECT 655.950 493.950 658.050 494.400 ;
        RECT 679.950 493.950 682.050 494.400 ;
        RECT 698.100 495.450 700.200 496.050 ;
        RECT 709.950 495.450 712.050 496.050 ;
        RECT 698.100 494.400 712.050 495.450 ;
        RECT 698.100 493.950 700.200 494.400 ;
        RECT 709.950 493.950 712.050 494.400 ;
        RECT 721.950 495.450 724.050 496.050 ;
        RECT 727.950 495.450 730.050 496.050 ;
        RECT 721.950 494.400 730.050 495.450 ;
        RECT 721.950 493.950 724.050 494.400 ;
        RECT 727.950 493.950 730.050 494.400 ;
        RECT 784.950 495.450 787.050 496.050 ;
        RECT 835.950 495.450 838.050 496.050 ;
        RECT 784.950 494.400 838.050 495.450 ;
        RECT 784.950 493.950 787.050 494.400 ;
        RECT 835.950 493.950 838.050 494.400 ;
        RECT 643.950 492.450 646.050 493.050 ;
        RECT 718.950 492.450 721.050 493.050 ;
        RECT 736.950 492.450 739.050 493.050 ;
        RECT 643.950 491.400 672.450 492.450 ;
        RECT 643.950 490.950 646.050 491.400 ;
        RECT 671.400 490.050 672.450 491.400 ;
        RECT 718.950 491.400 739.050 492.450 ;
        RECT 718.950 490.950 721.050 491.400 ;
        RECT 736.950 490.950 739.050 491.400 ;
        RECT 745.950 492.450 748.050 493.050 ;
        RECT 760.950 492.450 766.050 493.050 ;
        RECT 745.950 491.400 766.050 492.450 ;
        RECT 745.950 490.950 748.050 491.400 ;
        RECT 760.950 490.950 766.050 491.400 ;
        RECT 613.950 487.950 619.050 490.050 ;
        RECT 622.950 487.950 628.050 490.050 ;
        RECT 619.950 483.450 622.050 487.050 ;
        RECT 633.000 486.450 636.900 487.050 ;
        RECT 632.400 484.950 636.900 486.450 ;
        RECT 638.100 484.950 643.050 487.050 ;
        RECT 655.950 484.950 661.050 487.050 ;
        RECT 670.950 484.950 673.050 490.050 ;
        RECT 691.950 489.450 694.050 490.050 ;
        RECT 697.950 489.450 700.050 490.050 ;
        RECT 691.950 488.400 700.050 489.450 ;
        RECT 691.950 487.950 694.050 488.400 ;
        RECT 697.950 487.950 700.050 488.400 ;
        RECT 709.950 487.950 715.050 490.050 ;
        RECT 682.950 486.450 685.050 487.050 ;
        RECT 688.950 486.450 691.050 487.050 ;
        RECT 682.950 485.400 691.050 486.450 ;
        RECT 682.950 484.950 685.050 485.400 ;
        RECT 688.950 484.950 691.050 485.400 ;
        RECT 706.950 484.950 712.050 487.050 ;
        RECT 718.950 484.950 724.050 487.050 ;
        RECT 727.950 486.450 730.050 487.050 ;
        RECT 739.950 486.450 742.050 487.050 ;
        RECT 727.950 485.400 742.050 486.450 ;
        RECT 727.950 484.950 730.050 485.400 ;
        RECT 739.950 484.950 742.050 485.400 ;
        RECT 745.950 484.950 748.050 490.050 ;
        RECT 772.950 489.450 775.050 490.050 ;
        RECT 793.950 489.450 796.050 490.050 ;
        RECT 814.950 489.450 817.050 490.050 ;
        RECT 772.950 489.000 801.450 489.450 ;
        RECT 806.400 489.000 817.050 489.450 ;
        RECT 772.950 488.400 802.050 489.000 ;
        RECT 772.950 487.950 775.050 488.400 ;
        RECT 793.950 487.950 796.050 488.400 ;
        RECT 751.950 486.450 754.050 487.050 ;
        RECT 760.950 486.450 763.050 487.050 ;
        RECT 799.950 486.450 802.050 488.400 ;
        RECT 751.950 485.400 763.050 486.450 ;
        RECT 788.400 486.000 802.050 486.450 ;
        RECT 751.950 484.950 754.050 485.400 ;
        RECT 760.950 484.950 763.050 485.400 ;
        RECT 787.950 485.400 802.050 486.000 ;
        RECT 632.400 483.450 633.450 484.950 ;
        RECT 619.950 483.000 633.450 483.450 ;
        RECT 620.400 482.400 633.450 483.000 ;
        RECT 634.950 481.950 640.050 484.050 ;
        RECT 643.950 481.950 649.050 484.050 ;
        RECT 715.950 481.950 721.050 484.050 ;
        RECT 723.000 483.450 727.050 484.050 ;
        RECT 722.400 481.950 727.050 483.450 ;
        RECT 697.950 480.450 700.050 481.050 ;
        RECT 722.400 480.450 723.450 481.950 ;
        RECT 697.950 479.400 723.450 480.450 ;
        RECT 730.950 480.450 733.050 484.050 ;
        RECT 736.950 483.450 739.050 484.050 ;
        RECT 748.950 483.450 751.050 484.050 ;
        RECT 736.950 482.400 751.050 483.450 ;
        RECT 736.950 481.950 739.050 482.400 ;
        RECT 748.950 481.950 751.050 482.400 ;
        RECT 754.950 481.950 760.050 484.050 ;
        RECT 778.950 481.950 784.050 484.050 ;
        RECT 787.950 481.950 790.050 485.400 ;
        RECT 799.950 484.950 802.050 485.400 ;
        RECT 805.950 488.400 817.050 489.000 ;
        RECT 805.950 484.950 808.050 488.400 ;
        RECT 814.950 487.950 817.050 488.400 ;
        RECT 820.950 486.450 823.050 487.050 ;
        RECT 812.400 485.400 823.050 486.450 ;
        RECT 793.950 481.950 799.050 484.050 ;
        RECT 802.950 483.450 805.050 484.050 ;
        RECT 812.400 483.450 813.450 485.400 ;
        RECT 820.950 484.950 823.050 485.400 ;
        RECT 826.950 486.450 829.050 490.050 ;
        RECT 826.950 486.000 843.600 486.450 ;
        RECT 826.950 485.400 844.050 486.000 ;
        RECT 826.950 484.950 829.050 485.400 ;
        RECT 841.950 484.050 844.050 485.400 ;
        RECT 823.950 483.450 826.050 484.050 ;
        RECT 802.950 482.400 813.450 483.450 ;
        RECT 815.400 482.400 826.050 483.450 ;
        RECT 841.950 483.000 844.200 484.050 ;
        RECT 802.950 481.950 805.050 482.400 ;
        RECT 815.400 481.050 816.450 482.400 ;
        RECT 823.950 481.950 826.050 482.400 ;
        RECT 842.100 481.950 844.200 483.000 ;
        RECT 760.950 480.450 763.050 481.050 ;
        RECT 730.950 480.000 763.050 480.450 ;
        RECT 731.400 479.400 763.050 480.000 ;
        RECT 697.950 478.950 700.050 479.400 ;
        RECT 760.950 478.950 763.050 479.400 ;
        RECT 769.950 478.950 775.050 481.050 ;
        RECT 784.950 480.450 787.050 481.050 ;
        RECT 802.950 480.450 805.050 481.050 ;
        RECT 784.950 479.400 805.050 480.450 ;
        RECT 784.950 478.950 787.050 479.400 ;
        RECT 802.950 478.950 805.050 479.400 ;
        RECT 811.950 479.400 816.450 481.050 ;
        RECT 829.950 480.450 832.050 481.050 ;
        RECT 844.950 480.450 847.050 481.050 ;
        RECT 829.950 479.400 847.050 480.450 ;
        RECT 811.950 478.950 816.000 479.400 ;
        RECT 829.950 478.950 832.050 479.400 ;
        RECT 844.950 478.950 847.050 479.400 ;
        RECT 505.950 476.400 514.050 477.450 ;
        RECT 505.950 475.950 508.050 476.400 ;
        RECT 511.950 475.950 514.050 476.400 ;
        RECT 541.950 475.500 544.050 477.600 ;
        RECT 562.950 475.500 565.050 477.600 ;
        RECT 577.950 475.500 580.050 477.600 ;
        RECT 598.950 475.500 601.050 477.600 ;
        RECT 646.950 477.450 649.050 478.050 ;
        RECT 664.950 477.450 667.050 478.050 ;
        RECT 646.950 476.400 667.050 477.450 ;
        RECT 646.950 475.950 649.050 476.400 ;
        RECT 664.950 475.950 667.050 476.400 ;
        RECT 676.950 477.450 679.050 478.050 ;
        RECT 718.950 477.450 721.050 478.050 ;
        RECT 676.950 476.400 721.050 477.450 ;
        RECT 676.950 475.950 679.050 476.400 ;
        RECT 718.950 475.950 721.050 476.400 ;
        RECT 766.950 477.450 769.050 478.050 ;
        RECT 766.950 476.400 774.450 477.450 ;
        RECT 766.950 475.950 769.050 476.400 ;
        RECT 163.950 474.450 166.050 475.050 ;
        RECT 178.950 474.450 181.050 475.050 ;
        RECT 163.950 473.400 181.050 474.450 ;
        RECT 163.950 472.950 166.050 473.400 ;
        RECT 178.950 472.950 181.050 473.400 ;
        RECT 187.950 474.450 190.050 475.050 ;
        RECT 286.950 474.450 289.050 475.050 ;
        RECT 319.950 474.450 322.050 475.050 ;
        RECT 187.950 473.400 258.450 474.450 ;
        RECT 187.950 472.950 190.050 473.400 ;
        RECT 28.950 471.450 31.050 472.050 ;
        RECT 208.950 471.450 211.050 472.050 ;
        RECT 28.950 470.400 211.050 471.450 ;
        RECT 257.400 471.450 258.450 473.400 ;
        RECT 286.950 473.400 322.050 474.450 ;
        RECT 286.950 472.950 289.050 473.400 ;
        RECT 319.950 472.950 322.050 473.400 ;
        RECT 349.950 474.450 352.050 475.050 ;
        RECT 355.950 474.450 358.050 475.050 ;
        RECT 349.950 473.400 358.050 474.450 ;
        RECT 349.950 472.950 352.050 473.400 ;
        RECT 355.950 472.950 358.050 473.400 ;
        RECT 391.950 474.450 394.050 475.050 ;
        RECT 427.950 474.450 430.050 475.050 ;
        RECT 484.950 474.450 487.050 475.050 ;
        RECT 391.950 473.400 487.050 474.450 ;
        RECT 391.950 472.950 394.050 473.400 ;
        RECT 427.950 472.950 430.050 473.400 ;
        RECT 484.950 472.950 487.050 473.400 ;
        RECT 643.950 474.450 646.050 475.050 ;
        RECT 673.950 474.450 676.050 475.050 ;
        RECT 643.950 473.400 676.050 474.450 ;
        RECT 643.950 472.950 646.050 473.400 ;
        RECT 673.950 472.950 676.050 473.400 ;
        RECT 727.950 474.450 730.050 475.050 ;
        RECT 769.950 474.450 772.050 475.050 ;
        RECT 727.950 473.400 772.050 474.450 ;
        RECT 773.400 474.450 774.450 476.400 ;
        RECT 808.950 474.450 811.050 475.050 ;
        RECT 773.400 473.400 811.050 474.450 ;
        RECT 727.950 472.950 730.050 473.400 ;
        RECT 769.950 472.950 772.050 473.400 ;
        RECT 808.950 472.950 811.050 473.400 ;
        RECT 826.950 474.450 829.050 475.050 ;
        RECT 841.950 474.450 844.050 475.050 ;
        RECT 826.950 473.400 844.050 474.450 ;
        RECT 826.950 472.950 829.050 473.400 ;
        RECT 841.950 472.950 844.050 473.400 ;
        RECT 376.950 472.050 379.050 472.200 ;
        RECT 316.950 471.450 319.050 472.050 ;
        RECT 346.950 471.450 349.050 472.050 ;
        RECT 375.000 471.450 379.050 472.050 ;
        RECT 257.400 470.400 349.050 471.450 ;
        RECT 28.950 469.950 31.050 470.400 ;
        RECT 208.950 469.950 211.050 470.400 ;
        RECT 316.950 469.950 319.050 470.400 ;
        RECT 346.950 469.950 349.050 470.400 ;
        RECT 374.400 470.100 379.050 471.450 ;
        RECT 385.950 471.450 388.050 472.050 ;
        RECT 433.950 471.450 436.050 472.050 ;
        RECT 385.950 470.400 436.050 471.450 ;
        RECT 374.400 469.950 378.000 470.100 ;
        RECT 385.950 469.950 388.050 470.400 ;
        RECT 433.950 469.950 436.050 470.400 ;
        RECT 442.950 471.450 445.050 472.050 ;
        RECT 472.950 471.450 475.050 472.050 ;
        RECT 442.950 470.400 475.050 471.450 ;
        RECT 442.950 469.950 445.050 470.400 ;
        RECT 472.950 469.950 475.050 470.400 ;
        RECT 526.950 471.450 529.050 472.050 ;
        RECT 574.950 471.450 577.050 472.050 ;
        RECT 526.950 470.400 577.050 471.450 ;
        RECT 526.950 469.950 529.050 470.400 ;
        RECT 574.950 469.950 577.050 470.400 ;
        RECT 661.950 471.450 664.050 472.050 ;
        RECT 709.950 471.450 712.050 472.050 ;
        RECT 748.950 471.450 751.050 472.050 ;
        RECT 661.950 470.400 693.450 471.450 ;
        RECT 661.950 469.950 664.050 470.400 ;
        RECT 103.950 468.450 106.050 469.050 ;
        RECT 115.950 468.450 118.050 469.050 ;
        RECT 103.950 467.400 118.050 468.450 ;
        RECT 103.950 466.950 106.050 467.400 ;
        RECT 115.950 466.950 118.050 467.400 ;
        RECT 139.950 468.450 142.050 469.050 ;
        RECT 157.950 468.450 160.050 469.050 ;
        RECT 139.950 467.400 160.050 468.450 ;
        RECT 139.950 466.950 142.050 467.400 ;
        RECT 157.950 466.950 160.050 467.400 ;
        RECT 175.950 468.450 178.050 469.050 ;
        RECT 193.950 468.450 196.050 469.050 ;
        RECT 175.950 467.400 196.050 468.450 ;
        RECT 175.950 466.950 178.050 467.400 ;
        RECT 193.950 466.950 196.050 467.400 ;
        RECT 262.950 468.450 265.050 469.050 ;
        RECT 313.950 468.450 316.050 469.050 ;
        RECT 262.950 467.400 316.050 468.450 ;
        RECT 262.950 466.950 265.050 467.400 ;
        RECT 313.950 466.950 316.050 467.400 ;
        RECT 325.950 468.450 328.050 469.050 ;
        RECT 361.950 468.450 364.050 469.050 ;
        RECT 367.950 468.450 370.050 469.050 ;
        RECT 325.950 467.400 360.450 468.450 ;
        RECT 325.950 466.950 328.050 467.400 ;
        RECT 359.400 466.050 360.450 467.400 ;
        RECT 361.950 467.400 370.050 468.450 ;
        RECT 361.950 466.950 364.050 467.400 ;
        RECT 367.950 466.950 370.050 467.400 ;
        RECT 22.950 465.450 25.050 466.050 ;
        RECT 40.950 465.450 43.050 466.050 ;
        RECT 259.950 465.450 262.050 466.050 ;
        RECT 22.950 464.400 262.050 465.450 ;
        RECT 22.950 463.950 25.050 464.400 ;
        RECT 40.950 463.950 43.050 464.400 ;
        RECT 259.950 463.950 262.050 464.400 ;
        RECT 277.950 465.450 280.050 466.050 ;
        RECT 298.800 465.450 300.900 466.050 ;
        RECT 277.950 464.400 300.900 465.450 ;
        RECT 302.100 465.000 304.200 466.050 ;
        RECT 277.950 463.950 280.050 464.400 ;
        RECT 298.800 463.950 300.900 464.400 ;
        RECT 301.950 463.950 304.200 465.000 ;
        RECT 307.950 465.450 310.050 466.050 ;
        RECT 340.950 465.450 343.050 466.050 ;
        RECT 307.950 464.400 343.050 465.450 ;
        RECT 359.400 464.400 363.900 466.050 ;
        RECT 307.950 463.950 310.050 464.400 ;
        RECT 340.950 463.950 343.050 464.400 ;
        RECT 360.000 463.950 363.900 464.400 ;
        RECT 365.100 465.450 367.200 466.050 ;
        RECT 370.950 465.450 373.050 466.050 ;
        RECT 365.100 464.400 373.050 465.450 ;
        RECT 374.400 465.450 375.450 469.950 ;
        RECT 376.950 468.450 379.050 468.900 ;
        RECT 484.950 468.450 487.050 469.050 ;
        RECT 376.950 467.400 487.050 468.450 ;
        RECT 376.950 466.800 379.050 467.400 ;
        RECT 484.950 466.950 487.050 467.400 ;
        RECT 505.950 468.450 508.050 469.050 ;
        RECT 550.800 468.450 552.900 469.050 ;
        RECT 505.950 467.400 552.900 468.450 ;
        RECT 505.950 466.950 508.050 467.400 ;
        RECT 550.800 466.950 552.900 467.400 ;
        RECT 554.100 468.450 556.200 469.050 ;
        RECT 610.950 468.450 613.050 469.050 ;
        RECT 554.100 467.400 613.050 468.450 ;
        RECT 692.400 468.450 693.450 470.400 ;
        RECT 709.950 470.400 751.050 471.450 ;
        RECT 709.950 469.950 712.050 470.400 ;
        RECT 748.950 469.950 751.050 470.400 ;
        RECT 757.950 471.450 760.050 472.050 ;
        RECT 772.950 471.450 775.050 472.050 ;
        RECT 757.950 470.400 775.050 471.450 ;
        RECT 757.950 469.950 760.050 470.400 ;
        RECT 772.950 469.950 775.050 470.400 ;
        RECT 820.950 471.450 823.050 472.050 ;
        RECT 832.950 471.450 835.050 472.050 ;
        RECT 820.950 470.400 835.050 471.450 ;
        RECT 820.950 469.950 823.050 470.400 ;
        RECT 832.950 469.950 835.050 470.400 ;
        RECT 817.950 468.450 820.050 469.050 ;
        RECT 841.950 468.450 844.050 469.050 ;
        RECT 692.400 467.400 732.450 468.450 ;
        RECT 554.100 466.950 556.200 467.400 ;
        RECT 610.950 466.950 613.050 467.400 ;
        RECT 731.400 466.050 732.450 467.400 ;
        RECT 817.950 467.400 844.050 468.450 ;
        RECT 817.950 466.950 820.050 467.400 ;
        RECT 841.950 466.950 844.050 467.400 ;
        RECT 397.950 465.450 400.050 466.050 ;
        RECT 409.950 465.450 412.050 466.050 ;
        RECT 374.400 464.400 396.450 465.450 ;
        RECT 365.100 463.950 367.200 464.400 ;
        RECT 370.950 463.950 373.050 464.400 ;
        RECT 301.950 463.050 304.050 463.950 ;
        RECT 43.950 457.950 46.050 463.050 ;
        RECT 52.950 462.450 55.050 463.050 ;
        RECT 91.950 462.450 94.050 463.050 ;
        RECT 52.950 461.400 94.050 462.450 ;
        RECT 52.950 460.950 55.050 461.400 ;
        RECT 91.950 460.950 94.050 461.400 ;
        RECT 196.950 462.450 199.050 463.050 ;
        RECT 217.950 462.450 220.050 463.050 ;
        RECT 196.950 461.400 220.050 462.450 ;
        RECT 301.950 462.000 304.200 463.050 ;
        RECT 196.950 460.950 199.050 461.400 ;
        RECT 217.950 460.950 220.050 461.400 ;
        RECT 302.100 460.950 304.200 462.000 ;
        RECT 316.950 462.450 319.050 463.050 ;
        RECT 334.950 462.450 337.050 463.050 ;
        RECT 316.950 461.400 337.050 462.450 ;
        RECT 316.950 460.950 319.050 461.400 ;
        RECT 334.950 460.950 337.050 461.400 ;
        RECT 352.950 462.450 355.050 463.050 ;
        RECT 364.950 462.450 367.050 463.050 ;
        RECT 388.950 462.450 391.050 463.050 ;
        RECT 352.950 461.400 391.050 462.450 ;
        RECT 395.400 462.450 396.450 464.400 ;
        RECT 397.950 464.400 412.050 465.450 ;
        RECT 397.950 463.950 400.050 464.400 ;
        RECT 409.950 463.950 412.050 464.400 ;
        RECT 436.950 465.450 439.050 466.050 ;
        RECT 520.950 465.450 523.050 466.050 ;
        RECT 547.950 465.450 550.050 466.050 ;
        RECT 436.950 464.400 550.050 465.450 ;
        RECT 436.950 463.950 439.050 464.400 ;
        RECT 520.950 463.950 523.050 464.400 ;
        RECT 547.950 463.950 550.050 464.400 ;
        RECT 574.950 465.450 577.050 466.050 ;
        RECT 664.950 465.450 667.050 466.050 ;
        RECT 574.950 464.400 667.050 465.450 ;
        RECT 574.950 463.950 577.050 464.400 ;
        RECT 664.950 463.950 667.050 464.400 ;
        RECT 730.950 465.450 733.050 466.050 ;
        RECT 766.950 465.450 769.050 466.050 ;
        RECT 787.950 465.450 790.050 466.050 ;
        RECT 730.950 464.400 790.050 465.450 ;
        RECT 730.950 463.950 733.050 464.400 ;
        RECT 766.950 463.950 769.050 464.400 ;
        RECT 787.950 463.950 790.050 464.400 ;
        RECT 415.950 462.450 418.050 463.050 ;
        RECT 421.950 462.450 424.050 463.050 ;
        RECT 395.400 461.400 408.450 462.450 ;
        RECT 352.950 460.950 355.050 461.400 ;
        RECT 364.950 460.950 367.050 461.400 ;
        RECT 388.950 460.950 391.050 461.400 ;
        RECT 58.950 459.450 61.050 460.050 ;
        RECT 79.950 459.450 82.050 460.050 ;
        RECT 100.950 459.450 103.050 460.050 ;
        RECT 58.950 458.400 103.050 459.450 ;
        RECT 58.950 457.950 61.050 458.400 ;
        RECT 79.950 457.950 82.050 458.400 ;
        RECT 100.950 457.950 103.050 458.400 ;
        RECT 109.950 459.450 112.050 460.050 ;
        RECT 109.950 458.400 135.450 459.450 ;
        RECT 109.950 457.950 112.050 458.400 ;
        RECT 134.400 457.050 135.450 458.400 ;
        RECT 148.950 457.950 153.900 460.050 ;
        RECT 155.100 459.450 157.200 460.050 ;
        RECT 155.100 459.000 228.450 459.450 ;
        RECT 317.100 459.000 319.200 460.050 ;
        RECT 155.100 458.400 229.050 459.000 ;
        RECT 155.100 457.950 157.200 458.400 ;
        RECT 19.950 454.950 25.050 457.050 ;
        RECT 13.950 453.450 16.050 454.050 ;
        RECT 13.950 452.400 27.450 453.450 ;
        RECT 13.950 451.950 16.050 452.400 ;
        RECT 26.400 451.050 27.450 452.400 ;
        RECT 31.950 451.950 37.050 454.050 ;
        RECT 49.950 451.950 55.050 454.050 ;
        RECT 58.950 451.950 61.050 457.050 ;
        RECT 64.950 454.950 70.050 457.050 ;
        RECT 73.950 454.950 78.900 457.050 ;
        RECT 80.100 456.000 82.200 457.050 ;
        RECT 79.950 454.950 82.200 456.000 ;
        RECT 115.950 456.450 118.050 457.050 ;
        RECT 130.800 456.450 132.900 457.050 ;
        RECT 115.950 455.400 132.900 456.450 ;
        RECT 115.950 454.950 118.050 455.400 ;
        RECT 130.800 454.950 132.900 455.400 ;
        RECT 134.100 454.950 139.050 457.050 ;
        RECT 145.950 454.950 151.050 457.050 ;
        RECT 154.950 456.450 157.050 457.050 ;
        RECT 166.950 456.450 169.050 457.050 ;
        RECT 205.950 456.450 208.050 457.050 ;
        RECT 154.950 455.400 169.050 456.450 ;
        RECT 188.400 456.000 208.050 456.450 ;
        RECT 154.950 454.950 157.050 455.400 ;
        RECT 166.950 454.950 169.050 455.400 ;
        RECT 187.950 455.400 208.050 456.000 ;
        RECT 70.950 451.950 76.050 454.050 ;
        RECT 79.950 451.950 82.050 454.950 ;
        RECT 91.950 451.950 97.050 454.050 ;
        RECT 100.950 453.450 103.050 454.050 ;
        RECT 109.950 453.450 112.050 454.050 ;
        RECT 100.950 452.400 112.050 453.450 ;
        RECT 100.950 451.950 103.050 452.400 ;
        RECT 109.950 451.950 112.050 452.400 ;
        RECT 124.950 451.950 129.900 454.050 ;
        RECT 131.100 451.950 136.050 454.050 ;
        RECT 136.950 453.450 139.050 454.950 ;
        RECT 154.950 453.450 157.050 454.050 ;
        RECT 166.950 453.450 169.050 454.050 ;
        RECT 136.950 453.000 157.050 453.450 ;
        RECT 137.400 452.400 157.050 453.000 ;
        RECT 154.950 451.950 157.050 452.400 ;
        RECT 158.400 452.400 169.050 453.450 ;
        RECT 25.950 448.950 31.050 451.050 ;
        RECT 34.950 450.450 37.050 451.050 ;
        RECT 40.800 450.450 42.900 451.050 ;
        RECT 34.950 449.400 42.900 450.450 ;
        RECT 34.950 448.950 37.050 449.400 ;
        RECT 40.800 448.950 42.900 449.400 ;
        RECT 44.100 448.950 49.050 451.050 ;
        RECT 55.950 447.450 58.050 451.050 ;
        RECT 73.950 447.450 76.050 448.050 ;
        RECT 55.950 447.000 76.050 447.450 ;
        RECT 56.400 446.400 76.050 447.000 ;
        RECT 73.950 445.950 76.050 446.400 ;
        RECT 97.950 447.450 100.050 451.050 ;
        RECT 145.950 450.450 148.050 451.050 ;
        RECT 158.400 450.450 159.450 452.400 ;
        RECT 166.950 451.950 169.050 452.400 ;
        RECT 181.950 453.450 184.050 454.050 ;
        RECT 187.950 453.450 190.050 455.400 ;
        RECT 205.950 454.950 208.050 455.400 ;
        RECT 214.950 456.450 217.050 457.050 ;
        RECT 220.950 456.450 223.050 457.050 ;
        RECT 214.950 455.400 223.050 456.450 ;
        RECT 214.950 454.950 217.050 455.400 ;
        RECT 220.950 454.950 223.050 455.400 ;
        RECT 226.950 454.950 229.050 458.400 ;
        RECT 316.950 457.950 319.200 459.000 ;
        RECT 361.950 459.450 364.050 460.050 ;
        RECT 382.950 459.450 385.050 460.050 ;
        RECT 403.950 459.450 406.050 460.050 ;
        RECT 361.950 458.400 385.050 459.450 ;
        RECT 392.400 459.000 406.050 459.450 ;
        RECT 361.950 457.950 364.050 458.400 ;
        RECT 382.950 457.950 385.050 458.400 ;
        RECT 391.950 458.400 406.050 459.000 ;
        RECT 313.800 457.050 315.900 457.200 ;
        RECT 232.950 454.950 238.050 457.050 ;
        RECT 253.950 456.450 256.050 457.050 ;
        RECT 265.950 456.450 268.050 457.050 ;
        RECT 253.950 455.400 268.050 456.450 ;
        RECT 253.950 454.950 256.050 455.400 ;
        RECT 265.950 454.950 268.050 455.400 ;
        RECT 181.950 452.400 190.050 453.450 ;
        RECT 181.950 451.950 184.050 452.400 ;
        RECT 187.950 451.950 190.050 452.400 ;
        RECT 145.950 449.400 159.450 450.450 ;
        RECT 145.950 448.950 148.050 449.400 ;
        RECT 160.950 448.950 166.050 451.050 ;
        RECT 169.950 450.450 172.050 451.050 ;
        RECT 187.950 450.450 193.050 451.050 ;
        RECT 169.950 449.400 193.050 450.450 ;
        RECT 193.950 450.450 196.050 454.050 ;
        RECT 202.950 451.950 208.050 454.050 ;
        RECT 220.950 451.950 225.900 454.050 ;
        RECT 227.100 451.950 232.050 454.050 ;
        RECT 262.950 453.450 265.050 454.050 ;
        RECT 268.950 453.450 271.050 454.050 ;
        RECT 262.950 452.400 271.050 453.450 ;
        RECT 262.950 451.950 265.050 452.400 ;
        RECT 268.950 451.950 271.050 452.400 ;
        RECT 274.950 451.950 277.050 457.050 ;
        RECT 280.950 454.950 286.050 457.050 ;
        RECT 289.950 456.450 292.050 457.050 ;
        RECT 298.950 456.450 301.050 457.050 ;
        RECT 289.950 455.400 301.050 456.450 ;
        RECT 289.950 454.950 292.050 455.400 ;
        RECT 298.950 454.950 301.050 455.400 ;
        RECT 307.800 456.000 309.900 457.050 ;
        RECT 307.800 454.950 310.050 456.000 ;
        RECT 311.100 455.100 315.900 457.050 ;
        RECT 316.950 457.050 319.050 457.950 ;
        RECT 391.950 457.050 394.050 458.400 ;
        RECT 403.950 457.950 406.050 458.400 ;
        RECT 407.400 457.050 408.450 461.400 ;
        RECT 415.950 461.400 424.050 462.450 ;
        RECT 415.950 460.950 418.050 461.400 ;
        RECT 421.950 460.950 424.050 461.400 ;
        RECT 445.950 462.450 448.050 463.050 ;
        RECT 505.950 462.450 508.050 463.050 ;
        RECT 445.950 461.400 508.050 462.450 ;
        RECT 445.950 460.950 448.050 461.400 ;
        RECT 505.950 460.950 508.050 461.400 ;
        RECT 634.800 462.000 636.900 463.050 ;
        RECT 676.950 462.450 679.050 463.050 ;
        RECT 688.800 462.450 690.900 463.050 ;
        RECT 634.800 460.950 637.050 462.000 ;
        RECT 676.950 461.400 690.900 462.450 ;
        RECT 676.950 460.950 679.050 461.400 ;
        RECT 688.800 460.950 690.900 461.400 ;
        RECT 692.100 462.450 694.200 463.050 ;
        RECT 706.950 462.450 709.050 463.050 ;
        RECT 692.100 461.400 709.050 462.450 ;
        RECT 692.100 460.950 694.200 461.400 ;
        RECT 706.950 460.950 709.050 461.400 ;
        RECT 634.950 460.050 637.050 460.950 ;
        RECT 316.950 456.000 319.200 457.050 ;
        RECT 311.100 454.950 315.000 455.100 ;
        RECT 317.100 454.950 319.200 456.000 ;
        RECT 325.950 454.950 331.050 457.050 ;
        RECT 343.950 454.950 349.050 457.050 ;
        RECT 352.800 456.000 354.900 457.050 ;
        RECT 352.800 454.950 355.050 456.000 ;
        RECT 356.100 454.950 361.050 457.050 ;
        RECT 391.800 456.000 394.050 457.050 ;
        RECT 391.800 454.950 393.900 456.000 ;
        RECT 395.100 454.950 400.050 457.050 ;
        RECT 406.950 454.950 409.050 457.050 ;
        RECT 412.950 454.950 415.050 460.050 ;
        RECT 424.950 454.950 430.050 457.050 ;
        RECT 433.950 454.950 436.050 460.050 ;
        RECT 454.950 459.450 457.050 460.050 ;
        RECT 463.800 459.450 465.900 460.050 ;
        RECT 454.950 458.400 465.900 459.450 ;
        RECT 454.950 457.950 457.050 458.400 ;
        RECT 463.800 457.950 465.900 458.400 ;
        RECT 467.100 459.450 469.200 460.050 ;
        RECT 493.950 459.450 496.050 460.050 ;
        RECT 580.950 459.450 583.050 460.050 ;
        RECT 586.950 459.450 589.050 460.050 ;
        RECT 601.950 459.450 604.050 460.050 ;
        RECT 467.100 459.000 492.450 459.450 ;
        RECT 493.950 459.000 513.450 459.450 ;
        RECT 467.100 458.400 493.050 459.000 ;
        RECT 467.100 457.950 469.200 458.400 ;
        RECT 490.950 457.050 493.050 458.400 ;
        RECT 493.950 458.400 514.050 459.000 ;
        RECT 493.950 457.950 496.050 458.400 ;
        RECT 307.950 454.050 310.050 454.950 ;
        RECT 283.950 451.950 289.050 454.050 ;
        RECT 292.950 451.950 298.050 454.050 ;
        RECT 307.800 453.000 310.050 454.050 ;
        RECT 307.800 451.950 309.900 453.000 ;
        RECT 311.100 451.950 316.050 454.050 ;
        RECT 319.950 453.450 322.050 454.050 ;
        RECT 331.950 453.450 334.050 454.050 ;
        RECT 319.950 452.400 334.050 453.450 ;
        RECT 319.950 451.950 322.050 452.400 ;
        RECT 331.950 451.950 334.050 452.400 ;
        RECT 352.950 451.950 355.050 454.950 ;
        RECT 370.950 451.950 376.050 454.050 ;
        RECT 379.950 453.450 382.050 454.050 ;
        RECT 385.950 453.450 391.050 454.050 ;
        RECT 379.950 452.400 391.050 453.450 ;
        RECT 379.950 451.950 382.050 452.400 ;
        RECT 385.950 451.950 391.050 452.400 ;
        RECT 394.950 451.950 400.050 454.050 ;
        RECT 403.950 453.450 406.050 454.050 ;
        RECT 409.950 453.450 412.050 454.050 ;
        RECT 403.950 452.400 412.050 453.450 ;
        RECT 403.950 451.950 406.050 452.400 ;
        RECT 409.950 451.950 412.050 452.400 ;
        RECT 421.950 453.450 424.050 454.050 ;
        RECT 430.950 453.450 433.050 454.050 ;
        RECT 421.950 452.400 433.050 453.450 ;
        RECT 421.950 451.950 424.050 452.400 ;
        RECT 430.950 451.950 433.050 452.400 ;
        RECT 454.950 453.450 457.050 454.050 ;
        RECT 463.950 453.450 466.050 457.050 ;
        RECT 469.950 456.450 472.050 457.050 ;
        RECT 469.950 455.400 483.450 456.450 ;
        RECT 469.950 454.950 472.050 455.400 ;
        RECT 454.950 453.000 466.050 453.450 ;
        RECT 454.950 452.400 465.450 453.000 ;
        RECT 454.950 451.950 457.050 452.400 ;
        RECT 466.950 451.950 471.900 454.050 ;
        RECT 482.400 453.450 483.450 455.400 ;
        RECT 484.950 454.950 489.900 457.050 ;
        RECT 490.800 456.000 493.050 457.050 ;
        RECT 494.100 456.000 496.200 457.050 ;
        RECT 490.800 454.950 492.900 456.000 ;
        RECT 493.950 454.950 496.200 456.000 ;
        RECT 499.950 456.450 502.050 457.050 ;
        RECT 505.950 456.450 508.050 457.050 ;
        RECT 499.950 455.400 508.050 456.450 ;
        RECT 499.950 454.950 502.050 455.400 ;
        RECT 505.950 454.950 508.050 455.400 ;
        RECT 511.950 454.950 514.050 458.400 ;
        RECT 580.950 458.400 589.050 459.450 ;
        RECT 580.950 457.950 583.050 458.400 ;
        RECT 586.950 457.950 589.050 458.400 ;
        RECT 590.400 458.400 604.050 459.450 ;
        RECT 529.950 454.950 534.900 457.050 ;
        RECT 536.100 454.950 541.050 457.050 ;
        RECT 562.950 454.950 568.050 457.050 ;
        RECT 583.950 456.450 586.050 457.050 ;
        RECT 590.400 456.450 591.450 458.400 ;
        RECT 601.950 457.950 604.050 458.400 ;
        RECT 583.950 455.400 591.450 456.450 ;
        RECT 583.950 454.950 586.050 455.400 ;
        RECT 487.950 453.450 490.050 454.050 ;
        RECT 482.400 452.400 490.050 453.450 ;
        RECT 487.950 451.950 490.050 452.400 ;
        RECT 493.950 451.950 496.050 454.950 ;
        RECT 505.950 451.950 511.050 454.050 ;
        RECT 514.950 451.950 520.050 454.050 ;
        RECT 202.950 450.450 205.050 451.050 ;
        RECT 193.950 450.000 205.050 450.450 ;
        RECT 194.400 449.400 205.050 450.000 ;
        RECT 169.950 448.950 172.050 449.400 ;
        RECT 187.950 448.950 193.050 449.400 ;
        RECT 130.950 447.450 133.050 448.050 ;
        RECT 97.950 446.400 133.050 447.450 ;
        RECT 97.950 445.950 100.050 446.400 ;
        RECT 130.950 445.950 133.050 446.400 ;
        RECT 202.950 445.950 205.050 449.400 ;
        RECT 208.950 450.450 211.050 451.050 ;
        RECT 217.950 450.450 220.050 451.050 ;
        RECT 227.400 450.450 228.450 451.950 ;
        RECT 208.950 449.400 228.450 450.450 ;
        RECT 271.950 450.450 274.050 451.050 ;
        RECT 298.950 450.450 301.050 451.050 ;
        RECT 271.950 449.400 301.050 450.450 ;
        RECT 208.950 448.950 211.050 449.400 ;
        RECT 217.950 448.950 220.050 449.400 ;
        RECT 271.950 448.950 274.050 449.400 ;
        RECT 298.950 448.950 301.050 449.400 ;
        RECT 343.950 450.450 346.050 451.050 ;
        RECT 370.950 450.450 373.050 451.050 ;
        RECT 343.950 449.400 373.050 450.450 ;
        RECT 343.950 448.950 346.050 449.400 ;
        RECT 370.950 448.950 373.050 449.400 ;
        RECT 376.950 450.450 379.050 451.050 ;
        RECT 382.950 450.450 385.050 451.050 ;
        RECT 394.950 450.450 397.050 451.050 ;
        RECT 376.950 449.400 397.050 450.450 ;
        RECT 376.950 448.950 379.050 449.400 ;
        RECT 382.950 448.950 385.050 449.400 ;
        RECT 394.950 448.950 397.050 449.400 ;
        RECT 511.950 450.450 514.050 451.050 ;
        RECT 532.800 450.450 534.900 451.050 ;
        RECT 511.950 449.400 534.900 450.450 ;
        RECT 511.950 448.950 514.050 449.400 ;
        RECT 532.800 448.950 534.900 449.400 ;
        RECT 536.100 450.450 538.200 451.050 ;
        RECT 547.950 450.450 550.050 454.050 ;
        RECT 553.950 453.450 556.050 454.050 ;
        RECT 559.950 453.450 562.050 454.050 ;
        RECT 553.950 452.400 562.050 453.450 ;
        RECT 553.950 451.950 556.050 452.400 ;
        RECT 559.950 451.950 562.050 452.400 ;
        RECT 586.950 453.450 589.050 454.050 ;
        RECT 598.950 453.450 601.050 457.050 ;
        RECT 613.950 454.950 616.050 460.050 ;
        RECT 634.800 459.000 637.050 460.050 ;
        RECT 634.800 457.950 636.900 459.000 ;
        RECT 586.950 453.000 601.050 453.450 ;
        RECT 619.950 453.450 622.050 454.050 ;
        RECT 631.950 453.450 634.050 457.050 ;
        RECT 646.950 454.050 649.050 457.050 ;
        RECT 652.950 454.950 655.050 460.050 ;
        RECT 715.950 459.450 718.050 460.050 ;
        RECT 778.950 459.450 781.050 460.050 ;
        RECT 793.800 459.450 795.900 460.050 ;
        RECT 692.400 459.000 711.450 459.450 ;
        RECT 691.950 458.400 712.050 459.000 ;
        RECT 664.950 456.450 667.050 457.050 ;
        RECT 685.950 456.450 688.050 457.200 ;
        RECT 664.950 455.400 688.050 456.450 ;
        RECT 664.950 454.950 667.050 455.400 ;
        RECT 685.950 454.950 688.050 455.400 ;
        RECT 691.950 454.950 694.050 458.400 ;
        RECT 619.950 453.000 634.050 453.450 ;
        RECT 646.800 453.000 649.050 454.050 ;
        RECT 650.100 453.000 652.200 454.050 ;
        RECT 586.950 452.400 600.450 453.000 ;
        RECT 619.950 452.400 633.450 453.000 ;
        RECT 586.950 451.950 589.050 452.400 ;
        RECT 619.950 451.950 622.050 452.400 ;
        RECT 646.800 451.950 648.900 453.000 ;
        RECT 649.950 451.950 652.200 453.000 ;
        RECT 655.950 453.450 658.050 454.050 ;
        RECT 661.950 453.450 664.050 454.050 ;
        RECT 655.950 452.400 664.050 453.450 ;
        RECT 655.950 451.950 658.050 452.400 ;
        RECT 661.950 451.950 664.050 452.400 ;
        RECT 673.950 453.450 676.050 454.050 ;
        RECT 687.000 453.900 691.050 454.050 ;
        RECT 673.950 452.400 684.450 453.450 ;
        RECT 673.950 451.950 676.050 452.400 ;
        RECT 536.100 449.400 550.050 450.450 ;
        RECT 536.100 448.950 538.200 449.400 ;
        RECT 547.950 448.950 550.050 449.400 ;
        RECT 556.950 450.450 559.050 451.050 ;
        RECT 601.950 450.450 604.050 451.050 ;
        RECT 556.950 449.400 604.050 450.450 ;
        RECT 556.950 448.950 559.050 449.400 ;
        RECT 601.950 448.950 604.050 449.400 ;
        RECT 607.950 450.450 610.050 451.050 ;
        RECT 613.950 450.450 616.050 451.050 ;
        RECT 625.950 450.450 628.050 451.050 ;
        RECT 607.950 449.400 628.050 450.450 ;
        RECT 607.950 448.950 610.050 449.400 ;
        RECT 613.950 448.950 616.050 449.400 ;
        RECT 625.950 448.950 628.050 449.400 ;
        RECT 634.950 450.450 637.050 451.050 ;
        RECT 649.950 450.450 652.050 451.950 ;
        RECT 634.950 450.000 652.050 450.450 ;
        RECT 634.950 449.400 651.600 450.000 ;
        RECT 634.950 448.950 637.050 449.400 ;
        RECT 670.950 448.950 675.900 451.050 ;
        RECT 677.100 450.000 679.200 451.050 ;
        RECT 676.950 448.950 679.200 450.000 ;
        RECT 683.400 450.450 684.450 452.400 ;
        RECT 685.950 451.950 691.050 453.900 ;
        RECT 685.950 451.800 688.050 451.950 ;
        RECT 694.950 450.450 697.050 454.050 ;
        RECT 697.950 453.450 700.050 457.050 ;
        RECT 709.950 454.950 712.050 458.400 ;
        RECT 715.950 458.400 795.900 459.450 ;
        RECT 797.100 459.000 799.200 460.050 ;
        RECT 715.950 454.950 718.050 458.400 ;
        RECT 778.950 457.950 781.050 458.400 ;
        RECT 793.800 457.950 795.900 458.400 ;
        RECT 796.950 457.950 799.200 459.000 ;
        RECT 802.950 459.450 805.050 460.050 ;
        RECT 820.950 459.450 823.050 460.050 ;
        RECT 802.950 458.400 823.050 459.450 ;
        RECT 802.950 457.950 805.050 458.400 ;
        RECT 820.950 457.950 823.050 458.400 ;
        RECT 829.950 457.950 835.050 460.050 ;
        RECT 796.950 457.050 799.050 457.950 ;
        RECT 784.950 456.450 787.050 457.050 ;
        RECT 755.400 456.000 787.050 456.450 ;
        RECT 754.950 455.400 787.050 456.000 ;
        RECT 703.950 453.450 706.050 454.050 ;
        RECT 697.950 453.000 706.050 453.450 ;
        RECT 698.400 452.400 706.050 453.000 ;
        RECT 703.950 451.950 706.050 452.400 ;
        RECT 712.800 453.000 714.900 454.050 ;
        RECT 717.000 453.900 721.050 454.050 ;
        RECT 712.800 451.950 715.050 453.000 ;
        RECT 712.950 451.050 715.050 451.950 ;
        RECT 716.100 451.950 721.050 453.900 ;
        RECT 730.800 453.000 732.900 454.050 ;
        RECT 734.100 453.450 736.200 454.050 ;
        RECT 742.800 453.450 744.900 454.050 ;
        RECT 730.800 451.950 733.050 453.000 ;
        RECT 734.100 452.400 744.900 453.450 ;
        RECT 734.100 451.950 736.200 452.400 ;
        RECT 742.800 451.950 744.900 452.400 ;
        RECT 746.100 451.950 751.050 454.050 ;
        RECT 754.950 451.950 757.050 455.400 ;
        RECT 784.950 454.950 787.050 455.400 ;
        RECT 796.800 456.000 799.050 457.050 ;
        RECT 800.100 456.000 802.200 457.050 ;
        RECT 803.100 456.000 805.200 457.050 ;
        RECT 796.800 454.950 798.900 456.000 ;
        RECT 799.950 454.950 802.200 456.000 ;
        RECT 802.950 454.950 805.200 456.000 ;
        RECT 808.950 456.450 811.050 457.050 ;
        RECT 817.950 456.450 820.050 457.050 ;
        RECT 808.950 455.400 820.050 456.450 ;
        RECT 808.950 454.950 811.050 455.400 ;
        RECT 817.950 454.950 820.050 455.400 ;
        RECT 823.950 456.450 826.050 457.050 ;
        RECT 835.950 456.450 841.050 457.050 ;
        RECT 823.950 455.400 841.050 456.450 ;
        RECT 823.950 454.950 826.050 455.400 ;
        RECT 835.950 454.950 841.050 455.400 ;
        RECT 799.950 454.050 802.050 454.950 ;
        RECT 766.950 451.950 772.050 454.050 ;
        RECT 775.950 451.950 781.050 454.050 ;
        RECT 790.950 451.950 796.050 454.050 ;
        RECT 799.800 453.000 802.050 454.050 ;
        RECT 802.950 454.050 805.050 454.950 ;
        RECT 802.950 453.000 805.200 454.050 ;
        RECT 799.800 451.950 801.900 453.000 ;
        RECT 803.100 451.950 805.200 453.000 ;
        RECT 716.100 451.800 718.200 451.950 ;
        RECT 730.950 451.050 733.050 451.950 ;
        RECT 683.400 450.000 697.050 450.450 ;
        RECT 712.800 450.000 715.050 451.050 ;
        RECT 683.400 449.400 696.450 450.000 ;
        RECT 712.800 448.950 714.900 450.000 ;
        RECT 724.950 448.950 729.900 451.050 ;
        RECT 730.950 450.000 733.200 451.050 ;
        RECT 731.100 448.950 733.200 450.000 ;
        RECT 736.950 448.950 742.050 451.050 ;
        RECT 232.950 447.450 235.050 448.050 ;
        RECT 280.950 447.450 283.050 448.050 ;
        RECT 232.950 446.400 283.050 447.450 ;
        RECT 232.950 445.950 235.050 446.400 ;
        RECT 280.950 445.950 283.050 446.400 ;
        RECT 358.950 447.450 361.050 448.050 ;
        RECT 373.950 447.450 376.050 448.050 ;
        RECT 358.950 446.400 376.050 447.450 ;
        RECT 358.950 445.950 361.050 446.400 ;
        RECT 373.950 445.950 376.050 446.400 ;
        RECT 424.950 447.450 427.050 448.050 ;
        RECT 466.950 447.450 469.050 448.050 ;
        RECT 424.950 446.400 469.050 447.450 ;
        RECT 424.950 445.950 427.050 446.400 ;
        RECT 466.950 445.950 469.050 446.400 ;
        RECT 484.950 447.450 487.050 448.050 ;
        RECT 538.800 447.450 540.900 448.050 ;
        RECT 484.950 446.400 540.900 447.450 ;
        RECT 484.950 445.950 487.050 446.400 ;
        RECT 538.800 445.950 540.900 446.400 ;
        RECT 542.100 447.450 544.200 448.050 ;
        RECT 559.950 447.450 562.050 448.050 ;
        RECT 595.950 447.450 598.050 448.050 ;
        RECT 542.100 446.400 598.050 447.450 ;
        RECT 542.100 445.950 544.200 446.400 ;
        RECT 559.950 445.950 562.050 446.400 ;
        RECT 595.950 445.950 598.050 446.400 ;
        RECT 641.100 447.450 643.200 448.050 ;
        RECT 655.950 447.450 658.050 448.050 ;
        RECT 641.100 446.400 658.050 447.450 ;
        RECT 641.100 445.950 643.200 446.400 ;
        RECT 655.950 445.950 658.050 446.400 ;
        RECT 664.950 447.450 667.050 448.050 ;
        RECT 676.950 447.450 679.050 448.950 ;
        RECT 664.950 447.000 679.050 447.450 ;
        RECT 715.950 447.450 718.050 448.050 ;
        RECT 745.950 447.450 748.050 448.050 ;
        RECT 664.950 446.400 678.600 447.000 ;
        RECT 715.950 446.400 748.050 447.450 ;
        RECT 751.950 447.450 754.050 451.050 ;
        RECT 760.950 448.950 766.050 451.050 ;
        RECT 769.950 448.950 775.050 451.050 ;
        RECT 796.950 450.450 799.050 451.050 ;
        RECT 814.950 450.450 817.050 454.050 ;
        RECT 796.950 450.000 817.050 450.450 ;
        RECT 796.950 449.400 816.450 450.000 ;
        RECT 796.950 448.950 799.050 449.400 ;
        RECT 820.950 448.950 823.050 454.050 ;
        RECT 826.950 453.450 829.050 454.050 ;
        RECT 841.950 453.450 844.050 454.050 ;
        RECT 826.950 452.400 844.050 453.450 ;
        RECT 826.950 451.950 829.050 452.400 ;
        RECT 841.950 451.950 844.050 452.400 ;
        RECT 763.800 447.450 765.900 448.050 ;
        RECT 751.950 447.000 765.900 447.450 ;
        RECT 752.400 446.400 765.900 447.000 ;
        RECT 664.950 445.950 667.050 446.400 ;
        RECT 715.950 445.950 718.050 446.400 ;
        RECT 745.950 445.950 748.050 446.400 ;
        RECT 763.800 445.950 765.900 446.400 ;
        RECT 767.100 447.450 769.200 448.050 ;
        RECT 772.950 447.450 775.050 448.200 ;
        RECT 767.100 446.400 775.050 447.450 ;
        RECT 767.100 445.950 769.200 446.400 ;
        RECT 772.950 446.100 775.050 446.400 ;
        RECT 790.950 447.450 795.000 448.050 ;
        RECT 790.950 445.950 795.450 447.450 ;
        RECT 10.950 444.450 13.050 445.050 ;
        RECT 40.950 444.450 43.050 445.050 ;
        RECT 55.950 444.450 58.050 445.050 ;
        RECT 10.950 443.400 58.050 444.450 ;
        RECT 10.950 442.950 13.050 443.400 ;
        RECT 40.950 442.950 43.050 443.400 ;
        RECT 55.950 442.950 58.050 443.400 ;
        RECT 37.950 441.450 40.050 442.050 ;
        RECT 43.950 441.450 46.050 442.050 ;
        RECT 37.950 440.400 46.050 441.450 ;
        RECT 37.950 439.950 40.050 440.400 ;
        RECT 43.950 439.950 46.050 440.400 ;
        RECT 85.950 439.950 88.050 445.050 ;
        RECT 91.950 444.450 94.050 445.050 ;
        RECT 124.950 444.450 127.050 445.050 ;
        RECT 178.950 444.450 181.050 445.050 ;
        RECT 91.950 443.400 181.050 444.450 ;
        RECT 91.950 442.950 94.050 443.400 ;
        RECT 124.950 442.950 127.050 443.400 ;
        RECT 178.950 442.950 181.050 443.400 ;
        RECT 202.950 444.450 205.050 445.050 ;
        RECT 214.950 444.450 217.050 445.050 ;
        RECT 241.950 444.450 244.050 445.050 ;
        RECT 202.950 443.400 244.050 444.450 ;
        RECT 202.950 442.950 205.050 443.400 ;
        RECT 214.950 442.950 217.050 443.400 ;
        RECT 241.950 442.950 244.050 443.400 ;
        RECT 268.950 444.450 271.050 445.050 ;
        RECT 292.950 444.450 295.050 445.050 ;
        RECT 268.950 443.400 295.050 444.450 ;
        RECT 268.950 442.950 271.050 443.400 ;
        RECT 292.950 442.950 295.050 443.400 ;
        RECT 301.950 442.950 307.050 445.050 ;
        RECT 364.950 444.450 367.050 445.050 ;
        RECT 382.950 444.450 385.050 445.050 ;
        RECT 364.950 443.400 385.050 444.450 ;
        RECT 364.950 442.950 367.050 443.400 ;
        RECT 382.950 442.950 385.050 443.400 ;
        RECT 421.950 444.450 424.050 445.050 ;
        RECT 445.950 444.450 448.050 445.050 ;
        RECT 421.950 443.400 448.050 444.450 ;
        RECT 421.950 442.950 424.050 443.400 ;
        RECT 445.950 442.950 448.050 443.400 ;
        RECT 457.950 444.450 460.050 445.050 ;
        RECT 508.950 444.450 511.050 445.050 ;
        RECT 457.950 443.400 511.050 444.450 ;
        RECT 457.950 442.950 460.050 443.400 ;
        RECT 508.950 442.950 511.050 443.400 ;
        RECT 550.950 444.450 553.050 445.050 ;
        RECT 613.950 444.450 616.050 445.050 ;
        RECT 550.950 443.400 616.050 444.450 ;
        RECT 550.950 442.950 553.050 443.400 ;
        RECT 613.950 442.950 616.050 443.400 ;
        RECT 625.950 444.450 628.050 445.050 ;
        RECT 697.950 444.450 700.050 445.050 ;
        RECT 625.950 443.400 700.050 444.450 ;
        RECT 625.950 442.950 628.050 443.400 ;
        RECT 697.950 442.950 700.050 443.400 ;
        RECT 712.950 444.450 715.050 445.200 ;
        RECT 742.950 444.450 745.050 445.050 ;
        RECT 712.950 443.400 745.050 444.450 ;
        RECT 712.950 443.100 715.050 443.400 ;
        RECT 742.950 442.950 745.050 443.400 ;
        RECT 772.950 444.450 775.050 444.900 ;
        RECT 784.950 444.450 787.050 445.050 ;
        RECT 772.950 443.400 787.050 444.450 ;
        RECT 794.400 444.450 795.450 445.950 ;
        RECT 832.950 444.450 835.050 445.050 ;
        RECT 794.400 443.400 835.050 444.450 ;
        RECT 772.950 442.800 775.050 443.400 ;
        RECT 784.950 442.950 787.050 443.400 ;
        RECT 832.950 442.950 835.050 443.400 ;
        RECT 187.950 441.450 190.050 442.050 ;
        RECT 220.950 441.450 223.050 442.050 ;
        RECT 187.950 440.400 223.050 441.450 ;
        RECT 187.950 439.950 190.050 440.400 ;
        RECT 220.950 439.950 223.050 440.400 ;
        RECT 271.950 441.450 274.050 442.050 ;
        RECT 313.950 441.450 316.050 442.050 ;
        RECT 334.950 441.450 337.050 442.050 ;
        RECT 271.950 440.400 337.050 441.450 ;
        RECT 271.950 439.950 274.050 440.400 ;
        RECT 313.950 439.950 316.050 440.400 ;
        RECT 334.950 439.950 337.050 440.400 ;
        RECT 343.950 441.450 346.050 442.050 ;
        RECT 397.950 441.450 400.050 442.050 ;
        RECT 343.950 440.400 400.050 441.450 ;
        RECT 343.950 439.950 346.050 440.400 ;
        RECT 397.950 439.950 400.050 440.400 ;
        RECT 529.950 441.450 532.050 442.050 ;
        RECT 607.800 441.450 609.900 442.050 ;
        RECT 529.950 440.400 609.900 441.450 ;
        RECT 529.950 439.950 532.050 440.400 ;
        RECT 607.800 439.950 609.900 440.400 ;
        RECT 611.100 441.450 613.200 442.050 ;
        RECT 616.950 441.450 619.050 442.200 ;
        RECT 611.100 440.400 619.050 441.450 ;
        RECT 611.100 439.950 613.200 440.400 ;
        RECT 616.950 440.100 619.050 440.400 ;
        RECT 670.950 441.450 673.050 442.050 ;
        RECT 682.950 441.450 685.050 442.050 ;
        RECT 670.950 440.400 685.050 441.450 ;
        RECT 670.950 439.950 673.050 440.400 ;
        RECT 682.950 439.950 685.050 440.400 ;
        RECT 712.950 441.450 715.050 441.900 ;
        RECT 724.950 441.450 727.050 442.050 ;
        RECT 712.950 440.400 727.050 441.450 ;
        RECT 712.950 439.800 715.050 440.400 ;
        RECT 724.950 439.950 727.050 440.400 ;
        RECT 793.950 441.450 796.050 442.050 ;
        RECT 829.950 441.450 832.050 442.050 ;
        RECT 793.950 440.400 832.050 441.450 ;
        RECT 793.950 439.950 796.050 440.400 ;
        RECT 829.950 439.950 832.050 440.400 ;
        RECT 4.950 438.450 7.050 439.050 ;
        RECT 28.950 438.450 31.050 439.050 ;
        RECT 4.950 437.400 31.050 438.450 ;
        RECT 4.950 436.950 7.050 437.400 ;
        RECT 28.950 436.950 31.050 437.400 ;
        RECT 70.950 438.450 73.050 439.050 ;
        RECT 148.950 438.450 151.050 439.050 ;
        RECT 70.950 437.400 151.050 438.450 ;
        RECT 70.950 436.950 73.050 437.400 ;
        RECT 148.950 436.950 151.050 437.400 ;
        RECT 346.950 438.450 349.050 439.050 ;
        RECT 445.950 438.450 448.050 439.050 ;
        RECT 346.950 437.400 448.050 438.450 ;
        RECT 346.950 436.950 349.050 437.400 ;
        RECT 445.950 436.950 448.050 437.400 ;
        RECT 538.950 438.450 541.050 439.050 ;
        RECT 577.950 438.450 580.050 439.050 ;
        RECT 601.950 438.450 604.050 439.050 ;
        RECT 538.950 437.400 604.050 438.450 ;
        RECT 538.950 436.950 541.050 437.400 ;
        RECT 577.950 436.950 580.050 437.400 ;
        RECT 601.950 436.950 604.050 437.400 ;
        RECT 616.950 438.450 619.050 438.900 ;
        RECT 640.800 438.450 642.900 439.050 ;
        RECT 616.950 437.400 642.900 438.450 ;
        RECT 616.950 436.800 619.050 437.400 ;
        RECT 640.800 436.950 642.900 437.400 ;
        RECT 644.100 438.450 646.200 439.050 ;
        RECT 652.800 438.450 654.900 439.050 ;
        RECT 644.100 437.400 654.900 438.450 ;
        RECT 644.100 436.950 646.200 437.400 ;
        RECT 652.800 436.950 654.900 437.400 ;
        RECT 736.950 438.450 739.050 438.900 ;
        RECT 742.950 438.450 745.050 439.050 ;
        RECT 736.950 437.400 745.050 438.450 ;
        RECT 736.950 436.800 739.050 437.400 ;
        RECT 742.950 436.950 745.050 437.400 ;
        RECT 748.950 438.450 751.050 439.050 ;
        RECT 808.950 438.450 811.050 439.050 ;
        RECT 748.950 437.400 811.050 438.450 ;
        RECT 748.950 436.950 751.050 437.400 ;
        RECT 808.950 436.950 811.050 437.400 ;
        RECT 838.950 438.450 841.050 439.050 ;
        RECT 844.950 438.450 847.050 439.050 ;
        RECT 838.950 437.400 847.050 438.450 ;
        RECT 838.950 436.950 841.050 437.400 ;
        RECT 844.950 436.950 847.050 437.400 ;
        RECT 1.950 435.450 4.050 436.050 ;
        RECT 10.950 435.450 13.050 436.050 ;
        RECT 1.950 434.400 13.050 435.450 ;
        RECT 1.950 433.950 4.050 434.400 ;
        RECT 10.950 433.950 13.050 434.400 ;
        RECT 73.950 435.450 76.050 436.050 ;
        RECT 88.950 435.450 91.050 436.050 ;
        RECT 73.950 434.400 91.050 435.450 ;
        RECT 73.950 433.950 76.050 434.400 ;
        RECT 88.950 433.950 91.050 434.400 ;
        RECT 247.950 435.450 250.050 436.050 ;
        RECT 391.950 435.450 394.050 436.050 ;
        RECT 442.950 435.450 445.050 436.050 ;
        RECT 247.950 434.400 381.450 435.450 ;
        RECT 247.950 433.950 250.050 434.400 ;
        RECT 289.950 432.450 292.050 433.050 ;
        RECT 346.950 432.450 349.050 433.050 ;
        RECT 289.950 431.400 349.050 432.450 ;
        RECT 380.400 432.450 381.450 434.400 ;
        RECT 391.950 434.400 445.050 435.450 ;
        RECT 391.950 433.950 394.050 434.400 ;
        RECT 442.950 433.950 445.050 434.400 ;
        RECT 454.950 435.450 457.050 436.050 ;
        RECT 517.950 435.450 520.050 436.050 ;
        RECT 454.950 434.400 520.050 435.450 ;
        RECT 454.950 433.950 457.050 434.400 ;
        RECT 517.950 433.950 520.050 434.400 ;
        RECT 586.950 435.450 589.050 436.050 ;
        RECT 637.950 435.450 640.050 436.050 ;
        RECT 586.950 434.400 640.050 435.450 ;
        RECT 586.950 433.950 589.050 434.400 ;
        RECT 637.950 433.950 640.050 434.400 ;
        RECT 646.950 435.450 649.050 436.050 ;
        RECT 670.950 435.450 673.050 436.050 ;
        RECT 646.950 434.400 673.050 435.450 ;
        RECT 646.950 433.950 649.050 434.400 ;
        RECT 670.950 433.950 673.050 434.400 ;
        RECT 676.950 435.450 679.050 436.050 ;
        RECT 718.950 435.450 721.050 436.050 ;
        RECT 808.950 435.450 811.050 436.050 ;
        RECT 676.950 434.400 721.050 435.450 ;
        RECT 676.950 433.950 679.050 434.400 ;
        RECT 718.950 433.950 721.050 434.400 ;
        RECT 785.400 434.400 811.050 435.450 ;
        RECT 406.950 432.450 409.050 433.050 ;
        RECT 451.950 432.450 454.050 433.050 ;
        RECT 380.400 431.400 454.050 432.450 ;
        RECT 289.950 430.950 292.050 431.400 ;
        RECT 346.950 430.950 349.050 431.400 ;
        RECT 406.950 430.950 409.050 431.400 ;
        RECT 451.950 430.950 454.050 431.400 ;
        RECT 466.950 432.450 469.050 433.050 ;
        RECT 556.950 432.450 559.050 433.050 ;
        RECT 466.950 431.400 559.050 432.450 ;
        RECT 466.950 430.950 469.050 431.400 ;
        RECT 556.950 430.950 559.050 431.400 ;
        RECT 565.950 432.450 568.050 433.050 ;
        RECT 577.950 432.450 580.050 433.050 ;
        RECT 619.800 432.450 621.900 433.050 ;
        RECT 565.950 431.400 580.050 432.450 ;
        RECT 565.950 430.950 568.050 431.400 ;
        RECT 577.950 430.950 580.050 431.400 ;
        RECT 608.400 431.400 621.900 432.450 ;
        RECT 124.950 429.450 127.050 430.050 ;
        RECT 139.800 429.450 141.900 430.050 ;
        RECT 124.950 428.400 141.900 429.450 ;
        RECT 124.950 427.950 127.050 428.400 ;
        RECT 139.800 427.950 141.900 428.400 ;
        RECT 143.100 429.450 145.200 430.050 ;
        RECT 148.950 429.450 151.050 430.050 ;
        RECT 143.100 428.400 151.050 429.450 ;
        RECT 143.100 427.950 145.200 428.400 ;
        RECT 148.950 427.950 151.050 428.400 ;
        RECT 160.950 429.450 163.050 430.050 ;
        RECT 169.950 429.450 172.050 430.050 ;
        RECT 241.950 429.450 244.050 430.050 ;
        RECT 160.950 428.400 244.050 429.450 ;
        RECT 160.950 427.950 163.050 428.400 ;
        RECT 169.950 427.950 172.050 428.400 ;
        RECT 241.950 427.950 244.050 428.400 ;
        RECT 253.950 429.450 256.050 430.050 ;
        RECT 280.950 429.450 283.050 430.050 ;
        RECT 319.950 429.450 322.050 430.050 ;
        RECT 253.950 428.400 322.050 429.450 ;
        RECT 253.950 427.950 256.050 428.400 ;
        RECT 280.950 427.950 283.050 428.400 ;
        RECT 319.950 427.950 322.050 428.400 ;
        RECT 325.950 429.450 328.050 430.050 ;
        RECT 352.950 429.450 355.050 430.050 ;
        RECT 325.950 428.400 355.050 429.450 ;
        RECT 325.950 427.950 328.050 428.400 ;
        RECT 352.950 427.950 355.050 428.400 ;
        RECT 463.950 429.450 466.050 430.050 ;
        RECT 496.800 429.450 498.900 430.050 ;
        RECT 463.950 428.400 498.900 429.450 ;
        RECT 463.950 427.950 466.050 428.400 ;
        RECT 496.800 427.950 498.900 428.400 ;
        RECT 500.100 429.450 502.200 430.050 ;
        RECT 517.950 429.450 520.050 430.050 ;
        RECT 500.100 428.400 520.050 429.450 ;
        RECT 500.100 427.950 502.200 428.400 ;
        RECT 517.950 427.950 520.050 428.400 ;
        RECT 565.950 429.450 568.050 430.050 ;
        RECT 608.400 429.450 609.450 431.400 ;
        RECT 619.800 430.950 621.900 431.400 ;
        RECT 623.100 432.450 625.200 433.050 ;
        RECT 655.950 432.450 658.050 433.050 ;
        RECT 623.100 431.400 658.050 432.450 ;
        RECT 623.100 430.950 625.200 431.400 ;
        RECT 655.950 430.950 658.050 431.400 ;
        RECT 661.950 432.450 664.050 433.050 ;
        RECT 748.950 432.450 751.050 433.050 ;
        RECT 661.950 431.400 751.050 432.450 ;
        RECT 661.950 430.950 664.050 431.400 ;
        RECT 748.950 430.950 751.050 431.400 ;
        RECT 760.950 432.450 763.050 433.050 ;
        RECT 785.400 432.450 786.450 434.400 ;
        RECT 808.950 433.950 811.050 434.400 ;
        RECT 760.950 431.400 786.450 432.450 ;
        RECT 787.950 432.450 790.050 433.050 ;
        RECT 802.950 432.450 805.050 433.050 ;
        RECT 787.950 431.400 805.050 432.450 ;
        RECT 760.950 430.950 763.050 431.400 ;
        RECT 787.950 430.950 790.050 431.400 ;
        RECT 802.950 430.950 805.050 431.400 ;
        RECT 697.950 429.450 700.050 430.050 ;
        RECT 565.950 428.400 609.450 429.450 ;
        RECT 611.400 428.400 700.050 429.450 ;
        RECT 565.950 427.950 568.050 428.400 ;
        RECT 19.950 426.450 22.050 427.050 ;
        RECT 31.950 426.450 34.050 427.200 ;
        RECT 19.950 425.400 34.050 426.450 ;
        RECT 19.950 424.950 22.050 425.400 ;
        RECT 31.950 425.100 34.050 425.400 ;
        RECT 130.950 426.450 133.050 427.050 ;
        RECT 136.950 426.450 139.050 427.050 ;
        RECT 190.950 426.450 193.050 427.050 ;
        RECT 130.950 425.400 193.050 426.450 ;
        RECT 130.950 424.950 133.050 425.400 ;
        RECT 136.950 424.950 139.050 425.400 ;
        RECT 190.950 424.950 193.050 425.400 ;
        RECT 295.950 426.450 298.050 427.050 ;
        RECT 322.950 426.450 325.050 427.050 ;
        RECT 340.950 426.450 343.050 427.050 ;
        RECT 295.950 425.400 325.050 426.450 ;
        RECT 295.950 424.950 298.050 425.400 ;
        RECT 322.950 424.950 325.050 425.400 ;
        RECT 326.400 425.400 343.050 426.450 ;
        RECT 7.950 423.450 10.050 424.050 ;
        RECT 25.950 423.450 28.050 424.050 ;
        RECT 31.950 423.450 34.050 423.900 ;
        RECT 7.950 422.400 34.050 423.450 ;
        RECT 7.950 421.950 10.050 422.400 ;
        RECT 25.950 421.950 28.050 422.400 ;
        RECT 31.950 421.800 34.050 422.400 ;
        RECT 79.950 423.450 82.050 424.050 ;
        RECT 118.950 423.450 121.050 424.050 ;
        RECT 157.950 423.450 160.050 424.050 ;
        RECT 184.950 423.450 187.050 424.050 ;
        RECT 259.950 423.450 262.050 424.050 ;
        RECT 79.950 422.400 121.050 423.450 ;
        RECT 79.950 421.950 82.050 422.400 ;
        RECT 118.950 421.950 121.050 422.400 ;
        RECT 122.400 422.400 160.050 423.450 ;
        RECT 25.950 417.450 28.050 418.050 ;
        RECT 17.550 417.000 28.050 417.450 ;
        RECT 16.950 416.400 28.050 417.000 ;
        RECT 16.950 415.050 19.050 416.400 ;
        RECT 25.950 415.950 28.050 416.400 ;
        RECT 31.950 415.950 34.050 421.050 ;
        RECT 43.950 420.450 46.050 421.050 ;
        RECT 55.950 420.450 58.050 421.050 ;
        RECT 38.400 420.000 58.050 420.450 ;
        RECT 37.950 419.400 58.050 420.000 ;
        RECT 37.950 415.950 40.050 419.400 ;
        RECT 43.950 418.950 46.050 419.400 ;
        RECT 55.950 418.950 58.050 419.400 ;
        RECT 73.950 420.450 76.050 421.050 ;
        RECT 122.400 420.450 123.450 422.400 ;
        RECT 157.950 421.950 160.050 422.400 ;
        RECT 161.400 422.400 262.050 423.450 ;
        RECT 73.950 419.400 123.450 420.450 ;
        RECT 73.950 418.950 76.050 419.400 ;
        RECT 161.400 418.050 162.450 422.400 ;
        RECT 184.950 421.950 187.050 422.400 ;
        RECT 259.950 421.950 262.050 422.400 ;
        RECT 286.950 423.450 289.050 424.050 ;
        RECT 313.800 423.450 315.900 424.050 ;
        RECT 286.950 422.400 315.900 423.450 ;
        RECT 286.950 421.950 289.050 422.400 ;
        RECT 313.800 421.950 315.900 422.400 ;
        RECT 317.100 423.450 319.200 424.050 ;
        RECT 326.400 423.450 327.450 425.400 ;
        RECT 340.950 424.950 343.050 425.400 ;
        RECT 370.950 426.450 373.050 427.050 ;
        RECT 376.950 426.450 379.050 427.050 ;
        RECT 370.950 425.400 379.050 426.450 ;
        RECT 370.950 424.950 373.050 425.400 ;
        RECT 376.950 424.950 379.050 425.400 ;
        RECT 400.950 426.450 403.050 427.050 ;
        RECT 436.950 426.450 439.050 427.050 ;
        RECT 400.950 425.400 439.050 426.450 ;
        RECT 514.950 426.450 517.050 427.050 ;
        RECT 559.950 426.450 562.050 427.050 ;
        RECT 514.950 425.400 562.050 426.450 ;
        RECT 400.950 424.950 403.050 425.400 ;
        RECT 436.950 424.950 439.050 425.400 ;
        RECT 317.100 422.400 327.450 423.450 ;
        RECT 337.950 423.450 340.050 424.050 ;
        RECT 385.950 423.450 388.050 424.050 ;
        RECT 337.950 422.400 388.050 423.450 ;
        RECT 475.950 423.300 478.050 425.400 ;
        RECT 514.950 424.950 517.050 425.400 ;
        RECT 559.950 424.950 562.050 425.400 ;
        RECT 565.950 426.450 568.050 427.050 ;
        RECT 611.400 426.450 612.450 428.400 ;
        RECT 697.950 427.950 700.050 428.400 ;
        RECT 709.950 429.450 712.050 430.050 ;
        RECT 739.950 429.450 742.050 430.050 ;
        RECT 769.950 429.450 772.050 430.050 ;
        RECT 709.950 428.400 772.050 429.450 ;
        RECT 709.950 427.950 712.050 428.400 ;
        RECT 739.950 427.950 742.050 428.400 ;
        RECT 769.950 427.950 772.050 428.400 ;
        RECT 775.950 429.450 778.050 430.050 ;
        RECT 784.950 429.450 787.050 430.050 ;
        RECT 775.950 428.400 787.050 429.450 ;
        RECT 775.950 427.950 778.050 428.400 ;
        RECT 784.950 427.950 787.050 428.400 ;
        RECT 565.950 425.400 612.450 426.450 ;
        RECT 613.950 426.450 616.050 427.050 ;
        RECT 706.950 426.450 709.050 427.050 ;
        RECT 736.950 426.450 739.050 427.050 ;
        RECT 613.950 425.400 739.050 426.450 ;
        RECT 565.950 424.950 568.050 425.400 ;
        RECT 613.950 424.950 616.050 425.400 ;
        RECT 706.950 424.950 709.050 425.400 ;
        RECT 736.950 424.950 739.050 425.400 ;
        RECT 317.100 421.950 319.200 422.400 ;
        RECT 337.950 421.950 340.050 422.400 ;
        RECT 385.950 421.950 388.050 422.400 ;
        RECT 55.950 417.450 58.050 418.050 ;
        RECT 41.400 417.000 58.050 417.450 ;
        RECT 40.950 416.400 58.050 417.000 ;
        RECT 7.950 412.950 12.900 415.050 ;
        RECT 13.800 414.000 15.900 415.050 ;
        RECT 16.950 414.000 19.200 415.050 ;
        RECT 33.000 414.900 37.050 415.050 ;
        RECT 13.800 412.950 16.050 414.000 ;
        RECT 17.100 412.950 19.200 414.000 ;
        RECT 31.950 412.950 37.050 414.900 ;
        RECT 40.950 412.950 43.050 416.400 ;
        RECT 55.950 415.950 58.050 416.400 ;
        RECT 55.950 412.950 60.900 415.050 ;
        RECT 62.100 414.450 64.200 415.050 ;
        RECT 67.950 414.450 70.050 415.050 ;
        RECT 62.100 413.400 70.050 414.450 ;
        RECT 62.100 412.950 64.200 413.400 ;
        RECT 67.950 412.950 70.050 413.400 ;
        RECT 73.950 412.950 76.050 418.050 ;
        RECT 79.950 412.950 82.050 418.050 ;
        RECT 142.800 417.450 144.900 418.050 ;
        RECT 116.400 417.000 144.900 417.450 ;
        RECT 115.950 416.400 144.900 417.000 ;
        RECT 88.950 414.450 91.050 415.050 ;
        RECT 97.950 414.450 100.050 415.050 ;
        RECT 109.950 414.450 112.050 415.050 ;
        RECT 88.950 413.400 112.050 414.450 ;
        RECT 88.950 412.950 91.050 413.400 ;
        RECT 97.950 412.950 100.050 413.400 ;
        RECT 109.950 412.950 112.050 413.400 ;
        RECT 115.950 412.950 118.050 416.400 ;
        RECT 130.950 412.950 133.050 416.400 ;
        RECT 142.800 415.950 144.900 416.400 ;
        RECT 146.100 417.450 148.200 418.050 ;
        RECT 151.950 417.450 154.050 418.050 ;
        RECT 146.100 416.400 154.050 417.450 ;
        RECT 146.100 415.950 148.200 416.400 ;
        RECT 151.950 415.950 154.050 416.400 ;
        RECT 157.950 416.400 162.450 418.050 ;
        RECT 157.950 415.950 162.000 416.400 ;
        RECT 166.950 415.950 169.050 421.050 ;
        RECT 181.950 420.450 184.050 421.050 ;
        RECT 304.950 420.450 307.050 421.050 ;
        RECT 370.950 420.450 373.050 421.050 ;
        RECT 173.400 420.000 184.050 420.450 ;
        RECT 293.400 420.000 373.050 420.450 ;
        RECT 172.950 419.400 184.050 420.000 ;
        RECT 172.950 415.950 175.050 419.400 ;
        RECT 181.950 418.950 184.050 419.400 ;
        RECT 292.950 419.400 373.050 420.000 ;
        RECT 184.950 415.050 187.050 418.050 ;
        RECT 190.950 417.450 193.050 418.050 ;
        RECT 208.950 417.450 211.050 418.050 ;
        RECT 250.950 417.450 253.050 418.050 ;
        RECT 277.950 417.450 280.050 418.050 ;
        RECT 190.950 416.400 280.050 417.450 ;
        RECT 190.950 415.950 193.050 416.400 ;
        RECT 208.950 415.950 211.050 416.400 ;
        RECT 136.950 412.950 142.050 415.050 ;
        RECT 145.950 414.450 148.050 415.050 ;
        RECT 154.800 414.450 156.900 415.050 ;
        RECT 145.950 413.400 156.900 414.450 ;
        RECT 145.950 412.950 148.050 413.400 ;
        RECT 154.800 412.950 156.900 413.400 ;
        RECT 158.100 414.450 160.200 415.050 ;
        RECT 169.950 414.450 172.050 415.050 ;
        RECT 158.100 413.400 172.050 414.450 ;
        RECT 158.100 412.950 160.200 413.400 ;
        RECT 169.950 412.950 172.050 413.400 ;
        RECT 184.800 414.000 187.050 415.050 ;
        RECT 184.800 412.950 186.900 414.000 ;
        RECT 188.100 412.950 193.050 415.050 ;
        RECT 217.950 414.450 220.050 415.050 ;
        RECT 226.950 414.450 229.050 415.050 ;
        RECT 217.950 413.400 229.050 414.450 ;
        RECT 217.950 412.950 220.050 413.400 ;
        RECT 226.950 412.950 229.050 413.400 ;
        RECT 232.950 412.950 235.050 416.400 ;
        RECT 250.950 415.950 253.050 416.400 ;
        RECT 277.950 415.950 280.050 416.400 ;
        RECT 283.950 415.950 289.050 418.050 ;
        RECT 292.950 415.950 295.050 419.400 ;
        RECT 304.950 418.950 307.050 419.400 ;
        RECT 370.950 418.950 373.050 419.400 ;
        RECT 427.950 420.450 430.050 421.050 ;
        RECT 448.950 420.450 451.050 421.050 ;
        RECT 427.950 419.400 451.050 420.450 ;
        RECT 476.850 419.700 478.050 423.300 ;
        RECT 496.950 422.400 499.050 424.500 ;
        RECT 535.950 423.450 538.050 424.050 ;
        RECT 547.950 423.450 550.050 424.050 ;
        RECT 535.950 422.400 550.050 423.450 ;
        RECT 427.950 418.950 430.050 419.400 ;
        RECT 448.950 418.950 451.050 419.400 ;
        RECT 316.950 417.450 319.050 418.050 ;
        RECT 311.400 417.000 319.050 417.450 ;
        RECT 310.950 416.400 319.050 417.000 ;
        RECT 13.950 412.050 16.050 412.950 ;
        RECT 31.950 412.800 34.050 412.950 ;
        RECT 13.800 411.000 16.050 412.050 ;
        RECT 13.800 409.950 15.900 411.000 ;
        RECT 19.950 409.950 24.900 412.050 ;
        RECT 26.100 411.450 28.200 412.050 ;
        RECT 43.950 411.450 46.050 412.050 ;
        RECT 49.950 411.450 52.050 412.050 ;
        RECT 26.100 410.400 52.050 411.450 ;
        RECT 26.100 409.950 28.200 410.400 ;
        RECT 43.950 409.950 46.050 410.400 ;
        RECT 49.950 409.950 52.050 410.400 ;
        RECT 55.950 409.950 61.050 412.050 ;
        RECT 64.950 411.450 67.050 412.050 ;
        RECT 76.950 411.450 79.050 412.050 ;
        RECT 64.950 410.400 79.050 411.450 ;
        RECT 64.950 409.950 67.050 410.400 ;
        RECT 76.950 409.950 79.050 410.400 ;
        RECT 82.950 406.950 85.050 412.050 ;
        RECT 97.950 406.950 100.050 412.050 ;
        RECT 109.950 409.950 115.050 412.050 ;
        RECT 118.950 411.450 121.050 412.050 ;
        RECT 127.950 411.450 132.900 412.050 ;
        RECT 118.950 410.400 132.900 411.450 ;
        RECT 134.100 411.000 136.200 412.050 ;
        RECT 118.950 409.950 121.050 410.400 ;
        RECT 127.950 409.950 132.900 410.400 ;
        RECT 133.950 409.950 136.200 411.000 ;
        RECT 202.950 411.450 205.050 412.050 ;
        RECT 214.950 411.450 217.050 412.050 ;
        RECT 223.800 411.450 225.900 412.050 ;
        RECT 202.950 410.400 225.900 411.450 ;
        RECT 202.950 409.950 205.050 410.400 ;
        RECT 214.950 409.950 217.050 410.400 ;
        RECT 223.800 409.950 225.900 410.400 ;
        RECT 227.100 409.950 232.050 412.050 ;
        RECT 133.950 408.450 136.050 409.950 ;
        RECT 101.400 408.000 136.050 408.450 ;
        RECT 145.950 408.450 148.050 409.050 ;
        RECT 151.800 408.450 153.900 409.050 ;
        RECT 101.400 407.400 135.450 408.000 ;
        RECT 145.950 407.400 153.900 408.450 ;
        RECT 34.950 405.450 37.050 406.050 ;
        RECT 67.950 405.450 70.050 406.050 ;
        RECT 101.400 405.450 102.450 407.400 ;
        RECT 145.950 406.950 148.050 407.400 ;
        RECT 151.800 406.950 153.900 407.400 ;
        RECT 155.100 408.450 157.200 409.050 ;
        RECT 166.950 408.450 169.050 409.050 ;
        RECT 199.950 408.450 202.050 409.050 ;
        RECT 155.100 407.400 202.050 408.450 ;
        RECT 235.950 408.450 238.050 412.050 ;
        RECT 247.950 409.950 250.050 415.050 ;
        RECT 253.950 414.450 256.050 415.050 ;
        RECT 280.950 414.450 283.050 415.050 ;
        RECT 253.950 413.400 283.050 414.450 ;
        RECT 253.950 412.950 256.050 413.400 ;
        RECT 280.950 412.950 283.050 413.400 ;
        RECT 252.000 411.450 256.050 412.050 ;
        RECT 251.400 409.950 256.050 411.450 ;
        RECT 241.950 408.450 244.050 409.050 ;
        RECT 251.400 408.450 252.450 409.950 ;
        RECT 256.950 408.450 259.050 409.050 ;
        RECT 235.950 408.000 259.050 408.450 ;
        RECT 236.400 407.400 259.050 408.000 ;
        RECT 155.100 406.950 157.200 407.400 ;
        RECT 166.950 406.950 169.050 407.400 ;
        RECT 199.950 406.950 202.050 407.400 ;
        RECT 241.950 406.950 244.050 407.400 ;
        RECT 256.950 406.950 259.050 407.400 ;
        RECT 265.950 406.950 268.050 412.050 ;
        RECT 271.950 409.950 277.050 412.050 ;
        RECT 289.950 409.950 292.050 415.050 ;
        RECT 298.950 414.450 301.050 415.050 ;
        RECT 304.950 414.450 307.050 415.050 ;
        RECT 298.950 413.400 307.050 414.450 ;
        RECT 298.950 412.950 301.050 413.400 ;
        RECT 304.950 412.950 307.050 413.400 ;
        RECT 310.950 412.950 313.050 416.400 ;
        RECT 316.950 415.950 319.050 416.400 ;
        RECT 322.950 415.950 327.900 418.050 ;
        RECT 329.100 417.450 331.200 418.050 ;
        RECT 337.950 417.450 340.050 418.050 ;
        RECT 329.100 416.400 340.050 417.450 ;
        RECT 329.100 415.950 331.200 416.400 ;
        RECT 337.950 415.950 340.050 416.400 ;
        RECT 355.950 417.450 358.050 418.050 ;
        RECT 361.800 417.450 363.900 418.050 ;
        RECT 355.950 416.400 363.900 417.450 ;
        RECT 355.950 415.950 358.050 416.400 ;
        RECT 361.800 415.950 363.900 416.400 ;
        RECT 365.100 415.950 370.050 418.050 ;
        RECT 379.950 417.450 382.050 418.050 ;
        RECT 388.950 417.450 391.050 418.050 ;
        RECT 379.950 416.400 391.050 417.450 ;
        RECT 379.950 415.950 382.050 416.400 ;
        RECT 388.950 415.950 391.050 416.400 ;
        RECT 322.950 412.950 328.050 415.050 ;
        RECT 298.950 411.450 301.050 412.050 ;
        RECT 307.950 411.450 310.050 412.050 ;
        RECT 298.950 410.400 310.050 411.450 ;
        RECT 298.950 409.950 301.050 410.400 ;
        RECT 307.950 409.950 310.050 410.400 ;
        RECT 313.950 409.950 319.050 412.050 ;
        RECT 346.950 409.950 349.050 415.050 ;
        RECT 364.950 414.450 367.050 415.050 ;
        RECT 379.950 414.450 382.050 415.050 ;
        RECT 364.950 413.400 382.050 414.450 ;
        RECT 364.950 412.950 367.050 413.400 ;
        RECT 379.950 412.950 382.050 413.400 ;
        RECT 385.950 412.050 388.050 415.050 ;
        RECT 412.950 414.450 415.050 415.050 ;
        RECT 421.950 414.450 424.050 415.050 ;
        RECT 412.950 413.400 424.050 414.450 ;
        RECT 412.950 412.950 415.050 413.400 ;
        RECT 421.950 412.950 424.050 413.400 ;
        RECT 427.950 412.950 430.050 418.050 ;
        RECT 439.950 412.950 445.050 415.050 ;
        RECT 448.950 414.450 451.050 415.050 ;
        RECT 454.950 414.450 457.050 415.050 ;
        RECT 448.950 413.400 457.050 414.450 ;
        RECT 448.950 412.950 451.050 413.400 ;
        RECT 454.950 412.950 457.050 413.400 ;
        RECT 463.950 412.950 466.050 418.050 ;
        RECT 475.950 417.600 478.050 419.700 ;
        RECT 352.950 409.950 358.050 412.050 ;
        RECT 379.950 409.950 384.900 412.050 ;
        RECT 385.950 411.000 388.200 412.050 ;
        RECT 386.100 409.950 388.200 411.000 ;
        RECT 280.950 408.450 283.050 409.050 ;
        RECT 292.950 408.450 295.050 409.050 ;
        RECT 280.950 407.400 295.050 408.450 ;
        RECT 280.950 406.950 283.050 407.400 ;
        RECT 292.950 406.950 295.050 407.400 ;
        RECT 409.950 406.950 412.050 412.050 ;
        RECT 415.950 409.950 421.050 412.050 ;
        RECT 424.950 409.950 427.050 412.050 ;
        RECT 433.950 411.450 436.050 412.050 ;
        RECT 439.950 411.450 442.050 412.050 ;
        RECT 433.950 410.400 442.050 411.450 ;
        RECT 433.950 409.950 436.050 410.400 ;
        RECT 439.950 409.950 442.050 410.400 ;
        RECT 445.950 409.950 451.050 412.050 ;
        RECT 34.950 404.400 102.450 405.450 ;
        RECT 298.950 405.450 301.050 406.050 ;
        RECT 328.950 405.450 331.050 406.050 ;
        RECT 298.950 404.400 331.050 405.450 ;
        RECT 34.950 403.950 37.050 404.400 ;
        RECT 67.950 403.950 70.050 404.400 ;
        RECT 298.950 403.950 301.050 404.400 ;
        RECT 328.950 403.950 331.050 404.400 ;
        RECT 340.950 405.450 343.050 406.050 ;
        RECT 358.950 405.450 361.050 406.050 ;
        RECT 340.950 404.400 361.050 405.450 ;
        RECT 340.950 403.950 343.050 404.400 ;
        RECT 358.950 403.950 361.050 404.400 ;
        RECT 394.950 405.450 397.050 406.050 ;
        RECT 415.950 405.450 418.050 406.050 ;
        RECT 394.950 404.400 418.050 405.450 ;
        RECT 425.400 405.450 426.450 409.950 ;
        RECT 427.950 408.450 430.050 409.050 ;
        RECT 466.950 408.450 469.050 409.050 ;
        RECT 472.950 408.450 475.050 409.050 ;
        RECT 427.950 407.400 475.050 408.450 ;
        RECT 427.950 406.950 430.050 407.400 ;
        RECT 466.950 406.950 469.050 407.400 ;
        RECT 472.950 406.950 475.050 407.400 ;
        RECT 442.950 405.450 445.050 406.050 ;
        RECT 476.850 405.600 478.050 417.600 ;
        RECT 484.950 406.950 487.050 412.050 ;
        RECT 490.950 406.950 493.050 412.050 ;
        RECT 497.100 405.600 498.300 422.400 ;
        RECT 535.950 421.950 538.050 422.400 ;
        RECT 547.950 421.950 550.050 422.400 ;
        RECT 556.950 423.450 559.050 424.050 ;
        RECT 571.950 423.450 574.050 424.050 ;
        RECT 556.950 422.400 574.050 423.450 ;
        RECT 556.950 421.950 559.050 422.400 ;
        RECT 571.950 421.950 574.050 422.400 ;
        RECT 601.950 423.450 604.050 424.050 ;
        RECT 721.950 423.450 724.050 424.050 ;
        RECT 733.950 423.450 736.050 424.050 ;
        RECT 601.950 422.400 657.450 423.450 ;
        RECT 601.950 421.950 604.050 422.400 ;
        RECT 499.950 420.450 502.050 421.050 ;
        RECT 505.950 420.450 508.050 421.050 ;
        RECT 499.950 419.400 508.050 420.450 ;
        RECT 499.950 418.950 502.050 419.400 ;
        RECT 505.950 418.950 508.050 419.400 ;
        RECT 532.950 420.450 535.050 421.050 ;
        RECT 541.950 420.450 544.050 421.050 ;
        RECT 532.950 419.400 544.050 420.450 ;
        RECT 532.950 418.950 535.050 419.400 ;
        RECT 541.950 418.950 544.050 419.400 ;
        RECT 550.950 420.450 553.050 421.050 ;
        RECT 580.950 420.450 583.050 421.050 ;
        RECT 550.950 419.400 583.050 420.450 ;
        RECT 550.950 418.950 553.050 419.400 ;
        RECT 580.950 418.950 583.050 419.400 ;
        RECT 589.950 420.450 592.050 421.050 ;
        RECT 607.950 420.450 610.050 421.050 ;
        RECT 589.950 419.400 610.050 420.450 ;
        RECT 589.950 418.950 592.050 419.400 ;
        RECT 607.950 418.950 610.050 419.400 ;
        RECT 613.950 420.450 616.050 421.050 ;
        RECT 656.400 420.450 657.450 422.400 ;
        RECT 721.950 422.400 736.050 423.450 ;
        RECT 721.950 421.950 724.050 422.400 ;
        RECT 733.950 421.950 736.050 422.400 ;
        RECT 799.950 423.450 802.050 424.050 ;
        RECT 805.950 423.450 808.050 424.050 ;
        RECT 832.950 423.450 835.050 424.050 ;
        RECT 799.950 422.400 808.050 423.450 ;
        RECT 799.950 421.950 802.050 422.400 ;
        RECT 805.950 421.950 808.050 422.400 ;
        RECT 809.400 422.400 835.050 423.450 ;
        RECT 667.950 420.450 670.050 421.050 ;
        RECT 676.950 420.450 679.050 421.050 ;
        RECT 613.950 419.400 642.450 420.450 ;
        RECT 656.400 419.400 660.450 420.450 ;
        RECT 613.950 418.950 616.050 419.400 ;
        RECT 529.950 417.450 532.050 418.050 ;
        RECT 515.400 417.000 532.050 417.450 ;
        RECT 514.950 416.400 532.050 417.000 ;
        RECT 514.950 412.950 517.050 416.400 ;
        RECT 529.950 415.950 532.050 416.400 ;
        RECT 538.950 415.050 541.050 418.050 ;
        RECT 583.950 417.450 586.050 418.050 ;
        RECT 589.950 417.450 592.050 418.050 ;
        RECT 583.950 416.400 592.050 417.450 ;
        RECT 583.950 415.950 586.050 416.400 ;
        RECT 589.950 415.950 592.050 416.400 ;
        RECT 520.950 414.450 523.050 415.050 ;
        RECT 535.800 414.450 537.900 415.050 ;
        RECT 520.950 413.400 537.900 414.450 ;
        RECT 538.950 414.000 541.200 415.050 ;
        RECT 520.950 412.950 523.050 413.400 ;
        RECT 535.800 412.950 537.900 413.400 ;
        RECT 539.100 412.950 541.200 414.000 ;
        RECT 499.950 411.450 502.050 412.050 ;
        RECT 517.950 411.450 520.050 412.050 ;
        RECT 499.950 410.400 520.050 411.450 ;
        RECT 499.950 409.950 502.050 410.400 ;
        RECT 517.950 409.950 520.050 410.400 ;
        RECT 547.950 411.450 550.050 412.200 ;
        RECT 553.950 411.450 556.050 412.050 ;
        RECT 547.950 410.400 556.050 411.450 ;
        RECT 547.950 410.100 550.050 410.400 ;
        RECT 553.950 409.950 556.050 410.400 ;
        RECT 559.950 409.950 562.050 415.050 ;
        RECT 589.950 412.950 595.050 415.050 ;
        RECT 595.950 414.450 598.050 418.050 ;
        RECT 601.950 414.450 604.050 415.050 ;
        RECT 595.950 414.000 604.050 414.450 ;
        RECT 596.400 413.400 604.050 414.000 ;
        RECT 601.950 412.050 604.050 413.400 ;
        RECT 607.950 412.950 610.050 418.050 ;
        RECT 613.950 412.950 619.050 415.050 ;
        RECT 628.950 412.950 634.050 415.050 ;
        RECT 637.950 412.950 640.050 418.050 ;
        RECT 641.400 417.450 642.450 419.400 ;
        RECT 659.400 417.450 660.450 419.400 ;
        RECT 667.950 419.400 679.050 420.450 ;
        RECT 667.950 418.950 670.050 419.400 ;
        RECT 676.950 418.950 679.050 419.400 ;
        RECT 700.950 420.450 703.050 421.050 ;
        RECT 778.950 420.450 781.050 421.050 ;
        RECT 809.400 420.450 810.450 422.400 ;
        RECT 832.950 421.950 835.050 422.400 ;
        RECT 856.950 423.450 859.050 424.050 ;
        RECT 856.950 422.400 867.450 423.450 ;
        RECT 856.950 421.950 859.050 422.400 ;
        RECT 700.950 419.400 744.450 420.450 ;
        RECT 700.950 418.950 703.050 419.400 ;
        RECT 673.950 417.450 676.050 418.050 ;
        RECT 641.400 416.400 657.450 417.450 ;
        RECT 659.400 416.400 676.050 417.450 ;
        RECT 743.400 417.450 744.450 419.400 ;
        RECT 778.950 419.400 810.450 420.450 ;
        RECT 811.950 420.450 814.050 421.050 ;
        RECT 811.950 420.000 822.450 420.450 ;
        RECT 811.950 419.400 823.050 420.000 ;
        RECT 778.950 418.950 781.050 419.400 ;
        RECT 811.950 418.950 814.050 419.400 ;
        RECT 754.800 417.450 756.900 418.050 ;
        RECT 743.400 416.400 756.900 417.450 ;
        RECT 649.950 412.950 655.050 415.050 ;
        RECT 656.400 412.050 657.450 416.400 ;
        RECT 673.950 415.950 676.050 416.400 ;
        RECT 754.800 415.950 756.900 416.400 ;
        RECT 758.100 415.950 763.050 418.050 ;
        RECT 802.950 415.950 808.050 418.050 ;
        RECT 820.950 415.950 823.050 419.400 ;
        RECT 826.950 415.950 829.050 421.050 ;
        RECT 658.950 414.450 661.050 415.050 ;
        RECT 676.950 414.450 679.050 415.050 ;
        RECT 658.950 413.400 679.050 414.450 ;
        RECT 658.950 412.950 661.050 413.400 ;
        RECT 676.950 412.950 679.050 413.400 ;
        RECT 691.800 414.000 693.900 415.050 ;
        RECT 691.800 412.950 694.050 414.000 ;
        RECT 695.100 412.950 700.050 415.050 ;
        RECT 703.950 414.450 706.050 415.050 ;
        RECT 712.950 414.450 715.050 415.050 ;
        RECT 703.950 413.400 715.050 414.450 ;
        RECT 703.950 412.950 706.050 413.400 ;
        RECT 712.950 412.950 715.050 413.400 ;
        RECT 718.950 412.950 724.050 415.050 ;
        RECT 739.950 414.450 742.050 415.050 ;
        RECT 754.800 414.450 756.900 415.050 ;
        RECT 739.950 413.400 756.900 414.450 ;
        RECT 739.950 412.950 742.050 413.400 ;
        RECT 754.800 412.950 756.900 413.400 ;
        RECT 758.100 414.450 760.200 415.050 ;
        RECT 775.800 414.450 777.900 415.050 ;
        RECT 758.100 413.400 777.900 414.450 ;
        RECT 758.100 412.950 760.200 413.400 ;
        RECT 775.800 412.950 777.900 413.400 ;
        RECT 808.950 412.950 814.050 415.050 ;
        RECT 817.950 414.450 820.050 415.050 ;
        RECT 823.800 414.450 825.900 415.050 ;
        RECT 817.950 413.400 825.900 414.450 ;
        RECT 817.950 412.950 820.050 413.400 ;
        RECT 823.800 412.950 825.900 413.400 ;
        RECT 827.100 414.450 829.200 415.050 ;
        RECT 844.950 414.450 850.050 415.050 ;
        RECT 827.100 413.400 850.050 414.450 ;
        RECT 827.100 412.950 829.200 413.400 ;
        RECT 844.950 412.950 850.050 413.400 ;
        RECT 691.950 412.050 694.050 412.950 ;
        RECT 565.950 409.950 571.050 412.050 ;
        RECT 574.950 409.950 580.050 412.050 ;
        RECT 601.950 411.000 606.900 412.050 ;
        RECT 602.400 410.400 606.900 411.000 ;
        RECT 603.000 409.950 606.900 410.400 ;
        RECT 608.100 409.950 613.050 412.050 ;
        RECT 625.950 409.950 631.050 412.050 ;
        RECT 633.000 411.450 637.050 412.050 ;
        RECT 632.400 409.950 637.050 411.450 ;
        RECT 547.950 408.450 550.050 408.900 ;
        RECT 556.950 408.450 559.050 409.050 ;
        RECT 547.950 407.400 559.050 408.450 ;
        RECT 547.950 406.800 550.050 407.400 ;
        RECT 556.950 406.950 559.050 407.400 ;
        RECT 619.950 408.450 622.050 409.050 ;
        RECT 632.400 408.450 633.450 409.950 ;
        RECT 619.950 407.400 633.450 408.450 ;
        RECT 619.950 406.950 622.050 407.400 ;
        RECT 640.950 406.950 643.050 412.050 ;
        RECT 649.950 408.450 652.050 412.050 ;
        RECT 655.950 409.950 658.050 412.050 ;
        RECT 679.950 411.450 682.050 412.050 ;
        RECT 688.800 411.450 690.900 412.050 ;
        RECT 679.950 410.400 690.900 411.450 ;
        RECT 679.950 409.950 682.050 410.400 ;
        RECT 688.800 409.950 690.900 410.400 ;
        RECT 691.800 411.000 694.050 412.050 ;
        RECT 695.100 411.450 697.200 412.050 ;
        RECT 700.950 411.450 703.050 412.050 ;
        RECT 691.800 409.950 693.900 411.000 ;
        RECT 695.100 410.400 703.050 411.450 ;
        RECT 695.100 409.950 697.200 410.400 ;
        RECT 700.950 409.950 703.050 410.400 ;
        RECT 709.950 411.450 712.050 412.050 ;
        RECT 715.950 411.450 718.050 412.050 ;
        RECT 709.950 410.400 718.050 411.450 ;
        RECT 734.100 411.000 736.200 412.050 ;
        RECT 709.950 409.950 712.050 410.400 ;
        RECT 715.950 409.950 718.050 410.400 ;
        RECT 733.950 409.950 736.200 411.000 ;
        RECT 751.950 411.450 754.050 412.050 ;
        RECT 772.950 411.450 775.050 412.050 ;
        RECT 778.950 411.450 781.050 412.050 ;
        RECT 751.950 410.400 781.050 411.450 ;
        RECT 751.950 409.950 754.050 410.400 ;
        RECT 772.950 409.950 775.050 410.400 ;
        RECT 778.950 409.950 781.050 410.400 ;
        RECT 790.950 411.450 793.050 412.050 ;
        RECT 802.950 411.450 805.050 412.050 ;
        RECT 790.950 410.400 805.050 411.450 ;
        RECT 790.950 409.950 793.050 410.400 ;
        RECT 802.950 409.950 805.050 410.400 ;
        RECT 832.950 411.450 835.050 412.050 ;
        RECT 838.950 411.450 841.050 412.050 ;
        RECT 866.400 411.450 867.450 422.400 ;
        RECT 832.950 410.400 841.050 411.450 ;
        RECT 832.950 409.950 835.050 410.400 ;
        RECT 838.950 409.950 841.050 410.400 ;
        RECT 863.400 410.400 867.450 411.450 ;
        RECT 661.950 408.450 664.050 409.050 ;
        RECT 649.950 408.000 664.050 408.450 ;
        RECT 650.400 407.400 664.050 408.000 ;
        RECT 680.400 408.450 681.450 409.950 ;
        RECT 703.950 408.450 706.050 409.050 ;
        RECT 680.400 407.400 706.050 408.450 ;
        RECT 661.950 406.950 664.050 407.400 ;
        RECT 703.950 406.950 706.050 407.400 ;
        RECT 718.950 408.450 721.050 409.050 ;
        RECT 733.950 408.450 736.050 409.950 ;
        RECT 718.950 408.000 736.050 408.450 ;
        RECT 844.950 408.450 847.050 409.050 ;
        RECT 850.950 408.450 853.050 409.050 ;
        RECT 718.950 407.400 735.600 408.000 ;
        RECT 844.950 407.400 853.050 408.450 ;
        RECT 718.950 406.950 721.050 407.400 ;
        RECT 844.950 406.950 847.050 407.400 ;
        RECT 850.950 406.950 853.050 407.400 ;
        RECT 425.400 404.400 445.050 405.450 ;
        RECT 394.950 403.950 397.050 404.400 ;
        RECT 415.950 403.950 418.050 404.400 ;
        RECT 442.950 403.950 445.050 404.400 ;
        RECT 475.950 403.500 478.050 405.600 ;
        RECT 496.950 403.500 499.050 405.600 ;
        RECT 511.950 405.450 514.050 406.050 ;
        RECT 565.950 405.450 568.050 406.050 ;
        RECT 511.950 404.400 568.050 405.450 ;
        RECT 511.950 403.950 514.050 404.400 ;
        RECT 565.950 403.950 568.050 404.400 ;
        RECT 589.950 405.450 592.050 406.050 ;
        RECT 625.950 405.450 628.050 406.050 ;
        RECT 589.950 404.400 628.050 405.450 ;
        RECT 589.950 403.950 592.050 404.400 ;
        RECT 625.950 403.950 628.050 404.400 ;
        RECT 706.950 403.950 712.050 406.050 ;
        RECT 778.950 405.450 781.050 406.050 ;
        RECT 784.950 405.450 787.050 406.050 ;
        RECT 778.950 404.400 787.050 405.450 ;
        RECT 778.950 403.950 781.050 404.400 ;
        RECT 784.950 403.950 787.050 404.400 ;
        RECT 409.950 402.450 412.050 403.050 ;
        RECT 427.950 402.450 430.050 403.050 ;
        RECT 409.950 401.400 430.050 402.450 ;
        RECT 409.950 400.950 412.050 401.400 ;
        RECT 427.950 400.950 430.050 401.400 ;
        RECT 439.950 402.450 442.050 403.050 ;
        RECT 457.950 402.450 460.050 403.050 ;
        RECT 439.950 401.400 460.050 402.450 ;
        RECT 439.950 400.950 442.050 401.400 ;
        RECT 457.950 400.950 460.050 401.400 ;
        RECT 508.950 402.450 511.050 403.050 ;
        RECT 574.950 402.450 577.050 403.050 ;
        RECT 508.950 401.400 577.050 402.450 ;
        RECT 508.950 400.950 511.050 401.400 ;
        RECT 574.950 400.950 577.050 401.400 ;
        RECT 607.950 402.450 610.050 403.050 ;
        RECT 637.800 402.450 639.900 403.050 ;
        RECT 607.950 401.400 639.900 402.450 ;
        RECT 607.950 400.950 610.050 401.400 ;
        RECT 637.800 400.950 639.900 401.400 ;
        RECT 641.100 402.450 643.200 403.050 ;
        RECT 688.950 402.450 691.050 403.050 ;
        RECT 641.100 401.400 691.050 402.450 ;
        RECT 641.100 400.950 643.200 401.400 ;
        RECT 688.950 400.950 691.050 401.400 ;
        RECT 694.950 402.450 697.050 403.050 ;
        RECT 718.950 402.450 721.050 403.050 ;
        RECT 694.950 401.400 721.050 402.450 ;
        RECT 694.950 400.950 697.050 401.400 ;
        RECT 718.950 400.950 721.050 401.400 ;
        RECT 748.950 402.450 751.050 403.050 ;
        RECT 799.800 402.450 801.900 403.050 ;
        RECT 748.950 401.400 801.900 402.450 ;
        RECT 748.950 400.950 751.050 401.400 ;
        RECT 799.800 400.950 801.900 401.400 ;
        RECT 803.100 402.450 805.200 403.050 ;
        RECT 817.950 402.450 820.050 403.050 ;
        RECT 803.100 401.400 820.050 402.450 ;
        RECT 803.100 400.950 805.200 401.400 ;
        RECT 817.950 400.950 820.050 401.400 ;
        RECT 850.950 400.950 856.050 403.050 ;
        RECT 247.950 399.450 250.050 400.050 ;
        RECT 271.950 399.450 274.050 400.050 ;
        RECT 247.950 398.400 274.050 399.450 ;
        RECT 247.950 397.950 250.050 398.400 ;
        RECT 271.950 397.950 274.050 398.400 ;
        RECT 277.950 399.450 280.050 400.050 ;
        RECT 346.950 399.450 349.050 400.050 ;
        RECT 277.950 398.400 349.050 399.450 ;
        RECT 277.950 397.950 280.050 398.400 ;
        RECT 346.950 397.950 349.050 398.400 ;
        RECT 385.950 399.450 388.050 400.050 ;
        RECT 493.950 399.450 496.050 400.050 ;
        RECT 385.950 398.400 496.050 399.450 ;
        RECT 385.950 397.950 388.050 398.400 ;
        RECT 493.950 397.950 496.050 398.400 ;
        RECT 514.950 399.450 517.050 400.050 ;
        RECT 565.950 399.450 568.050 400.050 ;
        RECT 514.950 398.400 568.050 399.450 ;
        RECT 514.950 397.950 517.050 398.400 ;
        RECT 565.950 397.950 568.050 398.400 ;
        RECT 628.950 399.450 631.050 400.050 ;
        RECT 646.950 399.450 649.050 400.050 ;
        RECT 703.950 399.450 706.050 400.050 ;
        RECT 628.950 398.400 706.050 399.450 ;
        RECT 628.950 397.950 631.050 398.400 ;
        RECT 646.950 397.950 649.050 398.400 ;
        RECT 703.950 397.950 706.050 398.400 ;
        RECT 712.950 399.450 715.050 400.050 ;
        RECT 730.950 399.450 733.050 400.050 ;
        RECT 712.950 398.400 733.050 399.450 ;
        RECT 712.950 397.950 715.050 398.400 ;
        RECT 730.950 397.950 733.050 398.400 ;
        RECT 742.950 399.450 745.050 400.050 ;
        RECT 772.800 399.450 774.900 400.050 ;
        RECT 742.950 398.400 774.900 399.450 ;
        RECT 742.950 397.950 745.050 398.400 ;
        RECT 772.800 397.950 774.900 398.400 ;
        RECT 776.100 399.450 778.200 400.050 ;
        RECT 787.950 399.450 790.050 400.050 ;
        RECT 776.100 398.400 790.050 399.450 ;
        RECT 776.100 397.950 778.200 398.400 ;
        RECT 787.950 397.950 790.050 398.400 ;
        RECT 94.950 396.450 97.050 397.050 ;
        RECT 50.400 396.000 97.050 396.450 ;
        RECT 49.950 395.400 97.050 396.000 ;
        RECT 49.950 391.950 52.050 395.400 ;
        RECT 94.950 394.950 97.050 395.400 ;
        RECT 106.950 396.450 109.050 397.050 ;
        RECT 124.950 396.450 127.050 397.050 ;
        RECT 106.950 395.400 127.050 396.450 ;
        RECT 106.950 394.950 109.050 395.400 ;
        RECT 124.950 394.950 127.050 395.400 ;
        RECT 151.950 396.450 154.050 397.050 ;
        RECT 217.950 396.450 220.050 397.050 ;
        RECT 253.950 396.450 256.050 397.050 ;
        RECT 151.950 395.400 256.050 396.450 ;
        RECT 151.950 394.950 154.050 395.400 ;
        RECT 217.950 394.950 220.050 395.400 ;
        RECT 253.950 394.950 256.050 395.400 ;
        RECT 265.950 396.450 268.050 397.050 ;
        RECT 373.950 396.450 376.050 397.050 ;
        RECT 265.950 395.400 376.050 396.450 ;
        RECT 265.950 394.950 268.050 395.400 ;
        RECT 373.950 394.950 376.050 395.400 ;
        RECT 436.950 396.450 439.050 397.050 ;
        RECT 454.950 396.450 457.050 397.050 ;
        RECT 436.950 395.400 457.050 396.450 ;
        RECT 436.950 394.950 439.050 395.400 ;
        RECT 454.950 394.950 457.050 395.400 ;
        RECT 460.950 396.450 463.050 397.050 ;
        RECT 484.950 396.450 487.050 397.050 ;
        RECT 460.950 395.400 487.050 396.450 ;
        RECT 460.950 394.950 463.050 395.400 ;
        RECT 484.950 394.950 487.050 395.400 ;
        RECT 490.950 396.450 493.050 397.050 ;
        RECT 499.950 396.450 502.050 397.050 ;
        RECT 511.950 396.450 514.050 397.050 ;
        RECT 490.950 395.400 502.050 396.450 ;
        RECT 490.950 394.950 493.050 395.400 ;
        RECT 499.950 394.950 502.050 395.400 ;
        RECT 503.400 395.400 514.050 396.450 ;
        RECT 64.950 393.450 67.050 394.050 ;
        RECT 85.950 393.450 88.050 394.050 ;
        RECT 64.950 392.400 88.050 393.450 ;
        RECT 64.950 391.950 67.050 392.400 ;
        RECT 85.950 391.950 88.050 392.400 ;
        RECT 118.950 393.450 121.050 394.050 ;
        RECT 145.950 393.450 148.050 394.050 ;
        RECT 118.950 392.400 148.050 393.450 ;
        RECT 118.950 391.950 121.050 392.400 ;
        RECT 145.950 391.950 148.050 392.400 ;
        RECT 178.950 391.950 184.050 394.050 ;
        RECT 208.950 393.450 211.050 394.050 ;
        RECT 226.950 393.450 229.050 394.050 ;
        RECT 208.950 392.400 229.050 393.450 ;
        RECT 208.950 391.950 211.050 392.400 ;
        RECT 226.950 391.950 229.050 392.400 ;
        RECT 241.950 393.450 244.050 394.050 ;
        RECT 322.950 393.450 325.050 394.050 ;
        RECT 241.950 392.400 325.050 393.450 ;
        RECT 241.950 391.950 244.050 392.400 ;
        RECT 322.950 391.950 325.050 392.400 ;
        RECT 352.950 391.950 358.050 394.050 ;
        RECT 367.950 393.450 370.050 394.050 ;
        RECT 418.950 393.450 421.050 394.050 ;
        RECT 367.950 392.400 421.050 393.450 ;
        RECT 367.950 391.950 370.050 392.400 ;
        RECT 418.950 391.950 421.050 392.400 ;
        RECT 424.950 393.450 427.050 394.050 ;
        RECT 430.950 393.450 433.050 394.050 ;
        RECT 424.950 392.400 433.050 393.450 ;
        RECT 424.950 391.950 427.050 392.400 ;
        RECT 430.950 391.950 433.050 392.400 ;
        RECT 481.950 393.450 484.050 394.050 ;
        RECT 503.400 393.450 504.450 395.400 ;
        RECT 511.950 394.950 514.050 395.400 ;
        RECT 529.950 396.450 532.050 397.050 ;
        RECT 643.950 396.450 646.050 397.050 ;
        RECT 529.950 395.400 646.050 396.450 ;
        RECT 529.950 394.950 532.050 395.400 ;
        RECT 643.950 394.950 646.050 395.400 ;
        RECT 808.950 396.450 811.050 397.050 ;
        RECT 820.950 396.450 823.050 397.050 ;
        RECT 808.950 395.400 823.050 396.450 ;
        RECT 808.950 394.950 811.050 395.400 ;
        RECT 820.950 394.950 823.050 395.400 ;
        RECT 481.950 392.400 504.450 393.450 ;
        RECT 505.950 393.450 508.050 394.050 ;
        RECT 514.950 393.450 517.050 394.050 ;
        RECT 505.950 392.400 517.050 393.450 ;
        RECT 481.950 391.950 484.050 392.400 ;
        RECT 505.950 391.950 508.050 392.400 ;
        RECT 514.950 391.950 517.050 392.400 ;
        RECT 535.950 393.450 538.050 394.050 ;
        RECT 544.950 393.450 547.050 394.200 ;
        RECT 535.950 392.400 547.050 393.450 ;
        RECT 535.950 391.950 538.050 392.400 ;
        RECT 544.950 392.100 547.050 392.400 ;
        RECT 589.950 393.450 592.050 394.050 ;
        RECT 607.800 393.450 609.900 394.050 ;
        RECT 589.950 392.400 609.900 393.450 ;
        RECT 589.950 391.950 592.050 392.400 ;
        RECT 607.800 391.950 609.900 392.400 ;
        RECT 611.100 393.450 613.200 394.050 ;
        RECT 658.950 393.450 661.050 394.050 ;
        RECT 611.100 392.400 661.050 393.450 ;
        RECT 611.100 391.950 613.200 392.400 ;
        RECT 658.950 391.950 661.050 392.400 ;
        RECT 688.950 393.450 691.050 394.050 ;
        RECT 760.950 393.450 763.050 394.050 ;
        RECT 688.950 392.400 763.050 393.450 ;
        RECT 688.950 391.950 691.050 392.400 ;
        RECT 760.950 391.950 763.050 392.400 ;
        RECT 853.950 393.450 856.050 394.050 ;
        RECT 863.400 393.450 864.450 410.400 ;
        RECT 853.950 392.400 864.450 393.450 ;
        RECT 853.950 391.950 856.050 392.400 ;
        RECT 19.950 390.450 22.050 391.050 ;
        RECT 25.950 390.450 28.050 391.050 ;
        RECT 19.950 389.400 28.050 390.450 ;
        RECT 19.950 388.950 22.050 389.400 ;
        RECT 25.950 388.950 28.050 389.400 ;
        RECT 73.950 390.450 76.050 391.050 ;
        RECT 73.950 389.400 87.450 390.450 ;
        RECT 73.950 388.950 76.050 389.400 ;
        RECT 13.950 387.450 16.050 388.050 ;
        RECT 13.950 386.400 30.450 387.450 ;
        RECT 13.950 385.950 16.050 386.400 ;
        RECT 29.400 385.050 30.450 386.400 ;
        RECT 43.950 385.950 48.900 388.050 ;
        RECT 50.100 387.450 52.200 388.050 ;
        RECT 50.100 386.400 78.450 387.450 ;
        RECT 50.100 385.950 52.200 386.400 ;
        RECT 77.400 385.050 78.450 386.400 ;
        RECT 86.400 385.050 87.450 389.400 ;
        RECT 127.950 388.950 133.050 391.050 ;
        RECT 253.950 390.450 256.050 391.050 ;
        RECT 265.950 390.450 268.050 391.050 ;
        RECT 212.400 390.000 268.050 390.450 ;
        RECT 211.950 389.400 268.050 390.000 ;
        RECT 112.950 387.450 115.050 388.050 ;
        RECT 104.400 387.000 115.050 387.450 ;
        RECT 103.950 386.400 115.050 387.000 ;
        RECT 13.950 379.950 16.050 385.050 ;
        RECT 19.950 381.450 22.050 385.050 ;
        RECT 28.800 384.000 30.900 385.050 ;
        RECT 32.100 384.000 34.200 385.050 ;
        RECT 28.800 382.950 31.050 384.000 ;
        RECT 28.950 382.050 31.050 382.950 ;
        RECT 25.800 381.450 27.900 382.050 ;
        RECT 19.950 380.400 27.900 381.450 ;
        RECT 19.950 379.950 22.050 380.400 ;
        RECT 25.800 379.950 27.900 380.400 ;
        RECT 28.800 381.000 31.050 382.050 ;
        RECT 31.950 382.950 34.200 384.000 ;
        RECT 40.950 384.450 43.050 385.050 ;
        RECT 46.800 384.450 48.900 385.050 ;
        RECT 40.950 383.400 48.900 384.450 ;
        RECT 40.950 382.950 43.050 383.400 ;
        RECT 46.800 382.950 48.900 383.400 ;
        RECT 50.100 384.450 52.200 385.050 ;
        RECT 58.950 384.450 61.050 385.050 ;
        RECT 70.950 384.450 76.050 385.050 ;
        RECT 50.100 384.000 57.450 384.450 ;
        RECT 50.100 383.400 58.050 384.000 ;
        RECT 50.100 382.950 52.200 383.400 ;
        RECT 31.950 382.050 34.050 382.950 ;
        RECT 31.950 381.000 34.200 382.050 ;
        RECT 28.800 379.950 30.900 381.000 ;
        RECT 32.100 379.950 34.200 381.000 ;
        RECT 35.100 381.450 37.200 382.050 ;
        RECT 49.950 381.450 52.050 382.050 ;
        RECT 35.100 380.400 52.050 381.450 ;
        RECT 35.100 379.950 37.200 380.400 ;
        RECT 49.950 379.950 52.050 380.400 ;
        RECT 55.950 379.950 58.050 383.400 ;
        RECT 58.950 383.400 76.050 384.450 ;
        RECT 77.400 383.400 82.050 385.050 ;
        RECT 58.950 382.950 61.050 383.400 ;
        RECT 70.950 382.950 76.050 383.400 ;
        RECT 78.000 382.950 82.050 383.400 ;
        RECT 85.950 382.950 88.050 385.050 ;
        RECT 91.950 382.950 97.050 385.050 ;
        RECT 103.950 382.950 106.050 386.400 ;
        RECT 112.950 385.950 115.050 386.400 ;
        RECT 118.950 385.950 124.050 388.050 ;
        RECT 139.950 387.450 142.050 388.050 ;
        RECT 172.950 387.450 175.050 388.050 ;
        RECT 139.950 386.400 175.050 387.450 ;
        RECT 139.950 385.950 142.050 386.400 ;
        RECT 172.950 385.950 175.050 386.400 ;
        RECT 205.950 387.450 208.050 388.050 ;
        RECT 211.950 387.450 214.050 389.400 ;
        RECT 253.950 388.950 256.050 389.400 ;
        RECT 265.950 388.950 268.050 389.400 ;
        RECT 280.950 390.450 283.050 391.050 ;
        RECT 295.950 390.450 298.050 391.050 ;
        RECT 280.950 389.400 298.050 390.450 ;
        RECT 280.950 388.950 283.050 389.400 ;
        RECT 295.950 388.950 298.050 389.400 ;
        RECT 319.950 390.450 322.050 391.050 ;
        RECT 334.950 390.450 337.050 391.050 ;
        RECT 319.950 389.400 337.050 390.450 ;
        RECT 319.950 388.950 322.050 389.400 ;
        RECT 334.950 388.950 337.050 389.400 ;
        RECT 364.950 390.450 367.050 391.050 ;
        RECT 382.950 390.450 385.050 391.050 ;
        RECT 364.950 389.400 385.050 390.450 ;
        RECT 454.950 389.400 457.050 391.500 ;
        RECT 475.950 389.400 478.050 391.500 ;
        RECT 502.950 390.450 505.050 391.050 ;
        RECT 517.950 390.450 520.050 391.050 ;
        RECT 502.950 389.400 520.050 390.450 ;
        RECT 364.950 388.950 367.050 389.400 ;
        RECT 382.950 388.950 385.050 389.400 ;
        RECT 205.950 386.400 214.050 387.450 ;
        RECT 205.950 385.950 208.050 386.400 ;
        RECT 211.950 385.950 214.050 386.400 ;
        RECT 226.950 385.950 232.050 388.050 ;
        RECT 265.950 385.050 268.050 388.050 ;
        RECT 286.950 387.450 292.050 388.050 ;
        RECT 328.950 387.450 331.050 388.050 ;
        RECT 286.950 386.400 309.450 387.450 ;
        RECT 323.400 387.000 331.050 387.450 ;
        RECT 286.950 385.950 292.050 386.400 ;
        RECT 61.950 381.450 67.050 382.050 ;
        RECT 76.950 381.450 79.050 382.050 ;
        RECT 61.950 380.400 79.050 381.450 ;
        RECT 61.950 379.950 67.050 380.400 ;
        RECT 76.950 379.950 79.050 380.400 ;
        RECT 4.950 376.950 10.050 379.050 ;
        RECT 16.950 378.450 19.050 379.050 ;
        RECT 31.950 378.450 34.050 379.050 ;
        RECT 49.950 378.450 52.050 379.050 ;
        RECT 16.950 377.400 52.050 378.450 ;
        RECT 16.950 376.950 19.050 377.400 ;
        RECT 31.950 376.950 34.050 377.400 ;
        RECT 49.950 376.950 52.050 377.400 ;
        RECT 46.950 370.950 49.050 376.050 ;
        RECT 58.950 373.950 61.050 379.050 ;
        RECT 82.950 376.950 85.050 382.050 ;
        RECT 100.950 376.950 103.050 382.050 ;
        RECT 106.950 376.950 109.050 382.050 ;
        RECT 127.950 381.450 130.050 382.050 ;
        RECT 136.950 381.450 139.050 382.050 ;
        RECT 127.950 380.400 139.050 381.450 ;
        RECT 127.950 379.950 130.050 380.400 ;
        RECT 136.950 379.950 139.050 380.400 ;
        RECT 154.950 379.950 157.050 385.050 ;
        RECT 169.950 382.950 174.900 385.050 ;
        RECT 176.100 384.450 178.200 385.050 ;
        RECT 196.950 384.450 199.050 385.050 ;
        RECT 176.100 383.400 199.050 384.450 ;
        RECT 176.100 382.950 178.200 383.400 ;
        RECT 196.950 382.950 199.050 383.400 ;
        RECT 160.950 381.450 163.050 382.050 ;
        RECT 169.950 381.450 172.050 382.050 ;
        RECT 160.950 380.400 172.050 381.450 ;
        RECT 160.950 379.950 163.050 380.400 ;
        RECT 169.950 379.950 172.050 380.400 ;
        RECT 178.950 381.450 181.050 382.050 ;
        RECT 193.950 381.450 196.050 382.050 ;
        RECT 178.950 380.400 196.050 381.450 ;
        RECT 178.950 379.950 181.050 380.400 ;
        RECT 193.950 379.950 196.050 380.400 ;
        RECT 211.950 379.950 217.050 382.050 ;
        RECT 223.950 379.950 229.050 382.050 ;
        RECT 241.950 379.950 244.050 385.050 ;
        RECT 259.950 384.450 264.900 385.050 ;
        RECT 248.400 384.000 264.900 384.450 ;
        RECT 265.950 384.000 268.200 385.050 ;
        RECT 247.950 383.400 264.900 384.000 ;
        RECT 247.950 379.950 250.050 383.400 ;
        RECT 259.950 382.950 264.900 383.400 ;
        RECT 266.100 382.950 268.200 384.000 ;
        RECT 271.950 382.950 277.050 385.050 ;
        RECT 308.400 382.050 309.450 386.400 ;
        RECT 322.950 386.400 331.050 387.000 ;
        RECT 322.950 385.050 325.050 386.400 ;
        RECT 328.950 385.950 331.050 386.400 ;
        RECT 340.950 387.450 343.050 388.050 ;
        RECT 346.950 387.450 349.050 388.050 ;
        RECT 340.950 386.400 349.050 387.450 ;
        RECT 340.950 385.950 343.050 386.400 ;
        RECT 346.950 385.950 349.050 386.400 ;
        RECT 313.950 382.950 319.050 385.050 ;
        RECT 322.800 384.000 325.050 385.050 ;
        RECT 326.100 384.450 328.200 385.050 ;
        RECT 337.950 384.450 340.050 385.050 ;
        RECT 326.100 384.000 340.050 384.450 ;
        RECT 322.800 382.950 324.900 384.000 ;
        RECT 325.950 383.400 340.050 384.000 ;
        RECT 325.950 382.950 328.200 383.400 ;
        RECT 337.950 382.950 340.050 383.400 ;
        RECT 349.950 384.450 355.050 385.050 ;
        RECT 361.950 384.450 364.050 385.050 ;
        RECT 349.950 383.400 364.050 384.450 ;
        RECT 349.950 382.950 355.050 383.400 ;
        RECT 361.950 382.950 364.050 383.400 ;
        RECT 325.950 382.050 328.050 382.950 ;
        RECT 259.950 379.950 265.050 382.050 ;
        RECT 268.950 379.950 274.050 382.050 ;
        RECT 298.950 379.950 304.050 382.050 ;
        RECT 307.950 379.950 310.050 382.050 ;
        RECT 319.950 379.950 324.900 382.050 ;
        RECT 325.950 381.000 328.200 382.050 ;
        RECT 326.100 379.950 328.200 381.000 ;
        RECT 343.950 379.950 349.050 382.050 ;
        RECT 367.950 379.950 370.050 385.050 ;
        RECT 376.950 382.950 379.050 388.050 ;
        RECT 385.950 382.950 388.050 388.050 ;
        RECT 412.950 387.450 415.050 388.050 ;
        RECT 407.400 387.000 450.450 387.450 ;
        RECT 406.950 386.400 450.450 387.000 ;
        RECT 406.950 382.950 409.050 386.400 ;
        RECT 412.950 385.950 415.050 386.400 ;
        RECT 449.400 385.050 450.450 386.400 ;
        RECT 382.950 381.450 385.050 382.050 ;
        RECT 388.950 381.450 391.050 382.050 ;
        RECT 382.950 380.400 391.050 381.450 ;
        RECT 382.950 379.950 385.050 380.400 ;
        RECT 388.950 379.950 391.050 380.400 ;
        RECT 421.950 381.450 424.050 382.050 ;
        RECT 430.950 381.450 433.050 385.050 ;
        RECT 436.800 384.000 438.900 385.050 ;
        RECT 436.800 382.950 439.050 384.000 ;
        RECT 442.950 382.950 448.050 385.050 ;
        RECT 449.400 383.400 454.050 385.050 ;
        RECT 450.000 382.950 454.050 383.400 ;
        RECT 436.950 382.050 439.050 382.950 ;
        RECT 421.950 381.000 433.050 381.450 ;
        RECT 433.800 381.000 435.900 382.050 ;
        RECT 436.800 381.000 439.050 382.050 ;
        RECT 440.100 381.450 442.200 382.050 ;
        RECT 448.950 381.450 451.050 382.050 ;
        RECT 421.950 380.400 432.450 381.000 ;
        RECT 421.950 379.950 424.050 380.400 ;
        RECT 433.800 379.950 436.050 381.000 ;
        RECT 436.800 379.950 438.900 381.000 ;
        RECT 440.100 380.400 451.050 381.450 ;
        RECT 440.100 379.950 442.200 380.400 ;
        RECT 448.950 379.950 451.050 380.400 ;
        RECT 118.950 378.450 121.050 379.050 ;
        RECT 124.950 378.450 127.050 379.050 ;
        RECT 118.950 377.400 127.050 378.450 ;
        RECT 118.950 376.950 121.050 377.400 ;
        RECT 124.950 376.950 127.050 377.400 ;
        RECT 130.950 376.950 136.050 379.050 ;
        RECT 100.950 375.450 103.050 376.050 ;
        RECT 136.950 375.450 139.050 376.050 ;
        RECT 100.950 374.400 139.050 375.450 ;
        RECT 139.950 375.450 142.050 379.050 ;
        RECT 151.950 378.450 154.050 379.050 ;
        RECT 157.950 378.450 160.050 379.050 ;
        RECT 151.950 377.400 160.050 378.450 ;
        RECT 151.950 376.950 154.050 377.400 ;
        RECT 157.950 376.950 160.050 377.400 ;
        RECT 187.950 376.950 193.050 379.050 ;
        RECT 154.950 375.450 157.050 376.050 ;
        RECT 178.950 375.450 181.050 376.050 ;
        RECT 139.950 375.000 181.050 375.450 ;
        RECT 140.400 374.400 181.050 375.000 ;
        RECT 100.950 373.950 103.050 374.400 ;
        RECT 136.950 373.950 139.050 374.400 ;
        RECT 154.950 373.950 157.050 374.400 ;
        RECT 178.950 373.950 181.050 374.400 ;
        RECT 196.950 373.950 199.050 379.050 ;
        RECT 232.950 376.950 238.050 379.050 ;
        RECT 244.950 378.450 247.050 379.050 ;
        RECT 260.400 378.450 261.450 379.950 ;
        RECT 244.950 377.400 261.450 378.450 ;
        RECT 265.950 378.450 268.050 379.050 ;
        RECT 280.950 378.450 283.050 379.050 ;
        RECT 265.950 377.400 283.050 378.450 ;
        RECT 244.950 376.950 247.050 377.400 ;
        RECT 265.950 376.950 268.050 377.400 ;
        RECT 280.950 376.950 283.050 377.400 ;
        RECT 286.950 378.450 289.050 379.050 ;
        RECT 295.950 378.450 298.050 379.050 ;
        RECT 286.950 377.400 298.050 378.450 ;
        RECT 286.950 376.950 289.050 377.400 ;
        RECT 295.950 376.950 298.050 377.400 ;
        RECT 304.950 376.950 310.050 379.050 ;
        RECT 400.950 378.450 403.050 379.050 ;
        RECT 430.950 378.450 433.050 379.050 ;
        RECT 433.950 378.450 436.050 379.950 ;
        RECT 400.950 378.000 436.050 378.450 ;
        RECT 400.950 377.400 435.300 378.000 ;
        RECT 455.850 377.400 457.050 389.400 ;
        RECT 460.950 382.950 466.050 385.050 ;
        RECT 469.950 379.950 472.050 385.050 ;
        RECT 400.950 376.950 403.050 377.400 ;
        RECT 430.950 376.950 433.050 377.400 ;
        RECT 229.950 375.450 232.050 376.050 ;
        RECT 283.950 375.450 286.050 376.050 ;
        RECT 229.950 374.400 286.050 375.450 ;
        RECT 229.950 373.950 232.050 374.400 ;
        RECT 283.950 373.950 286.050 374.400 ;
        RECT 292.950 375.450 295.050 376.050 ;
        RECT 313.950 375.450 316.050 376.050 ;
        RECT 292.950 374.400 316.050 375.450 ;
        RECT 292.950 373.950 295.050 374.400 ;
        RECT 313.950 373.950 316.050 374.400 ;
        RECT 322.950 375.450 325.050 376.050 ;
        RECT 343.950 375.450 346.050 376.050 ;
        RECT 322.950 374.400 346.050 375.450 ;
        RECT 454.950 375.300 457.050 377.400 ;
        RECT 322.950 373.950 325.050 374.400 ;
        RECT 343.950 373.950 346.050 374.400 ;
        RECT 73.950 372.450 76.050 373.050 ;
        RECT 112.950 372.450 115.050 373.050 ;
        RECT 73.950 371.400 115.050 372.450 ;
        RECT 73.950 370.950 76.050 371.400 ;
        RECT 112.950 370.950 115.050 371.400 ;
        RECT 133.950 372.450 136.050 373.050 ;
        RECT 148.950 372.450 151.050 373.050 ;
        RECT 133.950 371.400 151.050 372.450 ;
        RECT 133.950 370.950 136.050 371.400 ;
        RECT 148.950 370.950 151.050 371.400 ;
        RECT 367.950 372.450 370.050 373.050 ;
        RECT 421.950 372.450 424.050 373.200 ;
        RECT 367.950 371.400 424.050 372.450 ;
        RECT 455.850 371.700 457.050 375.300 ;
        RECT 476.100 372.600 477.300 389.400 ;
        RECT 502.950 388.950 505.050 389.400 ;
        RECT 517.950 388.950 520.050 389.400 ;
        RECT 526.950 390.450 529.050 391.050 ;
        RECT 544.950 390.450 547.050 390.900 ;
        RECT 526.950 389.400 547.050 390.450 ;
        RECT 526.950 388.950 529.050 389.400 ;
        RECT 544.950 388.800 547.050 389.400 ;
        RECT 625.950 390.450 628.050 391.050 ;
        RECT 685.950 390.450 688.050 391.050 ;
        RECT 802.950 390.450 805.050 391.050 ;
        RECT 817.950 390.450 820.050 391.050 ;
        RECT 625.950 389.400 688.050 390.450 ;
        RECT 740.400 390.000 805.050 390.450 ;
        RECT 625.950 388.950 628.050 389.400 ;
        RECT 685.950 388.950 688.050 389.400 ;
        RECT 739.950 389.400 805.050 390.000 ;
        RECT 529.950 387.450 532.050 388.050 ;
        RECT 509.400 386.400 532.050 387.450 ;
        RECT 493.800 384.000 495.900 385.050 ;
        RECT 497.100 384.450 499.200 385.050 ;
        RECT 509.400 384.450 510.450 386.400 ;
        RECT 529.950 385.950 532.050 386.400 ;
        RECT 493.800 382.950 496.050 384.000 ;
        RECT 497.100 383.400 510.450 384.450 ;
        RECT 497.100 382.950 499.200 383.400 ;
        RECT 511.950 382.950 517.050 385.050 ;
        RECT 538.950 382.950 541.050 388.050 ;
        RECT 544.950 382.950 547.050 388.050 ;
        RECT 610.950 387.450 613.050 388.050 ;
        RECT 661.950 387.450 664.050 388.050 ;
        RECT 610.950 387.000 618.300 387.450 ;
        RECT 644.400 387.000 664.050 387.450 ;
        RECT 610.950 386.400 619.050 387.000 ;
        RECT 610.950 385.950 613.050 386.400 ;
        RECT 616.950 385.050 619.050 386.400 ;
        RECT 643.950 386.400 664.050 387.000 ;
        RECT 550.950 384.450 553.050 385.050 ;
        RECT 559.950 384.450 562.050 385.050 ;
        RECT 550.950 383.400 562.050 384.450 ;
        RECT 550.950 382.950 553.050 383.400 ;
        RECT 559.950 382.950 562.050 383.400 ;
        RECT 574.950 382.950 580.050 385.050 ;
        RECT 583.950 382.950 589.050 385.050 ;
        RECT 607.950 384.450 610.050 385.050 ;
        RECT 613.800 384.450 615.900 385.050 ;
        RECT 593.400 383.400 615.900 384.450 ;
        RECT 493.950 379.950 496.050 382.950 ;
        RECT 593.400 382.050 594.450 383.400 ;
        RECT 607.950 382.950 610.050 383.400 ;
        RECT 613.800 382.950 615.900 383.400 ;
        RECT 616.800 384.000 619.050 385.050 ;
        RECT 619.800 384.000 621.900 385.050 ;
        RECT 623.100 384.450 625.200 385.050 ;
        RECT 631.800 384.450 633.900 385.050 ;
        RECT 616.800 382.950 618.900 384.000 ;
        RECT 619.800 382.950 622.050 384.000 ;
        RECT 623.100 383.400 633.900 384.450 ;
        RECT 623.100 382.950 625.200 383.400 ;
        RECT 631.800 382.950 633.900 383.400 ;
        RECT 635.100 382.950 640.050 385.050 ;
        RECT 643.950 382.950 646.050 386.400 ;
        RECT 661.950 385.950 664.050 386.400 ;
        RECT 667.950 387.450 670.050 388.200 ;
        RECT 667.950 386.400 678.450 387.450 ;
        RECT 667.950 386.100 670.050 386.400 ;
        RECT 677.400 385.050 678.450 386.400 ;
        RECT 718.950 385.950 724.050 388.050 ;
        RECT 739.950 385.950 742.050 389.400 ;
        RECT 802.950 388.950 805.050 389.400 ;
        RECT 812.400 389.400 820.050 390.450 ;
        RECT 799.950 387.450 802.050 388.200 ;
        RECT 812.400 387.450 813.450 389.400 ;
        RECT 817.950 388.950 820.050 389.400 ;
        RECT 826.950 390.450 829.050 391.050 ;
        RECT 832.950 390.450 835.050 391.200 ;
        RECT 826.950 389.400 835.050 390.450 ;
        RECT 826.950 388.950 829.050 389.400 ;
        RECT 832.950 389.100 835.050 389.400 ;
        RECT 844.950 390.450 847.050 391.050 ;
        RECT 850.950 390.450 853.050 391.050 ;
        RECT 844.950 389.400 853.050 390.450 ;
        RECT 844.950 388.950 847.050 389.400 ;
        RECT 850.950 388.950 853.050 389.400 ;
        RECT 799.950 386.400 813.450 387.450 ;
        RECT 799.950 386.100 802.050 386.400 ;
        RECT 806.400 385.050 807.450 386.400 ;
        RECT 649.950 384.450 652.050 385.050 ;
        RECT 658.950 384.450 661.050 385.050 ;
        RECT 649.950 383.400 661.050 384.450 ;
        RECT 649.950 382.950 652.050 383.400 ;
        RECT 658.950 382.950 661.050 383.400 ;
        RECT 667.950 384.450 670.050 384.900 ;
        RECT 667.950 384.000 675.450 384.450 ;
        RECT 667.950 383.400 676.050 384.000 ;
        RECT 677.400 383.400 682.050 385.050 ;
        RECT 487.950 378.450 490.050 379.050 ;
        RECT 499.950 378.450 502.050 382.050 ;
        RECT 505.950 381.450 508.050 382.050 ;
        RECT 511.800 381.450 513.900 382.050 ;
        RECT 505.950 380.400 513.900 381.450 ;
        RECT 505.950 379.950 508.050 380.400 ;
        RECT 511.800 379.950 513.900 380.400 ;
        RECT 515.100 379.950 520.050 382.050 ;
        RECT 529.950 381.450 532.050 382.050 ;
        RECT 535.950 381.450 538.050 382.050 ;
        RECT 529.950 380.400 538.050 381.450 ;
        RECT 529.950 379.950 532.050 380.400 ;
        RECT 535.950 379.950 538.050 380.400 ;
        RECT 487.950 378.000 502.050 378.450 ;
        RECT 502.950 378.450 505.050 379.050 ;
        RECT 517.800 378.450 519.900 379.050 ;
        RECT 487.950 377.400 501.450 378.000 ;
        RECT 502.950 377.400 519.900 378.450 ;
        RECT 487.950 376.950 490.050 377.400 ;
        RECT 502.950 376.950 505.050 377.400 ;
        RECT 517.800 376.950 519.900 377.400 ;
        RECT 521.100 378.450 523.200 379.050 ;
        RECT 532.950 378.450 535.050 379.050 ;
        RECT 521.100 377.400 535.050 378.450 ;
        RECT 541.950 378.450 544.050 382.050 ;
        RECT 547.950 381.450 550.050 382.050 ;
        RECT 556.950 381.450 559.050 382.050 ;
        RECT 547.950 380.400 559.050 381.450 ;
        RECT 547.950 379.950 550.050 380.400 ;
        RECT 556.950 379.950 559.050 380.400 ;
        RECT 580.950 381.450 583.050 382.050 ;
        RECT 580.950 380.400 588.450 381.450 ;
        RECT 580.950 379.950 583.050 380.400 ;
        RECT 550.950 378.450 553.050 379.050 ;
        RECT 541.950 378.000 553.050 378.450 ;
        RECT 542.400 377.400 553.050 378.000 ;
        RECT 587.400 378.450 588.450 380.400 ;
        RECT 589.950 380.400 594.450 382.050 ;
        RECT 589.950 379.950 594.000 380.400 ;
        RECT 598.950 379.950 604.050 382.050 ;
        RECT 619.950 379.950 622.050 382.950 ;
        RECT 667.950 382.800 670.050 383.400 ;
        RECT 625.950 379.950 631.050 382.050 ;
        RECT 640.950 379.950 645.900 382.050 ;
        RECT 647.100 381.000 649.200 382.050 ;
        RECT 646.950 379.950 649.200 381.000 ;
        RECT 661.950 381.450 664.050 382.050 ;
        RECT 667.950 381.450 670.050 382.050 ;
        RECT 661.950 380.400 670.050 381.450 ;
        RECT 661.950 379.950 664.050 380.400 ;
        RECT 667.950 379.950 670.050 380.400 ;
        RECT 673.950 379.950 676.050 383.400 ;
        RECT 678.000 382.950 682.050 383.400 ;
        RECT 703.950 384.450 706.050 385.050 ;
        RECT 709.950 384.450 712.050 385.050 ;
        RECT 703.950 383.400 712.050 384.450 ;
        RECT 703.950 382.950 706.050 383.400 ;
        RECT 709.950 382.950 712.050 383.400 ;
        RECT 760.950 384.450 763.050 385.050 ;
        RECT 766.950 384.450 769.050 385.050 ;
        RECT 760.950 383.400 769.050 384.450 ;
        RECT 760.950 382.950 763.050 383.400 ;
        RECT 766.950 382.950 769.050 383.400 ;
        RECT 781.950 384.450 784.050 385.050 ;
        RECT 793.950 384.450 796.050 385.050 ;
        RECT 781.950 383.400 796.050 384.450 ;
        RECT 781.950 382.950 784.050 383.400 ;
        RECT 793.950 382.950 796.050 383.400 ;
        RECT 799.950 382.950 805.050 385.050 ;
        RECT 806.400 383.400 811.050 385.050 ;
        RECT 807.000 382.950 811.050 383.400 ;
        RECT 814.950 382.950 817.050 388.050 ;
        RECT 832.950 387.450 835.050 387.900 ;
        RECT 853.950 387.450 856.050 388.050 ;
        RECT 832.950 386.400 856.050 387.450 ;
        RECT 832.950 385.800 835.050 386.400 ;
        RECT 853.950 385.950 856.050 386.400 ;
        RECT 820.950 384.450 825.000 385.050 ;
        RECT 826.950 384.450 829.050 385.050 ;
        RECT 847.950 384.450 850.050 385.050 ;
        RECT 820.950 382.950 825.450 384.450 ;
        RECT 826.950 383.400 850.050 384.450 ;
        RECT 826.950 382.950 829.050 383.400 ;
        RECT 847.950 382.950 850.050 383.400 ;
        RECT 685.950 381.450 688.050 382.050 ;
        RECT 706.950 381.450 709.050 382.050 ;
        RECT 685.950 380.400 709.050 381.450 ;
        RECT 685.950 379.950 688.050 380.400 ;
        RECT 706.950 379.950 709.050 380.400 ;
        RECT 715.950 379.950 721.050 382.050 ;
        RECT 730.950 381.450 733.050 382.050 ;
        RECT 736.950 381.450 739.050 382.050 ;
        RECT 730.950 380.400 739.050 381.450 ;
        RECT 730.950 379.950 733.050 380.400 ;
        RECT 736.950 379.950 739.050 380.400 ;
        RECT 772.950 381.450 775.050 382.050 ;
        RECT 790.950 381.450 793.050 382.050 ;
        RECT 772.950 380.400 793.050 381.450 ;
        RECT 772.950 379.950 775.050 380.400 ;
        RECT 790.950 379.950 793.050 380.400 ;
        RECT 646.950 379.050 649.050 379.950 ;
        RECT 598.950 378.450 601.050 379.050 ;
        RECT 587.400 377.400 601.050 378.450 ;
        RECT 521.100 376.950 523.200 377.400 ;
        RECT 532.950 376.950 535.050 377.400 ;
        RECT 550.950 376.950 553.050 377.400 ;
        RECT 598.950 376.950 601.050 377.400 ;
        RECT 604.950 378.450 607.050 379.050 ;
        RECT 610.950 378.450 613.050 379.050 ;
        RECT 604.950 377.400 613.050 378.450 ;
        RECT 646.950 378.000 649.200 379.050 ;
        RECT 670.950 378.450 673.050 379.050 ;
        RECT 604.950 376.950 607.050 377.400 ;
        RECT 610.950 376.950 613.050 377.400 ;
        RECT 647.100 376.950 649.200 378.000 ;
        RECT 659.400 377.400 673.050 378.450 ;
        RECT 484.950 375.450 487.050 376.050 ;
        RECT 514.950 375.450 517.050 376.050 ;
        RECT 553.950 375.450 556.050 376.050 ;
        RECT 484.950 374.400 556.050 375.450 ;
        RECT 484.950 373.950 487.050 374.400 ;
        RECT 514.950 373.950 517.050 374.400 ;
        RECT 553.950 373.950 556.050 374.400 ;
        RECT 640.950 375.450 643.050 376.050 ;
        RECT 659.400 375.450 660.450 377.400 ;
        RECT 670.950 376.950 673.050 377.400 ;
        RECT 691.950 378.450 694.050 379.050 ;
        RECT 700.950 378.450 706.050 379.050 ;
        RECT 691.950 377.400 706.050 378.450 ;
        RECT 691.950 376.950 694.050 377.400 ;
        RECT 700.950 376.950 706.050 377.400 ;
        RECT 773.100 376.950 778.050 379.050 ;
        RECT 796.950 378.450 799.050 382.050 ;
        RECT 808.950 378.450 811.050 379.050 ;
        RECT 796.950 378.000 811.050 378.450 ;
        RECT 811.950 378.450 814.050 382.050 ;
        RECT 817.950 379.950 823.050 382.050 ;
        RECT 824.400 381.450 825.450 382.950 ;
        RECT 835.950 381.450 838.050 382.050 ;
        RECT 824.400 380.400 838.050 381.450 ;
        RECT 835.950 379.950 838.050 380.400 ;
        RECT 826.950 378.450 829.050 379.050 ;
        RECT 811.950 378.000 829.050 378.450 ;
        RECT 797.400 377.400 811.050 378.000 ;
        RECT 812.400 377.400 829.050 378.000 ;
        RECT 808.950 376.950 811.050 377.400 ;
        RECT 826.950 376.950 829.050 377.400 ;
        RECT 640.950 374.400 660.450 375.450 ;
        RECT 661.950 375.450 664.050 376.050 ;
        RECT 670.950 375.450 673.050 376.050 ;
        RECT 682.950 375.450 685.050 376.050 ;
        RECT 661.950 374.400 685.050 375.450 ;
        RECT 640.950 373.950 643.050 374.400 ;
        RECT 661.950 373.950 664.050 374.400 ;
        RECT 670.950 373.950 673.050 374.400 ;
        RECT 682.950 373.950 685.050 374.400 ;
        RECT 706.950 375.450 709.050 376.050 ;
        RECT 712.950 375.450 715.050 376.050 ;
        RECT 706.950 374.400 715.050 375.450 ;
        RECT 706.950 373.950 709.050 374.400 ;
        RECT 712.950 373.950 715.050 374.400 ;
        RECT 733.950 375.450 736.050 376.050 ;
        RECT 745.950 375.450 748.050 376.050 ;
        RECT 733.950 374.400 748.050 375.450 ;
        RECT 832.950 375.450 835.050 379.050 ;
        RECT 838.950 378.450 841.050 379.050 ;
        RECT 844.950 378.450 847.050 379.050 ;
        RECT 850.950 378.450 853.050 379.050 ;
        RECT 838.950 377.400 853.050 378.450 ;
        RECT 838.950 376.950 841.050 377.400 ;
        RECT 844.950 376.950 847.050 377.400 ;
        RECT 850.950 376.950 853.050 377.400 ;
        RECT 841.950 375.450 844.050 376.050 ;
        RECT 853.950 375.450 856.050 376.050 ;
        RECT 832.950 375.000 856.050 375.450 ;
        RECT 833.400 374.400 856.050 375.000 ;
        RECT 733.950 373.950 736.050 374.400 ;
        RECT 745.950 373.950 748.050 374.400 ;
        RECT 841.950 373.950 844.050 374.400 ;
        RECT 853.950 373.950 856.050 374.400 ;
        RECT 367.950 370.950 370.050 371.400 ;
        RECT 421.950 371.100 424.050 371.400 ;
        RECT 187.950 369.450 190.050 370.050 ;
        RECT 214.950 369.450 217.050 370.050 ;
        RECT 187.950 368.400 217.050 369.450 ;
        RECT 187.950 367.950 190.050 368.400 ;
        RECT 214.950 367.950 217.050 368.400 ;
        RECT 259.950 369.450 262.050 370.050 ;
        RECT 277.950 369.450 280.050 370.050 ;
        RECT 259.950 368.400 280.050 369.450 ;
        RECT 259.950 367.950 262.050 368.400 ;
        RECT 277.950 367.950 280.050 368.400 ;
        RECT 304.950 369.450 307.050 370.050 ;
        RECT 328.950 369.450 331.050 370.050 ;
        RECT 423.000 369.900 427.050 370.050 ;
        RECT 304.950 368.400 331.050 369.450 ;
        RECT 304.950 367.950 307.050 368.400 ;
        RECT 328.950 367.950 331.050 368.400 ;
        RECT 421.950 367.950 427.050 369.900 ;
        RECT 421.950 367.800 424.050 367.950 ;
        RECT 13.950 366.450 16.050 367.050 ;
        RECT 25.950 366.450 28.050 367.050 ;
        RECT 13.950 365.400 28.050 366.450 ;
        RECT 13.950 364.950 16.050 365.400 ;
        RECT 25.950 364.950 28.050 365.400 ;
        RECT 112.950 364.950 118.050 367.050 ;
        RECT 130.950 366.450 133.050 367.050 ;
        RECT 145.950 366.450 148.050 367.050 ;
        RECT 130.950 365.400 148.050 366.450 ;
        RECT 130.950 364.950 133.050 365.400 ;
        RECT 145.950 364.950 148.050 365.400 ;
        RECT 178.950 364.950 184.050 367.050 ;
        RECT 211.950 366.450 214.050 367.050 ;
        RECT 292.950 366.450 295.050 367.050 ;
        RECT 211.950 365.400 295.050 366.450 ;
        RECT 211.950 364.950 214.050 365.400 ;
        RECT 292.950 364.950 295.050 365.400 ;
        RECT 370.950 366.450 373.050 367.050 ;
        RECT 409.950 366.450 412.050 367.050 ;
        RECT 370.950 365.400 412.050 366.450 ;
        RECT 436.950 366.450 439.050 370.050 ;
        RECT 454.950 369.600 457.050 371.700 ;
        RECT 475.950 370.500 478.050 372.600 ;
        RECT 487.950 372.450 490.050 373.050 ;
        RECT 511.950 372.450 514.050 373.050 ;
        RECT 487.950 371.400 514.050 372.450 ;
        RECT 487.950 370.950 490.050 371.400 ;
        RECT 511.950 370.950 514.050 371.400 ;
        RECT 613.950 372.450 616.050 373.050 ;
        RECT 622.950 372.450 625.050 373.050 ;
        RECT 613.950 371.400 625.050 372.450 ;
        RECT 613.950 370.950 616.050 371.400 ;
        RECT 622.950 370.950 625.050 371.400 ;
        RECT 673.950 372.450 676.050 373.050 ;
        RECT 694.950 372.450 697.050 373.050 ;
        RECT 673.950 371.400 697.050 372.450 ;
        RECT 673.950 370.950 676.050 371.400 ;
        RECT 694.950 370.950 697.050 371.400 ;
        RECT 709.950 372.450 712.050 373.050 ;
        RECT 844.950 372.450 847.050 373.050 ;
        RECT 709.950 371.400 847.050 372.450 ;
        RECT 709.950 370.950 712.050 371.400 ;
        RECT 844.950 370.950 847.050 371.400 ;
        RECT 496.950 369.450 499.050 370.050 ;
        RECT 505.950 369.450 508.050 370.050 ;
        RECT 496.950 368.400 508.050 369.450 ;
        RECT 496.950 367.950 499.050 368.400 ;
        RECT 505.950 367.950 508.050 368.400 ;
        RECT 571.950 369.450 574.050 370.050 ;
        RECT 601.950 369.450 604.050 370.050 ;
        RECT 730.950 369.450 733.050 370.050 ;
        RECT 772.950 369.450 775.050 370.050 ;
        RECT 571.950 368.400 733.050 369.450 ;
        RECT 571.950 367.950 574.050 368.400 ;
        RECT 601.950 367.950 604.050 368.400 ;
        RECT 730.950 367.950 733.050 368.400 ;
        RECT 761.400 368.400 775.050 369.450 ;
        RECT 469.950 366.450 472.050 367.050 ;
        RECT 436.950 366.000 472.050 366.450 ;
        RECT 437.400 365.400 472.050 366.000 ;
        RECT 370.950 364.950 373.050 365.400 ;
        RECT 409.950 364.950 412.050 365.400 ;
        RECT 469.950 364.950 472.050 365.400 ;
        RECT 481.950 366.450 484.050 367.050 ;
        RECT 526.950 366.450 529.050 367.050 ;
        RECT 481.950 365.400 529.050 366.450 ;
        RECT 481.950 364.950 484.050 365.400 ;
        RECT 526.950 364.950 529.050 365.400 ;
        RECT 559.950 366.450 562.050 367.050 ;
        RECT 571.950 366.450 574.050 367.050 ;
        RECT 559.950 365.400 574.050 366.450 ;
        RECT 559.950 364.950 562.050 365.400 ;
        RECT 571.950 364.950 574.050 365.400 ;
        RECT 625.950 366.450 628.050 367.050 ;
        RECT 631.950 366.450 634.050 367.050 ;
        RECT 625.950 365.400 634.050 366.450 ;
        RECT 625.950 364.950 628.050 365.400 ;
        RECT 631.950 364.950 634.050 365.400 ;
        RECT 646.950 366.450 649.050 367.050 ;
        RECT 676.950 366.450 679.050 367.050 ;
        RECT 646.950 365.400 679.050 366.450 ;
        RECT 646.950 364.950 649.050 365.400 ;
        RECT 676.950 364.950 679.050 365.400 ;
        RECT 694.950 366.450 697.050 367.050 ;
        RECT 700.950 366.450 703.050 367.050 ;
        RECT 694.950 365.400 703.050 366.450 ;
        RECT 694.950 364.950 697.050 365.400 ;
        RECT 700.950 364.950 703.050 365.400 ;
        RECT 730.950 366.450 733.050 367.050 ;
        RECT 761.400 366.450 762.450 368.400 ;
        RECT 772.950 367.950 775.050 368.400 ;
        RECT 796.950 369.450 799.050 370.050 ;
        RECT 820.950 369.450 823.050 370.050 ;
        RECT 796.950 368.400 823.050 369.450 ;
        RECT 796.950 367.950 799.050 368.400 ;
        RECT 820.950 367.950 823.050 368.400 ;
        RECT 826.950 367.950 832.050 370.050 ;
        RECT 853.950 367.950 859.050 370.050 ;
        RECT 799.950 366.450 802.050 367.050 ;
        RECT 730.950 365.400 762.450 366.450 ;
        RECT 788.400 365.400 802.050 366.450 ;
        RECT 730.950 364.950 733.050 365.400 ;
        RECT 73.950 363.450 76.050 364.050 ;
        RECT 124.950 363.450 127.050 364.050 ;
        RECT 145.950 363.450 148.050 364.050 ;
        RECT 73.950 362.400 148.050 363.450 ;
        RECT 73.950 361.950 76.050 362.400 ;
        RECT 124.950 361.950 127.050 362.400 ;
        RECT 145.950 361.950 148.050 362.400 ;
        RECT 373.950 363.450 376.050 364.050 ;
        RECT 508.950 363.450 511.050 364.050 ;
        RECT 373.950 362.400 511.050 363.450 ;
        RECT 373.950 361.950 376.050 362.400 ;
        RECT 508.950 361.950 511.050 362.400 ;
        RECT 637.950 363.450 640.050 364.050 ;
        RECT 706.950 363.450 709.050 364.050 ;
        RECT 637.950 362.400 709.050 363.450 ;
        RECT 637.950 361.950 640.050 362.400 ;
        RECT 706.950 361.950 709.050 362.400 ;
        RECT 715.950 363.450 718.050 364.050 ;
        RECT 788.400 363.450 789.450 365.400 ;
        RECT 799.950 364.950 802.050 365.400 ;
        RECT 715.950 362.400 789.450 363.450 ;
        RECT 715.950 361.950 718.050 362.400 ;
        RECT 37.950 360.450 40.050 361.050 ;
        RECT 67.950 360.450 70.050 361.050 ;
        RECT 37.950 359.400 70.050 360.450 ;
        RECT 37.950 358.950 40.050 359.400 ;
        RECT 67.950 358.950 70.050 359.400 ;
        RECT 97.950 360.450 100.050 361.050 ;
        RECT 136.950 360.450 139.050 361.050 ;
        RECT 97.950 359.400 139.050 360.450 ;
        RECT 97.950 358.950 100.050 359.400 ;
        RECT 136.950 358.950 139.050 359.400 ;
        RECT 238.950 360.450 241.050 361.050 ;
        RECT 250.950 360.450 253.050 361.200 ;
        RECT 238.950 359.400 253.050 360.450 ;
        RECT 238.950 358.950 241.050 359.400 ;
        RECT 250.950 359.100 253.050 359.400 ;
        RECT 79.950 357.450 82.050 358.050 ;
        RECT 103.950 357.450 106.050 358.050 ;
        RECT 172.950 357.450 175.050 358.050 ;
        RECT 250.950 357.450 253.050 357.900 ;
        RECT 79.950 356.400 135.450 357.450 ;
        RECT 79.950 355.950 82.050 356.400 ;
        RECT 103.950 355.950 106.050 356.400 ;
        RECT 134.400 355.050 135.450 356.400 ;
        RECT 172.950 356.400 253.050 357.450 ;
        RECT 172.950 355.950 175.050 356.400 ;
        RECT 250.950 355.800 253.050 356.400 ;
        RECT 262.950 357.450 265.050 358.050 ;
        RECT 271.950 357.450 274.050 358.050 ;
        RECT 262.950 356.400 274.050 357.450 ;
        RECT 283.950 357.450 286.050 361.050 ;
        RECT 430.950 360.450 433.050 361.050 ;
        RECT 436.950 360.450 439.050 361.050 ;
        RECT 430.950 359.400 439.050 360.450 ;
        RECT 430.950 358.950 433.050 359.400 ;
        RECT 436.950 358.950 439.050 359.400 ;
        RECT 463.950 360.450 466.050 361.050 ;
        RECT 556.800 360.450 558.900 361.050 ;
        RECT 463.950 359.400 558.900 360.450 ;
        RECT 463.950 358.950 466.050 359.400 ;
        RECT 556.800 358.950 558.900 359.400 ;
        RECT 560.100 360.450 562.200 361.050 ;
        RECT 586.950 360.450 589.050 361.050 ;
        RECT 560.100 359.400 589.050 360.450 ;
        RECT 560.100 358.950 562.200 359.400 ;
        RECT 586.950 358.950 589.050 359.400 ;
        RECT 640.950 360.450 643.050 361.050 ;
        RECT 679.950 360.450 682.050 361.050 ;
        RECT 640.950 359.400 682.050 360.450 ;
        RECT 640.950 358.950 643.050 359.400 ;
        RECT 679.950 358.950 682.050 359.400 ;
        RECT 703.950 360.450 706.050 361.050 ;
        RECT 757.950 360.450 760.050 361.050 ;
        RECT 781.950 360.450 784.050 361.050 ;
        RECT 703.950 359.400 760.050 360.450 ;
        RECT 703.950 358.950 706.050 359.400 ;
        RECT 757.950 358.950 760.050 359.400 ;
        RECT 764.400 359.400 784.050 360.450 ;
        RECT 400.950 357.450 403.050 358.050 ;
        RECT 283.950 357.000 403.050 357.450 ;
        RECT 284.400 356.400 403.050 357.000 ;
        RECT 262.950 355.950 265.050 356.400 ;
        RECT 271.950 355.950 274.050 356.400 ;
        RECT 400.950 355.950 403.050 356.400 ;
        RECT 496.950 357.450 499.050 358.050 ;
        RECT 547.950 357.450 550.050 358.050 ;
        RECT 496.950 356.400 550.050 357.450 ;
        RECT 496.950 355.950 499.050 356.400 ;
        RECT 547.950 355.950 550.050 356.400 ;
        RECT 571.950 357.450 574.050 358.050 ;
        RECT 577.950 357.450 580.050 358.050 ;
        RECT 571.950 356.400 580.050 357.450 ;
        RECT 571.950 355.950 574.050 356.400 ;
        RECT 577.950 355.950 580.050 356.400 ;
        RECT 598.950 357.450 601.050 358.200 ;
        RECT 607.950 357.450 610.050 358.050 ;
        RECT 598.950 356.400 610.050 357.450 ;
        RECT 598.950 356.100 601.050 356.400 ;
        RECT 607.950 355.950 610.050 356.400 ;
        RECT 643.950 357.450 646.050 358.050 ;
        RECT 655.950 357.450 658.050 358.050 ;
        RECT 643.950 356.400 658.050 357.450 ;
        RECT 643.950 355.950 646.050 356.400 ;
        RECT 655.950 355.950 658.050 356.400 ;
        RECT 691.950 357.450 694.050 358.050 ;
        RECT 764.400 357.450 765.450 359.400 ;
        RECT 781.950 358.950 784.050 359.400 ;
        RECT 823.950 360.450 826.050 361.050 ;
        RECT 856.950 360.450 859.050 361.050 ;
        RECT 823.950 359.400 859.050 360.450 ;
        RECT 823.950 358.950 826.050 359.400 ;
        RECT 856.950 358.950 859.050 359.400 ;
        RECT 691.950 356.400 765.450 357.450 ;
        RECT 772.950 357.450 775.050 358.050 ;
        RECT 796.950 357.450 799.050 358.050 ;
        RECT 772.950 356.400 799.050 357.450 ;
        RECT 691.950 355.950 694.050 356.400 ;
        RECT 772.950 355.950 775.050 356.400 ;
        RECT 796.950 355.950 799.050 356.400 ;
        RECT 805.950 357.450 808.050 358.050 ;
        RECT 817.950 357.450 820.050 358.050 ;
        RECT 805.950 356.400 820.050 357.450 ;
        RECT 805.950 355.950 808.050 356.400 ;
        RECT 817.950 355.950 820.050 356.400 ;
        RECT 844.950 357.450 847.050 358.050 ;
        RECT 850.950 357.450 853.050 358.050 ;
        RECT 844.950 356.400 853.050 357.450 ;
        RECT 844.950 355.950 847.050 356.400 ;
        RECT 850.950 355.950 853.050 356.400 ;
        RECT 64.950 354.450 67.050 355.050 ;
        RECT 82.950 354.450 85.050 355.050 ;
        RECT 118.950 354.450 121.050 355.050 ;
        RECT 64.950 353.400 121.050 354.450 ;
        RECT 64.950 352.950 67.050 353.400 ;
        RECT 82.950 352.950 85.050 353.400 ;
        RECT 118.950 352.950 121.050 353.400 ;
        RECT 133.950 354.450 136.050 355.050 ;
        RECT 208.950 354.450 211.050 355.050 ;
        RECT 376.950 354.450 379.050 355.050 ;
        RECT 133.950 353.400 211.050 354.450 ;
        RECT 133.950 352.950 136.050 353.400 ;
        RECT 208.950 352.950 211.050 353.400 ;
        RECT 353.400 353.400 379.050 354.450 ;
        RECT 353.400 352.200 354.450 353.400 ;
        RECT 376.950 352.950 379.050 353.400 ;
        RECT 382.950 354.450 385.050 355.050 ;
        RECT 388.950 354.450 391.050 355.050 ;
        RECT 382.950 353.400 391.050 354.450 ;
        RECT 382.950 352.950 385.050 353.400 ;
        RECT 388.950 352.950 391.050 353.400 ;
        RECT 430.950 354.450 433.050 355.050 ;
        RECT 475.950 354.450 478.050 355.050 ;
        RECT 430.950 353.400 478.050 354.450 ;
        RECT 430.950 352.950 433.050 353.400 ;
        RECT 475.950 352.950 478.050 353.400 ;
        RECT 550.950 354.450 553.050 355.050 ;
        RECT 565.950 354.450 568.050 355.050 ;
        RECT 550.950 353.400 568.050 354.450 ;
        RECT 550.950 352.950 553.050 353.400 ;
        RECT 565.950 352.950 568.050 353.400 ;
        RECT 583.950 354.450 586.050 355.050 ;
        RECT 598.950 354.450 601.050 354.900 ;
        RECT 613.950 354.450 616.050 355.050 ;
        RECT 583.950 353.400 616.050 354.450 ;
        RECT 583.950 352.950 586.050 353.400 ;
        RECT 598.950 352.800 601.050 353.400 ;
        RECT 613.950 352.950 616.050 353.400 ;
        RECT 661.950 354.450 664.050 355.050 ;
        RECT 691.950 354.450 694.050 355.050 ;
        RECT 661.950 353.400 694.050 354.450 ;
        RECT 661.950 352.950 664.050 353.400 ;
        RECT 691.950 352.950 694.050 353.400 ;
        RECT 724.950 354.450 727.050 355.050 ;
        RECT 739.950 354.450 742.050 355.050 ;
        RECT 856.950 354.450 859.050 355.050 ;
        RECT 724.950 353.400 742.050 354.450 ;
        RECT 724.950 352.950 727.050 353.400 ;
        RECT 739.950 352.950 742.050 353.400 ;
        RECT 815.400 353.400 859.050 354.450 ;
        RECT 76.950 351.450 79.050 352.050 ;
        RECT 85.950 351.450 88.050 352.050 ;
        RECT 127.950 351.450 130.050 352.050 ;
        RECT 76.950 350.400 130.050 351.450 ;
        RECT 76.950 349.950 79.050 350.400 ;
        RECT 85.950 349.950 88.050 350.400 ;
        RECT 127.950 349.950 130.050 350.400 ;
        RECT 184.950 351.450 187.050 352.050 ;
        RECT 247.950 351.450 250.050 352.050 ;
        RECT 184.950 350.400 250.050 351.450 ;
        RECT 184.950 349.950 187.050 350.400 ;
        RECT 247.950 349.950 250.050 350.400 ;
        RECT 298.950 351.450 301.050 352.050 ;
        RECT 319.950 351.450 322.050 352.050 ;
        RECT 298.950 350.400 322.050 351.450 ;
        RECT 298.950 349.950 301.050 350.400 ;
        RECT 319.950 349.950 322.050 350.400 ;
        RECT 325.950 351.450 328.050 352.050 ;
        RECT 352.950 351.450 355.050 352.200 ;
        RECT 325.950 350.400 355.050 351.450 ;
        RECT 325.950 349.950 328.050 350.400 ;
        RECT 352.950 350.100 355.050 350.400 ;
        RECT 436.950 351.450 439.050 352.050 ;
        RECT 457.950 351.450 460.050 352.050 ;
        RECT 496.950 351.450 499.050 352.050 ;
        RECT 436.950 350.400 499.050 351.450 ;
        RECT 436.950 349.950 439.050 350.400 ;
        RECT 457.950 349.950 460.050 350.400 ;
        RECT 496.950 349.950 499.050 350.400 ;
        RECT 514.950 351.450 517.050 352.050 ;
        RECT 595.950 351.450 598.050 352.050 ;
        RECT 622.950 351.450 625.050 352.050 ;
        RECT 514.950 350.400 625.050 351.450 ;
        RECT 514.950 349.950 517.050 350.400 ;
        RECT 595.950 349.950 598.050 350.400 ;
        RECT 622.950 349.950 625.050 350.400 ;
        RECT 631.950 351.450 634.050 352.050 ;
        RECT 652.950 351.450 655.050 352.050 ;
        RECT 631.950 350.400 655.050 351.450 ;
        RECT 631.950 349.950 634.050 350.400 ;
        RECT 652.950 349.950 655.050 350.400 ;
        RECT 664.950 351.450 667.050 352.050 ;
        RECT 682.950 351.450 685.050 352.050 ;
        RECT 700.950 351.450 703.050 352.050 ;
        RECT 664.950 350.400 703.050 351.450 ;
        RECT 664.950 349.950 667.050 350.400 ;
        RECT 682.950 349.950 685.050 350.400 ;
        RECT 700.950 349.950 703.050 350.400 ;
        RECT 706.950 351.450 709.050 352.050 ;
        RECT 778.950 351.450 781.050 352.050 ;
        RECT 802.950 351.450 805.050 352.050 ;
        RECT 815.400 351.450 816.450 353.400 ;
        RECT 856.950 352.950 859.050 353.400 ;
        RECT 706.950 350.400 756.450 351.450 ;
        RECT 706.950 349.950 709.050 350.400 ;
        RECT 755.400 349.050 756.450 350.400 ;
        RECT 778.950 350.400 816.450 351.450 ;
        RECT 817.950 351.450 820.050 352.050 ;
        RECT 832.800 351.450 834.900 352.050 ;
        RECT 817.950 350.400 834.900 351.450 ;
        RECT 778.950 349.950 781.050 350.400 ;
        RECT 802.950 349.950 805.050 350.400 ;
        RECT 817.950 349.950 820.050 350.400 ;
        RECT 832.800 349.950 834.900 350.400 ;
        RECT 836.100 351.450 838.200 352.050 ;
        RECT 850.950 351.450 853.050 352.050 ;
        RECT 836.100 350.400 853.050 351.450 ;
        RECT 836.100 349.950 838.200 350.400 ;
        RECT 850.950 349.950 853.050 350.400 ;
        RECT 22.950 348.450 25.050 349.050 ;
        RECT 91.950 348.450 94.050 349.050 ;
        RECT 115.800 348.450 117.900 349.050 ;
        RECT 22.950 347.400 60.600 348.450 ;
        RECT 22.950 346.950 25.050 347.400 ;
        RECT 14.100 346.050 16.200 346.200 ;
        RECT 7.950 343.950 12.900 346.050 ;
        RECT 14.100 344.100 19.050 346.050 ;
        RECT 15.000 343.950 19.050 344.100 ;
        RECT 28.950 343.050 31.050 343.200 ;
        RECT 13.950 337.950 16.050 343.050 ;
        RECT 19.950 340.950 25.050 343.050 ;
        RECT 28.950 341.100 34.050 343.050 ;
        RECT 30.000 340.950 34.050 341.100 ;
        RECT 37.950 342.450 40.050 343.050 ;
        RECT 46.950 342.450 49.050 343.200 ;
        RECT 59.550 343.050 60.600 347.400 ;
        RECT 91.950 348.000 117.900 348.450 ;
        RECT 119.100 348.450 123.000 349.050 ;
        RECT 144.000 348.450 148.050 349.050 ;
        RECT 119.100 348.000 123.450 348.450 ;
        RECT 91.950 347.400 118.050 348.000 ;
        RECT 91.950 346.950 94.050 347.400 ;
        RECT 115.800 346.950 118.050 347.400 ;
        RECT 119.100 346.950 124.050 348.000 ;
        RECT 73.950 345.450 76.050 346.200 ;
        RECT 79.950 345.450 82.050 346.050 ;
        RECT 106.950 345.450 111.000 346.050 ;
        RECT 73.950 344.400 82.050 345.450 ;
        RECT 83.400 345.000 111.450 345.450 ;
        RECT 73.950 344.100 76.050 344.400 ;
        RECT 79.950 343.950 82.050 344.400 ;
        RECT 82.950 344.400 111.450 345.000 ;
        RECT 52.800 342.450 54.900 343.050 ;
        RECT 37.950 341.400 54.900 342.450 ;
        RECT 37.950 340.950 40.050 341.400 ;
        RECT 46.950 341.100 49.050 341.400 ;
        RECT 52.800 340.950 54.900 341.400 ;
        RECT 55.800 342.000 57.900 343.050 ;
        RECT 55.800 340.950 58.050 342.000 ;
        RECT 59.100 340.950 61.200 343.050 ;
        RECT 75.000 342.900 79.050 343.050 ;
        RECT 73.950 340.950 79.050 342.900 ;
        RECT 82.950 340.950 85.050 344.400 ;
        RECT 106.950 343.950 111.450 344.400 ;
        RECT 115.950 343.950 118.050 346.950 ;
        RECT 121.950 343.950 124.050 346.950 ;
        RECT 143.400 346.950 148.050 348.450 ;
        RECT 154.950 348.450 157.050 349.050 ;
        RECT 175.950 348.450 178.050 349.050 ;
        RECT 184.950 348.450 187.050 349.050 ;
        RECT 154.950 347.400 178.050 348.450 ;
        RECT 154.950 346.950 157.050 347.400 ;
        RECT 175.950 346.950 178.050 347.400 ;
        RECT 179.400 347.400 187.050 348.450 ;
        RECT 137.100 345.000 139.200 346.050 ;
        RECT 136.950 343.950 139.200 345.000 ;
        RECT 98.100 343.050 100.200 343.200 ;
        RECT 110.400 343.050 111.450 343.950 ;
        RECT 136.950 343.050 139.050 343.950 ;
        RECT 143.400 343.050 144.450 346.950 ;
        RECT 148.950 345.450 151.050 346.050 ;
        RECT 154.950 345.450 157.050 346.050 ;
        RECT 148.950 344.400 157.050 345.450 ;
        RECT 148.950 343.950 151.050 344.400 ;
        RECT 154.950 343.950 157.050 344.400 ;
        RECT 163.950 345.450 166.050 346.050 ;
        RECT 179.400 345.450 180.450 347.400 ;
        RECT 163.950 344.400 180.450 345.450 ;
        RECT 163.950 343.950 166.050 344.400 ;
        RECT 184.950 343.950 187.050 347.400 ;
        RECT 196.950 348.450 199.050 349.050 ;
        RECT 226.950 348.450 229.050 349.050 ;
        RECT 196.950 347.400 229.050 348.450 ;
        RECT 196.950 343.950 199.050 347.400 ;
        RECT 226.950 346.950 229.050 347.400 ;
        RECT 232.950 348.450 235.050 349.050 ;
        RECT 265.950 348.450 268.050 349.050 ;
        RECT 352.950 348.450 355.050 348.900 ;
        RECT 232.950 347.400 268.050 348.450 ;
        RECT 232.950 346.950 235.050 347.400 ;
        RECT 265.950 346.950 268.050 347.400 ;
        RECT 275.400 347.400 285.450 348.450 ;
        RECT 202.950 343.950 208.050 346.050 ;
        RECT 223.950 345.450 226.050 346.050 ;
        RECT 241.950 345.450 244.050 346.050 ;
        RECT 275.400 345.450 276.450 347.400 ;
        RECT 223.950 344.400 276.450 345.450 ;
        RECT 91.950 340.950 96.900 343.050 ;
        RECT 98.100 341.100 102.900 343.050 ;
        RECT 104.100 342.000 106.200 343.050 ;
        RECT 99.000 340.950 102.900 341.100 ;
        RECT 103.950 340.950 106.200 342.000 ;
        RECT 110.400 341.400 115.050 343.050 ;
        RECT 111.000 340.950 115.050 341.400 ;
        RECT 55.950 340.050 58.050 340.950 ;
        RECT 73.950 340.800 76.050 340.950 ;
        RECT 103.950 340.050 106.050 340.950 ;
        RECT 28.950 339.450 31.050 339.900 ;
        RECT 34.950 339.450 37.050 340.050 ;
        RECT 28.950 338.400 37.050 339.450 ;
        RECT 28.950 337.800 31.050 338.400 ;
        RECT 34.950 337.950 37.050 338.400 ;
        RECT 40.950 339.450 43.050 340.050 ;
        RECT 48.000 339.900 52.050 340.050 ;
        RECT 46.950 339.450 52.050 339.900 ;
        RECT 40.950 338.400 52.050 339.450 ;
        RECT 40.950 337.950 43.050 338.400 ;
        RECT 46.950 337.950 52.050 338.400 ;
        RECT 55.800 339.000 58.050 340.050 ;
        RECT 55.800 337.950 57.900 339.000 ;
        RECT 97.950 337.950 102.900 340.050 ;
        RECT 103.950 339.000 106.200 340.050 ;
        RECT 118.950 339.450 121.050 343.050 ;
        RECT 133.800 342.000 135.900 343.050 ;
        RECT 136.950 342.000 139.200 343.050 ;
        RECT 133.800 340.950 136.050 342.000 ;
        RECT 137.100 340.950 139.200 342.000 ;
        RECT 142.950 340.950 145.050 343.050 ;
        RECT 154.950 342.450 157.050 343.050 ;
        RECT 160.950 342.450 163.050 343.050 ;
        RECT 154.950 341.400 163.050 342.450 ;
        RECT 154.950 340.950 157.050 341.400 ;
        RECT 160.950 340.950 163.050 341.400 ;
        RECT 166.950 340.950 172.050 343.050 ;
        RECT 175.950 342.450 178.050 343.050 ;
        RECT 181.950 342.450 184.050 343.050 ;
        RECT 175.950 341.400 184.050 342.450 ;
        RECT 175.950 340.950 178.050 341.400 ;
        RECT 181.950 340.950 184.050 341.400 ;
        RECT 127.950 339.450 130.050 340.050 ;
        RECT 118.950 339.000 130.050 339.450 ;
        RECT 104.100 337.950 106.200 339.000 ;
        RECT 119.400 338.400 130.050 339.000 ;
        RECT 127.950 337.950 130.050 338.400 ;
        RECT 133.950 337.950 136.050 340.950 ;
        RECT 138.000 339.450 142.050 340.050 ;
        RECT 137.400 337.950 142.050 339.450 ;
        RECT 187.950 337.950 190.050 343.050 ;
        RECT 199.950 340.950 205.050 343.050 ;
        RECT 214.950 340.950 220.050 343.050 ;
        RECT 223.950 340.950 226.050 344.400 ;
        RECT 241.950 343.950 244.050 344.400 ;
        RECT 46.950 337.800 49.050 337.950 ;
        RECT 124.950 336.450 127.050 337.050 ;
        RECT 137.400 336.450 138.450 337.950 ;
        RECT 124.950 335.400 138.450 336.450 ;
        RECT 157.950 336.450 160.050 337.050 ;
        RECT 172.950 336.450 175.050 337.050 ;
        RECT 157.950 335.400 175.050 336.450 ;
        RECT 124.950 334.950 127.050 335.400 ;
        RECT 157.950 334.950 160.050 335.400 ;
        RECT 172.950 334.950 175.050 335.400 ;
        RECT 202.950 336.450 205.050 337.050 ;
        RECT 220.950 336.450 223.050 340.050 ;
        RECT 226.950 339.450 229.050 340.050 ;
        RECT 232.950 339.450 238.050 340.050 ;
        RECT 226.950 338.400 238.050 339.450 ;
        RECT 226.950 337.950 229.050 338.400 ;
        RECT 232.950 337.950 238.050 338.400 ;
        RECT 241.950 337.950 244.050 343.050 ;
        RECT 253.950 340.950 259.050 343.050 ;
        RECT 262.950 340.950 265.050 344.400 ;
        RECT 284.400 343.050 285.450 347.400 ;
        RECT 296.400 347.400 355.050 348.450 ;
        RECT 296.400 346.050 297.450 347.400 ;
        RECT 352.950 346.800 355.050 347.400 ;
        RECT 358.950 348.450 361.050 349.050 ;
        RECT 364.950 348.450 367.050 349.050 ;
        RECT 358.950 347.400 367.050 348.450 ;
        RECT 358.950 346.950 361.050 347.400 ;
        RECT 364.950 346.950 367.050 347.400 ;
        RECT 376.950 348.450 379.050 349.050 ;
        RECT 409.950 348.450 412.050 349.050 ;
        RECT 439.950 348.450 442.050 349.050 ;
        RECT 376.950 348.000 390.450 348.450 ;
        RECT 376.950 347.400 391.050 348.000 ;
        RECT 376.950 346.950 379.050 347.400 ;
        RECT 328.950 346.050 331.050 346.200 ;
        RECT 388.950 346.050 391.050 347.400 ;
        RECT 409.950 347.400 442.050 348.450 ;
        RECT 409.950 346.950 412.050 347.400 ;
        RECT 439.950 346.950 442.050 347.400 ;
        RECT 547.950 348.450 550.050 349.050 ;
        RECT 559.950 348.450 562.050 349.050 ;
        RECT 547.950 347.400 562.050 348.450 ;
        RECT 547.950 346.950 550.050 347.400 ;
        RECT 559.950 346.950 562.050 347.400 ;
        RECT 583.800 348.000 585.900 349.050 ;
        RECT 587.100 348.450 589.200 349.050 ;
        RECT 610.950 348.450 613.050 349.050 ;
        RECT 616.950 348.450 619.050 349.050 ;
        RECT 583.800 346.950 586.050 348.000 ;
        RECT 587.100 347.400 619.050 348.450 ;
        RECT 587.100 346.950 589.200 347.400 ;
        RECT 610.950 346.950 613.050 347.400 ;
        RECT 616.950 346.950 619.050 347.400 ;
        RECT 628.950 348.450 631.050 349.050 ;
        RECT 634.950 348.450 637.050 349.050 ;
        RECT 628.950 347.400 637.050 348.450 ;
        RECT 628.950 346.950 631.050 347.400 ;
        RECT 634.950 346.950 637.050 347.400 ;
        RECT 295.800 345.450 297.900 346.050 ;
        RECT 287.550 344.400 297.900 345.450 ;
        RECT 299.100 345.000 301.200 346.050 ;
        RECT 271.950 342.450 274.050 343.050 ;
        RECT 277.950 342.450 280.050 343.050 ;
        RECT 271.950 341.400 280.050 342.450 ;
        RECT 271.950 340.950 274.050 341.400 ;
        RECT 277.950 340.050 280.050 341.400 ;
        RECT 283.950 340.950 286.050 343.050 ;
        RECT 287.550 340.050 288.600 344.400 ;
        RECT 295.800 343.950 297.900 344.400 ;
        RECT 298.950 343.950 301.200 345.000 ;
        RECT 307.950 345.450 310.050 346.050 ;
        RECT 319.950 345.450 322.050 346.050 ;
        RECT 307.950 344.400 322.050 345.450 ;
        RECT 307.950 343.950 310.050 344.400 ;
        RECT 319.950 343.950 322.050 344.400 ;
        RECT 325.950 344.100 331.050 346.050 ;
        RECT 364.950 345.450 367.050 346.050 ;
        RECT 373.950 345.450 376.050 346.050 ;
        RECT 364.950 344.400 376.050 345.450 ;
        RECT 325.950 343.950 330.000 344.100 ;
        RECT 364.950 343.950 367.050 344.400 ;
        RECT 373.950 343.950 376.050 344.400 ;
        RECT 385.950 343.950 391.050 346.050 ;
        RECT 397.950 343.950 403.050 346.050 ;
        RECT 484.950 345.450 487.050 346.050 ;
        RECT 470.400 345.000 487.050 345.450 ;
        RECT 469.950 344.400 487.050 345.000 ;
        RECT 289.950 342.450 292.050 343.050 ;
        RECT 298.950 342.450 301.050 343.950 ;
        RECT 289.950 341.400 301.050 342.450 ;
        RECT 289.950 340.950 292.050 341.400 ;
        RECT 298.950 340.950 301.050 341.400 ;
        RECT 304.950 342.450 307.050 343.050 ;
        RECT 322.950 342.450 325.050 343.050 ;
        RECT 328.950 342.450 331.050 342.900 ;
        RECT 304.950 341.400 331.050 342.450 ;
        RECT 304.950 340.950 307.050 341.400 ;
        RECT 322.950 340.950 325.050 341.400 ;
        RECT 328.950 340.800 331.050 341.400 ;
        RECT 340.950 340.050 343.050 343.050 ;
        RECT 355.950 342.450 358.050 343.050 ;
        RECT 361.950 342.450 364.050 343.050 ;
        RECT 355.950 341.400 364.050 342.450 ;
        RECT 355.950 340.950 358.050 341.400 ;
        RECT 361.950 340.950 364.050 341.400 ;
        RECT 247.950 339.450 250.050 340.050 ;
        RECT 259.950 339.450 262.050 340.050 ;
        RECT 247.950 338.400 262.050 339.450 ;
        RECT 247.950 337.950 250.050 338.400 ;
        RECT 259.950 337.950 262.050 338.400 ;
        RECT 202.950 336.000 223.050 336.450 ;
        RECT 226.950 336.450 229.050 337.050 ;
        RECT 238.950 336.450 241.050 337.050 ;
        RECT 202.950 335.400 222.450 336.000 ;
        RECT 226.950 335.400 241.050 336.450 ;
        RECT 202.950 334.950 205.050 335.400 ;
        RECT 226.950 334.950 229.050 335.400 ;
        RECT 238.950 334.950 241.050 335.400 ;
        RECT 265.950 334.950 268.050 340.050 ;
        RECT 277.800 339.000 280.050 340.050 ;
        RECT 277.800 337.950 279.900 339.000 ;
        RECT 281.100 337.950 285.900 340.050 ;
        RECT 287.100 337.950 289.200 340.050 ;
        RECT 292.950 337.950 298.050 340.050 ;
        RECT 300.000 339.450 304.050 340.050 ;
        RECT 299.400 337.950 304.050 339.450 ;
        RECT 307.950 339.450 310.050 340.050 ;
        RECT 340.950 339.450 345.900 340.050 ;
        RECT 307.950 338.400 345.900 339.450 ;
        RECT 307.950 337.950 310.050 338.400 ;
        RECT 342.000 337.950 345.900 338.400 ;
        RECT 347.100 339.450 352.050 340.050 ;
        RECT 373.950 339.450 376.050 343.050 ;
        RECT 388.950 340.950 394.050 343.050 ;
        RECT 347.100 339.000 376.050 339.450 ;
        RECT 347.100 338.400 375.450 339.000 ;
        RECT 347.100 337.950 352.050 338.400 ;
        RECT 271.950 336.450 274.050 337.050 ;
        RECT 299.400 336.450 300.450 337.950 ;
        RECT 271.950 335.400 300.450 336.450 ;
        RECT 271.950 334.950 274.050 335.400 ;
        RECT 376.950 334.950 379.050 340.050 ;
        RECT 406.950 337.950 409.050 343.050 ;
        RECT 421.950 340.950 427.050 343.050 ;
        RECT 445.950 342.450 448.050 343.050 ;
        RECT 463.950 342.450 466.050 343.050 ;
        RECT 445.950 341.400 466.050 342.450 ;
        RECT 445.950 340.950 448.050 341.400 ;
        RECT 463.950 340.950 466.050 341.400 ;
        RECT 469.950 340.950 472.050 344.400 ;
        RECT 484.950 343.950 487.050 344.400 ;
        RECT 490.950 345.450 493.050 346.050 ;
        RECT 514.950 345.450 517.050 346.050 ;
        RECT 528.000 345.450 532.050 346.050 ;
        RECT 490.950 344.400 517.050 345.450 ;
        RECT 490.950 343.950 493.050 344.400 ;
        RECT 514.950 343.950 517.050 344.400 ;
        RECT 527.550 343.950 532.050 345.450 ;
        RECT 523.950 340.050 526.050 343.050 ;
        RECT 527.550 340.050 528.600 343.950 ;
        RECT 577.950 343.050 580.050 346.050 ;
        RECT 583.950 343.950 586.050 346.950 ;
        RECT 415.950 339.450 418.050 340.050 ;
        RECT 427.950 339.450 430.050 340.050 ;
        RECT 415.950 338.400 430.050 339.450 ;
        RECT 415.950 337.950 418.050 338.400 ;
        RECT 427.950 337.950 430.050 338.400 ;
        RECT 436.950 339.450 439.050 340.050 ;
        RECT 442.950 339.450 445.050 340.050 ;
        RECT 436.950 338.400 445.050 339.450 ;
        RECT 436.950 337.950 439.050 338.400 ;
        RECT 442.950 337.950 445.050 338.400 ;
        RECT 442.950 334.950 448.050 337.050 ;
        RECT 448.950 336.450 451.050 340.050 ;
        RECT 454.950 339.450 457.050 340.050 ;
        RECT 460.800 339.450 462.900 340.050 ;
        RECT 454.950 338.400 462.900 339.450 ;
        RECT 454.950 337.950 457.050 338.400 ;
        RECT 460.800 337.950 462.900 338.400 ;
        RECT 464.100 337.950 469.050 340.050 ;
        RECT 472.950 337.950 478.050 340.050 ;
        RECT 490.950 339.450 493.050 340.050 ;
        RECT 505.800 339.450 507.900 340.050 ;
        RECT 490.950 338.400 507.900 339.450 ;
        RECT 490.950 337.950 493.050 338.400 ;
        RECT 505.800 337.950 507.900 338.400 ;
        RECT 509.100 339.450 511.200 340.050 ;
        RECT 514.950 339.450 517.050 340.050 ;
        RECT 509.100 338.400 517.050 339.450 ;
        RECT 509.100 337.950 511.200 338.400 ;
        RECT 514.950 337.950 517.050 338.400 ;
        RECT 523.800 339.000 526.050 340.050 ;
        RECT 523.800 337.950 525.900 339.000 ;
        RECT 527.100 337.950 529.200 340.050 ;
        RECT 529.950 339.450 532.050 343.050 ;
        RECT 538.950 342.450 541.050 343.050 ;
        RECT 556.800 342.450 558.900 343.050 ;
        RECT 538.950 341.400 558.900 342.450 ;
        RECT 538.950 340.950 541.050 341.400 ;
        RECT 556.800 340.950 558.900 341.400 ;
        RECT 560.100 340.950 565.050 343.050 ;
        RECT 577.800 342.000 580.050 343.050 ;
        RECT 577.800 340.950 579.900 342.000 ;
        RECT 581.100 340.950 586.050 343.050 ;
        RECT 595.950 340.950 598.050 346.050 ;
        RECT 616.950 345.450 619.050 346.050 ;
        RECT 646.950 345.450 649.050 346.050 ;
        RECT 616.950 344.400 649.050 345.450 ;
        RECT 553.950 339.450 556.050 340.050 ;
        RECT 529.950 339.000 556.050 339.450 ;
        RECT 530.400 338.400 556.050 339.000 ;
        RECT 484.950 337.050 487.050 337.200 ;
        RECT 457.950 336.450 460.050 337.050 ;
        RECT 448.950 336.000 460.050 336.450 ;
        RECT 449.400 335.400 460.050 336.000 ;
        RECT 457.950 334.950 460.050 335.400 ;
        RECT 484.950 335.100 490.050 337.050 ;
        RECT 486.000 334.950 490.050 335.100 ;
        RECT 505.950 336.450 508.050 337.050 ;
        RECT 511.950 336.450 514.050 337.050 ;
        RECT 505.950 335.400 514.050 336.450 ;
        RECT 505.950 334.950 508.050 335.400 ;
        RECT 511.950 334.950 514.050 335.400 ;
        RECT 523.950 336.450 526.050 337.050 ;
        RECT 529.950 336.450 532.050 337.050 ;
        RECT 543.000 336.450 547.050 337.050 ;
        RECT 523.950 335.400 532.050 336.450 ;
        RECT 523.950 334.950 526.050 335.400 ;
        RECT 529.950 334.950 532.050 335.400 ;
        RECT 542.400 334.950 547.050 336.450 ;
        RECT 553.950 334.950 556.050 338.400 ;
        RECT 559.950 339.450 562.050 340.050 ;
        RECT 571.950 339.450 574.050 340.050 ;
        RECT 559.950 338.400 574.050 339.450 ;
        RECT 559.950 337.950 562.050 338.400 ;
        RECT 571.950 337.950 574.050 338.400 ;
        RECT 586.950 339.450 589.050 340.050 ;
        RECT 592.950 339.450 595.050 340.050 ;
        RECT 597.000 339.450 601.050 340.050 ;
        RECT 586.950 338.400 595.050 339.450 ;
        RECT 586.950 337.950 589.050 338.400 ;
        RECT 592.950 337.950 595.050 338.400 ;
        RECT 596.400 337.950 601.050 339.450 ;
        RECT 601.950 339.450 604.050 343.050 ;
        RECT 616.950 340.950 619.050 344.400 ;
        RECT 646.950 343.950 649.050 344.400 ;
        RECT 652.950 343.950 658.050 346.050 ;
        RECT 661.950 343.950 664.050 349.050 ;
        RECT 622.950 342.450 628.050 343.050 ;
        RECT 658.950 342.450 661.050 343.050 ;
        RECT 622.950 342.000 636.300 342.450 ;
        RECT 658.950 342.000 675.300 342.450 ;
        RECT 622.950 341.400 637.050 342.000 ;
        RECT 622.950 340.950 628.050 341.400 ;
        RECT 634.950 340.050 637.050 341.400 ;
        RECT 658.950 341.400 676.050 342.000 ;
        RECT 658.950 340.950 661.050 341.400 ;
        RECT 673.950 340.050 676.050 341.400 ;
        RECT 676.950 340.950 679.050 346.050 ;
        RECT 682.950 340.950 685.050 346.050 ;
        RECT 691.950 343.950 694.050 349.050 ;
        RECT 712.950 348.450 715.050 349.050 ;
        RECT 724.950 348.450 727.050 349.050 ;
        RECT 712.950 347.400 727.050 348.450 ;
        RECT 712.950 346.950 715.050 347.400 ;
        RECT 724.950 346.950 727.050 347.400 ;
        RECT 754.950 348.450 757.050 349.050 ;
        RECT 775.950 348.450 778.050 349.050 ;
        RECT 805.950 348.450 808.050 349.050 ;
        RECT 754.950 347.400 808.050 348.450 ;
        RECT 754.950 346.950 757.050 347.400 ;
        RECT 775.950 346.950 778.050 347.400 ;
        RECT 805.950 346.950 808.050 347.400 ;
        RECT 814.950 348.450 817.050 349.050 ;
        RECT 844.950 348.450 847.050 349.050 ;
        RECT 814.950 347.400 847.050 348.450 ;
        RECT 814.950 346.950 817.050 347.400 ;
        RECT 844.950 346.950 847.050 347.400 ;
        RECT 706.950 345.450 709.050 346.050 ;
        RECT 695.400 344.400 709.050 345.450 ;
        RECT 695.400 340.050 696.450 344.400 ;
        RECT 706.950 343.950 709.050 344.400 ;
        RECT 700.800 343.050 702.900 343.200 ;
        RECT 721.950 343.050 724.050 346.050 ;
        RECT 727.950 343.950 733.050 346.050 ;
        RECT 745.950 345.450 748.050 346.050 ;
        RECT 781.950 345.450 784.050 346.050 ;
        RECT 796.950 345.450 799.050 346.050 ;
        RECT 745.950 344.400 784.050 345.450 ;
        RECT 791.250 345.000 799.050 345.450 ;
        RECT 745.950 343.950 748.050 344.400 ;
        RECT 697.950 341.100 702.900 343.050 ;
        RECT 704.100 342.450 706.200 343.050 ;
        RECT 715.950 342.450 718.050 343.050 ;
        RECT 704.100 341.400 718.050 342.450 ;
        RECT 697.950 340.950 702.000 341.100 ;
        RECT 704.100 340.950 706.200 341.400 ;
        RECT 715.950 340.950 718.050 341.400 ;
        RECT 721.800 342.000 724.050 343.050 ;
        RECT 721.800 340.950 723.900 342.000 ;
        RECT 725.100 340.950 730.050 343.050 ;
        RECT 736.950 342.450 739.050 343.050 ;
        RECT 742.950 342.450 745.050 343.050 ;
        RECT 736.950 341.400 745.050 342.450 ;
        RECT 736.950 340.950 739.050 341.400 ;
        RECT 742.950 340.950 745.050 341.400 ;
        RECT 760.950 340.950 763.050 344.400 ;
        RECT 781.950 343.950 784.050 344.400 ;
        RECT 790.950 344.400 799.050 345.000 ;
        RECT 790.950 343.050 793.050 344.400 ;
        RECT 796.950 343.950 799.050 344.400 ;
        RECT 811.950 345.450 816.000 346.050 ;
        RECT 829.950 345.450 832.050 346.050 ;
        RECT 811.950 345.000 816.450 345.450 ;
        RECT 829.950 345.000 837.450 345.450 ;
        RECT 811.950 343.950 817.050 345.000 ;
        RECT 829.950 344.400 838.050 345.000 ;
        RECT 829.950 343.950 832.050 344.400 ;
        RECT 766.950 342.450 769.050 343.050 ;
        RECT 772.950 342.450 775.050 343.050 ;
        RECT 766.950 341.400 775.050 342.450 ;
        RECT 766.950 340.950 769.050 341.400 ;
        RECT 772.950 340.950 775.050 341.400 ;
        RECT 784.950 340.950 789.900 343.050 ;
        RECT 790.800 342.000 793.050 343.050 ;
        RECT 794.100 342.450 796.200 343.050 ;
        RECT 808.950 342.450 811.050 343.050 ;
        RECT 790.800 340.950 792.900 342.000 ;
        RECT 794.100 341.400 811.050 342.450 ;
        RECT 794.100 340.950 796.200 341.400 ;
        RECT 808.950 340.950 811.050 341.400 ;
        RECT 814.950 340.950 817.050 343.950 ;
        RECT 823.950 342.450 828.000 343.050 ;
        RECT 823.950 342.000 828.300 342.450 ;
        RECT 823.950 340.950 829.050 342.000 ;
        RECT 761.100 340.050 763.200 340.200 ;
        RECT 826.950 340.050 829.050 340.950 ;
        RECT 829.950 340.050 832.050 343.050 ;
        RECT 835.950 340.950 838.050 344.400 ;
        RECT 610.950 339.450 613.050 340.050 ;
        RECT 619.950 339.450 622.050 340.050 ;
        RECT 601.950 339.000 622.050 339.450 ;
        RECT 602.400 338.400 622.050 339.000 ;
        RECT 610.950 337.950 613.050 338.400 ;
        RECT 619.950 337.950 622.050 338.400 ;
        RECT 625.950 337.950 628.050 340.050 ;
        RECT 634.800 339.000 637.050 340.050 ;
        RECT 637.800 339.000 639.900 340.050 ;
        RECT 641.100 339.450 643.200 340.050 ;
        RECT 646.950 339.450 649.050 340.050 ;
        RECT 634.800 337.950 636.900 339.000 ;
        RECT 637.800 337.950 640.050 339.000 ;
        RECT 641.100 338.400 649.050 339.450 ;
        RECT 641.100 337.950 643.200 338.400 ;
        RECT 646.950 337.950 649.050 338.400 ;
        RECT 673.800 339.000 676.050 340.050 ;
        RECT 678.000 339.900 682.050 340.050 ;
        RECT 673.800 337.950 675.900 339.000 ;
        RECT 677.100 337.950 682.050 339.900 ;
        RECT 577.950 336.450 580.050 337.050 ;
        RECT 596.400 336.450 597.450 337.950 ;
        RECT 577.950 335.400 597.450 336.450 ;
        RECT 604.950 336.450 607.050 337.050 ;
        RECT 613.950 336.450 616.050 337.050 ;
        RECT 604.950 335.400 616.050 336.450 ;
        RECT 577.950 334.950 580.050 335.400 ;
        RECT 604.950 334.950 607.050 335.400 ;
        RECT 613.950 334.950 616.050 335.400 ;
        RECT 118.950 333.450 121.050 334.050 ;
        RECT 211.950 333.450 214.050 334.050 ;
        RECT 118.950 332.400 214.050 333.450 ;
        RECT 118.950 331.950 121.050 332.400 ;
        RECT 211.950 331.950 214.050 332.400 ;
        RECT 46.950 330.450 49.050 331.050 ;
        RECT 67.950 330.450 70.050 331.050 ;
        RECT 46.950 329.400 70.050 330.450 ;
        RECT 46.950 328.950 49.050 329.400 ;
        RECT 67.950 328.950 70.050 329.400 ;
        RECT 112.950 330.450 115.050 331.050 ;
        RECT 235.950 330.450 238.050 331.050 ;
        RECT 112.950 329.400 238.050 330.450 ;
        RECT 112.950 328.950 115.050 329.400 ;
        RECT 235.950 328.950 238.050 329.400 ;
        RECT 277.950 330.450 280.050 331.050 ;
        RECT 331.950 330.450 337.050 331.050 ;
        RECT 277.950 329.400 337.050 330.450 ;
        RECT 277.950 328.950 280.050 329.400 ;
        RECT 331.950 328.950 337.050 329.400 ;
        RECT 382.950 328.950 385.050 334.050 ;
        RECT 430.950 333.450 433.050 334.050 ;
        RECT 484.950 333.450 487.050 333.900 ;
        RECT 430.950 332.400 487.050 333.450 ;
        RECT 430.950 331.950 433.050 332.400 ;
        RECT 484.950 331.800 487.050 332.400 ;
        RECT 514.950 333.450 517.050 334.050 ;
        RECT 542.400 333.450 543.450 334.950 ;
        RECT 626.400 334.050 627.450 337.950 ;
        RECT 637.950 337.050 640.050 337.950 ;
        RECT 677.100 337.800 679.200 337.950 ;
        RECT 637.800 336.000 640.050 337.050 ;
        RECT 637.800 334.950 639.900 336.000 ;
        RECT 685.950 334.950 688.050 340.050 ;
        RECT 694.950 337.950 697.050 340.050 ;
        RECT 700.950 334.950 703.050 340.050 ;
        RECT 706.950 339.450 709.050 340.050 ;
        RECT 712.950 339.450 715.050 340.050 ;
        RECT 706.950 338.400 715.050 339.450 ;
        RECT 706.950 337.950 709.050 338.400 ;
        RECT 712.950 337.950 715.050 338.400 ;
        RECT 721.950 339.450 724.050 340.050 ;
        RECT 736.950 339.450 739.050 340.050 ;
        RECT 721.950 338.400 739.050 339.450 ;
        RECT 721.950 337.950 724.050 338.400 ;
        RECT 736.950 337.950 739.050 338.400 ;
        RECT 745.950 337.950 753.900 340.050 ;
        RECT 755.100 337.950 759.900 340.050 ;
        RECT 761.100 338.100 766.050 340.050 ;
        RECT 762.000 337.950 766.050 338.100 ;
        RECT 724.950 336.450 727.050 337.050 ;
        RECT 742.950 336.450 745.050 337.050 ;
        RECT 724.950 335.400 745.050 336.450 ;
        RECT 724.950 334.950 727.050 335.400 ;
        RECT 742.950 334.950 745.050 335.400 ;
        RECT 760.950 336.450 763.050 336.900 ;
        RECT 769.950 336.450 772.050 340.050 ;
        RECT 775.950 339.450 778.050 340.050 ;
        RECT 781.950 339.450 784.050 340.050 ;
        RECT 775.950 338.400 784.050 339.450 ;
        RECT 775.950 337.950 778.050 338.400 ;
        RECT 781.950 337.950 784.050 338.400 ;
        RECT 787.950 337.050 790.050 340.050 ;
        RECT 793.950 337.950 799.050 340.050 ;
        RECT 802.950 339.450 805.050 340.050 ;
        RECT 811.950 339.450 814.050 340.050 ;
        RECT 802.950 338.400 814.050 339.450 ;
        RECT 802.950 337.950 805.050 338.400 ;
        RECT 811.950 337.950 814.050 338.400 ;
        RECT 817.950 337.950 823.050 340.050 ;
        RECT 826.800 339.000 829.050 340.050 ;
        RECT 829.800 339.000 832.050 340.050 ;
        RECT 826.800 337.950 828.900 339.000 ;
        RECT 829.800 337.950 831.900 339.000 ;
        RECT 833.100 337.950 838.050 340.050 ;
        RECT 760.950 336.000 772.050 336.450 ;
        RECT 784.950 336.000 790.050 337.050 ;
        RECT 799.950 336.450 802.050 337.050 ;
        RECT 817.950 336.450 820.050 337.050 ;
        RECT 760.950 335.400 771.450 336.000 ;
        RECT 784.950 335.400 789.450 336.000 ;
        RECT 799.950 335.400 820.050 336.450 ;
        RECT 827.400 336.450 828.450 337.950 ;
        RECT 827.400 335.400 834.450 336.450 ;
        RECT 760.950 334.800 763.050 335.400 ;
        RECT 784.950 334.950 789.000 335.400 ;
        RECT 799.950 334.950 802.050 335.400 ;
        RECT 817.950 334.950 820.050 335.400 ;
        RECT 514.950 332.400 543.450 333.450 ;
        RECT 544.950 333.450 547.050 334.050 ;
        RECT 589.950 333.450 592.050 334.050 ;
        RECT 544.950 332.400 592.050 333.450 ;
        RECT 514.950 331.950 517.050 332.400 ;
        RECT 544.950 331.950 547.050 332.400 ;
        RECT 589.950 331.950 592.050 332.400 ;
        RECT 610.950 331.050 613.050 334.050 ;
        RECT 626.400 332.400 631.050 334.050 ;
        RECT 627.000 331.950 631.050 332.400 ;
        RECT 697.950 333.450 700.050 334.050 ;
        RECT 736.950 333.450 739.050 334.050 ;
        RECT 697.950 332.400 739.050 333.450 ;
        RECT 697.950 331.950 700.050 332.400 ;
        RECT 736.950 331.950 739.050 332.400 ;
        RECT 754.950 333.450 757.050 334.050 ;
        RECT 775.950 333.450 778.050 334.050 ;
        RECT 754.950 332.400 778.050 333.450 ;
        RECT 754.950 331.950 757.050 332.400 ;
        RECT 775.950 331.950 778.050 332.400 ;
        RECT 820.950 333.450 823.050 334.050 ;
        RECT 829.950 333.450 832.050 334.050 ;
        RECT 820.950 332.400 832.050 333.450 ;
        RECT 820.950 331.950 823.050 332.400 ;
        RECT 829.950 331.950 832.050 332.400 ;
        RECT 412.950 330.450 415.050 331.050 ;
        RECT 424.950 330.450 427.050 331.050 ;
        RECT 412.950 329.400 427.050 330.450 ;
        RECT 412.950 328.950 415.050 329.400 ;
        RECT 424.950 328.950 427.050 329.400 ;
        RECT 478.950 330.450 481.050 331.050 ;
        RECT 520.950 330.450 523.050 331.050 ;
        RECT 574.950 330.450 577.050 331.050 ;
        RECT 478.950 329.400 577.050 330.450 ;
        RECT 478.950 328.950 481.050 329.400 ;
        RECT 520.950 328.950 523.050 329.400 ;
        RECT 574.950 328.950 577.050 329.400 ;
        RECT 604.950 328.950 609.900 331.050 ;
        RECT 610.950 330.000 613.200 331.050 ;
        RECT 611.100 328.950 613.200 330.000 ;
        RECT 673.950 330.450 676.050 331.050 ;
        RECT 715.950 330.450 718.050 331.050 ;
        RECT 769.950 330.450 772.050 331.050 ;
        RECT 673.950 329.400 772.050 330.450 ;
        RECT 673.950 328.950 676.050 329.400 ;
        RECT 715.950 328.950 718.050 329.400 ;
        RECT 769.950 328.950 772.050 329.400 ;
        RECT 787.950 330.450 790.050 331.050 ;
        RECT 802.950 330.450 805.050 331.050 ;
        RECT 787.950 329.400 805.050 330.450 ;
        RECT 787.950 328.950 790.050 329.400 ;
        RECT 802.950 328.950 805.050 329.400 ;
        RECT 808.950 330.450 811.050 331.050 ;
        RECT 833.400 330.450 834.450 335.400 ;
        RECT 808.950 329.400 834.450 330.450 ;
        RECT 808.950 328.950 811.050 329.400 ;
        RECT 181.950 325.050 184.050 328.050 ;
        RECT 187.950 327.450 190.050 328.050 ;
        RECT 214.950 327.450 217.050 328.050 ;
        RECT 355.950 327.450 358.050 328.050 ;
        RECT 187.950 326.400 358.050 327.450 ;
        RECT 187.950 325.950 190.050 326.400 ;
        RECT 214.950 325.950 217.050 326.400 ;
        RECT 355.950 325.950 358.050 326.400 ;
        RECT 370.950 327.450 373.050 328.050 ;
        RECT 376.950 327.450 379.050 328.050 ;
        RECT 370.950 326.400 379.050 327.450 ;
        RECT 370.950 325.950 373.050 326.400 ;
        RECT 376.950 325.950 379.050 326.400 ;
        RECT 436.950 327.450 439.050 328.050 ;
        RECT 442.950 327.450 445.050 328.050 ;
        RECT 511.950 327.450 514.050 328.050 ;
        RECT 436.950 326.400 514.050 327.450 ;
        RECT 436.950 325.950 439.050 326.400 ;
        RECT 442.950 325.950 445.050 326.400 ;
        RECT 511.950 325.950 514.050 326.400 ;
        RECT 526.950 327.450 529.050 328.050 ;
        RECT 622.950 327.450 625.050 328.050 ;
        RECT 748.950 327.450 751.050 328.050 ;
        RECT 526.950 326.400 555.450 327.450 ;
        RECT 526.950 325.950 529.050 326.400 ;
        RECT 181.950 324.000 187.050 325.050 ;
        RECT 182.400 323.400 187.050 324.000 ;
        RECT 183.000 322.950 187.050 323.400 ;
        RECT 190.950 324.450 193.050 325.050 ;
        RECT 202.950 324.450 205.050 325.050 ;
        RECT 190.950 323.400 205.050 324.450 ;
        RECT 190.950 322.950 193.050 323.400 ;
        RECT 202.950 322.950 205.050 323.400 ;
        RECT 295.950 324.450 298.050 325.050 ;
        RECT 310.950 324.450 313.050 325.050 ;
        RECT 371.400 324.450 372.450 325.950 ;
        RECT 554.400 325.050 555.450 326.400 ;
        RECT 622.950 326.400 751.050 327.450 ;
        RECT 622.950 325.950 625.050 326.400 ;
        RECT 748.950 325.950 751.050 326.400 ;
        RECT 784.950 327.450 787.050 328.050 ;
        RECT 811.950 327.450 814.050 328.050 ;
        RECT 784.950 326.400 814.050 327.450 ;
        RECT 784.950 325.950 787.050 326.400 ;
        RECT 811.950 325.950 814.050 326.400 ;
        RECT 841.950 325.950 844.050 331.050 ;
        RECT 295.950 323.400 372.450 324.450 ;
        RECT 295.950 322.950 298.050 323.400 ;
        RECT 310.950 322.950 313.050 323.400 ;
        RECT 4.950 321.450 7.050 322.050 ;
        RECT 16.950 321.450 19.050 322.050 ;
        RECT 4.950 320.400 19.050 321.450 ;
        RECT 4.950 319.950 7.050 320.400 ;
        RECT 16.950 319.950 19.050 320.400 ;
        RECT 64.950 319.950 70.050 322.050 ;
        RECT 247.950 321.450 250.050 322.050 ;
        RECT 283.950 321.450 286.050 322.050 ;
        RECT 247.950 320.400 286.050 321.450 ;
        RECT 247.950 319.950 250.050 320.400 ;
        RECT 283.950 319.950 286.050 320.400 ;
        RECT 301.950 321.450 304.050 322.050 ;
        RECT 421.950 321.450 424.050 322.050 ;
        RECT 301.950 320.400 424.050 321.450 ;
        RECT 301.950 319.950 304.050 320.400 ;
        RECT 421.950 319.950 424.050 320.400 ;
        RECT 10.950 318.450 13.050 319.050 ;
        RECT 22.950 318.450 25.050 319.050 ;
        RECT 10.950 317.400 25.050 318.450 ;
        RECT 10.950 316.950 13.050 317.400 ;
        RECT 22.950 316.950 25.050 317.400 ;
        RECT 34.950 318.450 37.050 319.050 ;
        RECT 55.950 318.450 58.050 319.050 ;
        RECT 34.950 317.400 58.050 318.450 ;
        RECT 34.950 316.950 37.050 317.400 ;
        RECT 55.950 316.950 58.050 317.400 ;
        RECT 61.950 318.450 64.050 319.050 ;
        RECT 106.950 318.450 109.050 319.050 ;
        RECT 142.950 318.450 145.050 319.050 ;
        RECT 61.950 317.400 145.050 318.450 ;
        RECT 61.950 316.950 64.050 317.400 ;
        RECT 106.950 316.950 109.050 317.400 ;
        RECT 142.950 316.950 145.050 317.400 ;
        RECT 172.950 318.450 175.050 319.050 ;
        RECT 190.950 318.450 193.050 319.050 ;
        RECT 172.950 317.400 193.050 318.450 ;
        RECT 172.950 316.950 175.050 317.400 ;
        RECT 190.950 316.950 193.050 317.400 ;
        RECT 223.950 318.450 226.050 319.050 ;
        RECT 256.950 318.450 259.050 319.050 ;
        RECT 223.950 317.400 259.050 318.450 ;
        RECT 223.950 316.950 226.050 317.400 ;
        RECT 256.950 316.950 259.050 317.400 ;
        RECT 313.950 318.450 316.050 319.050 ;
        RECT 337.950 318.450 340.050 319.050 ;
        RECT 313.950 317.400 340.050 318.450 ;
        RECT 313.950 316.950 316.050 317.400 ;
        RECT 337.950 316.950 340.050 317.400 ;
        RECT 364.950 318.450 367.050 319.050 ;
        RECT 376.950 318.450 379.050 319.050 ;
        RECT 364.950 317.400 379.050 318.450 ;
        RECT 364.950 316.950 367.050 317.400 ;
        RECT 376.950 316.950 379.050 317.400 ;
        RECT 439.950 316.950 442.050 322.050 ;
        RECT 463.950 321.450 466.050 322.050 ;
        RECT 490.950 321.450 493.050 322.050 ;
        RECT 463.950 320.400 493.050 321.450 ;
        RECT 463.950 319.950 466.050 320.400 ;
        RECT 490.950 319.950 493.050 320.400 ;
        RECT 496.950 319.950 499.050 325.050 ;
        RECT 505.950 324.450 508.050 325.050 ;
        RECT 547.950 324.450 550.050 325.050 ;
        RECT 505.950 323.400 550.050 324.450 ;
        RECT 505.950 322.950 508.050 323.400 ;
        RECT 547.950 322.950 550.050 323.400 ;
        RECT 553.950 324.450 556.050 325.050 ;
        RECT 586.950 324.450 589.050 325.050 ;
        RECT 553.950 323.400 589.050 324.450 ;
        RECT 553.950 322.950 556.050 323.400 ;
        RECT 586.950 322.950 589.050 323.400 ;
        RECT 595.950 324.450 598.050 325.050 ;
        RECT 601.950 324.450 604.050 325.050 ;
        RECT 595.950 323.400 604.050 324.450 ;
        RECT 595.950 322.950 598.050 323.400 ;
        RECT 601.950 322.950 604.050 323.400 ;
        RECT 607.950 324.450 610.050 325.050 ;
        RECT 667.950 324.450 670.050 325.200 ;
        RECT 607.950 323.400 670.050 324.450 ;
        RECT 607.950 322.950 610.050 323.400 ;
        RECT 667.950 323.100 670.050 323.400 ;
        RECT 731.100 324.450 733.200 325.050 ;
        RECT 736.950 324.450 739.050 325.050 ;
        RECT 769.950 324.450 772.050 325.050 ;
        RECT 731.100 323.400 739.050 324.450 ;
        RECT 731.100 322.950 733.200 323.400 ;
        RECT 736.950 322.950 739.050 323.400 ;
        RECT 743.400 323.400 772.050 324.450 ;
        RECT 538.950 321.450 541.050 322.050 ;
        RECT 622.950 321.450 625.050 322.050 ;
        RECT 538.950 320.400 625.050 321.450 ;
        RECT 538.950 319.950 541.050 320.400 ;
        RECT 622.950 319.950 625.050 320.400 ;
        RECT 640.950 319.950 646.050 322.050 ;
        RECT 667.950 321.450 670.050 321.900 ;
        RECT 691.950 321.450 694.050 322.050 ;
        RECT 667.950 320.400 694.050 321.450 ;
        RECT 667.950 319.800 670.050 320.400 ;
        RECT 691.950 319.950 694.050 320.400 ;
        RECT 697.950 319.950 703.050 322.050 ;
        RECT 721.950 321.450 724.050 322.050 ;
        RECT 743.400 321.450 744.450 323.400 ;
        RECT 769.950 322.950 772.050 323.400 ;
        RECT 796.950 321.450 799.050 322.050 ;
        RECT 805.950 321.450 808.050 322.050 ;
        RECT 721.950 320.400 744.450 321.450 ;
        RECT 746.400 320.400 795.450 321.450 ;
        RECT 721.950 319.950 724.050 320.400 ;
        RECT 481.950 318.450 484.050 319.050 ;
        RECT 499.950 318.450 502.050 319.050 ;
        RECT 481.950 317.400 502.050 318.450 ;
        RECT 481.950 316.950 484.050 317.400 ;
        RECT 499.950 316.950 502.050 317.400 ;
        RECT 556.950 318.450 559.050 319.050 ;
        RECT 571.950 318.450 574.050 319.050 ;
        RECT 556.950 317.400 574.050 318.450 ;
        RECT 556.950 316.950 559.050 317.400 ;
        RECT 571.950 316.950 574.050 317.400 ;
        RECT 595.800 318.000 597.900 319.050 ;
        RECT 599.100 318.450 601.200 319.050 ;
        RECT 664.950 318.450 667.050 319.200 ;
        RECT 746.400 319.050 747.450 320.400 ;
        RECT 673.950 318.450 676.050 319.050 ;
        RECT 595.800 316.950 598.050 318.000 ;
        RECT 599.100 317.400 633.450 318.450 ;
        RECT 599.100 316.950 601.200 317.400 ;
        RECT 17.100 315.000 19.200 316.050 ;
        RECT 16.950 313.950 19.200 315.000 ;
        RECT 25.950 315.450 28.050 316.050 ;
        RECT 35.400 315.450 36.450 316.950 ;
        RECT 118.950 315.450 121.050 316.050 ;
        RECT 25.950 314.400 36.450 315.450 ;
        RECT 104.400 315.000 121.050 315.450 ;
        RECT 103.950 314.400 121.050 315.000 ;
        RECT 25.950 313.950 28.050 314.400 ;
        RECT 16.950 313.050 19.050 313.950 ;
        RECT 61.950 313.050 64.050 313.200 ;
        RECT 10.950 310.950 15.900 313.050 ;
        RECT 16.950 312.450 19.200 313.050 ;
        RECT 16.950 312.000 30.600 312.450 ;
        RECT 17.100 311.400 31.050 312.000 ;
        RECT 17.100 310.950 19.200 311.400 ;
        RECT 28.950 310.050 31.050 311.400 ;
        RECT 4.950 309.450 7.050 310.050 ;
        RECT 13.950 309.450 16.050 310.050 ;
        RECT 4.950 308.400 16.050 309.450 ;
        RECT 4.950 307.950 7.050 308.400 ;
        RECT 13.950 307.950 16.050 308.400 ;
        RECT 19.950 309.450 22.050 310.050 ;
        RECT 25.800 309.450 27.900 310.050 ;
        RECT 19.950 308.400 27.900 309.450 ;
        RECT 28.950 309.000 31.200 310.050 ;
        RECT 19.950 307.950 22.050 308.400 ;
        RECT 25.800 307.950 27.900 308.400 ;
        RECT 29.100 307.950 31.200 309.000 ;
        RECT 34.950 307.950 37.050 313.050 ;
        RECT 40.950 312.450 43.050 313.050 ;
        RECT 49.950 312.450 52.050 313.050 ;
        RECT 40.950 311.400 52.050 312.450 ;
        RECT 40.950 310.950 43.050 311.400 ;
        RECT 49.950 310.950 52.050 311.400 ;
        RECT 58.950 311.100 64.050 313.050 ;
        RECT 67.950 312.450 70.050 313.050 ;
        RECT 76.950 312.450 79.050 313.050 ;
        RECT 67.950 311.400 79.050 312.450 ;
        RECT 58.950 310.950 63.000 311.100 ;
        RECT 67.950 310.950 70.050 311.400 ;
        RECT 76.950 310.950 79.050 311.400 ;
        RECT 82.950 310.950 88.050 313.050 ;
        RECT 103.950 310.950 106.050 314.400 ;
        RECT 118.950 313.950 121.050 314.400 ;
        RECT 127.950 315.450 130.050 316.050 ;
        RECT 148.950 315.450 151.050 316.050 ;
        RECT 127.950 314.400 151.050 315.450 ;
        RECT 127.950 313.950 130.050 314.400 ;
        RECT 148.950 313.950 151.050 314.400 ;
        RECT 166.950 315.450 169.050 316.050 ;
        RECT 199.950 315.450 202.050 316.050 ;
        RECT 214.950 315.450 220.050 316.050 ;
        RECT 166.950 314.400 177.450 315.450 ;
        RECT 166.950 313.950 169.050 314.400 ;
        RECT 43.950 309.450 46.050 310.050 ;
        RECT 55.800 309.450 57.900 310.050 ;
        RECT 43.950 308.400 57.900 309.450 ;
        RECT 43.950 307.950 46.050 308.400 ;
        RECT 55.800 307.950 57.900 308.400 ;
        RECT 59.100 307.950 64.050 310.050 ;
        RECT 4.950 303.450 7.050 304.050 ;
        RECT 31.950 303.450 34.050 307.050 ;
        RECT 40.950 306.450 43.050 307.050 ;
        RECT 70.950 306.450 73.050 307.050 ;
        RECT 73.950 306.450 76.050 310.050 ;
        RECT 40.950 306.000 76.050 306.450 ;
        RECT 40.950 305.400 75.450 306.000 ;
        RECT 40.950 304.950 43.050 305.400 ;
        RECT 70.950 304.950 73.050 305.400 ;
        RECT 79.950 304.950 82.050 310.050 ;
        RECT 97.800 309.000 99.900 310.050 ;
        RECT 101.100 309.450 103.200 310.050 ;
        RECT 115.950 309.450 118.050 310.050 ;
        RECT 97.800 307.950 100.050 309.000 ;
        RECT 101.100 308.400 118.050 309.450 ;
        RECT 101.100 307.950 103.200 308.400 ;
        RECT 115.950 307.950 118.050 308.400 ;
        RECT 124.950 309.450 127.050 310.050 ;
        RECT 133.950 309.450 136.050 310.050 ;
        RECT 124.950 308.400 136.050 309.450 ;
        RECT 124.950 307.950 127.050 308.400 ;
        RECT 133.950 307.950 136.050 308.400 ;
        RECT 142.950 309.450 145.050 310.050 ;
        RECT 154.950 309.450 157.050 310.050 ;
        RECT 142.950 308.400 157.050 309.450 ;
        RECT 142.950 307.950 145.050 308.400 ;
        RECT 154.950 307.950 157.050 308.400 ;
        RECT 172.950 307.950 175.050 313.050 ;
        RECT 176.400 312.450 177.450 314.400 ;
        RECT 199.950 314.400 220.050 315.450 ;
        RECT 199.950 313.950 202.050 314.400 ;
        RECT 214.950 313.950 220.050 314.400 ;
        RECT 176.400 311.400 207.450 312.450 ;
        RECT 178.950 307.950 181.050 311.400 ;
        RECT 206.400 310.050 207.450 311.400 ;
        RECT 223.950 310.950 229.050 313.050 ;
        RECT 232.950 310.950 235.050 316.050 ;
        RECT 247.950 315.450 250.050 316.050 ;
        RECT 253.950 315.450 256.050 316.050 ;
        RECT 239.400 315.000 256.050 315.450 ;
        RECT 238.950 314.400 256.050 315.000 ;
        RECT 238.950 310.950 241.050 314.400 ;
        RECT 247.950 313.950 250.050 314.400 ;
        RECT 253.950 313.950 256.050 314.400 ;
        RECT 271.950 315.450 276.000 316.050 ;
        RECT 280.950 315.450 283.050 316.050 ;
        RECT 271.950 315.000 276.450 315.450 ;
        RECT 271.950 313.950 277.050 315.000 ;
        RECT 280.950 314.400 297.450 315.450 ;
        RECT 280.950 313.950 283.050 314.400 ;
        RECT 256.950 312.450 259.050 313.050 ;
        RECT 268.950 312.450 271.050 313.050 ;
        RECT 256.950 311.400 271.050 312.450 ;
        RECT 256.950 310.950 259.050 311.400 ;
        RECT 268.950 310.950 271.050 311.400 ;
        RECT 274.950 310.950 277.050 313.950 ;
        RECT 280.950 310.950 286.050 313.050 ;
        RECT 296.400 310.050 297.450 314.400 ;
        RECT 310.950 310.950 313.050 316.050 ;
        RECT 316.950 310.950 319.050 316.050 ;
        RECT 338.400 315.450 339.450 316.950 ;
        RECT 412.950 315.450 415.050 316.050 ;
        RECT 421.950 315.450 424.050 316.050 ;
        RECT 338.400 314.400 375.450 315.450 ;
        RECT 367.950 310.950 373.050 313.050 ;
        RECT 374.400 310.050 375.450 314.400 ;
        RECT 412.950 314.400 424.050 315.450 ;
        RECT 412.950 313.950 415.050 314.400 ;
        RECT 421.950 313.950 424.050 314.400 ;
        RECT 451.950 315.450 454.050 316.050 ;
        RECT 469.950 315.450 472.050 316.050 ;
        RECT 451.950 314.400 504.450 315.450 ;
        RECT 451.950 313.950 454.050 314.400 ;
        RECT 469.950 313.950 472.050 314.400 ;
        RECT 376.950 310.950 382.050 313.050 ;
        RECT 385.950 312.450 388.050 313.200 ;
        RECT 466.800 313.050 468.900 313.200 ;
        RECT 503.400 313.050 504.450 314.400 ;
        RECT 547.950 313.950 553.050 316.050 ;
        RECT 595.950 313.950 598.050 316.950 ;
        RECT 601.950 315.450 604.050 316.050 ;
        RECT 607.950 315.450 610.050 316.050 ;
        RECT 601.950 314.400 610.050 315.450 ;
        RECT 601.950 313.950 604.050 314.400 ;
        RECT 607.950 313.950 610.050 314.400 ;
        RECT 391.950 312.450 394.050 313.050 ;
        RECT 385.950 311.400 394.050 312.450 ;
        RECT 385.950 311.100 388.050 311.400 ;
        RECT 391.950 310.950 394.050 311.400 ;
        RECT 400.950 310.950 406.050 313.050 ;
        RECT 454.950 312.450 457.050 313.050 ;
        RECT 463.950 312.450 468.900 313.050 ;
        RECT 454.950 311.400 468.900 312.450 ;
        RECT 454.950 310.950 457.050 311.400 ;
        RECT 463.950 311.100 468.900 311.400 ;
        RECT 470.100 312.450 472.200 313.050 ;
        RECT 470.100 311.400 501.450 312.450 ;
        RECT 503.400 311.400 508.050 313.050 ;
        RECT 463.950 310.950 468.000 311.100 ;
        RECT 470.100 310.950 472.200 311.400 ;
        RECT 500.400 310.050 501.450 311.400 ;
        RECT 504.000 310.950 508.050 311.400 ;
        RECT 523.950 310.950 528.900 313.050 ;
        RECT 530.100 310.950 535.050 313.050 ;
        RECT 572.100 312.450 574.200 313.050 ;
        RECT 592.950 312.450 595.050 313.050 ;
        RECT 572.100 311.400 595.050 312.450 ;
        RECT 572.100 310.950 574.200 311.400 ;
        RECT 592.950 310.950 595.050 311.400 ;
        RECT 625.950 310.950 631.050 313.050 ;
        RECT 632.400 310.050 633.450 317.400 ;
        RECT 664.950 317.400 676.050 318.450 ;
        RECT 664.950 317.100 667.050 317.400 ;
        RECT 673.950 316.950 676.050 317.400 ;
        RECT 685.950 318.450 688.050 319.050 ;
        RECT 706.950 318.450 709.050 319.050 ;
        RECT 745.950 318.450 748.050 319.050 ;
        RECT 685.950 317.400 709.050 318.450 ;
        RECT 685.950 316.950 688.050 317.400 ;
        RECT 706.950 316.950 709.050 317.400 ;
        RECT 710.400 317.400 748.050 318.450 ;
        RECT 664.950 315.450 667.050 315.900 ;
        RECT 710.400 315.450 711.450 317.400 ;
        RECT 745.950 316.950 748.050 317.400 ;
        RECT 763.950 318.450 766.050 319.050 ;
        RECT 784.950 318.450 787.050 319.050 ;
        RECT 763.950 317.400 787.050 318.450 ;
        RECT 794.400 318.450 795.450 320.400 ;
        RECT 796.950 320.400 808.050 321.450 ;
        RECT 820.950 321.450 823.050 325.050 ;
        RECT 841.950 321.450 844.050 322.050 ;
        RECT 820.950 321.000 844.050 321.450 ;
        RECT 821.400 320.400 844.050 321.000 ;
        RECT 796.950 319.950 799.050 320.400 ;
        RECT 805.950 319.950 808.050 320.400 ;
        RECT 841.950 319.950 844.050 320.400 ;
        RECT 799.800 318.450 801.900 319.050 ;
        RECT 794.400 317.400 801.900 318.450 ;
        RECT 763.950 316.950 766.050 317.400 ;
        RECT 784.950 316.950 787.050 317.400 ;
        RECT 799.800 316.950 801.900 317.400 ;
        RECT 803.100 318.450 805.200 319.050 ;
        RECT 817.950 318.450 820.050 319.050 ;
        RECT 803.100 317.400 820.050 318.450 ;
        RECT 803.100 316.950 805.200 317.400 ;
        RECT 817.950 316.950 820.050 317.400 ;
        RECT 826.950 318.450 829.050 319.050 ;
        RECT 838.950 318.450 841.050 319.050 ;
        RECT 826.950 317.400 841.050 318.450 ;
        RECT 826.950 316.950 829.050 317.400 ;
        RECT 838.950 316.950 841.050 317.400 ;
        RECT 644.400 314.400 667.050 315.450 ;
        RECT 634.950 310.950 640.050 313.050 ;
        RECT 644.400 310.050 645.450 314.400 ;
        RECT 664.950 313.800 667.050 314.400 ;
        RECT 680.400 314.400 711.450 315.450 ;
        RECT 712.950 315.450 715.050 316.050 ;
        RECT 721.950 315.450 724.050 316.050 ;
        RECT 832.950 315.450 835.050 316.050 ;
        RECT 856.950 315.450 859.050 316.050 ;
        RECT 712.950 314.400 724.050 315.450 ;
        RECT 755.400 315.000 768.450 315.450 ;
        RECT 680.400 313.050 681.450 314.400 ;
        RECT 712.950 313.950 715.050 314.400 ;
        RECT 721.950 313.950 724.050 314.400 ;
        RECT 754.950 314.400 768.450 315.000 ;
        RECT 646.950 310.950 652.050 313.050 ;
        RECT 655.950 312.450 658.050 313.050 ;
        RECT 661.950 312.450 664.050 313.050 ;
        RECT 655.950 311.400 664.050 312.450 ;
        RECT 655.950 310.950 658.050 311.400 ;
        RECT 661.950 310.950 664.050 311.400 ;
        RECT 670.950 312.450 673.050 313.050 ;
        RECT 676.950 312.450 681.450 313.050 ;
        RECT 670.950 311.400 681.450 312.450 ;
        RECT 670.950 310.950 673.050 311.400 ;
        RECT 676.950 310.950 681.000 311.400 ;
        RECT 682.950 310.950 688.050 313.050 ;
        RECT 691.950 312.450 694.050 313.050 ;
        RECT 706.950 312.450 709.050 313.050 ;
        RECT 691.950 311.400 709.050 312.450 ;
        RECT 691.950 310.950 694.050 311.400 ;
        RECT 706.950 310.950 709.050 311.400 ;
        RECT 721.950 310.950 727.050 313.050 ;
        RECT 742.950 312.450 745.050 313.050 ;
        RECT 748.950 312.450 751.050 313.050 ;
        RECT 742.950 311.400 751.050 312.450 ;
        RECT 742.950 310.950 745.050 311.400 ;
        RECT 748.950 310.950 751.050 311.400 ;
        RECT 754.950 310.950 757.050 314.400 ;
        RECT 767.400 313.050 768.450 314.400 ;
        RECT 832.950 314.400 859.050 315.450 ;
        RECT 832.950 313.950 835.050 314.400 ;
        RECT 856.950 313.950 859.050 314.400 ;
        RECT 762.000 312.450 766.050 313.050 ;
        RECT 761.400 310.950 766.050 312.450 ;
        RECT 767.400 311.400 772.050 313.050 ;
        RECT 768.000 310.950 772.050 311.400 ;
        RECT 775.950 312.450 778.050 313.050 ;
        RECT 784.800 312.450 786.900 313.050 ;
        RECT 775.950 311.400 786.900 312.450 ;
        RECT 775.950 310.950 778.050 311.400 ;
        RECT 784.800 310.950 786.900 311.400 ;
        RECT 788.100 310.950 792.900 313.050 ;
        RECT 794.100 312.000 796.200 313.050 ;
        RECT 793.950 310.950 796.200 312.000 ;
        RECT 799.950 312.450 802.050 313.050 ;
        RECT 817.950 312.450 820.050 313.050 ;
        RECT 826.950 312.450 829.050 313.050 ;
        RECT 799.950 311.400 829.050 312.450 ;
        RECT 799.950 310.950 802.050 311.400 ;
        RECT 817.950 310.950 820.050 311.400 ;
        RECT 826.950 310.950 829.050 311.400 ;
        RECT 190.950 307.950 196.050 310.050 ;
        RECT 199.950 307.950 205.050 310.050 ;
        RECT 206.400 308.400 211.050 310.050 ;
        RECT 207.000 307.950 211.050 308.400 ;
        RECT 220.950 309.450 223.050 310.050 ;
        RECT 226.950 309.450 232.050 310.050 ;
        RECT 220.950 308.400 232.050 309.450 ;
        RECT 220.950 307.950 223.050 308.400 ;
        RECT 226.950 307.950 232.050 308.400 ;
        RECT 97.950 306.450 100.050 307.950 ;
        RECT 109.950 306.450 115.050 307.050 ;
        RECT 97.950 306.000 115.050 306.450 ;
        RECT 98.250 305.400 115.050 306.000 ;
        RECT 109.950 304.950 115.050 305.400 ;
        RECT 118.950 304.950 124.050 307.050 ;
        RECT 127.950 304.950 133.050 307.050 ;
        RECT 4.950 303.000 34.050 303.450 ;
        RECT 4.950 302.400 33.450 303.000 ;
        RECT 4.950 301.950 7.050 302.400 ;
        RECT 136.950 301.950 139.050 307.050 ;
        RECT 151.950 303.450 154.050 307.050 ;
        RECT 157.950 304.950 163.050 307.050 ;
        RECT 165.000 306.450 169.050 307.050 ;
        RECT 164.400 304.950 169.050 306.450 ;
        RECT 175.950 306.450 178.050 307.050 ;
        RECT 196.950 306.900 201.000 307.050 ;
        RECT 196.950 306.450 202.050 306.900 ;
        RECT 175.950 305.400 202.050 306.450 ;
        RECT 235.950 306.450 238.050 310.050 ;
        RECT 250.950 307.950 256.050 310.050 ;
        RECT 262.950 309.450 265.050 310.050 ;
        RECT 271.950 309.450 276.900 310.050 ;
        RECT 262.950 308.400 276.900 309.450 ;
        RECT 278.100 309.000 280.200 310.050 ;
        RECT 262.950 307.950 265.050 308.400 ;
        RECT 271.950 307.950 276.900 308.400 ;
        RECT 277.950 307.950 280.200 309.000 ;
        RECT 295.950 307.950 298.050 310.050 ;
        RECT 301.950 307.950 307.050 310.050 ;
        RECT 244.950 306.450 247.050 307.050 ;
        RECT 250.800 306.450 252.900 307.050 ;
        RECT 235.950 306.000 252.900 306.450 ;
        RECT 236.400 305.400 252.900 306.000 ;
        RECT 175.950 304.950 178.050 305.400 ;
        RECT 196.950 304.950 202.050 305.400 ;
        RECT 244.950 304.950 247.050 305.400 ;
        RECT 250.800 304.950 252.900 305.400 ;
        RECT 254.100 304.950 259.050 307.050 ;
        RECT 277.950 306.450 280.050 307.950 ;
        RECT 283.950 306.450 286.050 307.050 ;
        RECT 277.950 306.000 286.050 306.450 ;
        RECT 278.550 305.400 286.050 306.000 ;
        RECT 283.950 304.950 286.050 305.400 ;
        RECT 292.950 304.950 297.900 307.050 ;
        RECT 299.100 306.450 303.000 307.050 ;
        RECT 299.100 304.950 303.450 306.450 ;
        RECT 313.950 304.950 316.050 310.050 ;
        RECT 319.950 304.950 322.050 310.050 ;
        RECT 337.950 309.450 340.050 310.050 ;
        RECT 355.950 309.450 358.050 310.050 ;
        RECT 337.950 308.400 358.050 309.450 ;
        RECT 337.950 307.950 340.050 308.400 ;
        RECT 355.950 307.950 358.050 308.400 ;
        RECT 361.950 307.950 367.050 310.050 ;
        RECT 373.950 307.950 376.050 310.050 ;
        RECT 379.950 309.450 382.050 310.050 ;
        RECT 388.950 309.450 391.050 310.050 ;
        RECT 379.950 308.400 391.050 309.450 ;
        RECT 379.950 307.950 382.050 308.400 ;
        RECT 388.950 307.950 391.050 308.400 ;
        RECT 394.950 307.950 400.050 310.050 ;
        RECT 406.950 309.450 409.050 310.050 ;
        RECT 418.800 309.450 420.900 310.050 ;
        RECT 406.950 308.400 420.900 309.450 ;
        RECT 406.950 307.950 409.050 308.400 ;
        RECT 418.800 307.950 420.900 308.400 ;
        RECT 422.100 309.450 424.200 310.050 ;
        RECT 430.950 309.450 433.050 310.050 ;
        RECT 422.100 308.400 433.050 309.450 ;
        RECT 422.100 307.950 424.200 308.400 ;
        RECT 430.950 307.950 433.050 308.400 ;
        RECT 439.950 309.450 442.050 310.050 ;
        RECT 448.950 309.450 451.050 310.050 ;
        RECT 465.000 309.900 469.050 310.050 ;
        RECT 439.950 308.400 451.050 309.450 ;
        RECT 439.950 307.950 442.050 308.400 ;
        RECT 448.950 307.950 451.050 308.400 ;
        RECT 463.950 307.950 469.050 309.900 ;
        RECT 472.950 309.450 475.050 310.050 ;
        RECT 487.800 309.450 489.900 310.050 ;
        RECT 472.950 308.400 489.900 309.450 ;
        RECT 491.100 309.000 493.200 310.050 ;
        RECT 472.950 307.950 475.050 308.400 ;
        RECT 487.800 307.950 489.900 308.400 ;
        RECT 490.950 307.950 493.200 309.000 ;
        RECT 500.400 308.400 505.050 310.050 ;
        RECT 501.000 307.950 505.050 308.400 ;
        RECT 508.950 307.950 514.050 310.050 ;
        RECT 463.950 307.800 466.050 307.950 ;
        RECT 331.950 304.950 337.050 307.050 ;
        RECT 358.950 306.450 361.050 307.050 ;
        RECT 409.950 306.450 412.050 307.050 ;
        RECT 358.950 305.400 412.050 306.450 ;
        RECT 358.950 304.950 361.050 305.400 ;
        RECT 409.950 304.950 412.050 305.400 ;
        RECT 427.950 306.450 430.050 307.050 ;
        RECT 445.950 306.450 451.050 307.050 ;
        RECT 427.950 305.400 451.050 306.450 ;
        RECT 427.950 304.950 430.050 305.400 ;
        RECT 445.950 304.950 451.050 305.400 ;
        RECT 481.950 304.950 487.050 307.050 ;
        RECT 490.950 304.950 493.050 307.950 ;
        RECT 526.950 304.950 529.050 310.050 ;
        RECT 532.950 306.450 535.050 310.050 ;
        RECT 538.950 309.450 541.050 310.050 ;
        RECT 568.950 309.450 571.050 310.050 ;
        RECT 538.950 308.400 571.050 309.450 ;
        RECT 538.950 307.950 541.050 308.400 ;
        RECT 568.950 307.950 571.050 308.400 ;
        RECT 574.950 307.950 580.050 310.050 ;
        RECT 583.800 309.000 585.900 310.050 ;
        RECT 583.800 307.950 586.050 309.000 ;
        RECT 587.100 307.950 592.050 310.050 ;
        RECT 604.950 307.950 609.900 310.050 ;
        RECT 611.100 309.450 616.050 310.050 ;
        RECT 625.950 309.450 628.050 310.050 ;
        RECT 611.100 308.400 628.050 309.450 ;
        RECT 611.100 307.950 616.050 308.400 ;
        RECT 625.950 307.950 628.050 308.400 ;
        RECT 631.950 307.950 634.050 310.050 ;
        RECT 644.400 308.400 649.050 310.050 ;
        RECT 645.000 307.950 649.050 308.400 ;
        RECT 652.950 309.450 655.050 310.050 ;
        RECT 661.950 309.450 664.050 310.050 ;
        RECT 652.950 308.400 664.050 309.450 ;
        RECT 652.950 307.950 655.050 308.400 ;
        RECT 661.950 307.950 664.050 308.400 ;
        RECT 670.950 307.950 676.050 310.050 ;
        RECT 679.950 309.450 682.050 310.050 ;
        RECT 688.950 309.450 691.050 310.050 ;
        RECT 679.950 308.400 691.050 309.450 ;
        RECT 679.950 307.950 682.050 308.400 ;
        RECT 688.950 307.950 691.050 308.400 ;
        RECT 694.950 309.450 697.050 310.050 ;
        RECT 709.950 309.450 712.050 310.050 ;
        RECT 694.950 308.400 712.050 309.450 ;
        RECT 694.950 307.950 697.050 308.400 ;
        RECT 709.950 307.950 712.050 308.400 ;
        RECT 730.950 309.450 733.050 310.050 ;
        RECT 745.950 309.450 748.050 310.050 ;
        RECT 730.950 308.400 748.050 309.450 ;
        RECT 730.950 307.950 733.050 308.400 ;
        RECT 745.950 307.950 748.050 308.400 ;
        RECT 751.950 309.450 754.050 310.050 ;
        RECT 757.950 309.450 760.050 310.050 ;
        RECT 751.950 308.400 760.050 309.450 ;
        RECT 751.950 307.950 754.050 308.400 ;
        RECT 757.950 307.950 760.050 308.400 ;
        RECT 538.950 306.450 541.050 307.050 ;
        RECT 532.950 306.000 541.050 306.450 ;
        RECT 533.400 305.400 541.050 306.000 ;
        RECT 164.400 303.450 165.450 304.950 ;
        RECT 199.950 304.800 202.050 304.950 ;
        RECT 151.950 303.000 165.450 303.450 ;
        RECT 152.400 302.400 165.450 303.000 ;
        RECT 302.400 303.450 303.450 304.950 ;
        RECT 316.800 303.450 318.900 304.050 ;
        RECT 302.400 302.400 318.900 303.450 ;
        RECT 316.800 301.950 318.900 302.400 ;
        RECT 320.100 303.450 322.200 304.050 ;
        RECT 340.950 303.450 343.050 304.050 ;
        RECT 320.100 302.400 343.050 303.450 ;
        RECT 320.100 301.950 322.200 302.400 ;
        RECT 340.950 301.950 343.050 302.400 ;
        RECT 415.950 303.450 418.050 304.050 ;
        RECT 451.950 303.450 454.050 304.050 ;
        RECT 415.950 302.400 454.050 303.450 ;
        RECT 415.950 301.950 418.050 302.400 ;
        RECT 451.950 301.950 454.050 302.400 ;
        RECT 484.950 303.450 487.050 304.050 ;
        RECT 505.950 303.450 508.050 304.050 ;
        RECT 484.950 302.400 508.050 303.450 ;
        RECT 533.400 303.000 534.450 305.400 ;
        RECT 538.950 304.950 541.050 305.400 ;
        RECT 559.950 304.950 565.050 307.050 ;
        RECT 571.950 306.900 576.000 307.050 ;
        RECT 571.950 304.950 577.050 306.900 ;
        RECT 583.950 304.950 586.050 307.950 ;
        RECT 589.950 304.950 592.050 307.050 ;
        RECT 574.950 304.800 577.050 304.950 ;
        RECT 536.100 303.450 538.200 304.050 ;
        RECT 544.950 303.450 547.050 304.050 ;
        RECT 484.950 301.950 487.050 302.400 ;
        RECT 505.950 301.950 508.050 302.400 ;
        RECT 85.950 300.450 88.050 301.050 ;
        RECT 124.950 300.450 127.050 301.050 ;
        RECT 85.950 299.400 127.050 300.450 ;
        RECT 85.950 298.950 88.050 299.400 ;
        RECT 124.950 298.950 127.050 299.400 ;
        RECT 136.950 300.450 139.050 301.050 ;
        RECT 184.950 300.450 187.050 301.050 ;
        RECT 136.950 299.400 187.050 300.450 ;
        RECT 136.950 298.950 139.050 299.400 ;
        RECT 184.950 298.950 187.050 299.400 ;
        RECT 235.950 300.450 238.050 301.050 ;
        RECT 250.950 300.450 253.050 301.050 ;
        RECT 235.950 299.400 253.050 300.450 ;
        RECT 235.950 298.950 238.050 299.400 ;
        RECT 250.950 298.950 253.050 299.400 ;
        RECT 283.950 300.450 286.050 301.050 ;
        RECT 298.950 300.450 301.050 301.050 ;
        RECT 283.950 299.400 301.050 300.450 ;
        RECT 341.400 300.450 342.450 301.950 ;
        RECT 400.950 300.450 403.050 301.050 ;
        RECT 341.400 299.400 403.050 300.450 ;
        RECT 283.950 298.950 286.050 299.400 ;
        RECT 298.950 298.950 301.050 299.400 ;
        RECT 400.950 298.950 403.050 299.400 ;
        RECT 421.950 300.450 424.050 301.050 ;
        RECT 427.950 300.450 433.050 301.050 ;
        RECT 421.950 299.400 433.050 300.450 ;
        RECT 421.950 298.950 424.050 299.400 ;
        RECT 427.950 298.950 433.050 299.400 ;
        RECT 532.950 298.950 535.050 303.000 ;
        RECT 536.100 302.400 547.050 303.450 ;
        RECT 536.100 301.950 538.200 302.400 ;
        RECT 544.950 301.950 547.050 302.400 ;
        RECT 590.400 300.450 591.450 304.950 ;
        RECT 595.950 301.950 598.050 307.050 ;
        RECT 604.950 306.450 609.000 307.050 ;
        RECT 610.950 306.450 613.050 307.050 ;
        RECT 622.950 306.450 625.050 307.050 ;
        RECT 604.950 304.950 609.450 306.450 ;
        RECT 610.950 305.400 625.050 306.450 ;
        RECT 610.950 304.950 613.050 305.400 ;
        RECT 622.950 304.950 625.050 305.400 ;
        RECT 628.950 306.450 631.050 307.050 ;
        RECT 655.950 306.450 658.050 307.050 ;
        RECT 628.950 305.400 658.050 306.450 ;
        RECT 628.950 304.950 631.050 305.400 ;
        RECT 655.950 304.950 658.050 305.400 ;
        RECT 712.950 306.450 715.050 307.050 ;
        RECT 718.800 306.450 720.900 307.050 ;
        RECT 712.950 305.400 720.900 306.450 ;
        RECT 712.950 304.950 715.050 305.400 ;
        RECT 718.800 304.950 720.900 305.400 ;
        RECT 722.100 306.450 724.200 307.050 ;
        RECT 727.800 306.450 729.900 307.050 ;
        RECT 722.100 305.400 729.900 306.450 ;
        RECT 722.100 304.950 724.200 305.400 ;
        RECT 727.800 304.950 729.900 305.400 ;
        RECT 737.100 306.450 739.200 307.050 ;
        RECT 761.400 306.450 762.450 310.950 ;
        RECT 766.950 307.950 771.900 310.050 ;
        RECT 773.100 309.000 775.200 310.050 ;
        RECT 772.950 307.950 775.200 309.000 ;
        RECT 737.100 305.400 762.450 306.450 ;
        RECT 772.950 306.450 775.050 307.950 ;
        RECT 787.950 306.450 790.050 310.050 ;
        RECT 793.950 307.950 796.050 310.950 ;
        RECT 832.950 310.050 835.050 313.050 ;
        RECT 802.950 309.450 805.050 310.050 ;
        RECT 811.950 309.450 814.050 310.050 ;
        RECT 802.950 308.400 814.050 309.450 ;
        RECT 802.950 307.950 805.050 308.400 ;
        RECT 811.950 307.950 814.050 308.400 ;
        RECT 832.950 307.950 838.050 310.050 ;
        RECT 799.950 306.450 805.050 307.050 ;
        RECT 772.950 306.000 780.450 306.450 ;
        RECT 787.950 306.000 805.050 306.450 ;
        RECT 773.550 305.400 780.450 306.000 ;
        RECT 788.400 305.400 805.050 306.000 ;
        RECT 737.100 304.950 739.200 305.400 ;
        RECT 608.400 303.450 609.450 304.950 ;
        RECT 637.950 303.450 640.050 304.050 ;
        RECT 608.400 302.400 640.050 303.450 ;
        RECT 637.950 301.950 640.050 302.400 ;
        RECT 649.950 303.450 652.050 304.050 ;
        RECT 685.950 303.450 688.050 304.050 ;
        RECT 649.950 302.400 688.050 303.450 ;
        RECT 649.950 301.950 652.050 302.400 ;
        RECT 685.950 301.950 688.050 302.400 ;
        RECT 697.950 303.450 700.050 304.050 ;
        RECT 721.950 303.450 724.050 304.050 ;
        RECT 697.950 302.400 724.050 303.450 ;
        RECT 697.950 301.950 700.050 302.400 ;
        RECT 721.950 301.950 724.050 302.400 ;
        RECT 727.950 303.450 730.050 304.050 ;
        RECT 775.950 303.450 778.050 304.200 ;
        RECT 727.950 302.400 778.050 303.450 ;
        RECT 779.400 303.450 780.450 305.400 ;
        RECT 799.950 304.950 805.050 305.400 ;
        RECT 850.950 304.950 853.050 310.050 ;
        RECT 793.950 303.450 796.050 304.050 ;
        RECT 841.950 303.450 844.050 304.050 ;
        RECT 779.400 302.400 844.050 303.450 ;
        RECT 727.950 301.950 730.050 302.400 ;
        RECT 775.950 302.100 778.050 302.400 ;
        RECT 793.950 301.950 796.050 302.400 ;
        RECT 841.950 301.950 844.050 302.400 ;
        RECT 847.950 303.450 850.050 304.050 ;
        RECT 853.950 303.450 856.050 304.050 ;
        RECT 847.950 302.400 856.050 303.450 ;
        RECT 847.950 301.950 850.050 302.400 ;
        RECT 853.950 301.950 856.050 302.400 ;
        RECT 604.950 300.450 607.050 301.050 ;
        RECT 590.400 299.400 607.050 300.450 ;
        RECT 604.950 298.950 607.050 299.400 ;
        RECT 625.950 300.450 628.050 301.200 ;
        RECT 646.950 300.450 649.050 301.050 ;
        RECT 625.950 299.400 649.050 300.450 ;
        RECT 625.950 299.100 628.050 299.400 ;
        RECT 646.950 298.950 649.050 299.400 ;
        RECT 670.950 300.450 673.050 301.050 ;
        RECT 688.950 300.450 691.050 301.050 ;
        RECT 670.950 299.400 691.050 300.450 ;
        RECT 670.950 298.950 673.050 299.400 ;
        RECT 688.950 298.950 691.050 299.400 ;
        RECT 700.950 298.950 706.050 301.050 ;
        RECT 769.950 298.950 774.900 301.050 ;
        RECT 776.100 300.450 778.200 300.900 ;
        RECT 781.950 300.450 784.050 301.050 ;
        RECT 802.950 300.450 805.050 301.050 ;
        RECT 776.100 299.400 805.050 300.450 ;
        RECT 226.950 297.450 229.050 298.050 ;
        RECT 284.400 297.450 285.450 298.950 ;
        RECT 776.100 298.800 778.200 299.400 ;
        RECT 781.950 298.950 784.050 299.400 ;
        RECT 802.950 298.950 805.050 299.400 ;
        RECT 844.950 300.450 847.050 301.050 ;
        RECT 853.950 300.450 856.050 301.050 ;
        RECT 844.950 299.400 856.050 300.450 ;
        RECT 844.950 298.950 847.050 299.400 ;
        RECT 853.950 298.950 856.050 299.400 ;
        RECT 226.950 296.400 285.450 297.450 ;
        RECT 370.950 297.450 373.050 298.050 ;
        RECT 376.950 297.450 379.050 298.050 ;
        RECT 370.950 296.400 379.050 297.450 ;
        RECT 226.950 295.950 229.050 296.400 ;
        RECT 370.950 295.950 373.050 296.400 ;
        RECT 376.950 295.950 379.050 296.400 ;
        RECT 427.950 297.450 430.050 298.050 ;
        RECT 466.950 297.450 469.050 298.050 ;
        RECT 427.950 296.400 469.050 297.450 ;
        RECT 427.950 295.950 430.050 296.400 ;
        RECT 466.950 295.950 469.050 296.400 ;
        RECT 472.950 297.450 475.050 298.050 ;
        RECT 496.950 297.450 499.050 298.050 ;
        RECT 472.950 296.400 499.050 297.450 ;
        RECT 472.950 295.950 475.050 296.400 ;
        RECT 496.950 295.950 499.050 296.400 ;
        RECT 556.950 297.450 559.050 298.050 ;
        RECT 598.950 297.450 601.050 298.050 ;
        RECT 556.950 296.400 601.050 297.450 ;
        RECT 556.950 295.950 559.050 296.400 ;
        RECT 598.950 295.950 601.050 296.400 ;
        RECT 640.950 295.950 646.050 298.050 ;
        RECT 55.950 294.450 58.050 295.050 ;
        RECT 67.950 294.450 70.050 295.050 ;
        RECT 55.950 293.400 70.050 294.450 ;
        RECT 55.950 292.950 58.050 293.400 ;
        RECT 67.950 292.950 70.050 293.400 ;
        RECT 82.950 294.450 85.050 295.050 ;
        RECT 88.950 294.450 91.050 295.050 ;
        RECT 82.950 293.400 91.050 294.450 ;
        RECT 82.950 292.950 85.050 293.400 ;
        RECT 88.950 292.950 91.050 293.400 ;
        RECT 253.950 294.450 256.050 295.050 ;
        RECT 310.950 294.450 313.050 295.050 ;
        RECT 346.950 294.450 349.050 295.050 ;
        RECT 253.950 293.400 349.050 294.450 ;
        RECT 253.950 292.950 256.050 293.400 ;
        RECT 310.950 292.950 313.050 293.400 ;
        RECT 346.950 292.950 349.050 293.400 ;
        RECT 373.950 294.450 376.050 295.050 ;
        RECT 421.950 294.450 424.050 295.050 ;
        RECT 373.950 293.400 424.050 294.450 ;
        RECT 373.950 292.950 376.050 293.400 ;
        RECT 421.950 292.950 424.050 293.400 ;
        RECT 439.950 294.450 442.050 295.050 ;
        RECT 469.950 294.450 472.050 295.050 ;
        RECT 439.950 293.400 472.050 294.450 ;
        RECT 439.950 292.950 442.050 293.400 ;
        RECT 469.950 292.950 472.050 293.400 ;
        RECT 475.950 294.450 478.050 295.050 ;
        RECT 496.950 294.450 499.050 295.050 ;
        RECT 475.950 293.400 499.050 294.450 ;
        RECT 475.950 292.950 478.050 293.400 ;
        RECT 496.950 292.950 499.050 293.400 ;
        RECT 517.950 294.450 520.050 295.050 ;
        RECT 550.950 294.450 553.050 295.050 ;
        RECT 517.950 293.400 553.050 294.450 ;
        RECT 517.950 292.950 520.050 293.400 ;
        RECT 550.950 292.950 553.050 293.400 ;
        RECT 574.950 294.450 577.050 295.050 ;
        RECT 616.950 294.450 619.050 294.900 ;
        RECT 574.950 293.400 619.050 294.450 ;
        RECT 574.950 292.950 577.050 293.400 ;
        RECT 616.950 292.800 619.050 293.400 ;
        RECT 640.950 294.450 643.050 295.050 ;
        RECT 658.950 294.450 661.050 295.050 ;
        RECT 640.950 293.400 661.050 294.450 ;
        RECT 664.950 294.450 667.050 298.050 ;
        RECT 679.950 297.450 682.050 298.050 ;
        RECT 727.950 297.450 730.050 298.050 ;
        RECT 754.950 297.450 757.050 298.050 ;
        RECT 679.950 296.400 720.450 297.450 ;
        RECT 679.950 295.950 682.050 296.400 ;
        RECT 719.400 295.050 720.450 296.400 ;
        RECT 727.950 296.400 757.050 297.450 ;
        RECT 727.950 295.950 730.050 296.400 ;
        RECT 754.950 295.950 757.050 296.400 ;
        RECT 832.950 297.450 835.050 298.050 ;
        RECT 841.950 297.450 844.050 298.050 ;
        RECT 832.950 296.400 844.050 297.450 ;
        RECT 832.950 295.950 835.050 296.400 ;
        RECT 841.950 295.950 844.050 296.400 ;
        RECT 847.950 295.950 853.050 298.050 ;
        RECT 718.950 294.450 721.050 295.050 ;
        RECT 844.950 294.450 847.050 295.050 ;
        RECT 852.000 294.900 856.050 295.050 ;
        RECT 664.950 294.000 717.450 294.450 ;
        RECT 665.400 293.400 717.450 294.000 ;
        RECT 640.950 292.950 643.050 293.400 ;
        RECT 658.950 292.950 661.050 293.400 ;
        RECT 34.950 291.450 37.050 292.050 ;
        RECT 100.950 291.450 103.050 292.050 ;
        RECT 105.000 291.450 109.050 292.050 ;
        RECT 34.950 290.400 103.050 291.450 ;
        RECT 104.400 291.000 109.050 291.450 ;
        RECT 34.950 289.950 37.050 290.400 ;
        RECT 100.950 289.950 103.050 290.400 ;
        RECT 103.950 289.950 109.050 291.000 ;
        RECT 268.950 291.450 271.050 292.050 ;
        RECT 334.950 291.450 337.050 292.050 ;
        RECT 268.950 290.400 337.050 291.450 ;
        RECT 268.950 289.950 271.050 290.400 ;
        RECT 334.950 289.950 337.050 290.400 ;
        RECT 403.950 291.450 406.050 292.050 ;
        RECT 436.950 291.450 439.050 292.050 ;
        RECT 403.950 290.400 439.050 291.450 ;
        RECT 403.950 289.950 406.050 290.400 ;
        RECT 436.950 289.950 439.050 290.400 ;
        RECT 448.950 291.450 451.050 292.050 ;
        RECT 484.950 291.450 487.050 292.050 ;
        RECT 448.950 290.400 487.050 291.450 ;
        RECT 448.950 289.950 451.050 290.400 ;
        RECT 484.950 289.950 487.050 290.400 ;
        RECT 490.950 291.450 493.050 292.050 ;
        RECT 601.950 291.450 604.050 292.050 ;
        RECT 661.950 291.450 664.050 292.050 ;
        RECT 490.950 290.400 604.050 291.450 ;
        RECT 490.950 289.950 493.050 290.400 ;
        RECT 601.950 289.950 604.050 290.400 ;
        RECT 608.400 290.400 664.050 291.450 ;
        RECT 716.400 291.450 717.450 293.400 ;
        RECT 718.950 293.400 847.050 294.450 ;
        RECT 718.950 292.950 721.050 293.400 ;
        RECT 844.950 292.950 847.050 293.400 ;
        RECT 850.950 292.950 856.050 294.900 ;
        RECT 850.950 292.800 853.050 292.950 ;
        RECT 733.950 291.450 736.050 292.050 ;
        RECT 716.400 290.400 736.050 291.450 ;
        RECT 13.950 288.450 16.050 289.050 ;
        RECT 49.950 288.450 52.050 289.050 ;
        RECT 79.950 288.450 82.050 289.050 ;
        RECT 13.950 287.400 82.050 288.450 ;
        RECT 13.950 286.950 16.050 287.400 ;
        RECT 49.950 286.950 52.050 287.400 ;
        RECT 79.950 286.950 82.050 287.400 ;
        RECT 85.950 288.450 88.050 289.050 ;
        RECT 97.950 288.450 100.050 289.050 ;
        RECT 85.950 287.400 100.050 288.450 ;
        RECT 85.950 286.950 88.050 287.400 ;
        RECT 97.950 286.950 100.050 287.400 ;
        RECT 103.950 286.950 106.050 289.950 ;
        RECT 109.950 288.450 112.050 289.050 ;
        RECT 232.950 288.450 235.050 289.050 ;
        RECT 109.950 287.400 235.050 288.450 ;
        RECT 109.950 286.950 112.050 287.400 ;
        RECT 232.950 286.950 235.050 287.400 ;
        RECT 307.950 288.450 310.050 289.050 ;
        RECT 316.950 288.450 319.050 289.050 ;
        RECT 439.950 288.450 442.050 289.050 ;
        RECT 307.950 287.400 442.050 288.450 ;
        RECT 307.950 286.950 310.050 287.400 ;
        RECT 316.950 286.950 319.050 287.400 ;
        RECT 439.950 286.950 442.050 287.400 ;
        RECT 454.950 288.450 457.050 289.050 ;
        RECT 502.950 288.450 505.050 289.050 ;
        RECT 454.950 287.400 505.050 288.450 ;
        RECT 454.950 286.950 457.050 287.400 ;
        RECT 502.950 286.950 505.050 287.400 ;
        RECT 511.950 288.450 514.050 289.050 ;
        RECT 608.400 288.450 609.450 290.400 ;
        RECT 661.950 289.950 664.050 290.400 ;
        RECT 733.950 289.950 736.050 290.400 ;
        RECT 745.950 291.450 748.050 292.050 ;
        RECT 793.950 291.450 796.050 292.050 ;
        RECT 745.950 290.400 796.050 291.450 ;
        RECT 745.950 289.950 748.050 290.400 ;
        RECT 793.950 289.950 796.050 290.400 ;
        RECT 511.950 287.400 609.450 288.450 ;
        RECT 682.950 288.450 685.050 289.050 ;
        RECT 715.800 288.450 717.900 289.050 ;
        RECT 682.950 287.400 717.900 288.450 ;
        RECT 511.950 286.950 514.050 287.400 ;
        RECT 682.950 286.950 685.050 287.400 ;
        RECT 715.800 286.950 717.900 287.400 ;
        RECT 719.100 288.450 721.200 289.050 ;
        RECT 760.950 288.450 763.050 289.050 ;
        RECT 719.100 287.400 763.050 288.450 ;
        RECT 719.100 286.950 721.200 287.400 ;
        RECT 760.950 286.950 763.050 287.400 ;
        RECT 814.950 288.450 817.050 289.050 ;
        RECT 841.950 288.450 844.050 289.050 ;
        RECT 814.950 287.400 844.050 288.450 ;
        RECT 814.950 286.950 817.050 287.400 ;
        RECT 841.950 286.950 844.050 287.400 ;
        RECT 43.950 285.450 46.050 286.050 ;
        RECT 61.950 285.450 64.050 286.050 ;
        RECT 94.950 285.450 97.050 286.050 ;
        RECT 112.950 285.450 115.050 286.050 ;
        RECT 43.950 284.400 115.050 285.450 ;
        RECT 43.950 283.950 46.050 284.400 ;
        RECT 61.950 283.950 64.050 284.400 ;
        RECT 94.950 283.950 97.050 284.400 ;
        RECT 112.950 283.950 115.050 284.400 ;
        RECT 178.950 285.450 181.050 286.050 ;
        RECT 193.950 285.450 196.050 286.050 ;
        RECT 178.950 284.400 196.050 285.450 ;
        RECT 178.950 283.950 181.050 284.400 ;
        RECT 193.950 283.950 196.050 284.400 ;
        RECT 289.950 285.450 292.050 286.050 ;
        RECT 307.950 285.450 310.050 286.050 ;
        RECT 289.950 284.400 310.050 285.450 ;
        RECT 289.950 283.950 292.050 284.400 ;
        RECT 307.950 283.950 310.050 284.400 ;
        RECT 322.950 285.450 325.050 286.050 ;
        RECT 337.950 285.450 340.050 286.050 ;
        RECT 322.950 284.400 340.050 285.450 ;
        RECT 322.950 283.950 325.050 284.400 ;
        RECT 337.950 283.950 340.050 284.400 ;
        RECT 343.950 285.450 346.050 286.050 ;
        RECT 352.950 285.450 355.050 286.050 ;
        RECT 343.950 284.400 355.050 285.450 ;
        RECT 343.950 283.950 346.050 284.400 ;
        RECT 352.950 283.950 355.050 284.400 ;
        RECT 457.950 285.450 460.050 286.050 ;
        RECT 478.950 285.450 481.050 286.050 ;
        RECT 457.950 284.400 481.050 285.450 ;
        RECT 457.950 283.950 460.050 284.400 ;
        RECT 478.950 283.950 481.050 284.400 ;
        RECT 484.950 285.450 487.050 286.050 ;
        RECT 526.950 285.450 529.050 286.050 ;
        RECT 484.950 284.400 529.050 285.450 ;
        RECT 484.950 283.950 487.050 284.400 ;
        RECT 526.950 283.950 529.050 284.400 ;
        RECT 532.950 283.950 538.050 286.050 ;
        RECT 556.950 283.950 562.050 286.050 ;
        RECT 583.950 285.450 586.050 286.050 ;
        RECT 721.950 285.450 724.050 286.050 ;
        RECT 583.950 284.400 724.050 285.450 ;
        RECT 583.950 283.950 586.050 284.400 ;
        RECT 721.950 283.950 724.050 284.400 ;
        RECT 733.950 285.450 736.050 286.050 ;
        RECT 769.950 285.450 772.050 286.050 ;
        RECT 733.950 284.400 772.050 285.450 ;
        RECT 733.950 283.950 736.050 284.400 ;
        RECT 769.950 283.950 772.050 284.400 ;
        RECT 799.950 285.450 802.050 286.050 ;
        RECT 853.950 285.450 856.050 286.050 ;
        RECT 799.950 284.400 856.050 285.450 ;
        RECT 799.950 283.950 802.050 284.400 ;
        RECT 853.950 283.950 856.050 284.400 ;
        RECT 70.950 282.450 73.050 283.050 ;
        RECT 97.950 282.450 100.050 283.050 ;
        RECT 118.950 282.450 121.050 283.050 ;
        RECT 70.950 281.400 121.050 282.450 ;
        RECT 70.950 280.950 73.050 281.400 ;
        RECT 97.950 280.950 100.050 281.400 ;
        RECT 118.950 280.950 121.050 281.400 ;
        RECT 133.950 282.450 136.050 283.050 ;
        RECT 169.950 282.450 172.050 283.050 ;
        RECT 133.950 281.400 172.050 282.450 ;
        RECT 133.950 280.950 136.050 281.400 ;
        RECT 169.950 280.950 172.050 281.400 ;
        RECT 259.950 282.450 262.050 283.050 ;
        RECT 292.950 282.450 295.050 283.050 ;
        RECT 259.950 281.400 295.050 282.450 ;
        RECT 259.950 280.950 262.050 281.400 ;
        RECT 292.950 280.950 295.050 281.400 ;
        RECT 298.950 282.450 301.050 283.050 ;
        RECT 415.950 282.450 418.050 283.050 ;
        RECT 298.950 281.400 418.050 282.450 ;
        RECT 298.950 280.950 301.050 281.400 ;
        RECT 415.950 280.950 418.050 281.400 ;
        RECT 469.950 282.450 472.050 283.050 ;
        RECT 511.950 282.450 514.050 283.050 ;
        RECT 469.950 281.400 514.050 282.450 ;
        RECT 469.950 280.950 472.050 281.400 ;
        RECT 511.950 280.950 514.050 281.400 ;
        RECT 520.950 282.450 523.050 283.050 ;
        RECT 529.950 282.450 532.050 283.050 ;
        RECT 520.950 281.400 532.050 282.450 ;
        RECT 520.950 280.950 523.050 281.400 ;
        RECT 529.950 280.950 532.050 281.400 ;
        RECT 550.950 282.450 553.050 283.050 ;
        RECT 556.950 282.450 559.050 283.050 ;
        RECT 550.950 281.400 559.050 282.450 ;
        RECT 550.950 280.950 553.050 281.400 ;
        RECT 556.950 280.950 559.050 281.400 ;
        RECT 604.950 282.450 607.050 283.050 ;
        RECT 622.950 282.450 625.050 283.050 ;
        RECT 604.950 281.400 625.050 282.450 ;
        RECT 604.950 280.950 607.050 281.400 ;
        RECT 622.950 280.950 625.050 281.400 ;
        RECT 661.950 282.450 664.050 283.050 ;
        RECT 700.950 282.450 703.050 283.050 ;
        RECT 736.800 282.450 738.900 283.050 ;
        RECT 661.950 281.400 738.900 282.450 ;
        RECT 661.950 280.950 664.050 281.400 ;
        RECT 700.950 280.950 703.050 281.400 ;
        RECT 736.800 280.950 738.900 281.400 ;
        RECT 740.100 282.450 742.200 283.050 ;
        RECT 766.950 282.450 769.050 283.050 ;
        RECT 740.100 281.400 769.050 282.450 ;
        RECT 740.100 280.950 742.200 281.400 ;
        RECT 766.950 280.950 769.050 281.400 ;
        RECT 790.950 280.950 796.050 283.050 ;
        RECT 820.950 282.450 823.050 283.050 ;
        RECT 826.800 282.450 828.900 283.050 ;
        RECT 820.950 281.400 828.900 282.450 ;
        RECT 820.950 280.950 823.050 281.400 ;
        RECT 826.800 280.950 828.900 281.400 ;
        RECT 830.100 280.950 835.050 283.050 ;
        RECT 13.950 279.450 16.050 280.050 ;
        RECT 43.950 279.450 46.050 280.050 ;
        RECT 73.950 279.450 76.050 280.050 ;
        RECT 136.950 279.450 139.050 280.050 ;
        RECT 13.950 278.400 76.050 279.450 ;
        RECT 13.950 277.950 16.050 278.400 ;
        RECT 43.950 277.950 46.050 278.400 ;
        RECT 73.950 277.950 76.050 278.400 ;
        RECT 92.400 278.400 139.050 279.450 ;
        RECT 10.950 276.450 13.050 277.050 ;
        RECT 22.950 276.450 25.050 277.050 ;
        RECT 10.950 275.400 25.050 276.450 ;
        RECT 10.950 274.950 13.050 275.400 ;
        RECT 22.950 274.950 25.050 275.400 ;
        RECT 49.950 276.450 52.050 277.050 ;
        RECT 64.950 276.450 67.050 277.050 ;
        RECT 49.950 275.400 67.050 276.450 ;
        RECT 49.950 274.950 52.050 275.400 ;
        RECT 64.950 274.950 67.050 275.400 ;
        RECT 70.950 276.450 73.050 277.050 ;
        RECT 92.400 276.450 93.450 278.400 ;
        RECT 136.950 277.950 139.050 278.400 ;
        RECT 226.950 279.450 229.050 280.050 ;
        RECT 262.800 279.450 264.900 280.050 ;
        RECT 226.950 278.400 264.900 279.450 ;
        RECT 226.950 277.950 229.050 278.400 ;
        RECT 262.800 277.950 264.900 278.400 ;
        RECT 266.100 279.450 268.200 280.050 ;
        RECT 271.950 279.450 274.050 280.050 ;
        RECT 266.100 278.400 274.050 279.450 ;
        RECT 266.100 277.950 268.200 278.400 ;
        RECT 271.950 277.950 274.050 278.400 ;
        RECT 322.950 279.450 325.050 280.050 ;
        RECT 361.950 279.450 364.050 280.050 ;
        RECT 388.950 279.450 391.050 280.050 ;
        RECT 322.950 278.400 391.050 279.450 ;
        RECT 322.950 277.950 325.050 278.400 ;
        RECT 361.950 277.950 364.050 278.400 ;
        RECT 388.950 277.950 391.050 278.400 ;
        RECT 424.950 279.450 427.050 280.050 ;
        RECT 466.950 279.450 469.050 280.050 ;
        RECT 490.950 279.450 493.050 280.050 ;
        RECT 424.950 278.400 493.050 279.450 ;
        RECT 424.950 277.950 427.050 278.400 ;
        RECT 466.950 277.950 469.050 278.400 ;
        RECT 490.950 277.950 493.050 278.400 ;
        RECT 508.950 279.450 511.050 280.050 ;
        RECT 565.950 279.450 568.050 280.050 ;
        RECT 508.950 278.400 568.050 279.450 ;
        RECT 508.950 277.950 511.050 278.400 ;
        RECT 565.950 277.950 568.050 278.400 ;
        RECT 694.950 279.450 697.050 280.050 ;
        RECT 703.950 279.450 706.050 280.050 ;
        RECT 694.950 278.400 706.050 279.450 ;
        RECT 694.950 277.950 697.050 278.400 ;
        RECT 703.950 277.950 706.050 278.400 ;
        RECT 70.950 275.400 93.450 276.450 ;
        RECT 136.950 276.450 139.050 277.050 ;
        RECT 154.950 276.450 157.050 277.050 ;
        RECT 136.950 275.400 157.050 276.450 ;
        RECT 70.950 274.950 73.050 275.400 ;
        RECT 28.950 273.450 34.050 274.050 ;
        RECT 20.250 273.000 34.050 273.450 ;
        RECT 19.950 272.400 34.050 273.000 ;
        RECT 19.950 271.050 22.050 272.400 ;
        RECT 28.950 271.950 34.050 272.400 ;
        RECT 43.950 273.450 46.050 274.050 ;
        RECT 43.950 273.000 54.600 273.450 ;
        RECT 43.950 272.400 55.050 273.000 ;
        RECT 43.950 271.950 46.050 272.400 ;
        RECT 52.950 271.050 55.050 272.400 ;
        RECT 13.950 268.950 18.900 271.050 ;
        RECT 19.800 270.000 22.050 271.050 ;
        RECT 23.100 270.450 25.200 271.050 ;
        RECT 28.950 270.450 31.050 271.050 ;
        RECT 19.800 268.950 21.900 270.000 ;
        RECT 23.100 269.400 31.050 270.450 ;
        RECT 23.100 268.950 25.200 269.400 ;
        RECT 28.950 268.950 31.050 269.400 ;
        RECT 10.950 265.950 15.900 268.050 ;
        RECT 16.800 267.000 18.900 268.050 ;
        RECT 20.100 267.450 22.200 268.050 ;
        RECT 28.950 267.450 31.050 268.050 ;
        RECT 34.950 267.450 37.050 271.050 ;
        RECT 49.800 270.000 51.900 271.050 ;
        RECT 52.950 270.000 55.200 271.050 ;
        RECT 49.800 268.950 52.050 270.000 ;
        RECT 53.100 268.950 55.200 270.000 ;
        RECT 58.950 268.950 64.050 271.050 ;
        RECT 73.950 268.950 76.050 274.050 ;
        RECT 91.950 271.950 97.050 274.050 ;
        RECT 103.950 273.450 106.050 274.050 ;
        RECT 103.950 272.400 111.450 273.450 ;
        RECT 103.950 271.950 106.050 272.400 ;
        RECT 110.400 271.050 111.450 272.400 ;
        RECT 112.950 271.950 118.050 274.050 ;
        RECT 136.950 271.950 139.050 275.400 ;
        RECT 154.950 274.950 157.050 275.400 ;
        RECT 145.950 271.950 151.050 274.050 ;
        RECT 253.950 273.450 256.050 277.050 ;
        RECT 239.400 273.000 256.050 273.450 ;
        RECT 238.950 272.400 256.050 273.000 ;
        RECT 79.950 270.450 82.050 271.050 ;
        RECT 88.950 270.450 94.050 271.050 ;
        RECT 79.950 269.400 94.050 270.450 ;
        RECT 79.950 268.950 82.050 269.400 ;
        RECT 88.950 268.950 94.050 269.400 ;
        RECT 97.950 268.950 103.050 271.050 ;
        RECT 110.400 270.450 115.050 271.050 ;
        RECT 104.400 269.400 115.050 270.450 ;
        RECT 20.100 267.000 37.050 267.450 ;
        RECT 16.800 265.950 19.050 267.000 ;
        RECT 20.100 266.400 36.450 267.000 ;
        RECT 20.100 265.950 22.200 266.400 ;
        RECT 28.950 265.950 31.050 266.400 ;
        RECT 49.950 265.950 52.050 268.950 ;
        RECT 10.950 264.450 13.050 265.050 ;
        RECT 16.950 264.450 19.050 265.950 ;
        RECT 10.950 264.000 19.050 264.450 ;
        RECT 55.950 264.450 58.050 268.050 ;
        RECT 64.950 267.450 67.050 268.050 ;
        RECT 70.950 267.450 73.050 268.050 ;
        RECT 64.950 266.400 73.050 267.450 ;
        RECT 64.950 265.950 67.050 266.400 ;
        RECT 70.950 265.950 73.050 266.400 ;
        RECT 70.950 264.450 73.050 265.050 ;
        RECT 55.950 264.000 73.050 264.450 ;
        RECT 10.950 263.400 18.300 264.000 ;
        RECT 56.400 263.400 73.050 264.000 ;
        RECT 10.950 262.950 13.050 263.400 ;
        RECT 70.950 262.950 73.050 263.400 ;
        RECT 76.950 262.950 79.050 268.050 ;
        RECT 85.950 267.450 88.050 268.050 ;
        RECT 104.400 267.450 105.450 269.400 ;
        RECT 111.000 268.950 115.050 269.400 ;
        RECT 85.950 266.400 105.450 267.450 ;
        RECT 85.950 265.950 88.050 266.400 ;
        RECT 118.950 265.950 121.050 271.050 ;
        RECT 133.950 265.950 136.050 271.050 ;
        RECT 139.950 265.950 142.050 271.050 ;
        RECT 151.950 268.950 157.050 271.050 ;
        RECT 160.950 268.050 163.050 271.050 ;
        RECT 172.950 270.450 175.050 271.050 ;
        RECT 178.950 270.450 181.050 271.050 ;
        RECT 172.950 269.400 181.050 270.450 ;
        RECT 172.950 268.950 175.050 269.400 ;
        RECT 178.950 268.950 181.050 269.400 ;
        RECT 184.950 270.450 187.050 271.050 ;
        RECT 196.950 270.450 199.050 271.050 ;
        RECT 201.000 270.450 205.050 271.050 ;
        RECT 184.950 269.400 199.050 270.450 ;
        RECT 184.950 268.950 187.050 269.400 ;
        RECT 196.950 268.950 199.050 269.400 ;
        RECT 200.400 268.950 205.050 270.450 ;
        RECT 208.950 270.450 211.050 271.050 ;
        RECT 217.950 270.450 220.050 271.050 ;
        RECT 208.950 269.400 220.050 270.450 ;
        RECT 208.950 268.950 211.050 269.400 ;
        RECT 217.950 268.950 220.050 269.400 ;
        RECT 238.950 268.950 241.050 272.400 ;
        RECT 253.950 271.950 256.050 272.400 ;
        RECT 259.950 271.950 262.050 277.050 ;
        RECT 349.950 276.450 352.050 277.050 ;
        RECT 439.950 276.450 442.050 277.050 ;
        RECT 472.950 276.450 475.050 277.050 ;
        RECT 349.950 276.000 390.450 276.450 ;
        RECT 349.950 275.400 391.050 276.000 ;
        RECT 349.950 274.950 352.050 275.400 ;
        RECT 280.950 273.450 283.050 274.050 ;
        RECT 292.950 273.450 295.050 274.050 ;
        RECT 280.950 272.400 295.050 273.450 ;
        RECT 280.950 271.950 283.050 272.400 ;
        RECT 292.950 271.950 295.050 272.400 ;
        RECT 298.950 271.050 301.050 274.050 ;
        RECT 370.950 273.450 373.050 274.050 ;
        RECT 382.950 273.450 385.050 274.050 ;
        RECT 370.950 272.400 385.050 273.450 ;
        RECT 370.950 271.950 373.050 272.400 ;
        RECT 382.950 271.950 385.050 272.400 ;
        RECT 388.950 271.950 391.050 275.400 ;
        RECT 439.950 275.400 475.050 276.450 ;
        RECT 439.950 274.950 442.050 275.400 ;
        RECT 472.950 274.950 475.050 275.400 ;
        RECT 394.950 273.450 400.050 274.050 ;
        RECT 424.950 273.450 427.050 274.050 ;
        RECT 394.950 272.400 427.050 273.450 ;
        RECT 394.950 271.950 400.050 272.400 ;
        RECT 424.950 271.950 427.050 272.400 ;
        RECT 430.950 273.450 433.050 274.050 ;
        RECT 436.950 273.450 439.050 274.050 ;
        RECT 430.950 272.400 439.050 273.450 ;
        RECT 430.950 271.950 433.050 272.400 ;
        RECT 436.950 271.950 439.050 272.400 ;
        RECT 448.950 273.450 451.050 274.050 ;
        RECT 457.950 273.450 460.050 274.050 ;
        RECT 448.950 272.400 460.050 273.450 ;
        RECT 448.950 271.950 451.050 272.400 ;
        RECT 457.950 271.950 460.050 272.400 ;
        RECT 463.950 271.050 466.050 271.200 ;
        RECT 244.950 270.450 247.050 271.050 ;
        RECT 256.950 270.450 259.050 271.050 ;
        RECT 244.950 269.400 259.050 270.450 ;
        RECT 244.950 268.950 247.050 269.400 ;
        RECT 256.950 268.950 259.050 269.400 ;
        RECT 268.950 268.950 274.050 271.050 ;
        RECT 289.950 270.450 292.050 271.050 ;
        RECT 295.800 270.450 297.900 271.050 ;
        RECT 289.950 269.400 297.900 270.450 ;
        RECT 298.950 270.000 301.200 271.050 ;
        RECT 289.950 268.950 292.050 269.400 ;
        RECT 295.800 268.950 297.900 269.400 ;
        RECT 299.100 268.950 301.200 270.000 ;
        RECT 310.950 268.950 316.050 271.050 ;
        RECT 319.950 270.450 322.050 271.050 ;
        RECT 328.950 270.450 331.050 271.050 ;
        RECT 319.950 269.400 331.050 270.450 ;
        RECT 319.950 268.950 322.050 269.400 ;
        RECT 328.950 268.950 331.050 269.400 ;
        RECT 148.950 267.450 151.050 268.050 ;
        RECT 157.800 267.450 159.900 268.050 ;
        RECT 148.950 266.400 159.900 267.450 ;
        RECT 160.950 267.000 163.200 268.050 ;
        RECT 148.950 265.950 151.050 266.400 ;
        RECT 157.800 265.950 159.900 266.400 ;
        RECT 161.100 265.950 163.200 267.000 ;
        RECT 166.950 265.950 172.050 268.050 ;
        RECT 130.950 264.450 133.050 265.050 ;
        RECT 139.950 264.450 142.050 265.050 ;
        RECT 160.950 264.450 163.050 265.050 ;
        RECT 130.950 263.400 163.050 264.450 ;
        RECT 130.950 262.950 133.050 263.400 ;
        RECT 139.950 262.950 142.050 263.400 ;
        RECT 160.950 262.950 163.050 263.400 ;
        RECT 175.950 262.950 178.050 268.050 ;
        RECT 181.950 267.450 184.050 268.050 ;
        RECT 190.950 267.450 193.050 268.050 ;
        RECT 200.400 267.450 201.450 268.950 ;
        RECT 181.950 266.400 189.450 267.450 ;
        RECT 181.950 265.950 184.050 266.400 ;
        RECT 188.400 264.450 189.450 266.400 ;
        RECT 190.950 266.400 201.450 267.450 ;
        RECT 190.950 265.950 193.050 266.400 ;
        RECT 202.950 265.950 208.050 268.050 ;
        RECT 229.950 265.950 235.050 268.050 ;
        RECT 244.950 267.450 247.050 268.050 ;
        RECT 259.950 267.450 262.050 268.050 ;
        RECT 244.950 266.400 262.050 267.450 ;
        RECT 244.950 265.950 247.050 266.400 ;
        RECT 259.950 265.950 262.050 266.400 ;
        RECT 280.950 265.050 283.050 268.050 ;
        RECT 298.950 267.450 301.050 268.050 ;
        RECT 316.950 267.450 319.050 268.050 ;
        RECT 298.950 266.400 319.050 267.450 ;
        RECT 298.950 265.950 301.050 266.400 ;
        RECT 316.950 265.950 319.050 266.400 ;
        RECT 322.950 265.950 328.050 268.050 ;
        RECT 334.950 265.950 337.050 271.050 ;
        RECT 343.950 270.450 346.050 271.050 ;
        RECT 352.950 270.450 355.050 271.050 ;
        RECT 343.950 269.400 355.050 270.450 ;
        RECT 343.950 268.950 346.050 269.400 ;
        RECT 352.950 268.950 355.050 269.400 ;
        RECT 358.950 268.950 364.050 271.050 ;
        RECT 340.950 267.450 343.050 268.050 ;
        RECT 346.950 267.450 349.050 268.050 ;
        RECT 352.800 267.450 354.900 268.050 ;
        RECT 340.950 266.400 354.900 267.450 ;
        RECT 340.950 265.950 343.050 266.400 ;
        RECT 346.950 265.950 349.050 266.400 ;
        RECT 352.800 265.950 354.900 266.400 ;
        RECT 355.800 267.000 357.900 268.050 ;
        RECT 359.100 267.450 361.200 268.050 ;
        RECT 370.950 267.450 373.050 268.050 ;
        RECT 355.800 265.950 358.050 267.000 ;
        RECT 359.100 266.400 373.050 267.450 ;
        RECT 359.100 265.950 361.200 266.400 ;
        RECT 370.950 265.950 373.050 266.400 ;
        RECT 376.950 265.950 379.050 271.050 ;
        RECT 388.950 268.950 394.050 271.050 ;
        RECT 382.950 267.450 385.050 268.050 ;
        RECT 409.950 267.450 412.050 271.050 ;
        RECT 418.950 270.450 421.050 271.050 ;
        RECT 427.800 270.450 429.900 271.050 ;
        RECT 418.950 269.400 429.900 270.450 ;
        RECT 418.950 268.950 421.050 269.400 ;
        RECT 427.800 268.950 429.900 269.400 ;
        RECT 431.100 270.450 433.200 271.050 ;
        RECT 442.950 270.450 448.050 271.050 ;
        RECT 431.100 269.400 448.050 270.450 ;
        RECT 431.100 268.950 433.200 269.400 ;
        RECT 442.950 268.950 448.050 269.400 ;
        RECT 451.950 268.950 457.050 271.050 ;
        RECT 463.950 269.100 469.050 271.050 ;
        RECT 465.000 268.950 469.050 269.100 ;
        RECT 472.950 268.950 475.050 274.050 ;
        RECT 478.800 273.000 480.900 274.050 ;
        RECT 478.800 271.950 481.050 273.000 ;
        RECT 482.100 271.950 487.050 274.050 ;
        RECT 490.950 271.950 493.050 277.050 ;
        RECT 544.950 276.450 547.050 277.050 ;
        RECT 553.950 276.450 556.050 277.050 ;
        RECT 583.800 276.450 585.900 277.050 ;
        RECT 544.950 275.400 556.050 276.450 ;
        RECT 544.950 274.950 547.050 275.400 ;
        RECT 553.950 274.950 556.050 275.400 ;
        RECT 557.400 275.400 585.900 276.450 ;
        RECT 499.950 273.450 502.050 274.050 ;
        RECT 514.950 273.450 517.050 274.050 ;
        RECT 499.950 272.400 517.050 273.450 ;
        RECT 499.950 271.950 502.050 272.400 ;
        RECT 514.950 271.950 517.050 272.400 ;
        RECT 523.950 273.450 526.050 274.050 ;
        RECT 535.950 273.450 538.050 274.050 ;
        RECT 550.950 273.450 553.050 274.050 ;
        RECT 557.400 273.450 558.450 275.400 ;
        RECT 583.800 274.950 585.900 275.400 ;
        RECT 613.950 276.450 616.050 277.050 ;
        RECT 640.950 276.450 643.050 277.050 ;
        RECT 613.950 275.400 643.050 276.450 ;
        RECT 613.950 274.950 616.050 275.400 ;
        RECT 640.950 274.950 643.050 275.400 ;
        RECT 685.950 276.450 688.050 277.050 ;
        RECT 718.950 276.450 721.050 277.200 ;
        RECT 685.950 275.400 721.050 276.450 ;
        RECT 685.950 274.950 688.050 275.400 ;
        RECT 718.950 275.100 721.050 275.400 ;
        RECT 736.950 276.450 739.050 277.050 ;
        RECT 751.950 276.450 754.050 277.050 ;
        RECT 736.950 275.400 754.050 276.450 ;
        RECT 736.950 274.950 739.050 275.400 ;
        RECT 751.950 274.950 754.050 275.400 ;
        RECT 523.950 273.000 549.300 273.450 ;
        RECT 523.950 272.400 550.050 273.000 ;
        RECT 523.950 271.950 526.050 272.400 ;
        RECT 535.950 271.950 538.050 272.400 ;
        RECT 478.950 270.450 481.050 271.950 ;
        RECT 547.950 271.050 550.050 272.400 ;
        RECT 550.950 272.400 558.450 273.450 ;
        RECT 571.950 273.450 574.050 274.050 ;
        RECT 580.950 273.450 583.050 274.050 ;
        RECT 571.950 272.400 583.050 273.450 ;
        RECT 550.950 271.950 553.050 272.400 ;
        RECT 571.950 271.950 574.050 272.400 ;
        RECT 580.950 271.950 583.050 272.400 ;
        RECT 584.250 271.050 585.300 274.950 ;
        RECT 769.950 274.050 772.050 274.200 ;
        RECT 619.950 273.450 622.050 274.050 ;
        RECT 634.950 273.450 637.050 274.050 ;
        RECT 608.400 273.000 622.050 273.450 ;
        RECT 629.400 273.000 637.050 273.450 ;
        RECT 607.950 272.400 622.050 273.000 ;
        RECT 478.950 270.000 483.450 270.450 ;
        RECT 479.250 269.400 483.450 270.000 ;
        RECT 382.950 267.000 412.050 267.450 ;
        RECT 382.950 266.400 411.450 267.000 ;
        RECT 382.950 265.950 385.050 266.400 ;
        RECT 433.950 265.950 439.050 268.050 ;
        RECT 442.950 265.950 448.050 268.050 ;
        RECT 457.950 267.450 460.050 268.050 ;
        RECT 463.950 267.450 466.050 268.050 ;
        RECT 468.000 267.450 472.050 268.050 ;
        RECT 457.950 266.400 466.050 267.450 ;
        RECT 457.950 265.950 460.050 266.400 ;
        RECT 193.950 264.450 196.050 265.050 ;
        RECT 188.400 263.400 196.050 264.450 ;
        RECT 193.950 262.950 196.050 263.400 ;
        RECT 223.950 264.450 226.050 265.050 ;
        RECT 229.950 264.450 232.050 265.050 ;
        RECT 223.950 263.400 232.050 264.450 ;
        RECT 223.950 262.950 226.050 263.400 ;
        RECT 229.950 262.950 232.050 263.400 ;
        RECT 280.800 264.000 283.050 265.050 ;
        RECT 284.100 264.450 286.200 265.050 ;
        RECT 299.400 264.450 300.450 265.950 ;
        RECT 337.950 264.450 340.050 265.050 ;
        RECT 280.800 262.950 282.900 264.000 ;
        RECT 284.100 263.400 300.450 264.450 ;
        RECT 302.400 263.400 340.050 264.450 ;
        RECT 284.100 262.950 286.200 263.400 ;
        RECT 61.950 261.450 64.050 262.050 ;
        RECT 85.950 261.450 88.050 262.050 ;
        RECT 61.950 260.400 88.050 261.450 ;
        RECT 61.950 259.950 64.050 260.400 ;
        RECT 85.950 259.950 88.050 260.400 ;
        RECT 106.950 261.450 109.050 262.050 ;
        RECT 133.950 261.450 136.050 262.050 ;
        RECT 148.800 261.450 150.900 262.050 ;
        RECT 106.950 260.400 150.900 261.450 ;
        RECT 106.950 259.950 109.050 260.400 ;
        RECT 133.950 259.950 136.050 260.400 ;
        RECT 148.800 259.950 150.900 260.400 ;
        RECT 152.100 261.450 154.200 262.050 ;
        RECT 169.950 261.450 172.050 262.050 ;
        RECT 152.100 260.400 172.050 261.450 ;
        RECT 152.100 259.950 154.200 260.400 ;
        RECT 169.950 259.950 172.050 260.400 ;
        RECT 259.950 261.450 262.050 262.050 ;
        RECT 265.950 261.450 268.050 262.050 ;
        RECT 259.950 260.400 268.050 261.450 ;
        RECT 259.950 259.950 262.050 260.400 ;
        RECT 265.950 259.950 268.050 260.400 ;
        RECT 280.950 261.450 283.050 262.050 ;
        RECT 302.400 261.450 303.450 263.400 ;
        RECT 337.950 262.950 340.050 263.400 ;
        RECT 355.950 262.950 358.050 265.950 ;
        RECT 463.950 265.800 466.050 266.400 ;
        RECT 467.400 265.950 472.050 267.450 ;
        RECT 475.950 265.950 481.050 268.050 ;
        RECT 373.950 264.450 376.050 265.050 ;
        RECT 388.950 264.450 391.050 265.050 ;
        RECT 373.950 263.400 391.050 264.450 ;
        RECT 373.950 262.950 376.050 263.400 ;
        RECT 388.950 262.950 391.050 263.400 ;
        RECT 412.950 264.450 415.050 265.050 ;
        RECT 418.950 264.450 421.050 265.050 ;
        RECT 412.950 263.400 421.050 264.450 ;
        RECT 412.950 262.950 415.050 263.400 ;
        RECT 418.950 262.950 421.050 263.400 ;
        RECT 427.950 264.450 430.050 265.050 ;
        RECT 439.950 264.450 442.050 265.050 ;
        RECT 427.950 263.400 442.050 264.450 ;
        RECT 427.950 262.950 430.050 263.400 ;
        RECT 439.950 262.950 442.050 263.400 ;
        RECT 448.950 262.950 453.900 265.050 ;
        RECT 455.100 264.450 457.200 265.050 ;
        RECT 467.400 264.450 468.450 265.950 ;
        RECT 455.100 263.400 468.450 264.450 ;
        RECT 482.400 264.450 483.450 269.400 ;
        RECT 484.950 268.950 490.050 271.050 ;
        RECT 535.950 270.450 538.050 271.050 ;
        RECT 541.950 270.450 544.050 271.050 ;
        RECT 535.950 269.400 544.050 270.450 ;
        RECT 535.950 268.950 538.050 269.400 ;
        RECT 541.950 268.950 544.050 269.400 ;
        RECT 547.800 270.000 550.050 271.050 ;
        RECT 551.100 270.000 553.200 271.050 ;
        RECT 547.800 268.950 549.900 270.000 ;
        RECT 550.950 268.950 553.200 270.000 ;
        RECT 556.950 270.450 559.050 271.050 ;
        RECT 565.800 270.450 567.900 271.050 ;
        RECT 556.950 269.400 567.900 270.450 ;
        RECT 556.950 268.950 559.050 269.400 ;
        RECT 565.800 268.950 567.900 269.400 ;
        RECT 569.100 268.950 574.050 271.050 ;
        RECT 583.800 268.950 585.900 271.050 ;
        RECT 587.100 268.950 592.050 271.050 ;
        RECT 607.950 268.950 610.050 272.400 ;
        RECT 619.950 271.950 622.050 272.400 ;
        RECT 628.950 272.400 637.050 273.000 ;
        RECT 511.950 268.050 514.050 268.200 ;
        RECT 508.950 266.100 514.050 268.050 ;
        RECT 544.950 267.450 549.000 268.050 ;
        RECT 508.950 265.950 513.000 266.100 ;
        RECT 544.950 265.950 549.450 267.450 ;
        RECT 550.950 265.950 553.050 268.950 ;
        RECT 613.950 268.050 616.050 271.050 ;
        RECT 628.950 270.450 631.050 272.400 ;
        RECT 634.950 271.950 637.050 272.400 ;
        RECT 673.950 273.450 676.050 274.050 ;
        RECT 688.950 273.450 691.050 274.050 ;
        RECT 718.950 273.450 721.050 273.900 ;
        RECT 673.950 273.000 687.450 273.450 ;
        RECT 673.950 272.400 688.050 273.000 ;
        RECT 673.950 271.950 676.050 272.400 ;
        RECT 617.250 270.000 631.050 270.450 ;
        RECT 616.950 269.400 631.050 270.000 ;
        RECT 616.950 268.050 619.050 269.400 ;
        RECT 628.950 268.950 631.050 269.400 ;
        RECT 634.950 268.050 637.050 271.050 ;
        RECT 649.950 268.950 655.050 271.050 ;
        RECT 658.950 268.950 664.050 271.050 ;
        RECT 676.950 268.950 682.050 271.050 ;
        RECT 685.950 270.450 688.050 272.400 ;
        RECT 688.950 272.400 721.050 273.450 ;
        RECT 688.950 271.950 691.050 272.400 ;
        RECT 697.950 271.050 700.050 272.400 ;
        RECT 718.950 271.800 721.050 272.400 ;
        RECT 739.950 273.450 742.050 274.050 ;
        RECT 751.950 273.450 754.050 274.050 ;
        RECT 739.950 272.400 754.050 273.450 ;
        RECT 739.950 271.950 742.050 272.400 ;
        RECT 751.950 271.950 754.050 272.400 ;
        RECT 685.950 269.400 696.450 270.450 ;
        RECT 685.950 268.950 688.050 269.400 ;
        RECT 559.950 265.950 564.900 268.050 ;
        RECT 566.100 265.950 571.050 268.050 ;
        RECT 505.950 264.450 508.050 265.050 ;
        RECT 482.400 263.400 508.050 264.450 ;
        RECT 455.100 262.950 457.200 263.400 ;
        RECT 505.950 262.950 508.050 263.400 ;
        RECT 517.950 264.450 520.050 265.200 ;
        RECT 523.950 264.450 526.050 265.050 ;
        RECT 517.950 263.400 526.050 264.450 ;
        RECT 548.400 264.450 549.450 265.950 ;
        RECT 548.400 263.400 573.450 264.450 ;
        RECT 517.950 263.100 520.050 263.400 ;
        RECT 523.950 262.950 526.050 263.400 ;
        RECT 280.950 260.400 303.450 261.450 ;
        RECT 409.950 261.450 412.050 262.050 ;
        RECT 418.950 261.450 421.050 262.050 ;
        RECT 409.950 260.400 421.050 261.450 ;
        RECT 280.950 259.950 283.050 260.400 ;
        RECT 409.950 259.950 412.050 260.400 ;
        RECT 418.950 259.950 421.050 260.400 ;
        RECT 514.950 261.900 519.000 262.050 ;
        RECT 514.950 259.950 520.050 261.900 ;
        RECT 535.950 261.450 538.050 262.050 ;
        RECT 556.950 261.450 559.050 262.050 ;
        RECT 535.950 260.400 559.050 261.450 ;
        RECT 572.400 261.450 573.450 263.400 ;
        RECT 574.950 262.950 577.050 268.050 ;
        RECT 583.950 265.950 589.050 268.050 ;
        RECT 595.950 267.450 598.050 268.050 ;
        RECT 604.950 267.450 607.050 268.050 ;
        RECT 610.800 267.450 612.900 268.050 ;
        RECT 595.950 266.400 603.450 267.450 ;
        RECT 595.950 265.950 598.050 266.400 ;
        RECT 602.400 264.450 603.450 266.400 ;
        RECT 604.950 266.400 612.900 267.450 ;
        RECT 604.950 265.950 607.050 266.400 ;
        RECT 610.800 265.950 612.900 266.400 ;
        RECT 613.800 267.000 616.050 268.050 ;
        RECT 616.800 267.000 619.050 268.050 ;
        RECT 620.100 267.450 622.200 268.050 ;
        RECT 631.800 267.450 633.900 268.050 ;
        RECT 613.800 265.950 615.900 267.000 ;
        RECT 616.800 265.950 618.900 267.000 ;
        RECT 620.100 266.400 633.900 267.450 ;
        RECT 620.100 265.950 622.200 266.400 ;
        RECT 631.800 265.950 633.900 266.400 ;
        RECT 634.800 267.000 637.050 268.050 ;
        RECT 638.100 267.450 640.200 268.050 ;
        RECT 655.950 267.450 658.050 268.050 ;
        RECT 634.800 265.950 636.900 267.000 ;
        RECT 638.100 266.400 658.050 267.450 ;
        RECT 638.100 265.950 640.200 266.400 ;
        RECT 655.950 265.950 658.050 266.400 ;
        RECT 664.950 267.450 667.050 268.050 ;
        RECT 670.800 267.450 672.900 268.050 ;
        RECT 664.950 266.400 672.900 267.450 ;
        RECT 664.950 265.950 667.050 266.400 ;
        RECT 670.800 265.950 672.900 266.400 ;
        RECT 674.100 267.450 676.200 268.050 ;
        RECT 682.950 267.450 685.050 268.050 ;
        RECT 674.100 266.400 685.050 267.450 ;
        RECT 674.100 265.950 676.200 266.400 ;
        RECT 682.950 265.950 685.050 266.400 ;
        RECT 688.950 265.950 694.050 268.050 ;
        RECT 695.400 267.450 696.450 269.400 ;
        RECT 697.800 270.000 700.050 271.050 ;
        RECT 697.800 268.950 699.900 270.000 ;
        RECT 701.100 268.950 706.050 271.050 ;
        RECT 736.950 268.950 742.050 271.050 ;
        RECT 745.950 268.950 751.050 271.050 ;
        RECT 757.950 268.950 760.050 274.050 ;
        RECT 763.950 268.950 766.050 274.050 ;
        RECT 769.950 272.100 775.050 274.050 ;
        RECT 771.000 271.950 775.050 272.100 ;
        RECT 784.950 273.450 787.050 274.050 ;
        RECT 790.800 273.450 792.900 274.050 ;
        RECT 784.950 272.400 792.900 273.450 ;
        RECT 784.950 271.950 787.050 272.400 ;
        RECT 790.800 271.950 792.900 272.400 ;
        RECT 794.100 273.450 796.200 274.050 ;
        RECT 838.950 273.450 843.000 274.050 ;
        RECT 850.950 273.450 853.050 274.050 ;
        RECT 794.100 273.000 837.450 273.450 ;
        RECT 794.100 272.400 838.050 273.000 ;
        RECT 794.100 271.950 796.200 272.400 ;
        RECT 769.950 270.450 772.050 270.900 ;
        RECT 769.950 270.000 786.450 270.450 ;
        RECT 769.950 269.400 787.050 270.000 ;
        RECT 769.950 268.800 772.050 269.400 ;
        RECT 784.950 268.050 787.050 269.400 ;
        RECT 835.950 268.950 838.050 272.400 ;
        RECT 838.950 272.400 853.050 273.450 ;
        RECT 838.950 271.950 844.050 272.400 ;
        RECT 850.950 271.950 853.050 272.400 ;
        RECT 841.950 268.950 844.050 271.950 ;
        RECT 700.950 267.450 703.050 268.050 ;
        RECT 695.400 266.400 703.050 267.450 ;
        RECT 700.950 265.950 703.050 266.400 ;
        RECT 709.950 265.950 714.900 268.050 ;
        RECT 722.100 265.950 727.050 268.050 ;
        RECT 613.950 264.450 616.050 265.050 ;
        RECT 634.950 264.450 637.050 265.050 ;
        RECT 646.950 264.450 649.050 265.050 ;
        RECT 602.400 263.400 649.050 264.450 ;
        RECT 613.950 262.950 616.050 263.400 ;
        RECT 634.950 262.950 637.050 263.400 ;
        RECT 646.950 262.950 649.050 263.400 ;
        RECT 652.950 264.450 655.050 265.050 ;
        RECT 661.950 264.450 664.050 265.050 ;
        RECT 652.950 263.400 664.050 264.450 ;
        RECT 652.950 262.950 655.050 263.400 ;
        RECT 661.950 262.950 664.050 263.400 ;
        RECT 694.950 264.450 697.050 265.050 ;
        RECT 700.950 264.450 703.050 265.050 ;
        RECT 694.950 263.400 703.050 264.450 ;
        RECT 694.950 262.950 697.050 263.400 ;
        RECT 700.950 262.950 703.050 263.400 ;
        RECT 736.950 262.950 739.050 268.050 ;
        RECT 742.950 267.450 745.050 268.050 ;
        RECT 751.950 267.450 754.050 268.050 ;
        RECT 760.800 267.450 762.900 268.050 ;
        RECT 765.000 267.900 769.050 268.050 ;
        RECT 742.950 266.400 750.450 267.450 ;
        RECT 742.950 265.950 745.050 266.400 ;
        RECT 749.400 264.450 750.450 266.400 ;
        RECT 751.950 266.400 762.900 267.450 ;
        RECT 751.950 265.950 754.050 266.400 ;
        RECT 760.800 265.950 762.900 266.400 ;
        RECT 764.100 265.950 769.050 267.900 ;
        RECT 784.950 267.000 787.200 268.050 ;
        RECT 785.100 265.950 787.200 267.000 ;
        RECT 793.950 267.450 796.050 268.050 ;
        RECT 799.950 267.450 802.050 268.050 ;
        RECT 793.950 266.400 802.050 267.450 ;
        RECT 793.950 265.950 796.050 266.400 ;
        RECT 799.950 265.950 802.050 266.400 ;
        RECT 805.950 267.450 808.050 268.050 ;
        RECT 814.950 267.450 817.050 268.050 ;
        RECT 805.950 266.400 817.050 267.450 ;
        RECT 805.950 265.950 808.050 266.400 ;
        RECT 814.950 265.950 817.050 266.400 ;
        RECT 764.100 265.800 766.200 265.950 ;
        RECT 760.950 264.450 763.050 265.050 ;
        RECT 749.400 263.400 763.050 264.450 ;
        RECT 760.950 262.950 763.050 263.400 ;
        RECT 589.950 261.450 592.050 262.200 ;
        RECT 572.400 260.400 592.050 261.450 ;
        RECT 535.950 259.950 538.050 260.400 ;
        RECT 556.950 259.950 559.050 260.400 ;
        RECT 589.950 260.100 592.050 260.400 ;
        RECT 676.950 261.450 679.050 262.050 ;
        RECT 757.950 261.450 760.050 262.050 ;
        RECT 769.800 261.450 771.900 262.050 ;
        RECT 676.950 260.400 693.450 261.450 ;
        RECT 676.950 259.950 679.050 260.400 ;
        RECT 517.950 259.800 520.050 259.950 ;
        RECT 55.950 258.450 58.050 259.050 ;
        RECT 103.950 258.450 106.050 259.050 ;
        RECT 55.950 257.400 106.050 258.450 ;
        RECT 55.950 256.950 58.050 257.400 ;
        RECT 103.950 256.950 106.050 257.400 ;
        RECT 127.950 258.450 130.050 259.050 ;
        RECT 175.950 258.450 178.050 259.050 ;
        RECT 223.950 258.450 226.050 259.050 ;
        RECT 229.950 258.450 232.050 259.050 ;
        RECT 289.950 258.450 292.050 259.050 ;
        RECT 127.950 257.400 138.450 258.450 ;
        RECT 127.950 256.950 130.050 257.400 ;
        RECT 61.950 255.450 64.050 256.050 ;
        RECT 85.950 255.450 88.050 256.050 ;
        RECT 61.950 254.400 88.050 255.450 ;
        RECT 137.400 255.450 138.450 257.400 ;
        RECT 175.950 257.400 292.050 258.450 ;
        RECT 175.950 256.950 178.050 257.400 ;
        RECT 223.950 256.950 226.050 257.400 ;
        RECT 229.950 256.950 232.050 257.400 ;
        RECT 289.950 256.950 292.050 257.400 ;
        RECT 307.950 256.950 313.050 259.050 ;
        RECT 457.950 258.450 460.050 259.050 ;
        RECT 526.950 258.450 529.050 259.050 ;
        RECT 457.950 257.400 529.050 258.450 ;
        RECT 457.950 256.950 460.050 257.400 ;
        RECT 526.950 256.950 529.050 257.400 ;
        RECT 532.950 258.450 535.050 259.050 ;
        RECT 589.950 258.450 592.050 258.900 ;
        RECT 532.950 257.400 592.050 258.450 ;
        RECT 532.950 256.950 535.050 257.400 ;
        RECT 589.950 256.800 592.050 257.400 ;
        RECT 598.950 258.450 601.050 259.050 ;
        RECT 619.950 258.450 622.050 259.050 ;
        RECT 598.950 257.400 622.050 258.450 ;
        RECT 598.950 256.950 601.050 257.400 ;
        RECT 619.950 256.950 622.050 257.400 ;
        RECT 679.950 258.450 682.050 259.050 ;
        RECT 688.950 258.450 691.050 259.050 ;
        RECT 679.950 257.400 691.050 258.450 ;
        RECT 692.400 258.450 693.450 260.400 ;
        RECT 757.950 260.400 771.900 261.450 ;
        RECT 757.950 259.950 760.050 260.400 ;
        RECT 769.800 259.950 771.900 260.400 ;
        RECT 773.100 261.450 775.200 262.200 ;
        RECT 790.950 261.450 793.050 262.050 ;
        RECT 773.100 260.400 793.050 261.450 ;
        RECT 773.100 260.100 775.200 260.400 ;
        RECT 790.950 259.950 793.050 260.400 ;
        RECT 802.950 259.950 805.050 265.050 ;
        RECT 838.950 262.950 841.050 268.050 ;
        RECT 844.950 262.950 847.050 268.050 ;
        RECT 850.950 262.950 853.050 268.050 ;
        RECT 811.950 261.450 814.050 262.050 ;
        RECT 817.950 261.450 820.050 262.050 ;
        RECT 811.950 260.400 820.050 261.450 ;
        RECT 811.950 259.950 814.050 260.400 ;
        RECT 817.950 259.950 820.050 260.400 ;
        RECT 829.950 261.450 832.050 262.050 ;
        RECT 853.950 261.450 856.050 262.200 ;
        RECT 829.950 260.400 856.050 261.450 ;
        RECT 829.950 259.950 832.050 260.400 ;
        RECT 853.950 260.100 856.050 260.400 ;
        RECT 706.950 258.450 709.050 259.200 ;
        RECT 715.950 258.450 718.050 259.050 ;
        RECT 692.400 257.400 699.450 258.450 ;
        RECT 679.950 256.950 682.050 257.400 ;
        RECT 688.950 256.950 691.050 257.400 ;
        RECT 157.950 255.450 160.050 256.050 ;
        RECT 137.400 254.400 160.050 255.450 ;
        RECT 61.950 253.950 64.050 254.400 ;
        RECT 85.950 253.950 88.050 254.400 ;
        RECT 157.950 253.950 160.050 254.400 ;
        RECT 178.950 255.450 181.050 256.050 ;
        RECT 184.950 255.450 187.050 256.050 ;
        RECT 178.950 254.400 187.050 255.450 ;
        RECT 178.950 253.950 181.050 254.400 ;
        RECT 184.950 253.950 187.050 254.400 ;
        RECT 205.950 255.450 208.050 256.050 ;
        RECT 244.950 255.450 247.050 256.050 ;
        RECT 205.950 254.400 247.050 255.450 ;
        RECT 205.950 253.950 208.050 254.400 ;
        RECT 244.950 253.950 247.050 254.400 ;
        RECT 364.950 255.450 367.050 256.050 ;
        RECT 436.950 255.450 439.050 256.200 ;
        RECT 364.950 254.400 439.050 255.450 ;
        RECT 364.950 253.950 367.050 254.400 ;
        RECT 436.950 254.100 439.050 254.400 ;
        RECT 502.950 255.450 505.050 256.050 ;
        RECT 565.950 255.450 568.050 256.050 ;
        RECT 604.950 255.450 607.050 256.050 ;
        RECT 502.950 254.400 531.450 255.450 ;
        RECT 502.950 253.950 505.050 254.400 ;
        RECT 52.950 252.450 55.050 253.050 ;
        RECT 82.950 252.450 85.050 253.050 ;
        RECT 52.950 251.400 85.050 252.450 ;
        RECT 52.950 250.950 55.050 251.400 ;
        RECT 82.950 250.950 85.050 251.400 ;
        RECT 145.950 252.450 148.050 253.050 ;
        RECT 202.950 252.450 205.050 253.050 ;
        RECT 241.950 252.450 244.050 253.050 ;
        RECT 283.950 252.450 286.050 253.050 ;
        RECT 145.950 251.400 286.050 252.450 ;
        RECT 145.950 250.950 148.050 251.400 ;
        RECT 202.950 250.950 205.050 251.400 ;
        RECT 241.950 250.950 244.050 251.400 ;
        RECT 283.950 250.950 286.050 251.400 ;
        RECT 307.950 252.450 310.050 253.050 ;
        RECT 403.950 252.450 406.050 253.050 ;
        RECT 307.950 251.400 406.050 252.450 ;
        RECT 307.950 250.950 310.050 251.400 ;
        RECT 403.950 250.950 406.050 251.400 ;
        RECT 412.950 252.450 415.050 253.050 ;
        RECT 436.950 252.450 439.050 252.900 ;
        RECT 412.950 251.400 439.050 252.450 ;
        RECT 412.950 250.950 415.050 251.400 ;
        RECT 436.950 250.800 439.050 251.400 ;
        RECT 442.950 252.450 445.050 253.050 ;
        RECT 484.950 252.450 487.050 253.050 ;
        RECT 442.950 251.400 487.050 252.450 ;
        RECT 530.400 252.450 531.450 254.400 ;
        RECT 565.950 254.400 607.050 255.450 ;
        RECT 565.950 253.950 568.050 254.400 ;
        RECT 604.950 253.950 607.050 254.400 ;
        RECT 655.950 255.450 658.050 256.050 ;
        RECT 691.950 255.450 694.050 256.050 ;
        RECT 655.950 254.400 694.050 255.450 ;
        RECT 698.400 255.450 699.450 257.400 ;
        RECT 706.950 257.400 718.050 258.450 ;
        RECT 706.950 257.100 709.050 257.400 ;
        RECT 715.950 256.950 718.050 257.400 ;
        RECT 742.950 258.450 745.050 259.050 ;
        RECT 774.000 258.900 778.050 259.050 ;
        RECT 742.950 257.400 753.450 258.450 ;
        RECT 742.950 256.950 745.050 257.400 ;
        RECT 706.950 255.450 709.050 255.900 ;
        RECT 748.950 255.450 751.050 256.050 ;
        RECT 698.400 254.400 751.050 255.450 ;
        RECT 752.400 255.450 753.450 257.400 ;
        RECT 772.950 256.950 778.050 258.900 ;
        RECT 781.950 258.450 784.050 259.050 ;
        RECT 790.800 258.450 792.900 259.050 ;
        RECT 781.950 257.400 792.900 258.450 ;
        RECT 781.950 256.950 784.050 257.400 ;
        RECT 790.800 256.950 792.900 257.400 ;
        RECT 794.100 256.950 799.050 259.050 ;
        RECT 829.950 256.950 835.050 259.050 ;
        RECT 850.950 258.900 855.000 259.050 ;
        RECT 850.950 256.950 856.050 258.900 ;
        RECT 772.950 256.800 775.050 256.950 ;
        RECT 853.950 256.800 856.050 256.950 ;
        RECT 802.950 255.450 805.050 256.050 ;
        RECT 811.800 255.450 813.900 256.050 ;
        RECT 752.400 254.400 813.900 255.450 ;
        RECT 655.950 253.950 658.050 254.400 ;
        RECT 691.950 253.950 694.050 254.400 ;
        RECT 706.950 253.800 709.050 254.400 ;
        RECT 748.950 253.950 751.050 254.400 ;
        RECT 802.950 253.950 805.050 254.400 ;
        RECT 811.800 253.950 813.900 254.400 ;
        RECT 815.100 255.450 817.200 256.200 ;
        RECT 826.950 255.450 829.050 256.050 ;
        RECT 844.950 255.450 847.050 256.050 ;
        RECT 815.100 254.400 847.050 255.450 ;
        RECT 815.100 254.100 817.200 254.400 ;
        RECT 826.950 253.950 829.050 254.400 ;
        RECT 844.950 253.950 847.050 254.400 ;
        RECT 547.950 252.450 550.050 253.050 ;
        RECT 530.400 251.400 550.050 252.450 ;
        RECT 442.950 250.950 445.050 251.400 ;
        RECT 484.950 250.950 487.050 251.400 ;
        RECT 547.950 250.950 550.050 251.400 ;
        RECT 568.950 252.450 571.050 253.050 ;
        RECT 592.950 252.450 595.050 253.050 ;
        RECT 568.950 251.400 595.050 252.450 ;
        RECT 568.950 250.950 571.050 251.400 ;
        RECT 592.950 250.950 595.050 251.400 ;
        RECT 673.950 252.450 676.050 253.050 ;
        RECT 694.950 252.450 697.050 253.200 ;
        RECT 673.950 251.400 697.050 252.450 ;
        RECT 673.950 250.950 676.050 251.400 ;
        RECT 694.950 251.100 697.050 251.400 ;
        RECT 718.950 252.450 721.050 253.050 ;
        RECT 754.950 252.450 757.050 253.050 ;
        RECT 790.950 252.450 793.050 253.050 ;
        RECT 814.950 252.450 817.050 252.900 ;
        RECT 718.950 252.000 780.450 252.450 ;
        RECT 718.950 251.400 781.050 252.000 ;
        RECT 718.950 250.950 721.050 251.400 ;
        RECT 754.950 250.950 757.050 251.400 ;
        RECT 25.950 247.950 31.050 250.050 ;
        RECT 79.950 249.450 82.050 250.050 ;
        RECT 148.950 249.450 151.050 250.050 ;
        RECT 79.950 248.400 151.050 249.450 ;
        RECT 79.950 247.950 82.050 248.400 ;
        RECT 148.950 247.950 151.050 248.400 ;
        RECT 190.950 249.450 193.050 250.050 ;
        RECT 196.950 249.450 199.050 250.050 ;
        RECT 247.950 249.450 250.050 250.050 ;
        RECT 286.950 249.450 289.050 250.050 ;
        RECT 190.950 248.400 289.050 249.450 ;
        RECT 190.950 247.950 193.050 248.400 ;
        RECT 196.950 247.950 199.050 248.400 ;
        RECT 247.950 247.950 250.050 248.400 ;
        RECT 286.950 247.950 289.050 248.400 ;
        RECT 367.950 249.450 370.050 250.050 ;
        RECT 415.950 249.450 418.050 250.050 ;
        RECT 469.950 249.450 472.050 250.050 ;
        RECT 523.950 249.450 526.050 250.050 ;
        RECT 583.950 249.450 586.050 250.050 ;
        RECT 367.950 248.400 472.050 249.450 ;
        RECT 367.950 247.950 370.050 248.400 ;
        RECT 415.950 247.950 418.050 248.400 ;
        RECT 469.950 247.950 472.050 248.400 ;
        RECT 506.400 248.400 586.050 249.450 ;
        RECT 235.950 247.050 238.050 247.200 ;
        RECT 16.950 246.450 19.050 247.050 ;
        RECT 97.950 246.450 100.050 247.050 ;
        RECT 124.950 246.450 127.050 247.050 ;
        RECT 16.950 245.400 75.450 246.450 ;
        RECT 16.950 244.950 19.050 245.400 ;
        RECT 46.950 243.450 49.050 244.050 ;
        RECT 70.950 243.450 73.050 244.050 ;
        RECT 46.950 242.400 73.050 243.450 ;
        RECT 74.400 243.450 75.450 245.400 ;
        RECT 97.950 245.400 127.050 246.450 ;
        RECT 97.950 244.950 100.050 245.400 ;
        RECT 124.950 244.950 127.050 245.400 ;
        RECT 157.950 246.450 160.050 247.050 ;
        RECT 169.950 246.450 172.050 247.050 ;
        RECT 157.950 245.400 172.050 246.450 ;
        RECT 157.950 244.950 160.050 245.400 ;
        RECT 169.950 244.950 172.050 245.400 ;
        RECT 232.950 245.100 238.050 247.050 ;
        RECT 253.950 246.450 256.050 247.050 ;
        RECT 262.950 246.450 265.050 247.050 ;
        RECT 253.950 245.400 265.050 246.450 ;
        RECT 232.950 244.950 237.000 245.100 ;
        RECT 253.950 244.950 256.050 245.400 ;
        RECT 262.950 244.950 265.050 245.400 ;
        RECT 316.950 246.450 319.050 247.050 ;
        RECT 343.950 246.450 346.050 247.050 ;
        RECT 433.950 246.450 436.050 247.200 ;
        RECT 506.400 246.450 507.450 248.400 ;
        RECT 523.950 247.950 526.050 248.400 ;
        RECT 583.950 247.950 586.050 248.400 ;
        RECT 649.950 249.450 652.050 250.050 ;
        RECT 679.950 249.450 682.050 250.050 ;
        RECT 694.800 249.450 696.900 249.900 ;
        RECT 649.950 248.400 696.900 249.450 ;
        RECT 649.950 247.950 652.050 248.400 ;
        RECT 679.950 247.950 682.050 248.400 ;
        RECT 694.800 247.800 696.900 248.400 ;
        RECT 698.100 249.450 700.200 250.050 ;
        RECT 706.950 249.450 709.050 250.050 ;
        RECT 698.100 248.400 709.050 249.450 ;
        RECT 698.100 247.950 700.200 248.400 ;
        RECT 706.950 247.950 709.050 248.400 ;
        RECT 727.950 249.450 730.050 250.050 ;
        RECT 742.950 249.450 745.050 250.050 ;
        RECT 727.950 248.400 745.050 249.450 ;
        RECT 727.950 247.950 730.050 248.400 ;
        RECT 742.950 247.950 745.050 248.400 ;
        RECT 778.950 247.950 781.050 251.400 ;
        RECT 790.950 251.400 817.050 252.450 ;
        RECT 790.950 250.950 793.050 251.400 ;
        RECT 814.950 250.800 817.050 251.400 ;
        RECT 832.950 252.450 835.050 253.050 ;
        RECT 850.950 252.450 853.050 253.050 ;
        RECT 856.950 252.450 859.050 253.050 ;
        RECT 832.950 251.400 849.450 252.450 ;
        RECT 832.950 250.950 835.050 251.400 ;
        RECT 848.400 250.050 849.450 251.400 ;
        RECT 850.950 251.400 859.050 252.450 ;
        RECT 850.950 250.950 853.050 251.400 ;
        RECT 856.950 250.950 859.050 251.400 ;
        RECT 799.950 249.450 802.050 250.050 ;
        RECT 820.950 249.450 823.050 250.050 ;
        RECT 799.950 248.400 823.050 249.450 ;
        RECT 799.950 247.950 802.050 248.400 ;
        RECT 820.950 247.950 823.050 248.400 ;
        RECT 838.950 247.950 844.050 250.050 ;
        RECT 848.400 248.400 853.050 250.050 ;
        RECT 849.000 247.950 853.050 248.400 ;
        RECT 316.950 246.000 393.450 246.450 ;
        RECT 316.950 245.400 394.050 246.000 ;
        RECT 316.950 244.950 319.050 245.400 ;
        RECT 343.950 244.950 346.050 245.400 ;
        RECT 109.950 243.450 112.050 244.050 ;
        RECT 74.400 242.400 102.450 243.450 ;
        RECT 46.950 241.950 49.050 242.400 ;
        RECT 56.400 241.050 57.450 242.400 ;
        RECT 70.950 241.950 73.050 242.400 ;
        RECT 4.950 240.450 7.050 241.050 ;
        RECT 13.950 240.450 16.050 241.050 ;
        RECT 4.950 239.400 16.050 240.450 ;
        RECT 4.950 238.950 7.050 239.400 ;
        RECT 13.950 238.950 16.050 239.400 ;
        RECT 19.950 240.450 22.050 241.050 ;
        RECT 28.950 240.450 31.050 241.050 ;
        RECT 34.800 240.450 36.900 241.050 ;
        RECT 19.950 239.400 36.900 240.450 ;
        RECT 19.950 238.950 22.050 239.400 ;
        RECT 28.950 238.950 31.050 239.400 ;
        RECT 34.800 238.950 36.900 239.400 ;
        RECT 38.100 240.450 40.200 241.050 ;
        RECT 52.950 240.450 55.050 241.050 ;
        RECT 38.100 239.400 55.050 240.450 ;
        RECT 56.400 239.400 61.050 241.050 ;
        RECT 38.100 238.950 40.200 239.400 ;
        RECT 52.950 238.950 55.050 239.400 ;
        RECT 57.000 238.950 61.050 239.400 ;
        RECT 10.950 232.950 13.050 238.050 ;
        RECT 16.950 235.950 22.050 238.050 ;
        RECT 16.950 234.450 19.050 234.900 ;
        RECT 34.950 234.450 37.050 238.050 ;
        RECT 40.950 237.450 43.050 238.050 ;
        RECT 49.950 237.450 52.050 238.050 ;
        RECT 40.950 236.400 52.050 237.450 ;
        RECT 40.950 235.950 43.050 236.400 ;
        RECT 49.950 235.950 52.050 236.400 ;
        RECT 46.950 234.450 49.050 235.050 ;
        RECT 16.950 233.400 49.050 234.450 ;
        RECT 16.950 232.800 19.050 233.400 ;
        RECT 46.950 232.950 49.050 233.400 ;
        RECT 55.950 232.950 58.050 238.050 ;
        RECT 61.950 235.950 67.050 238.050 ;
        RECT 70.950 235.950 73.050 241.050 ;
        RECT 85.950 240.450 88.050 241.050 ;
        RECT 77.400 240.000 88.050 240.450 ;
        RECT 76.950 239.400 88.050 240.000 ;
        RECT 76.950 235.950 79.050 239.400 ;
        RECT 85.950 238.950 88.050 239.400 ;
        RECT 97.950 235.950 100.050 241.050 ;
        RECT 101.400 240.450 102.450 242.400 ;
        RECT 109.950 243.000 135.450 243.450 ;
        RECT 109.950 242.400 136.050 243.000 ;
        RECT 109.950 241.950 112.050 242.400 ;
        RECT 112.800 240.450 114.900 241.050 ;
        RECT 101.400 239.400 114.900 240.450 ;
        RECT 112.800 238.950 114.900 239.400 ;
        RECT 116.100 240.450 118.200 241.050 ;
        RECT 121.800 240.450 123.900 241.050 ;
        RECT 116.100 239.400 123.900 240.450 ;
        RECT 125.100 240.000 127.200 241.050 ;
        RECT 116.100 238.950 118.200 239.400 ;
        RECT 121.800 238.950 123.900 239.400 ;
        RECT 124.950 238.950 127.200 240.000 ;
        RECT 133.950 238.950 136.050 242.400 ;
        RECT 139.950 238.950 142.050 244.050 ;
        RECT 169.950 243.450 172.050 244.050 ;
        RECT 190.950 243.450 193.050 244.050 ;
        RECT 217.950 243.450 220.050 244.050 ;
        RECT 235.950 243.450 238.050 243.900 ;
        RECT 169.950 242.400 216.450 243.450 ;
        RECT 169.950 241.950 172.050 242.400 ;
        RECT 190.950 241.950 193.050 242.400 ;
        RECT 151.800 240.450 153.900 241.050 ;
        RECT 146.400 239.400 153.900 240.450 ;
        RECT 103.950 237.450 106.050 238.050 ;
        RECT 118.950 237.450 121.050 238.050 ;
        RECT 103.950 236.400 121.050 237.450 ;
        RECT 103.950 235.950 106.050 236.400 ;
        RECT 65.400 234.450 66.450 235.950 ;
        RECT 73.800 234.450 75.900 235.050 ;
        RECT 65.400 233.400 75.900 234.450 ;
        RECT 73.800 232.950 75.900 233.400 ;
        RECT 77.100 232.950 82.050 235.050 ;
        RECT 100.950 234.450 106.050 235.050 ;
        RECT 115.950 234.450 118.050 235.050 ;
        RECT 100.950 233.400 118.050 234.450 ;
        RECT 118.950 234.450 121.050 236.400 ;
        RECT 124.950 235.950 127.050 238.950 ;
        RECT 146.400 238.050 147.450 239.400 ;
        RECT 151.800 238.950 153.900 239.400 ;
        RECT 155.100 238.950 160.050 241.050 ;
        RECT 166.950 240.450 169.050 241.050 ;
        RECT 172.950 240.450 175.050 241.050 ;
        RECT 166.950 239.400 189.450 240.450 ;
        RECT 166.950 238.950 169.050 239.400 ;
        RECT 172.950 238.950 175.050 239.400 ;
        RECT 136.950 235.050 139.050 238.050 ;
        RECT 142.950 236.400 147.450 238.050 ;
        RECT 148.950 237.450 151.050 238.050 ;
        RECT 154.950 237.450 157.050 238.050 ;
        RECT 148.950 236.400 157.050 237.450 ;
        RECT 142.950 235.950 147.000 236.400 ;
        RECT 148.950 235.950 151.050 236.400 ;
        RECT 154.950 235.950 157.050 236.400 ;
        RECT 133.800 234.450 135.900 235.050 ;
        RECT 118.950 234.000 135.900 234.450 ;
        RECT 136.950 234.000 139.200 235.050 ;
        RECT 119.400 233.400 135.900 234.000 ;
        RECT 100.950 232.950 106.050 233.400 ;
        RECT 115.950 232.950 118.050 233.400 ;
        RECT 133.800 232.950 135.900 233.400 ;
        RECT 137.100 232.950 139.200 234.000 ;
        RECT 160.950 232.950 163.050 238.050 ;
        RECT 169.950 237.450 172.050 238.050 ;
        RECT 175.950 237.450 178.050 238.050 ;
        RECT 169.950 236.400 178.050 237.450 ;
        RECT 169.950 235.950 172.050 236.400 ;
        RECT 175.950 235.950 178.050 236.400 ;
        RECT 181.950 235.950 187.050 238.050 ;
        RECT 188.400 237.450 189.450 239.400 ;
        RECT 196.950 238.950 199.050 242.400 ;
        RECT 215.400 241.050 216.450 242.400 ;
        RECT 217.950 242.400 238.050 243.450 ;
        RECT 217.950 241.950 220.050 242.400 ;
        RECT 235.950 241.800 238.050 242.400 ;
        RECT 280.950 243.450 283.050 244.050 ;
        RECT 289.950 243.450 292.050 244.050 ;
        RECT 280.950 242.400 292.050 243.450 ;
        RECT 280.950 241.950 283.050 242.400 ;
        RECT 289.950 241.950 292.050 242.400 ;
        RECT 319.950 243.450 322.050 244.050 ;
        RECT 328.950 243.450 331.050 244.050 ;
        RECT 319.950 242.400 331.050 243.450 ;
        RECT 319.950 241.950 322.050 242.400 ;
        RECT 328.950 241.950 331.050 242.400 ;
        RECT 391.950 243.450 394.050 245.400 ;
        RECT 433.950 245.400 507.450 246.450 ;
        RECT 508.950 246.450 511.050 247.050 ;
        RECT 514.950 246.450 517.050 247.050 ;
        RECT 508.950 245.400 517.050 246.450 ;
        RECT 589.950 245.400 592.050 247.500 ;
        RECT 610.950 245.400 613.050 247.500 ;
        RECT 631.950 247.050 634.050 247.200 ;
        RECT 433.950 245.100 436.050 245.400 ;
        RECT 508.950 244.950 511.050 245.400 ;
        RECT 514.950 244.950 517.050 245.400 ;
        RECT 391.950 243.000 423.450 243.450 ;
        RECT 391.950 242.400 424.050 243.000 ;
        RECT 391.950 241.950 394.050 242.400 ;
        RECT 202.950 240.450 205.050 241.050 ;
        RECT 211.950 240.450 214.050 241.050 ;
        RECT 202.950 239.400 214.050 240.450 ;
        RECT 215.400 239.400 219.900 241.050 ;
        RECT 202.950 238.950 205.050 239.400 ;
        RECT 211.950 238.950 214.050 239.400 ;
        RECT 216.000 238.950 219.900 239.400 ;
        RECT 221.100 238.950 226.050 241.050 ;
        RECT 253.950 240.450 256.050 241.050 ;
        RECT 262.950 240.450 265.050 241.050 ;
        RECT 253.950 239.400 265.050 240.450 ;
        RECT 253.950 238.950 256.050 239.400 ;
        RECT 262.950 238.950 265.050 239.400 ;
        RECT 199.950 237.450 202.050 238.050 ;
        RECT 188.400 236.400 202.050 237.450 ;
        RECT 199.950 235.950 202.050 236.400 ;
        RECT 58.950 231.450 61.050 232.050 ;
        RECT 85.950 231.450 88.050 232.050 ;
        RECT 58.950 230.400 88.050 231.450 ;
        RECT 58.950 229.950 61.050 230.400 ;
        RECT 85.950 229.950 88.050 230.400 ;
        RECT 148.950 231.450 151.050 232.050 ;
        RECT 178.950 231.450 181.050 235.050 ;
        RECT 205.950 234.450 208.050 238.050 ;
        RECT 217.950 235.950 223.050 238.050 ;
        RECT 226.950 237.450 229.050 238.050 ;
        RECT 235.950 237.450 240.900 238.050 ;
        RECT 226.950 236.400 240.900 237.450 ;
        RECT 226.950 235.950 229.050 236.400 ;
        RECT 235.950 235.950 240.900 236.400 ;
        RECT 241.800 237.000 243.900 238.050 ;
        RECT 241.800 235.950 244.050 237.000 ;
        RECT 245.100 235.950 250.050 238.050 ;
        RECT 256.950 235.950 262.050 238.050 ;
        RECT 223.950 234.450 226.050 235.050 ;
        RECT 205.950 234.000 226.050 234.450 ;
        RECT 206.400 233.400 226.050 234.000 ;
        RECT 223.950 232.950 226.050 233.400 ;
        RECT 241.950 232.950 244.050 235.950 ;
        RECT 265.950 232.950 268.050 238.050 ;
        RECT 280.950 235.950 283.050 241.050 ;
        RECT 286.950 235.950 289.050 241.050 ;
        RECT 301.950 238.950 307.050 241.050 ;
        RECT 337.950 240.450 340.050 241.050 ;
        RECT 343.950 240.450 346.050 241.050 ;
        RECT 337.950 239.400 346.050 240.450 ;
        RECT 337.950 238.950 340.050 239.400 ;
        RECT 343.950 238.950 346.050 239.400 ;
        RECT 352.950 240.450 355.050 241.050 ;
        RECT 352.950 239.400 363.450 240.450 ;
        RECT 352.950 238.950 355.050 239.400 ;
        RECT 362.400 238.050 363.450 239.400 ;
        RECT 295.950 237.450 298.050 238.050 ;
        RECT 301.950 237.450 304.050 238.050 ;
        RECT 295.950 236.400 304.050 237.450 ;
        RECT 295.950 235.950 298.050 236.400 ;
        RECT 301.950 235.950 304.050 236.400 ;
        RECT 307.950 237.450 310.050 238.050 ;
        RECT 319.950 237.450 325.050 238.050 ;
        RECT 307.950 236.400 325.050 237.450 ;
        RECT 307.950 235.950 310.050 236.400 ;
        RECT 319.950 235.950 325.050 236.400 ;
        RECT 328.950 235.950 334.050 238.050 ;
        RECT 343.950 237.450 346.050 238.050 ;
        RECT 349.950 237.450 352.050 238.050 ;
        RECT 343.950 236.400 352.050 237.450 ;
        RECT 343.950 235.950 346.050 236.400 ;
        RECT 349.950 235.950 352.050 236.400 ;
        RECT 355.950 235.950 361.050 238.050 ;
        RECT 362.400 235.950 367.050 238.050 ;
        RECT 370.950 235.950 373.050 241.050 ;
        RECT 403.950 238.950 409.050 241.050 ;
        RECT 412.950 238.950 418.050 241.050 ;
        RECT 421.950 238.950 424.050 242.400 ;
        RECT 427.950 241.050 430.050 244.050 ;
        RECT 433.950 243.450 436.050 243.900 ;
        RECT 454.950 243.450 457.050 244.200 ;
        RECT 484.950 243.450 487.050 244.050 ;
        RECT 433.950 242.400 457.050 243.450 ;
        RECT 479.400 243.000 489.450 243.450 ;
        RECT 506.400 243.000 522.450 243.450 ;
        RECT 433.950 241.800 436.050 242.400 ;
        RECT 454.950 242.100 457.050 242.400 ;
        RECT 478.950 242.400 489.450 243.000 ;
        RECT 427.800 240.000 430.050 241.050 ;
        RECT 431.100 240.450 433.200 241.050 ;
        RECT 454.950 240.450 457.050 240.900 ;
        RECT 427.800 238.950 429.900 240.000 ;
        RECT 431.100 239.400 457.050 240.450 ;
        RECT 458.400 240.000 474.450 240.450 ;
        RECT 431.100 238.950 433.200 239.400 ;
        RECT 391.950 237.450 394.050 238.050 ;
        RECT 403.950 237.450 406.050 238.050 ;
        RECT 391.950 236.400 406.050 237.450 ;
        RECT 391.950 235.950 394.050 236.400 ;
        RECT 403.950 235.950 406.050 236.400 ;
        RECT 148.950 231.000 181.050 231.450 ;
        RECT 199.950 231.450 202.050 232.050 ;
        RECT 217.950 231.450 220.050 232.050 ;
        RECT 148.950 230.400 180.450 231.000 ;
        RECT 199.950 230.400 220.050 231.450 ;
        RECT 148.950 229.950 151.050 230.400 ;
        RECT 199.950 229.950 202.050 230.400 ;
        RECT 217.950 229.950 220.050 230.400 ;
        RECT 283.950 229.950 286.050 235.050 ;
        RECT 292.950 234.450 295.050 235.050 ;
        RECT 304.950 234.450 307.050 235.050 ;
        RECT 325.950 234.450 328.050 235.050 ;
        RECT 292.950 233.400 328.050 234.450 ;
        RECT 292.950 232.950 295.050 233.400 ;
        RECT 304.950 232.950 307.050 233.400 ;
        RECT 325.950 232.950 328.050 233.400 ;
        RECT 334.950 234.450 337.050 235.050 ;
        RECT 362.400 234.450 363.450 235.950 ;
        RECT 409.950 235.050 412.050 238.050 ;
        RECT 416.400 237.450 417.450 238.950 ;
        RECT 454.950 238.800 457.050 239.400 ;
        RECT 457.950 239.400 474.450 240.000 ;
        RECT 424.950 237.450 427.050 238.050 ;
        RECT 416.400 236.400 427.050 237.450 ;
        RECT 424.950 235.950 427.050 236.400 ;
        RECT 334.950 233.400 363.450 234.450 ;
        RECT 334.950 232.950 337.050 233.400 ;
        RECT 367.950 231.450 370.050 235.050 ;
        RECT 406.950 234.000 412.050 235.050 ;
        RECT 406.950 233.400 411.450 234.000 ;
        RECT 406.950 232.950 411.000 233.400 ;
        RECT 430.950 232.950 433.050 238.050 ;
        RECT 439.950 237.450 442.050 238.050 ;
        RECT 445.950 237.450 448.050 238.050 ;
        RECT 439.950 236.400 448.050 237.450 ;
        RECT 439.950 235.950 442.050 236.400 ;
        RECT 445.950 235.950 448.050 236.400 ;
        RECT 457.950 235.950 460.050 239.400 ;
        RECT 466.950 238.050 469.050 239.400 ;
        RECT 463.800 237.000 465.900 238.050 ;
        RECT 466.800 237.000 469.050 238.050 ;
        RECT 470.100 237.000 472.200 238.050 ;
        RECT 463.800 235.950 466.050 237.000 ;
        RECT 466.800 235.950 468.900 237.000 ;
        RECT 469.950 235.950 472.200 237.000 ;
        RECT 473.400 237.450 474.450 239.400 ;
        RECT 478.950 238.950 481.050 242.400 ;
        RECT 484.950 241.950 487.050 242.400 ;
        RECT 488.400 240.450 489.450 242.400 ;
        RECT 505.950 242.400 523.050 243.000 ;
        RECT 499.950 240.450 502.050 241.050 ;
        RECT 488.400 239.400 502.050 240.450 ;
        RECT 499.950 238.950 502.050 239.400 ;
        RECT 505.950 238.950 508.050 242.400 ;
        RECT 520.950 238.950 523.050 242.400 ;
        RECT 526.950 238.950 529.050 244.050 ;
        RECT 562.950 241.950 571.050 244.050 ;
        RECT 580.950 243.450 583.050 244.050 ;
        RECT 580.950 243.000 588.450 243.450 ;
        RECT 580.950 242.400 589.050 243.000 ;
        RECT 580.950 241.950 583.050 242.400 ;
        RECT 535.950 240.450 538.050 241.050 ;
        RECT 535.950 240.000 564.450 240.450 ;
        RECT 535.950 239.400 565.050 240.000 ;
        RECT 535.950 238.950 538.050 239.400 ;
        RECT 484.950 237.450 487.050 238.050 ;
        RECT 502.950 237.450 505.050 238.050 ;
        RECT 473.400 236.400 505.050 237.450 ;
        RECT 484.950 235.950 487.050 236.400 ;
        RECT 502.950 235.950 505.050 236.400 ;
        RECT 520.950 235.950 526.050 238.050 ;
        RECT 529.950 237.450 532.050 238.050 ;
        RECT 544.950 237.450 547.050 238.050 ;
        RECT 529.950 236.400 547.050 237.450 ;
        RECT 529.950 235.950 532.050 236.400 ;
        RECT 544.950 235.950 547.050 236.400 ;
        RECT 562.950 235.950 565.050 239.400 ;
        RECT 586.950 238.950 589.050 242.400 ;
        RECT 571.950 235.950 577.050 238.050 ;
        RECT 442.800 234.000 444.900 235.050 ;
        RECT 442.800 232.950 445.050 234.000 ;
        RECT 446.100 232.950 451.050 235.050 ;
        RECT 463.950 232.950 466.050 235.950 ;
        RECT 469.950 232.950 472.050 235.950 ;
        RECT 505.950 234.450 508.050 235.050 ;
        RECT 532.950 234.450 535.050 235.050 ;
        RECT 505.950 233.400 535.050 234.450 ;
        RECT 505.950 232.950 508.050 233.400 ;
        RECT 532.950 232.950 535.050 233.400 ;
        RECT 538.950 234.450 541.050 235.050 ;
        RECT 547.950 234.450 553.050 235.050 ;
        RECT 538.950 233.400 553.050 234.450 ;
        RECT 590.850 233.400 592.050 245.400 ;
        RECT 595.950 238.950 601.050 241.050 ;
        RECT 604.950 238.950 607.050 244.050 ;
        RECT 538.950 232.950 541.050 233.400 ;
        RECT 547.950 232.950 553.050 233.400 ;
        RECT 403.950 231.450 406.050 232.050 ;
        RECT 367.950 231.000 406.050 231.450 ;
        RECT 368.400 230.400 406.050 231.000 ;
        RECT 403.950 229.950 406.050 230.400 ;
        RECT 427.950 231.450 430.050 232.050 ;
        RECT 442.950 231.450 445.050 232.950 ;
        RECT 427.950 231.000 445.050 231.450 ;
        RECT 493.950 231.450 496.050 232.050 ;
        RECT 523.950 231.450 526.050 232.050 ;
        RECT 427.950 230.400 444.300 231.000 ;
        RECT 493.950 230.400 526.050 231.450 ;
        RECT 589.950 231.300 592.050 233.400 ;
        RECT 427.950 229.950 430.050 230.400 ;
        RECT 493.950 229.950 496.050 230.400 ;
        RECT 523.950 229.950 526.050 230.400 ;
        RECT 160.950 228.450 163.050 229.050 ;
        RECT 181.950 228.450 184.050 229.050 ;
        RECT 160.950 227.400 184.050 228.450 ;
        RECT 160.950 226.950 163.050 227.400 ;
        RECT 181.950 226.950 184.050 227.400 ;
        RECT 211.950 228.450 214.050 229.050 ;
        RECT 256.950 228.450 259.050 229.050 ;
        RECT 211.950 227.400 259.050 228.450 ;
        RECT 211.950 226.950 214.050 227.400 ;
        RECT 256.950 226.950 259.050 227.400 ;
        RECT 274.950 228.450 277.050 229.050 ;
        RECT 412.950 228.450 415.050 229.050 ;
        RECT 274.950 227.400 415.050 228.450 ;
        RECT 274.950 226.950 277.050 227.400 ;
        RECT 412.950 226.950 415.050 227.400 ;
        RECT 418.950 228.450 421.050 229.050 ;
        RECT 463.950 228.450 466.050 229.050 ;
        RECT 418.950 227.400 466.050 228.450 ;
        RECT 590.850 227.700 592.050 231.300 ;
        RECT 611.100 228.600 612.300 245.400 ;
        RECT 631.950 245.100 637.050 247.050 ;
        RECT 633.000 244.950 637.050 245.100 ;
        RECT 736.950 246.450 739.050 247.050 ;
        RECT 772.950 246.450 775.050 247.050 ;
        RECT 793.950 246.450 796.050 247.050 ;
        RECT 736.950 245.400 775.050 246.450 ;
        RECT 736.950 244.950 739.050 245.400 ;
        RECT 772.950 244.950 775.050 245.400 ;
        RECT 776.400 245.400 796.050 246.450 ;
        RECT 619.950 243.450 622.050 244.050 ;
        RECT 625.950 243.450 628.050 244.050 ;
        RECT 631.950 243.450 634.050 243.900 ;
        RECT 619.950 242.400 634.050 243.450 ;
        RECT 619.950 241.950 622.050 242.400 ;
        RECT 625.950 241.950 628.050 242.400 ;
        RECT 631.950 241.800 634.050 242.400 ;
        RECT 637.950 243.450 640.050 244.050 ;
        RECT 646.950 243.450 649.050 244.050 ;
        RECT 637.950 242.400 649.050 243.450 ;
        RECT 637.950 241.950 640.050 242.400 ;
        RECT 646.950 241.950 649.050 242.400 ;
        RECT 658.950 243.450 661.050 244.050 ;
        RECT 667.950 243.450 670.050 244.050 ;
        RECT 658.950 242.400 670.050 243.450 ;
        RECT 658.950 241.950 661.050 242.400 ;
        RECT 667.950 241.950 670.050 242.400 ;
        RECT 628.950 240.450 631.050 241.050 ;
        RECT 628.950 240.000 678.450 240.450 ;
        RECT 628.950 239.400 679.050 240.000 ;
        RECT 628.950 238.950 631.050 239.400 ;
        RECT 619.950 237.450 622.050 238.050 ;
        RECT 628.800 237.450 630.900 238.050 ;
        RECT 619.950 236.400 630.900 237.450 ;
        RECT 619.950 235.950 622.050 236.400 ;
        RECT 628.800 235.950 630.900 236.400 ;
        RECT 632.100 237.450 634.200 238.050 ;
        RECT 643.800 237.450 645.900 238.050 ;
        RECT 632.100 236.400 645.900 237.450 ;
        RECT 647.100 237.000 649.200 238.050 ;
        RECT 632.100 235.950 634.200 236.400 ;
        RECT 643.800 235.950 645.900 236.400 ;
        RECT 646.950 235.950 649.200 237.000 ;
        RECT 652.950 237.450 655.050 238.050 ;
        RECT 664.950 237.450 670.050 238.050 ;
        RECT 652.950 236.400 670.050 237.450 ;
        RECT 652.950 235.950 655.050 236.400 ;
        RECT 664.950 235.950 670.050 236.400 ;
        RECT 676.950 235.950 679.050 239.400 ;
        RECT 679.950 238.950 682.050 244.050 ;
        RECT 715.950 243.450 718.050 244.050 ;
        RECT 724.950 243.450 729.000 244.050 ;
        RECT 715.950 243.000 723.600 243.450 ;
        RECT 724.950 243.000 729.450 243.450 ;
        RECT 742.800 243.000 744.900 244.050 ;
        RECT 715.950 242.400 724.050 243.000 ;
        RECT 715.950 241.950 718.050 242.400 ;
        RECT 721.950 241.050 724.050 242.400 ;
        RECT 724.950 241.950 730.050 243.000 ;
        RECT 742.800 241.950 745.050 243.000 ;
        RECT 688.950 240.450 691.050 241.050 ;
        RECT 706.950 240.450 709.050 241.050 ;
        RECT 688.950 239.400 709.050 240.450 ;
        RECT 688.950 238.950 691.050 239.400 ;
        RECT 706.950 238.950 709.050 239.400 ;
        RECT 712.950 240.450 715.050 241.050 ;
        RECT 718.800 240.450 720.900 241.050 ;
        RECT 712.950 239.400 720.900 240.450 ;
        RECT 712.950 238.950 715.050 239.400 ;
        RECT 718.800 238.950 720.900 239.400 ;
        RECT 721.950 238.950 724.200 241.050 ;
        RECT 727.950 238.950 730.050 241.950 ;
        RECT 742.950 241.050 745.050 241.950 ;
        RECT 742.800 240.000 745.050 241.050 ;
        RECT 742.800 238.950 744.900 240.000 ;
        RECT 746.100 238.950 751.050 241.050 ;
        RECT 754.950 240.450 757.050 241.050 ;
        RECT 763.950 240.450 766.050 241.050 ;
        RECT 754.950 239.400 766.050 240.450 ;
        RECT 754.950 238.950 757.050 239.400 ;
        RECT 763.950 238.950 766.050 239.400 ;
        RECT 769.950 238.950 772.050 244.050 ;
        RECT 721.950 238.050 724.050 238.950 ;
        RECT 776.400 238.050 777.450 245.400 ;
        RECT 793.950 244.950 796.050 245.400 ;
        RECT 841.950 246.450 844.050 247.050 ;
        RECT 850.950 246.450 853.050 247.050 ;
        RECT 841.950 245.400 853.050 246.450 ;
        RECT 841.950 244.950 844.050 245.400 ;
        RECT 850.950 244.950 853.050 245.400 ;
        RECT 799.950 243.450 802.050 244.050 ;
        RECT 808.950 243.450 811.050 244.050 ;
        RECT 799.950 242.400 811.050 243.450 ;
        RECT 799.950 241.950 802.050 242.400 ;
        RECT 808.950 241.950 811.050 242.400 ;
        RECT 844.950 243.450 847.050 244.050 ;
        RECT 856.950 243.450 859.050 244.050 ;
        RECT 844.950 242.400 859.050 243.450 ;
        RECT 844.950 241.950 847.050 242.400 ;
        RECT 856.950 241.950 859.050 242.400 ;
        RECT 778.950 240.450 781.050 241.050 ;
        RECT 787.950 240.450 790.050 241.050 ;
        RECT 778.950 239.400 790.050 240.450 ;
        RECT 778.950 238.950 781.050 239.400 ;
        RECT 787.950 238.950 790.050 239.400 ;
        RECT 814.950 240.450 817.050 241.050 ;
        RECT 814.950 239.400 822.450 240.450 ;
        RECT 814.950 238.950 817.050 239.400 ;
        RECT 685.950 237.450 688.050 238.050 ;
        RECT 680.400 236.400 688.050 237.450 ;
        RECT 646.950 235.050 649.050 235.950 ;
        RECT 613.950 231.450 616.050 232.050 ;
        RECT 622.950 231.450 625.050 232.050 ;
        RECT 613.950 230.400 625.050 231.450 ;
        RECT 613.950 229.950 616.050 230.400 ;
        RECT 622.950 229.950 625.050 230.400 ;
        RECT 631.950 231.450 634.050 232.050 ;
        RECT 640.950 231.450 643.050 235.050 ;
        RECT 646.800 234.000 649.050 235.050 ;
        RECT 650.100 234.450 652.200 235.050 ;
        RECT 661.950 234.450 664.050 235.050 ;
        RECT 646.800 232.950 648.900 234.000 ;
        RECT 650.100 233.400 664.050 234.450 ;
        RECT 650.100 232.950 652.200 233.400 ;
        RECT 661.950 232.950 664.050 233.400 ;
        RECT 667.950 234.450 673.050 235.050 ;
        RECT 680.400 234.450 681.450 236.400 ;
        RECT 685.950 235.950 688.050 236.400 ;
        RECT 694.950 237.450 697.050 238.050 ;
        RECT 703.950 237.450 706.050 238.050 ;
        RECT 694.950 236.400 706.050 237.450 ;
        RECT 694.950 235.950 697.050 236.400 ;
        RECT 703.950 235.950 706.050 236.400 ;
        RECT 709.950 237.450 712.050 238.050 ;
        RECT 715.950 237.450 718.050 238.050 ;
        RECT 709.950 236.400 718.050 237.450 ;
        RECT 709.950 235.950 712.050 236.400 ;
        RECT 715.950 235.950 718.050 236.400 ;
        RECT 721.800 237.000 724.050 238.050 ;
        RECT 725.100 237.000 727.200 238.050 ;
        RECT 721.800 235.950 723.900 237.000 ;
        RECT 724.950 235.950 727.200 237.000 ;
        RECT 730.950 237.450 733.050 238.050 ;
        RECT 742.800 237.450 744.900 238.050 ;
        RECT 730.950 236.400 744.900 237.450 ;
        RECT 746.100 237.000 748.200 238.050 ;
        RECT 730.950 235.950 733.050 236.400 ;
        RECT 742.800 235.950 744.900 236.400 ;
        RECT 745.950 235.950 748.200 237.000 ;
        RECT 751.950 237.450 754.050 238.050 ;
        RECT 757.950 237.450 760.050 238.050 ;
        RECT 751.950 236.400 760.050 237.450 ;
        RECT 751.950 235.950 754.050 236.400 ;
        RECT 757.950 235.950 760.050 236.400 ;
        RECT 700.950 234.450 703.050 235.050 ;
        RECT 667.950 233.400 681.450 234.450 ;
        RECT 689.400 233.400 703.050 234.450 ;
        RECT 667.950 232.950 673.050 233.400 ;
        RECT 652.950 231.450 655.050 232.050 ;
        RECT 631.950 230.400 655.050 231.450 ;
        RECT 631.950 229.950 634.050 230.400 ;
        RECT 652.950 229.950 655.050 230.400 ;
        RECT 673.950 231.450 676.050 232.050 ;
        RECT 689.400 231.450 690.450 233.400 ;
        RECT 700.950 232.950 703.050 233.400 ;
        RECT 709.950 234.450 712.050 235.050 ;
        RECT 724.950 234.450 727.050 235.950 ;
        RECT 745.950 234.450 748.050 235.950 ;
        RECT 709.950 234.000 748.050 234.450 ;
        RECT 766.950 234.450 769.050 238.050 ;
        RECT 772.950 236.400 777.450 238.050 ;
        RECT 778.950 237.450 781.050 238.050 ;
        RECT 784.950 237.450 787.050 238.050 ;
        RECT 778.950 236.400 787.050 237.450 ;
        RECT 772.950 235.950 777.000 236.400 ;
        RECT 778.950 235.950 781.050 236.400 ;
        RECT 784.950 235.950 787.050 236.400 ;
        RECT 775.950 234.450 778.050 235.050 ;
        RECT 766.950 234.000 778.050 234.450 ;
        RECT 709.950 233.400 747.600 234.000 ;
        RECT 767.400 233.400 778.050 234.000 ;
        RECT 709.950 232.950 712.050 233.400 ;
        RECT 775.950 232.950 778.050 233.400 ;
        RECT 790.950 232.950 793.050 238.050 ;
        RECT 811.950 235.950 814.050 238.050 ;
        RECT 673.950 230.400 690.450 231.450 ;
        RECT 721.950 231.450 724.050 232.050 ;
        RECT 757.950 231.450 760.050 232.050 ;
        RECT 721.950 230.400 760.050 231.450 ;
        RECT 673.950 229.950 676.050 230.400 ;
        RECT 721.950 229.950 724.050 230.400 ;
        RECT 757.950 229.950 760.050 230.400 ;
        RECT 766.950 231.450 769.050 232.050 ;
        RECT 812.400 231.450 813.450 235.950 ;
        RECT 817.950 234.450 820.050 238.050 ;
        RECT 821.400 237.450 822.450 239.400 ;
        RECT 823.950 238.950 829.050 241.050 ;
        RECT 832.950 240.450 835.050 241.050 ;
        RECT 841.950 240.450 844.050 241.050 ;
        RECT 832.950 239.400 844.050 240.450 ;
        RECT 832.950 238.950 835.050 239.400 ;
        RECT 841.950 238.950 844.050 239.400 ;
        RECT 828.000 237.900 831.900 238.050 ;
        RECT 826.950 237.450 831.900 237.900 ;
        RECT 821.400 236.400 831.900 237.450 ;
        RECT 826.950 235.950 831.900 236.400 ;
        RECT 833.100 235.950 838.050 238.050 ;
        RECT 826.950 235.800 829.050 235.950 ;
        RECT 823.950 234.450 826.050 235.050 ;
        RECT 817.950 234.000 826.050 234.450 ;
        RECT 818.400 233.400 826.050 234.000 ;
        RECT 823.950 232.950 826.050 233.400 ;
        RECT 838.950 234.450 841.050 235.050 ;
        RECT 853.950 234.450 856.050 235.050 ;
        RECT 838.950 233.400 856.050 234.450 ;
        RECT 838.950 232.950 841.050 233.400 ;
        RECT 853.950 232.950 856.050 233.400 ;
        RECT 841.950 231.450 844.050 232.050 ;
        RECT 766.950 230.400 810.450 231.450 ;
        RECT 812.400 230.400 844.050 231.450 ;
        RECT 766.950 229.950 769.050 230.400 ;
        RECT 418.950 226.950 421.050 227.400 ;
        RECT 463.950 226.950 466.050 227.400 ;
        RECT 10.950 225.450 13.050 226.050 ;
        RECT 46.950 225.450 49.050 226.050 ;
        RECT 88.950 225.450 91.050 226.050 ;
        RECT 10.950 224.400 91.050 225.450 ;
        RECT 10.950 223.950 13.050 224.400 ;
        RECT 46.950 223.950 49.050 224.400 ;
        RECT 88.950 223.950 91.050 224.400 ;
        RECT 232.950 223.950 238.050 226.050 ;
        RECT 277.950 225.450 280.050 226.050 ;
        RECT 307.950 225.450 310.050 226.050 ;
        RECT 277.950 224.400 310.050 225.450 ;
        RECT 277.950 223.950 280.050 224.400 ;
        RECT 307.950 223.950 310.050 224.400 ;
        RECT 346.950 225.450 349.050 226.050 ;
        RECT 406.950 225.450 409.050 226.050 ;
        RECT 430.950 225.450 433.050 226.050 ;
        RECT 346.950 224.400 433.050 225.450 ;
        RECT 346.950 223.950 349.050 224.400 ;
        RECT 406.950 223.950 409.050 224.400 ;
        RECT 430.950 223.950 433.050 224.400 ;
        RECT 481.950 225.450 484.050 226.050 ;
        RECT 499.950 225.450 502.050 226.050 ;
        RECT 481.950 224.400 502.050 225.450 ;
        RECT 481.950 223.950 484.050 224.400 ;
        RECT 499.950 223.950 502.050 224.400 ;
        RECT 514.950 225.450 517.050 226.050 ;
        RECT 529.950 225.450 532.050 226.050 ;
        RECT 589.950 225.600 592.050 227.700 ;
        RECT 610.950 226.500 613.050 228.600 ;
        RECT 697.950 228.450 700.050 229.050 ;
        RECT 715.800 228.450 717.900 229.050 ;
        RECT 697.950 227.400 717.900 228.450 ;
        RECT 697.950 226.950 700.050 227.400 ;
        RECT 715.800 226.950 717.900 227.400 ;
        RECT 719.100 228.450 721.200 229.050 ;
        RECT 802.950 228.450 805.050 229.050 ;
        RECT 719.100 227.400 805.050 228.450 ;
        RECT 809.400 228.450 810.450 230.400 ;
        RECT 841.950 229.950 844.050 230.400 ;
        RECT 823.950 228.450 826.050 229.050 ;
        RECT 809.400 227.400 826.050 228.450 ;
        RECT 719.100 226.950 721.200 227.400 ;
        RECT 802.950 226.950 805.050 227.400 ;
        RECT 823.950 226.950 826.050 227.400 ;
        RECT 830.100 228.450 832.200 229.050 ;
        RECT 847.950 228.450 850.050 229.050 ;
        RECT 830.100 227.400 850.050 228.450 ;
        RECT 830.100 226.950 832.200 227.400 ;
        RECT 847.950 226.950 850.050 227.400 ;
        RECT 514.950 224.400 532.050 225.450 ;
        RECT 514.950 223.950 517.050 224.400 ;
        RECT 529.950 223.950 532.050 224.400 ;
        RECT 622.950 225.450 625.050 226.050 ;
        RECT 640.950 225.450 643.050 226.050 ;
        RECT 622.950 224.400 643.050 225.450 ;
        RECT 622.950 223.950 625.050 224.400 ;
        RECT 640.950 223.950 643.050 224.400 ;
        RECT 664.950 225.450 667.050 226.050 ;
        RECT 700.950 225.450 703.050 226.050 ;
        RECT 664.950 224.400 703.050 225.450 ;
        RECT 664.950 223.950 667.050 224.400 ;
        RECT 700.950 223.950 703.050 224.400 ;
        RECT 769.950 225.450 772.050 226.050 ;
        RECT 790.950 225.450 793.050 226.050 ;
        RECT 769.950 224.400 793.050 225.450 ;
        RECT 800.100 225.000 802.200 226.050 ;
        RECT 769.950 223.950 772.050 224.400 ;
        RECT 790.950 223.950 793.050 224.400 ;
        RECT 799.950 223.950 802.200 225.000 ;
        RECT 835.950 225.450 838.050 226.050 ;
        RECT 841.950 225.450 844.050 226.050 ;
        RECT 835.950 224.400 844.050 225.450 ;
        RECT 835.950 223.950 838.050 224.400 ;
        RECT 841.950 223.950 844.050 224.400 ;
        RECT 799.950 223.050 802.050 223.950 ;
        RECT 220.950 222.450 223.050 223.050 ;
        RECT 295.950 222.450 298.050 223.050 ;
        RECT 331.950 222.450 334.050 223.050 ;
        RECT 220.950 221.400 334.050 222.450 ;
        RECT 220.950 220.950 223.050 221.400 ;
        RECT 295.950 220.950 298.050 221.400 ;
        RECT 331.950 220.950 334.050 221.400 ;
        RECT 379.950 222.450 382.050 223.050 ;
        RECT 448.950 222.450 451.050 223.050 ;
        RECT 379.950 221.400 451.050 222.450 ;
        RECT 379.950 220.950 382.050 221.400 ;
        RECT 448.950 220.950 451.050 221.400 ;
        RECT 469.950 222.450 472.050 223.050 ;
        RECT 568.950 222.450 571.050 223.050 ;
        RECT 619.950 222.450 622.050 223.050 ;
        RECT 469.950 221.400 525.450 222.450 ;
        RECT 469.950 220.950 472.050 221.400 ;
        RECT 166.950 219.450 169.050 220.050 ;
        RECT 181.950 219.450 184.050 220.050 ;
        RECT 268.950 219.450 271.050 220.050 ;
        RECT 166.950 218.400 271.050 219.450 ;
        RECT 166.950 217.950 169.050 218.400 ;
        RECT 181.950 217.950 184.050 218.400 ;
        RECT 268.950 217.950 271.050 218.400 ;
        RECT 382.950 219.450 385.050 220.050 ;
        RECT 466.950 219.450 469.050 220.050 ;
        RECT 382.950 218.400 469.050 219.450 ;
        RECT 382.950 217.950 385.050 218.400 ;
        RECT 466.950 217.950 469.050 218.400 ;
        RECT 472.950 219.450 475.050 220.050 ;
        RECT 508.950 219.450 511.050 220.050 ;
        RECT 472.950 218.400 511.050 219.450 ;
        RECT 524.400 219.450 525.450 221.400 ;
        RECT 568.950 221.400 622.050 222.450 ;
        RECT 568.950 220.950 571.050 221.400 ;
        RECT 619.950 220.950 622.050 221.400 ;
        RECT 634.950 222.450 637.050 223.050 ;
        RECT 646.950 222.450 649.050 223.050 ;
        RECT 634.950 221.400 649.050 222.450 ;
        RECT 634.950 220.950 637.050 221.400 ;
        RECT 646.950 220.950 649.050 221.400 ;
        RECT 658.950 222.450 661.050 223.050 ;
        RECT 706.950 222.450 709.050 223.050 ;
        RECT 658.950 221.400 709.050 222.450 ;
        RECT 658.950 220.950 661.050 221.400 ;
        RECT 706.950 220.950 709.050 221.400 ;
        RECT 736.950 222.450 742.050 223.050 ;
        RECT 757.950 222.450 760.050 223.050 ;
        RECT 736.950 221.400 760.050 222.450 ;
        RECT 736.950 220.950 742.050 221.400 ;
        RECT 757.950 220.950 760.050 221.400 ;
        RECT 772.950 222.450 775.050 223.050 ;
        RECT 796.800 222.450 798.900 223.050 ;
        RECT 772.950 221.400 798.900 222.450 ;
        RECT 799.950 222.000 802.200 223.050 ;
        RECT 844.950 222.450 847.050 223.050 ;
        RECT 772.950 220.950 775.050 221.400 ;
        RECT 796.800 220.950 798.900 221.400 ;
        RECT 800.100 220.950 802.200 222.000 ;
        RECT 803.400 221.400 847.050 222.450 ;
        RECT 652.950 219.450 655.050 220.050 ;
        RECT 524.400 218.400 655.050 219.450 ;
        RECT 472.950 217.950 475.050 218.400 ;
        RECT 508.950 217.950 511.050 218.400 ;
        RECT 652.950 217.950 655.050 218.400 ;
        RECT 697.950 219.450 700.050 220.050 ;
        RECT 742.950 219.450 745.050 220.050 ;
        RECT 697.950 218.400 745.050 219.450 ;
        RECT 697.950 217.950 700.050 218.400 ;
        RECT 742.950 217.950 745.050 218.400 ;
        RECT 784.950 219.450 787.050 220.050 ;
        RECT 803.400 219.450 804.450 221.400 ;
        RECT 844.950 220.950 847.050 221.400 ;
        RECT 850.950 220.950 856.050 223.050 ;
        RECT 817.950 219.450 820.050 220.050 ;
        RECT 784.950 218.400 804.450 219.450 ;
        RECT 806.400 218.400 820.050 219.450 ;
        RECT 784.950 217.950 787.050 218.400 ;
        RECT 127.950 216.450 130.050 217.050 ;
        RECT 92.400 215.400 130.050 216.450 ;
        RECT 67.950 213.450 70.050 214.050 ;
        RECT 92.400 213.450 93.450 215.400 ;
        RECT 127.950 214.950 130.050 215.400 ;
        RECT 178.950 216.450 181.050 217.050 ;
        RECT 211.950 216.450 214.050 217.050 ;
        RECT 349.800 216.450 351.900 217.050 ;
        RECT 178.950 215.400 351.900 216.450 ;
        RECT 178.950 214.950 181.050 215.400 ;
        RECT 211.950 214.950 214.050 215.400 ;
        RECT 349.800 214.950 351.900 215.400 ;
        RECT 353.100 216.450 355.200 217.050 ;
        RECT 418.950 216.450 421.050 217.050 ;
        RECT 353.100 215.400 421.050 216.450 ;
        RECT 353.100 214.950 355.200 215.400 ;
        RECT 418.950 214.950 421.050 215.400 ;
        RECT 517.950 216.450 520.050 217.050 ;
        RECT 598.950 216.450 601.050 217.050 ;
        RECT 517.950 215.400 601.050 216.450 ;
        RECT 517.950 214.950 520.050 215.400 ;
        RECT 598.950 214.950 601.050 215.400 ;
        RECT 640.950 216.450 643.050 217.050 ;
        RECT 649.950 216.450 652.050 217.050 ;
        RECT 640.950 215.400 652.050 216.450 ;
        RECT 640.950 214.950 643.050 215.400 ;
        RECT 649.950 214.950 652.050 215.400 ;
        RECT 688.950 216.450 691.050 217.200 ;
        RECT 703.950 216.450 706.050 217.050 ;
        RECT 688.950 215.400 706.050 216.450 ;
        RECT 688.950 215.100 691.050 215.400 ;
        RECT 703.950 214.950 706.050 215.400 ;
        RECT 736.950 216.450 739.050 217.050 ;
        RECT 766.950 216.450 769.050 217.050 ;
        RECT 736.950 215.400 769.050 216.450 ;
        RECT 736.950 214.950 739.050 215.400 ;
        RECT 766.950 214.950 769.050 215.400 ;
        RECT 796.950 216.450 799.050 217.050 ;
        RECT 806.400 216.450 807.450 218.400 ;
        RECT 817.950 217.950 820.050 218.400 ;
        RECT 796.950 215.400 807.450 216.450 ;
        RECT 811.950 216.450 814.050 217.050 ;
        RECT 832.950 216.450 835.050 217.050 ;
        RECT 811.950 215.400 835.050 216.450 ;
        RECT 796.950 214.950 799.050 215.400 ;
        RECT 811.950 214.950 814.050 215.400 ;
        RECT 832.950 214.950 835.050 215.400 ;
        RECT 67.950 212.400 93.450 213.450 ;
        RECT 103.950 213.450 106.050 214.050 ;
        RECT 136.950 213.450 139.050 214.050 ;
        RECT 184.800 213.450 186.900 214.050 ;
        RECT 103.950 212.400 186.900 213.450 ;
        RECT 67.950 211.950 70.050 212.400 ;
        RECT 103.950 211.950 106.050 212.400 ;
        RECT 136.950 211.950 139.050 212.400 ;
        RECT 184.800 211.950 186.900 212.400 ;
        RECT 188.100 213.450 190.200 214.050 ;
        RECT 229.950 213.450 232.050 214.050 ;
        RECT 188.100 212.400 232.050 213.450 ;
        RECT 188.100 211.950 190.200 212.400 ;
        RECT 229.950 211.950 232.050 212.400 ;
        RECT 358.950 213.450 361.050 214.050 ;
        RECT 367.950 213.450 373.050 214.050 ;
        RECT 358.950 212.400 373.050 213.450 ;
        RECT 358.950 211.950 361.050 212.400 ;
        RECT 367.950 211.950 373.050 212.400 ;
        RECT 439.950 213.450 442.050 214.050 ;
        RECT 511.950 213.450 514.050 213.900 ;
        RECT 544.950 213.450 547.050 214.050 ;
        RECT 439.950 212.400 547.050 213.450 ;
        RECT 439.950 211.950 442.050 212.400 ;
        RECT 511.950 211.800 514.050 212.400 ;
        RECT 544.950 211.950 547.050 212.400 ;
        RECT 613.950 213.450 616.050 214.050 ;
        RECT 655.950 213.450 658.050 214.050 ;
        RECT 613.950 212.400 658.050 213.450 ;
        RECT 613.950 211.950 616.050 212.400 ;
        RECT 655.950 211.950 658.050 212.400 ;
        RECT 688.950 213.450 691.050 213.900 ;
        RECT 727.800 213.450 729.900 214.050 ;
        RECT 688.950 212.400 729.900 213.450 ;
        RECT 688.950 211.800 691.050 212.400 ;
        RECT 727.800 211.950 729.900 212.400 ;
        RECT 731.100 213.450 733.200 214.050 ;
        RECT 739.950 213.450 742.050 214.050 ;
        RECT 731.100 212.400 742.050 213.450 ;
        RECT 731.100 211.950 733.200 212.400 ;
        RECT 739.950 211.950 742.050 212.400 ;
        RECT 751.950 213.450 754.050 214.050 ;
        RECT 790.950 213.450 793.050 214.050 ;
        RECT 751.950 212.400 793.050 213.450 ;
        RECT 751.950 211.950 754.050 212.400 ;
        RECT 790.950 211.950 793.050 212.400 ;
        RECT 808.950 213.450 811.050 214.200 ;
        RECT 841.950 213.450 844.050 214.050 ;
        RECT 808.950 212.400 844.050 213.450 ;
        RECT 808.950 212.100 811.050 212.400 ;
        RECT 841.950 211.950 844.050 212.400 ;
        RECT 94.950 210.450 97.050 211.050 ;
        RECT 139.950 210.450 142.050 211.050 ;
        RECT 94.950 209.400 142.050 210.450 ;
        RECT 94.950 208.950 97.050 209.400 ;
        RECT 139.950 208.950 142.050 209.400 ;
        RECT 190.950 210.450 193.050 211.050 ;
        RECT 226.950 210.450 229.050 211.050 ;
        RECT 190.950 209.400 229.050 210.450 ;
        RECT 190.950 208.950 193.050 209.400 ;
        RECT 226.950 208.950 229.050 209.400 ;
        RECT 349.950 210.450 352.050 211.050 ;
        RECT 364.950 210.450 367.050 211.050 ;
        RECT 349.950 209.400 367.050 210.450 ;
        RECT 619.950 210.450 622.050 211.050 ;
        RECT 670.950 210.450 673.050 211.050 ;
        RECT 619.950 209.400 673.050 210.450 ;
        RECT 349.950 208.950 352.050 209.400 ;
        RECT 364.950 208.950 367.050 209.400 ;
        RECT 34.950 207.450 37.050 208.050 ;
        RECT 85.950 207.450 88.050 208.050 ;
        RECT 151.950 207.450 154.050 208.050 ;
        RECT 34.950 206.400 51.450 207.450 ;
        RECT 34.950 205.950 37.050 206.400 ;
        RECT 50.400 205.050 51.450 206.400 ;
        RECT 85.950 206.400 154.050 207.450 ;
        RECT 85.950 205.950 88.050 206.400 ;
        RECT 151.950 205.950 154.050 206.400 ;
        RECT 259.950 207.450 262.050 208.050 ;
        RECT 274.950 207.450 277.050 208.050 ;
        RECT 259.950 206.400 277.050 207.450 ;
        RECT 259.950 205.950 262.050 206.400 ;
        RECT 274.950 205.950 277.050 206.400 ;
        RECT 304.950 207.450 307.050 208.050 ;
        RECT 358.950 207.450 361.050 208.050 ;
        RECT 304.950 206.400 361.050 207.450 ;
        RECT 304.950 205.950 307.050 206.400 ;
        RECT 358.950 205.950 361.050 206.400 ;
        RECT 391.950 207.450 394.050 208.050 ;
        RECT 442.950 207.450 445.050 208.050 ;
        RECT 391.950 206.400 445.050 207.450 ;
        RECT 502.950 207.300 505.050 209.400 ;
        RECT 619.950 208.950 622.050 209.400 ;
        RECT 670.950 208.950 673.050 209.400 ;
        RECT 682.950 210.450 685.050 211.050 ;
        RECT 724.950 210.450 727.050 211.050 ;
        RECT 682.950 209.400 727.050 210.450 ;
        RECT 682.950 208.950 685.050 209.400 ;
        RECT 724.950 208.950 727.050 209.400 ;
        RECT 742.950 210.450 745.050 211.050 ;
        RECT 766.950 210.450 769.050 211.050 ;
        RECT 742.950 209.400 769.050 210.450 ;
        RECT 742.950 208.950 745.050 209.400 ;
        RECT 766.950 208.950 769.050 209.400 ;
        RECT 808.950 210.450 811.050 210.900 ;
        RECT 814.950 210.450 817.050 211.050 ;
        RECT 808.950 209.400 817.050 210.450 ;
        RECT 808.950 208.800 811.050 209.400 ;
        RECT 814.950 208.950 817.050 209.400 ;
        RECT 826.950 210.450 829.050 211.050 ;
        RECT 856.950 210.450 859.050 211.050 ;
        RECT 826.950 209.400 859.050 210.450 ;
        RECT 826.950 208.950 829.050 209.400 ;
        RECT 856.950 208.950 859.050 209.400 ;
        RECT 391.950 205.950 394.050 206.400 ;
        RECT 442.950 205.950 445.050 206.400 ;
        RECT 46.800 204.450 48.900 205.050 ;
        RECT 32.550 204.000 48.900 204.450 ;
        RECT 31.950 203.400 48.900 204.000 ;
        RECT 31.950 202.050 34.050 203.400 ;
        RECT 46.800 202.950 48.900 203.400 ;
        RECT 50.100 204.450 54.000 205.050 ;
        RECT 76.950 204.450 79.050 205.050 ;
        RECT 50.100 203.400 79.050 204.450 ;
        RECT 50.100 202.950 55.050 203.400 ;
        RECT 76.950 202.950 79.050 203.400 ;
        RECT 118.950 204.450 121.050 205.050 ;
        RECT 118.950 204.000 138.450 204.450 ;
        RECT 118.950 203.400 139.050 204.000 ;
        RECT 118.950 202.950 121.050 203.400 ;
        RECT 28.800 201.450 30.900 202.050 ;
        RECT 11.400 201.000 30.900 201.450 ;
        RECT 31.950 201.000 34.200 202.050 ;
        RECT 10.950 200.400 31.050 201.000 ;
        RECT 10.950 196.950 13.050 200.400 ;
        RECT 28.800 199.950 31.050 200.400 ;
        RECT 32.100 199.950 34.200 201.000 ;
        RECT 40.950 199.950 46.050 202.050 ;
        RECT 52.950 199.950 55.050 202.950 ;
        RECT 61.950 201.450 64.050 202.050 ;
        RECT 73.950 201.450 76.050 202.050 ;
        RECT 61.950 200.400 76.050 201.450 ;
        RECT 61.950 199.950 64.050 200.400 ;
        RECT 73.950 199.950 76.050 200.400 ;
        RECT 16.950 196.050 19.050 199.050 ;
        RECT 28.950 196.950 31.050 199.950 ;
        RECT 34.950 196.950 40.050 199.050 ;
        RECT 46.950 196.950 51.900 199.050 ;
        RECT 53.100 196.950 58.050 199.050 ;
        RECT 64.950 198.450 67.050 199.050 ;
        RECT 76.800 198.450 78.900 199.050 ;
        RECT 64.950 197.400 78.900 198.450 ;
        RECT 64.950 196.950 67.050 197.400 ;
        RECT 76.800 196.950 78.900 197.400 ;
        RECT 80.100 196.950 85.050 199.050 ;
        RECT 94.950 196.950 97.050 202.050 ;
        RECT 136.950 199.950 139.050 203.400 ;
        RECT 145.950 199.950 151.050 202.050 ;
        RECT 175.950 199.950 178.050 205.050 ;
        RECT 181.950 199.950 184.050 205.050 ;
        RECT 217.950 204.450 220.050 205.050 ;
        RECT 316.950 204.450 319.050 205.050 ;
        RECT 331.950 204.450 334.050 205.050 ;
        RECT 349.950 204.450 352.050 205.050 ;
        RECT 217.950 203.400 352.050 204.450 ;
        RECT 217.950 202.950 220.050 203.400 ;
        RECT 316.950 202.950 319.050 203.400 ;
        RECT 331.950 202.950 334.050 203.400 ;
        RECT 349.950 202.950 352.050 203.400 ;
        RECT 367.950 204.450 370.050 205.050 ;
        RECT 454.950 204.450 457.050 205.050 ;
        RECT 478.950 204.450 481.050 205.050 ;
        RECT 490.950 204.450 493.050 205.050 ;
        RECT 367.950 204.000 381.450 204.450 ;
        RECT 367.950 203.400 382.050 204.000 ;
        RECT 367.950 202.950 370.050 203.400 ;
        RECT 190.950 201.450 193.050 202.050 ;
        RECT 196.950 201.450 199.050 202.050 ;
        RECT 190.950 200.400 199.050 201.450 ;
        RECT 190.950 199.950 193.050 200.400 ;
        RECT 196.950 199.950 199.050 200.400 ;
        RECT 202.950 201.450 205.050 202.050 ;
        RECT 208.950 201.450 214.050 202.050 ;
        RECT 202.950 200.400 214.050 201.450 ;
        RECT 202.950 199.950 205.050 200.400 ;
        RECT 208.950 199.950 214.050 200.400 ;
        RECT 229.950 199.950 235.050 202.050 ;
        RECT 238.950 201.450 241.050 202.050 ;
        RECT 262.950 201.450 265.050 202.050 ;
        RECT 310.950 201.450 313.050 202.050 ;
        RECT 238.950 200.400 265.050 201.450 ;
        RECT 299.250 201.000 313.050 201.450 ;
        RECT 238.950 199.950 241.050 200.400 ;
        RECT 262.950 199.950 265.050 200.400 ;
        RECT 298.950 200.400 313.050 201.000 ;
        RECT 298.950 199.050 301.050 200.400 ;
        RECT 310.950 199.950 313.050 200.400 ;
        RECT 337.950 199.950 343.050 202.050 ;
        RECT 352.950 201.450 355.050 202.200 ;
        RECT 361.800 201.450 363.900 202.050 ;
        RECT 352.950 200.400 363.900 201.450 ;
        RECT 352.950 200.100 355.050 200.400 ;
        RECT 361.800 199.950 363.900 200.400 ;
        RECT 365.100 201.450 367.200 202.050 ;
        RECT 373.950 201.450 376.050 202.050 ;
        RECT 365.100 200.400 376.050 201.450 ;
        RECT 365.100 199.950 367.200 200.400 ;
        RECT 373.950 199.950 376.050 200.400 ;
        RECT 379.950 199.950 382.050 203.400 ;
        RECT 454.950 203.400 493.050 204.450 ;
        RECT 503.850 203.700 505.050 207.300 ;
        RECT 523.950 206.400 526.050 208.500 ;
        RECT 592.950 207.450 595.050 208.050 ;
        RECT 601.950 207.450 604.050 208.050 ;
        RECT 592.950 206.400 604.050 207.450 ;
        RECT 454.950 202.950 457.050 203.400 ;
        RECT 478.950 202.950 481.050 203.400 ;
        RECT 490.950 202.950 493.050 203.400 ;
        RECT 433.950 201.450 436.050 202.050 ;
        RECT 438.000 201.450 442.050 202.050 ;
        RECT 502.950 201.600 505.050 203.700 ;
        RECT 392.400 201.000 411.300 201.450 ;
        RECT 416.550 201.000 436.050 201.450 ;
        RECT 437.400 201.000 442.050 201.450 ;
        RECT 392.400 200.400 412.050 201.000 ;
        RECT 392.400 199.050 393.450 200.400 ;
        RECT 409.950 199.050 412.050 200.400 ;
        RECT 415.950 200.400 436.050 201.000 ;
        RECT 415.950 199.050 418.050 200.400 ;
        RECT 433.950 199.950 436.050 200.400 ;
        RECT 436.950 199.950 442.050 201.000 ;
        RECT 100.950 196.050 103.050 199.050 ;
        RECT 115.950 196.950 120.900 199.050 ;
        RECT 122.100 196.950 127.050 199.050 ;
        RECT 130.950 196.950 136.050 199.050 ;
        RECT 13.800 195.000 15.900 196.050 ;
        RECT 16.800 195.000 19.050 196.050 ;
        RECT 13.800 193.950 16.050 195.000 ;
        RECT 16.800 193.950 18.900 195.000 ;
        RECT 20.100 193.950 25.050 196.050 ;
        RECT 13.950 190.950 16.050 193.950 ;
        RECT 79.950 192.450 82.050 196.050 ;
        RECT 97.800 195.000 99.900 196.050 ;
        RECT 100.800 195.000 103.050 196.050 ;
        RECT 104.100 195.450 106.200 196.050 ;
        RECT 112.950 195.450 115.050 196.050 ;
        RECT 97.800 193.950 100.050 195.000 ;
        RECT 100.800 193.950 102.900 195.000 ;
        RECT 104.100 194.400 115.050 195.450 ;
        RECT 104.100 193.950 106.200 194.400 ;
        RECT 112.950 193.950 115.050 194.400 ;
        RECT 94.950 192.450 97.050 193.050 ;
        RECT 79.950 192.000 97.050 192.450 ;
        RECT 97.950 192.450 100.050 193.950 ;
        RECT 118.950 192.450 121.050 196.050 ;
        RECT 124.950 193.950 130.050 196.050 ;
        RECT 139.950 195.450 142.050 199.050 ;
        RECT 160.950 198.450 163.050 199.050 ;
        RECT 175.800 198.450 177.900 199.050 ;
        RECT 160.950 197.400 177.900 198.450 ;
        RECT 160.950 196.950 163.050 197.400 ;
        RECT 175.800 196.950 177.900 197.400 ;
        RECT 179.100 196.950 183.900 199.050 ;
        RECT 185.100 198.450 187.200 199.050 ;
        RECT 199.950 198.450 202.050 199.050 ;
        RECT 185.100 197.400 202.050 198.450 ;
        RECT 185.100 196.950 187.200 197.400 ;
        RECT 199.950 196.950 202.050 197.400 ;
        RECT 214.950 198.450 217.050 199.050 ;
        RECT 226.950 198.450 229.050 199.050 ;
        RECT 214.950 197.400 229.050 198.450 ;
        RECT 214.950 196.950 217.050 197.400 ;
        RECT 226.950 196.950 229.050 197.400 ;
        RECT 235.950 198.450 238.050 199.050 ;
        RECT 244.950 198.450 247.050 199.050 ;
        RECT 235.950 197.400 247.050 198.450 ;
        RECT 235.950 196.950 238.050 197.400 ;
        RECT 244.950 196.950 247.050 197.400 ;
        RECT 256.950 198.450 259.050 199.050 ;
        RECT 268.950 198.450 271.050 199.050 ;
        RECT 256.950 197.400 271.050 198.450 ;
        RECT 256.950 196.950 259.050 197.400 ;
        RECT 268.950 196.950 271.050 197.400 ;
        RECT 286.950 198.450 289.050 199.050 ;
        RECT 286.950 198.000 297.450 198.450 ;
        RECT 298.800 198.000 301.050 199.050 ;
        RECT 286.950 197.400 298.050 198.000 ;
        RECT 286.950 196.950 289.050 197.400 ;
        RECT 154.950 195.450 157.050 196.050 ;
        RECT 139.950 195.000 157.050 195.450 ;
        RECT 140.400 194.400 157.050 195.000 ;
        RECT 154.950 193.950 157.050 194.400 ;
        RECT 166.950 193.950 172.050 196.050 ;
        RECT 252.000 195.900 255.000 196.050 ;
        RECT 250.950 193.950 256.050 195.900 ;
        RECT 295.950 193.950 298.050 197.400 ;
        RECT 298.800 196.950 300.900 198.000 ;
        RECT 302.100 196.950 307.050 199.050 ;
        RECT 322.950 198.450 325.050 199.050 ;
        RECT 331.950 198.450 334.050 199.050 ;
        RECT 352.950 198.450 355.050 198.900 ;
        RECT 322.950 197.400 355.050 198.450 ;
        RECT 322.950 196.950 325.050 197.400 ;
        RECT 331.950 196.950 334.050 197.400 ;
        RECT 352.950 196.800 355.050 197.400 ;
        RECT 358.950 196.950 364.050 199.050 ;
        RECT 367.950 196.950 373.050 199.050 ;
        RECT 250.950 193.800 253.050 193.950 ;
        RECT 253.950 193.800 256.050 193.950 ;
        RECT 160.950 192.450 163.050 193.050 ;
        RECT 97.950 192.000 117.450 192.450 ;
        RECT 118.950 192.000 163.050 192.450 ;
        RECT 80.400 191.400 97.050 192.000 ;
        RECT 98.400 191.400 117.450 192.000 ;
        RECT 119.400 191.400 163.050 192.000 ;
        RECT 94.950 190.950 97.050 191.400 ;
        RECT 31.950 189.450 34.050 190.050 ;
        RECT 82.950 189.450 85.050 190.050 ;
        RECT 31.950 188.400 85.050 189.450 ;
        RECT 116.400 189.450 117.450 191.400 ;
        RECT 160.950 190.950 163.050 191.400 ;
        RECT 259.800 192.000 261.900 193.050 ;
        RECT 263.100 192.450 265.200 193.050 ;
        RECT 280.950 192.450 283.050 193.050 ;
        RECT 259.800 190.950 262.050 192.000 ;
        RECT 263.100 191.400 283.050 192.450 ;
        RECT 301.950 192.450 304.050 196.050 ;
        RECT 310.950 192.450 313.050 193.050 ;
        RECT 301.950 192.000 313.050 192.450 ;
        RECT 302.400 191.400 313.050 192.000 ;
        RECT 263.100 190.950 265.200 191.400 ;
        RECT 280.950 190.950 283.050 191.400 ;
        RECT 310.950 190.950 313.050 191.400 ;
        RECT 322.950 190.950 328.050 193.050 ;
        RECT 334.950 190.950 337.050 196.050 ;
        RECT 343.950 193.950 349.050 196.050 ;
        RECT 376.950 193.950 379.050 199.050 ;
        RECT 391.950 193.950 394.050 199.050 ;
        RECT 397.950 195.450 400.050 199.050 ;
        RECT 409.800 198.000 412.050 199.050 ;
        RECT 412.800 198.000 414.900 199.050 ;
        RECT 415.950 198.000 418.200 199.050 ;
        RECT 409.800 196.950 411.900 198.000 ;
        RECT 412.800 196.950 415.050 198.000 ;
        RECT 416.100 196.950 418.200 198.000 ;
        RECT 436.950 196.950 439.050 199.950 ;
        RECT 451.950 198.450 454.050 199.050 ;
        RECT 440.400 197.400 454.050 198.450 ;
        RECT 412.950 196.050 415.050 196.950 ;
        RECT 406.950 195.450 409.050 196.050 ;
        RECT 397.950 194.400 409.050 195.450 ;
        RECT 397.950 193.950 400.050 194.400 ;
        RECT 406.950 193.950 409.050 194.400 ;
        RECT 412.800 195.000 415.050 196.050 ;
        RECT 412.800 193.950 414.900 195.000 ;
        RECT 394.950 192.450 397.050 193.050 ;
        RECT 394.950 191.400 411.450 192.450 ;
        RECT 394.950 190.950 397.050 191.400 ;
        RECT 154.950 189.450 157.050 190.050 ;
        RECT 116.400 188.400 157.050 189.450 ;
        RECT 31.950 187.950 34.050 188.400 ;
        RECT 82.950 187.950 85.050 188.400 ;
        RECT 154.950 187.950 157.050 188.400 ;
        RECT 184.950 187.950 190.050 190.050 ;
        RECT 250.950 189.450 253.050 190.050 ;
        RECT 259.950 189.450 262.050 190.950 ;
        RECT 250.950 189.000 262.050 189.450 ;
        RECT 289.950 189.450 292.050 190.050 ;
        RECT 334.950 189.450 337.050 190.050 ;
        RECT 373.950 189.450 376.050 190.050 ;
        RECT 250.950 188.400 261.300 189.000 ;
        RECT 289.950 188.400 376.050 189.450 ;
        RECT 410.400 189.450 411.450 191.400 ;
        RECT 418.950 190.950 421.050 196.050 ;
        RECT 433.950 195.450 436.050 196.050 ;
        RECT 440.400 195.450 441.450 197.400 ;
        RECT 451.950 196.950 454.050 197.400 ;
        RECT 469.800 196.950 471.900 199.050 ;
        RECT 472.800 198.000 474.900 199.050 ;
        RECT 472.800 196.950 475.050 198.000 ;
        RECT 476.100 196.950 481.050 199.050 ;
        RECT 487.950 198.450 490.050 199.050 ;
        RECT 482.400 197.400 490.050 198.450 ;
        RECT 433.950 194.400 441.450 195.450 ;
        RECT 433.950 193.950 436.050 194.400 ;
        RECT 442.950 193.950 448.050 196.050 ;
        RECT 451.950 195.450 454.050 196.050 ;
        RECT 457.950 195.450 460.050 196.050 ;
        RECT 451.950 194.400 460.050 195.450 ;
        RECT 451.950 193.950 454.050 194.400 ;
        RECT 457.950 193.950 460.050 194.400 ;
        RECT 463.950 193.950 469.050 196.050 ;
        RECT 427.950 189.450 430.050 190.050 ;
        RECT 410.400 188.400 430.050 189.450 ;
        RECT 448.950 189.450 451.050 193.050 ;
        RECT 470.250 192.450 471.300 196.950 ;
        RECT 472.950 196.050 475.050 196.950 ;
        RECT 482.400 196.050 483.450 197.400 ;
        RECT 487.950 196.950 490.050 197.400 ;
        RECT 472.800 195.000 475.050 196.050 ;
        RECT 472.800 193.950 474.900 195.000 ;
        RECT 478.950 194.400 483.450 196.050 ;
        RECT 478.950 193.950 483.000 194.400 ;
        RECT 484.950 192.450 487.050 193.050 ;
        RECT 470.250 191.400 487.050 192.450 ;
        RECT 484.950 190.950 487.050 191.400 ;
        RECT 493.950 192.450 499.050 193.050 ;
        RECT 499.950 192.450 502.050 196.050 ;
        RECT 493.950 192.000 502.050 192.450 ;
        RECT 493.950 191.400 501.450 192.000 ;
        RECT 493.950 190.950 499.050 191.400 ;
        RECT 457.950 189.450 460.050 190.050 ;
        RECT 503.850 189.600 505.050 201.600 ;
        RECT 511.950 193.950 516.900 196.050 ;
        RECT 518.100 195.000 520.200 196.050 ;
        RECT 517.950 193.950 520.200 195.000 ;
        RECT 508.950 192.450 511.050 193.050 ;
        RECT 517.950 192.450 520.050 193.950 ;
        RECT 508.950 192.000 520.050 192.450 ;
        RECT 508.950 191.400 519.600 192.000 ;
        RECT 508.950 190.950 511.050 191.400 ;
        RECT 524.100 189.600 525.300 206.400 ;
        RECT 592.950 205.950 595.050 206.400 ;
        RECT 601.950 205.950 604.050 206.400 ;
        RECT 694.950 207.450 697.050 208.050 ;
        RECT 718.950 207.450 721.050 208.050 ;
        RECT 694.950 206.400 721.050 207.450 ;
        RECT 694.950 205.950 697.050 206.400 ;
        RECT 718.950 205.950 721.050 206.400 ;
        RECT 733.950 207.450 736.050 208.050 ;
        RECT 745.950 207.450 748.050 208.050 ;
        RECT 733.950 206.400 748.050 207.450 ;
        RECT 733.950 205.950 736.050 206.400 ;
        RECT 745.950 205.950 748.050 206.400 ;
        RECT 763.950 207.450 766.050 208.050 ;
        RECT 775.950 207.450 778.050 208.050 ;
        RECT 763.950 206.400 778.050 207.450 ;
        RECT 763.950 205.950 766.050 206.400 ;
        RECT 775.950 205.950 778.050 206.400 ;
        RECT 823.950 207.450 826.050 208.050 ;
        RECT 823.950 206.400 837.450 207.450 ;
        RECT 823.950 205.950 826.050 206.400 ;
        RECT 541.950 204.450 544.050 205.050 ;
        RECT 583.950 204.450 586.050 205.050 ;
        RECT 541.950 203.400 586.050 204.450 ;
        RECT 541.950 202.950 544.050 203.400 ;
        RECT 583.950 202.950 586.050 203.400 ;
        RECT 595.950 204.450 598.050 205.050 ;
        RECT 640.950 204.450 643.050 205.050 ;
        RECT 724.950 204.450 727.050 205.050 ;
        RECT 730.950 204.450 733.050 205.050 ;
        RECT 595.950 203.400 643.050 204.450 ;
        RECT 644.400 204.000 733.050 204.450 ;
        RECT 595.950 202.950 598.050 203.400 ;
        RECT 640.950 202.950 643.050 203.400 ;
        RECT 643.950 203.400 733.050 204.000 ;
        RECT 544.950 198.450 547.050 199.050 ;
        RECT 559.950 198.450 562.050 199.050 ;
        RECT 544.950 197.400 562.050 198.450 ;
        RECT 544.950 196.950 547.050 197.400 ;
        RECT 559.950 196.950 562.050 197.400 ;
        RECT 565.950 196.950 570.900 199.050 ;
        RECT 572.100 198.450 574.200 199.050 ;
        RECT 577.950 198.450 580.050 199.050 ;
        RECT 572.100 197.400 580.050 198.450 ;
        RECT 572.100 196.950 574.200 197.400 ;
        RECT 577.950 196.950 580.050 197.400 ;
        RECT 583.950 196.950 589.050 199.050 ;
        RECT 619.950 196.950 622.050 202.050 ;
        RECT 631.950 199.950 637.050 202.050 ;
        RECT 643.950 199.950 646.050 203.400 ;
        RECT 724.950 202.950 727.050 203.400 ;
        RECT 730.950 202.950 733.050 203.400 ;
        RECT 742.950 202.950 748.050 205.050 ;
        RECT 760.950 204.450 763.050 205.050 ;
        RECT 787.950 204.450 790.050 205.050 ;
        RECT 817.950 204.450 820.050 205.050 ;
        RECT 831.000 204.450 835.050 205.050 ;
        RECT 760.950 203.400 790.050 204.450 ;
        RECT 794.400 204.000 820.050 204.450 ;
        RECT 830.400 204.000 835.050 204.450 ;
        RECT 760.950 202.950 763.050 203.400 ;
        RECT 787.950 202.950 790.050 203.400 ;
        RECT 793.950 203.400 820.050 204.000 ;
        RECT 652.950 199.950 658.050 202.050 ;
        RECT 661.950 201.450 664.050 202.050 ;
        RECT 667.950 201.450 670.050 202.050 ;
        RECT 681.000 201.450 685.050 202.050 ;
        RECT 661.950 200.400 670.050 201.450 ;
        RECT 661.950 199.950 664.050 200.400 ;
        RECT 667.950 199.950 670.050 200.400 ;
        RECT 680.400 199.950 685.050 201.450 ;
        RECT 631.950 198.450 634.050 199.050 ;
        RECT 640.950 198.450 643.050 199.050 ;
        RECT 631.950 197.400 643.050 198.450 ;
        RECT 631.950 196.950 634.050 197.400 ;
        RECT 640.950 196.950 643.050 197.400 ;
        RECT 646.950 198.450 649.050 199.050 ;
        RECT 653.400 198.450 654.450 199.950 ;
        RECT 646.950 197.400 654.450 198.450 ;
        RECT 658.950 198.450 661.050 199.050 ;
        RECT 670.950 198.450 673.050 199.050 ;
        RECT 658.950 197.400 673.050 198.450 ;
        RECT 646.950 196.950 649.050 197.400 ;
        RECT 658.950 196.950 661.050 197.400 ;
        RECT 670.950 196.950 673.050 197.400 ;
        RECT 680.400 196.050 681.450 199.950 ;
        RECT 694.950 196.950 697.050 202.050 ;
        RECT 745.950 201.450 748.050 202.050 ;
        RECT 751.950 201.450 754.050 202.050 ;
        RECT 763.950 201.450 766.050 202.050 ;
        RECT 745.950 200.400 754.050 201.450 ;
        RECT 758.400 201.000 766.050 201.450 ;
        RECT 745.950 199.950 748.050 200.400 ;
        RECT 751.950 199.950 754.050 200.400 ;
        RECT 757.950 200.400 766.050 201.000 ;
        RECT 718.800 199.050 720.900 199.200 ;
        RECT 700.950 198.450 703.050 199.050 ;
        RECT 706.950 198.450 709.050 199.050 ;
        RECT 700.950 197.400 709.050 198.450 ;
        RECT 700.950 196.950 703.050 197.400 ;
        RECT 706.950 196.950 709.050 197.400 ;
        RECT 715.950 197.100 720.900 199.050 ;
        RECT 715.950 196.950 720.000 197.100 ;
        RECT 722.100 196.950 727.050 199.050 ;
        RECT 739.950 198.450 745.050 199.050 ;
        RECT 751.950 198.450 754.050 199.050 ;
        RECT 739.950 197.400 754.050 198.450 ;
        RECT 739.950 196.950 745.050 197.400 ;
        RECT 751.950 196.950 754.050 197.400 ;
        RECT 757.950 196.950 760.050 200.400 ;
        RECT 763.950 199.950 766.050 200.400 ;
        RECT 776.250 200.400 786.450 201.450 ;
        RECT 553.950 193.950 559.050 196.050 ;
        RECT 562.950 192.450 565.050 196.050 ;
        RECT 577.950 193.950 583.050 196.050 ;
        RECT 571.950 192.450 574.050 193.050 ;
        RECT 562.950 191.400 574.050 192.450 ;
        RECT 586.950 192.450 589.050 196.050 ;
        RECT 595.950 193.950 601.050 196.050 ;
        RECT 604.950 195.450 607.050 196.050 ;
        RECT 619.950 195.450 622.050 196.050 ;
        RECT 604.950 194.400 622.050 195.450 ;
        RECT 604.950 193.950 607.050 194.400 ;
        RECT 619.950 193.950 622.050 194.400 ;
        RECT 625.950 195.450 628.050 196.050 ;
        RECT 640.950 195.450 643.050 196.050 ;
        RECT 625.950 194.400 643.050 195.450 ;
        RECT 625.950 193.950 628.050 194.400 ;
        RECT 640.950 193.950 643.050 194.400 ;
        RECT 661.950 195.450 664.050 196.050 ;
        RECT 673.950 195.450 676.050 196.050 ;
        RECT 661.950 194.400 676.050 195.450 ;
        RECT 661.950 193.950 664.050 194.400 ;
        RECT 673.950 193.950 676.050 194.400 ;
        RECT 679.950 193.950 682.050 196.050 ;
        RECT 688.950 193.950 693.900 196.050 ;
        RECT 695.100 193.950 700.050 196.050 ;
        RECT 707.400 195.450 708.450 196.950 ;
        RECT 776.250 196.050 777.300 200.400 ;
        RECT 785.400 198.450 786.450 200.400 ;
        RECT 793.950 199.950 796.050 203.400 ;
        RECT 817.950 202.950 820.050 203.400 ;
        RECT 829.950 202.950 835.050 204.000 ;
        RECT 799.950 201.450 802.050 202.050 ;
        RECT 811.950 201.450 814.050 202.050 ;
        RECT 799.950 200.400 814.050 201.450 ;
        RECT 799.950 199.950 802.050 200.400 ;
        RECT 811.950 199.950 814.050 200.400 ;
        RECT 829.950 199.950 832.050 202.950 ;
        RECT 836.400 202.050 837.450 206.400 ;
        RECT 835.950 199.950 838.050 202.050 ;
        RECT 796.950 198.450 799.050 199.050 ;
        RECT 814.800 198.450 816.900 199.050 ;
        RECT 785.400 197.400 799.050 198.450 ;
        RECT 796.950 196.950 799.050 197.400 ;
        RECT 803.400 197.400 816.900 198.450 ;
        RECT 712.950 195.450 715.050 196.050 ;
        RECT 707.400 194.400 715.050 195.450 ;
        RECT 712.950 193.950 715.050 194.400 ;
        RECT 718.950 193.950 724.050 196.050 ;
        RECT 601.950 192.450 604.050 193.050 ;
        RECT 586.950 192.000 604.050 192.450 ;
        RECT 587.400 191.400 604.050 192.000 ;
        RECT 562.950 190.950 565.050 191.400 ;
        RECT 571.950 190.950 574.050 191.400 ;
        RECT 601.950 190.950 604.050 191.400 ;
        RECT 646.950 192.450 649.050 193.050 ;
        RECT 655.950 192.450 658.050 193.050 ;
        RECT 646.950 191.400 658.050 192.450 ;
        RECT 646.950 190.950 649.050 191.400 ;
        RECT 655.950 190.950 658.050 191.400 ;
        RECT 676.950 190.950 681.900 193.050 ;
        RECT 683.100 192.450 685.200 193.050 ;
        RECT 691.950 192.450 694.050 193.050 ;
        RECT 683.100 191.400 694.050 192.450 ;
        RECT 683.100 190.950 685.200 191.400 ;
        RECT 691.950 190.950 694.050 191.400 ;
        RECT 697.950 192.450 700.050 193.050 ;
        RECT 724.950 192.450 727.050 193.050 ;
        RECT 697.950 191.400 727.050 192.450 ;
        RECT 697.950 190.950 700.050 191.400 ;
        RECT 724.950 190.950 727.050 191.400 ;
        RECT 733.950 190.950 736.050 196.050 ;
        RECT 739.950 195.450 742.050 196.050 ;
        RECT 748.950 195.450 751.050 196.050 ;
        RECT 739.950 194.400 751.050 195.450 ;
        RECT 739.950 193.950 742.050 194.400 ;
        RECT 748.950 193.950 751.050 194.400 ;
        RECT 754.950 192.450 757.050 196.050 ;
        RECT 760.950 195.450 763.050 196.050 ;
        RECT 772.800 195.450 774.900 196.050 ;
        RECT 760.950 194.400 774.900 195.450 ;
        RECT 760.950 193.950 763.050 194.400 ;
        RECT 772.800 193.950 774.900 194.400 ;
        RECT 775.800 193.950 777.900 196.050 ;
        RECT 779.100 193.950 784.050 196.050 ;
        RECT 796.950 195.450 799.050 196.050 ;
        RECT 803.400 195.450 804.450 197.400 ;
        RECT 814.800 196.950 816.900 197.400 ;
        RECT 818.100 198.450 823.050 199.050 ;
        RECT 832.950 198.450 835.050 199.050 ;
        RECT 847.950 198.450 850.050 199.050 ;
        RECT 818.100 197.400 835.050 198.450 ;
        RECT 818.100 196.950 823.050 197.400 ;
        RECT 832.950 196.950 835.050 197.400 ;
        RECT 839.400 197.400 850.050 198.450 ;
        RECT 796.950 194.400 804.450 195.450 ;
        RECT 796.950 193.950 799.050 194.400 ;
        RECT 805.950 193.950 810.900 196.050 ;
        RECT 812.100 195.450 814.200 196.050 ;
        RECT 817.950 195.450 820.050 196.050 ;
        RECT 839.400 195.450 840.450 197.400 ;
        RECT 847.950 196.950 850.050 197.400 ;
        RECT 812.100 194.400 840.450 195.450 ;
        RECT 812.100 193.950 814.200 194.400 ;
        RECT 817.950 193.950 820.050 194.400 ;
        RECT 769.950 192.450 772.050 193.050 ;
        RECT 754.950 192.000 772.050 192.450 ;
        RECT 755.400 191.400 772.050 192.000 ;
        RECT 769.950 190.950 772.050 191.400 ;
        RECT 778.950 192.450 781.050 193.050 ;
        RECT 847.950 192.450 850.050 193.050 ;
        RECT 853.950 192.450 856.050 193.050 ;
        RECT 778.950 191.400 816.450 192.450 ;
        RECT 778.950 190.950 781.050 191.400 ;
        RECT 448.950 189.000 460.050 189.450 ;
        RECT 449.400 188.400 460.050 189.000 ;
        RECT 250.950 187.950 253.050 188.400 ;
        RECT 289.950 187.950 292.050 188.400 ;
        RECT 334.950 187.950 337.050 188.400 ;
        RECT 373.950 187.950 376.050 188.400 ;
        RECT 427.950 187.950 430.050 188.400 ;
        RECT 457.950 187.950 460.050 188.400 ;
        RECT 4.950 186.450 7.050 187.050 ;
        RECT 52.950 186.450 55.050 187.050 ;
        RECT 4.950 185.400 55.050 186.450 ;
        RECT 83.400 186.450 84.450 187.950 ;
        RECT 502.950 187.500 505.050 189.600 ;
        RECT 523.950 187.500 526.050 189.600 ;
        RECT 685.950 189.450 688.050 190.200 ;
        RECT 736.950 189.450 739.050 190.050 ;
        RECT 685.950 188.400 739.050 189.450 ;
        RECT 685.950 188.100 688.050 188.400 ;
        RECT 736.950 187.950 739.050 188.400 ;
        RECT 751.950 189.450 754.050 190.200 ;
        RECT 763.950 189.450 766.050 190.050 ;
        RECT 778.950 189.450 781.050 190.050 ;
        RECT 793.950 189.450 796.050 190.050 ;
        RECT 751.950 188.400 796.050 189.450 ;
        RECT 815.400 189.450 816.450 191.400 ;
        RECT 847.950 191.400 856.050 192.450 ;
        RECT 847.950 190.950 850.050 191.400 ;
        RECT 853.950 190.950 856.050 191.400 ;
        RECT 820.950 189.450 823.050 190.050 ;
        RECT 815.400 188.400 823.050 189.450 ;
        RECT 751.950 188.100 754.050 188.400 ;
        RECT 763.950 187.950 766.050 188.400 ;
        RECT 778.950 187.950 781.050 188.400 ;
        RECT 793.950 187.950 796.050 188.400 ;
        RECT 820.950 187.950 823.050 188.400 ;
        RECT 133.950 186.450 136.050 187.050 ;
        RECT 83.400 185.400 136.050 186.450 ;
        RECT 4.950 184.950 7.050 185.400 ;
        RECT 52.950 184.950 55.050 185.400 ;
        RECT 133.950 184.950 136.050 185.400 ;
        RECT 160.950 186.450 163.050 187.050 ;
        RECT 259.950 186.450 262.050 187.050 ;
        RECT 268.800 186.450 270.900 187.050 ;
        RECT 160.950 185.400 270.900 186.450 ;
        RECT 160.950 184.950 163.050 185.400 ;
        RECT 259.950 184.950 262.050 185.400 ;
        RECT 268.800 184.950 270.900 185.400 ;
        RECT 272.100 186.450 274.200 187.050 ;
        RECT 337.950 186.450 340.050 187.050 ;
        RECT 272.100 185.400 340.050 186.450 ;
        RECT 272.100 184.950 274.200 185.400 ;
        RECT 337.950 184.950 340.050 185.400 ;
        RECT 343.950 186.450 346.050 187.050 ;
        RECT 355.800 186.450 357.900 187.050 ;
        RECT 343.950 185.400 357.900 186.450 ;
        RECT 343.950 184.950 346.050 185.400 ;
        RECT 355.800 184.950 357.900 185.400 ;
        RECT 359.100 186.450 361.200 187.050 ;
        RECT 397.950 186.450 400.050 187.050 ;
        RECT 359.100 185.400 400.050 186.450 ;
        RECT 359.100 184.950 361.200 185.400 ;
        RECT 397.950 184.950 400.050 185.400 ;
        RECT 412.950 186.450 415.050 187.050 ;
        RECT 442.950 186.450 445.050 187.050 ;
        RECT 412.950 185.400 445.050 186.450 ;
        RECT 412.950 184.950 415.050 185.400 ;
        RECT 442.950 184.950 445.050 185.400 ;
        RECT 586.950 186.450 589.050 187.050 ;
        RECT 610.950 186.450 613.050 187.050 ;
        RECT 685.950 186.450 688.050 186.900 ;
        RECT 586.950 185.400 688.050 186.450 ;
        RECT 586.950 184.950 589.050 185.400 ;
        RECT 610.950 184.950 613.050 185.400 ;
        RECT 685.950 184.800 688.050 185.400 ;
        RECT 712.950 186.450 715.050 187.050 ;
        RECT 733.950 186.450 736.050 187.050 ;
        RECT 712.950 185.400 736.050 186.450 ;
        RECT 712.950 184.950 715.050 185.400 ;
        RECT 733.950 184.950 736.050 185.400 ;
        RECT 742.950 186.450 745.050 187.050 ;
        RECT 751.950 186.450 754.050 186.900 ;
        RECT 742.950 185.400 754.050 186.450 ;
        RECT 742.950 184.950 745.050 185.400 ;
        RECT 751.950 184.800 754.050 185.400 ;
        RECT 844.950 186.450 847.050 187.050 ;
        RECT 850.950 186.450 853.050 187.050 ;
        RECT 844.950 185.400 853.050 186.450 ;
        RECT 844.950 184.950 847.050 185.400 ;
        RECT 850.950 184.950 853.050 185.400 ;
        RECT 100.950 183.450 103.050 184.050 ;
        RECT 124.800 183.450 126.900 184.050 ;
        RECT 100.950 182.400 126.900 183.450 ;
        RECT 100.950 181.950 103.050 182.400 ;
        RECT 124.800 181.950 126.900 182.400 ;
        RECT 128.100 183.450 130.200 184.050 ;
        RECT 181.950 183.450 184.050 184.050 ;
        RECT 128.100 182.400 184.050 183.450 ;
        RECT 128.100 181.950 130.200 182.400 ;
        RECT 181.950 181.950 184.050 182.400 ;
        RECT 193.950 183.450 196.050 184.050 ;
        RECT 295.950 183.450 298.050 184.050 ;
        RECT 193.950 182.400 298.050 183.450 ;
        RECT 193.950 181.950 196.050 182.400 ;
        RECT 295.950 181.950 298.050 182.400 ;
        RECT 352.950 183.450 355.050 184.050 ;
        RECT 382.950 183.450 385.050 184.050 ;
        RECT 352.950 182.400 385.050 183.450 ;
        RECT 352.950 181.950 355.050 182.400 ;
        RECT 382.950 181.950 385.050 182.400 ;
        RECT 406.950 183.450 409.050 184.050 ;
        RECT 505.950 183.450 508.050 184.050 ;
        RECT 517.950 183.450 520.050 184.200 ;
        RECT 556.950 183.450 559.050 184.050 ;
        RECT 631.950 183.450 634.050 184.050 ;
        RECT 406.950 182.400 435.450 183.450 ;
        RECT 406.950 181.950 409.050 182.400 ;
        RECT 13.950 180.450 16.050 181.050 ;
        RECT 82.950 180.450 85.050 181.050 ;
        RECT 13.950 179.400 85.050 180.450 ;
        RECT 13.950 178.950 16.050 179.400 ;
        RECT 82.950 178.950 85.050 179.400 ;
        RECT 187.950 180.450 190.050 181.050 ;
        RECT 235.950 180.450 238.050 181.200 ;
        RECT 434.400 181.050 435.450 182.400 ;
        RECT 505.950 182.400 555.450 183.450 ;
        RECT 505.950 181.950 508.050 182.400 ;
        RECT 517.950 182.100 520.050 182.400 ;
        RECT 187.950 179.400 238.050 180.450 ;
        RECT 187.950 178.950 190.050 179.400 ;
        RECT 235.950 179.100 238.050 179.400 ;
        RECT 349.950 180.450 352.050 181.050 ;
        RECT 412.950 180.450 415.050 181.050 ;
        RECT 349.950 179.400 415.050 180.450 ;
        RECT 349.950 178.950 352.050 179.400 ;
        RECT 412.950 178.950 415.050 179.400 ;
        RECT 433.950 180.450 436.050 181.050 ;
        RECT 466.950 180.450 469.050 181.050 ;
        RECT 433.950 179.400 469.050 180.450 ;
        RECT 433.950 178.950 436.050 179.400 ;
        RECT 466.950 178.950 469.050 179.400 ;
        RECT 496.950 180.450 499.050 181.050 ;
        RECT 517.950 180.450 520.050 180.900 ;
        RECT 526.950 180.450 529.050 181.050 ;
        RECT 496.950 179.400 516.450 180.450 ;
        RECT 496.950 178.950 499.050 179.400 ;
        RECT 16.950 177.450 19.050 178.050 ;
        RECT 25.950 177.450 28.050 178.050 ;
        RECT 16.950 176.400 28.050 177.450 ;
        RECT 16.950 175.950 19.050 176.400 ;
        RECT 25.950 175.950 28.050 176.400 ;
        RECT 64.950 177.450 67.050 178.050 ;
        RECT 112.950 177.450 115.050 178.050 ;
        RECT 64.950 176.400 115.050 177.450 ;
        RECT 64.950 175.950 67.050 176.400 ;
        RECT 112.950 175.950 115.050 176.400 ;
        RECT 169.950 177.450 172.050 178.050 ;
        RECT 205.950 177.450 208.050 178.050 ;
        RECT 169.950 176.400 208.050 177.450 ;
        RECT 169.950 175.950 172.050 176.400 ;
        RECT 205.950 175.950 208.050 176.400 ;
        RECT 235.950 177.450 238.050 177.900 ;
        RECT 277.950 177.450 280.050 178.050 ;
        RECT 235.950 176.400 280.050 177.450 ;
        RECT 235.950 175.800 238.050 176.400 ;
        RECT 277.950 175.950 280.050 176.400 ;
        RECT 343.950 177.450 346.050 178.050 ;
        RECT 352.950 177.450 355.050 178.050 ;
        RECT 343.950 176.400 355.050 177.450 ;
        RECT 343.950 175.950 346.050 176.400 ;
        RECT 352.950 175.950 355.050 176.400 ;
        RECT 481.950 177.450 484.050 178.050 ;
        RECT 499.950 177.450 502.050 178.050 ;
        RECT 481.950 176.400 502.050 177.450 ;
        RECT 515.400 177.450 516.450 179.400 ;
        RECT 517.950 179.400 529.050 180.450 ;
        RECT 554.400 180.450 555.450 182.400 ;
        RECT 556.950 182.400 634.050 183.450 ;
        RECT 556.950 181.950 559.050 182.400 ;
        RECT 631.950 181.950 634.050 182.400 ;
        RECT 691.950 183.450 694.050 184.050 ;
        RECT 739.950 183.450 742.050 184.050 ;
        RECT 691.950 182.400 742.050 183.450 ;
        RECT 691.950 181.950 694.050 182.400 ;
        RECT 739.950 181.950 742.050 182.400 ;
        RECT 748.950 183.450 751.050 184.050 ;
        RECT 784.950 183.450 787.050 184.050 ;
        RECT 748.950 182.400 787.050 183.450 ;
        RECT 748.950 181.950 751.050 182.400 ;
        RECT 784.950 181.950 787.050 182.400 ;
        RECT 799.950 183.450 802.050 184.050 ;
        RECT 826.950 183.450 829.050 184.050 ;
        RECT 799.950 182.400 829.050 183.450 ;
        RECT 799.950 181.950 802.050 182.400 ;
        RECT 826.950 181.950 829.050 182.400 ;
        RECT 562.950 180.450 565.050 181.050 ;
        RECT 554.400 179.400 565.050 180.450 ;
        RECT 517.950 178.800 520.050 179.400 ;
        RECT 526.950 178.950 529.050 179.400 ;
        RECT 562.950 178.950 565.050 179.400 ;
        RECT 742.950 180.450 745.050 181.050 ;
        RECT 796.950 180.450 799.050 181.050 ;
        RECT 742.950 179.400 799.050 180.450 ;
        RECT 742.950 178.950 745.050 179.400 ;
        RECT 796.950 178.950 799.050 179.400 ;
        RECT 838.950 180.450 841.050 181.050 ;
        RECT 853.950 180.450 856.050 181.050 ;
        RECT 838.950 179.400 856.050 180.450 ;
        RECT 838.950 178.950 841.050 179.400 ;
        RECT 853.950 178.950 856.050 179.400 ;
        RECT 520.950 177.450 523.050 178.050 ;
        RECT 515.400 176.400 523.050 177.450 ;
        RECT 481.950 175.950 484.050 176.400 ;
        RECT 499.950 175.950 502.050 176.400 ;
        RECT 520.950 175.950 523.050 176.400 ;
        RECT 700.950 177.450 703.050 178.050 ;
        RECT 727.950 177.450 730.050 178.050 ;
        RECT 700.950 176.400 730.050 177.450 ;
        RECT 700.950 175.950 703.050 176.400 ;
        RECT 727.950 175.950 730.050 176.400 ;
        RECT 769.950 177.450 772.050 178.050 ;
        RECT 784.950 177.450 787.050 178.050 ;
        RECT 769.950 176.400 787.050 177.450 ;
        RECT 769.950 175.950 772.050 176.400 ;
        RECT 784.950 175.950 787.050 176.400 ;
        RECT 823.950 177.450 826.050 178.050 ;
        RECT 835.950 177.450 838.050 178.050 ;
        RECT 823.950 176.400 838.050 177.450 ;
        RECT 823.950 175.950 826.050 176.400 ;
        RECT 835.950 175.950 838.050 176.400 ;
        RECT 13.950 174.450 16.050 175.050 ;
        RECT 25.950 174.450 28.050 175.050 ;
        RECT 43.950 174.450 46.050 175.050 ;
        RECT 13.950 173.400 46.050 174.450 ;
        RECT 13.950 172.950 16.050 173.400 ;
        RECT 25.950 172.950 28.050 173.400 ;
        RECT 43.950 172.950 46.050 173.400 ;
        RECT 85.950 174.450 88.050 175.050 ;
        RECT 100.950 174.450 103.050 175.050 ;
        RECT 106.950 174.450 109.050 175.050 ;
        RECT 85.950 173.400 109.050 174.450 ;
        RECT 85.950 172.950 88.050 173.400 ;
        RECT 100.950 172.950 103.050 173.400 ;
        RECT 106.950 172.950 109.050 173.400 ;
        RECT 118.950 174.450 121.050 175.050 ;
        RECT 139.950 174.450 142.050 175.050 ;
        RECT 118.950 173.400 142.050 174.450 ;
        RECT 118.950 172.950 121.050 173.400 ;
        RECT 139.950 172.950 142.050 173.400 ;
        RECT 148.950 174.450 151.050 175.050 ;
        RECT 178.950 174.450 181.050 175.050 ;
        RECT 202.950 174.450 205.050 175.050 ;
        RECT 148.950 173.400 205.050 174.450 ;
        RECT 148.950 172.950 151.050 173.400 ;
        RECT 178.950 172.950 181.050 173.400 ;
        RECT 202.950 172.950 205.050 173.400 ;
        RECT 214.950 174.450 217.050 175.050 ;
        RECT 250.950 174.450 256.050 175.050 ;
        RECT 214.950 173.400 256.050 174.450 ;
        RECT 214.950 172.950 217.050 173.400 ;
        RECT 250.950 172.950 256.050 173.400 ;
        RECT 271.950 172.950 277.050 175.050 ;
        RECT 376.950 174.450 379.050 175.050 ;
        RECT 418.950 174.450 421.050 175.050 ;
        RECT 454.950 174.450 457.050 175.050 ;
        RECT 490.950 174.450 493.050 175.050 ;
        RECT 526.950 174.450 529.050 175.050 ;
        RECT 376.950 174.000 438.450 174.450 ;
        RECT 376.950 173.400 439.050 174.000 ;
        RECT 376.950 172.950 379.050 173.400 ;
        RECT 418.950 172.950 421.050 173.400 ;
        RECT 13.950 166.950 16.050 172.050 ;
        RECT 19.950 166.950 22.050 172.050 ;
        RECT 73.950 171.450 76.050 172.050 ;
        RECT 91.950 171.450 94.050 172.050 ;
        RECT 151.950 171.450 154.050 172.050 ;
        RECT 73.950 170.400 94.050 171.450 ;
        RECT 24.000 168.450 28.050 169.050 ;
        RECT 23.400 166.950 28.050 168.450 ;
        RECT 40.950 168.450 43.050 169.050 ;
        RECT 52.950 168.450 55.050 169.050 ;
        RECT 40.950 167.400 55.050 168.450 ;
        RECT 4.950 165.450 7.050 166.050 ;
        RECT 10.950 165.450 13.050 166.050 ;
        RECT 4.950 164.400 13.050 165.450 ;
        RECT 4.950 163.950 7.050 164.400 ;
        RECT 10.950 163.950 13.050 164.400 ;
        RECT 16.950 165.450 19.050 166.050 ;
        RECT 23.400 165.450 24.450 166.950 ;
        RECT 40.950 166.050 43.050 167.400 ;
        RECT 52.950 166.950 55.050 167.400 ;
        RECT 61.950 166.950 67.050 169.050 ;
        RECT 73.950 166.950 76.050 170.400 ;
        RECT 91.950 169.950 94.050 170.400 ;
        RECT 137.400 170.400 154.050 171.450 ;
        RECT 80.400 167.400 102.450 168.450 ;
        RECT 80.400 166.050 81.450 167.400 ;
        RECT 101.400 166.050 102.450 167.400 ;
        RECT 109.950 166.950 115.050 169.050 ;
        RECT 118.950 168.450 121.050 169.050 ;
        RECT 137.400 168.450 138.450 170.400 ;
        RECT 151.950 169.950 154.050 170.400 ;
        RECT 202.950 171.450 205.050 172.050 ;
        RECT 217.950 171.450 220.050 172.050 ;
        RECT 202.950 170.400 220.050 171.450 ;
        RECT 118.950 167.400 138.450 168.450 ;
        RECT 118.950 166.950 121.050 167.400 ;
        RECT 16.950 164.400 24.450 165.450 ;
        RECT 25.950 165.450 28.050 166.050 ;
        RECT 34.950 165.450 37.050 166.050 ;
        RECT 25.950 164.400 37.050 165.450 ;
        RECT 16.950 163.950 19.050 164.400 ;
        RECT 25.950 163.950 28.050 164.400 ;
        RECT 34.950 163.950 37.050 164.400 ;
        RECT 40.800 165.000 43.050 166.050 ;
        RECT 44.100 165.450 46.200 166.050 ;
        RECT 49.950 165.450 52.050 166.050 ;
        RECT 40.800 163.950 42.900 165.000 ;
        RECT 44.100 164.400 52.050 165.450 ;
        RECT 44.100 163.950 46.200 164.400 ;
        RECT 49.950 163.950 52.050 164.400 ;
        RECT 31.950 160.950 36.900 163.050 ;
        RECT 38.100 162.450 40.200 163.050 ;
        RECT 46.950 162.450 49.050 163.050 ;
        RECT 55.950 162.450 58.050 166.050 ;
        RECT 38.100 162.000 58.050 162.450 ;
        RECT 70.950 162.450 73.050 166.050 ;
        RECT 76.950 164.400 81.450 166.050 ;
        RECT 76.950 163.950 81.000 164.400 ;
        RECT 88.950 163.950 94.050 166.050 ;
        RECT 97.950 163.950 103.050 166.050 ;
        RECT 106.950 165.450 109.050 166.050 ;
        RECT 115.950 165.450 118.050 166.050 ;
        RECT 106.950 164.400 118.050 165.450 ;
        RECT 106.950 163.950 109.050 164.400 ;
        RECT 115.950 163.950 118.050 164.400 ;
        RECT 121.950 165.450 124.050 166.050 ;
        RECT 127.950 165.450 130.050 166.050 ;
        RECT 133.950 165.450 136.050 166.050 ;
        RECT 121.950 164.400 136.050 165.450 ;
        RECT 121.950 163.950 124.050 164.400 ;
        RECT 127.950 163.950 130.050 164.400 ;
        RECT 133.950 163.950 136.050 164.400 ;
        RECT 139.950 163.950 142.050 169.050 ;
        RECT 154.950 166.950 159.900 169.050 ;
        RECT 161.100 166.950 165.900 169.050 ;
        RECT 167.100 166.950 172.050 169.050 ;
        RECT 202.950 166.950 205.050 170.400 ;
        RECT 217.950 169.950 220.050 170.400 ;
        RECT 253.950 171.450 256.050 172.050 ;
        RECT 268.950 171.450 271.050 172.050 ;
        RECT 277.950 171.450 283.050 172.050 ;
        RECT 253.950 170.400 283.050 171.450 ;
        RECT 253.950 169.950 256.050 170.400 ;
        RECT 268.950 169.950 271.050 170.400 ;
        RECT 277.950 169.950 283.050 170.400 ;
        RECT 343.950 171.450 346.050 172.050 ;
        RECT 361.950 171.450 364.050 172.050 ;
        RECT 343.950 170.400 364.050 171.450 ;
        RECT 343.950 169.950 346.050 170.400 ;
        RECT 361.950 169.950 364.050 170.400 ;
        RECT 421.950 169.950 427.050 172.050 ;
        RECT 436.950 171.450 439.050 173.400 ;
        RECT 454.950 173.400 529.050 174.450 ;
        RECT 454.950 172.950 457.050 173.400 ;
        RECT 490.950 172.950 493.050 173.400 ;
        RECT 526.950 172.950 529.050 173.400 ;
        RECT 535.950 174.450 538.050 175.050 ;
        RECT 541.950 174.450 544.050 175.050 ;
        RECT 535.950 173.400 544.050 174.450 ;
        RECT 553.950 173.400 556.050 175.500 ;
        RECT 574.950 173.400 577.050 175.500 ;
        RECT 622.950 174.450 625.050 175.050 ;
        RECT 643.950 174.450 646.050 175.050 ;
        RECT 622.950 173.400 646.050 174.450 ;
        RECT 535.950 172.950 538.050 173.400 ;
        RECT 541.950 172.950 544.050 173.400 ;
        RECT 451.950 171.450 454.050 172.050 ;
        RECT 463.950 171.450 466.050 172.050 ;
        RECT 487.950 171.450 490.050 172.050 ;
        RECT 496.800 171.450 498.900 172.050 ;
        RECT 436.950 170.400 454.050 171.450 ;
        RECT 458.400 171.000 477.450 171.450 ;
        RECT 436.950 169.950 439.050 170.400 ;
        RECT 451.950 169.950 454.050 170.400 ;
        RECT 457.950 170.400 478.050 171.000 ;
        RECT 233.400 168.000 246.450 168.450 ;
        RECT 233.400 167.400 247.050 168.000 ;
        RECT 82.950 162.450 85.050 163.050 ;
        RECT 94.950 162.450 97.050 163.050 ;
        RECT 70.950 162.000 97.050 162.450 ;
        RECT 38.100 161.400 57.450 162.000 ;
        RECT 71.400 161.400 97.050 162.000 ;
        RECT 38.100 160.950 40.200 161.400 ;
        RECT 46.950 160.950 49.050 161.400 ;
        RECT 82.950 160.950 85.050 161.400 ;
        RECT 94.950 160.950 97.050 161.400 ;
        RECT 103.950 162.450 106.050 163.050 ;
        RECT 118.950 162.450 121.050 163.050 ;
        RECT 103.950 161.400 121.050 162.450 ;
        RECT 103.950 160.950 106.050 161.400 ;
        RECT 118.950 160.950 121.050 161.400 ;
        RECT 133.950 160.950 139.050 163.050 ;
        RECT 145.950 162.450 148.050 163.050 ;
        RECT 160.950 162.450 163.050 166.050 ;
        RECT 145.950 162.000 163.050 162.450 ;
        RECT 166.950 162.450 169.050 166.050 ;
        RECT 175.950 163.950 180.900 166.050 ;
        RECT 182.100 163.950 187.050 166.050 ;
        RECT 196.950 163.950 202.050 166.050 ;
        RECT 172.950 162.450 175.050 163.050 ;
        RECT 166.950 162.000 175.050 162.450 ;
        RECT 145.950 161.400 162.450 162.000 ;
        RECT 167.400 161.400 175.050 162.000 ;
        RECT 145.950 160.950 148.050 161.400 ;
        RECT 172.950 160.950 175.050 161.400 ;
        RECT 100.950 159.450 103.050 160.050 ;
        RECT 145.950 159.450 148.050 160.050 ;
        RECT 100.950 158.400 148.050 159.450 ;
        RECT 100.950 157.950 103.050 158.400 ;
        RECT 145.950 157.950 148.050 158.400 ;
        RECT 151.950 159.450 154.050 160.050 ;
        RECT 181.950 159.450 184.050 163.050 ;
        RECT 190.950 160.950 196.050 163.050 ;
        RECT 205.950 160.950 208.050 166.050 ;
        RECT 223.950 165.450 226.050 166.050 ;
        RECT 233.400 165.450 234.450 167.400 ;
        RECT 223.950 164.400 234.450 165.450 ;
        RECT 223.950 163.950 226.050 164.400 ;
        RECT 238.950 163.050 241.050 166.050 ;
        RECT 244.950 163.950 247.050 167.400 ;
        RECT 256.950 166.950 262.050 169.050 ;
        RECT 265.950 168.450 268.050 169.050 ;
        RECT 289.950 168.450 292.050 169.050 ;
        RECT 265.950 167.400 292.050 168.450 ;
        RECT 265.950 166.950 268.050 167.400 ;
        RECT 289.950 166.950 292.050 167.400 ;
        RECT 295.950 168.450 298.050 169.050 ;
        RECT 319.950 168.450 322.050 169.050 ;
        RECT 295.950 167.400 322.050 168.450 ;
        RECT 217.950 160.950 223.050 163.050 ;
        RECT 196.950 159.450 199.050 160.050 ;
        RECT 226.950 159.450 229.050 163.050 ;
        RECT 238.800 162.000 241.050 163.050 ;
        RECT 242.100 162.000 244.200 163.050 ;
        RECT 238.800 160.950 240.900 162.000 ;
        RECT 241.950 160.950 244.200 162.000 ;
        RECT 151.950 159.000 229.050 159.450 ;
        RECT 232.950 159.450 235.050 160.050 ;
        RECT 241.950 159.450 244.050 160.950 ;
        RECT 232.950 159.000 244.050 159.450 ;
        RECT 247.950 159.450 250.050 163.050 ;
        RECT 253.950 162.450 256.050 163.050 ;
        RECT 262.950 162.450 265.050 166.050 ;
        RECT 253.950 162.000 265.050 162.450 ;
        RECT 253.950 161.400 264.450 162.000 ;
        RECT 253.950 160.950 256.050 161.400 ;
        RECT 268.950 160.950 271.050 166.050 ;
        RECT 286.950 165.450 289.050 166.050 ;
        RECT 286.950 164.400 294.450 165.450 ;
        RECT 286.950 163.950 289.050 164.400 ;
        RECT 293.400 162.450 294.450 164.400 ;
        RECT 295.950 163.950 298.050 167.400 ;
        RECT 319.950 166.950 322.050 167.400 ;
        RECT 328.950 168.450 333.000 169.050 ;
        RECT 328.950 166.950 333.450 168.450 ;
        RECT 334.950 166.950 340.050 169.050 ;
        RECT 343.950 168.450 346.050 169.050 ;
        RECT 349.950 168.450 352.050 169.050 ;
        RECT 357.000 168.450 361.050 169.050 ;
        RECT 343.950 167.400 352.050 168.450 ;
        RECT 343.950 166.950 346.050 167.400 ;
        RECT 349.950 166.950 352.050 167.400 ;
        RECT 356.400 166.950 361.050 168.450 ;
        RECT 364.950 168.450 367.050 169.050 ;
        RECT 370.950 168.450 373.050 169.050 ;
        RECT 364.950 167.400 373.050 168.450 ;
        RECT 364.950 166.950 367.050 167.400 ;
        RECT 370.950 166.950 373.050 167.400 ;
        RECT 406.950 168.450 409.050 169.050 ;
        RECT 418.950 168.450 421.050 169.050 ;
        RECT 406.950 167.400 421.050 168.450 ;
        RECT 406.950 166.950 409.050 167.400 ;
        RECT 418.950 166.950 421.050 167.400 ;
        RECT 424.950 166.950 430.050 169.050 ;
        RECT 457.950 166.950 460.050 170.400 ;
        RECT 463.950 169.950 466.050 170.400 ;
        RECT 463.950 166.950 469.050 169.050 ;
        RECT 475.950 166.950 478.050 170.400 ;
        RECT 487.950 170.400 498.900 171.450 ;
        RECT 500.100 171.000 502.200 172.050 ;
        RECT 487.950 169.950 490.050 170.400 ;
        RECT 496.800 169.950 498.900 170.400 ;
        RECT 499.950 169.950 502.200 171.000 ;
        RECT 511.950 171.450 514.050 172.050 ;
        RECT 544.950 171.450 549.000 172.050 ;
        RECT 511.950 170.400 522.450 171.450 ;
        RECT 511.950 169.950 514.050 170.400 ;
        RECT 499.950 169.050 502.050 169.950 ;
        RECT 521.400 169.050 522.450 170.400 ;
        RECT 544.950 169.950 549.450 171.450 ;
        RECT 548.400 169.050 549.450 169.950 ;
        RECT 484.950 168.450 487.050 169.050 ;
        RECT 493.800 168.450 495.900 169.050 ;
        RECT 484.950 167.400 495.900 168.450 ;
        RECT 484.950 166.950 487.050 167.400 ;
        RECT 493.800 166.950 495.900 167.400 ;
        RECT 496.800 168.000 498.900 169.050 ;
        RECT 499.950 168.000 502.200 169.050 ;
        RECT 496.800 166.950 499.050 168.000 ;
        RECT 500.100 166.950 502.200 168.000 ;
        RECT 508.950 168.450 511.050 169.050 ;
        RECT 517.950 168.450 520.050 169.050 ;
        RECT 508.950 167.400 520.050 168.450 ;
        RECT 521.400 167.400 526.050 169.050 ;
        RECT 508.950 166.950 511.050 167.400 ;
        RECT 517.950 166.950 520.050 167.400 ;
        RECT 522.000 166.950 526.050 167.400 ;
        RECT 529.950 168.450 534.000 169.050 ;
        RECT 541.950 168.450 544.050 169.050 ;
        RECT 548.400 168.450 553.050 169.050 ;
        RECT 529.950 166.950 534.450 168.450 ;
        RECT 541.950 167.400 553.050 168.450 ;
        RECT 541.950 166.950 544.050 167.400 ;
        RECT 549.000 166.950 553.050 167.400 ;
        RECT 301.950 165.450 307.050 166.050 ;
        RECT 316.950 165.450 319.050 166.050 ;
        RECT 301.950 164.400 319.050 165.450 ;
        RECT 301.950 163.950 307.050 164.400 ;
        RECT 316.950 163.950 319.050 164.400 ;
        RECT 298.950 162.450 301.050 163.050 ;
        RECT 322.950 162.450 325.050 166.050 ;
        RECT 332.400 165.450 333.450 166.950 ;
        RECT 340.950 165.450 345.900 166.050 ;
        RECT 332.400 164.400 345.900 165.450 ;
        RECT 347.100 165.450 349.200 166.050 ;
        RECT 356.400 165.450 357.450 166.950 ;
        RECT 347.100 165.000 357.450 165.450 ;
        RECT 340.950 163.950 345.900 164.400 ;
        RECT 346.950 164.400 357.450 165.000 ;
        RECT 346.950 163.950 349.200 164.400 ;
        RECT 358.950 163.950 364.050 166.050 ;
        RECT 293.400 162.000 325.050 162.450 ;
        RECT 325.950 162.450 328.050 163.050 ;
        RECT 334.950 162.450 337.050 163.050 ;
        RECT 346.950 162.450 349.050 163.950 ;
        RECT 325.950 162.000 349.050 162.450 ;
        RECT 367.950 162.450 370.050 166.050 ;
        RECT 373.950 165.450 376.050 166.050 ;
        RECT 379.800 165.450 381.900 166.050 ;
        RECT 373.950 164.400 381.900 165.450 ;
        RECT 373.950 163.950 376.050 164.400 ;
        RECT 379.800 163.950 381.900 164.400 ;
        RECT 383.100 163.950 388.050 166.050 ;
        RECT 391.950 165.450 394.050 166.050 ;
        RECT 403.950 165.450 406.050 166.050 ;
        RECT 412.950 165.450 415.050 166.050 ;
        RECT 391.950 164.400 406.050 165.450 ;
        RECT 407.400 165.000 415.050 165.450 ;
        RECT 391.950 163.950 394.050 164.400 ;
        RECT 403.950 163.950 406.050 164.400 ;
        RECT 406.950 164.400 415.050 165.000 ;
        RECT 382.950 162.450 385.050 163.050 ;
        RECT 367.950 162.000 385.050 162.450 ;
        RECT 293.400 161.400 324.450 162.000 ;
        RECT 325.950 161.400 348.600 162.000 ;
        RECT 368.400 161.400 385.050 162.000 ;
        RECT 298.950 160.950 301.050 161.400 ;
        RECT 325.950 160.950 328.050 161.400 ;
        RECT 334.950 160.950 337.050 161.400 ;
        RECT 304.950 159.450 307.050 160.050 ;
        RECT 247.950 159.000 307.050 159.450 ;
        RECT 151.950 158.400 228.450 159.000 ;
        RECT 232.950 158.400 243.600 159.000 ;
        RECT 248.400 158.400 307.050 159.000 ;
        RECT 151.950 157.950 154.050 158.400 ;
        RECT 196.950 157.950 199.050 158.400 ;
        RECT 232.950 157.950 235.050 158.400 ;
        RECT 304.950 157.950 307.050 158.400 ;
        RECT 310.950 159.450 313.050 160.050 ;
        RECT 382.950 159.450 385.050 161.400 ;
        RECT 391.950 162.450 394.050 163.050 ;
        RECT 400.950 162.450 403.050 163.050 ;
        RECT 391.950 161.400 403.050 162.450 ;
        RECT 391.950 160.950 394.050 161.400 ;
        RECT 400.950 160.950 403.050 161.400 ;
        RECT 406.950 160.950 409.050 164.400 ;
        RECT 412.950 163.950 415.050 164.400 ;
        RECT 430.950 165.450 433.050 166.050 ;
        RECT 436.950 165.450 439.050 166.050 ;
        RECT 430.950 164.400 439.050 165.450 ;
        RECT 430.950 163.950 433.050 164.400 ;
        RECT 436.950 163.950 439.050 164.400 ;
        RECT 451.950 163.950 457.050 166.050 ;
        RECT 460.950 160.950 463.050 166.050 ;
        RECT 472.950 160.950 475.050 166.050 ;
        RECT 478.950 160.950 481.050 166.050 ;
        RECT 496.950 163.950 499.050 166.950 ;
        RECT 514.950 165.450 517.050 166.050 ;
        RECT 520.800 165.450 522.900 166.050 ;
        RECT 514.950 164.400 522.900 165.450 ;
        RECT 514.950 163.950 517.050 164.400 ;
        RECT 520.800 163.950 522.900 164.400 ;
        RECT 524.100 163.950 529.050 166.050 ;
        RECT 533.400 165.450 534.450 166.950 ;
        RECT 538.950 165.450 541.050 166.050 ;
        RECT 533.400 164.400 541.050 165.450 ;
        RECT 538.950 163.950 541.050 164.400 ;
        RECT 554.850 161.400 556.050 173.400 ;
        RECT 559.950 166.950 565.050 169.050 ;
        RECT 562.950 165.450 565.050 165.900 ;
        RECT 568.950 165.450 571.050 169.050 ;
        RECT 562.950 165.000 571.050 165.450 ;
        RECT 562.950 164.400 570.450 165.000 ;
        RECT 562.950 163.800 565.050 164.400 ;
        RECT 310.950 159.000 385.050 159.450 ;
        RECT 457.950 159.450 460.050 160.050 ;
        RECT 478.950 159.450 481.050 160.050 ;
        RECT 310.950 158.400 384.450 159.000 ;
        RECT 457.950 158.400 481.050 159.450 ;
        RECT 310.950 157.950 313.050 158.400 ;
        RECT 457.950 157.950 460.050 158.400 ;
        RECT 478.950 157.950 481.050 158.400 ;
        RECT 508.950 159.450 511.050 160.050 ;
        RECT 535.950 159.450 538.050 160.050 ;
        RECT 508.950 158.400 538.050 159.450 ;
        RECT 553.950 159.300 556.050 161.400 ;
        RECT 508.950 157.950 511.050 158.400 ;
        RECT 535.950 157.950 538.050 158.400 ;
        RECT 166.950 156.450 169.050 157.050 ;
        RECT 238.950 156.450 241.050 157.050 ;
        RECT 166.950 155.400 241.050 156.450 ;
        RECT 166.950 154.950 169.050 155.400 ;
        RECT 238.950 154.950 241.050 155.400 ;
        RECT 403.950 156.450 406.050 157.050 ;
        RECT 409.950 156.450 412.050 157.050 ;
        RECT 403.950 155.400 412.050 156.450 ;
        RECT 403.950 154.950 406.050 155.400 ;
        RECT 409.950 154.950 412.050 155.400 ;
        RECT 427.950 156.450 430.050 157.050 ;
        RECT 460.950 156.450 463.050 157.050 ;
        RECT 427.950 155.400 463.050 156.450 ;
        RECT 554.850 155.700 556.050 159.300 ;
        RECT 575.100 156.600 576.300 173.400 ;
        RECT 622.950 172.950 625.050 173.400 ;
        RECT 643.950 172.950 646.050 173.400 ;
        RECT 679.950 174.450 682.050 175.050 ;
        RECT 748.950 174.450 751.050 175.050 ;
        RECT 679.950 173.400 751.050 174.450 ;
        RECT 679.950 172.950 682.050 173.400 ;
        RECT 748.950 172.950 751.050 173.400 ;
        RECT 595.950 169.950 601.050 172.050 ;
        RECT 652.950 171.450 655.050 172.050 ;
        RECT 667.950 171.450 670.050 172.050 ;
        RECT 652.950 170.400 670.050 171.450 ;
        RECT 652.950 169.950 655.050 170.400 ;
        RECT 667.950 169.950 670.050 170.400 ;
        RECT 577.950 168.450 580.050 169.050 ;
        RECT 592.800 168.450 594.900 169.050 ;
        RECT 577.950 167.400 594.900 168.450 ;
        RECT 577.950 166.950 580.050 167.400 ;
        RECT 592.800 166.950 594.900 167.400 ;
        RECT 596.100 166.950 601.050 169.050 ;
        RECT 610.950 166.950 616.050 169.050 ;
        RECT 681.000 168.450 685.050 169.050 ;
        RECT 680.400 166.950 685.050 168.450 ;
        RECT 688.950 166.950 691.050 172.050 ;
        RECT 697.950 171.450 700.050 172.050 ;
        RECT 709.950 171.450 712.050 172.050 ;
        RECT 697.950 170.400 712.050 171.450 ;
        RECT 697.950 169.950 700.050 170.400 ;
        RECT 709.950 169.950 712.050 170.400 ;
        RECT 718.950 171.450 721.050 172.050 ;
        RECT 730.950 171.450 733.050 172.050 ;
        RECT 718.950 170.400 733.050 171.450 ;
        RECT 718.950 169.950 721.050 170.400 ;
        RECT 730.950 169.950 733.050 170.400 ;
        RECT 751.950 169.950 757.050 172.050 ;
        RECT 763.950 169.950 766.050 175.050 ;
        RECT 772.950 174.450 775.050 175.050 ;
        RECT 787.950 174.450 790.050 175.050 ;
        RECT 805.950 174.450 808.050 175.050 ;
        RECT 832.950 174.450 835.050 175.050 ;
        RECT 772.950 173.400 790.050 174.450 ;
        RECT 772.950 172.950 775.050 173.400 ;
        RECT 787.950 172.950 790.050 173.400 ;
        RECT 791.400 173.400 835.050 174.450 ;
        RECT 736.950 168.450 739.050 169.050 ;
        RECT 692.250 168.000 739.050 168.450 ;
        RECT 691.950 167.400 739.050 168.000 ;
        RECT 616.950 163.950 622.050 166.050 ;
        RECT 631.950 163.950 637.050 166.050 ;
        RECT 640.950 163.050 643.050 166.050 ;
        RECT 649.950 163.950 655.050 166.050 ;
        RECT 673.950 165.450 676.050 166.050 ;
        RECT 680.400 165.450 681.450 166.950 ;
        RECT 691.950 166.050 694.050 167.400 ;
        RECT 728.400 166.050 729.450 167.400 ;
        RECT 736.950 166.950 739.050 167.400 ;
        RECT 742.950 166.950 748.050 169.050 ;
        RECT 766.950 166.950 772.050 169.050 ;
        RECT 775.950 166.950 778.050 172.050 ;
        RECT 791.400 169.050 792.450 173.400 ;
        RECT 805.950 172.950 808.050 173.400 ;
        RECT 790.950 166.950 793.050 169.050 ;
        RECT 796.950 166.950 799.050 172.050 ;
        RECT 811.950 169.950 817.050 172.050 ;
        RECT 827.400 169.050 828.450 173.400 ;
        RECT 832.950 172.950 835.050 173.400 ;
        RECT 847.950 172.950 850.050 178.050 ;
        RECT 829.950 171.450 832.050 172.050 ;
        RECT 835.950 171.450 838.050 172.050 ;
        RECT 829.950 170.400 838.050 171.450 ;
        RECT 829.950 169.950 832.050 170.400 ;
        RECT 835.950 169.950 838.050 170.400 ;
        RECT 805.950 168.450 808.050 169.050 ;
        RECT 811.950 168.450 814.050 169.050 ;
        RECT 805.950 167.400 814.050 168.450 ;
        RECT 805.950 166.950 808.050 167.400 ;
        RECT 811.950 166.950 814.050 167.400 ;
        RECT 817.950 166.950 823.050 169.050 ;
        RECT 827.400 167.400 832.050 169.050 ;
        RECT 828.000 166.950 832.050 167.400 ;
        RECT 835.950 168.450 838.050 169.050 ;
        RECT 841.950 168.450 847.050 169.050 ;
        RECT 835.950 167.400 847.050 168.450 ;
        RECT 835.950 166.950 838.050 167.400 ;
        RECT 841.950 166.950 847.050 167.400 ;
        RECT 673.950 164.400 681.450 165.450 ;
        RECT 673.950 163.950 676.050 164.400 ;
        RECT 682.950 163.950 688.050 166.050 ;
        RECT 691.800 165.000 694.050 166.050 ;
        RECT 695.100 165.450 697.200 166.050 ;
        RECT 703.950 165.450 706.050 166.050 ;
        RECT 691.800 163.950 693.900 165.000 ;
        RECT 695.100 164.400 706.050 165.450 ;
        RECT 695.100 163.950 697.200 164.400 ;
        RECT 703.950 163.950 706.050 164.400 ;
        RECT 724.950 164.400 729.450 166.050 ;
        RECT 724.950 163.950 729.000 164.400 ;
        RECT 730.950 163.950 736.050 166.050 ;
        RECT 739.950 165.450 742.050 166.050 ;
        RECT 754.950 165.450 757.050 166.050 ;
        RECT 739.950 164.400 757.050 165.450 ;
        RECT 739.950 163.950 742.050 164.400 ;
        RECT 754.950 163.950 757.050 164.400 ;
        RECT 769.950 163.950 775.050 166.050 ;
        RECT 778.950 163.950 784.050 166.050 ;
        RECT 787.950 165.450 790.050 166.050 ;
        RECT 793.950 165.450 796.050 166.050 ;
        RECT 787.950 164.400 796.050 165.450 ;
        RECT 787.950 163.950 790.050 164.400 ;
        RECT 793.950 163.950 796.050 164.400 ;
        RECT 595.950 162.450 598.050 163.050 ;
        RECT 610.950 162.450 613.050 163.050 ;
        RECT 595.950 161.400 613.050 162.450 ;
        RECT 595.950 160.950 598.050 161.400 ;
        RECT 610.950 160.950 613.050 161.400 ;
        RECT 625.950 160.950 631.050 163.050 ;
        RECT 634.950 160.950 639.900 163.050 ;
        RECT 640.950 162.000 643.200 163.050 ;
        RECT 641.100 160.950 643.200 162.000 ;
        RECT 646.950 160.950 652.050 163.050 ;
        RECT 655.950 162.450 658.050 163.050 ;
        RECT 688.950 162.450 691.050 163.050 ;
        RECT 655.950 161.400 691.050 162.450 ;
        RECT 655.950 160.950 658.050 161.400 ;
        RECT 688.950 160.950 691.050 161.400 ;
        RECT 703.950 162.450 706.050 163.050 ;
        RECT 724.950 162.450 727.050 163.050 ;
        RECT 703.950 161.400 727.050 162.450 ;
        RECT 703.950 160.950 706.050 161.400 ;
        RECT 724.950 160.950 727.050 161.400 ;
        RECT 766.950 162.450 769.050 163.050 ;
        RECT 790.950 162.450 793.050 163.050 ;
        RECT 799.950 162.450 802.050 166.050 ;
        RECT 826.950 165.450 829.050 166.050 ;
        RECT 832.950 165.450 835.050 166.050 ;
        RECT 826.950 164.400 835.050 165.450 ;
        RECT 826.950 163.950 829.050 164.400 ;
        RECT 832.950 163.950 835.050 164.400 ;
        RECT 766.950 162.000 802.050 162.450 ;
        RECT 766.950 161.400 801.450 162.000 ;
        RECT 766.950 160.950 769.050 161.400 ;
        RECT 790.950 160.950 793.050 161.400 ;
        RECT 838.950 160.950 841.050 166.050 ;
        RECT 640.950 159.450 643.050 160.050 ;
        RECT 655.950 159.450 658.050 160.050 ;
        RECT 640.950 158.400 658.050 159.450 ;
        RECT 640.950 157.950 643.050 158.400 ;
        RECT 655.950 157.950 658.050 158.400 ;
        RECT 706.950 159.450 709.050 160.050 ;
        RECT 763.950 159.450 766.050 160.050 ;
        RECT 706.950 158.400 766.050 159.450 ;
        RECT 706.950 157.950 709.050 158.400 ;
        RECT 763.950 157.950 766.050 158.400 ;
        RECT 778.950 159.450 781.050 160.050 ;
        RECT 796.950 159.450 799.050 160.050 ;
        RECT 778.950 158.400 799.050 159.450 ;
        RECT 778.950 157.950 781.050 158.400 ;
        RECT 796.950 157.950 799.050 158.400 ;
        RECT 814.950 159.450 817.050 160.050 ;
        RECT 844.950 159.450 847.050 160.050 ;
        RECT 814.950 158.400 847.050 159.450 ;
        RECT 814.950 157.950 817.050 158.400 ;
        RECT 844.950 157.950 847.050 158.400 ;
        RECT 427.950 154.950 430.050 155.400 ;
        RECT 460.950 154.950 463.050 155.400 ;
        RECT 40.950 153.450 43.050 154.050 ;
        RECT 181.950 153.450 184.050 154.050 ;
        RECT 205.950 153.450 208.050 154.050 ;
        RECT 40.950 152.400 208.050 153.450 ;
        RECT 40.950 151.950 43.050 152.400 ;
        RECT 181.950 151.950 184.050 152.400 ;
        RECT 205.950 151.950 208.050 152.400 ;
        RECT 274.950 148.950 277.050 154.050 ;
        RECT 331.950 153.450 334.050 154.050 ;
        RECT 499.950 153.450 502.050 154.050 ;
        RECT 553.950 153.600 556.050 155.700 ;
        RECT 574.950 154.500 577.050 156.600 ;
        RECT 622.950 154.950 628.050 157.050 ;
        RECT 634.950 156.450 637.050 157.050 ;
        RECT 646.950 156.450 649.050 157.050 ;
        RECT 634.950 155.400 649.050 156.450 ;
        RECT 634.950 154.950 637.050 155.400 ;
        RECT 646.950 154.950 649.050 155.400 ;
        RECT 670.950 156.450 673.050 157.050 ;
        RECT 730.950 156.450 733.050 157.050 ;
        RECT 670.950 155.400 733.050 156.450 ;
        RECT 670.950 154.950 673.050 155.400 ;
        RECT 730.950 154.950 733.050 155.400 ;
        RECT 748.950 156.450 751.050 157.050 ;
        RECT 754.950 156.450 757.050 157.050 ;
        RECT 748.950 155.400 757.050 156.450 ;
        RECT 748.950 154.950 751.050 155.400 ;
        RECT 754.950 154.950 757.050 155.400 ;
        RECT 817.950 156.450 820.050 157.050 ;
        RECT 823.950 156.450 826.050 157.050 ;
        RECT 817.950 155.400 826.050 156.450 ;
        RECT 817.950 154.950 820.050 155.400 ;
        RECT 823.950 154.950 826.050 155.400 ;
        RECT 331.950 152.400 502.050 153.450 ;
        RECT 331.950 151.950 334.050 152.400 ;
        RECT 499.950 151.950 502.050 152.400 ;
        RECT 751.950 153.450 754.050 154.050 ;
        RECT 760.950 153.450 763.050 154.050 ;
        RECT 751.950 152.400 763.050 153.450 ;
        RECT 751.950 151.950 754.050 152.400 ;
        RECT 760.950 151.950 763.050 152.400 ;
        RECT 805.950 153.450 808.050 154.050 ;
        RECT 832.950 153.450 835.050 154.050 ;
        RECT 805.950 152.400 835.050 153.450 ;
        RECT 805.950 151.950 808.050 152.400 ;
        RECT 832.950 151.950 835.050 152.400 ;
        RECT 364.950 150.450 367.050 151.050 ;
        RECT 388.950 150.450 391.050 151.050 ;
        RECT 364.950 149.400 391.050 150.450 ;
        RECT 364.950 148.950 367.050 149.400 ;
        RECT 388.950 148.950 391.050 149.400 ;
        RECT 409.950 150.450 412.050 151.050 ;
        RECT 487.950 150.450 490.050 151.050 ;
        RECT 409.950 149.400 490.050 150.450 ;
        RECT 409.950 148.950 412.050 149.400 ;
        RECT 487.950 148.950 490.050 149.400 ;
        RECT 511.950 150.450 514.050 151.050 ;
        RECT 541.950 150.450 544.050 151.050 ;
        RECT 547.800 150.450 549.900 151.050 ;
        RECT 511.950 149.400 540.450 150.450 ;
        RECT 511.950 148.950 514.050 149.400 ;
        RECT 539.400 147.450 540.450 149.400 ;
        RECT 541.950 149.400 549.900 150.450 ;
        RECT 541.950 148.950 544.050 149.400 ;
        RECT 547.800 148.950 549.900 149.400 ;
        RECT 673.950 150.450 676.050 151.050 ;
        RECT 766.950 150.450 769.050 151.050 ;
        RECT 673.950 149.400 769.050 150.450 ;
        RECT 673.950 148.950 676.050 149.400 ;
        RECT 766.950 148.950 769.050 149.400 ;
        RECT 784.950 150.450 787.050 151.050 ;
        RECT 838.950 150.450 841.050 151.200 ;
        RECT 784.950 149.400 841.050 150.450 ;
        RECT 784.950 148.950 787.050 149.400 ;
        RECT 838.950 149.100 841.050 149.400 ;
        RECT 562.950 147.450 565.050 148.050 ;
        RECT 539.400 146.400 565.050 147.450 ;
        RECT 562.950 145.950 565.050 146.400 ;
        RECT 610.950 147.450 613.050 148.050 ;
        RECT 622.950 147.450 625.050 148.050 ;
        RECT 610.950 146.400 625.050 147.450 ;
        RECT 610.950 145.950 613.050 146.400 ;
        RECT 622.950 145.950 625.050 146.400 ;
        RECT 646.950 147.450 649.050 148.050 ;
        RECT 655.950 147.450 658.050 148.050 ;
        RECT 646.950 146.400 658.050 147.450 ;
        RECT 646.950 145.950 649.050 146.400 ;
        RECT 655.950 145.950 658.050 146.400 ;
        RECT 748.950 147.450 751.050 148.050 ;
        RECT 763.950 147.450 766.050 148.050 ;
        RECT 748.950 146.400 766.050 147.450 ;
        RECT 748.950 145.950 751.050 146.400 ;
        RECT 763.950 145.950 766.050 146.400 ;
        RECT 823.950 147.450 826.050 148.050 ;
        RECT 829.950 147.450 832.050 148.050 ;
        RECT 823.950 146.400 832.050 147.450 ;
        RECT 823.950 145.950 826.050 146.400 ;
        RECT 829.950 145.950 832.050 146.400 ;
        RECT 838.950 147.450 841.050 147.900 ;
        RECT 847.950 147.450 850.050 151.050 ;
        RECT 838.950 147.000 850.050 147.450 ;
        RECT 838.950 146.400 849.450 147.000 ;
        RECT 838.950 145.800 841.050 146.400 ;
        RECT 397.950 144.450 400.050 145.050 ;
        RECT 475.950 144.450 478.050 145.050 ;
        RECT 397.950 143.400 478.050 144.450 ;
        RECT 397.950 142.950 400.050 143.400 ;
        RECT 475.950 142.950 478.050 143.400 ;
        RECT 568.950 144.450 571.050 145.050 ;
        RECT 604.950 144.450 607.050 145.050 ;
        RECT 649.950 144.450 652.050 145.050 ;
        RECT 568.950 143.400 652.050 144.450 ;
        RECT 568.950 142.950 571.050 143.400 ;
        RECT 604.950 142.950 607.050 143.400 ;
        RECT 649.950 142.950 652.050 143.400 ;
        RECT 661.950 144.450 664.050 145.050 ;
        RECT 718.950 144.450 721.050 145.050 ;
        RECT 661.950 143.400 721.050 144.450 ;
        RECT 661.950 142.950 664.050 143.400 ;
        RECT 718.950 142.950 721.050 143.400 ;
        RECT 724.950 144.450 727.050 145.050 ;
        RECT 769.950 144.450 772.050 145.050 ;
        RECT 724.950 143.400 772.050 144.450 ;
        RECT 724.950 142.950 727.050 143.400 ;
        RECT 769.950 142.950 772.050 143.400 ;
        RECT 37.950 141.450 40.050 142.050 ;
        RECT 55.950 141.450 58.050 142.050 ;
        RECT 37.950 140.400 58.050 141.450 ;
        RECT 37.950 139.950 40.050 140.400 ;
        RECT 55.950 139.950 58.050 140.400 ;
        RECT 103.950 141.450 106.050 142.050 ;
        RECT 145.950 141.450 148.050 142.050 ;
        RECT 103.950 140.400 148.050 141.450 ;
        RECT 103.950 139.950 106.050 140.400 ;
        RECT 145.950 139.950 148.050 140.400 ;
        RECT 151.950 141.450 154.050 142.050 ;
        RECT 172.950 141.450 175.050 142.050 ;
        RECT 232.950 141.450 235.050 142.050 ;
        RECT 151.950 140.400 235.050 141.450 ;
        RECT 151.950 139.950 154.050 140.400 ;
        RECT 172.950 139.950 175.050 140.400 ;
        RECT 232.950 139.950 235.050 140.400 ;
        RECT 454.950 141.450 457.050 142.050 ;
        RECT 484.950 141.450 487.050 142.050 ;
        RECT 454.950 140.400 487.050 141.450 ;
        RECT 454.950 139.950 457.050 140.400 ;
        RECT 484.950 139.950 487.050 140.400 ;
        RECT 532.950 141.450 535.050 142.050 ;
        RECT 574.950 141.450 577.050 142.050 ;
        RECT 532.950 140.400 577.050 141.450 ;
        RECT 532.950 139.950 535.050 140.400 ;
        RECT 574.950 139.950 577.050 140.400 ;
        RECT 616.950 141.450 619.050 142.050 ;
        RECT 655.950 141.450 658.050 142.050 ;
        RECT 616.950 140.400 658.050 141.450 ;
        RECT 616.950 139.950 619.050 140.400 ;
        RECT 655.950 139.950 658.050 140.400 ;
        RECT 700.950 141.450 703.050 142.050 ;
        RECT 757.950 141.450 760.050 142.050 ;
        RECT 700.950 140.400 760.050 141.450 ;
        RECT 700.950 139.950 703.050 140.400 ;
        RECT 757.950 139.950 760.050 140.400 ;
        RECT 793.950 141.450 796.050 142.050 ;
        RECT 808.950 141.450 811.050 142.050 ;
        RECT 793.950 140.400 811.050 141.450 ;
        RECT 793.950 139.950 796.050 140.400 ;
        RECT 808.950 139.950 811.050 140.400 ;
        RECT 817.950 139.950 823.050 142.050 ;
        RECT 832.950 141.450 835.050 142.050 ;
        RECT 844.950 141.450 847.050 142.050 ;
        RECT 832.950 140.400 847.050 141.450 ;
        RECT 832.950 139.950 835.050 140.400 ;
        RECT 844.950 139.950 847.050 140.400 ;
        RECT 49.950 138.450 52.050 139.050 ;
        RECT 88.950 138.450 91.050 139.050 ;
        RECT 103.950 138.450 106.050 139.050 ;
        RECT 49.950 137.400 106.050 138.450 ;
        RECT 49.950 136.950 52.050 137.400 ;
        RECT 88.950 136.950 91.050 137.400 ;
        RECT 103.950 136.950 106.050 137.400 ;
        RECT 196.950 138.450 199.050 139.050 ;
        RECT 274.950 138.450 277.050 139.050 ;
        RECT 196.950 137.400 277.050 138.450 ;
        RECT 196.950 136.950 199.050 137.400 ;
        RECT 274.950 136.950 277.050 137.400 ;
        RECT 298.950 138.450 301.050 139.050 ;
        RECT 346.950 138.450 349.050 139.050 ;
        RECT 298.950 137.400 349.050 138.450 ;
        RECT 298.950 136.950 301.050 137.400 ;
        RECT 346.950 136.950 349.050 137.400 ;
        RECT 529.950 138.450 532.050 139.050 ;
        RECT 559.950 138.450 562.050 139.050 ;
        RECT 529.950 137.400 562.050 138.450 ;
        RECT 529.950 136.950 532.050 137.400 ;
        RECT 559.950 136.950 562.050 137.400 ;
        RECT 613.950 138.450 616.050 139.050 ;
        RECT 625.950 138.450 628.050 139.050 ;
        RECT 613.950 137.400 628.050 138.450 ;
        RECT 613.950 136.950 616.050 137.400 ;
        RECT 625.950 136.950 628.050 137.400 ;
        RECT 676.950 138.450 679.050 139.050 ;
        RECT 721.950 138.450 724.050 139.050 ;
        RECT 676.950 137.400 724.050 138.450 ;
        RECT 676.950 136.950 679.050 137.400 ;
        RECT 721.950 136.950 724.050 137.400 ;
        RECT 727.950 138.450 730.050 139.050 ;
        RECT 745.950 138.450 748.050 139.050 ;
        RECT 727.950 137.400 748.050 138.450 ;
        RECT 727.950 136.950 730.050 137.400 ;
        RECT 745.950 136.950 748.050 137.400 ;
        RECT 757.950 138.450 760.050 139.050 ;
        RECT 775.950 138.450 778.050 139.050 ;
        RECT 757.950 137.400 778.050 138.450 ;
        RECT 757.950 136.950 760.050 137.400 ;
        RECT 775.950 136.950 778.050 137.400 ;
        RECT 784.950 138.450 787.050 139.050 ;
        RECT 853.950 138.450 856.050 139.050 ;
        RECT 784.950 137.400 856.050 138.450 ;
        RECT 784.950 136.950 787.050 137.400 ;
        RECT 853.950 136.950 856.050 137.400 ;
        RECT 13.950 135.450 16.050 136.050 ;
        RECT 37.950 135.450 40.050 136.050 ;
        RECT 106.950 135.450 109.050 136.050 ;
        RECT 121.950 135.450 124.050 136.050 ;
        RECT 13.950 134.400 124.050 135.450 ;
        RECT 13.950 133.950 16.050 134.400 ;
        RECT 37.950 133.950 40.050 134.400 ;
        RECT 106.950 133.950 109.050 134.400 ;
        RECT 121.950 133.950 124.050 134.400 ;
        RECT 271.950 135.450 274.050 136.050 ;
        RECT 307.950 135.450 310.050 136.050 ;
        RECT 271.950 134.400 310.050 135.450 ;
        RECT 271.950 133.950 274.050 134.400 ;
        RECT 307.950 133.950 310.050 134.400 ;
        RECT 427.950 135.450 430.050 136.050 ;
        RECT 466.950 135.450 469.050 136.050 ;
        RECT 472.950 135.450 475.050 136.050 ;
        RECT 427.950 134.400 475.050 135.450 ;
        RECT 427.950 133.950 430.050 134.400 ;
        RECT 466.950 133.950 469.050 134.400 ;
        RECT 472.950 133.950 475.050 134.400 ;
        RECT 586.950 135.450 589.050 136.050 ;
        RECT 646.950 135.450 649.050 136.050 ;
        RECT 664.950 135.450 667.050 136.050 ;
        RECT 586.950 134.400 636.450 135.450 ;
        RECT 586.950 133.950 589.050 134.400 ;
        RECT 22.950 132.450 25.050 133.050 ;
        RECT 34.950 132.450 37.050 133.050 ;
        RECT 103.950 132.450 106.050 133.050 ;
        RECT 178.950 132.450 181.050 133.050 ;
        RECT 235.950 132.450 238.050 133.050 ;
        RECT 253.950 132.450 256.050 133.050 ;
        RECT 22.950 131.400 37.050 132.450 ;
        RECT 22.950 130.950 25.050 131.400 ;
        RECT 34.950 130.950 37.050 131.400 ;
        RECT 92.400 131.400 108.600 132.450 ;
        RECT 13.950 126.450 16.050 127.050 ;
        RECT 22.950 126.450 25.050 127.050 ;
        RECT 13.950 125.400 25.050 126.450 ;
        RECT 13.950 124.950 16.050 125.400 ;
        RECT 22.950 124.950 25.050 125.400 ;
        RECT 28.950 124.950 31.050 130.050 ;
        RECT 46.950 127.950 52.050 130.050 ;
        RECT 55.950 127.950 61.050 130.050 ;
        RECT 67.950 127.050 70.050 130.050 ;
        RECT 76.950 129.450 79.050 130.050 ;
        RECT 92.400 129.450 93.450 131.400 ;
        RECT 103.950 130.950 106.050 131.400 ;
        RECT 76.950 128.400 93.450 129.450 ;
        RECT 76.950 127.950 79.050 128.400 ;
        RECT 91.800 127.050 93.900 127.200 ;
        RECT 107.550 127.050 108.600 131.400 ;
        RECT 178.950 131.400 256.050 132.450 ;
        RECT 178.950 130.950 181.050 131.400 ;
        RECT 235.950 130.950 238.050 131.400 ;
        RECT 253.950 130.950 256.050 131.400 ;
        RECT 280.950 132.450 283.050 133.050 ;
        RECT 301.950 132.450 304.050 133.050 ;
        RECT 340.950 132.450 343.050 133.050 ;
        RECT 361.950 132.450 364.050 133.050 ;
        RECT 280.950 131.400 343.050 132.450 ;
        RECT 280.950 130.950 283.050 131.400 ;
        RECT 301.950 130.950 304.050 131.400 ;
        RECT 340.950 130.950 343.050 131.400 ;
        RECT 344.400 131.400 364.050 132.450 ;
        RECT 109.950 127.950 115.050 130.050 ;
        RECT 118.950 129.450 121.050 130.050 ;
        RECT 127.950 129.450 130.050 130.050 ;
        RECT 184.950 129.450 187.050 130.050 ;
        RECT 118.950 128.400 130.050 129.450 ;
        RECT 134.400 129.000 187.050 129.450 ;
        RECT 118.950 127.950 121.050 128.400 ;
        RECT 127.950 127.950 130.050 128.400 ;
        RECT 133.950 128.400 187.050 129.000 ;
        RECT 34.950 126.450 37.050 127.050 ;
        RECT 43.950 126.450 46.050 127.050 ;
        RECT 34.950 125.400 46.050 126.450 ;
        RECT 34.950 124.950 37.050 125.400 ;
        RECT 43.950 124.950 46.050 125.400 ;
        RECT 13.950 118.950 19.050 121.050 ;
        RECT 25.950 118.950 28.050 124.050 ;
        RECT 49.950 123.450 52.050 127.050 ;
        RECT 61.950 124.950 66.900 127.050 ;
        RECT 67.950 126.000 70.200 127.050 ;
        RECT 71.100 126.000 73.200 127.050 ;
        RECT 68.100 124.950 70.200 126.000 ;
        RECT 70.950 124.950 73.200 126.000 ;
        RECT 88.950 125.100 93.900 127.050 ;
        RECT 95.100 126.450 97.200 127.050 ;
        RECT 103.800 126.450 105.900 127.050 ;
        RECT 95.100 125.400 105.900 126.450 ;
        RECT 88.950 124.950 93.000 125.100 ;
        RECT 95.100 124.950 97.200 125.400 ;
        RECT 103.800 124.950 105.900 125.400 ;
        RECT 107.100 124.950 109.200 127.050 ;
        RECT 70.950 123.450 73.050 124.950 ;
        RECT 85.950 123.450 88.050 124.050 ;
        RECT 49.950 123.000 88.050 123.450 ;
        RECT 50.400 122.400 88.050 123.000 ;
        RECT 85.950 121.950 88.050 122.400 ;
        RECT 91.950 121.950 96.900 124.050 ;
        RECT 98.100 123.000 100.200 124.050 ;
        RECT 112.950 123.450 115.050 127.050 ;
        RECT 121.950 126.450 124.050 127.050 ;
        RECT 127.950 126.450 130.050 127.050 ;
        RECT 133.950 126.450 136.050 128.400 ;
        RECT 184.950 127.950 187.050 128.400 ;
        RECT 196.950 129.450 199.050 130.050 ;
        RECT 202.950 129.450 205.050 130.050 ;
        RECT 196.950 128.400 205.050 129.450 ;
        RECT 121.950 125.400 130.050 126.450 ;
        RECT 121.950 124.950 124.050 125.400 ;
        RECT 127.950 124.950 130.050 125.400 ;
        RECT 131.400 125.400 136.050 126.450 ;
        RECT 131.400 123.450 132.450 125.400 ;
        RECT 133.950 124.950 136.050 125.400 ;
        RECT 139.950 126.450 142.050 127.050 ;
        RECT 151.950 126.450 154.050 127.050 ;
        RECT 139.950 125.400 154.050 126.450 ;
        RECT 139.950 124.950 142.050 125.400 ;
        RECT 151.950 124.950 154.050 125.400 ;
        RECT 157.950 124.050 160.050 127.050 ;
        RECT 187.800 126.450 189.900 127.050 ;
        RECT 173.550 126.000 189.900 126.450 ;
        RECT 191.100 126.000 193.200 127.050 ;
        RECT 172.950 125.400 189.900 126.000 ;
        RECT 172.950 124.050 175.050 125.400 ;
        RECT 187.800 124.950 189.900 125.400 ;
        RECT 190.950 124.950 193.200 126.000 ;
        RECT 196.950 124.950 199.050 128.400 ;
        RECT 202.950 127.950 205.050 128.400 ;
        RECT 244.950 129.450 247.050 130.050 ;
        RECT 265.950 129.450 268.050 130.050 ;
        RECT 286.950 129.450 289.050 130.050 ;
        RECT 298.950 129.450 301.050 130.050 ;
        RECT 325.950 129.450 328.050 130.050 ;
        RECT 344.400 129.450 345.450 131.400 ;
        RECT 361.950 130.950 364.050 131.400 ;
        RECT 244.950 128.400 301.050 129.450 ;
        RECT 314.400 129.000 345.450 129.450 ;
        RECT 244.950 127.950 247.050 128.400 ;
        RECT 265.950 127.950 268.050 128.400 ;
        RECT 286.950 127.950 289.050 128.400 ;
        RECT 298.950 127.950 301.050 128.400 ;
        RECT 313.950 128.400 345.450 129.000 ;
        RECT 370.950 129.450 373.050 130.050 ;
        RECT 385.950 129.450 388.050 130.050 ;
        RECT 370.950 128.400 388.050 129.450 ;
        RECT 214.950 124.950 219.900 127.050 ;
        RECT 221.100 124.950 226.050 127.050 ;
        RECT 289.950 124.950 295.050 127.050 ;
        RECT 304.950 124.950 310.050 127.050 ;
        RECT 313.950 124.950 316.050 128.400 ;
        RECT 325.950 127.950 328.050 128.400 ;
        RECT 370.950 127.950 373.050 128.400 ;
        RECT 385.950 127.950 388.050 128.400 ;
        RECT 421.950 127.950 427.050 130.050 ;
        RECT 430.950 127.950 433.050 133.050 ;
        RECT 436.950 132.450 439.050 133.200 ;
        RECT 635.400 133.050 636.450 134.400 ;
        RECT 646.950 134.400 667.050 135.450 ;
        RECT 646.950 133.950 649.050 134.400 ;
        RECT 664.950 133.950 667.050 134.400 ;
        RECT 706.950 133.950 712.050 136.050 ;
        RECT 718.950 135.450 721.050 136.050 ;
        RECT 727.800 135.450 729.900 136.050 ;
        RECT 718.950 134.400 729.900 135.450 ;
        RECT 718.950 133.950 721.050 134.400 ;
        RECT 727.800 133.950 729.900 134.400 ;
        RECT 731.100 135.450 733.200 136.050 ;
        RECT 754.950 135.450 757.050 136.050 ;
        RECT 731.100 134.400 757.050 135.450 ;
        RECT 731.100 133.950 733.200 134.400 ;
        RECT 754.950 133.950 757.050 134.400 ;
        RECT 778.950 135.450 781.050 136.050 ;
        RECT 790.950 135.450 793.050 136.050 ;
        RECT 778.950 134.400 793.050 135.450 ;
        RECT 778.950 133.950 781.050 134.400 ;
        RECT 790.950 133.950 793.050 134.400 ;
        RECT 796.950 133.950 802.050 136.050 ;
        RECT 808.950 135.450 811.050 136.050 ;
        RECT 814.950 135.450 817.050 136.050 ;
        RECT 808.950 134.400 817.050 135.450 ;
        RECT 808.950 133.950 811.050 134.400 ;
        RECT 814.950 133.950 817.050 134.400 ;
        RECT 445.950 132.450 448.050 133.050 ;
        RECT 436.950 131.400 448.050 132.450 ;
        RECT 436.950 131.100 439.050 131.400 ;
        RECT 445.950 130.950 448.050 131.400 ;
        RECT 463.800 132.000 465.900 133.050 ;
        RECT 463.800 130.950 466.050 132.000 ;
        RECT 463.950 130.050 466.050 130.950 ;
        RECT 436.950 129.450 439.050 129.900 ;
        RECT 445.950 129.450 448.050 130.050 ;
        RECT 436.950 128.400 448.050 129.450 ;
        RECT 436.950 127.800 439.050 128.400 ;
        RECT 445.950 127.950 448.050 128.400 ;
        RECT 463.800 129.000 466.050 130.050 ;
        RECT 467.100 129.000 469.200 130.050 ;
        RECT 463.800 127.950 465.900 129.000 ;
        RECT 466.950 127.950 469.200 129.000 ;
        RECT 497.100 129.450 499.200 130.050 ;
        RECT 505.950 129.450 508.050 130.050 ;
        RECT 497.100 128.400 508.050 129.450 ;
        RECT 497.100 127.950 499.200 128.400 ;
        RECT 505.950 127.950 508.050 128.400 ;
        RECT 511.950 129.450 514.050 130.050 ;
        RECT 511.950 129.000 528.600 129.450 ;
        RECT 511.950 128.400 529.050 129.000 ;
        RECT 511.950 127.950 514.050 128.400 ;
        RECT 379.950 127.050 382.050 127.200 ;
        RECT 190.950 124.050 193.050 124.950 ;
        RECT 112.950 123.000 132.450 123.450 ;
        RECT 97.950 121.950 100.200 123.000 ;
        RECT 113.400 122.400 132.450 123.000 ;
        RECT 145.950 123.450 148.050 124.050 ;
        RECT 154.800 123.450 156.900 124.050 ;
        RECT 145.950 122.400 156.900 123.450 ;
        RECT 145.950 121.950 148.050 122.400 ;
        RECT 154.800 121.950 156.900 122.400 ;
        RECT 157.800 123.000 160.050 124.050 ;
        RECT 161.100 123.450 163.200 124.050 ;
        RECT 169.800 123.450 171.900 124.050 ;
        RECT 157.800 121.950 159.900 123.000 ;
        RECT 161.100 122.400 171.900 123.450 ;
        RECT 172.950 123.000 175.200 124.050 ;
        RECT 161.100 121.950 163.200 122.400 ;
        RECT 169.800 121.950 171.900 122.400 ;
        RECT 173.100 121.950 175.200 123.000 ;
        RECT 178.950 121.950 184.050 124.050 ;
        RECT 190.800 123.000 193.050 124.050 ;
        RECT 194.100 123.000 196.200 124.050 ;
        RECT 190.800 121.950 192.900 123.000 ;
        RECT 193.950 121.950 196.200 123.000 ;
        RECT 34.950 120.450 37.050 121.050 ;
        RECT 64.950 120.450 67.050 121.050 ;
        RECT 34.950 119.400 67.050 120.450 ;
        RECT 97.950 120.450 100.050 121.950 ;
        RECT 121.950 120.450 124.050 121.050 ;
        RECT 97.950 120.000 124.050 120.450 ;
        RECT 98.550 119.400 124.050 120.000 ;
        RECT 34.950 118.950 37.050 119.400 ;
        RECT 64.950 118.950 67.050 119.400 ;
        RECT 121.950 118.950 124.050 119.400 ;
        RECT 130.950 120.450 133.050 121.050 ;
        RECT 145.950 120.450 148.050 121.050 ;
        RECT 175.950 120.450 178.050 121.050 ;
        RECT 130.950 119.400 148.050 120.450 ;
        RECT 130.950 118.950 133.050 119.400 ;
        RECT 145.950 118.950 148.050 119.400 ;
        RECT 149.400 119.400 178.050 120.450 ;
        RECT 31.950 117.450 34.050 118.050 ;
        RECT 103.950 117.450 106.050 118.050 ;
        RECT 149.400 117.450 150.450 119.400 ;
        RECT 175.950 118.950 178.050 119.400 ;
        RECT 184.950 120.450 187.050 121.050 ;
        RECT 193.950 120.450 196.050 121.950 ;
        RECT 199.950 121.050 202.050 124.050 ;
        RECT 232.950 121.950 238.050 124.050 ;
        RECT 184.950 120.000 196.050 120.450 ;
        RECT 196.950 120.450 202.050 121.050 ;
        RECT 214.950 120.450 217.050 121.050 ;
        RECT 226.950 120.450 229.050 121.050 ;
        RECT 184.950 119.400 195.450 120.000 ;
        RECT 196.950 119.400 229.050 120.450 ;
        RECT 184.950 118.950 187.050 119.400 ;
        RECT 196.950 118.950 201.000 119.400 ;
        RECT 214.950 118.950 217.050 119.400 ;
        RECT 226.950 118.950 229.050 119.400 ;
        RECT 238.950 120.450 241.050 121.050 ;
        RECT 244.950 120.450 247.050 124.050 ;
        RECT 250.950 121.950 256.050 124.050 ;
        RECT 262.950 121.950 268.050 124.050 ;
        RECT 274.950 123.450 277.050 124.050 ;
        RECT 280.800 123.450 282.900 124.050 ;
        RECT 274.950 123.000 282.900 123.450 ;
        RECT 274.950 122.400 283.050 123.000 ;
        RECT 274.950 121.950 277.050 122.400 ;
        RECT 280.800 121.950 283.050 122.400 ;
        RECT 284.100 121.950 289.050 124.050 ;
        RECT 238.950 120.000 247.050 120.450 ;
        RECT 238.950 119.400 246.450 120.000 ;
        RECT 238.950 118.950 241.050 119.400 ;
        RECT 31.950 116.400 150.450 117.450 ;
        RECT 190.950 117.450 193.050 118.050 ;
        RECT 238.950 117.450 241.050 118.050 ;
        RECT 247.950 117.450 250.050 121.050 ;
        RECT 268.950 118.950 274.050 121.050 ;
        RECT 280.950 118.950 283.050 121.950 ;
        RECT 304.950 120.450 307.050 124.050 ;
        RECT 310.950 123.450 316.050 124.050 ;
        RECT 322.950 123.450 325.050 127.050 ;
        RECT 328.950 124.950 334.050 127.050 ;
        RECT 346.950 124.950 352.050 127.050 ;
        RECT 379.950 125.100 385.050 127.050 ;
        RECT 381.000 124.950 385.050 125.100 ;
        RECT 392.100 126.450 394.200 127.050 ;
        RECT 403.950 126.450 406.050 127.050 ;
        RECT 392.100 125.400 406.050 126.450 ;
        RECT 392.100 124.950 394.200 125.400 ;
        RECT 403.950 124.950 406.050 125.400 ;
        RECT 409.950 126.450 412.050 127.050 ;
        RECT 415.950 126.450 418.050 127.050 ;
        RECT 409.950 125.400 418.050 126.450 ;
        RECT 409.950 124.950 412.050 125.400 ;
        RECT 415.950 124.950 418.050 125.400 ;
        RECT 427.950 124.950 433.050 127.050 ;
        RECT 310.950 123.000 325.050 123.450 ;
        RECT 310.950 122.400 324.450 123.000 ;
        RECT 310.950 121.950 316.050 122.400 ;
        RECT 340.950 121.950 346.050 124.050 ;
        RECT 352.950 123.450 355.050 124.050 ;
        RECT 361.950 123.450 364.050 124.050 ;
        RECT 352.950 122.400 364.050 123.450 ;
        RECT 352.950 121.950 355.050 122.400 ;
        RECT 361.950 121.950 364.050 122.400 ;
        RECT 376.950 121.950 382.050 124.050 ;
        RECT 319.950 120.450 322.050 121.050 ;
        RECT 304.950 120.000 322.050 120.450 ;
        RECT 305.400 119.400 322.050 120.000 ;
        RECT 319.950 118.950 322.050 119.400 ;
        RECT 385.950 118.950 388.050 124.050 ;
        RECT 397.950 121.950 403.050 124.050 ;
        RECT 406.950 123.450 409.050 124.050 ;
        RECT 439.950 123.450 442.050 127.050 ;
        RECT 445.950 126.450 448.050 127.050 ;
        RECT 451.950 126.450 454.050 127.050 ;
        RECT 445.950 125.400 454.050 126.450 ;
        RECT 445.950 124.950 448.050 125.400 ;
        RECT 451.950 124.950 454.050 125.400 ;
        RECT 457.950 124.950 463.050 127.050 ;
        RECT 466.950 124.950 469.050 127.950 ;
        RECT 475.950 126.450 478.050 127.050 ;
        RECT 484.950 126.450 489.900 127.050 ;
        RECT 475.950 125.400 489.900 126.450 ;
        RECT 475.950 124.950 478.050 125.400 ;
        RECT 484.950 124.950 489.900 125.400 ;
        RECT 406.950 123.000 442.050 123.450 ;
        RECT 442.950 123.450 445.050 124.050 ;
        RECT 448.950 123.450 451.050 124.050 ;
        RECT 406.950 122.400 441.450 123.000 ;
        RECT 442.950 122.400 451.050 123.450 ;
        RECT 406.950 121.950 409.050 122.400 ;
        RECT 442.950 121.950 445.050 122.400 ;
        RECT 448.950 121.950 451.050 122.400 ;
        RECT 472.950 123.450 475.050 124.050 ;
        RECT 499.950 123.450 502.050 127.050 ;
        RECT 505.950 126.450 508.050 127.050 ;
        RECT 517.950 126.450 520.050 127.050 ;
        RECT 523.800 126.450 525.900 127.200 ;
        RECT 505.950 125.400 525.900 126.450 ;
        RECT 526.950 127.050 529.050 128.400 ;
        RECT 535.950 127.950 541.050 130.050 ;
        RECT 562.950 129.450 565.050 130.050 ;
        RECT 580.950 129.450 583.050 130.050 ;
        RECT 562.950 128.400 583.050 129.450 ;
        RECT 562.950 127.950 565.050 128.400 ;
        RECT 580.950 127.950 583.050 128.400 ;
        RECT 598.950 127.950 601.050 133.050 ;
        RECT 604.950 127.950 607.050 133.050 ;
        RECT 616.950 127.950 619.050 133.050 ;
        RECT 634.950 132.450 637.050 133.050 ;
        RECT 742.950 132.450 745.050 133.050 ;
        RECT 775.950 132.450 778.050 133.050 ;
        RECT 634.950 131.400 745.050 132.450 ;
        RECT 634.950 130.950 637.050 131.400 ;
        RECT 742.950 130.950 745.050 131.400 ;
        RECT 746.400 131.400 778.050 132.450 ;
        RECT 622.950 127.950 628.050 130.050 ;
        RECT 709.950 129.450 712.050 130.050 ;
        RECT 695.400 129.000 712.050 129.450 ;
        RECT 694.950 128.400 712.050 129.000 ;
        RECT 526.950 126.000 529.200 127.050 ;
        RECT 505.950 124.950 508.050 125.400 ;
        RECT 517.950 124.950 520.050 125.400 ;
        RECT 523.800 125.100 525.900 125.400 ;
        RECT 527.100 124.950 529.200 126.000 ;
        RECT 532.950 126.450 535.050 127.050 ;
        RECT 538.800 126.450 540.900 127.050 ;
        RECT 532.950 125.400 540.900 126.450 ;
        RECT 542.100 126.000 544.200 127.050 ;
        RECT 532.950 124.950 535.050 125.400 ;
        RECT 538.800 124.950 540.900 125.400 ;
        RECT 541.950 124.950 544.200 126.000 ;
        RECT 559.950 126.450 562.050 127.050 ;
        RECT 577.950 126.450 580.050 127.050 ;
        RECT 559.950 125.400 580.050 126.450 ;
        RECT 559.950 124.950 562.050 125.400 ;
        RECT 577.950 124.950 580.050 125.400 ;
        RECT 583.950 124.950 589.050 127.050 ;
        RECT 601.950 126.450 604.050 127.050 ;
        RECT 607.950 126.450 610.050 127.050 ;
        RECT 601.950 125.400 610.050 126.450 ;
        RECT 601.950 124.950 604.050 125.400 ;
        RECT 607.950 124.950 610.050 125.400 ;
        RECT 619.950 124.950 622.050 127.050 ;
        RECT 628.950 124.950 633.900 127.050 ;
        RECT 634.800 126.000 636.900 127.050 ;
        RECT 638.100 126.450 640.200 127.050 ;
        RECT 652.950 126.450 655.050 127.050 ;
        RECT 634.800 124.950 637.050 126.000 ;
        RECT 638.100 125.400 655.050 126.450 ;
        RECT 638.100 124.950 640.200 125.400 ;
        RECT 652.950 124.950 655.050 125.400 ;
        RECT 658.950 124.950 664.050 127.050 ;
        RECT 667.950 124.950 672.900 127.050 ;
        RECT 674.100 124.950 679.050 127.050 ;
        RECT 694.950 124.950 697.050 128.400 ;
        RECT 709.950 127.950 712.050 128.400 ;
        RECT 715.950 127.950 721.050 130.050 ;
        RECT 736.950 129.450 739.050 130.050 ;
        RECT 746.400 129.450 747.450 131.400 ;
        RECT 775.950 130.950 778.050 131.400 ;
        RECT 778.950 129.450 781.050 130.050 ;
        RECT 736.950 128.400 747.450 129.450 ;
        RECT 770.400 129.000 781.050 129.450 ;
        RECT 769.950 128.400 781.050 129.000 ;
        RECT 736.950 127.950 739.050 128.400 ;
        RECT 715.950 126.900 720.000 127.050 ;
        RECT 715.950 124.950 720.900 126.900 ;
        RECT 722.100 126.450 727.050 127.050 ;
        RECT 748.800 126.450 750.900 127.050 ;
        RECT 722.100 125.400 750.900 126.450 ;
        RECT 722.100 124.950 727.050 125.400 ;
        RECT 748.800 124.950 750.900 125.400 ;
        RECT 752.100 126.450 754.200 127.050 ;
        RECT 763.950 126.450 766.050 127.050 ;
        RECT 752.100 125.400 766.050 126.450 ;
        RECT 752.100 124.950 754.200 125.400 ;
        RECT 763.950 124.950 766.050 125.400 ;
        RECT 769.950 124.950 772.050 128.400 ;
        RECT 778.950 127.950 781.050 128.400 ;
        RECT 784.950 127.950 787.050 133.050 ;
        RECT 802.950 132.450 805.050 133.050 ;
        RECT 820.950 132.450 823.050 133.050 ;
        RECT 802.950 131.400 823.050 132.450 ;
        RECT 802.950 130.950 805.050 131.400 ;
        RECT 820.950 130.950 823.050 131.400 ;
        RECT 829.950 132.450 832.050 133.050 ;
        RECT 850.950 132.450 853.050 133.050 ;
        RECT 829.950 131.400 853.050 132.450 ;
        RECT 829.950 130.950 832.050 131.400 ;
        RECT 850.950 130.950 853.050 131.400 ;
        RECT 790.950 127.950 796.050 130.050 ;
        RECT 775.950 126.450 778.050 127.050 ;
        RECT 787.950 126.450 790.050 127.050 ;
        RECT 775.950 125.400 790.050 126.450 ;
        RECT 775.950 124.950 778.050 125.400 ;
        RECT 787.950 124.950 790.050 125.400 ;
        RECT 802.950 124.950 805.050 130.050 ;
        RECT 814.950 129.450 817.050 130.050 ;
        RECT 838.950 129.450 841.050 130.050 ;
        RECT 809.400 129.000 817.050 129.450 ;
        RECT 830.400 129.000 846.450 129.450 ;
        RECT 808.950 128.400 817.050 129.000 ;
        RECT 808.950 124.950 811.050 128.400 ;
        RECT 814.950 127.950 817.050 128.400 ;
        RECT 829.950 128.400 846.450 129.000 ;
        RECT 820.950 124.950 826.050 127.050 ;
        RECT 829.950 124.950 832.050 128.400 ;
        RECT 838.950 127.950 841.050 128.400 ;
        RECT 845.400 127.050 846.450 128.400 ;
        RECT 844.950 126.450 847.050 127.050 ;
        RECT 850.950 126.450 853.050 127.050 ;
        RECT 844.950 125.400 853.050 126.450 ;
        RECT 844.950 124.950 847.050 125.400 ;
        RECT 850.950 124.950 853.050 125.400 ;
        RECT 472.950 123.000 502.050 123.450 ;
        RECT 472.950 122.400 501.450 123.000 ;
        RECT 472.950 121.950 475.050 122.400 ;
        RECT 502.950 121.050 505.050 124.050 ;
        RECT 511.950 121.950 517.050 124.050 ;
        RECT 523.950 121.950 528.900 124.050 ;
        RECT 530.100 123.450 532.200 124.050 ;
        RECT 541.950 123.450 544.050 124.950 ;
        RECT 530.100 123.000 544.050 123.450 ;
        RECT 568.950 123.450 571.050 124.050 ;
        RECT 574.950 123.450 577.050 124.050 ;
        RECT 530.100 122.400 543.450 123.000 ;
        RECT 568.950 122.400 577.050 123.450 ;
        RECT 530.100 121.950 532.200 122.400 ;
        RECT 568.950 121.950 571.050 122.400 ;
        RECT 574.950 121.950 577.050 122.400 ;
        RECT 580.950 123.450 583.050 124.050 ;
        RECT 592.950 123.450 595.050 124.050 ;
        RECT 580.950 122.400 595.050 123.450 ;
        RECT 580.950 121.950 583.050 122.400 ;
        RECT 592.950 121.950 595.050 122.400 ;
        RECT 421.950 120.450 424.050 121.050 ;
        RECT 442.950 120.450 445.050 121.050 ;
        RECT 421.950 119.400 445.050 120.450 ;
        RECT 421.950 118.950 424.050 119.400 ;
        RECT 442.950 118.950 445.050 119.400 ;
        RECT 502.800 120.000 505.050 121.050 ;
        RECT 506.100 120.450 508.200 121.050 ;
        RECT 517.950 120.450 520.050 121.050 ;
        RECT 502.800 118.950 504.900 120.000 ;
        RECT 506.100 119.400 520.050 120.450 ;
        RECT 506.100 118.950 508.200 119.400 ;
        RECT 517.950 118.950 520.050 119.400 ;
        RECT 550.950 120.450 553.050 121.050 ;
        RECT 604.950 120.450 607.050 121.050 ;
        RECT 620.400 120.450 621.450 124.950 ;
        RECT 634.950 121.950 637.050 124.950 ;
        RECT 718.800 124.800 720.900 124.950 ;
        RECT 640.950 121.950 646.050 124.050 ;
        RECT 673.950 123.450 676.050 124.050 ;
        RECT 668.400 122.400 676.050 123.450 ;
        RECT 668.400 121.050 669.450 122.400 ;
        RECT 673.950 121.950 676.050 122.400 ;
        RECT 550.950 119.400 621.450 120.450 ;
        RECT 622.950 120.450 625.050 121.050 ;
        RECT 646.950 120.450 649.050 121.050 ;
        RECT 622.950 119.400 649.050 120.450 ;
        RECT 550.950 118.950 553.050 119.400 ;
        RECT 604.950 118.950 607.050 119.400 ;
        RECT 622.950 118.950 625.050 119.400 ;
        RECT 646.950 118.950 649.050 119.400 ;
        RECT 652.950 120.450 655.050 121.050 ;
        RECT 658.950 120.450 663.900 121.050 ;
        RECT 652.950 119.400 663.900 120.450 ;
        RECT 652.950 118.950 655.050 119.400 ;
        RECT 658.950 118.950 663.900 119.400 ;
        RECT 665.100 119.400 669.450 121.050 ;
        RECT 679.950 120.450 682.050 124.050 ;
        RECT 700.950 121.950 706.050 124.050 ;
        RECT 757.950 123.450 760.050 124.050 ;
        RECT 766.950 123.450 769.050 124.050 ;
        RECT 757.950 122.400 769.050 123.450 ;
        RECT 757.950 121.950 760.050 122.400 ;
        RECT 766.950 121.950 769.050 122.400 ;
        RECT 772.950 123.450 775.050 124.050 ;
        RECT 805.800 123.450 807.900 124.050 ;
        RECT 772.950 122.400 807.900 123.450 ;
        RECT 772.950 121.950 775.050 122.400 ;
        RECT 805.800 121.950 807.900 122.400 ;
        RECT 809.100 121.950 813.900 124.050 ;
        RECT 815.100 123.450 817.200 124.050 ;
        RECT 826.800 123.450 828.900 124.050 ;
        RECT 815.100 122.400 828.900 123.450 ;
        RECT 815.100 121.950 817.200 122.400 ;
        RECT 826.800 121.950 828.900 122.400 ;
        RECT 830.100 121.950 835.050 124.050 ;
        RECT 841.950 121.950 846.900 124.050 ;
        RECT 848.100 123.000 850.200 124.050 ;
        RECT 847.950 121.950 850.200 123.000 ;
        RECT 694.950 120.450 697.050 121.050 ;
        RECT 679.950 120.000 697.050 120.450 ;
        RECT 680.400 119.400 697.050 120.000 ;
        RECT 665.100 118.950 669.000 119.400 ;
        RECT 694.950 118.950 697.050 119.400 ;
        RECT 268.950 117.450 271.050 118.050 ;
        RECT 190.950 116.400 225.450 117.450 ;
        RECT 31.950 115.950 34.050 116.400 ;
        RECT 103.950 115.950 106.050 116.400 ;
        RECT 190.950 115.950 193.050 116.400 ;
        RECT 224.400 115.050 225.450 116.400 ;
        RECT 238.950 116.400 271.050 117.450 ;
        RECT 238.950 115.950 241.050 116.400 ;
        RECT 268.950 115.950 271.050 116.400 ;
        RECT 292.950 117.450 295.050 118.050 ;
        RECT 331.950 117.450 334.050 118.050 ;
        RECT 292.950 116.400 334.050 117.450 ;
        RECT 292.950 115.950 295.050 116.400 ;
        RECT 331.950 115.950 334.050 116.400 ;
        RECT 337.950 117.450 340.050 118.050 ;
        RECT 364.950 117.450 367.050 118.050 ;
        RECT 337.950 116.400 367.050 117.450 ;
        RECT 337.950 115.950 340.050 116.400 ;
        RECT 364.950 115.950 367.050 116.400 ;
        RECT 370.950 117.450 373.050 118.050 ;
        RECT 400.950 117.450 403.050 118.050 ;
        RECT 370.950 116.400 403.050 117.450 ;
        RECT 370.950 115.950 373.050 116.400 ;
        RECT 400.950 115.950 403.050 116.400 ;
        RECT 409.950 117.450 412.050 118.050 ;
        RECT 424.950 117.450 427.050 118.050 ;
        RECT 409.950 116.400 427.050 117.450 ;
        RECT 409.950 115.950 412.050 116.400 ;
        RECT 424.950 115.950 427.050 116.400 ;
        RECT 448.950 117.450 451.050 118.050 ;
        RECT 532.950 117.450 535.050 118.050 ;
        RECT 448.950 116.400 535.050 117.450 ;
        RECT 448.950 115.950 451.050 116.400 ;
        RECT 532.950 115.950 535.050 116.400 ;
        RECT 667.950 117.450 670.050 118.050 ;
        RECT 688.950 117.450 691.050 118.050 ;
        RECT 667.950 116.400 691.050 117.450 ;
        RECT 736.950 117.450 739.050 121.050 ;
        RECT 748.950 118.950 754.050 121.050 ;
        RECT 778.950 120.450 781.050 121.050 ;
        RECT 802.950 120.450 805.050 121.050 ;
        RECT 778.950 119.400 805.050 120.450 ;
        RECT 778.950 118.950 781.050 119.400 ;
        RECT 802.950 118.950 805.050 119.400 ;
        RECT 823.950 120.450 826.050 121.050 ;
        RECT 847.950 120.450 850.050 121.950 ;
        RECT 823.950 120.000 850.050 120.450 ;
        RECT 823.950 119.400 849.450 120.000 ;
        RECT 823.950 118.950 826.050 119.400 ;
        RECT 772.950 117.450 775.050 118.050 ;
        RECT 736.950 117.000 775.050 117.450 ;
        RECT 737.400 116.400 775.050 117.000 ;
        RECT 667.950 115.950 670.050 116.400 ;
        RECT 688.950 115.950 691.050 116.400 ;
        RECT 772.950 115.950 775.050 116.400 ;
        RECT 25.950 114.450 28.050 115.050 ;
        RECT 67.950 114.450 70.050 115.050 ;
        RECT 25.950 113.400 70.050 114.450 ;
        RECT 25.950 112.950 28.050 113.400 ;
        RECT 67.950 112.950 70.050 113.400 ;
        RECT 91.950 114.450 94.050 115.050 ;
        RECT 109.950 114.450 112.050 115.050 ;
        RECT 121.950 114.450 124.050 115.050 ;
        RECT 91.950 113.400 124.050 114.450 ;
        RECT 91.950 112.950 94.050 113.400 ;
        RECT 109.950 112.950 112.050 113.400 ;
        RECT 121.950 112.950 124.050 113.400 ;
        RECT 127.950 114.450 130.050 115.050 ;
        RECT 139.800 114.450 141.900 115.050 ;
        RECT 127.950 113.400 141.900 114.450 ;
        RECT 127.950 112.950 130.050 113.400 ;
        RECT 139.800 112.950 141.900 113.400 ;
        RECT 143.100 114.450 145.200 115.050 ;
        RECT 157.950 114.450 160.050 115.050 ;
        RECT 172.950 114.450 175.050 115.050 ;
        RECT 143.100 113.400 175.050 114.450 ;
        RECT 143.100 112.950 145.200 113.400 ;
        RECT 157.950 112.950 160.050 113.400 ;
        RECT 172.950 112.950 175.050 113.400 ;
        RECT 223.950 114.450 226.050 115.050 ;
        RECT 295.950 114.450 298.050 115.050 ;
        RECT 223.950 113.400 298.050 114.450 ;
        RECT 223.950 112.950 226.050 113.400 ;
        RECT 295.950 112.950 298.050 113.400 ;
        RECT 304.950 114.450 307.050 115.050 ;
        RECT 379.950 114.450 382.050 115.050 ;
        RECT 304.950 113.400 382.050 114.450 ;
        RECT 304.950 112.950 307.050 113.400 ;
        RECT 379.950 112.950 382.050 113.400 ;
        RECT 418.950 114.450 421.050 115.050 ;
        RECT 436.950 114.450 439.050 115.050 ;
        RECT 418.950 113.400 439.050 114.450 ;
        RECT 418.950 112.950 421.050 113.400 ;
        RECT 436.950 112.950 439.050 113.400 ;
        RECT 475.950 114.450 478.050 115.050 ;
        RECT 481.950 114.450 484.050 115.050 ;
        RECT 475.950 113.400 484.050 114.450 ;
        RECT 475.950 112.950 478.050 113.400 ;
        RECT 481.950 112.950 484.050 113.400 ;
        RECT 517.950 112.950 523.050 115.050 ;
        RECT 526.950 114.450 529.050 115.050 ;
        RECT 538.950 114.450 541.050 115.050 ;
        RECT 526.950 113.400 541.050 114.450 ;
        RECT 526.950 112.950 529.050 113.400 ;
        RECT 538.950 112.950 541.050 113.400 ;
        RECT 580.950 114.450 583.050 115.050 ;
        RECT 685.950 114.450 688.050 115.050 ;
        RECT 580.950 113.400 688.050 114.450 ;
        RECT 580.950 112.950 583.050 113.400 ;
        RECT 685.950 112.950 688.050 113.400 ;
        RECT 706.950 114.450 709.050 115.050 ;
        RECT 733.950 114.450 736.050 115.050 ;
        RECT 706.950 113.400 736.050 114.450 ;
        RECT 706.950 112.950 709.050 113.400 ;
        RECT 733.950 112.950 736.050 113.400 ;
        RECT 748.950 114.450 751.050 115.050 ;
        RECT 796.950 114.450 799.050 115.050 ;
        RECT 748.950 113.400 799.050 114.450 ;
        RECT 748.950 112.950 751.050 113.400 ;
        RECT 796.950 112.950 799.050 113.400 ;
        RECT 817.950 114.450 820.050 115.050 ;
        RECT 841.950 114.450 844.050 115.050 ;
        RECT 817.950 113.400 844.050 114.450 ;
        RECT 817.950 112.950 820.050 113.400 ;
        RECT 841.950 112.950 844.050 113.400 ;
        RECT 52.950 111.450 55.050 112.050 ;
        RECT 73.950 111.450 76.050 112.050 ;
        RECT 232.950 111.450 235.050 112.050 ;
        RECT 289.950 111.450 292.050 112.050 ;
        RECT 52.950 110.400 235.050 111.450 ;
        RECT 52.950 109.950 55.050 110.400 ;
        RECT 73.950 109.950 76.050 110.400 ;
        RECT 232.950 109.950 235.050 110.400 ;
        RECT 236.400 110.400 292.050 111.450 ;
        RECT 136.950 108.450 139.050 109.050 ;
        RECT 151.950 108.450 154.050 109.050 ;
        RECT 136.950 107.400 154.050 108.450 ;
        RECT 136.950 106.950 139.050 107.400 ;
        RECT 151.950 106.950 154.050 107.400 ;
        RECT 196.950 108.450 199.050 109.050 ;
        RECT 236.400 108.450 237.450 110.400 ;
        RECT 289.950 109.950 292.050 110.400 ;
        RECT 307.950 111.450 310.050 112.050 ;
        RECT 385.950 111.450 388.050 112.050 ;
        RECT 472.950 111.450 475.050 112.050 ;
        RECT 307.950 110.400 360.450 111.450 ;
        RECT 307.950 109.950 310.050 110.400 ;
        RECT 196.950 107.400 237.450 108.450 ;
        RECT 359.400 108.450 360.450 110.400 ;
        RECT 385.950 110.400 475.050 111.450 ;
        RECT 385.950 109.950 388.050 110.400 ;
        RECT 472.950 109.950 475.050 110.400 ;
        RECT 484.950 111.450 487.050 112.050 ;
        RECT 496.950 111.450 499.050 112.050 ;
        RECT 484.950 110.400 499.050 111.450 ;
        RECT 484.950 109.950 487.050 110.400 ;
        RECT 496.950 109.950 499.050 110.400 ;
        RECT 502.950 111.450 505.050 112.050 ;
        RECT 523.950 111.450 526.050 112.050 ;
        RECT 502.950 110.400 526.050 111.450 ;
        RECT 502.950 109.950 505.050 110.400 ;
        RECT 523.950 109.950 526.050 110.400 ;
        RECT 592.950 111.450 595.050 112.050 ;
        RECT 664.950 111.450 667.050 112.050 ;
        RECT 592.950 110.400 667.050 111.450 ;
        RECT 592.950 109.950 595.050 110.400 ;
        RECT 664.950 109.950 667.050 110.400 ;
        RECT 670.950 111.450 673.050 112.050 ;
        RECT 679.950 111.450 682.050 112.050 ;
        RECT 670.950 110.400 682.050 111.450 ;
        RECT 670.950 109.950 673.050 110.400 ;
        RECT 679.950 109.950 682.050 110.400 ;
        RECT 739.950 111.450 742.050 112.050 ;
        RECT 811.950 111.450 814.050 112.050 ;
        RECT 739.950 110.400 814.050 111.450 ;
        RECT 739.950 109.950 742.050 110.400 ;
        RECT 811.950 109.950 814.050 110.400 ;
        RECT 409.950 108.450 412.050 109.050 ;
        RECT 359.400 107.400 412.050 108.450 ;
        RECT 196.950 106.950 199.050 107.400 ;
        RECT 409.950 106.950 412.050 107.400 ;
        RECT 415.950 108.450 418.050 109.050 ;
        RECT 511.950 108.450 514.050 109.050 ;
        RECT 415.950 107.400 514.050 108.450 ;
        RECT 415.950 106.950 418.050 107.400 ;
        RECT 511.950 106.950 514.050 107.400 ;
        RECT 589.950 108.450 592.050 109.050 ;
        RECT 598.950 108.450 601.050 109.050 ;
        RECT 589.950 107.400 601.050 108.450 ;
        RECT 589.950 106.950 592.050 107.400 ;
        RECT 598.950 106.950 601.050 107.400 ;
        RECT 655.950 108.450 658.050 109.050 ;
        RECT 712.950 108.450 715.050 109.050 ;
        RECT 655.950 107.400 715.050 108.450 ;
        RECT 655.950 106.950 658.050 107.400 ;
        RECT 712.950 106.950 715.050 107.400 ;
        RECT 730.950 108.450 733.050 109.050 ;
        RECT 790.950 108.450 793.050 109.050 ;
        RECT 730.950 107.400 793.050 108.450 ;
        RECT 730.950 106.950 733.050 107.400 ;
        RECT 790.950 106.950 793.050 107.400 ;
        RECT 799.950 108.450 802.050 109.050 ;
        RECT 847.950 108.450 850.050 109.050 ;
        RECT 799.950 107.400 850.050 108.450 ;
        RECT 799.950 106.950 802.050 107.400 ;
        RECT 847.950 106.950 850.050 107.400 ;
        RECT 13.950 105.450 16.050 106.050 ;
        RECT 49.950 105.450 52.050 106.050 ;
        RECT 13.950 104.400 52.050 105.450 ;
        RECT 13.950 103.950 16.050 104.400 ;
        RECT 49.950 103.950 52.050 104.400 ;
        RECT 112.950 105.450 115.050 106.050 ;
        RECT 148.950 105.450 151.050 106.050 ;
        RECT 184.950 105.450 187.050 106.050 ;
        RECT 112.950 104.400 187.050 105.450 ;
        RECT 112.950 103.950 115.050 104.400 ;
        RECT 148.950 103.950 151.050 104.400 ;
        RECT 184.950 103.950 187.050 104.400 ;
        RECT 217.950 105.450 220.050 106.050 ;
        RECT 244.950 105.450 247.050 106.050 ;
        RECT 217.950 104.400 247.050 105.450 ;
        RECT 217.950 103.950 220.050 104.400 ;
        RECT 244.950 103.950 247.050 104.400 ;
        RECT 262.950 105.450 265.050 106.050 ;
        RECT 322.950 105.450 325.050 106.050 ;
        RECT 262.950 104.400 325.050 105.450 ;
        RECT 262.950 103.950 265.050 104.400 ;
        RECT 322.950 103.950 325.050 104.400 ;
        RECT 331.950 105.450 334.050 106.050 ;
        RECT 391.950 105.450 394.050 106.050 ;
        RECT 331.950 104.400 394.050 105.450 ;
        RECT 331.950 103.950 334.050 104.400 ;
        RECT 391.950 103.950 394.050 104.400 ;
        RECT 397.950 105.450 400.050 106.050 ;
        RECT 403.950 105.450 406.050 106.050 ;
        RECT 451.950 105.450 454.050 106.050 ;
        RECT 397.950 104.400 406.050 105.450 ;
        RECT 397.950 103.950 400.050 104.400 ;
        RECT 403.950 103.950 406.050 104.400 ;
        RECT 428.400 104.400 454.050 105.450 ;
        RECT 428.400 103.050 429.450 104.400 ;
        RECT 451.950 103.950 454.050 104.400 ;
        RECT 499.950 105.450 502.050 106.050 ;
        RECT 508.950 105.450 511.050 106.050 ;
        RECT 499.950 104.400 511.050 105.450 ;
        RECT 499.950 103.950 502.050 104.400 ;
        RECT 508.950 103.950 511.050 104.400 ;
        RECT 574.950 105.450 577.050 106.050 ;
        RECT 625.950 105.450 628.050 106.050 ;
        RECT 574.950 104.400 628.050 105.450 ;
        RECT 574.950 103.950 577.050 104.400 ;
        RECT 625.950 103.950 628.050 104.400 ;
        RECT 640.950 105.450 643.050 106.050 ;
        RECT 676.950 105.450 679.050 106.050 ;
        RECT 700.950 105.450 703.050 106.050 ;
        RECT 640.950 104.400 703.050 105.450 ;
        RECT 640.950 103.950 643.050 104.400 ;
        RECT 676.950 103.950 679.050 104.400 ;
        RECT 700.950 103.950 703.050 104.400 ;
        RECT 718.950 105.450 721.050 106.050 ;
        RECT 727.950 105.450 730.050 106.050 ;
        RECT 718.950 104.400 730.050 105.450 ;
        RECT 718.950 103.950 721.050 104.400 ;
        RECT 727.950 103.950 730.050 104.400 ;
        RECT 754.950 105.450 757.050 106.050 ;
        RECT 766.950 105.450 769.050 106.050 ;
        RECT 754.950 104.400 769.050 105.450 ;
        RECT 754.950 103.950 757.050 104.400 ;
        RECT 766.950 103.950 769.050 104.400 ;
        RECT 796.950 105.450 799.050 106.050 ;
        RECT 808.950 105.450 811.050 106.050 ;
        RECT 796.950 104.400 811.050 105.450 ;
        RECT 796.950 103.950 799.050 104.400 ;
        RECT 808.950 103.950 811.050 104.400 ;
        RECT 13.950 97.950 16.050 103.050 ;
        RECT 46.950 102.450 49.050 103.050 ;
        RECT 82.950 102.450 85.050 103.050 ;
        RECT 46.950 101.400 85.050 102.450 ;
        RECT 46.950 100.950 49.050 101.400 ;
        RECT 82.950 100.950 85.050 101.400 ;
        RECT 88.950 102.450 91.050 103.050 ;
        RECT 160.950 102.450 163.050 103.050 ;
        RECT 88.950 101.400 163.050 102.450 ;
        RECT 88.950 100.950 91.050 101.400 ;
        RECT 160.950 100.950 163.050 101.400 ;
        RECT 169.950 102.450 172.050 103.050 ;
        RECT 181.950 102.450 184.050 103.050 ;
        RECT 169.950 101.400 184.050 102.450 ;
        RECT 169.950 100.950 172.050 101.400 ;
        RECT 181.950 100.950 184.050 101.400 ;
        RECT 208.950 102.450 211.050 103.050 ;
        RECT 238.950 102.450 241.050 103.050 ;
        RECT 208.950 101.400 241.050 102.450 ;
        RECT 208.950 100.950 211.050 101.400 ;
        RECT 238.950 100.950 241.050 101.400 ;
        RECT 28.950 94.950 31.050 100.050 ;
        RECT 36.000 99.450 40.050 100.050 ;
        RECT 112.950 99.450 115.050 100.050 ;
        RECT 35.400 99.000 40.050 99.450 ;
        RECT 95.400 99.000 115.050 99.450 ;
        RECT 34.950 97.950 40.050 99.000 ;
        RECT 94.950 98.400 115.050 99.000 ;
        RECT 34.950 94.950 37.050 97.950 ;
        RECT 55.950 96.450 58.050 97.050 ;
        RECT 67.950 96.450 70.050 97.050 ;
        RECT 55.950 95.400 70.050 96.450 ;
        RECT 52.800 94.050 54.900 94.200 ;
        RECT 13.950 93.450 16.050 94.050 ;
        RECT 25.950 93.450 28.050 94.050 ;
        RECT 13.950 92.400 28.050 93.450 ;
        RECT 13.950 91.950 16.050 92.400 ;
        RECT 25.950 91.950 28.050 92.400 ;
        RECT 31.950 91.950 37.050 94.050 ;
        RECT 49.950 92.100 54.900 94.050 ;
        RECT 55.950 94.050 58.050 95.400 ;
        RECT 67.950 94.950 70.050 95.400 ;
        RECT 76.950 96.450 79.050 97.050 ;
        RECT 88.950 96.450 91.050 97.050 ;
        RECT 76.950 96.000 93.300 96.450 ;
        RECT 76.950 95.400 94.050 96.000 ;
        RECT 76.950 94.950 79.050 95.400 ;
        RECT 88.950 94.950 91.050 95.400 ;
        RECT 91.950 94.050 94.050 95.400 ;
        RECT 94.950 94.950 97.050 98.400 ;
        RECT 112.950 97.950 115.050 98.400 ;
        RECT 100.950 96.450 103.050 97.050 ;
        RECT 154.950 96.450 157.050 97.050 ;
        RECT 100.950 95.400 157.050 96.450 ;
        RECT 100.950 94.950 103.050 95.400 ;
        RECT 154.950 94.950 157.050 95.400 ;
        RECT 160.950 96.450 163.050 100.050 ;
        RECT 184.950 99.450 187.050 100.050 ;
        RECT 176.400 99.000 187.050 99.450 ;
        RECT 175.950 98.400 187.050 99.000 ;
        RECT 169.950 96.450 172.050 97.050 ;
        RECT 160.950 95.400 172.050 96.450 ;
        RECT 160.950 94.950 163.050 95.400 ;
        RECT 169.950 94.950 172.050 95.400 ;
        RECT 175.950 94.950 178.050 98.400 ;
        RECT 184.950 97.950 187.050 98.400 ;
        RECT 187.950 96.450 190.050 97.050 ;
        RECT 196.950 96.450 199.050 97.050 ;
        RECT 187.950 95.400 199.050 96.450 ;
        RECT 187.950 94.950 190.050 95.400 ;
        RECT 196.950 94.950 199.050 95.400 ;
        RECT 202.950 94.950 205.050 100.050 ;
        RECT 229.950 99.450 232.050 100.050 ;
        RECT 250.950 99.450 253.050 100.050 ;
        RECT 229.950 98.400 253.050 99.450 ;
        RECT 229.950 97.950 232.050 98.400 ;
        RECT 241.950 97.050 244.050 98.400 ;
        RECT 250.950 97.950 253.050 98.400 ;
        RECT 274.950 97.950 277.050 103.050 ;
        RECT 364.950 102.450 367.050 103.050 ;
        RECT 427.950 102.450 430.050 103.050 ;
        RECT 364.950 101.400 430.050 102.450 ;
        RECT 364.950 100.950 367.050 101.400 ;
        RECT 427.950 100.950 430.050 101.400 ;
        RECT 445.950 102.450 448.050 103.050 ;
        RECT 466.950 102.450 469.050 103.050 ;
        RECT 445.950 101.400 469.050 102.450 ;
        RECT 445.950 100.950 448.050 101.400 ;
        RECT 466.950 100.950 469.050 101.400 ;
        RECT 490.950 102.450 493.050 103.050 ;
        RECT 502.950 102.450 505.050 103.050 ;
        RECT 538.950 102.450 541.050 103.050 ;
        RECT 559.950 102.450 562.050 103.050 ;
        RECT 490.950 101.400 562.050 102.450 ;
        RECT 490.950 100.950 493.050 101.400 ;
        RECT 502.950 100.950 505.050 101.400 ;
        RECT 538.950 100.950 541.050 101.400 ;
        RECT 559.950 100.950 562.050 101.400 ;
        RECT 595.950 102.450 598.050 103.050 ;
        RECT 646.950 102.450 649.050 103.200 ;
        RECT 670.950 102.450 673.050 103.050 ;
        RECT 595.950 101.400 612.450 102.450 ;
        RECT 595.950 100.950 598.050 101.400 ;
        RECT 322.950 99.450 325.050 100.050 ;
        RECT 355.950 99.450 358.050 100.050 ;
        RECT 367.950 99.450 373.050 100.050 ;
        RECT 322.950 99.000 336.450 99.450 ;
        RECT 322.950 98.400 337.050 99.000 ;
        RECT 322.950 97.950 325.050 98.400 ;
        RECT 223.950 96.450 226.050 97.050 ;
        RECT 218.400 96.000 226.050 96.450 ;
        RECT 217.950 95.400 226.050 96.000 ;
        RECT 55.950 93.000 58.200 94.050 ;
        RECT 49.950 91.950 54.000 92.100 ;
        RECT 56.100 91.950 58.200 93.000 ;
        RECT 46.950 90.450 51.000 91.050 ;
        RECT 52.950 90.450 58.050 91.050 ;
        RECT 64.950 90.450 67.050 94.050 ;
        RECT 70.950 91.950 76.050 94.050 ;
        RECT 91.800 93.000 94.050 94.050 ;
        RECT 91.800 91.950 93.900 93.000 ;
        RECT 95.100 91.950 100.050 94.050 ;
        RECT 109.950 91.950 115.050 94.050 ;
        RECT 118.950 93.450 121.050 94.050 ;
        RECT 127.950 93.450 130.050 94.050 ;
        RECT 118.950 92.400 130.050 93.450 ;
        RECT 118.950 91.950 121.050 92.400 ;
        RECT 127.950 91.950 130.050 92.400 ;
        RECT 46.950 88.950 51.450 90.450 ;
        RECT 52.950 90.000 67.050 90.450 ;
        RECT 52.950 89.400 66.450 90.000 ;
        RECT 52.950 88.950 58.050 89.400 ;
        RECT 103.950 88.950 109.050 91.050 ;
        RECT 28.950 87.450 31.050 88.050 ;
        RECT 46.950 87.450 49.050 88.050 ;
        RECT 28.950 86.400 49.050 87.450 ;
        RECT 50.400 87.450 51.450 88.950 ;
        RECT 94.950 87.450 97.050 88.050 ;
        RECT 115.950 87.450 118.050 91.050 ;
        RECT 133.950 90.450 136.050 94.050 ;
        RECT 139.950 93.450 142.050 94.050 ;
        RECT 145.800 93.450 147.900 94.050 ;
        RECT 139.950 92.400 147.900 93.450 ;
        RECT 139.950 91.950 142.050 92.400 ;
        RECT 145.800 91.950 147.900 92.400 ;
        RECT 149.100 91.950 154.050 94.050 ;
        RECT 125.400 90.000 136.050 90.450 ;
        RECT 125.400 89.400 135.450 90.000 ;
        RECT 125.400 87.450 126.450 89.400 ;
        RECT 50.400 86.400 126.450 87.450 ;
        RECT 127.950 87.450 130.050 88.050 ;
        RECT 136.950 87.450 139.050 91.050 ;
        RECT 157.950 90.450 160.050 94.050 ;
        RECT 172.950 91.950 177.900 94.050 ;
        RECT 179.100 91.950 184.050 94.050 ;
        RECT 173.400 90.450 174.450 91.950 ;
        RECT 157.950 90.000 174.450 90.450 ;
        RECT 158.400 89.400 174.450 90.000 ;
        RECT 193.950 88.950 196.050 94.050 ;
        RECT 199.950 93.450 202.050 94.050 ;
        RECT 208.950 93.450 211.050 94.050 ;
        RECT 199.950 92.400 211.050 93.450 ;
        RECT 199.950 91.950 202.050 92.400 ;
        RECT 208.950 91.950 211.050 92.400 ;
        RECT 217.950 91.950 220.050 95.400 ;
        RECT 223.950 94.950 226.050 95.400 ;
        RECT 229.950 94.950 235.050 97.050 ;
        RECT 238.800 96.000 240.900 97.050 ;
        RECT 241.950 96.000 244.200 97.050 ;
        RECT 238.800 94.950 241.050 96.000 ;
        RECT 242.100 94.950 244.200 96.000 ;
        RECT 259.950 94.950 264.900 97.050 ;
        RECT 266.100 96.450 268.200 97.050 ;
        RECT 274.950 96.450 277.050 97.050 ;
        RECT 266.100 95.400 277.050 96.450 ;
        RECT 266.100 94.950 268.200 95.400 ;
        RECT 274.950 94.950 277.050 95.400 ;
        RECT 223.950 93.450 226.050 94.050 ;
        RECT 229.950 93.450 232.050 94.050 ;
        RECT 223.950 92.400 232.050 93.450 ;
        RECT 223.950 91.950 226.050 92.400 ;
        RECT 229.950 91.950 232.050 92.400 ;
        RECT 238.950 91.950 241.050 94.950 ;
        RECT 244.950 93.450 250.050 94.050 ;
        RECT 256.950 93.450 259.050 94.050 ;
        RECT 244.950 92.400 259.050 93.450 ;
        RECT 244.950 91.950 250.050 92.400 ;
        RECT 256.950 91.950 259.050 92.400 ;
        RECT 262.950 93.450 265.050 94.050 ;
        RECT 268.950 93.450 271.050 94.050 ;
        RECT 262.950 92.400 271.050 93.450 ;
        RECT 262.950 91.950 265.050 92.400 ;
        RECT 268.950 91.950 271.050 92.400 ;
        RECT 280.950 93.450 283.050 94.050 ;
        RECT 280.950 92.400 288.450 93.450 ;
        RECT 280.950 91.950 283.050 92.400 ;
        RECT 220.950 88.950 226.050 91.050 ;
        RECT 250.950 90.450 253.050 91.050 ;
        RECT 287.400 90.450 288.450 92.400 ;
        RECT 289.950 91.950 292.050 97.050 ;
        RECT 295.950 91.950 298.050 97.050 ;
        RECT 320.400 96.000 333.450 96.450 ;
        RECT 320.400 95.400 334.050 96.000 ;
        RECT 316.950 93.450 319.050 94.050 ;
        RECT 320.400 93.450 321.450 95.400 ;
        RECT 308.400 92.400 321.450 93.450 ;
        RECT 292.950 90.450 295.050 91.050 ;
        RECT 250.950 89.400 295.050 90.450 ;
        RECT 250.950 88.950 253.050 89.400 ;
        RECT 292.950 88.950 295.050 89.400 ;
        RECT 301.950 90.450 304.050 91.050 ;
        RECT 308.400 90.450 309.450 92.400 ;
        RECT 316.950 91.950 319.050 92.400 ;
        RECT 322.950 91.950 328.050 94.050 ;
        RECT 331.950 91.950 334.050 95.400 ;
        RECT 334.950 94.950 337.050 98.400 ;
        RECT 355.950 98.400 373.050 99.450 ;
        RECT 355.950 97.950 358.050 98.400 ;
        RECT 367.950 97.950 373.050 98.400 ;
        RECT 340.950 94.950 346.050 97.050 ;
        RECT 352.950 94.050 355.050 97.050 ;
        RECT 358.800 96.000 360.900 97.050 ;
        RECT 364.950 96.450 367.050 97.050 ;
        RECT 370.950 96.450 373.050 97.200 ;
        RECT 358.800 94.950 361.050 96.000 ;
        RECT 364.950 95.400 373.050 96.450 ;
        RECT 364.950 94.950 367.050 95.400 ;
        RECT 370.950 95.100 373.050 95.400 ;
        RECT 385.950 96.450 388.050 97.050 ;
        RECT 394.950 96.450 397.050 97.050 ;
        RECT 385.950 95.400 397.050 96.450 ;
        RECT 385.950 94.950 388.050 95.400 ;
        RECT 394.950 94.950 397.050 95.400 ;
        RECT 400.950 94.950 403.050 100.050 ;
        RECT 436.950 99.450 439.050 100.050 ;
        RECT 481.950 99.450 484.050 100.050 ;
        RECT 490.950 99.450 493.050 100.050 ;
        RECT 416.400 99.000 447.450 99.450 ;
        RECT 415.950 98.400 447.450 99.000 ;
        RECT 406.950 97.050 409.050 97.200 ;
        RECT 406.950 95.100 412.050 97.050 ;
        RECT 408.000 94.950 412.050 95.100 ;
        RECT 415.950 94.950 418.050 98.400 ;
        RECT 436.950 97.950 439.050 98.400 ;
        RECT 358.950 94.050 361.050 94.950 ;
        RECT 301.950 89.400 309.450 90.450 ;
        RECT 316.950 90.450 322.050 91.050 ;
        RECT 337.950 90.450 340.050 94.050 ;
        RECT 352.950 93.000 357.900 94.050 ;
        RECT 353.400 92.400 357.900 93.000 ;
        RECT 354.000 91.950 357.900 92.400 ;
        RECT 358.800 93.000 361.050 94.050 ;
        RECT 362.100 93.450 364.200 94.050 ;
        RECT 372.000 93.900 376.050 94.050 ;
        RECT 370.950 93.450 376.050 93.900 ;
        RECT 358.800 91.950 360.900 93.000 ;
        RECT 362.100 92.400 376.050 93.450 ;
        RECT 362.100 91.950 364.200 92.400 ;
        RECT 370.950 91.950 376.050 92.400 ;
        RECT 388.950 91.950 394.050 94.050 ;
        RECT 370.950 91.800 373.050 91.950 ;
        RECT 397.950 91.050 400.050 94.050 ;
        RECT 406.950 93.450 409.050 93.900 ;
        RECT 412.950 93.450 415.050 94.050 ;
        RECT 406.950 92.400 415.050 93.450 ;
        RECT 406.950 91.800 409.050 92.400 ;
        RECT 412.950 91.950 415.050 92.400 ;
        RECT 316.950 90.000 340.050 90.450 ;
        RECT 361.950 90.450 364.050 91.050 ;
        RECT 397.800 90.450 400.050 91.050 ;
        RECT 361.950 90.000 400.050 90.450 ;
        RECT 401.100 90.450 403.200 91.050 ;
        RECT 418.950 90.450 421.050 94.050 ;
        RECT 427.950 93.450 430.050 94.050 ;
        RECT 436.950 93.450 439.050 94.050 ;
        RECT 427.950 92.400 439.050 93.450 ;
        RECT 427.950 91.950 430.050 92.400 ;
        RECT 436.950 91.950 439.050 92.400 ;
        RECT 442.950 91.950 445.050 97.050 ;
        RECT 446.400 96.450 447.450 98.400 ;
        RECT 481.950 98.400 493.050 99.450 ;
        RECT 481.950 97.950 484.050 98.400 ;
        RECT 490.950 97.950 493.050 98.400 ;
        RECT 499.950 99.450 502.050 100.050 ;
        RECT 520.950 99.450 523.050 100.050 ;
        RECT 499.950 98.400 523.050 99.450 ;
        RECT 499.950 97.950 502.050 98.400 ;
        RECT 520.950 97.950 523.050 98.400 ;
        RECT 454.800 96.450 456.900 97.050 ;
        RECT 446.400 95.400 456.900 96.450 ;
        RECT 454.800 94.950 456.900 95.400 ;
        RECT 458.100 94.950 463.050 97.050 ;
        RECT 520.950 94.950 526.050 97.050 ;
        RECT 532.950 94.950 535.050 100.050 ;
        RECT 538.950 96.450 541.050 97.050 ;
        RECT 544.950 96.450 547.050 97.050 ;
        RECT 538.950 95.400 547.050 96.450 ;
        RECT 538.950 94.950 541.050 95.400 ;
        RECT 544.950 94.950 547.050 95.400 ;
        RECT 550.950 94.950 553.050 100.050 ;
        RECT 559.950 99.450 562.050 100.050 ;
        RECT 592.950 99.450 595.050 100.050 ;
        RECT 607.950 99.450 610.050 100.050 ;
        RECT 559.950 99.000 588.450 99.450 ;
        RECT 559.950 98.400 589.050 99.000 ;
        RECT 559.950 97.950 562.050 98.400 ;
        RECT 554.400 96.000 573.450 96.450 ;
        RECT 553.950 95.400 574.050 96.000 ;
        RECT 448.950 91.950 454.050 94.050 ;
        RECT 401.100 90.000 421.050 90.450 ;
        RECT 316.950 89.400 339.450 90.000 ;
        RECT 361.950 89.400 399.900 90.000 ;
        RECT 301.950 88.950 304.050 89.400 ;
        RECT 316.950 88.950 322.050 89.400 ;
        RECT 361.950 88.950 364.050 89.400 ;
        RECT 397.800 88.950 399.900 89.400 ;
        RECT 401.100 89.400 420.450 90.000 ;
        RECT 401.100 88.950 403.200 89.400 ;
        RECT 436.950 88.950 441.900 91.050 ;
        RECT 443.100 90.450 445.200 91.050 ;
        RECT 457.950 90.450 460.050 94.050 ;
        RECT 469.950 93.450 472.050 94.050 ;
        RECT 478.800 93.450 480.900 94.050 ;
        RECT 469.950 92.400 480.900 93.450 ;
        RECT 482.100 93.000 484.200 94.050 ;
        RECT 469.950 91.950 472.050 92.400 ;
        RECT 478.800 91.950 480.900 92.400 ;
        RECT 481.950 91.950 484.200 93.000 ;
        RECT 511.950 91.950 516.900 94.050 ;
        RECT 518.100 93.450 520.200 94.050 ;
        RECT 529.950 93.450 532.050 94.050 ;
        RECT 518.100 92.400 532.050 93.450 ;
        RECT 518.100 91.950 520.200 92.400 ;
        RECT 529.950 91.950 532.050 92.400 ;
        RECT 443.100 90.000 460.050 90.450 ;
        RECT 460.950 90.450 463.050 91.050 ;
        RECT 475.950 90.450 478.050 91.050 ;
        RECT 443.100 89.400 459.450 90.000 ;
        RECT 460.950 89.400 478.050 90.450 ;
        RECT 443.100 88.950 445.200 89.400 ;
        RECT 460.950 88.950 463.050 89.400 ;
        RECT 475.950 88.950 478.050 89.400 ;
        RECT 481.950 88.950 484.050 91.950 ;
        RECT 535.950 91.050 538.050 94.050 ;
        RECT 544.950 91.950 550.050 94.050 ;
        RECT 553.950 91.950 556.050 95.400 ;
        RECT 571.950 91.950 574.050 95.400 ;
        RECT 586.950 94.950 589.050 98.400 ;
        RECT 592.950 98.400 610.050 99.450 ;
        RECT 611.400 99.450 612.450 101.400 ;
        RECT 646.950 101.400 673.050 102.450 ;
        RECT 646.950 101.100 649.050 101.400 ;
        RECT 670.950 100.950 673.050 101.400 ;
        RECT 688.950 102.450 691.050 103.050 ;
        RECT 742.950 102.450 745.050 103.050 ;
        RECT 688.950 101.400 745.050 102.450 ;
        RECT 688.950 100.950 691.050 101.400 ;
        RECT 742.950 100.950 745.050 101.400 ;
        RECT 769.950 102.450 772.050 103.050 ;
        RECT 832.950 102.450 835.050 103.050 ;
        RECT 769.950 101.400 835.050 102.450 ;
        RECT 769.950 100.950 772.050 101.400 ;
        RECT 832.950 100.950 835.050 101.400 ;
        RECT 628.950 99.450 631.050 100.050 ;
        RECT 611.400 98.400 631.050 99.450 ;
        RECT 592.950 97.950 595.050 98.400 ;
        RECT 607.950 97.950 610.050 98.400 ;
        RECT 628.950 97.950 631.050 98.400 ;
        RECT 640.800 99.000 642.900 100.050 ;
        RECT 644.100 99.900 648.000 100.050 ;
        RECT 640.800 97.950 643.050 99.000 ;
        RECT 644.100 97.950 649.050 99.900 ;
        RECT 661.800 99.450 663.900 100.050 ;
        RECT 595.950 94.950 601.050 97.050 ;
        RECT 604.950 94.050 607.050 97.050 ;
        RECT 610.950 96.450 613.050 97.050 ;
        RECT 616.950 96.450 619.050 97.050 ;
        RECT 610.950 95.400 619.050 96.450 ;
        RECT 610.950 94.950 613.050 95.400 ;
        RECT 616.950 94.950 619.050 95.400 ;
        RECT 622.950 94.950 628.050 97.050 ;
        RECT 589.950 91.950 595.050 94.050 ;
        RECT 604.950 93.000 610.050 94.050 ;
        RECT 605.400 92.400 610.050 93.000 ;
        RECT 606.000 91.950 610.050 92.400 ;
        RECT 631.950 91.950 634.050 97.050 ;
        RECT 640.950 94.950 643.050 97.950 ;
        RECT 646.950 97.800 649.050 97.950 ;
        RECT 650.400 98.400 663.900 99.450 ;
        RECT 665.100 99.450 667.200 100.050 ;
        RECT 676.950 99.450 679.050 100.050 ;
        RECT 665.100 99.000 679.050 99.450 ;
        RECT 650.400 97.050 651.450 98.400 ;
        RECT 661.800 97.950 663.900 98.400 ;
        RECT 664.950 98.400 679.050 99.000 ;
        RECT 664.950 97.950 667.200 98.400 ;
        RECT 676.950 97.950 679.050 98.400 ;
        RECT 664.950 97.050 667.050 97.950 ;
        RECT 646.950 95.400 651.450 97.050 ;
        RECT 646.950 94.950 651.000 95.400 ;
        RECT 658.950 94.950 663.900 97.050 ;
        RECT 664.950 96.000 667.200 97.050 ;
        RECT 679.950 96.450 682.050 97.050 ;
        RECT 665.100 94.950 667.200 96.000 ;
        RECT 674.400 95.400 682.050 96.450 ;
        RECT 659.400 93.450 660.450 94.950 ;
        RECT 674.400 93.450 675.450 95.400 ;
        RECT 679.950 94.950 682.050 95.400 ;
        RECT 694.950 94.950 700.050 97.050 ;
        RECT 703.950 94.950 709.050 97.050 ;
        RECT 742.950 96.450 745.050 100.050 ;
        RECT 778.950 99.450 781.050 100.050 ;
        RECT 761.400 98.400 781.050 99.450 ;
        RECT 761.400 97.050 762.450 98.400 ;
        RECT 778.950 97.950 781.050 98.400 ;
        RECT 808.950 99.450 811.050 100.050 ;
        RECT 814.950 99.450 819.900 100.050 ;
        RECT 808.950 98.400 819.900 99.450 ;
        RECT 808.950 97.950 811.050 98.400 ;
        RECT 814.950 97.950 819.900 98.400 ;
        RECT 821.100 99.450 823.200 100.050 ;
        RECT 853.950 99.450 856.050 100.050 ;
        RECT 821.100 98.400 856.050 99.450 ;
        RECT 821.100 97.950 823.200 98.400 ;
        RECT 853.950 97.950 856.050 98.400 ;
        RECT 751.950 96.450 756.900 97.050 ;
        RECT 742.950 96.000 756.900 96.450 ;
        RECT 743.400 95.400 756.900 96.000 ;
        RECT 751.950 94.950 756.900 95.400 ;
        RECT 758.100 94.950 763.050 97.050 ;
        RECT 790.950 96.450 793.050 97.200 ;
        RECT 796.950 96.450 799.050 97.050 ;
        RECT 764.400 95.400 799.050 96.450 ;
        RECT 659.400 92.400 675.450 93.450 ;
        RECT 502.950 90.450 505.050 91.050 ;
        RECT 508.950 90.450 511.050 91.050 ;
        RECT 502.950 89.400 511.050 90.450 ;
        RECT 502.950 88.950 505.050 89.400 ;
        RECT 508.950 88.950 511.050 89.400 ;
        RECT 535.800 90.000 538.050 91.050 ;
        RECT 539.100 90.450 541.200 91.050 ;
        RECT 547.950 90.450 550.050 91.050 ;
        RECT 535.800 88.950 537.900 90.000 ;
        RECT 539.100 89.400 550.050 90.450 ;
        RECT 539.100 88.950 541.200 89.400 ;
        RECT 547.950 88.950 550.050 89.400 ;
        RECT 559.950 90.450 562.050 91.050 ;
        RECT 568.950 90.450 571.050 91.050 ;
        RECT 559.950 89.400 571.050 90.450 ;
        RECT 559.950 88.950 562.050 89.400 ;
        RECT 568.950 88.950 571.050 89.400 ;
        RECT 577.950 90.450 580.050 91.050 ;
        RECT 616.950 90.450 619.050 91.050 ;
        RECT 646.950 90.450 649.050 91.050 ;
        RECT 577.950 89.400 649.050 90.450 ;
        RECT 577.950 88.950 580.050 89.400 ;
        RECT 616.950 88.950 619.050 89.400 ;
        RECT 646.950 88.950 649.050 89.400 ;
        RECT 676.950 88.950 679.050 94.050 ;
        RECT 682.950 93.450 685.050 94.050 ;
        RECT 695.400 93.450 696.450 94.950 ;
        RECT 764.400 94.050 765.450 95.400 ;
        RECT 790.950 95.100 793.050 95.400 ;
        RECT 796.950 94.950 799.050 95.400 ;
        RECT 802.950 94.950 808.050 97.050 ;
        RECT 812.400 96.000 834.450 96.450 ;
        RECT 812.400 95.400 835.050 96.000 ;
        RECT 682.950 92.400 696.450 93.450 ;
        RECT 682.950 91.950 685.050 92.400 ;
        RECT 697.950 91.950 703.050 94.050 ;
        RECT 706.950 90.450 709.050 94.050 ;
        RECT 712.950 93.450 715.050 94.050 ;
        RECT 721.800 93.450 723.900 94.050 ;
        RECT 712.950 92.400 723.900 93.450 ;
        RECT 712.950 91.950 715.050 92.400 ;
        RECT 721.800 91.950 723.900 92.400 ;
        RECT 725.100 93.450 727.200 94.050 ;
        RECT 736.950 93.450 739.050 94.050 ;
        RECT 725.100 92.400 739.050 93.450 ;
        RECT 725.100 91.950 727.200 92.400 ;
        RECT 736.950 91.950 739.050 92.400 ;
        RECT 742.950 93.450 745.050 94.050 ;
        RECT 748.950 93.450 751.050 94.050 ;
        RECT 742.950 92.400 751.050 93.450 ;
        RECT 742.950 91.950 745.050 92.400 ;
        RECT 748.950 91.950 751.050 92.400 ;
        RECT 718.950 90.450 723.900 91.050 ;
        RECT 706.950 90.000 723.900 90.450 ;
        RECT 725.100 90.450 727.200 91.050 ;
        RECT 754.950 90.450 757.050 94.050 ;
        RECT 760.950 92.400 765.450 94.050 ;
        RECT 760.950 91.950 765.000 92.400 ;
        RECT 766.950 91.950 772.050 94.050 ;
        RECT 775.950 91.950 781.050 94.050 ;
        RECT 784.950 91.050 787.050 94.050 ;
        RECT 792.000 93.900 796.050 94.050 ;
        RECT 790.950 91.950 796.050 93.900 ;
        RECT 799.950 93.450 802.050 94.050 ;
        RECT 812.400 93.450 813.450 95.400 ;
        RECT 799.950 92.400 813.450 93.450 ;
        RECT 820.950 93.450 823.050 94.050 ;
        RECT 820.950 93.000 831.450 93.450 ;
        RECT 820.950 92.400 832.050 93.000 ;
        RECT 799.950 91.950 802.050 92.400 ;
        RECT 820.950 91.950 823.050 92.400 ;
        RECT 790.950 91.800 793.050 91.950 ;
        RECT 772.950 90.450 775.050 91.050 ;
        RECT 725.100 90.000 757.050 90.450 ;
        RECT 707.400 89.400 723.900 90.000 ;
        RECT 718.950 88.950 723.900 89.400 ;
        RECT 724.950 89.400 756.450 90.000 ;
        RECT 758.400 89.400 775.050 90.450 ;
        RECT 724.950 88.950 727.200 89.400 ;
        RECT 127.950 87.000 139.050 87.450 ;
        RECT 145.950 87.450 148.050 88.050 ;
        RECT 178.950 87.450 181.050 88.050 ;
        RECT 127.950 86.400 138.450 87.000 ;
        RECT 145.950 86.400 181.050 87.450 ;
        RECT 28.950 85.950 31.050 86.400 ;
        RECT 46.950 85.950 49.050 86.400 ;
        RECT 94.950 85.950 97.050 86.400 ;
        RECT 127.950 85.950 130.050 86.400 ;
        RECT 145.950 85.950 148.050 86.400 ;
        RECT 178.950 85.950 181.050 86.400 ;
        RECT 325.950 87.450 328.050 88.050 ;
        RECT 358.950 87.450 361.050 88.050 ;
        RECT 325.950 86.400 361.050 87.450 ;
        RECT 325.950 85.950 328.050 86.400 ;
        RECT 358.950 85.950 361.050 86.400 ;
        RECT 397.950 87.450 400.050 88.050 ;
        RECT 406.950 87.450 409.050 88.050 ;
        RECT 397.950 86.400 409.050 87.450 ;
        RECT 397.950 85.950 400.050 86.400 ;
        RECT 406.950 85.950 409.050 86.400 ;
        RECT 535.950 87.450 538.050 88.050 ;
        RECT 550.950 87.450 553.050 88.050 ;
        RECT 535.950 86.400 553.050 87.450 ;
        RECT 535.950 85.950 538.050 86.400 ;
        RECT 550.950 85.950 553.050 86.400 ;
        RECT 691.950 87.450 694.050 88.050 ;
        RECT 724.950 87.450 727.050 88.950 ;
        RECT 691.950 87.000 727.050 87.450 ;
        RECT 727.950 87.450 730.050 88.050 ;
        RECT 758.400 87.450 759.450 89.400 ;
        RECT 772.950 88.950 775.050 89.400 ;
        RECT 781.800 90.000 783.900 91.050 ;
        RECT 784.950 90.000 787.200 91.050 ;
        RECT 781.800 88.950 784.050 90.000 ;
        RECT 785.100 88.950 787.200 90.000 ;
        RECT 829.950 88.950 832.050 92.400 ;
        RECT 832.950 91.950 835.050 95.400 ;
        RECT 847.950 93.450 850.050 94.050 ;
        RECT 839.400 92.400 850.050 93.450 ;
        RECT 839.400 91.050 840.450 92.400 ;
        RECT 847.950 91.950 850.050 92.400 ;
        RECT 835.950 89.400 840.450 91.050 ;
        RECT 835.950 88.950 840.000 89.400 ;
        RECT 781.950 88.050 784.050 88.950 ;
        RECT 691.950 86.400 726.600 87.000 ;
        RECT 727.950 86.400 759.450 87.450 ;
        RECT 781.800 87.000 784.050 88.050 ;
        RECT 785.100 87.450 787.200 88.050 ;
        RECT 835.950 87.450 838.050 88.050 ;
        RECT 691.950 85.950 694.050 86.400 ;
        RECT 727.950 85.950 730.050 86.400 ;
        RECT 781.800 85.950 783.900 87.000 ;
        RECT 785.100 86.400 838.050 87.450 ;
        RECT 785.100 85.950 787.200 86.400 ;
        RECT 835.950 85.950 838.050 86.400 ;
        RECT 40.950 84.450 43.050 85.050 ;
        RECT 52.950 84.450 55.050 85.050 ;
        RECT 40.950 83.400 55.050 84.450 ;
        RECT 40.950 82.950 43.050 83.400 ;
        RECT 52.950 82.950 55.050 83.400 ;
        RECT 82.950 84.450 85.050 85.050 ;
        RECT 124.950 84.450 127.050 85.050 ;
        RECT 82.950 83.400 127.050 84.450 ;
        RECT 82.950 82.950 85.050 83.400 ;
        RECT 124.950 82.950 127.050 83.400 ;
        RECT 157.950 84.450 160.050 85.050 ;
        RECT 208.950 84.450 211.050 85.050 ;
        RECT 157.950 83.400 211.050 84.450 ;
        RECT 157.950 82.950 160.050 83.400 ;
        RECT 208.950 82.950 211.050 83.400 ;
        RECT 247.950 84.450 250.050 85.050 ;
        RECT 355.950 84.450 358.050 85.050 ;
        RECT 247.950 83.400 358.050 84.450 ;
        RECT 247.950 82.950 250.050 83.400 ;
        RECT 355.950 82.950 358.050 83.400 ;
        RECT 391.950 84.450 394.050 85.050 ;
        RECT 424.950 84.450 427.050 85.050 ;
        RECT 487.950 84.450 490.050 85.050 ;
        RECT 391.950 83.400 490.050 84.450 ;
        RECT 391.950 82.950 394.050 83.400 ;
        RECT 424.950 82.950 427.050 83.400 ;
        RECT 487.950 82.950 490.050 83.400 ;
        RECT 514.950 84.450 517.050 85.050 ;
        RECT 601.950 84.450 604.050 85.050 ;
        RECT 514.950 83.400 604.050 84.450 ;
        RECT 514.950 82.950 517.050 83.400 ;
        RECT 601.950 82.950 604.050 83.400 ;
        RECT 754.950 84.450 757.050 85.050 ;
        RECT 785.400 84.450 786.450 85.950 ;
        RECT 754.950 83.400 786.450 84.450 ;
        RECT 805.950 84.450 808.050 85.050 ;
        RECT 850.950 84.450 853.050 85.050 ;
        RECT 805.950 83.400 853.050 84.450 ;
        RECT 754.950 82.950 757.050 83.400 ;
        RECT 805.950 82.950 808.050 83.400 ;
        RECT 850.950 82.950 853.050 83.400 ;
        RECT 91.950 81.450 94.050 82.050 ;
        RECT 163.950 81.450 166.050 82.050 ;
        RECT 91.950 80.400 166.050 81.450 ;
        RECT 91.950 79.950 94.050 80.400 ;
        RECT 163.950 79.950 166.050 80.400 ;
        RECT 169.950 81.450 172.050 82.050 ;
        RECT 220.950 81.450 223.050 82.050 ;
        RECT 307.950 81.450 310.050 82.050 ;
        RECT 169.950 80.400 210.450 81.450 ;
        RECT 169.950 79.950 172.050 80.400 ;
        RECT 25.950 78.450 28.050 79.050 ;
        RECT 184.950 78.450 187.050 79.050 ;
        RECT 25.950 77.400 187.050 78.450 ;
        RECT 209.400 78.450 210.450 80.400 ;
        RECT 220.950 80.400 310.050 81.450 ;
        RECT 220.950 79.950 223.050 80.400 ;
        RECT 307.950 79.950 310.050 80.400 ;
        RECT 358.950 81.450 361.050 82.050 ;
        RECT 427.950 81.450 430.050 82.050 ;
        RECT 358.950 80.400 430.050 81.450 ;
        RECT 358.950 79.950 361.050 80.400 ;
        RECT 427.950 79.950 430.050 80.400 ;
        RECT 721.950 81.450 724.050 82.050 ;
        RECT 793.950 81.450 796.050 82.050 ;
        RECT 721.950 80.400 796.050 81.450 ;
        RECT 721.950 79.950 724.050 80.400 ;
        RECT 793.950 79.950 796.050 80.400 ;
        RECT 385.950 78.450 388.050 79.050 ;
        RECT 209.400 77.400 388.050 78.450 ;
        RECT 25.950 76.950 28.050 77.400 ;
        RECT 184.950 76.950 187.050 77.400 ;
        RECT 385.950 76.950 388.050 77.400 ;
        RECT 451.950 78.450 454.050 79.050 ;
        RECT 466.950 78.450 469.050 79.050 ;
        RECT 451.950 77.400 469.050 78.450 ;
        RECT 451.950 76.950 454.050 77.400 ;
        RECT 466.950 76.950 469.050 77.400 ;
        RECT 670.950 78.450 673.050 79.050 ;
        RECT 682.950 78.450 685.050 79.050 ;
        RECT 670.950 77.400 685.050 78.450 ;
        RECT 670.950 76.950 673.050 77.400 ;
        RECT 682.950 76.950 685.050 77.400 ;
        RECT 736.950 78.450 739.050 79.050 ;
        RECT 802.950 78.450 805.050 79.050 ;
        RECT 736.950 77.400 805.050 78.450 ;
        RECT 736.950 76.950 739.050 77.400 ;
        RECT 802.950 76.950 805.050 77.400 ;
        RECT 118.950 75.450 121.050 76.050 ;
        RECT 193.950 75.450 196.050 76.050 ;
        RECT 118.950 74.400 196.050 75.450 ;
        RECT 118.950 73.950 121.050 74.400 ;
        RECT 193.950 73.950 196.050 74.400 ;
        RECT 274.950 75.450 277.050 76.050 ;
        RECT 463.800 75.450 465.900 76.050 ;
        RECT 274.950 74.400 465.900 75.450 ;
        RECT 274.950 73.950 277.050 74.400 ;
        RECT 463.800 73.950 465.900 74.400 ;
        RECT 467.100 75.450 469.200 76.050 ;
        RECT 484.950 75.450 487.050 76.050 ;
        RECT 467.100 74.400 487.050 75.450 ;
        RECT 467.100 73.950 469.200 74.400 ;
        RECT 484.950 73.950 487.050 74.400 ;
        RECT 688.950 75.450 691.050 76.050 ;
        RECT 748.950 75.450 751.050 76.050 ;
        RECT 760.950 75.450 763.050 76.050 ;
        RECT 688.950 74.400 763.050 75.450 ;
        RECT 688.950 73.950 691.050 74.400 ;
        RECT 748.950 73.950 751.050 74.400 ;
        RECT 760.950 73.950 763.050 74.400 ;
        RECT 772.950 75.450 775.050 76.050 ;
        RECT 781.950 75.450 784.050 76.050 ;
        RECT 829.950 75.450 832.050 76.050 ;
        RECT 772.950 74.400 832.050 75.450 ;
        RECT 772.950 73.950 775.050 74.400 ;
        RECT 781.950 73.950 784.050 74.400 ;
        RECT 829.950 73.950 832.050 74.400 ;
        RECT 133.950 72.450 136.050 73.050 ;
        RECT 178.950 72.450 181.050 73.050 ;
        RECT 325.950 72.450 328.050 73.050 ;
        RECT 133.950 71.400 328.050 72.450 ;
        RECT 133.950 70.950 136.050 71.400 ;
        RECT 178.950 70.950 181.050 71.400 ;
        RECT 325.950 70.950 328.050 71.400 ;
        RECT 430.950 72.450 433.050 73.050 ;
        RECT 568.950 72.450 571.050 73.050 ;
        RECT 430.950 71.400 571.050 72.450 ;
        RECT 430.950 70.950 433.050 71.400 ;
        RECT 568.950 70.950 571.050 71.400 ;
        RECT 700.950 72.450 703.050 73.050 ;
        RECT 784.950 72.450 787.050 73.050 ;
        RECT 700.950 71.400 787.050 72.450 ;
        RECT 700.950 70.950 703.050 71.400 ;
        RECT 784.950 70.950 787.050 71.400 ;
        RECT 94.950 69.450 97.050 70.050 ;
        RECT 100.950 69.450 103.050 70.050 ;
        RECT 94.950 68.400 103.050 69.450 ;
        RECT 94.950 67.950 97.050 68.400 ;
        RECT 100.950 67.950 103.050 68.400 ;
        RECT 175.950 69.450 178.050 70.050 ;
        RECT 187.950 69.450 190.050 70.050 ;
        RECT 175.950 68.400 190.050 69.450 ;
        RECT 175.950 67.950 178.050 68.400 ;
        RECT 187.950 67.950 190.050 68.400 ;
        RECT 196.950 69.450 199.050 70.050 ;
        RECT 226.950 69.450 229.050 70.050 ;
        RECT 340.950 69.450 343.050 70.050 ;
        RECT 196.950 68.400 343.050 69.450 ;
        RECT 196.950 67.950 199.050 68.400 ;
        RECT 226.950 67.950 229.050 68.400 ;
        RECT 340.950 67.950 343.050 68.400 ;
        RECT 409.950 69.450 412.050 70.050 ;
        RECT 460.800 69.450 462.900 70.050 ;
        RECT 409.950 68.400 462.900 69.450 ;
        RECT 409.950 67.950 412.050 68.400 ;
        RECT 460.800 67.950 462.900 68.400 ;
        RECT 464.100 69.450 466.200 70.050 ;
        RECT 544.950 69.450 547.050 70.050 ;
        RECT 464.100 68.400 547.050 69.450 ;
        RECT 464.100 67.950 466.200 68.400 ;
        RECT 544.950 67.950 547.050 68.400 ;
        RECT 562.950 69.450 565.050 70.050 ;
        RECT 583.950 69.450 586.050 70.050 ;
        RECT 562.950 68.400 586.050 69.450 ;
        RECT 562.950 67.950 565.050 68.400 ;
        RECT 583.950 67.950 586.050 68.400 ;
        RECT 670.950 69.450 673.050 70.050 ;
        RECT 697.950 69.450 700.050 70.050 ;
        RECT 670.950 68.400 700.050 69.450 ;
        RECT 670.950 67.950 673.050 68.400 ;
        RECT 697.950 67.950 700.050 68.400 ;
        RECT 706.950 69.450 709.050 70.050 ;
        RECT 721.950 69.450 724.050 70.050 ;
        RECT 820.950 69.450 823.050 70.050 ;
        RECT 706.950 68.400 724.050 69.450 ;
        RECT 706.950 67.950 709.050 68.400 ;
        RECT 721.950 67.950 724.050 68.400 ;
        RECT 740.400 68.400 823.050 69.450 ;
        RECT 740.400 67.050 741.450 68.400 ;
        RECT 820.950 67.950 823.050 68.400 ;
        RECT 31.950 66.450 34.050 67.050 ;
        RECT 109.800 66.450 111.900 67.050 ;
        RECT 31.950 65.400 111.900 66.450 ;
        RECT 31.950 64.950 34.050 65.400 ;
        RECT 109.800 64.950 111.900 65.400 ;
        RECT 113.100 66.450 115.200 67.050 ;
        RECT 217.950 66.450 220.050 67.050 ;
        RECT 113.100 65.400 220.050 66.450 ;
        RECT 113.100 64.950 115.200 65.400 ;
        RECT 217.950 64.950 220.050 65.400 ;
        RECT 295.950 66.450 298.050 67.050 ;
        RECT 304.950 66.450 307.050 67.050 ;
        RECT 295.950 65.400 307.050 66.450 ;
        RECT 295.950 64.950 298.050 65.400 ;
        RECT 304.950 64.950 307.050 65.400 ;
        RECT 316.950 66.450 319.050 67.050 ;
        RECT 328.950 66.450 331.050 67.050 ;
        RECT 316.950 65.400 331.050 66.450 ;
        RECT 316.950 64.950 319.050 65.400 ;
        RECT 328.950 64.950 331.050 65.400 ;
        RECT 37.950 63.450 40.050 64.050 ;
        RECT 103.950 63.450 106.050 64.050 ;
        RECT 37.950 62.400 106.050 63.450 ;
        RECT 37.950 61.950 40.050 62.400 ;
        RECT 103.950 61.950 106.050 62.400 ;
        RECT 124.950 63.450 127.050 64.050 ;
        RECT 316.950 63.450 319.050 64.050 ;
        RECT 334.950 63.450 337.050 67.050 ;
        RECT 625.950 66.450 628.050 67.050 ;
        RECT 664.950 66.450 667.050 67.050 ;
        RECT 625.950 65.400 667.050 66.450 ;
        RECT 124.950 62.400 174.450 63.450 ;
        RECT 124.950 61.950 127.050 62.400 ;
        RECT 173.400 61.050 174.450 62.400 ;
        RECT 316.950 63.000 337.050 63.450 ;
        RECT 349.950 63.450 352.050 64.050 ;
        RECT 364.800 63.450 366.900 64.050 ;
        RECT 316.950 62.400 336.450 63.000 ;
        RECT 349.950 62.400 366.900 63.450 ;
        RECT 316.950 61.950 319.050 62.400 ;
        RECT 349.950 61.950 352.050 62.400 ;
        RECT 364.800 61.950 366.900 62.400 ;
        RECT 368.100 63.450 370.200 64.050 ;
        RECT 403.950 63.450 406.050 64.050 ;
        RECT 368.100 62.400 406.050 63.450 ;
        RECT 460.950 63.300 463.050 65.400 ;
        RECT 625.950 64.950 628.050 65.400 ;
        RECT 664.950 64.950 667.050 65.400 ;
        RECT 682.950 66.450 685.050 67.050 ;
        RECT 694.950 66.450 697.050 67.050 ;
        RECT 739.950 66.450 742.050 67.050 ;
        RECT 682.950 65.400 742.050 66.450 ;
        RECT 682.950 64.950 685.050 65.400 ;
        RECT 694.950 64.950 697.050 65.400 ;
        RECT 739.950 64.950 742.050 65.400 ;
        RECT 745.950 66.450 748.050 67.050 ;
        RECT 811.950 66.450 814.050 67.050 ;
        RECT 745.950 65.400 814.050 66.450 ;
        RECT 745.950 64.950 748.050 65.400 ;
        RECT 811.950 64.950 814.050 65.400 ;
        RECT 368.100 61.950 370.200 62.400 ;
        RECT 403.950 61.950 406.050 62.400 ;
        RECT 17.400 60.000 27.450 60.450 ;
        RECT 16.950 59.400 27.450 60.000 ;
        RECT 16.950 55.950 19.050 59.400 ;
        RECT 26.400 58.050 27.450 59.400 ;
        RECT 25.950 57.450 30.000 58.050 ;
        RECT 43.950 57.450 46.050 58.050 ;
        RECT 25.950 57.000 30.300 57.450 ;
        RECT 43.950 57.000 54.450 57.450 ;
        RECT 25.950 55.950 31.050 57.000 ;
        RECT 43.950 56.400 55.050 57.000 ;
        RECT 43.950 55.950 46.050 56.400 ;
        RECT 28.950 55.050 31.050 55.950 ;
        RECT 13.950 49.950 16.050 55.050 ;
        RECT 19.950 51.450 22.050 55.050 ;
        RECT 28.800 54.000 31.050 55.050 ;
        RECT 28.800 52.950 30.900 54.000 ;
        RECT 32.100 52.950 37.050 55.050 ;
        RECT 31.950 51.450 34.050 52.050 ;
        RECT 37.950 51.450 40.050 52.050 ;
        RECT 19.950 51.000 40.050 51.450 ;
        RECT 20.400 50.400 40.050 51.000 ;
        RECT 31.950 49.950 34.050 50.400 ;
        RECT 37.950 49.950 40.050 50.400 ;
        RECT 46.950 49.950 49.050 55.050 ;
        RECT 52.950 52.950 55.050 56.400 ;
        RECT 70.950 55.950 76.050 58.050 ;
        RECT 79.950 55.950 82.050 61.050 ;
        RECT 163.950 60.450 166.050 61.050 ;
        RECT 169.800 60.450 171.900 61.050 ;
        RECT 155.400 59.400 171.900 60.450 ;
        RECT 88.950 57.450 91.050 58.050 ;
        RECT 112.950 57.450 115.050 58.050 ;
        RECT 88.950 56.400 115.050 57.450 ;
        RECT 88.950 55.950 91.050 56.400 ;
        RECT 112.950 55.950 115.050 56.400 ;
        RECT 118.950 57.450 121.050 58.050 ;
        RECT 136.950 57.450 139.050 58.050 ;
        RECT 118.950 56.400 139.050 57.450 ;
        RECT 58.950 52.950 64.050 55.050 ;
        RECT 52.950 49.950 58.050 52.050 ;
        RECT 76.950 51.450 79.050 55.050 ;
        RECT 82.950 54.450 88.050 55.050 ;
        RECT 97.800 54.450 99.900 55.050 ;
        RECT 82.950 53.400 99.900 54.450 ;
        RECT 82.950 52.950 88.050 53.400 ;
        RECT 97.800 52.950 99.900 53.400 ;
        RECT 101.100 52.950 106.050 55.050 ;
        RECT 118.950 54.450 121.050 56.400 ;
        RECT 136.950 55.950 139.050 56.400 ;
        RECT 145.950 57.450 148.050 58.050 ;
        RECT 155.400 57.450 156.450 59.400 ;
        RECT 163.950 58.950 166.050 59.400 ;
        RECT 169.800 58.950 171.900 59.400 ;
        RECT 173.100 60.450 175.200 61.050 ;
        RECT 187.950 60.450 190.050 61.050 ;
        RECT 220.950 60.450 223.050 61.050 ;
        RECT 173.100 59.400 190.050 60.450 ;
        RECT 209.400 60.000 223.050 60.450 ;
        RECT 173.100 58.950 175.200 59.400 ;
        RECT 187.950 58.950 190.050 59.400 ;
        RECT 208.950 59.400 223.050 60.000 ;
        RECT 145.950 56.400 156.450 57.450 ;
        RECT 145.950 55.950 148.050 56.400 ;
        RECT 107.250 54.000 121.050 54.450 ;
        RECT 106.950 53.400 121.050 54.000 ;
        RECT 106.950 52.050 109.050 53.400 ;
        RECT 118.950 52.950 121.050 53.400 ;
        RECT 124.950 52.950 130.050 55.050 ;
        RECT 88.950 51.450 91.050 52.050 ;
        RECT 76.950 51.000 91.050 51.450 ;
        RECT 77.400 50.400 91.050 51.000 ;
        RECT 88.950 49.950 91.050 50.400 ;
        RECT 94.800 51.000 96.900 52.050 ;
        RECT 94.800 49.950 97.050 51.000 ;
        RECT 98.100 49.950 103.050 52.050 ;
        RECT 106.800 51.000 109.050 52.050 ;
        RECT 110.100 51.450 112.200 52.050 ;
        RECT 121.950 51.450 124.050 52.050 ;
        RECT 106.800 49.950 108.900 51.000 ;
        RECT 110.100 50.400 124.050 51.450 ;
        RECT 110.100 49.950 112.200 50.400 ;
        RECT 121.950 49.950 124.050 50.400 ;
        RECT 127.950 51.450 130.050 52.050 ;
        RECT 133.950 51.450 136.050 52.050 ;
        RECT 127.950 50.400 136.050 51.450 ;
        RECT 142.950 51.450 145.050 55.050 ;
        RECT 148.950 52.950 154.050 55.050 ;
        RECT 157.950 54.450 160.050 58.050 ;
        RECT 155.400 53.400 160.050 54.450 ;
        RECT 155.400 51.450 156.450 53.400 ;
        RECT 157.950 52.950 160.050 53.400 ;
        RECT 163.950 52.950 166.050 58.050 ;
        RECT 193.950 57.450 198.000 58.050 ;
        RECT 193.950 55.950 198.450 57.450 ;
        RECT 199.950 55.950 205.050 58.050 ;
        RECT 208.950 55.950 211.050 59.400 ;
        RECT 220.950 58.950 223.050 59.400 ;
        RECT 244.950 60.450 247.050 61.050 ;
        RECT 244.950 60.000 264.450 60.450 ;
        RECT 244.950 59.400 265.050 60.000 ;
        RECT 244.950 58.950 247.050 59.400 ;
        RECT 262.950 55.950 265.050 59.400 ;
        RECT 268.950 55.950 274.050 58.050 ;
        RECT 277.950 57.450 283.050 58.050 ;
        RECT 277.950 56.400 300.450 57.450 ;
        RECT 277.950 55.950 283.050 56.400 ;
        RECT 178.950 52.950 184.050 55.050 ;
        RECT 187.950 52.950 193.050 55.050 ;
        RECT 197.400 54.450 198.450 55.950 ;
        RECT 299.400 55.050 300.450 56.400 ;
        RECT 304.950 55.950 307.050 61.050 ;
        RECT 334.950 60.450 337.050 61.050 ;
        RECT 359.100 60.450 361.200 61.050 ;
        RECT 436.950 60.450 439.050 61.050 ;
        RECT 334.950 59.400 361.200 60.450 ;
        RECT 334.950 58.950 337.050 59.400 ;
        RECT 358.950 58.950 361.200 59.400 ;
        RECT 419.400 59.400 439.050 60.450 ;
        RECT 461.850 59.700 463.050 63.300 ;
        RECT 481.950 62.400 484.050 64.500 ;
        RECT 700.950 63.450 703.050 64.050 ;
        RECT 650.250 62.400 703.050 63.450 ;
        RECT 358.950 58.050 361.050 58.950 ;
        RECT 419.400 58.050 420.450 59.400 ;
        RECT 436.950 58.950 439.050 59.400 ;
        RECT 316.950 57.450 319.050 58.050 ;
        RECT 322.950 57.450 325.050 58.050 ;
        RECT 316.950 56.400 325.050 57.450 ;
        RECT 316.950 55.950 319.050 56.400 ;
        RECT 322.950 55.950 325.050 56.400 ;
        RECT 328.950 57.450 331.050 58.050 ;
        RECT 355.800 57.450 357.900 58.050 ;
        RECT 328.950 57.000 357.900 57.450 ;
        RECT 358.950 57.000 361.200 58.050 ;
        RECT 328.950 56.400 358.050 57.000 ;
        RECT 328.950 55.950 331.050 56.400 ;
        RECT 355.800 55.950 358.050 56.400 ;
        RECT 359.100 55.950 361.200 57.000 ;
        RECT 373.950 55.950 379.050 58.050 ;
        RECT 382.950 57.450 388.050 58.050 ;
        RECT 397.950 57.450 400.050 58.050 ;
        RECT 382.950 56.400 400.050 57.450 ;
        RECT 382.950 55.950 388.050 56.400 ;
        RECT 397.950 55.950 400.050 56.400 ;
        RECT 403.950 55.950 409.050 58.050 ;
        RECT 418.950 57.450 423.000 58.050 ;
        RECT 430.950 57.450 433.050 58.050 ;
        RECT 460.950 57.600 463.050 59.700 ;
        RECT 418.950 57.000 423.450 57.450 ;
        RECT 430.950 57.000 447.600 57.450 ;
        RECT 418.950 55.950 424.050 57.000 ;
        RECT 430.950 56.400 448.050 57.000 ;
        RECT 430.950 55.950 433.050 56.400 ;
        RECT 205.950 54.450 208.050 55.050 ;
        RECT 197.400 53.400 208.050 54.450 ;
        RECT 205.950 52.950 208.050 53.400 ;
        RECT 142.950 51.000 156.450 51.450 ;
        RECT 143.400 50.400 156.450 51.000 ;
        RECT 160.950 51.450 163.050 52.050 ;
        RECT 175.950 51.450 178.050 52.050 ;
        RECT 160.950 50.400 178.050 51.450 ;
        RECT 127.950 49.950 130.050 50.400 ;
        RECT 133.950 49.950 136.050 50.400 ;
        RECT 160.950 49.950 163.050 50.400 ;
        RECT 175.950 49.950 178.050 50.400 ;
        RECT 181.950 49.950 187.050 52.050 ;
        RECT 190.950 51.450 193.050 52.050 ;
        RECT 196.950 51.450 199.050 52.050 ;
        RECT 190.950 50.400 199.050 51.450 ;
        RECT 190.950 49.950 193.050 50.400 ;
        RECT 196.950 49.950 199.050 50.400 ;
        RECT 211.950 49.950 214.050 55.050 ;
        RECT 226.950 52.950 231.900 55.050 ;
        RECT 233.100 54.000 235.200 55.050 ;
        RECT 232.950 52.950 235.200 54.000 ;
        RECT 247.950 52.950 253.050 55.050 ;
        RECT 265.950 54.450 268.050 55.050 ;
        RECT 274.950 54.450 277.050 55.050 ;
        RECT 265.950 53.400 277.050 54.450 ;
        RECT 265.950 52.950 268.050 53.400 ;
        RECT 274.950 52.950 277.050 53.400 ;
        RECT 220.950 51.450 223.050 52.050 ;
        RECT 229.950 51.450 232.050 52.050 ;
        RECT 220.950 50.400 232.050 51.450 ;
        RECT 232.950 51.450 235.050 52.950 ;
        RECT 241.950 51.450 244.050 52.050 ;
        RECT 232.950 51.000 244.050 51.450 ;
        RECT 220.950 49.950 223.050 50.400 ;
        RECT 229.950 49.950 232.050 50.400 ;
        RECT 233.400 50.400 244.050 51.000 ;
        RECT 94.950 49.050 97.050 49.950 ;
        RECT 13.950 48.450 16.050 49.050 ;
        RECT 31.950 48.450 34.050 49.050 ;
        RECT 13.950 47.400 34.050 48.450 ;
        RECT 13.950 46.950 16.050 47.400 ;
        RECT 31.950 46.950 34.050 47.400 ;
        RECT 79.950 48.450 82.050 49.050 ;
        RECT 94.800 48.450 97.050 49.050 ;
        RECT 79.950 48.000 97.050 48.450 ;
        RECT 148.950 48.450 151.050 49.050 ;
        RECT 160.950 48.450 163.050 49.050 ;
        RECT 79.950 47.400 96.900 48.000 ;
        RECT 79.950 46.950 82.050 47.400 ;
        RECT 94.800 46.950 96.900 47.400 ;
        RECT 148.950 47.400 163.050 48.450 ;
        RECT 148.950 46.950 151.050 47.400 ;
        RECT 160.950 46.950 163.050 47.400 ;
        RECT 211.950 48.450 214.050 49.050 ;
        RECT 233.400 48.450 234.450 50.400 ;
        RECT 241.950 49.950 244.050 50.400 ;
        RECT 211.950 47.400 234.450 48.450 ;
        RECT 211.950 46.950 214.050 47.400 ;
        RECT 253.950 46.950 256.050 52.050 ;
        RECT 271.950 51.450 274.050 52.050 ;
        RECT 280.950 51.450 283.050 55.050 ;
        RECT 286.950 54.450 289.050 55.050 ;
        RECT 292.950 54.450 295.050 55.050 ;
        RECT 286.950 53.400 295.050 54.450 ;
        RECT 299.400 53.400 304.050 55.050 ;
        RECT 286.950 52.950 289.050 53.400 ;
        RECT 292.950 52.950 295.050 53.400 ;
        RECT 300.000 52.950 304.050 53.400 ;
        RECT 271.950 51.000 283.050 51.450 ;
        RECT 271.950 50.400 282.450 51.000 ;
        RECT 271.950 49.950 274.050 50.400 ;
        RECT 283.950 49.950 286.050 52.050 ;
        RECT 293.400 51.450 294.450 52.950 ;
        RECT 307.950 51.450 310.050 55.050 ;
        RECT 293.400 51.000 310.050 51.450 ;
        RECT 313.950 51.450 316.050 52.050 ;
        RECT 325.950 51.450 328.050 55.050 ;
        RECT 355.950 52.950 358.050 55.950 ;
        RECT 361.950 52.950 367.050 55.050 ;
        RECT 373.950 54.450 376.050 55.050 ;
        RECT 382.950 54.450 385.050 55.050 ;
        RECT 373.950 53.400 385.050 54.450 ;
        RECT 373.950 52.950 376.050 53.400 ;
        RECT 382.950 52.950 385.050 53.400 ;
        RECT 388.950 52.950 394.050 55.050 ;
        RECT 400.950 54.450 403.050 55.050 ;
        RECT 409.800 54.450 411.900 55.050 ;
        RECT 400.950 53.400 411.900 54.450 ;
        RECT 400.950 52.950 403.050 53.400 ;
        RECT 409.800 52.950 411.900 53.400 ;
        RECT 413.100 52.950 418.050 55.050 ;
        RECT 421.950 52.950 424.050 55.950 ;
        RECT 445.950 55.050 448.050 56.400 ;
        RECT 436.950 52.950 441.900 55.050 ;
        RECT 442.800 54.000 444.900 55.050 ;
        RECT 445.950 54.000 448.200 55.050 ;
        RECT 442.800 52.950 445.050 54.000 ;
        RECT 446.100 52.950 448.200 54.000 ;
        RECT 313.950 51.000 328.050 51.450 ;
        RECT 383.400 51.450 384.450 52.950 ;
        RECT 442.950 52.050 445.050 52.950 ;
        RECT 406.950 51.450 409.050 52.050 ;
        RECT 293.400 50.400 309.450 51.000 ;
        RECT 313.950 50.400 327.450 51.000 ;
        RECT 383.400 50.400 409.050 51.450 ;
        RECT 313.950 49.950 316.050 50.400 ;
        RECT 406.950 49.950 409.050 50.400 ;
        RECT 418.950 49.950 424.050 52.050 ;
        RECT 284.400 48.450 285.450 49.950 ;
        RECT 304.950 48.450 307.050 49.050 ;
        RECT 284.400 47.400 307.050 48.450 ;
        RECT 43.950 45.450 46.050 46.050 ;
        RECT 67.950 45.450 70.050 46.050 ;
        RECT 43.950 44.400 70.050 45.450 ;
        RECT 43.950 43.950 46.050 44.400 ;
        RECT 67.950 43.950 70.050 44.400 ;
        RECT 118.950 45.450 121.050 46.050 ;
        RECT 284.400 45.450 285.450 47.400 ;
        RECT 304.950 46.950 307.050 47.400 ;
        RECT 118.950 44.400 285.450 45.450 ;
        RECT 286.950 45.450 289.050 46.050 ;
        RECT 310.950 45.450 313.050 46.050 ;
        RECT 346.950 45.450 349.050 49.050 ;
        RECT 403.950 48.450 406.050 49.050 ;
        RECT 436.950 48.450 439.050 52.050 ;
        RECT 442.800 51.000 445.050 52.050 ;
        RECT 442.800 49.950 444.900 51.000 ;
        RECT 448.950 49.950 453.900 52.050 ;
        RECT 455.100 49.950 460.050 52.050 ;
        RECT 457.950 48.450 460.050 49.050 ;
        RECT 403.950 48.000 439.050 48.450 ;
        RECT 403.950 47.400 438.450 48.000 ;
        RECT 452.400 47.400 460.050 48.450 ;
        RECT 403.950 46.950 406.050 47.400 ;
        RECT 452.400 45.450 453.450 47.400 ;
        RECT 457.950 46.950 460.050 47.400 ;
        RECT 461.850 45.600 463.050 57.600 ;
        RECT 466.950 49.950 471.900 52.050 ;
        RECT 473.100 49.950 478.050 52.050 ;
        RECT 482.100 45.600 483.300 62.400 ;
        RECT 511.950 60.450 514.050 61.050 ;
        RECT 517.950 60.450 520.050 61.050 ;
        RECT 631.950 60.450 634.050 61.050 ;
        RECT 511.950 59.400 520.050 60.450 ;
        RECT 581.400 60.000 634.050 60.450 ;
        RECT 511.950 58.950 514.050 59.400 ;
        RECT 517.950 58.950 520.050 59.400 ;
        RECT 580.950 59.400 634.050 60.000 ;
        RECT 502.950 54.450 505.050 55.050 ;
        RECT 502.950 53.400 510.450 54.450 ;
        RECT 502.950 52.950 505.050 53.400 ;
        RECT 509.400 52.050 510.450 53.400 ;
        RECT 511.950 52.950 517.050 55.050 ;
        RECT 520.950 52.950 523.050 58.050 ;
        RECT 568.950 55.950 574.050 58.050 ;
        RECT 580.950 55.950 583.050 59.400 ;
        RECT 601.950 57.450 604.050 58.050 ;
        RECT 625.950 57.450 628.050 58.050 ;
        RECT 601.950 56.400 628.050 57.450 ;
        RECT 574.950 52.950 580.050 55.050 ;
        RECT 601.950 52.950 604.050 56.400 ;
        RECT 625.950 55.950 628.050 56.400 ;
        RECT 631.950 55.950 634.050 59.400 ;
        RECT 650.250 58.050 651.300 62.400 ;
        RECT 700.950 61.950 703.050 62.400 ;
        RECT 712.950 63.450 715.050 64.050 ;
        RECT 754.950 63.450 757.050 64.050 ;
        RECT 712.950 62.400 757.050 63.450 ;
        RECT 712.950 61.950 715.050 62.400 ;
        RECT 754.950 61.950 757.050 62.400 ;
        RECT 763.950 63.450 766.050 64.050 ;
        RECT 802.950 63.450 805.050 64.050 ;
        RECT 763.950 62.400 805.050 63.450 ;
        RECT 763.950 61.950 766.050 62.400 ;
        RECT 802.950 61.950 805.050 62.400 ;
        RECT 823.950 63.450 826.050 64.050 ;
        RECT 844.950 63.450 847.050 64.050 ;
        RECT 823.950 62.400 847.050 63.450 ;
        RECT 823.950 61.950 826.050 62.400 ;
        RECT 844.950 61.950 847.050 62.400 ;
        RECT 688.800 60.000 690.900 61.050 ;
        RECT 688.800 58.950 691.050 60.000 ;
        RECT 688.950 58.050 691.050 58.950 ;
        RECT 637.950 57.450 640.050 58.050 ;
        RECT 646.800 57.450 648.900 58.050 ;
        RECT 637.950 56.400 648.900 57.450 ;
        RECT 637.950 55.950 640.050 56.400 ;
        RECT 646.800 55.950 648.900 56.400 ;
        RECT 649.800 55.950 651.900 58.050 ;
        RECT 653.100 55.950 658.050 58.050 ;
        RECT 664.950 57.450 667.050 58.050 ;
        RECT 670.950 57.450 673.050 58.050 ;
        RECT 664.950 56.400 673.050 57.450 ;
        RECT 664.950 55.950 667.050 56.400 ;
        RECT 670.950 55.950 673.050 56.400 ;
        RECT 676.950 57.450 679.050 58.050 ;
        RECT 682.950 57.450 685.050 58.050 ;
        RECT 676.950 56.400 685.050 57.450 ;
        RECT 676.950 55.950 679.050 56.400 ;
        RECT 682.950 55.950 685.050 56.400 ;
        RECT 688.800 57.000 691.050 58.050 ;
        RECT 688.800 55.950 690.900 57.000 ;
        RECT 692.100 55.950 697.050 58.050 ;
        RECT 712.950 55.950 715.050 61.050 ;
        RECT 736.950 60.450 739.050 61.050 ;
        RECT 742.950 60.450 745.050 61.050 ;
        RECT 736.950 59.400 745.050 60.450 ;
        RECT 736.950 58.950 739.050 59.400 ;
        RECT 742.950 58.950 745.050 59.400 ;
        RECT 748.950 55.950 751.050 61.050 ;
        RECT 754.950 55.950 760.050 58.050 ;
        RECT 772.950 55.950 775.050 61.050 ;
        RECT 796.950 60.450 799.050 61.050 ;
        RECT 850.950 60.450 853.050 61.050 ;
        RECT 796.950 59.400 853.050 60.450 ;
        RECT 796.950 58.950 799.050 59.400 ;
        RECT 850.950 58.950 853.050 59.400 ;
        RECT 781.950 55.950 787.050 58.050 ;
        RECT 793.950 57.450 796.050 58.050 ;
        RECT 808.950 57.450 811.050 58.050 ;
        RECT 793.950 56.400 811.050 57.450 ;
        RECT 793.950 55.950 796.050 56.400 ;
        RECT 619.950 54.450 622.050 55.050 ;
        RECT 634.950 54.450 637.050 55.050 ;
        RECT 619.950 53.400 637.050 54.450 ;
        RECT 619.950 52.950 622.050 53.400 ;
        RECT 634.950 52.950 637.050 53.400 ;
        RECT 640.950 54.450 643.050 55.050 ;
        RECT 650.400 54.450 651.450 55.950 ;
        RECT 640.950 53.400 651.450 54.450 ;
        RECT 640.950 52.950 643.050 53.400 ;
        RECT 509.400 50.400 514.050 52.050 ;
        RECT 510.000 49.950 514.050 50.400 ;
        RECT 484.950 48.450 487.050 49.050 ;
        RECT 493.950 48.450 496.050 49.050 ;
        RECT 484.950 47.400 496.050 48.450 ;
        RECT 484.950 46.950 487.050 47.400 ;
        RECT 493.950 46.950 496.050 47.400 ;
        RECT 517.950 46.950 520.050 52.050 ;
        RECT 523.950 49.950 529.050 52.050 ;
        RECT 535.950 49.950 541.050 52.050 ;
        RECT 562.950 46.950 565.050 52.050 ;
        RECT 592.950 51.450 595.050 52.050 ;
        RECT 598.950 51.450 601.050 52.050 ;
        RECT 592.950 50.400 601.050 51.450 ;
        RECT 592.950 49.950 595.050 50.400 ;
        RECT 598.950 49.950 601.050 50.400 ;
        RECT 604.950 48.450 607.050 52.050 ;
        RECT 625.950 51.450 628.050 52.050 ;
        RECT 652.950 51.450 655.050 55.050 ;
        RECT 655.950 54.450 658.050 55.950 ;
        RECT 670.800 54.450 672.900 55.050 ;
        RECT 655.950 54.000 672.900 54.450 ;
        RECT 674.100 54.000 676.200 55.050 ;
        RECT 656.400 53.400 672.900 54.000 ;
        RECT 670.800 52.950 672.900 53.400 ;
        RECT 673.950 52.950 676.200 54.000 ;
        RECT 679.950 54.450 682.050 55.050 ;
        RECT 691.950 54.450 694.050 55.050 ;
        RECT 679.950 53.400 694.050 54.450 ;
        RECT 679.950 52.950 682.050 53.400 ;
        RECT 691.950 52.950 694.050 53.400 ;
        RECT 703.950 54.450 706.050 55.050 ;
        RECT 709.950 54.450 712.050 55.050 ;
        RECT 703.950 53.400 712.050 54.450 ;
        RECT 703.950 52.950 706.050 53.400 ;
        RECT 709.950 52.950 712.050 53.400 ;
        RECT 625.950 51.000 655.050 51.450 ;
        RECT 664.950 51.450 667.050 52.050 ;
        RECT 673.950 51.450 676.050 52.950 ;
        RECT 664.950 51.000 676.050 51.450 ;
        RECT 715.950 51.450 718.050 55.050 ;
        RECT 721.950 52.950 727.050 55.050 ;
        RECT 730.950 54.450 733.050 55.050 ;
        RECT 739.950 54.450 742.050 55.050 ;
        RECT 730.950 53.400 742.050 54.450 ;
        RECT 730.950 52.950 733.050 53.400 ;
        RECT 739.950 52.950 742.050 53.400 ;
        RECT 724.950 51.450 730.050 52.050 ;
        RECT 715.950 51.000 730.050 51.450 ;
        RECT 751.950 51.450 754.050 55.050 ;
        RECT 769.950 52.950 774.900 55.050 ;
        RECT 775.800 54.000 777.900 55.050 ;
        RECT 779.100 54.450 781.200 55.050 ;
        RECT 790.800 54.450 792.900 55.050 ;
        RECT 775.800 52.950 778.050 54.000 ;
        RECT 779.100 53.400 792.900 54.450 ;
        RECT 779.100 52.950 781.200 53.400 ;
        RECT 790.800 52.950 792.900 53.400 ;
        RECT 794.100 52.950 799.050 55.050 ;
        RECT 808.950 52.950 811.050 56.400 ;
        RECT 814.950 52.950 817.050 58.050 ;
        RECT 829.950 52.950 832.050 58.050 ;
        RECT 837.000 57.450 841.050 58.050 ;
        RECT 836.400 57.000 841.050 57.450 ;
        RECT 835.950 55.950 841.050 57.000 ;
        RECT 835.950 52.950 838.050 55.950 ;
        RECT 844.950 54.450 850.050 55.050 ;
        RECT 839.400 54.000 850.050 54.450 ;
        RECT 838.950 53.400 850.050 54.000 ;
        RECT 769.950 51.450 772.050 52.950 ;
        RECT 751.950 51.000 772.050 51.450 ;
        RECT 775.950 51.450 778.050 52.950 ;
        RECT 794.400 51.450 795.450 52.950 ;
        RECT 811.950 51.450 814.050 52.050 ;
        RECT 775.950 51.000 795.450 51.450 ;
        RECT 625.950 50.400 654.450 51.000 ;
        RECT 664.950 50.400 675.600 51.000 ;
        RECT 716.400 50.400 730.050 51.000 ;
        RECT 752.400 50.400 771.450 51.000 ;
        RECT 776.250 50.400 795.450 51.000 ;
        RECT 797.400 50.400 814.050 51.450 ;
        RECT 625.950 49.950 628.050 50.400 ;
        RECT 664.950 49.950 667.050 50.400 ;
        RECT 724.950 49.950 730.050 50.400 ;
        RECT 613.950 48.450 616.050 49.050 ;
        RECT 604.950 47.400 616.050 48.450 ;
        RECT 604.950 46.950 607.050 47.400 ;
        RECT 613.950 46.950 616.050 47.400 ;
        RECT 751.950 48.450 754.050 49.050 ;
        RECT 757.950 48.450 760.050 49.050 ;
        RECT 751.950 47.400 760.050 48.450 ;
        RECT 751.950 46.950 754.050 47.400 ;
        RECT 757.950 46.950 760.050 47.400 ;
        RECT 763.950 48.450 766.050 49.050 ;
        RECT 797.400 48.450 798.450 50.400 ;
        RECT 811.950 49.950 814.050 50.400 ;
        RECT 817.950 51.450 820.050 52.050 ;
        RECT 823.950 51.450 826.050 52.050 ;
        RECT 832.950 51.450 835.050 52.050 ;
        RECT 817.950 50.400 826.050 51.450 ;
        RECT 817.950 49.950 820.050 50.400 ;
        RECT 823.950 49.950 826.050 50.400 ;
        RECT 827.400 50.400 835.050 51.450 ;
        RECT 763.950 47.400 798.450 48.450 ;
        RECT 802.950 48.450 805.050 49.050 ;
        RECT 808.950 48.450 811.050 49.050 ;
        RECT 802.950 47.400 811.050 48.450 ;
        RECT 763.950 46.950 766.050 47.400 ;
        RECT 802.950 46.950 805.050 47.400 ;
        RECT 808.950 46.950 811.050 47.400 ;
        RECT 814.950 48.450 817.050 49.050 ;
        RECT 827.400 48.450 828.450 50.400 ;
        RECT 832.950 49.950 835.050 50.400 ;
        RECT 838.950 49.950 841.050 53.400 ;
        RECT 844.950 52.950 850.050 53.400 ;
        RECT 814.950 47.400 828.450 48.450 ;
        RECT 814.950 46.950 817.050 47.400 ;
        RECT 850.950 46.950 856.050 49.050 ;
        RECT 286.950 44.400 453.450 45.450 ;
        RECT 118.950 43.950 121.050 44.400 ;
        RECT 286.950 43.950 289.050 44.400 ;
        RECT 310.950 43.950 313.050 44.400 ;
        RECT 460.950 43.500 463.050 45.600 ;
        RECT 481.950 43.500 484.050 45.600 ;
        RECT 691.950 45.450 694.050 46.050 ;
        RECT 700.950 45.450 703.050 46.050 ;
        RECT 691.950 44.400 703.050 45.450 ;
        RECT 691.950 43.950 694.050 44.400 ;
        RECT 700.950 43.950 703.050 44.400 ;
        RECT 739.950 45.450 742.050 46.050 ;
        RECT 817.950 45.450 820.050 46.050 ;
        RECT 838.950 45.450 841.050 46.200 ;
        RECT 739.950 44.400 841.050 45.450 ;
        RECT 739.950 43.950 742.050 44.400 ;
        RECT 817.950 43.950 820.050 44.400 ;
        RECT 838.950 44.100 841.050 44.400 ;
        RECT 4.950 42.450 7.050 43.050 ;
        RECT 25.950 42.450 28.050 43.050 ;
        RECT 58.950 42.450 61.050 43.050 ;
        RECT 91.950 42.450 94.050 43.050 ;
        RECT 4.950 41.400 94.050 42.450 ;
        RECT 4.950 40.950 7.050 41.400 ;
        RECT 25.950 40.950 28.050 41.400 ;
        RECT 58.950 40.950 61.050 41.400 ;
        RECT 91.950 40.950 94.050 41.400 ;
        RECT 103.950 42.450 106.050 43.050 ;
        RECT 199.950 42.450 202.050 43.050 ;
        RECT 313.800 42.450 315.900 43.050 ;
        RECT 103.950 41.400 202.050 42.450 ;
        RECT 103.950 40.950 106.050 41.400 ;
        RECT 199.950 40.950 202.050 41.400 ;
        RECT 254.400 41.400 315.900 42.450 ;
        RECT 254.400 40.050 255.450 41.400 ;
        RECT 313.800 40.950 315.900 41.400 ;
        RECT 317.100 42.450 319.200 43.050 ;
        RECT 385.950 42.450 388.050 43.050 ;
        RECT 317.100 41.400 388.050 42.450 ;
        RECT 317.100 40.950 319.200 41.400 ;
        RECT 385.950 40.950 388.050 41.400 ;
        RECT 421.950 42.450 424.050 43.050 ;
        RECT 454.950 42.450 457.050 43.050 ;
        RECT 421.950 41.400 457.050 42.450 ;
        RECT 421.950 40.950 424.050 41.400 ;
        RECT 454.950 40.950 457.050 41.400 ;
        RECT 682.950 42.450 685.050 43.050 ;
        RECT 724.950 42.450 727.050 43.050 ;
        RECT 760.950 42.450 763.050 43.050 ;
        RECT 682.950 41.400 763.050 42.450 ;
        RECT 682.950 40.950 685.050 41.400 ;
        RECT 724.950 40.950 727.050 41.400 ;
        RECT 760.950 40.950 763.050 41.400 ;
        RECT 766.950 42.450 769.050 43.050 ;
        RECT 838.950 42.450 841.050 42.900 ;
        RECT 766.950 41.400 841.050 42.450 ;
        RECT 766.950 40.950 769.050 41.400 ;
        RECT 838.950 40.800 841.050 41.400 ;
        RECT 76.950 39.450 79.050 40.050 ;
        RECT 253.950 39.450 256.050 40.050 ;
        RECT 76.950 38.400 256.050 39.450 ;
        RECT 76.950 37.950 79.050 38.400 ;
        RECT 253.950 37.950 256.050 38.400 ;
        RECT 322.950 39.450 325.050 40.050 ;
        RECT 370.950 39.450 373.050 40.050 ;
        RECT 322.950 38.400 373.050 39.450 ;
        RECT 322.950 37.950 325.050 38.400 ;
        RECT 370.950 37.950 373.050 38.400 ;
        RECT 442.950 39.450 445.050 40.050 ;
        RECT 475.950 39.450 478.050 40.050 ;
        RECT 442.950 38.400 478.050 39.450 ;
        RECT 442.950 37.950 445.050 38.400 ;
        RECT 475.950 37.950 478.050 38.400 ;
        RECT 664.950 39.450 667.050 40.050 ;
        RECT 718.950 39.450 721.050 40.050 ;
        RECT 763.950 39.450 766.050 40.050 ;
        RECT 664.950 38.400 766.050 39.450 ;
        RECT 664.950 37.950 667.050 38.400 ;
        RECT 718.950 37.950 721.050 38.400 ;
        RECT 763.950 37.950 766.050 38.400 ;
        RECT 775.950 39.450 778.050 40.050 ;
        RECT 856.950 39.450 859.050 40.050 ;
        RECT 775.950 38.400 859.050 39.450 ;
        RECT 775.950 37.950 778.050 38.400 ;
        RECT 856.950 37.950 859.050 38.400 ;
        RECT 127.950 36.450 130.050 37.050 ;
        RECT 136.950 36.450 139.050 37.050 ;
        RECT 127.950 35.400 139.050 36.450 ;
        RECT 127.950 34.950 130.050 35.400 ;
        RECT 136.950 34.950 139.050 35.400 ;
        RECT 277.950 36.450 280.050 37.050 ;
        RECT 295.950 36.450 298.050 37.050 ;
        RECT 334.950 36.450 337.050 37.050 ;
        RECT 277.950 35.400 337.050 36.450 ;
        RECT 277.950 34.950 280.050 35.400 ;
        RECT 295.950 34.950 298.050 35.400 ;
        RECT 334.950 34.950 337.050 35.400 ;
        RECT 340.950 36.450 343.050 37.050 ;
        RECT 469.950 36.450 472.050 37.050 ;
        RECT 340.950 35.400 472.050 36.450 ;
        RECT 340.950 34.950 343.050 35.400 ;
        RECT 469.950 34.950 472.050 35.400 ;
        RECT 697.950 36.450 700.050 37.050 ;
        RECT 790.950 36.450 793.050 37.050 ;
        RECT 697.950 35.400 793.050 36.450 ;
        RECT 697.950 34.950 700.050 35.400 ;
        RECT 790.950 34.950 793.050 35.400 ;
        RECT 808.950 36.450 811.050 37.050 ;
        RECT 817.950 36.450 820.050 37.050 ;
        RECT 808.950 35.400 820.050 36.450 ;
        RECT 808.950 34.950 811.050 35.400 ;
        RECT 817.950 34.950 820.050 35.400 ;
        RECT 172.950 33.450 175.050 34.050 ;
        RECT 181.950 33.450 184.050 34.050 ;
        RECT 172.950 32.400 184.050 33.450 ;
        RECT 172.950 31.950 175.050 32.400 ;
        RECT 181.950 31.950 184.050 32.400 ;
        RECT 214.950 33.450 217.050 34.050 ;
        RECT 247.950 33.450 250.050 34.050 ;
        RECT 358.950 33.450 361.050 34.050 ;
        RECT 415.950 33.450 418.050 34.050 ;
        RECT 214.950 32.400 333.450 33.450 ;
        RECT 214.950 31.950 217.050 32.400 ;
        RECT 247.950 31.950 250.050 32.400 ;
        RECT 332.400 31.050 333.450 32.400 ;
        RECT 358.950 32.400 418.050 33.450 ;
        RECT 358.950 31.950 361.050 32.400 ;
        RECT 415.950 31.950 418.050 32.400 ;
        RECT 802.950 31.950 808.050 34.050 ;
        RECT 832.950 33.450 835.050 34.050 ;
        RECT 809.400 32.400 835.050 33.450 ;
        RECT 46.950 30.450 49.050 31.050 ;
        RECT 76.950 30.450 79.050 31.050 ;
        RECT 14.400 30.000 79.050 30.450 ;
        RECT 13.950 29.400 79.050 30.000 ;
        RECT 13.950 25.950 16.050 29.400 ;
        RECT 46.950 28.950 49.050 29.400 ;
        RECT 76.950 28.950 79.050 29.400 ;
        RECT 211.950 30.450 214.050 31.050 ;
        RECT 217.950 30.450 220.050 31.050 ;
        RECT 220.950 30.450 223.050 31.050 ;
        RECT 211.950 29.400 223.050 30.450 ;
        RECT 211.950 28.950 214.050 29.400 ;
        RECT 19.950 27.450 22.050 28.050 ;
        RECT 43.950 27.450 46.050 28.050 ;
        RECT 19.950 26.400 46.050 27.450 ;
        RECT 19.950 25.950 22.050 26.400 ;
        RECT 43.950 25.950 46.050 26.400 ;
        RECT 49.950 22.950 52.050 28.050 ;
        RECT 97.950 27.450 100.050 28.050 ;
        RECT 65.400 27.000 100.050 27.450 ;
        RECT 64.950 26.400 100.050 27.000 ;
        RECT 55.950 24.450 58.050 25.050 ;
        RECT 64.950 24.450 67.050 26.400 ;
        RECT 97.950 25.950 100.050 26.400 ;
        RECT 106.950 27.450 109.050 28.050 ;
        RECT 148.950 27.450 151.050 28.050 ;
        RECT 160.950 27.450 163.050 28.050 ;
        RECT 181.950 27.450 184.050 28.050 ;
        RECT 199.950 27.450 202.050 28.050 ;
        RECT 106.950 26.400 163.050 27.450 ;
        RECT 106.950 25.950 109.050 26.400 ;
        RECT 148.950 25.950 151.050 26.400 ;
        RECT 160.950 25.950 163.050 26.400 ;
        RECT 173.400 26.400 184.050 27.450 ;
        RECT 188.400 27.000 202.050 27.450 ;
        RECT 55.950 23.400 67.050 24.450 ;
        RECT 55.950 22.950 58.050 23.400 ;
        RECT 64.950 22.950 67.050 23.400 ;
        RECT 70.950 24.450 73.050 25.050 ;
        RECT 82.950 24.450 85.050 25.050 ;
        RECT 70.950 23.400 85.050 24.450 ;
        RECT 70.950 22.950 73.050 23.400 ;
        RECT 82.950 22.950 85.050 23.400 ;
        RECT 13.950 21.450 16.050 22.050 ;
        RECT 19.950 21.450 24.900 22.050 ;
        RECT 13.950 20.400 24.900 21.450 ;
        RECT 13.950 19.950 16.050 20.400 ;
        RECT 19.950 19.950 24.900 20.400 ;
        RECT 26.100 19.950 31.050 22.050 ;
        RECT 43.950 19.950 49.050 22.050 ;
        RECT 25.950 15.450 28.050 19.050 ;
        RECT 52.950 18.450 55.050 22.050 ;
        RECT 64.950 19.950 70.050 22.050 ;
        RECT 73.950 21.450 79.050 22.050 ;
        RECT 85.950 21.450 88.050 22.050 ;
        RECT 73.950 20.400 88.050 21.450 ;
        RECT 73.950 19.950 79.050 20.400 ;
        RECT 85.950 19.950 88.050 20.400 ;
        RECT 91.950 19.950 97.050 22.050 ;
        RECT 106.950 19.950 109.050 25.050 ;
        RECT 112.950 19.950 115.050 25.050 ;
        RECT 130.950 24.450 133.050 25.050 ;
        RECT 173.400 24.450 174.450 26.400 ;
        RECT 181.950 25.950 184.050 26.400 ;
        RECT 187.950 26.400 202.050 27.000 ;
        RECT 187.950 24.450 190.050 26.400 ;
        RECT 199.950 25.950 202.050 26.400 ;
        RECT 217.950 25.950 220.050 29.400 ;
        RECT 220.950 28.950 223.050 29.400 ;
        RECT 229.950 30.450 232.050 31.050 ;
        RECT 292.800 30.450 294.900 31.050 ;
        RECT 229.950 29.400 294.900 30.450 ;
        RECT 296.100 30.000 298.200 31.050 ;
        RECT 229.950 28.950 232.050 29.400 ;
        RECT 130.950 23.400 174.450 24.450 ;
        RECT 176.550 24.000 190.050 24.450 ;
        RECT 175.950 23.400 190.050 24.000 ;
        RECT 130.950 22.950 133.050 23.400 ;
        RECT 124.950 19.950 130.050 22.050 ;
        RECT 133.950 19.950 139.050 22.050 ;
        RECT 143.400 21.450 144.450 23.400 ;
        RECT 172.800 22.050 174.900 22.200 ;
        RECT 148.950 21.450 151.050 22.050 ;
        RECT 143.400 20.400 151.050 21.450 ;
        RECT 148.950 19.950 151.050 20.400 ;
        RECT 166.950 20.100 174.900 22.050 ;
        RECT 175.950 22.050 178.050 23.400 ;
        RECT 187.950 22.950 190.050 23.400 ;
        RECT 196.950 24.600 199.050 25.200 ;
        RECT 208.950 25.050 211.050 25.200 ;
        RECT 205.950 24.600 211.050 25.050 ;
        RECT 196.950 23.550 211.050 24.600 ;
        RECT 196.950 23.100 199.050 23.550 ;
        RECT 205.950 23.100 211.050 23.550 ;
        RECT 205.950 22.950 210.000 23.100 ;
        RECT 235.950 22.950 241.050 25.050 ;
        RECT 244.950 22.950 247.050 28.050 ;
        RECT 259.950 25.950 262.050 29.400 ;
        RECT 292.800 28.950 294.900 29.400 ;
        RECT 295.950 28.950 298.200 30.000 ;
        RECT 301.950 30.450 304.050 31.050 ;
        RECT 322.950 30.450 325.050 31.050 ;
        RECT 301.950 29.400 325.050 30.450 ;
        RECT 301.950 28.950 304.050 29.400 ;
        RECT 322.950 28.950 325.050 29.400 ;
        RECT 331.950 30.450 334.050 31.050 ;
        RECT 373.950 30.450 376.050 31.050 ;
        RECT 331.950 29.400 376.050 30.450 ;
        RECT 436.950 29.400 439.050 31.500 ;
        RECT 457.950 29.400 460.050 31.500 ;
        RECT 508.950 30.450 511.050 31.050 ;
        RECT 742.950 30.450 745.050 31.050 ;
        RECT 508.950 29.400 745.050 30.450 ;
        RECT 751.950 29.400 754.050 31.500 ;
        RECT 772.950 29.400 775.050 31.500 ;
        RECT 796.950 30.450 799.050 31.050 ;
        RECT 809.400 30.450 810.450 32.400 ;
        RECT 832.950 31.950 835.050 32.400 ;
        RECT 796.950 29.400 810.450 30.450 ;
        RECT 811.950 30.450 814.050 31.050 ;
        RECT 823.950 30.450 826.050 31.050 ;
        RECT 811.950 29.400 826.050 30.450 ;
        RECT 331.950 28.950 334.050 29.400 ;
        RECT 373.950 28.950 376.050 29.400 ;
        RECT 268.950 27.450 271.050 28.050 ;
        RECT 268.950 27.000 282.450 27.450 ;
        RECT 268.950 26.400 283.050 27.000 ;
        RECT 268.950 25.950 271.050 26.400 ;
        RECT 280.950 22.950 283.050 26.400 ;
        RECT 295.950 25.950 298.050 28.950 ;
        RECT 286.950 24.450 289.050 25.050 ;
        RECT 301.950 24.450 304.050 25.050 ;
        RECT 286.950 23.400 304.050 24.450 ;
        RECT 286.950 22.950 289.050 23.400 ;
        RECT 301.950 22.950 304.050 23.400 ;
        RECT 310.950 22.950 313.050 28.050 ;
        RECT 316.950 22.950 319.050 28.050 ;
        RECT 357.000 27.450 361.050 28.050 ;
        RECT 356.400 27.000 361.050 27.450 ;
        RECT 355.950 25.950 361.050 27.000 ;
        RECT 397.950 27.450 400.050 28.050 ;
        RECT 421.950 27.450 424.050 28.050 ;
        RECT 397.950 26.400 424.050 27.450 ;
        RECT 397.950 25.950 400.050 26.400 ;
        RECT 355.950 22.950 358.050 25.950 ;
        RECT 403.950 25.050 406.050 26.400 ;
        RECT 421.950 25.950 424.050 26.400 ;
        RECT 427.950 25.950 433.050 28.050 ;
        RECT 361.950 24.450 364.050 25.050 ;
        RECT 367.950 24.450 370.050 25.050 ;
        RECT 361.950 23.400 370.050 24.450 ;
        RECT 361.950 22.950 364.050 23.400 ;
        RECT 367.950 22.950 370.050 23.400 ;
        RECT 403.800 24.000 406.050 25.050 ;
        RECT 403.800 22.950 405.900 24.000 ;
        RECT 175.950 21.000 178.200 22.050 ;
        RECT 166.950 19.950 174.000 20.100 ;
        RECT 176.100 19.950 178.200 21.000 ;
        RECT 181.950 19.950 187.050 22.050 ;
        RECT 190.950 21.450 193.050 22.050 ;
        RECT 196.950 21.450 199.050 22.050 ;
        RECT 190.950 20.400 199.050 21.450 ;
        RECT 190.950 19.950 193.050 20.400 ;
        RECT 196.950 19.950 199.050 20.400 ;
        RECT 214.950 19.950 220.050 22.050 ;
        RECT 65.400 18.450 66.450 19.950 ;
        RECT 52.950 18.000 66.450 18.450 ;
        RECT 53.400 17.400 66.450 18.000 ;
        RECT 73.950 18.450 76.050 19.050 ;
        RECT 88.950 18.450 91.050 19.050 ;
        RECT 73.950 17.400 91.050 18.450 ;
        RECT 73.950 16.950 76.050 17.400 ;
        RECT 88.950 16.950 91.050 17.400 ;
        RECT 97.950 18.450 100.050 19.050 ;
        RECT 109.950 18.450 112.050 19.050 ;
        RECT 97.950 17.400 112.050 18.450 ;
        RECT 97.950 16.950 100.050 17.400 ;
        RECT 109.950 16.950 112.050 17.400 ;
        RECT 118.950 16.950 124.050 19.050 ;
        RECT 130.950 16.950 136.050 19.050 ;
        RECT 172.950 16.950 178.050 19.050 ;
        RECT 193.950 18.450 196.050 19.050 ;
        RECT 211.950 18.450 214.050 19.050 ;
        RECT 241.950 18.450 244.050 22.050 ;
        RECT 247.950 19.950 253.050 22.050 ;
        RECT 265.950 19.950 271.050 22.050 ;
        RECT 277.950 19.950 282.900 22.050 ;
        RECT 284.100 19.950 289.050 22.050 ;
        RECT 301.950 21.450 304.050 22.050 ;
        RECT 313.950 21.450 316.050 22.050 ;
        RECT 301.950 20.400 316.050 21.450 ;
        RECT 301.950 19.950 304.050 20.400 ;
        RECT 313.950 19.950 316.050 20.400 ;
        RECT 319.950 19.950 325.050 22.050 ;
        RECT 334.950 21.450 337.050 22.050 ;
        RECT 349.800 21.450 351.900 22.050 ;
        RECT 334.950 20.400 351.900 21.450 ;
        RECT 334.950 19.950 337.050 20.400 ;
        RECT 349.800 19.950 351.900 20.400 ;
        RECT 352.800 21.000 354.900 22.050 ;
        RECT 352.800 19.950 355.050 21.000 ;
        RECT 356.100 19.950 361.050 22.050 ;
        RECT 376.950 21.450 379.050 22.050 ;
        RECT 362.400 20.400 379.050 21.450 ;
        RECT 193.950 18.000 244.050 18.450 ;
        RECT 193.950 17.400 243.450 18.000 ;
        RECT 193.950 16.950 196.050 17.400 ;
        RECT 211.950 16.950 214.050 17.400 ;
        RECT 331.950 16.950 336.900 19.050 ;
        RECT 338.100 16.950 343.050 19.050 ;
        RECT 352.950 18.450 355.050 19.950 ;
        RECT 362.400 18.450 363.450 20.400 ;
        RECT 376.950 19.950 379.050 20.400 ;
        RECT 394.950 21.450 397.050 22.050 ;
        RECT 403.950 21.450 406.050 22.050 ;
        RECT 394.950 20.400 406.050 21.450 ;
        RECT 394.950 19.950 397.050 20.400 ;
        RECT 403.950 19.950 406.050 20.400 ;
        RECT 352.950 18.000 363.450 18.450 ;
        RECT 353.250 17.400 363.450 18.000 ;
        RECT 367.950 18.450 370.050 19.050 ;
        RECT 373.950 18.450 376.050 19.050 ;
        RECT 367.950 17.400 376.050 18.450 ;
        RECT 367.950 16.950 370.050 17.400 ;
        RECT 373.950 16.950 376.050 17.400 ;
        RECT 382.950 18.450 385.050 19.050 ;
        RECT 424.950 18.450 427.050 22.050 ;
        RECT 382.950 18.000 427.050 18.450 ;
        RECT 382.950 17.400 426.450 18.000 ;
        RECT 382.950 16.950 385.050 17.400 ;
        RECT 74.400 15.450 75.450 16.950 ;
        RECT 25.950 15.000 75.450 15.450 ;
        RECT 26.400 14.400 75.450 15.000 ;
        RECT 166.950 15.450 169.050 16.050 ;
        RECT 181.950 15.450 184.050 16.050 ;
        RECT 166.950 14.400 184.050 15.450 ;
        RECT 166.950 13.950 169.050 14.400 ;
        RECT 181.950 13.950 184.050 14.400 ;
        RECT 196.950 15.450 199.050 16.050 ;
        RECT 268.950 15.450 271.050 16.050 ;
        RECT 196.950 14.400 271.050 15.450 ;
        RECT 196.950 13.950 199.050 14.400 ;
        RECT 268.950 13.950 271.050 14.400 ;
        RECT 49.950 12.450 52.050 13.050 ;
        RECT 112.950 12.450 115.050 13.050 ;
        RECT 49.950 11.400 115.050 12.450 ;
        RECT 49.950 10.950 52.050 11.400 ;
        RECT 112.950 10.950 115.050 11.400 ;
        RECT 142.950 12.450 145.050 13.050 ;
        RECT 271.950 12.450 274.050 13.050 ;
        RECT 437.700 12.600 438.900 29.400 ;
        RECT 442.950 19.950 445.050 25.050 ;
        RECT 448.950 19.950 451.050 25.050 ;
        RECT 457.950 17.400 459.150 29.400 ;
        RECT 508.950 28.950 511.050 29.400 ;
        RECT 742.950 28.950 745.050 29.400 ;
        RECT 461.400 27.000 486.450 27.450 ;
        RECT 460.950 26.400 486.450 27.000 ;
        RECT 460.950 22.950 463.050 26.400 ;
        RECT 485.400 25.050 486.450 26.400 ;
        RECT 481.950 22.950 487.050 25.050 ;
        RECT 499.950 22.950 502.050 28.050 ;
        RECT 652.950 27.450 655.050 28.050 ;
        RECT 593.550 27.000 655.050 27.450 ;
        RECT 592.950 26.400 655.050 27.000 ;
        RECT 592.950 25.050 595.050 26.400 ;
        RECT 652.950 25.950 655.050 26.400 ;
        RECT 658.950 27.450 661.050 28.050 ;
        RECT 691.950 27.450 694.050 28.050 ;
        RECT 658.950 26.400 694.050 27.450 ;
        RECT 658.950 25.950 661.050 26.400 ;
        RECT 691.950 25.950 694.050 26.400 ;
        RECT 703.950 27.450 706.050 28.050 ;
        RECT 715.950 27.450 718.050 28.050 ;
        RECT 739.950 27.450 742.050 28.050 ;
        RECT 703.950 26.400 742.050 27.450 ;
        RECT 703.950 25.950 706.050 26.400 ;
        RECT 715.950 25.950 718.050 26.400 ;
        RECT 739.950 25.950 742.050 26.400 ;
        RECT 586.950 24.450 591.900 25.050 ;
        RECT 551.400 23.400 591.900 24.450 ;
        RECT 592.950 24.000 595.200 25.050 ;
        RECT 505.950 19.950 511.050 22.050 ;
        RECT 520.950 21.450 523.050 22.050 ;
        RECT 529.950 21.450 532.050 22.050 ;
        RECT 520.950 20.400 532.050 21.450 ;
        RECT 520.950 19.950 523.050 20.400 ;
        RECT 529.950 19.950 532.050 20.400 ;
        RECT 538.950 21.450 541.050 22.050 ;
        RECT 547.950 21.450 550.050 22.050 ;
        RECT 538.950 20.400 550.050 21.450 ;
        RECT 538.950 19.950 541.050 20.400 ;
        RECT 547.950 19.950 550.050 20.400 ;
        RECT 551.400 19.050 552.450 23.400 ;
        RECT 586.950 22.950 591.900 23.400 ;
        RECT 593.100 22.950 595.200 24.000 ;
        RECT 613.950 22.950 619.050 25.050 ;
        RECT 565.800 21.000 567.900 22.050 ;
        RECT 568.800 21.000 570.900 22.050 ;
        RECT 572.100 21.450 574.200 22.050 ;
        RECT 580.950 21.450 586.050 22.050 ;
        RECT 565.800 19.950 568.050 21.000 ;
        RECT 568.800 19.950 571.050 21.000 ;
        RECT 572.100 20.400 586.050 21.450 ;
        RECT 572.100 19.950 574.200 20.400 ;
        RECT 580.950 19.950 586.050 20.400 ;
        RECT 589.950 19.950 595.050 22.050 ;
        RECT 565.950 19.050 568.050 19.950 ;
        RECT 457.950 15.300 460.050 17.400 ;
        RECT 142.950 11.400 274.050 12.450 ;
        RECT 142.950 10.950 145.050 11.400 ;
        RECT 271.950 10.950 274.050 11.400 ;
        RECT 436.950 10.500 439.050 12.600 ;
        RECT 457.950 11.700 459.150 15.300 ;
        RECT 526.950 13.950 529.050 19.050 ;
        RECT 532.950 15.450 535.050 19.050 ;
        RECT 541.950 16.950 547.050 19.050 ;
        RECT 550.950 16.950 553.050 19.050 ;
        RECT 559.950 18.450 562.050 19.050 ;
        RECT 554.400 17.400 562.050 18.450 ;
        RECT 554.400 15.450 555.450 17.400 ;
        RECT 559.950 16.950 562.050 17.400 ;
        RECT 565.800 18.000 568.050 19.050 ;
        RECT 568.950 19.050 571.050 19.950 ;
        RECT 568.950 18.000 571.200 19.050 ;
        RECT 565.800 16.950 567.900 18.000 ;
        RECT 569.100 16.950 571.200 18.000 ;
        RECT 625.950 16.950 628.050 22.050 ;
        RECT 631.950 19.950 634.050 25.050 ;
        RECT 637.950 24.450 640.050 25.050 ;
        RECT 685.950 24.450 688.050 25.050 ;
        RECT 637.950 24.000 645.450 24.450 ;
        RECT 637.950 23.400 646.050 24.000 ;
        RECT 637.950 22.950 640.050 23.400 ;
        RECT 643.950 19.950 646.050 23.400 ;
        RECT 685.950 23.400 696.450 24.450 ;
        RECT 685.950 22.950 688.050 23.400 ;
        RECT 695.400 22.050 696.450 23.400 ;
        RECT 652.950 21.450 655.050 22.050 ;
        RECT 661.950 21.450 664.050 22.050 ;
        RECT 652.950 20.400 664.050 21.450 ;
        RECT 652.950 19.950 655.050 20.400 ;
        RECT 661.950 19.950 664.050 20.400 ;
        RECT 679.950 19.950 684.900 22.050 ;
        RECT 685.800 21.000 687.900 22.050 ;
        RECT 685.800 19.950 688.050 21.000 ;
        RECT 689.100 19.950 694.050 22.050 ;
        RECT 695.400 20.400 700.050 22.050 ;
        RECT 696.000 19.950 700.050 20.400 ;
        RECT 718.950 19.950 721.050 25.050 ;
        RECT 742.950 24.450 745.050 25.050 ;
        RECT 748.950 24.450 751.050 25.050 ;
        RECT 742.950 23.400 751.050 24.450 ;
        RECT 742.950 22.950 745.050 23.400 ;
        RECT 748.950 22.950 751.050 23.400 ;
        RECT 724.950 19.950 730.050 22.050 ;
        RECT 736.950 19.950 742.050 22.050 ;
        RECT 631.950 18.450 634.050 19.050 ;
        RECT 640.950 18.450 643.050 19.050 ;
        RECT 631.950 17.400 643.050 18.450 ;
        RECT 631.950 16.950 634.050 17.400 ;
        RECT 640.950 16.050 643.050 17.400 ;
        RECT 532.950 15.000 555.450 15.450 ;
        RECT 533.400 14.400 555.450 15.000 ;
        RECT 565.950 15.450 568.050 16.050 ;
        RECT 637.800 15.450 639.900 16.050 ;
        RECT 565.950 14.400 639.900 15.450 ;
        RECT 640.950 15.000 643.200 16.050 ;
        RECT 565.950 13.950 568.050 14.400 ;
        RECT 637.800 13.950 639.900 14.400 ;
        RECT 641.100 13.950 643.200 15.000 ;
        RECT 646.950 15.450 649.050 19.050 ;
        RECT 655.950 16.950 661.050 19.050 ;
        RECT 664.950 18.450 667.050 19.050 ;
        RECT 680.400 18.450 681.450 19.950 ;
        RECT 664.950 17.400 681.450 18.450 ;
        RECT 664.950 16.950 667.050 17.400 ;
        RECT 685.950 16.950 688.050 19.950 ;
        RECT 715.950 18.450 718.050 19.050 ;
        RECT 721.950 18.450 724.050 19.050 ;
        RECT 715.950 17.400 724.050 18.450 ;
        RECT 715.950 16.950 718.050 17.400 ;
        RECT 721.950 16.950 724.050 17.400 ;
        RECT 730.950 16.950 736.050 19.050 ;
        RECT 673.950 15.450 676.050 16.050 ;
        RECT 646.950 14.400 676.050 15.450 ;
        RECT 739.950 15.450 742.050 19.050 ;
        RECT 752.850 17.400 754.050 29.400 ;
        RECT 757.950 22.950 763.050 25.050 ;
        RECT 766.950 19.950 769.050 25.050 ;
        RECT 745.950 15.450 748.050 16.050 ;
        RECT 739.950 15.000 748.050 15.450 ;
        RECT 751.950 15.300 754.050 17.400 ;
        RECT 740.400 14.400 748.050 15.000 ;
        RECT 646.950 13.950 649.050 14.400 ;
        RECT 673.950 13.950 676.050 14.400 ;
        RECT 745.950 13.950 748.050 14.400 ;
        RECT 526.950 12.450 529.050 13.050 ;
        RECT 538.950 12.450 541.050 13.050 ;
        RECT 82.950 9.450 85.050 10.050 ;
        RECT 136.950 9.450 139.050 10.050 ;
        RECT 82.950 8.400 139.050 9.450 ;
        RECT 82.950 7.950 85.050 8.400 ;
        RECT 136.950 7.950 139.050 8.400 ;
        RECT 172.950 9.450 175.050 10.050 ;
        RECT 196.950 9.450 199.050 10.050 ;
        RECT 172.950 8.400 199.050 9.450 ;
        RECT 172.950 7.950 175.050 8.400 ;
        RECT 196.950 7.950 199.050 8.400 ;
        RECT 205.950 9.450 208.050 10.050 ;
        RECT 238.950 9.450 241.050 10.050 ;
        RECT 457.950 9.600 460.050 11.700 ;
        RECT 526.950 11.400 541.050 12.450 ;
        RECT 526.950 10.950 529.050 11.400 ;
        RECT 538.950 10.950 541.050 11.400 ;
        RECT 544.950 12.450 547.050 13.200 ;
        RECT 616.950 12.450 619.050 13.050 ;
        RECT 544.950 11.400 619.050 12.450 ;
        RECT 544.950 11.100 547.050 11.400 ;
        RECT 616.950 10.950 619.050 11.400 ;
        RECT 640.950 12.450 643.050 13.050 ;
        RECT 709.950 12.450 712.050 13.050 ;
        RECT 640.950 11.400 712.050 12.450 ;
        RECT 752.850 11.700 754.050 15.300 ;
        RECT 773.100 12.600 774.300 29.400 ;
        RECT 796.950 28.950 799.050 29.400 ;
        RECT 811.950 28.950 814.050 29.400 ;
        RECT 823.950 28.950 826.050 29.400 ;
        RECT 838.950 30.450 841.050 31.050 ;
        RECT 838.950 29.400 846.450 30.450 ;
        RECT 838.950 28.950 841.050 29.400 ;
        RECT 845.400 28.050 846.450 29.400 ;
        RECT 790.950 22.950 793.050 28.050 ;
        RECT 802.950 27.450 805.050 28.050 ;
        RECT 802.950 26.400 813.450 27.450 ;
        RECT 845.400 26.400 850.050 28.050 ;
        RECT 802.950 25.950 805.050 26.400 ;
        RECT 812.400 25.050 813.450 26.400 ;
        RECT 846.000 25.950 850.050 26.400 ;
        RECT 796.950 24.450 799.050 25.050 ;
        RECT 808.950 24.450 811.050 25.050 ;
        RECT 796.950 23.400 811.050 24.450 ;
        RECT 812.400 23.400 817.050 25.050 ;
        RECT 796.950 22.950 799.050 23.400 ;
        RECT 808.950 22.950 811.050 23.400 ;
        RECT 813.000 22.950 817.050 23.400 ;
        RECT 826.950 24.450 829.050 25.050 ;
        RECT 835.950 24.450 838.050 25.050 ;
        RECT 826.950 23.400 838.050 24.450 ;
        RECT 826.950 22.950 829.050 23.400 ;
        RECT 835.950 22.950 838.050 23.400 ;
        RECT 775.950 21.450 778.050 22.050 ;
        RECT 787.950 21.450 790.050 22.050 ;
        RECT 775.950 20.400 790.050 21.450 ;
        RECT 775.950 19.950 778.050 20.400 ;
        RECT 787.950 19.950 790.050 20.400 ;
        RECT 793.950 16.950 796.050 22.050 ;
        RECT 799.950 21.450 802.050 22.050 ;
        RECT 811.950 21.450 814.050 22.050 ;
        RECT 799.950 20.400 814.050 21.450 ;
        RECT 799.950 19.950 802.050 20.400 ;
        RECT 811.950 19.950 814.050 20.400 ;
        RECT 817.950 16.950 820.050 22.050 ;
        RECT 832.950 21.450 835.050 22.050 ;
        RECT 847.950 21.450 850.050 22.050 ;
        RECT 832.950 20.400 850.050 21.450 ;
        RECT 832.950 19.950 835.050 20.400 ;
        RECT 847.950 19.950 850.050 20.400 ;
        RECT 793.950 15.450 796.050 16.050 ;
        RECT 841.950 15.450 844.050 16.050 ;
        RECT 793.950 14.400 844.050 15.450 ;
        RECT 793.950 13.950 796.050 14.400 ;
        RECT 841.950 13.950 844.050 14.400 ;
        RECT 640.950 10.950 643.050 11.400 ;
        RECT 709.950 10.950 712.050 11.400 ;
        RECT 205.950 8.400 241.050 9.450 ;
        RECT 205.950 7.950 208.050 8.400 ;
        RECT 238.950 7.950 241.050 8.400 ;
        RECT 625.950 9.450 628.050 10.050 ;
        RECT 646.950 9.450 649.050 10.050 ;
        RECT 751.950 9.600 754.050 11.700 ;
        RECT 772.950 10.500 775.050 12.600 ;
        RECT 784.950 12.450 787.050 13.050 ;
        RECT 826.950 12.450 829.050 13.050 ;
        RECT 784.950 11.400 829.050 12.450 ;
        RECT 784.950 10.950 787.050 11.400 ;
        RECT 826.950 10.950 829.050 11.400 ;
        RECT 625.950 8.400 649.050 9.450 ;
        RECT 625.950 7.950 628.050 8.400 ;
        RECT 646.950 7.950 649.050 8.400 ;
        RECT 37.950 6.450 40.050 7.050 ;
        RECT 127.950 6.450 130.050 7.050 ;
        RECT 37.950 5.400 130.050 6.450 ;
        RECT 37.950 4.950 40.050 5.400 ;
        RECT 127.950 4.950 130.050 5.400 ;
        RECT 442.950 6.450 445.050 7.050 ;
        RECT 517.950 6.450 520.050 7.050 ;
        RECT 442.950 5.400 520.050 6.450 ;
        RECT 442.950 4.950 445.050 5.400 ;
        RECT 517.950 4.950 520.050 5.400 ;
        RECT 610.950 6.450 613.050 7.050 ;
        RECT 766.950 6.450 769.050 7.050 ;
        RECT 610.950 5.400 769.050 6.450 ;
        RECT 610.950 4.950 613.050 5.400 ;
        RECT 766.950 4.950 769.050 5.400 ;
        RECT 772.950 6.450 775.050 7.050 ;
        RECT 853.950 6.450 856.050 7.050 ;
        RECT 772.950 5.400 856.050 6.450 ;
        RECT 772.950 4.950 775.050 5.400 ;
        RECT 853.950 4.950 856.050 5.400 ;
        RECT 448.950 3.450 451.050 4.050 ;
        RECT 463.950 3.450 466.050 4.050 ;
        RECT 448.950 2.400 466.050 3.450 ;
        RECT 448.950 1.950 451.050 2.400 ;
        RECT 463.950 1.950 466.050 2.400 ;
        RECT 679.950 3.450 682.050 4.050 ;
        RECT 814.950 3.450 817.050 4.050 ;
        RECT 679.950 2.400 817.050 3.450 ;
        RECT 679.950 1.950 682.050 2.400 ;
        RECT 814.950 1.950 817.050 2.400 ;
      LAYER metal3 ;
        RECT 640.950 865.950 643.050 868.050 ;
        RECT 718.950 865.950 721.050 868.050 ;
        RECT 739.950 865.950 742.050 868.050 ;
        RECT 814.950 865.950 817.050 868.050 ;
        RECT 601.950 862.950 604.050 865.050 ;
        RECT 634.950 862.950 637.050 865.050 ;
        RECT 226.950 859.950 229.050 862.050 ;
        RECT 283.950 859.950 286.050 862.050 ;
        RECT 88.950 856.950 91.050 859.050 ;
        RECT 196.950 856.950 199.050 859.050 ;
        RECT 46.950 850.950 49.050 853.050 ;
        RECT 47.400 847.050 48.600 850.950 ;
        RECT 7.950 844.950 10.050 847.050 ;
        RECT 46.950 844.950 49.050 847.050 ;
        RECT 58.950 844.950 61.050 847.050 ;
        RECT 77.100 844.950 79.200 847.050 ;
        RECT 8.400 823.050 9.600 844.950 ;
        RECT 28.950 841.950 31.050 844.050 ;
        RECT 34.950 841.950 37.050 844.050 ;
        RECT 49.950 841.950 52.050 844.050 ;
        RECT 29.400 835.050 30.600 841.950 ;
        RECT 35.400 838.050 36.600 841.950 ;
        RECT 34.950 835.950 37.050 838.050 ;
        RECT 50.400 835.050 51.600 841.950 ;
        RECT 59.400 838.050 60.600 844.950 ;
        RECT 72.000 843.600 75.900 844.050 ;
        RECT 71.400 841.950 75.900 843.600 ;
        RECT 58.950 835.950 61.050 838.050 ;
        RECT 28.950 832.950 31.050 835.050 ;
        RECT 49.950 832.950 52.050 835.050 ;
        RECT 34.950 829.950 37.050 832.050 ;
        RECT 7.950 820.950 10.050 823.050 ;
        RECT 8.400 817.050 9.600 820.950 ;
        RECT 7.950 814.950 10.050 817.050 ;
        RECT 13.950 814.950 16.050 817.050 ;
        RECT 14.400 787.050 15.600 814.950 ;
        RECT 35.400 814.050 36.600 829.950 ;
        RECT 40.950 823.950 43.050 826.050 ;
        RECT 21.000 813.600 25.050 814.050 ;
        RECT 20.400 811.950 25.050 813.600 ;
        RECT 31.950 812.400 36.600 814.050 ;
        RECT 41.400 814.050 42.600 823.950 ;
        RECT 41.400 812.400 46.050 814.050 ;
        RECT 31.950 811.950 36.000 812.400 ;
        RECT 42.000 811.950 46.050 812.400 ;
        RECT 16.950 808.950 19.050 811.050 ;
        RECT 17.400 790.050 18.600 808.950 ;
        RECT 16.950 787.950 19.050 790.050 ;
        RECT 13.950 784.950 16.050 787.050 ;
        RECT 20.400 784.050 21.600 811.950 ;
        RECT 52.950 805.950 55.050 811.050 ;
        RECT 59.400 808.050 60.600 835.950 ;
        RECT 71.400 826.050 72.600 841.950 ;
        RECT 77.400 841.050 78.600 844.950 ;
        RECT 76.950 838.950 79.050 841.050 ;
        RECT 82.950 838.950 85.050 841.050 ;
        RECT 77.400 829.050 78.600 838.950 ;
        RECT 83.400 835.050 84.600 838.950 ;
        RECT 82.950 832.950 85.050 835.050 ;
        RECT 76.950 826.950 79.050 829.050 ;
        RECT 70.950 823.950 73.050 826.050 ;
        RECT 89.400 817.050 90.600 856.950 ;
        RECT 91.950 853.950 94.050 856.050 ;
        RECT 92.400 844.050 93.600 853.950 ;
        RECT 130.950 850.950 133.050 853.050 ;
        RECT 118.950 847.950 121.050 850.050 ;
        RECT 119.400 844.050 120.600 847.950 ;
        RECT 131.400 847.050 132.600 850.950 ;
        RECT 138.000 849.600 142.050 850.050 ;
        RECT 137.400 847.950 142.050 849.600 ;
        RECT 151.950 847.950 154.050 853.050 ;
        RECT 130.800 844.950 132.900 847.050 ;
        RECT 91.800 841.950 93.900 844.050 ;
        RECT 95.100 841.950 97.200 844.050 ;
        RECT 118.950 841.950 121.050 844.050 ;
        RECT 134.100 841.950 136.200 844.050 ;
        RECT 95.400 835.050 96.600 841.950 ;
        RECT 103.950 838.950 106.050 841.050 ;
        RECT 94.950 832.950 97.050 835.050 ;
        RECT 104.400 832.050 105.600 838.950 ;
        RECT 134.400 838.050 135.600 841.950 ;
        RECT 133.950 835.950 136.050 838.050 ;
        RECT 124.950 832.950 127.050 835.050 ;
        RECT 103.950 829.950 106.050 832.050 ;
        RECT 109.950 826.950 112.050 829.050 ;
        RECT 100.950 820.950 103.050 823.050 ;
        RECT 79.800 814.950 81.900 817.050 ;
        RECT 88.950 814.950 91.050 817.050 ;
        RECT 80.400 808.050 81.600 814.950 ;
        RECT 101.400 814.050 102.600 820.950 ;
        RECT 103.950 817.950 106.050 820.050 ;
        RECT 104.400 814.050 105.600 817.950 ;
        RECT 100.800 811.950 102.900 814.050 ;
        RECT 104.100 811.950 106.200 814.050 ;
        RECT 110.400 811.050 111.600 826.950 ;
        RECT 112.950 817.950 115.050 820.050 ;
        RECT 106.950 809.400 111.600 811.050 ;
        RECT 106.950 808.950 111.000 809.400 ;
        RECT 58.950 805.950 61.050 808.050 ;
        RECT 79.950 805.950 82.050 808.050 ;
        RECT 19.950 781.950 22.050 784.050 ;
        RECT 49.950 781.950 52.050 784.050 ;
        RECT 50.400 778.050 51.600 781.950 ;
        RECT 10.950 772.950 13.050 778.050 ;
        RECT 25.950 777.600 30.000 778.050 ;
        RECT 36.000 777.600 40.050 778.050 ;
        RECT 25.950 775.950 30.600 777.600 ;
        RECT 19.950 771.600 22.050 772.050 ;
        RECT 14.400 770.400 22.050 771.600 ;
        RECT 14.400 763.050 15.600 770.400 ;
        RECT 19.950 769.950 22.050 770.400 ;
        RECT 22.950 766.950 25.050 769.050 ;
        RECT 13.950 760.950 16.050 763.050 ;
        RECT 14.400 742.050 15.600 760.950 ;
        RECT 23.400 748.050 24.600 766.950 ;
        RECT 29.400 754.050 30.600 775.950 ;
        RECT 35.400 775.950 40.050 777.600 ;
        RECT 49.950 775.950 52.050 778.050 ;
        RECT 35.400 763.050 36.600 775.950 ;
        RECT 43.950 771.600 48.000 772.050 ;
        RECT 43.950 769.950 48.600 771.600 ;
        RECT 53.400 771.000 57.600 771.600 ;
        RECT 34.950 760.950 37.050 763.050 ;
        RECT 28.950 751.950 31.050 754.050 ;
        RECT 47.400 751.050 48.600 769.950 ;
        RECT 52.950 770.400 57.600 771.000 ;
        RECT 52.950 766.950 55.050 770.400 ;
        RECT 46.950 748.950 49.050 751.050 ;
        RECT 22.950 745.950 25.050 748.050 ;
        RECT 25.950 742.950 28.050 745.050 ;
        RECT 48.000 744.600 51.900 745.050 ;
        RECT 47.400 742.950 51.900 744.600 ;
        RECT 4.950 739.950 7.050 742.050 ;
        RECT 10.950 740.400 15.600 742.050 ;
        RECT 10.950 739.950 15.000 740.400 ;
        RECT 5.400 670.050 6.600 739.950 ;
        RECT 26.400 739.050 27.600 742.950 ;
        RECT 30.000 741.600 33.900 742.050 ;
        RECT 29.400 739.950 33.900 741.600 ;
        RECT 25.950 736.950 28.050 739.050 ;
        RECT 10.950 733.950 13.050 736.050 ;
        RECT 16.950 733.950 19.050 736.050 ;
        RECT 11.400 727.050 12.600 733.950 ;
        RECT 10.950 724.950 13.050 727.050 ;
        RECT 7.950 721.950 10.050 724.050 ;
        RECT 8.400 703.050 9.600 721.950 ;
        RECT 17.400 709.050 18.600 733.950 ;
        RECT 29.400 733.050 30.600 739.950 ;
        RECT 28.950 730.950 31.050 733.050 ;
        RECT 22.950 724.950 25.050 727.050 ;
        RECT 16.950 706.950 19.050 709.050 ;
        RECT 23.400 703.050 24.600 724.950 ;
        RECT 32.400 703.050 33.600 739.950 ;
        RECT 47.400 733.050 48.600 742.950 ;
        RECT 56.400 742.050 57.600 770.400 ;
        RECT 59.400 745.050 60.600 805.950 ;
        RECT 61.950 802.950 64.050 805.050 ;
        RECT 62.400 760.050 63.600 802.950 ;
        RECT 113.400 796.050 114.600 817.950 ;
        RECT 125.400 814.050 126.600 832.950 ;
        RECT 137.400 826.050 138.600 847.950 ;
        RECT 142.950 844.950 145.050 847.050 ;
        RECT 160.950 844.950 163.050 847.050 ;
        RECT 166.950 846.600 171.000 847.050 ;
        RECT 166.950 844.950 171.600 846.600 ;
        RECT 178.950 844.950 181.050 847.050 ;
        RECT 143.400 835.050 144.600 844.950 ;
        RECT 148.950 838.950 151.050 841.050 ;
        RECT 142.950 832.950 145.050 835.050 ;
        RECT 136.950 823.950 139.050 826.050 ;
        RECT 133.950 816.600 138.000 817.050 ;
        RECT 133.950 814.950 138.600 816.600 ;
        RECT 115.950 811.950 118.050 814.050 ;
        RECT 124.950 811.950 127.050 814.050 ;
        RECT 130.950 811.950 133.050 814.050 ;
        RECT 116.400 808.050 117.600 811.950 ;
        RECT 115.950 805.950 118.050 808.050 ;
        RECT 131.400 799.050 132.600 811.950 ;
        RECT 137.400 808.050 138.600 814.950 ;
        RECT 136.950 805.950 139.050 808.050 ;
        RECT 130.950 796.950 133.050 799.050 ;
        RECT 112.950 793.950 115.050 796.050 ;
        RECT 133.950 793.950 136.050 796.050 ;
        RECT 70.950 781.950 73.050 784.050 ;
        RECT 71.400 775.050 72.600 781.950 ;
        RECT 115.950 778.050 118.050 781.050 ;
        RECT 85.950 775.950 88.050 778.050 ;
        RECT 115.950 777.000 118.200 778.050 ;
        RECT 116.100 775.950 118.200 777.000 ;
        RECT 70.950 772.950 73.050 775.050 ;
        RECT 64.950 766.950 67.050 772.050 ;
        RECT 61.950 757.950 64.050 760.050 ;
        RECT 86.400 745.050 87.600 775.950 ;
        RECT 134.400 775.050 135.600 793.950 ;
        RECT 143.400 790.050 144.600 832.950 ;
        RECT 149.400 799.050 150.600 838.950 ;
        RECT 161.400 835.050 162.600 844.950 ;
        RECT 170.400 838.050 171.600 844.950 ;
        RECT 169.950 835.950 172.050 838.050 ;
        RECT 160.950 832.950 163.050 835.050 ;
        RECT 170.400 823.050 171.600 835.950 ;
        RECT 179.400 832.050 180.600 844.950 ;
        RECT 193.950 841.950 196.050 844.050 ;
        RECT 181.950 838.950 184.050 841.050 ;
        RECT 182.400 835.050 183.600 838.950 ;
        RECT 181.950 832.950 184.050 835.050 ;
        RECT 178.950 829.950 181.050 832.050 ;
        RECT 169.950 820.950 172.050 823.050 ;
        RECT 175.950 817.950 178.050 820.050 ;
        RECT 157.950 808.950 160.050 814.050 ;
        RECT 163.950 811.950 166.050 814.050 ;
        RECT 164.400 808.050 165.600 811.950 ;
        RECT 176.400 808.050 177.600 817.950 ;
        RECT 163.950 805.950 166.050 808.050 ;
        RECT 169.950 805.950 172.050 808.050 ;
        RECT 166.950 799.950 169.050 802.050 ;
        RECT 148.950 796.950 151.050 799.050 ;
        RECT 142.950 787.950 145.050 790.050 ;
        RECT 167.400 781.050 168.600 799.950 ;
        RECT 170.400 787.050 171.600 805.950 ;
        RECT 175.950 802.950 178.050 808.050 ;
        RECT 169.950 784.950 172.050 787.050 ;
        RECT 166.950 778.950 169.050 781.050 ;
        RECT 91.950 772.950 94.050 775.050 ;
        RECT 111.000 774.600 114.900 775.050 ;
        RECT 110.400 772.950 114.900 774.600 ;
        RECT 133.800 774.000 135.900 775.050 ;
        RECT 133.800 772.950 136.050 774.000 ;
        RECT 145.950 772.950 148.050 775.050 ;
        RECT 92.400 754.050 93.600 772.950 ;
        RECT 100.800 769.950 102.900 772.050 ;
        RECT 101.400 763.050 102.600 769.950 ;
        RECT 100.950 760.950 103.050 763.050 ;
        RECT 110.400 757.050 111.600 772.950 ;
        RECT 133.950 771.000 136.050 772.950 ;
        RECT 134.400 770.400 135.600 771.000 ;
        RECT 118.950 763.950 121.050 769.050 ;
        RECT 127.950 766.950 130.050 769.050 ;
        RECT 115.950 760.950 118.050 763.050 ;
        RECT 109.950 754.950 112.050 757.050 ;
        RECT 91.950 751.950 94.050 754.050 ;
        RECT 58.950 742.950 61.050 745.050 ;
        RECT 73.950 744.600 78.000 745.050 ;
        RECT 73.950 742.950 78.600 744.600 ;
        RECT 85.950 742.950 88.050 745.050 ;
        RECT 94.950 742.950 97.050 745.050 ;
        RECT 55.950 739.950 58.050 742.050 ;
        RECT 70.950 739.950 73.050 742.050 ;
        RECT 52.950 736.950 55.050 739.050 ;
        RECT 46.950 730.950 49.050 733.050 ;
        RECT 53.400 715.050 54.600 736.950 ;
        RECT 58.950 727.950 61.050 730.050 ;
        RECT 67.950 727.950 70.050 730.050 ;
        RECT 52.950 712.950 55.050 715.050 ;
        RECT 49.950 703.950 52.050 706.050 ;
        RECT 7.950 700.950 10.050 703.050 ;
        RECT 22.950 700.950 25.050 703.050 ;
        RECT 32.100 700.950 34.200 703.050 ;
        RECT 50.400 700.050 51.600 703.950 ;
        RECT 59.400 703.050 60.600 727.950 ;
        RECT 55.800 701.400 60.600 703.050 ;
        RECT 55.800 700.950 60.000 701.400 ;
        RECT 61.950 700.950 64.050 703.050 ;
        RECT 13.950 697.950 16.050 700.050 ;
        RECT 49.950 697.950 52.050 700.050 ;
        RECT 10.950 691.950 13.050 694.050 ;
        RECT 11.400 673.050 12.600 691.950 ;
        RECT 14.400 682.050 15.600 697.950 ;
        RECT 55.950 694.950 58.050 697.050 ;
        RECT 49.950 691.950 52.050 694.050 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 34.950 676.950 37.050 679.050 ;
        RECT 19.950 673.950 22.050 676.050 ;
        RECT 10.950 670.950 13.050 673.050 ;
        RECT 4.950 667.950 7.050 670.050 ;
        RECT 20.400 667.050 21.600 673.950 ;
        RECT 31.800 667.950 33.900 670.050 ;
        RECT 19.950 664.950 22.050 667.050 ;
        RECT 13.950 631.950 16.050 637.050 ;
        RECT 25.950 631.950 28.050 634.050 ;
        RECT 21.000 630.600 25.050 631.050 ;
        RECT 20.400 628.950 25.050 630.600 ;
        RECT 20.400 625.050 21.600 628.950 ;
        RECT 20.100 622.950 22.200 625.050 ;
        RECT 16.950 607.950 19.050 610.050 ;
        RECT 17.400 604.050 18.600 607.950 ;
        RECT 26.400 607.050 27.600 631.950 ;
        RECT 32.400 628.050 33.600 667.950 ;
        RECT 35.400 667.050 36.600 676.950 ;
        RECT 40.950 673.050 43.050 673.200 ;
        RECT 39.000 672.750 43.050 673.050 ;
        RECT 38.400 671.100 43.050 672.750 ;
        RECT 38.400 670.950 42.000 671.100 ;
        RECT 35.100 664.950 37.200 667.050 ;
        RECT 38.400 664.050 39.600 670.950 ;
        RECT 42.000 669.600 46.050 670.050 ;
        RECT 41.400 667.950 46.050 669.600 ;
        RECT 37.950 661.950 40.050 664.050 ;
        RECT 41.400 646.050 42.600 667.950 ;
        RECT 40.950 643.950 43.050 646.050 ;
        RECT 37.950 634.950 40.050 640.050 ;
        RECT 42.000 630.600 46.050 631.050 ;
        RECT 41.400 628.950 46.050 630.600 ;
        RECT 31.950 627.600 34.050 628.050 ;
        RECT 31.950 626.400 36.600 627.600 ;
        RECT 31.950 625.950 34.050 626.400 ;
        RECT 25.950 604.950 28.050 607.050 ;
        RECT 16.950 601.950 19.050 604.050 ;
        RECT 7.950 594.600 12.000 595.050 ;
        RECT 7.950 592.950 12.600 594.600 ;
        RECT 1.950 556.950 4.050 559.050 ;
        RECT 2.400 436.050 3.600 556.950 ;
        RECT 11.400 538.050 12.600 592.950 ;
        RECT 17.400 592.050 18.600 601.950 ;
        RECT 26.400 598.050 27.600 604.950 ;
        RECT 28.800 598.950 30.900 601.050 ;
        RECT 25.950 595.950 28.050 598.050 ;
        RECT 16.950 589.950 19.050 592.050 ;
        RECT 22.950 589.950 25.050 592.050 ;
        RECT 16.950 577.950 19.050 580.050 ;
        RECT 17.400 556.050 18.600 577.950 ;
        RECT 23.400 559.050 24.600 589.950 ;
        RECT 29.400 589.050 30.600 598.950 ;
        RECT 28.950 586.950 31.050 589.050 ;
        RECT 28.950 571.950 31.050 574.050 ;
        RECT 22.950 556.950 25.050 559.050 ;
        RECT 17.400 554.400 22.050 556.050 ;
        RECT 18.000 553.950 22.050 554.400 ;
        RECT 25.950 553.950 28.050 556.050 ;
        RECT 10.950 535.950 13.050 538.050 ;
        RECT 26.400 532.050 27.600 553.950 ;
        RECT 25.950 529.950 28.050 532.050 ;
        RECT 29.400 529.050 30.600 571.950 ;
        RECT 35.400 571.050 36.600 626.400 ;
        RECT 41.400 622.050 42.600 628.950 ;
        RECT 40.950 619.950 43.050 622.050 ;
        RECT 41.400 616.050 42.600 619.950 ;
        RECT 40.950 613.950 43.050 616.050 ;
        RECT 50.400 613.050 51.600 691.950 ;
        RECT 56.400 679.050 57.600 694.950 ;
        RECT 62.400 694.050 63.600 700.950 ;
        RECT 68.400 700.050 69.600 727.950 ;
        RECT 71.400 724.050 72.600 739.950 ;
        RECT 77.400 736.050 78.600 742.950 ;
        RECT 81.000 741.600 85.050 742.050 ;
        RECT 80.400 739.950 85.050 741.600 ;
        RECT 91.950 739.950 94.050 742.050 ;
        RECT 76.950 733.950 79.050 736.050 ;
        RECT 80.400 727.050 81.600 739.950 ;
        RECT 79.950 724.950 82.050 727.050 ;
        RECT 92.400 724.050 93.600 739.950 ;
        RECT 70.950 721.950 73.050 724.050 ;
        RECT 91.950 721.950 94.050 724.050 ;
        RECT 91.950 712.950 94.050 715.050 ;
        RECT 92.400 706.050 93.600 712.950 ;
        RECT 95.400 709.050 96.600 742.950 ;
        RECT 106.950 739.950 109.050 742.050 ;
        RECT 101.100 736.950 103.200 739.050 ;
        RECT 97.800 733.950 99.900 736.050 ;
        RECT 98.400 718.050 99.600 733.950 ;
        RECT 101.400 727.050 102.600 736.950 ;
        RECT 107.400 733.050 108.600 739.950 ;
        RECT 116.400 739.050 117.600 760.950 ;
        RECT 128.400 757.050 129.600 766.950 ;
        RECT 127.950 754.950 130.050 757.050 ;
        RECT 128.400 748.050 129.600 754.950 ;
        RECT 128.400 746.400 133.050 748.050 ;
        RECT 129.000 745.950 133.050 746.400 ;
        RECT 146.400 745.050 147.600 772.950 ;
        RECT 179.400 772.050 180.600 829.950 ;
        RECT 194.400 826.050 195.600 841.950 ;
        RECT 193.950 823.950 196.050 826.050 ;
        RECT 181.950 820.950 184.050 823.050 ;
        RECT 182.400 796.050 183.600 820.950 ;
        RECT 184.950 814.950 187.050 817.050 ;
        RECT 181.950 793.950 184.050 796.050 ;
        RECT 185.400 790.050 186.600 814.950 ;
        RECT 194.400 811.050 195.600 823.950 ;
        RECT 197.400 820.050 198.600 856.950 ;
        RECT 211.950 847.950 214.050 850.050 ;
        RECT 220.950 847.950 223.050 850.050 ;
        RECT 212.400 838.050 213.600 847.950 ;
        RECT 214.950 838.950 217.050 841.050 ;
        RECT 211.950 835.950 214.050 838.050 ;
        RECT 196.950 817.950 199.050 820.050 ;
        RECT 201.000 813.600 205.050 814.050 ;
        RECT 200.400 811.950 205.050 813.600 ;
        RECT 208.950 811.950 211.050 814.050 ;
        RECT 193.950 808.950 196.050 811.050 ;
        RECT 194.400 799.050 195.600 808.950 ;
        RECT 193.950 796.950 196.050 799.050 ;
        RECT 184.950 787.950 187.050 790.050 ;
        RECT 193.950 784.950 196.050 787.050 ;
        RECT 184.950 778.950 187.050 781.050 ;
        RECT 154.950 769.950 157.050 772.050 ;
        RECT 166.950 771.600 171.000 772.050 ;
        RECT 166.950 769.950 171.600 771.600 ;
        RECT 179.100 769.950 181.200 772.050 ;
        RECT 155.400 750.600 156.600 769.950 ;
        RECT 160.950 766.950 163.050 769.050 ;
        RECT 157.950 750.600 160.050 751.050 ;
        RECT 155.400 749.400 160.050 750.600 ;
        RECT 157.950 748.950 160.050 749.400 ;
        RECT 145.950 742.050 148.050 745.050 ;
        RECT 145.800 741.000 148.050 742.050 ;
        RECT 145.800 739.950 147.900 741.000 ;
        RECT 151.950 739.950 154.050 742.050 ;
        RECT 115.950 736.950 118.050 739.050 ;
        RECT 152.400 733.050 153.600 739.950 ;
        RECT 158.400 739.050 159.600 748.950 ;
        RECT 161.400 748.050 162.600 766.950 ;
        RECT 170.400 751.050 171.600 769.950 ;
        RECT 176.100 766.950 178.200 769.050 ;
        RECT 176.400 754.050 177.600 766.950 ;
        RECT 175.950 751.950 178.050 754.050 ;
        RECT 169.950 748.950 172.050 751.050 ;
        RECT 160.950 745.950 163.050 748.050 ;
        RECT 172.950 739.950 175.050 742.050 ;
        RECT 157.950 736.950 160.050 739.050 ;
        RECT 173.400 733.050 174.600 739.950 ;
        RECT 106.950 730.950 109.050 733.050 ;
        RECT 151.950 730.950 154.050 733.050 ;
        RECT 172.950 730.950 175.050 733.050 ;
        RECT 100.950 724.950 103.050 727.050 ;
        RECT 103.950 721.950 106.050 724.050 ;
        RECT 97.950 715.950 100.050 718.050 ;
        RECT 95.100 706.950 97.200 709.050 ;
        RECT 91.800 703.950 93.900 706.050 ;
        RECT 82.950 700.950 85.050 703.050 ;
        RECT 67.950 697.950 70.050 700.050 ;
        RECT 77.400 699.000 78.600 699.600 ;
        RECT 76.950 694.950 79.050 699.000 ;
        RECT 61.950 691.950 64.050 694.050 ;
        RECT 77.400 685.050 78.600 694.950 ;
        RECT 83.400 694.050 84.600 700.950 ;
        RECT 97.950 697.950 100.050 700.050 ;
        RECT 98.400 694.050 99.600 697.950 ;
        RECT 82.950 691.950 85.050 694.050 ;
        RECT 97.950 691.950 100.050 694.050 ;
        RECT 76.950 682.950 79.050 685.050 ;
        RECT 55.950 676.950 58.050 679.050 ;
        RECT 73.950 670.950 76.050 673.050 ;
        RECT 52.950 664.950 55.050 670.050 ;
        RECT 58.950 667.950 61.050 670.050 ;
        RECT 53.400 637.050 54.600 664.950 ;
        RECT 59.400 643.050 60.600 667.950 ;
        RECT 64.950 664.950 67.050 667.050 ;
        RECT 58.950 640.950 61.050 643.050 ;
        RECT 52.950 634.950 55.050 637.050 ;
        RECT 59.100 628.950 61.200 631.050 ;
        RECT 49.950 610.950 52.050 613.050 ;
        RECT 52.950 607.950 55.050 610.050 ;
        RECT 49.950 604.950 52.050 607.050 ;
        RECT 50.400 598.050 51.600 604.950 ;
        RECT 46.950 596.400 51.600 598.050 ;
        RECT 46.950 595.950 51.000 596.400 ;
        RECT 53.400 595.050 54.600 607.950 ;
        RECT 59.400 607.050 60.600 628.950 ;
        RECT 58.950 604.950 61.050 607.050 ;
        RECT 53.400 593.400 58.050 595.050 ;
        RECT 54.000 592.950 58.050 593.400 ;
        RECT 40.950 586.950 43.050 589.050 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 35.400 562.050 36.600 568.950 ;
        RECT 34.950 559.950 37.050 562.050 ;
        RECT 41.400 559.050 42.600 586.950 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 53.400 559.050 54.600 568.950 ;
        RECT 40.950 556.950 43.050 559.050 ;
        RECT 53.100 556.950 55.200 559.050 ;
        RECT 47.100 553.950 49.200 556.050 ;
        RECT 55.800 553.950 57.900 556.050 ;
        RECT 47.400 547.050 48.600 553.950 ;
        RECT 56.400 550.050 57.600 553.950 ;
        RECT 55.950 547.950 58.050 550.050 ;
        RECT 46.950 544.950 49.050 547.050 ;
        RECT 34.950 535.950 37.050 538.050 ;
        RECT 35.400 529.050 36.600 535.950 ;
        RECT 7.950 528.600 12.000 529.050 ;
        RECT 7.950 526.950 12.600 528.600 ;
        RECT 14.100 526.950 16.200 529.050 ;
        RECT 20.100 528.000 22.200 529.050 ;
        RECT 19.950 526.950 22.200 528.000 ;
        RECT 28.950 526.950 31.050 529.050 ;
        RECT 34.950 526.950 37.050 529.050 ;
        RECT 11.400 493.050 12.600 526.950 ;
        RECT 14.400 520.050 15.600 526.950 ;
        RECT 19.950 526.050 22.050 526.950 ;
        RECT 16.800 525.000 22.050 526.050 ;
        RECT 16.800 524.400 21.600 525.000 ;
        RECT 16.800 523.950 21.000 524.400 ;
        RECT 28.800 522.600 30.900 523.050 ;
        RECT 35.400 522.600 36.600 526.950 ;
        RECT 28.800 521.400 36.600 522.600 ;
        RECT 28.800 520.950 30.900 521.400 ;
        RECT 13.950 517.950 16.050 520.050 ;
        RECT 43.950 514.950 46.050 517.050 ;
        RECT 28.950 508.950 31.050 511.050 ;
        RECT 16.950 502.950 19.050 505.050 ;
        RECT 10.950 490.950 13.050 493.050 ;
        RECT 7.950 486.600 12.000 487.050 ;
        RECT 7.950 484.950 12.600 486.600 ;
        RECT 11.400 445.050 12.600 484.950 ;
        RECT 17.400 484.050 18.600 502.950 ;
        RECT 29.400 487.050 30.600 508.950 ;
        RECT 34.950 490.950 37.050 493.050 ;
        RECT 35.400 487.050 36.600 490.950 ;
        RECT 44.400 487.050 45.600 514.950 ;
        RECT 28.800 484.950 30.900 487.050 ;
        RECT 34.800 484.950 36.900 487.050 ;
        RECT 43.950 484.950 46.050 487.050 ;
        RECT 16.800 481.950 18.900 484.050 ;
        RECT 28.950 469.950 31.050 472.050 ;
        RECT 22.950 463.950 25.050 466.050 ;
        RECT 23.400 457.050 24.600 463.950 ;
        RECT 22.950 454.950 25.050 457.050 ;
        RECT 29.400 451.050 30.600 469.950 ;
        RECT 44.400 463.050 45.600 484.950 ;
        RECT 43.950 460.950 46.050 463.050 ;
        RECT 33.000 453.600 37.050 454.050 ;
        RECT 25.950 449.400 30.600 451.050 ;
        RECT 32.400 451.950 37.050 453.600 ;
        RECT 25.950 448.950 30.000 449.400 ;
        RECT 10.950 442.950 13.050 445.050 ;
        RECT 28.950 436.950 31.050 439.050 ;
        RECT 1.950 433.950 4.050 436.050 ;
        RECT 10.950 433.950 13.050 436.050 ;
        RECT 11.400 429.600 12.600 433.950 ;
        RECT 11.400 428.400 15.600 429.600 ;
        RECT 7.950 421.950 10.050 424.050 ;
        RECT 8.400 415.050 9.600 421.950 ;
        RECT 14.400 415.050 15.600 428.400 ;
        RECT 19.950 424.950 22.050 427.050 ;
        RECT 7.950 412.950 10.050 415.050 ;
        RECT 13.800 414.000 15.900 415.050 ;
        RECT 13.800 412.950 16.050 414.000 ;
        RECT 13.950 411.000 16.050 412.950 ;
        RECT 20.400 412.050 21.600 424.950 ;
        RECT 25.950 421.950 28.050 424.050 ;
        RECT 14.400 410.400 15.600 411.000 ;
        RECT 20.400 410.400 24.900 412.050 ;
        RECT 21.000 409.950 24.900 410.400 ;
        RECT 19.950 388.950 22.050 391.050 ;
        RECT 13.950 382.950 16.050 388.050 ;
        RECT 20.400 385.050 21.600 388.950 ;
        RECT 19.950 382.950 22.050 385.050 ;
        RECT 4.950 376.950 7.050 379.050 ;
        RECT 16.950 376.950 19.050 379.050 ;
        RECT 5.400 322.050 6.600 376.950 ;
        RECT 13.950 364.950 16.050 367.050 ;
        RECT 14.400 346.200 15.600 364.950 ;
        RECT 7.950 345.600 12.000 346.050 ;
        RECT 7.950 343.950 12.600 345.600 ;
        RECT 14.100 344.100 16.200 346.200 ;
        RECT 4.950 319.950 7.050 322.050 ;
        RECT 11.400 319.050 12.600 343.950 ;
        RECT 17.400 342.600 18.600 376.950 ;
        RECT 23.400 349.050 24.600 409.950 ;
        RECT 26.400 391.050 27.600 421.950 ;
        RECT 25.950 388.950 28.050 391.050 ;
        RECT 29.400 385.050 30.600 436.950 ;
        RECT 32.400 427.200 33.600 451.950 ;
        RECT 44.100 448.950 46.200 451.050 ;
        RECT 40.950 442.950 43.050 445.050 ;
        RECT 37.950 439.950 40.050 442.050 ;
        RECT 31.950 425.100 34.050 427.200 ;
        RECT 31.950 421.800 34.050 423.900 ;
        RECT 32.400 421.050 33.600 421.800 ;
        RECT 31.950 417.000 34.050 421.050 ;
        RECT 32.400 416.400 33.600 417.000 ;
        RECT 33.000 414.900 36.000 415.050 ;
        RECT 31.950 414.450 36.000 414.900 ;
        RECT 31.950 412.950 36.600 414.450 ;
        RECT 31.950 412.800 34.050 412.950 ;
        RECT 35.400 406.050 36.600 412.950 ;
        RECT 34.950 403.950 37.050 406.050 ;
        RECT 28.800 382.950 30.900 385.050 ;
        RECT 25.800 379.950 27.900 382.050 ;
        RECT 26.400 367.050 27.600 379.950 ;
        RECT 25.950 364.950 28.050 367.050 ;
        RECT 22.950 346.950 25.050 349.050 ;
        RECT 23.400 343.050 24.600 346.950 ;
        RECT 29.400 343.200 30.600 382.950 ;
        RECT 32.100 381.000 34.200 382.050 ;
        RECT 31.950 379.950 34.200 381.000 ;
        RECT 31.950 376.950 34.050 379.950 ;
        RECT 38.400 361.050 39.600 439.950 ;
        RECT 37.950 358.950 40.050 361.050 ;
        RECT 14.400 342.000 18.600 342.600 ;
        RECT 13.950 341.400 18.600 342.000 ;
        RECT 13.950 337.950 16.050 341.400 ;
        RECT 22.950 340.950 25.050 343.050 ;
        RECT 28.950 341.100 31.050 343.200 ;
        RECT 28.950 337.800 31.050 339.900 ;
        RECT 16.950 319.950 19.050 322.050 ;
        RECT 10.950 316.950 13.050 319.050 ;
        RECT 17.400 316.050 18.600 319.950 ;
        RECT 22.950 316.950 25.050 319.050 ;
        RECT 17.100 313.950 19.200 316.050 ;
        RECT 13.800 310.950 15.900 313.050 ;
        RECT 4.950 307.950 7.050 310.050 ;
        RECT 5.400 304.050 6.600 307.950 ;
        RECT 4.950 301.950 7.050 304.050 ;
        RECT 5.400 241.050 6.600 301.950 ;
        RECT 14.400 289.050 15.600 310.950 ;
        RECT 13.950 286.950 16.050 289.050 ;
        RECT 13.950 277.950 16.050 280.050 ;
        RECT 10.950 274.950 13.050 277.050 ;
        RECT 11.400 265.050 12.600 274.950 ;
        RECT 14.400 268.050 15.600 277.950 ;
        RECT 23.400 277.050 24.600 316.950 ;
        RECT 25.950 313.950 28.050 316.050 ;
        RECT 26.400 310.050 27.600 313.950 ;
        RECT 25.800 307.950 27.900 310.050 ;
        RECT 22.950 274.950 25.050 277.050 ;
        RECT 23.400 271.050 24.600 274.950 ;
        RECT 29.400 274.050 30.600 337.800 ;
        RECT 34.950 316.950 37.050 319.050 ;
        RECT 35.400 313.050 36.600 316.950 ;
        RECT 41.400 313.050 42.600 442.950 ;
        RECT 44.400 421.050 45.600 448.950 ;
        RECT 43.950 418.950 46.050 421.050 ;
        RECT 43.950 409.950 46.050 412.050 ;
        RECT 44.400 388.050 45.600 409.950 ;
        RECT 43.950 385.950 46.050 388.050 ;
        RECT 47.400 385.050 48.600 544.950 ;
        RECT 49.950 526.950 52.050 529.050 ;
        RECT 50.400 523.050 51.600 526.950 ;
        RECT 49.800 520.950 51.900 523.050 ;
        RECT 56.100 520.950 58.200 523.050 ;
        RECT 50.400 490.050 51.600 520.950 ;
        RECT 56.400 517.050 57.600 520.950 ;
        RECT 55.950 514.950 58.050 517.050 ;
        RECT 49.800 487.950 51.900 490.050 ;
        RECT 55.950 481.950 58.050 484.050 ;
        RECT 52.950 460.950 55.050 463.050 ;
        RECT 53.400 454.050 54.600 460.950 ;
        RECT 49.950 452.400 54.600 454.050 ;
        RECT 49.950 451.950 54.000 452.400 ;
        RECT 56.400 445.050 57.600 481.950 ;
        RECT 58.950 454.950 61.050 460.050 ;
        RECT 65.400 457.050 66.600 664.950 ;
        RECT 74.400 664.050 75.600 670.950 ;
        RECT 73.800 663.600 75.900 664.050 ;
        RECT 71.400 662.400 75.900 663.600 ;
        RECT 71.400 649.050 72.600 662.400 ;
        RECT 73.800 661.950 75.900 662.400 ;
        RECT 77.100 661.950 79.200 664.050 ;
        RECT 70.950 646.950 73.050 649.050 ;
        RECT 71.400 637.050 72.600 646.950 ;
        RECT 77.400 643.050 78.600 661.950 ;
        RECT 76.950 640.950 79.050 643.050 ;
        RECT 83.400 639.600 84.600 691.950 ;
        RECT 91.950 688.950 94.050 691.050 ;
        RECT 88.950 676.950 91.050 679.050 ;
        RECT 89.400 667.050 90.600 676.950 ;
        RECT 92.400 673.050 93.600 688.950 ;
        RECT 91.950 670.950 94.050 673.050 ;
        RECT 97.950 670.950 100.050 676.050 ;
        RECT 88.950 664.950 91.050 667.050 ;
        RECT 104.400 664.050 105.600 721.950 ;
        RECT 112.950 712.950 115.050 715.050 ;
        RECT 124.950 712.950 127.050 715.050 ;
        RECT 113.400 706.050 114.600 712.950 ;
        RECT 118.950 709.950 121.050 712.050 ;
        RECT 112.950 703.950 115.050 706.050 ;
        RECT 119.400 703.050 120.600 709.950 ;
        RECT 125.400 703.050 126.600 712.950 ;
        RECT 139.950 709.950 142.050 712.050 ;
        RECT 178.950 709.950 181.050 712.050 ;
        RECT 140.400 703.050 141.600 709.950 ;
        RECT 179.400 706.050 180.600 709.950 ;
        RECT 175.950 704.400 180.600 706.050 ;
        RECT 185.400 706.050 186.600 778.950 ;
        RECT 194.400 778.050 195.600 784.950 ;
        RECT 200.400 784.050 201.600 811.950 ;
        RECT 209.400 802.050 210.600 811.950 ;
        RECT 215.400 802.050 216.600 838.950 ;
        RECT 221.400 832.050 222.600 847.950 ;
        RECT 227.400 847.050 228.600 859.950 ;
        RECT 241.950 850.950 244.050 853.050 ;
        RECT 256.950 850.950 259.050 853.050 ;
        RECT 232.950 847.950 235.050 850.050 ;
        RECT 226.950 844.950 229.050 847.050 ;
        RECT 220.950 829.950 223.050 832.050 ;
        RECT 226.950 826.950 229.050 829.050 ;
        RECT 217.950 814.950 220.050 817.050 ;
        RECT 218.400 811.050 219.600 814.950 ;
        RECT 227.400 814.050 228.600 826.950 ;
        RECT 233.400 820.050 234.600 847.950 ;
        RECT 242.400 847.050 243.600 850.950 ;
        RECT 241.800 844.950 243.900 847.050 ;
        RECT 247.950 841.950 250.050 844.050 ;
        RECT 248.400 838.050 249.600 841.950 ;
        RECT 247.950 835.950 250.050 838.050 ;
        RECT 241.950 832.950 244.050 835.050 ;
        RECT 235.950 820.950 238.050 823.050 ;
        RECT 232.950 817.950 235.050 820.050 ;
        RECT 236.400 814.050 237.600 820.950 ;
        RECT 226.950 811.950 229.050 814.050 ;
        RECT 236.400 812.400 241.050 814.050 ;
        RECT 237.000 811.950 241.050 812.400 ;
        RECT 242.400 811.050 243.600 832.950 ;
        RECT 250.950 814.950 253.050 820.050 ;
        RECT 257.400 817.050 258.600 850.950 ;
        RECT 284.400 847.050 285.600 859.950 ;
        RECT 316.950 853.950 319.050 856.050 ;
        RECT 343.950 853.950 346.050 856.050 ;
        RECT 439.950 853.950 442.050 856.050 ;
        RECT 283.950 844.950 286.050 847.050 ;
        RECT 297.000 843.600 301.050 844.050 ;
        RECT 290.400 843.000 291.600 843.600 ;
        RECT 289.950 838.950 292.050 843.000 ;
        RECT 296.400 841.950 301.050 843.600 ;
        RECT 274.950 829.950 277.050 832.050 ;
        RECT 256.950 814.950 259.050 817.050 ;
        RECT 217.950 808.950 220.050 811.050 ;
        RECT 223.950 808.950 226.050 811.050 ;
        RECT 241.950 808.950 244.050 811.050 ;
        RECT 208.950 799.950 211.050 802.050 ;
        RECT 214.950 799.950 217.050 802.050 ;
        RECT 205.950 796.950 208.050 799.050 ;
        RECT 199.950 781.950 202.050 784.050 ;
        RECT 206.400 778.050 207.600 796.950 ;
        RECT 224.400 793.050 225.600 808.950 ;
        RECT 275.400 808.050 276.600 829.950 ;
        RECT 277.950 820.950 280.050 823.050 ;
        RECT 278.400 817.050 279.600 820.950 ;
        RECT 277.950 813.000 280.050 817.050 ;
        RECT 290.400 814.050 291.600 838.950 ;
        RECT 296.400 838.050 297.600 841.950 ;
        RECT 304.950 838.950 307.050 841.050 ;
        RECT 295.950 835.950 298.050 838.050 ;
        RECT 296.400 829.050 297.600 835.950 ;
        RECT 295.950 826.950 298.050 829.050 ;
        RECT 305.400 820.050 306.600 838.950 ;
        RECT 310.950 829.950 313.050 832.050 ;
        RECT 304.950 817.950 307.050 820.050 ;
        RECT 311.400 817.050 312.600 829.950 ;
        RECT 317.400 817.050 318.600 853.950 ;
        RECT 319.950 850.950 322.050 853.050 ;
        RECT 320.400 847.050 321.600 850.950 ;
        RECT 344.400 847.050 345.600 853.950 ;
        RECT 421.950 850.950 424.050 853.050 ;
        RECT 358.950 847.950 361.050 850.050 ;
        RECT 319.800 844.950 321.900 847.050 ;
        RECT 337.950 844.950 340.050 847.050 ;
        RECT 343.950 844.950 346.050 847.050 ;
        RECT 328.800 840.000 330.900 841.050 ;
        RECT 328.800 838.950 331.050 840.000 ;
        RECT 328.950 835.950 331.050 838.950 ;
        RECT 338.400 835.050 339.600 844.950 ;
        RECT 344.400 841.050 345.600 844.950 ;
        RECT 351.000 843.600 355.050 844.050 ;
        RECT 350.400 841.950 355.050 843.600 ;
        RECT 343.800 838.950 345.900 841.050 ;
        RECT 350.400 838.050 351.600 841.950 ;
        RECT 359.400 841.050 360.600 847.950 ;
        RECT 422.400 847.050 423.600 850.950 ;
        RECT 433.950 849.600 438.000 850.050 ;
        RECT 433.950 847.950 438.600 849.600 ;
        RECT 364.800 846.600 366.900 847.050 ;
        RECT 373.950 846.600 376.050 847.050 ;
        RECT 364.800 845.400 376.050 846.600 ;
        RECT 364.800 844.950 366.900 845.400 ;
        RECT 373.950 844.950 376.050 845.400 ;
        RECT 406.950 844.950 409.050 847.050 ;
        RECT 418.950 845.400 423.600 847.050 ;
        RECT 429.000 846.600 433.050 847.050 ;
        RECT 418.950 844.950 423.000 845.400 ;
        RECT 428.400 844.950 433.050 846.600 ;
        RECT 376.950 841.950 379.050 844.050 ;
        RECT 403.950 841.950 406.050 844.050 ;
        RECT 358.950 838.950 361.050 841.050 ;
        RECT 364.950 838.950 367.050 841.050 ;
        RECT 349.950 835.950 352.050 838.050 ;
        RECT 337.950 832.950 340.050 835.050 ;
        RECT 311.100 814.950 313.200 817.050 ;
        RECT 316.950 814.950 319.050 817.050 ;
        RECT 278.400 812.400 279.600 813.000 ;
        RECT 289.950 811.950 292.050 814.050 ;
        RECT 307.800 811.950 309.900 814.050 ;
        RECT 295.950 810.600 300.000 811.050 ;
        RECT 295.950 808.950 300.600 810.600 ;
        RECT 274.950 805.950 277.050 808.050 ;
        RECT 299.400 805.050 300.600 808.950 ;
        RECT 232.950 802.950 235.050 805.050 ;
        RECT 298.950 802.950 301.050 805.050 ;
        RECT 223.950 790.950 226.050 793.050 ;
        RECT 214.950 784.950 217.050 787.050 ;
        RECT 193.950 775.950 196.050 778.050 ;
        RECT 205.950 775.950 208.050 778.050 ;
        RECT 215.400 775.050 216.600 784.950 ;
        RECT 233.400 781.050 234.600 802.950 ;
        RECT 308.400 802.050 309.600 811.950 ;
        RECT 322.950 808.950 325.050 811.050 ;
        RECT 329.100 810.600 333.000 811.050 ;
        RECT 329.100 808.950 333.600 810.600 ;
        RECT 307.950 799.950 310.050 802.050 ;
        RECT 292.950 796.950 295.050 799.050 ;
        RECT 238.950 793.950 241.050 796.050 ;
        RECT 232.950 778.950 235.050 781.050 ;
        RECT 219.000 777.600 223.050 778.050 ;
        RECT 211.950 773.400 216.600 775.050 ;
        RECT 218.400 775.950 223.050 777.600 ;
        RECT 211.950 772.950 216.000 773.400 ;
        RECT 218.400 766.050 219.600 775.950 ;
        RECT 233.400 772.050 234.600 778.950 ;
        RECT 236.100 772.950 238.200 775.050 ;
        RECT 220.950 769.950 223.050 772.050 ;
        RECT 232.950 769.950 235.050 772.050 ;
        RECT 217.950 763.950 220.050 766.050 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 194.400 712.050 195.600 757.950 ;
        RECT 208.950 754.950 211.050 757.050 ;
        RECT 199.950 745.950 202.050 748.050 ;
        RECT 200.400 720.600 201.600 745.950 ;
        RECT 209.400 745.050 210.600 754.950 ;
        RECT 208.950 741.000 211.050 745.050 ;
        RECT 209.400 740.400 210.600 741.000 ;
        RECT 205.950 733.950 208.050 736.050 ;
        RECT 211.950 733.950 214.050 736.050 ;
        RECT 206.400 724.050 207.600 733.950 ;
        RECT 205.950 721.950 208.050 724.050 ;
        RECT 200.400 719.400 204.600 720.600 ;
        RECT 193.950 709.950 196.050 712.050 ;
        RECT 185.400 704.400 190.050 706.050 ;
        RECT 175.950 703.950 180.000 704.400 ;
        RECT 186.000 703.950 190.050 704.400 ;
        RECT 194.400 703.050 195.600 709.950 ;
        RECT 119.400 701.400 123.900 703.050 ;
        RECT 120.000 700.950 123.900 701.400 ;
        RECT 125.100 700.950 127.200 703.050 ;
        RECT 140.400 701.400 145.050 703.050 ;
        RECT 165.000 702.600 169.050 703.050 ;
        RECT 180.000 702.900 183.000 703.050 ;
        RECT 141.000 700.950 145.050 701.400 ;
        RECT 164.400 700.950 169.050 702.600 ;
        RECT 178.950 702.600 183.000 702.900 ;
        RECT 178.950 700.950 183.600 702.600 ;
        RECT 190.950 701.400 195.600 703.050 ;
        RECT 190.950 700.950 195.000 701.400 ;
        RECT 140.100 697.800 142.200 699.900 ;
        RECT 112.950 688.950 115.050 691.050 ;
        RECT 106.950 679.950 109.050 682.050 ;
        RECT 107.400 673.050 108.600 679.950 ;
        RECT 113.400 673.050 114.600 688.950 ;
        RECT 140.400 682.050 141.600 697.800 ;
        RECT 164.400 691.050 165.600 700.950 ;
        RECT 178.950 700.800 181.050 700.950 ;
        RECT 145.950 688.950 148.050 691.050 ;
        RECT 163.950 688.950 166.050 691.050 ;
        RECT 139.950 679.950 142.050 682.050 ;
        RECT 106.950 670.950 109.050 673.050 ;
        RECT 112.950 670.950 115.050 673.050 ;
        RECT 140.400 670.050 141.600 679.950 ;
        RECT 139.950 667.950 142.050 670.050 ;
        RECT 146.400 667.050 147.600 688.950 ;
        RECT 148.950 682.950 151.050 685.050 ;
        RECT 149.400 679.050 150.600 682.950 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 148.950 676.950 151.050 679.050 ;
        RECT 149.400 673.050 150.600 676.950 ;
        RECT 161.400 676.050 162.600 679.950 ;
        RECT 169.950 676.950 172.050 679.050 ;
        RECT 160.950 673.950 163.050 676.050 ;
        RECT 148.950 670.950 151.050 673.050 ;
        RECT 161.400 670.050 162.600 673.950 ;
        RECT 170.400 673.050 171.600 676.950 ;
        RECT 182.400 676.050 183.600 700.950 ;
        RECT 199.950 694.950 202.050 700.050 ;
        RECT 184.950 688.950 187.050 691.050 ;
        RECT 181.950 673.950 184.050 676.050 ;
        RECT 169.950 670.950 172.050 673.050 ;
        RECT 185.400 670.050 186.600 688.950 ;
        RECT 199.950 679.950 202.050 682.050 ;
        RECT 190.950 670.950 193.050 676.050 ;
        RECT 160.950 667.950 163.050 670.050 ;
        RECT 181.950 668.400 186.600 670.050 ;
        RECT 181.950 667.950 186.000 668.400 ;
        RECT 146.400 665.400 151.050 667.050 ;
        RECT 147.000 664.950 151.050 665.400 ;
        RECT 172.950 664.950 175.050 667.050 ;
        RECT 94.950 661.950 97.050 664.050 ;
        RECT 103.950 661.950 106.050 664.050 ;
        RECT 91.950 640.950 94.050 643.050 ;
        RECT 80.400 638.400 84.600 639.600 ;
        RECT 70.950 634.950 73.050 637.050 ;
        RECT 67.950 631.950 70.050 634.050 ;
        RECT 68.400 610.050 69.600 631.950 ;
        RECT 80.400 622.050 81.600 638.400 ;
        RECT 79.950 619.950 82.050 622.050 ;
        RECT 85.950 616.950 88.050 619.050 ;
        RECT 79.950 610.950 82.050 613.050 ;
        RECT 67.950 607.950 70.050 610.050 ;
        RECT 80.400 601.050 81.600 610.950 ;
        RECT 72.000 600.600 75.900 601.050 ;
        RECT 71.400 598.950 75.900 600.600 ;
        RECT 79.950 598.950 82.050 601.050 ;
        RECT 71.400 586.050 72.600 598.950 ;
        RECT 79.950 589.950 82.050 595.050 ;
        RECT 70.950 583.950 73.050 586.050 ;
        RECT 71.400 574.050 72.600 583.950 ;
        RECT 70.950 571.950 73.050 574.050 ;
        RECT 80.400 568.050 81.600 589.950 ;
        RECT 79.950 565.950 82.050 568.050 ;
        RECT 70.950 559.950 73.050 562.050 ;
        RECT 71.400 556.050 72.600 559.950 ;
        RECT 86.400 556.050 87.600 616.950 ;
        RECT 88.950 613.950 91.050 616.050 ;
        RECT 89.400 601.050 90.600 613.950 ;
        RECT 88.950 598.950 91.050 601.050 ;
        RECT 92.400 598.050 93.600 640.950 ;
        RECT 95.400 637.050 96.600 661.950 ;
        RECT 160.950 658.950 163.050 661.050 ;
        RECT 145.950 652.950 148.050 655.050 ;
        RECT 109.950 646.950 112.050 649.050 ;
        RECT 94.950 634.950 97.050 637.050 ;
        RECT 100.950 634.950 103.050 637.050 ;
        RECT 94.800 628.950 96.900 631.050 ;
        RECT 95.400 622.050 96.600 628.950 ;
        RECT 101.400 628.050 102.600 634.950 ;
        RECT 110.400 628.050 111.600 646.950 ;
        RECT 127.950 637.950 130.050 640.050 ;
        RECT 128.400 631.050 129.600 637.950 ;
        RECT 127.950 628.950 130.050 631.050 ;
        RECT 140.100 630.000 142.200 631.050 ;
        RECT 139.950 628.950 142.200 630.000 ;
        RECT 97.800 626.400 102.600 628.050 ;
        RECT 97.800 625.950 102.000 626.400 ;
        RECT 103.950 625.950 106.050 628.050 ;
        RECT 109.950 625.950 112.050 628.050 ;
        RECT 115.800 625.950 117.900 628.050 ;
        RECT 121.800 625.950 123.900 628.050 ;
        RECT 94.950 619.950 97.050 622.050 ;
        RECT 104.400 610.050 105.600 625.950 ;
        RECT 116.400 622.050 117.600 625.950 ;
        RECT 115.950 619.950 118.050 622.050 ;
        RECT 109.950 616.950 112.050 619.050 ;
        RECT 103.950 607.950 106.050 610.050 ;
        RECT 110.400 607.050 111.600 616.950 ;
        RECT 109.950 604.950 112.050 607.050 ;
        RECT 91.800 595.950 93.900 598.050 ;
        RECT 103.950 592.950 106.050 595.050 ;
        RECT 100.950 580.950 103.050 583.050 ;
        RECT 71.400 555.900 75.000 556.050 ;
        RECT 71.400 554.400 76.050 555.900 ;
        RECT 72.000 553.950 76.050 554.400 ;
        RECT 85.950 553.950 88.050 556.050 ;
        RECT 73.950 553.800 76.050 553.950 ;
        RECT 76.950 552.600 81.000 553.050 ;
        RECT 76.950 550.950 81.600 552.600 ;
        RECT 80.400 547.050 81.600 550.950 ;
        RECT 79.950 544.950 82.050 547.050 ;
        RECT 73.950 541.950 76.050 544.050 ;
        RECT 74.400 532.050 75.600 541.950 ;
        RECT 73.950 529.950 76.050 532.050 ;
        RECT 74.400 520.050 75.600 529.950 ;
        RECT 101.400 529.050 102.600 580.950 ;
        RECT 94.800 526.950 96.900 529.050 ;
        RECT 100.950 526.950 103.050 529.050 ;
        RECT 73.950 517.950 76.050 520.050 ;
        RECT 70.950 493.950 73.050 496.050 ;
        RECT 71.400 481.050 72.600 493.950 ;
        RECT 74.400 493.050 75.600 517.950 ;
        RECT 73.950 490.950 76.050 493.050 ;
        RECT 79.950 490.950 82.050 496.050 ;
        RECT 95.400 487.050 96.600 526.950 ;
        RECT 76.950 486.600 79.050 487.050 ;
        RECT 86.100 486.600 88.200 487.050 ;
        RECT 76.950 485.400 88.200 486.600 ;
        RECT 76.950 484.950 79.050 485.400 ;
        RECT 86.100 484.950 88.200 485.400 ;
        RECT 95.100 484.950 97.200 487.050 ;
        RECT 95.400 484.050 96.600 484.950 ;
        RECT 91.800 482.400 96.600 484.050 ;
        RECT 91.800 481.950 96.000 482.400 ;
        RECT 70.950 478.950 73.050 481.050 ;
        RECT 104.400 469.050 105.600 592.950 ;
        RECT 122.400 562.050 123.600 625.950 ;
        RECT 128.400 610.050 129.600 628.950 ;
        RECT 139.950 625.950 142.050 628.950 ;
        RECT 130.950 619.950 133.050 622.050 ;
        RECT 127.950 607.950 130.050 610.050 ;
        RECT 131.400 601.050 132.600 619.950 ;
        RECT 130.950 597.000 133.050 601.050 ;
        RECT 131.400 596.400 132.600 597.000 ;
        RECT 136.950 595.950 139.050 598.050 ;
        RECT 129.000 594.900 132.000 595.050 ;
        RECT 129.000 594.600 132.900 594.900 ;
        RECT 128.400 592.950 132.900 594.600 ;
        RECT 128.400 589.050 129.600 592.950 ;
        RECT 130.800 592.800 132.900 592.950 ;
        RECT 127.950 586.950 130.050 589.050 ;
        RECT 137.400 586.050 138.600 595.950 ;
        RECT 136.950 583.950 139.050 586.050 ;
        RECT 146.400 571.050 147.600 652.950 ;
        RECT 161.400 601.050 162.600 658.950 ;
        RECT 169.950 652.950 172.050 655.050 ;
        RECT 170.400 604.050 171.600 652.950 ;
        RECT 169.950 601.950 172.050 604.050 ;
        RECT 160.950 598.950 163.050 601.050 ;
        RECT 173.400 598.050 174.600 664.950 ;
        RECT 185.100 631.950 187.200 634.050 ;
        RECT 175.950 628.950 178.050 631.050 ;
        RECT 176.400 619.050 177.600 628.950 ;
        RECT 185.400 628.050 186.600 631.950 ;
        RECT 184.950 625.950 187.050 628.050 ;
        RECT 175.950 616.950 178.050 619.050 ;
        RECT 196.950 607.950 199.050 610.050 ;
        RECT 184.950 601.950 187.050 604.050 ;
        RECT 166.950 595.950 169.050 598.050 ;
        RECT 173.100 595.950 175.200 598.050 ;
        RECT 148.950 589.950 151.050 592.050 ;
        RECT 154.950 589.950 157.050 592.050 ;
        RECT 145.950 568.950 148.050 571.050 ;
        RECT 127.950 565.950 130.050 568.050 ;
        RECT 128.400 562.050 129.600 565.950 ;
        RECT 149.400 565.050 150.600 589.950 ;
        RECT 155.400 568.050 156.600 589.950 ;
        RECT 167.400 583.050 168.600 595.950 ;
        RECT 166.950 580.950 169.050 583.050 ;
        RECT 154.950 565.950 157.050 568.050 ;
        RECT 172.950 565.950 175.050 568.050 ;
        RECT 148.950 562.950 151.050 565.050 ;
        RECT 157.950 562.950 160.050 565.050 ;
        RECT 121.950 559.950 124.050 562.050 ;
        RECT 127.950 559.950 130.050 562.050 ;
        RECT 145.950 559.050 148.050 562.050 ;
        RECT 151.800 559.050 153.900 559.200 ;
        RECT 130.800 556.950 132.900 559.050 ;
        RECT 145.800 558.000 148.050 559.050 ;
        RECT 150.000 558.600 153.900 559.050 ;
        RECT 145.800 556.950 147.900 558.000 ;
        RECT 149.400 557.100 153.900 558.600 ;
        RECT 149.400 556.950 153.000 557.100 ;
        RECT 109.950 547.950 112.050 553.050 ;
        RECT 131.400 550.050 132.600 556.950 ;
        RECT 149.400 553.050 150.600 556.950 ;
        RECT 158.400 556.050 159.600 562.950 ;
        RECT 173.400 562.050 174.600 565.950 ;
        RECT 172.950 559.950 175.050 562.050 ;
        RECT 178.950 556.950 181.050 562.050 ;
        RECT 152.400 555.000 153.600 555.600 ;
        RECT 151.950 553.050 154.050 555.000 ;
        RECT 158.400 554.400 163.050 556.050 ;
        RECT 159.000 553.950 163.050 554.400 ;
        RECT 148.800 550.950 150.900 553.050 ;
        RECT 151.950 552.000 154.200 553.050 ;
        RECT 152.100 550.950 154.200 552.000 ;
        RECT 130.950 547.950 133.050 550.050 ;
        RECT 106.950 532.950 109.050 535.050 ;
        RECT 118.950 532.950 121.050 535.050 ;
        RECT 107.400 523.050 108.600 532.950 ;
        RECT 119.400 529.050 120.600 532.950 ;
        RECT 112.950 526.950 115.050 529.050 ;
        RECT 118.950 526.950 121.050 529.050 ;
        RECT 138.000 528.600 142.050 529.050 ;
        RECT 137.400 526.950 142.050 528.600 ;
        RECT 106.950 520.950 109.050 523.050 ;
        RECT 107.400 499.050 108.600 520.950 ;
        RECT 113.400 517.050 114.600 526.950 ;
        RECT 133.950 520.950 136.050 523.050 ;
        RECT 115.950 517.950 118.050 520.050 ;
        RECT 112.950 514.950 115.050 517.050 ;
        RECT 116.400 505.050 117.600 517.950 ;
        RECT 134.400 517.050 135.600 520.950 ;
        RECT 133.950 514.950 136.050 517.050 ;
        RECT 115.950 502.950 118.050 505.050 ;
        RECT 124.950 502.950 127.050 505.050 ;
        RECT 106.950 496.950 109.050 499.050 ;
        RECT 125.400 484.050 126.600 502.950 ;
        RECT 127.950 496.950 130.050 499.050 ;
        RECT 128.400 487.050 129.600 496.950 ;
        RECT 134.400 490.050 135.600 514.950 ;
        RECT 137.400 505.050 138.600 526.950 ;
        RECT 152.400 511.050 153.600 550.950 ;
        RECT 175.950 529.950 178.050 532.050 ;
        RECT 176.400 522.600 177.600 529.950 ;
        RECT 185.400 526.050 186.600 601.950 ;
        RECT 190.950 592.950 193.050 595.050 ;
        RECT 191.400 583.050 192.600 592.950 ;
        RECT 190.950 580.950 193.050 583.050 ;
        RECT 187.950 568.950 190.050 571.050 ;
        RECT 188.400 529.050 189.600 568.950 ;
        RECT 193.950 553.950 196.050 556.050 ;
        RECT 194.400 550.050 195.600 553.950 ;
        RECT 193.950 547.950 196.050 550.050 ;
        RECT 193.950 541.950 196.050 544.050 ;
        RECT 194.400 535.050 195.600 541.950 ;
        RECT 193.950 532.950 196.050 535.050 ;
        RECT 187.950 528.600 190.050 529.050 ;
        RECT 187.950 527.400 192.600 528.600 ;
        RECT 187.950 526.950 190.050 527.400 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 191.400 523.050 192.600 527.400 ;
        RECT 173.400 521.400 177.600 522.600 ;
        RECT 151.950 508.950 154.050 511.050 ;
        RECT 173.400 505.050 174.600 521.400 ;
        RECT 190.950 520.950 193.050 523.050 ;
        RECT 175.950 517.950 178.050 520.050 ;
        RECT 136.950 502.950 139.050 505.050 ;
        RECT 172.950 502.950 175.050 505.050 ;
        RECT 169.950 493.950 172.050 496.050 ;
        RECT 133.950 487.950 136.050 490.050 ;
        RECT 151.950 487.950 154.050 493.050 ;
        RECT 170.400 490.050 171.600 493.950 ;
        RECT 176.400 490.200 177.600 517.950 ;
        RECT 197.400 493.050 198.600 607.950 ;
        RECT 200.400 583.050 201.600 679.950 ;
        RECT 203.400 631.050 204.600 719.400 ;
        RECT 208.950 697.950 211.050 700.050 ;
        RECT 209.400 667.050 210.600 697.950 ;
        RECT 212.400 684.600 213.600 733.950 ;
        RECT 218.400 718.050 219.600 763.950 ;
        RECT 217.950 715.950 220.050 718.050 ;
        RECT 218.400 706.050 219.600 715.950 ;
        RECT 217.950 703.950 220.050 706.050 ;
        RECT 212.400 683.400 216.600 684.600 ;
        RECT 208.800 666.600 213.000 667.050 ;
        RECT 208.800 664.950 213.600 666.600 ;
        RECT 202.950 628.950 205.050 631.050 ;
        RECT 202.950 622.950 205.050 625.050 ;
        RECT 203.400 616.050 204.600 622.950 ;
        RECT 202.950 613.950 205.050 616.050 ;
        RECT 205.950 601.950 208.050 604.050 ;
        RECT 202.950 598.950 205.050 601.050 ;
        RECT 199.950 580.950 202.050 583.050 ;
        RECT 199.950 562.950 202.050 565.050 ;
        RECT 200.400 502.050 201.600 562.950 ;
        RECT 203.400 544.050 204.600 598.950 ;
        RECT 202.950 541.950 205.050 544.050 ;
        RECT 206.400 541.050 207.600 601.950 ;
        RECT 212.400 601.050 213.600 664.950 ;
        RECT 211.950 598.950 214.050 601.050 ;
        RECT 211.950 592.950 214.050 595.050 ;
        RECT 208.950 583.950 211.050 586.050 ;
        RECT 209.400 547.050 210.600 583.950 ;
        RECT 208.950 544.950 211.050 547.050 ;
        RECT 205.950 538.950 208.050 541.050 ;
        RECT 212.400 538.050 213.600 592.950 ;
        RECT 215.400 544.050 216.600 683.400 ;
        RECT 221.400 670.050 222.600 769.950 ;
        RECT 236.400 766.050 237.600 772.950 ;
        RECT 239.400 772.050 240.600 793.950 ;
        RECT 262.950 790.950 265.050 793.050 ;
        RECT 253.950 781.950 256.050 784.050 ;
        RECT 254.400 775.050 255.600 781.950 ;
        RECT 254.400 773.400 259.050 775.050 ;
        RECT 255.000 772.950 259.050 773.400 ;
        RECT 263.400 772.050 264.600 790.950 ;
        RECT 289.950 784.950 292.050 787.050 ;
        RECT 265.950 778.950 268.050 781.050 ;
        RECT 274.950 778.950 277.050 781.050 ;
        RECT 266.400 775.050 267.600 778.950 ;
        RECT 265.950 772.950 268.050 775.050 ;
        RECT 238.950 769.950 241.050 772.050 ;
        RECT 262.950 769.950 265.050 772.050 ;
        RECT 235.950 763.950 238.050 766.050 ;
        RECT 256.950 763.950 259.050 766.050 ;
        RECT 257.400 745.050 258.600 763.950 ;
        RECT 223.950 739.950 226.050 742.050 ;
        RECT 229.950 739.950 232.050 742.050 ;
        RECT 256.950 739.950 259.050 745.050 ;
        RECT 224.400 733.050 225.600 739.950 ;
        RECT 223.950 730.950 226.050 733.050 ;
        RECT 224.100 694.950 226.200 697.050 ;
        RECT 224.400 676.050 225.600 694.950 ;
        RECT 230.400 682.050 231.600 739.950 ;
        RECT 263.400 739.050 264.600 769.950 ;
        RECT 275.400 763.050 276.600 778.950 ;
        RECT 280.950 778.050 283.050 781.050 ;
        RECT 280.950 777.000 283.200 778.050 ;
        RECT 281.100 775.950 283.200 777.000 ;
        RECT 290.400 775.050 291.600 784.950 ;
        RECT 289.950 772.950 292.050 775.050 ;
        RECT 286.950 769.950 289.050 772.050 ;
        RECT 287.400 763.050 288.600 769.950 ;
        RECT 274.950 760.950 277.050 763.050 ;
        RECT 286.950 760.950 289.050 763.050 ;
        RECT 235.950 736.950 238.050 739.050 ;
        RECT 262.950 736.950 265.050 739.050 ;
        RECT 277.800 738.000 279.900 739.050 ;
        RECT 277.800 736.950 280.050 738.000 ;
        RECT 236.400 724.050 237.600 736.950 ;
        RECT 241.950 733.950 244.050 736.050 ;
        RECT 277.950 733.950 280.050 736.950 ;
        RECT 235.950 721.950 238.050 724.050 ;
        RECT 238.950 709.950 241.050 712.050 ;
        RECT 239.400 706.050 240.600 709.950 ;
        RECT 238.800 703.950 240.900 706.050 ;
        RECT 242.400 688.050 243.600 733.950 ;
        RECT 259.950 724.950 262.050 727.050 ;
        RECT 246.000 702.600 250.050 703.050 ;
        RECT 245.400 700.950 250.050 702.600 ;
        RECT 245.400 694.050 246.600 700.950 ;
        RECT 260.400 700.050 261.600 724.950 ;
        RECT 293.400 721.050 294.600 796.950 ;
        RECT 301.950 772.950 304.050 775.050 ;
        RECT 302.400 742.050 303.600 772.950 ;
        RECT 308.400 772.050 309.600 799.950 ;
        RECT 316.950 784.950 319.050 787.050 ;
        RECT 317.400 775.050 318.600 784.950 ;
        RECT 317.400 773.400 322.050 775.050 ;
        RECT 318.000 772.950 322.050 773.400 ;
        RECT 307.950 769.950 310.050 772.050 ;
        RECT 319.950 763.950 322.050 769.050 ;
        RECT 313.950 748.950 316.050 751.050 ;
        RECT 314.400 745.050 315.600 748.950 ;
        RECT 319.950 745.950 322.050 748.050 ;
        RECT 313.950 742.950 316.050 745.050 ;
        RECT 301.950 739.950 304.050 742.050 ;
        RECT 314.400 739.050 315.600 742.950 ;
        RECT 320.400 739.050 321.600 745.950 ;
        RECT 310.950 737.400 315.600 739.050 ;
        RECT 310.950 736.950 315.000 737.400 ;
        RECT 319.950 736.950 322.050 739.050 ;
        RECT 292.950 718.950 295.050 721.050 ;
        RECT 323.400 712.050 324.600 808.950 ;
        RECT 332.400 805.050 333.600 808.950 ;
        RECT 331.950 802.950 334.050 805.050 ;
        RECT 350.400 790.050 351.600 835.950 ;
        RECT 365.400 814.050 366.600 838.950 ;
        RECT 377.400 820.050 378.600 841.950 ;
        RECT 404.400 820.050 405.600 841.950 ;
        RECT 407.400 835.050 408.600 844.950 ;
        RECT 412.950 838.950 415.050 841.050 ;
        RECT 406.950 832.950 409.050 835.050 ;
        RECT 376.950 817.950 379.050 820.050 ;
        RECT 403.950 817.950 406.050 820.050 ;
        RECT 355.950 811.950 358.050 814.050 ;
        RECT 362.100 811.950 366.600 814.050 ;
        RECT 349.950 787.950 352.050 790.050 ;
        RECT 356.400 787.050 357.600 811.950 ;
        RECT 355.950 784.950 358.050 787.050 ;
        RECT 331.950 781.950 334.050 784.050 ;
        RECT 340.950 781.950 343.050 784.050 ;
        RECT 352.950 781.950 355.050 784.050 ;
        RECT 332.400 772.050 333.600 781.950 ;
        RECT 341.400 772.050 342.600 781.950 ;
        RECT 353.400 772.050 354.600 781.950 ;
        RECT 365.400 781.050 366.600 811.950 ;
        RECT 407.400 811.050 408.600 832.950 ;
        RECT 413.400 813.600 414.600 838.950 ;
        RECT 428.400 838.050 429.600 844.950 ;
        RECT 437.400 841.050 438.600 847.950 ;
        RECT 440.400 847.050 441.600 853.950 ;
        RECT 484.950 850.950 487.050 853.050 ;
        RECT 574.950 850.950 577.050 853.050 ;
        RECT 440.400 845.400 445.050 847.050 ;
        RECT 441.000 844.950 445.050 845.400 ;
        RECT 475.950 844.950 478.050 847.050 ;
        RECT 469.950 841.950 472.050 844.050 ;
        RECT 436.950 838.950 439.050 841.050 ;
        RECT 427.950 835.950 430.050 838.050 ;
        RECT 424.950 817.950 427.050 820.050 ;
        RECT 445.950 817.950 448.050 820.050 ;
        RECT 425.400 814.050 426.600 817.950 ;
        RECT 415.950 813.600 418.050 814.050 ;
        RECT 413.400 812.400 418.050 813.600 ;
        RECT 415.950 811.950 418.050 812.400 ;
        RECT 424.950 811.950 427.050 814.050 ;
        RECT 400.950 808.950 403.050 811.050 ;
        RECT 406.950 808.950 409.050 811.050 ;
        RECT 401.400 784.050 402.600 808.950 ;
        RECT 407.400 793.050 408.600 808.950 ;
        RECT 416.400 807.600 417.600 811.950 ;
        RECT 421.950 808.950 424.050 811.050 ;
        RECT 434.100 808.950 436.200 811.050 ;
        RECT 416.400 806.400 420.600 807.600 ;
        RECT 406.950 790.950 409.050 793.050 ;
        RECT 400.950 781.950 403.050 784.050 ;
        RECT 364.950 778.950 367.050 781.050 ;
        RECT 358.950 775.950 361.050 778.050 ;
        RECT 394.950 777.600 399.000 778.050 ;
        RECT 394.950 775.950 399.600 777.600 ;
        RECT 331.950 769.950 334.050 772.050 ;
        RECT 341.400 770.400 346.050 772.050 ;
        RECT 342.000 769.950 346.050 770.400 ;
        RECT 352.800 771.000 354.900 772.050 ;
        RECT 352.800 769.950 355.050 771.000 ;
        RECT 346.950 766.950 349.050 769.050 ;
        RECT 352.950 768.000 355.050 769.950 ;
        RECT 359.400 769.050 360.600 775.950 ;
        RECT 370.950 774.600 375.000 775.050 ;
        RECT 370.950 772.950 375.600 774.600 ;
        RECT 391.950 772.950 394.050 775.050 ;
        RECT 364.950 769.950 367.050 772.050 ;
        RECT 353.400 767.400 354.600 768.000 ;
        RECT 358.950 766.950 361.050 769.050 ;
        RECT 340.950 760.950 343.050 763.050 ;
        RECT 341.400 745.050 342.600 760.950 ;
        RECT 347.400 751.050 348.600 766.950 ;
        RECT 346.950 748.950 349.050 751.050 ;
        RECT 358.950 748.950 361.050 751.050 ;
        RECT 359.400 745.050 360.600 748.950 ;
        RECT 325.950 742.950 328.050 745.050 ;
        RECT 335.100 742.950 337.200 745.050 ;
        RECT 341.100 742.950 343.200 745.050 ;
        RECT 358.800 742.950 360.900 745.050 ;
        RECT 326.400 730.050 327.600 742.950 ;
        RECT 335.400 733.050 336.600 742.950 ;
        RECT 365.400 736.050 366.600 769.950 ;
        RECT 374.400 766.050 375.600 772.950 ;
        RECT 388.950 766.950 391.050 769.050 ;
        RECT 373.950 763.950 376.050 766.050 ;
        RECT 389.400 739.050 390.600 766.950 ;
        RECT 392.400 742.050 393.600 772.950 ;
        RECT 398.400 754.050 399.600 775.950 ;
        RECT 415.950 754.950 418.050 757.050 ;
        RECT 397.950 751.950 400.050 754.050 ;
        RECT 416.400 745.050 417.600 754.950 ;
        RECT 419.400 754.050 420.600 806.400 ;
        RECT 422.400 760.050 423.600 808.950 ;
        RECT 434.400 799.050 435.600 808.950 ;
        RECT 446.400 808.050 447.600 817.950 ;
        RECT 466.950 811.950 469.050 814.050 ;
        RECT 445.950 805.950 448.050 808.050 ;
        RECT 460.950 802.950 463.050 805.050 ;
        RECT 433.950 796.950 436.050 799.050 ;
        RECT 454.950 790.950 457.050 793.050 ;
        RECT 448.950 784.950 451.050 787.050 ;
        RECT 430.950 778.950 433.050 784.050 ;
        RECT 449.400 778.050 450.600 784.950 ;
        RECT 446.100 776.400 450.600 778.050 ;
        RECT 446.100 775.950 450.000 776.400 ;
        RECT 455.400 775.050 456.600 790.950 ;
        RECT 454.950 772.950 457.050 775.050 ;
        RECT 442.950 769.950 445.050 772.050 ;
        RECT 421.950 757.950 424.050 760.050 ;
        RECT 418.950 751.950 421.050 754.050 ;
        RECT 433.950 751.950 436.050 754.050 ;
        RECT 418.950 745.950 421.050 748.050 ;
        RECT 397.800 742.950 399.900 745.050 ;
        RECT 403.800 742.950 405.900 745.050 ;
        RECT 415.950 744.600 418.050 745.050 ;
        RECT 413.400 743.400 418.050 744.600 ;
        RECT 391.950 739.950 394.050 742.050 ;
        RECT 388.950 736.950 391.050 739.050 ;
        RECT 355.950 733.950 358.050 736.050 ;
        RECT 364.950 733.950 367.050 736.050 ;
        RECT 334.950 730.950 337.050 733.050 ;
        RECT 325.950 727.950 328.050 730.050 ;
        RECT 328.950 718.950 331.050 721.050 ;
        RECT 292.950 709.950 295.050 712.050 ;
        RECT 322.950 709.950 325.050 712.050 ;
        RECT 268.950 703.950 271.050 706.050 ;
        RECT 256.800 699.000 258.900 700.050 ;
        RECT 256.800 697.950 259.050 699.000 ;
        RECT 260.400 698.400 264.900 700.050 ;
        RECT 261.000 697.950 264.900 698.400 ;
        RECT 256.950 694.950 259.050 697.950 ;
        RECT 244.950 691.950 247.050 694.050 ;
        RECT 262.950 691.950 265.050 694.050 ;
        RECT 247.950 688.950 250.050 691.050 ;
        RECT 241.950 685.950 244.050 688.050 ;
        RECT 244.950 682.950 247.050 685.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 223.950 673.950 226.050 676.050 ;
        RECT 232.950 673.950 235.050 676.050 ;
        RECT 220.800 667.950 222.900 670.050 ;
        RECT 217.950 664.950 220.050 667.050 ;
        RECT 218.400 598.050 219.600 664.950 ;
        RECT 229.950 640.950 232.050 643.050 ;
        RECT 223.950 630.600 228.000 631.050 ;
        RECT 223.950 628.950 228.600 630.600 ;
        RECT 227.400 619.050 228.600 628.950 ;
        RECT 226.950 616.950 229.050 619.050 ;
        RECT 230.400 601.050 231.600 640.950 ;
        RECT 230.100 598.950 232.200 601.050 ;
        RECT 233.400 598.050 234.600 673.950 ;
        RECT 241.950 667.950 244.050 670.050 ;
        RECT 235.950 646.950 238.050 649.050 ;
        RECT 236.400 631.050 237.600 646.950 ;
        RECT 235.950 628.950 238.050 631.050 ;
        RECT 236.400 625.050 237.600 628.950 ;
        RECT 238.950 625.950 241.050 628.050 ;
        RECT 235.950 622.950 238.050 625.050 ;
        RECT 239.400 616.050 240.600 625.950 ;
        RECT 242.400 625.200 243.600 667.950 ;
        RECT 241.950 623.100 244.050 625.200 ;
        RECT 241.950 619.800 244.050 621.900 ;
        RECT 238.950 613.950 241.050 616.050 ;
        RECT 236.100 600.000 238.200 601.050 ;
        RECT 235.950 598.950 238.200 600.000 ;
        RECT 235.950 598.050 238.050 598.950 ;
        RECT 218.400 596.400 223.050 598.050 ;
        RECT 219.000 595.950 223.050 596.400 ;
        RECT 232.800 597.000 238.050 598.050 ;
        RECT 232.800 596.400 237.600 597.000 ;
        RECT 232.800 595.950 237.000 596.400 ;
        RECT 229.950 592.950 232.050 595.050 ;
        RECT 238.950 592.950 241.050 595.050 ;
        RECT 226.950 583.950 229.050 586.050 ;
        RECT 217.950 580.950 220.050 583.050 ;
        RECT 218.400 556.050 219.600 580.950 ;
        RECT 227.400 562.050 228.600 583.950 ;
        RECT 226.950 559.950 229.050 562.050 ;
        RECT 217.950 553.950 220.050 556.050 ;
        RECT 214.950 541.950 217.050 544.050 ;
        RECT 220.950 541.950 223.050 544.050 ;
        RECT 217.950 538.950 220.050 541.050 ;
        RECT 211.950 535.950 214.050 538.050 ;
        RECT 205.950 526.950 208.050 529.050 ;
        RECT 202.950 523.950 205.050 526.050 ;
        RECT 203.400 517.050 204.600 523.950 ;
        RECT 202.950 514.950 205.050 517.050 ;
        RECT 199.950 499.950 202.050 502.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 169.800 487.950 171.900 490.050 ;
        RECT 175.950 488.100 178.050 490.200 ;
        RECT 127.950 484.950 130.050 487.050 ;
        RECT 124.950 481.950 127.050 484.050 ;
        RECT 134.400 481.050 135.600 487.950 ;
        RECT 163.950 484.950 166.050 487.050 ;
        RECT 177.000 486.600 181.050 487.050 ;
        RECT 176.400 484.950 181.050 486.600 ;
        RECT 190.950 486.600 195.000 487.050 ;
        RECT 190.950 484.950 195.600 486.600 ;
        RECT 158.100 481.950 160.200 484.050 ;
        RECT 127.950 478.950 130.050 481.050 ;
        RECT 133.950 478.950 136.050 481.050 ;
        RECT 103.950 466.950 106.050 469.050 ;
        RECT 115.950 466.950 118.050 469.050 ;
        RECT 91.950 460.950 94.050 463.050 ;
        RECT 79.950 457.050 82.050 460.050 ;
        RECT 64.950 454.950 67.050 457.050 ;
        RECT 73.950 454.950 76.050 457.050 ;
        RECT 79.950 456.000 82.200 457.050 ;
        RECT 80.100 454.950 82.200 456.000 ;
        RECT 70.950 451.950 73.050 454.050 ;
        RECT 55.950 442.950 58.050 445.050 ;
        RECT 71.400 439.050 72.600 451.950 ;
        RECT 74.400 448.050 75.600 454.950 ;
        RECT 92.400 454.050 93.600 460.950 ;
        RECT 100.950 457.950 103.050 460.050 ;
        RECT 101.400 454.050 102.600 457.950 ;
        RECT 116.400 457.050 117.600 466.950 ;
        RECT 115.950 454.950 118.050 457.050 ;
        RECT 91.950 451.950 94.050 454.050 ;
        RECT 100.950 451.950 103.050 454.050 ;
        RECT 124.950 451.950 127.050 454.050 ;
        RECT 73.950 445.950 76.050 448.050 ;
        RECT 70.950 436.950 73.050 439.050 ;
        RECT 74.400 436.050 75.600 445.950 ;
        RECT 92.400 445.050 93.600 451.950 ;
        RECT 97.950 445.950 100.050 448.050 ;
        RECT 91.950 442.950 94.050 445.050 ;
        RECT 85.950 439.950 88.050 442.050 ;
        RECT 73.950 433.950 76.050 436.050 ;
        RECT 79.950 421.950 82.050 424.050 ;
        RECT 55.950 418.950 58.050 421.050 ;
        RECT 56.400 412.050 57.600 418.950 ;
        RECT 73.950 415.950 76.050 421.050 ;
        RECT 80.400 418.050 81.600 421.950 ;
        RECT 79.950 415.950 82.050 418.050 ;
        RECT 58.800 414.600 63.000 415.050 ;
        RECT 58.800 412.950 63.600 414.600 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 62.400 412.050 63.600 412.950 ;
        RECT 55.950 409.950 58.050 412.050 ;
        RECT 62.400 410.400 67.050 412.050 ;
        RECT 63.000 409.950 67.050 410.400 ;
        RECT 68.400 406.050 69.600 412.950 ;
        RECT 67.950 403.950 70.050 406.050 ;
        RECT 64.950 391.950 67.050 394.050 ;
        RECT 50.100 385.950 52.200 388.050 ;
        RECT 46.800 382.950 48.900 385.050 ;
        RECT 50.400 382.050 51.600 385.950 ;
        RECT 58.950 382.950 61.050 385.050 ;
        RECT 49.950 379.950 52.050 382.050 ;
        RECT 46.950 370.950 49.050 373.050 ;
        RECT 47.400 343.200 48.600 370.950 ;
        RECT 46.950 341.100 49.050 343.200 ;
        RECT 50.400 340.050 51.600 379.950 ;
        RECT 59.400 376.050 60.600 382.950 ;
        RECT 65.400 382.050 66.600 391.950 ;
        RECT 74.400 391.050 75.600 415.950 ;
        RECT 82.950 406.950 85.050 409.050 ;
        RECT 73.950 388.950 76.050 391.050 ;
        RECT 83.400 390.600 84.600 406.950 ;
        RECT 86.400 394.050 87.600 439.950 ;
        RECT 88.950 433.950 91.050 436.050 ;
        RECT 89.400 415.050 90.600 433.950 ;
        RECT 88.950 412.950 91.050 415.050 ;
        RECT 98.400 412.050 99.600 445.950 ;
        RECT 125.400 445.050 126.600 451.950 ;
        RECT 124.950 442.950 127.050 445.050 ;
        RECT 124.950 427.950 127.050 430.050 ;
        RECT 118.950 421.950 121.050 424.050 ;
        RECT 97.950 409.950 100.050 412.050 ;
        RECT 109.950 411.600 114.000 412.050 ;
        RECT 109.950 409.950 114.600 411.600 ;
        RECT 94.950 394.950 97.050 397.050 ;
        RECT 106.950 394.950 109.050 397.050 ;
        RECT 85.950 391.950 88.050 394.050 ;
        RECT 80.400 389.400 84.600 390.600 ;
        RECT 70.950 384.600 75.000 385.050 ;
        RECT 70.950 382.950 75.600 384.600 ;
        RECT 64.950 379.950 67.050 382.050 ;
        RECT 58.950 373.950 61.050 376.050 ;
        RECT 74.400 373.050 75.600 382.950 ;
        RECT 73.950 370.950 76.050 373.050 ;
        RECT 73.950 361.950 76.050 364.050 ;
        RECT 67.950 358.950 70.050 361.050 ;
        RECT 64.950 352.950 67.050 355.050 ;
        RECT 55.800 340.950 57.900 343.050 ;
        RECT 48.000 339.900 51.600 340.050 ;
        RECT 46.950 338.250 51.600 339.900 ;
        RECT 46.950 337.950 51.000 338.250 ;
        RECT 46.950 337.800 49.050 337.950 ;
        RECT 46.950 328.950 49.050 331.050 ;
        RECT 34.950 310.950 37.050 313.050 ;
        RECT 40.950 310.950 43.050 313.050 ;
        RECT 43.950 307.950 46.050 310.050 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 28.950 271.950 31.050 274.050 ;
        RECT 16.800 270.600 21.000 271.050 ;
        RECT 16.800 270.000 21.600 270.600 ;
        RECT 16.800 268.950 22.050 270.000 ;
        RECT 23.100 268.950 25.200 271.050 ;
        RECT 19.950 268.050 22.050 268.950 ;
        RECT 13.800 265.950 15.900 268.050 ;
        RECT 19.950 267.000 22.200 268.050 ;
        RECT 20.100 265.950 22.200 267.000 ;
        RECT 28.950 265.950 31.050 268.050 ;
        RECT 10.950 262.950 13.050 265.050 ;
        RECT 29.400 250.050 30.600 265.950 ;
        RECT 28.950 247.950 31.050 250.050 ;
        RECT 16.950 244.950 19.050 247.050 ;
        RECT 4.950 238.950 7.050 241.050 ;
        RECT 17.400 238.050 18.600 244.950 ;
        RECT 35.400 241.050 36.600 289.950 ;
        RECT 44.400 280.050 45.600 307.950 ;
        RECT 43.950 277.950 46.050 280.050 ;
        RECT 44.400 274.050 45.600 277.950 ;
        RECT 43.950 271.950 46.050 274.050 ;
        RECT 47.400 244.050 48.600 328.950 ;
        RECT 56.400 319.050 57.600 340.950 ;
        RECT 65.400 322.050 66.600 352.950 ;
        RECT 64.950 319.950 67.050 322.050 ;
        RECT 55.950 316.950 58.050 319.050 ;
        RECT 61.950 316.950 64.050 319.050 ;
        RECT 62.400 313.200 63.600 316.950 ;
        RECT 61.950 311.100 64.050 313.200 ;
        RECT 68.400 313.050 69.600 358.950 ;
        RECT 74.400 346.200 75.600 361.950 ;
        RECT 80.400 358.050 81.600 389.400 ;
        RECT 95.400 385.050 96.600 394.950 ;
        RECT 85.950 382.950 88.050 385.050 ;
        RECT 94.950 382.950 97.050 385.050 ;
        RECT 82.950 376.950 85.050 379.050 ;
        RECT 79.950 355.950 82.050 358.050 ;
        RECT 83.400 355.050 84.600 376.950 ;
        RECT 82.950 352.950 85.050 355.050 ;
        RECT 86.400 352.050 87.600 382.950 ;
        RECT 107.400 379.050 108.600 394.950 ;
        RECT 100.950 373.950 103.050 379.050 ;
        RECT 106.950 376.950 109.050 379.050 ;
        RECT 97.950 358.950 100.050 361.050 ;
        RECT 76.950 349.950 79.050 352.050 ;
        RECT 85.950 349.950 88.050 352.050 ;
        RECT 73.950 344.100 76.050 346.200 ;
        RECT 77.400 343.050 78.600 349.950 ;
        RECT 91.950 346.950 94.050 349.050 ;
        RECT 92.400 343.050 93.600 346.950 ;
        RECT 98.400 343.200 99.600 358.950 ;
        RECT 103.950 355.950 106.050 358.050 ;
        RECT 75.000 342.900 78.600 343.050 ;
        RECT 73.950 341.250 78.600 342.900 ;
        RECT 73.950 340.950 78.000 341.250 ;
        RECT 91.950 340.950 94.050 343.050 ;
        RECT 98.100 341.100 100.200 343.200 ;
        RECT 104.400 343.050 105.600 355.950 ;
        RECT 107.400 346.050 108.600 376.950 ;
        RECT 113.400 373.050 114.600 409.950 ;
        RECT 119.400 394.050 120.600 421.950 ;
        RECT 125.400 397.050 126.600 427.950 ;
        RECT 124.950 394.950 127.050 397.050 ;
        RECT 118.950 391.950 121.050 394.050 ;
        RECT 119.400 388.050 120.600 391.950 ;
        RECT 128.400 391.050 129.600 478.950 ;
        RECT 158.400 469.050 159.600 481.950 ;
        RECT 164.400 475.050 165.600 484.950 ;
        RECT 166.950 475.950 169.050 478.050 ;
        RECT 163.950 472.950 166.050 475.050 ;
        RECT 139.950 466.950 142.050 469.050 ;
        RECT 157.950 466.950 160.050 469.050 ;
        RECT 134.100 454.950 136.200 457.050 ;
        RECT 131.100 451.950 133.200 454.050 ;
        RECT 131.400 448.050 132.600 451.950 ;
        RECT 130.950 445.950 133.050 448.050 ;
        RECT 131.400 427.050 132.600 445.950 ;
        RECT 130.950 424.950 133.050 427.050 ;
        RECT 134.400 412.050 135.600 454.950 ;
        RECT 140.400 430.050 141.600 466.950 ;
        RECT 148.950 457.950 151.050 460.050 ;
        RECT 155.100 457.950 157.200 460.050 ;
        RECT 145.950 454.950 148.050 457.050 ;
        RECT 146.400 451.050 147.600 454.950 ;
        RECT 145.950 448.950 148.050 451.050 ;
        RECT 149.400 439.050 150.600 457.950 ;
        RECT 155.400 454.050 156.600 457.950 ;
        RECT 167.400 457.050 168.600 475.950 ;
        RECT 176.400 469.050 177.600 484.950 ;
        RECT 191.400 478.050 192.600 484.950 ;
        RECT 194.400 481.050 195.600 484.950 ;
        RECT 193.950 478.950 196.050 481.050 ;
        RECT 202.950 478.950 205.050 481.050 ;
        RECT 190.950 475.950 193.050 478.050 ;
        RECT 178.950 472.950 181.050 475.050 ;
        RECT 175.950 466.950 178.050 469.050 ;
        RECT 166.950 454.950 169.050 457.050 ;
        RECT 154.950 451.950 157.050 454.050 ;
        RECT 160.950 448.950 163.050 451.050 ;
        RECT 148.950 436.950 151.050 439.050 ;
        RECT 149.400 430.050 150.600 436.950 ;
        RECT 161.400 430.050 162.600 448.950 ;
        RECT 139.800 427.950 141.900 430.050 ;
        RECT 143.100 427.950 145.200 430.050 ;
        RECT 148.950 427.950 151.050 430.050 ;
        RECT 160.950 427.950 163.050 430.050 ;
        RECT 169.950 427.950 172.050 430.050 ;
        RECT 136.950 424.950 139.050 427.050 ;
        RECT 137.400 415.050 138.600 424.950 ;
        RECT 143.400 418.050 144.600 427.950 ;
        RECT 157.950 421.950 160.050 424.050 ;
        RECT 142.800 415.950 144.900 418.050 ;
        RECT 158.400 415.050 159.600 421.950 ;
        RECT 166.950 418.950 169.050 421.050 ;
        RECT 137.400 413.400 142.050 415.050 ;
        RECT 138.000 412.950 142.050 413.400 ;
        RECT 145.950 412.950 148.050 415.050 ;
        RECT 158.100 412.950 160.200 415.050 ;
        RECT 130.800 410.400 135.600 412.050 ;
        RECT 130.800 409.950 135.000 410.400 ;
        RECT 146.400 394.050 147.600 412.950 ;
        RECT 167.400 409.050 168.600 418.950 ;
        RECT 151.800 406.950 153.900 409.050 ;
        RECT 155.100 406.950 157.200 409.050 ;
        RECT 166.950 406.950 169.050 409.050 ;
        RECT 152.400 397.050 153.600 406.950 ;
        RECT 151.950 394.950 154.050 397.050 ;
        RECT 145.950 391.950 148.050 394.050 ;
        RECT 127.950 388.950 130.050 391.050 ;
        RECT 118.950 385.950 121.050 388.050 ;
        RECT 139.950 385.950 142.050 388.050 ;
        RECT 119.400 379.050 120.600 385.950 ;
        RECT 140.400 381.600 141.600 385.950 ;
        RECT 137.400 380.400 141.600 381.600 ;
        RECT 118.950 376.950 121.050 379.050 ;
        RECT 124.950 376.950 127.050 379.050 ;
        RECT 133.950 376.950 136.050 379.050 ;
        RECT 112.950 370.950 115.050 373.050 ;
        RECT 115.950 364.950 118.050 367.050 ;
        RECT 116.400 349.050 117.600 364.950 ;
        RECT 125.400 364.050 126.600 376.950 ;
        RECT 134.400 373.050 135.600 376.950 ;
        RECT 137.400 376.050 138.600 380.400 ;
        RECT 152.400 379.050 153.600 394.950 ;
        RECT 155.400 385.050 156.600 406.950 ;
        RECT 154.950 382.950 157.050 385.050 ;
        RECT 170.400 382.050 171.600 427.950 ;
        RECT 179.400 394.050 180.600 472.950 ;
        RECT 193.950 466.950 196.050 469.050 ;
        RECT 181.950 451.950 184.050 454.050 ;
        RECT 182.400 421.050 183.600 451.950 ;
        RECT 187.950 448.950 190.050 451.050 ;
        RECT 188.400 442.050 189.600 448.950 ;
        RECT 187.950 439.950 190.050 442.050 ;
        RECT 190.950 424.950 193.050 427.050 ;
        RECT 181.950 418.950 184.050 421.050 ;
        RECT 191.400 415.050 192.600 424.950 ;
        RECT 184.800 412.950 186.900 415.050 ;
        RECT 190.950 412.950 193.050 415.050 ;
        RECT 178.950 391.950 181.050 394.050 ;
        RECT 172.800 382.950 174.900 385.050 ;
        RECT 169.950 379.950 172.050 382.050 ;
        RECT 151.950 376.950 154.050 379.050 ;
        RECT 136.950 373.950 139.050 376.050 ;
        RECT 154.950 373.950 157.050 376.050 ;
        RECT 133.950 370.950 136.050 373.050 ;
        RECT 130.950 364.950 133.050 367.050 ;
        RECT 124.950 361.950 127.050 364.050 ;
        RECT 118.950 352.950 121.050 355.050 ;
        RECT 119.400 349.050 120.600 352.950 ;
        RECT 127.950 349.950 130.050 352.050 ;
        RECT 115.800 346.950 117.900 349.050 ;
        RECT 119.100 346.950 121.200 349.050 ;
        RECT 106.950 343.950 109.050 346.050 ;
        RECT 104.100 340.950 106.200 343.050 ;
        RECT 73.950 340.800 76.050 340.950 ;
        RECT 128.400 340.050 129.600 349.950 ;
        RECT 99.000 339.600 102.900 340.050 ;
        RECT 98.400 337.950 102.900 339.600 ;
        RECT 127.950 337.950 130.050 340.050 ;
        RECT 67.950 310.950 70.050 313.050 ;
        RECT 85.950 310.950 88.050 313.050 ;
        RECT 59.100 309.600 63.000 310.050 ;
        RECT 59.100 307.950 63.600 309.600 ;
        RECT 55.950 292.950 58.050 295.050 ;
        RECT 49.950 286.950 52.050 289.050 ;
        RECT 50.400 277.050 51.600 286.950 ;
        RECT 49.950 274.950 52.050 277.050 ;
        RECT 50.400 271.050 51.600 274.950 ;
        RECT 49.800 268.950 51.900 271.050 ;
        RECT 56.400 259.050 57.600 292.950 ;
        RECT 62.400 286.050 63.600 307.950 ;
        RECT 70.950 304.950 73.050 307.050 ;
        RECT 79.950 304.950 82.050 307.050 ;
        RECT 61.950 283.950 64.050 286.050 ;
        RECT 71.400 283.050 72.600 304.950 ;
        RECT 80.400 289.050 81.600 304.950 ;
        RECT 86.400 301.050 87.600 310.950 ;
        RECT 85.950 300.600 88.050 301.050 ;
        RECT 85.950 299.400 90.600 300.600 ;
        RECT 85.950 298.950 88.050 299.400 ;
        RECT 82.950 292.950 85.050 295.050 ;
        RECT 79.950 286.950 82.050 289.050 ;
        RECT 70.950 280.950 73.050 283.050 ;
        RECT 73.950 277.950 76.050 280.050 ;
        RECT 70.950 274.950 73.050 277.050 ;
        RECT 61.950 268.950 64.050 271.050 ;
        RECT 62.400 262.050 63.600 268.950 ;
        RECT 71.400 265.050 72.600 274.950 ;
        RECT 74.400 274.050 75.600 277.950 ;
        RECT 73.950 271.950 76.050 274.050 ;
        RECT 77.400 267.000 78.600 267.600 ;
        RECT 70.950 262.950 73.050 265.050 ;
        RECT 76.950 262.950 79.050 267.000 ;
        RECT 61.950 259.950 64.050 262.050 ;
        RECT 55.950 256.950 58.050 259.050 ;
        RECT 61.950 253.950 64.050 256.050 ;
        RECT 52.950 250.950 55.050 253.050 ;
        RECT 46.950 241.950 49.050 244.050 ;
        RECT 53.400 241.050 54.600 250.950 ;
        RECT 28.950 238.950 31.050 241.050 ;
        RECT 34.800 238.950 36.900 241.050 ;
        RECT 52.950 238.950 55.050 241.050 ;
        RECT 17.400 236.400 22.050 238.050 ;
        RECT 18.000 235.950 22.050 236.400 ;
        RECT 10.950 232.950 13.050 235.050 ;
        RECT 11.400 226.050 12.600 232.950 ;
        RECT 16.950 232.800 19.050 234.900 ;
        RECT 10.950 223.950 13.050 226.050 ;
        RECT 17.400 196.050 18.600 232.800 ;
        RECT 20.400 196.050 21.600 235.950 ;
        RECT 29.400 202.050 30.600 238.950 ;
        RECT 49.950 235.950 52.050 238.050 ;
        RECT 46.950 223.950 49.050 226.050 ;
        RECT 34.950 205.950 37.050 208.050 ;
        RECT 28.800 199.950 30.900 202.050 ;
        RECT 35.400 199.050 36.600 205.950 ;
        RECT 47.400 205.050 48.600 223.950 ;
        RECT 50.400 205.050 51.600 235.950 ;
        RECT 46.800 202.950 48.900 205.050 ;
        RECT 50.100 202.950 52.200 205.050 ;
        RECT 40.950 199.950 43.050 202.050 ;
        RECT 35.400 197.400 40.050 199.050 ;
        RECT 36.000 196.950 40.050 197.400 ;
        RECT 14.400 195.000 15.600 195.600 ;
        RECT 13.950 190.950 16.050 195.000 ;
        RECT 16.800 193.950 18.900 196.050 ;
        RECT 20.400 193.950 25.050 196.050 ;
        RECT 4.950 184.950 7.050 187.050 ;
        RECT 5.400 166.050 6.600 184.950 ;
        RECT 14.400 181.050 15.600 190.950 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 17.400 178.050 18.600 193.950 ;
        RECT 16.950 175.950 19.050 178.050 ;
        RECT 13.950 172.950 16.050 175.050 ;
        RECT 14.400 172.050 15.600 172.950 ;
        RECT 20.400 172.050 21.600 193.950 ;
        RECT 31.950 187.950 34.050 190.050 ;
        RECT 25.950 172.950 28.050 175.050 ;
        RECT 13.950 168.000 16.050 172.050 ;
        RECT 19.950 169.950 22.050 172.050 ;
        RECT 14.400 167.400 15.600 168.000 ;
        RECT 26.400 166.050 27.600 172.950 ;
        RECT 4.950 163.950 7.050 166.050 ;
        RECT 25.950 163.950 28.050 166.050 ;
        RECT 32.400 163.050 33.600 187.950 ;
        RECT 41.400 169.050 42.600 199.950 ;
        RECT 47.400 199.050 48.600 202.950 ;
        RECT 53.400 199.050 54.600 238.950 ;
        RECT 62.400 238.050 63.600 253.950 ;
        RECT 77.400 252.600 78.600 262.950 ;
        RECT 83.400 253.050 84.600 292.950 ;
        RECT 85.950 286.950 88.050 289.050 ;
        RECT 86.400 256.050 87.600 286.950 ;
        RECT 89.400 271.050 90.600 299.400 ;
        RECT 98.400 289.050 99.600 337.950 ;
        RECT 124.950 334.950 127.050 337.050 ;
        RECT 118.950 331.950 121.050 334.050 ;
        RECT 112.950 328.950 115.050 331.050 ;
        RECT 106.950 316.950 109.050 319.050 ;
        RECT 101.100 307.950 103.200 310.050 ;
        RECT 101.400 292.050 102.600 307.950 ;
        RECT 107.400 292.050 108.600 316.950 ;
        RECT 113.400 307.050 114.600 328.950 ;
        RECT 119.400 316.050 120.600 331.950 ;
        RECT 118.950 313.950 121.050 316.050 ;
        RECT 109.950 305.400 114.600 307.050 ;
        RECT 119.400 307.050 120.600 313.950 ;
        RECT 119.400 305.400 124.050 307.050 ;
        RECT 109.950 304.950 114.000 305.400 ;
        RECT 120.000 304.950 124.050 305.400 ;
        RECT 100.950 289.950 103.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 97.950 286.950 100.050 289.050 ;
        RECT 103.950 286.950 106.050 289.050 ;
        RECT 109.950 286.950 112.050 289.050 ;
        RECT 94.950 283.950 97.050 286.050 ;
        RECT 95.400 274.050 96.600 283.950 ;
        RECT 97.950 280.950 100.050 283.050 ;
        RECT 91.950 272.400 96.600 274.050 ;
        RECT 91.950 271.950 96.000 272.400 ;
        RECT 98.400 271.050 99.600 280.950 ;
        RECT 104.400 274.050 105.600 286.950 ;
        RECT 103.950 271.950 106.050 274.050 ;
        RECT 88.950 268.950 91.050 271.050 ;
        RECT 98.400 269.400 103.050 271.050 ;
        RECT 99.000 268.950 103.050 269.400 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 85.950 253.950 88.050 256.050 ;
        RECT 77.400 252.000 81.600 252.600 ;
        RECT 77.400 251.400 82.050 252.000 ;
        RECT 79.950 247.950 82.050 251.400 ;
        RECT 82.950 250.950 85.050 253.050 ;
        RECT 97.950 244.950 100.050 247.050 ;
        RECT 70.950 238.950 73.050 244.050 ;
        RECT 98.400 241.050 99.600 244.950 ;
        RECT 85.950 238.950 88.050 241.050 ;
        RECT 97.950 238.950 100.050 241.050 ;
        RECT 56.400 237.000 60.600 237.600 ;
        RECT 55.950 236.400 60.600 237.000 ;
        RECT 62.400 236.400 67.050 238.050 ;
        RECT 55.950 232.950 58.050 236.400 ;
        RECT 59.400 232.050 60.600 236.400 ;
        RECT 63.000 235.950 67.050 236.400 ;
        RECT 77.100 232.950 79.200 235.050 ;
        RECT 58.950 229.950 61.050 232.050 ;
        RECT 46.950 196.950 49.050 199.050 ;
        RECT 53.100 196.950 55.200 199.050 ;
        RECT 53.400 187.050 54.600 196.950 ;
        RECT 52.950 184.950 55.050 187.050 ;
        RECT 43.950 172.950 46.050 175.050 ;
        RECT 40.950 166.950 43.050 169.050 ;
        RECT 44.400 166.050 45.600 172.950 ;
        RECT 44.100 163.950 46.200 166.050 ;
        RECT 32.400 161.400 36.900 163.050 ;
        RECT 33.000 160.950 36.900 161.400 ;
        RECT 46.950 160.950 49.050 163.050 ;
        RECT 40.950 151.950 43.050 154.050 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 14.400 121.050 15.600 133.950 ;
        RECT 22.950 130.950 25.050 133.050 ;
        RECT 34.950 130.950 37.050 133.050 ;
        RECT 23.400 127.050 24.600 130.950 ;
        RECT 22.950 124.950 25.050 127.050 ;
        RECT 28.950 126.600 31.050 130.050 ;
        RECT 35.400 127.050 36.600 130.950 ;
        RECT 28.950 126.000 33.600 126.600 ;
        RECT 29.400 125.400 33.600 126.000 ;
        RECT 14.400 119.400 19.050 121.050 ;
        RECT 15.000 118.950 19.050 119.400 ;
        RECT 25.950 118.950 28.050 121.050 ;
        RECT 26.400 115.050 27.600 118.950 ;
        RECT 32.400 118.050 33.600 125.400 ;
        RECT 34.950 124.950 37.050 127.050 ;
        RECT 35.400 121.050 36.600 124.950 ;
        RECT 34.950 118.950 37.050 121.050 ;
        RECT 31.950 115.950 34.050 118.050 ;
        RECT 25.950 112.950 28.050 115.050 ;
        RECT 13.950 100.950 16.050 106.050 ;
        RECT 26.400 94.050 27.600 112.950 ;
        RECT 28.950 97.950 31.050 100.050 ;
        RECT 25.950 91.950 28.050 94.050 ;
        RECT 29.400 88.050 30.600 97.950 ;
        RECT 32.400 94.050 33.600 115.950 ;
        RECT 38.400 100.050 39.600 133.950 ;
        RECT 37.950 97.950 40.050 100.050 ;
        RECT 32.400 92.400 37.050 94.050 ;
        RECT 33.000 91.950 37.050 92.400 ;
        RECT 28.950 85.950 31.050 88.050 ;
        RECT 41.400 85.050 42.600 151.950 ;
        RECT 47.400 103.050 48.600 160.950 ;
        RECT 59.400 153.600 60.600 229.950 ;
        RECT 77.400 205.050 78.600 232.950 ;
        RECT 86.400 232.050 87.600 238.950 ;
        RECT 104.400 235.050 105.600 256.950 ;
        RECT 110.400 244.050 111.600 286.950 ;
        RECT 112.950 283.950 115.050 286.050 ;
        RECT 113.400 274.050 114.600 283.950 ;
        RECT 118.950 280.950 121.050 283.050 ;
        RECT 112.950 271.950 115.050 274.050 ;
        RECT 119.400 268.050 120.600 280.950 ;
        RECT 118.950 265.950 121.050 268.050 ;
        RECT 125.400 247.050 126.600 334.950 ;
        RECT 127.950 313.950 130.050 316.050 ;
        RECT 128.400 307.050 129.600 313.950 ;
        RECT 131.400 309.600 132.600 364.950 ;
        RECT 137.400 361.050 138.600 373.950 ;
        RECT 148.950 370.950 151.050 373.050 ;
        RECT 145.950 361.950 148.050 364.050 ;
        RECT 136.950 358.950 139.050 361.050 ;
        RECT 133.950 352.950 136.050 355.050 ;
        RECT 134.400 343.050 135.600 352.950 ;
        RECT 137.400 346.050 138.600 358.950 ;
        RECT 146.400 349.050 147.600 361.950 ;
        RECT 145.950 346.950 148.050 349.050 ;
        RECT 149.400 346.050 150.600 370.950 ;
        RECT 155.400 349.050 156.600 373.950 ;
        RECT 173.400 358.050 174.600 382.950 ;
        RECT 178.950 379.950 181.050 382.050 ;
        RECT 185.400 381.600 186.600 412.950 ;
        RECT 182.400 380.400 186.600 381.600 ;
        RECT 179.400 376.050 180.600 379.950 ;
        RECT 178.950 373.950 181.050 376.050 ;
        RECT 182.400 375.600 183.600 380.400 ;
        RECT 187.950 376.950 190.050 379.050 ;
        RECT 182.400 374.400 186.600 375.600 ;
        RECT 178.950 364.950 181.050 367.050 ;
        RECT 172.950 355.950 175.050 358.050 ;
        RECT 154.950 346.950 157.050 349.050 ;
        RECT 175.950 346.950 178.050 349.050 ;
        RECT 137.100 343.950 139.200 346.050 ;
        RECT 148.950 343.950 151.050 346.050 ;
        RECT 133.800 340.950 135.900 343.050 ;
        RECT 142.950 316.950 145.050 319.050 ;
        RECT 143.400 310.050 144.600 316.950 ;
        RECT 149.400 316.050 150.600 343.950 ;
        RECT 155.400 343.050 156.600 346.950 ;
        RECT 176.400 343.050 177.600 346.950 ;
        RECT 154.950 340.950 157.050 343.050 ;
        RECT 168.000 342.600 172.050 343.050 ;
        RECT 167.400 340.950 172.050 342.600 ;
        RECT 175.950 340.950 178.050 343.050 ;
        RECT 157.950 334.950 160.050 337.050 ;
        RECT 148.950 313.950 151.050 316.050 ;
        RECT 131.400 308.400 135.600 309.600 ;
        RECT 127.950 304.950 130.050 307.050 ;
        RECT 134.400 283.050 135.600 308.400 ;
        RECT 142.950 307.950 145.050 310.050 ;
        RECT 158.400 307.050 159.600 334.950 ;
        RECT 167.400 316.050 168.600 340.950 ;
        RECT 172.950 316.950 175.050 319.050 ;
        RECT 166.950 313.950 169.050 316.050 ;
        RECT 173.400 313.050 174.600 316.950 ;
        RECT 172.950 310.950 175.050 313.050 ;
        RECT 158.400 305.400 163.050 307.050 ;
        RECT 159.000 304.950 163.050 305.400 ;
        RECT 136.950 298.950 139.050 304.050 ;
        RECT 179.400 286.050 180.600 364.950 ;
        RECT 185.400 363.600 186.600 374.400 ;
        RECT 188.400 370.050 189.600 376.950 ;
        RECT 187.950 367.950 190.050 370.050 ;
        RECT 182.400 362.400 186.600 363.600 ;
        RECT 182.400 328.050 183.600 362.400 ;
        RECT 184.950 346.950 187.050 352.050 ;
        RECT 187.950 337.950 190.050 340.050 ;
        RECT 188.400 328.050 189.600 337.950 ;
        RECT 181.950 325.950 184.050 328.050 ;
        RECT 187.950 325.950 190.050 328.050 ;
        RECT 184.950 322.950 187.050 325.050 ;
        RECT 190.950 322.950 193.050 325.050 ;
        RECT 178.950 283.950 181.050 286.050 ;
        RECT 133.950 280.950 136.050 283.050 ;
        RECT 136.950 274.950 139.050 280.050 ;
        RECT 154.950 274.950 157.050 277.050 ;
        RECT 145.950 271.950 148.050 274.050 ;
        RECT 133.950 265.950 136.050 268.050 ;
        RECT 130.950 262.950 133.050 265.050 ;
        RECT 124.950 244.950 127.050 247.050 ;
        RECT 109.950 243.600 112.050 244.050 ;
        RECT 107.400 242.400 112.050 243.600 ;
        RECT 103.950 232.950 106.050 235.050 ;
        RECT 85.950 229.950 88.050 232.050 ;
        RECT 103.950 211.950 106.050 214.050 ;
        RECT 94.950 208.950 97.050 211.050 ;
        RECT 85.950 205.950 88.050 208.050 ;
        RECT 76.950 202.950 79.050 205.050 ;
        RECT 73.950 199.950 76.050 202.050 ;
        RECT 64.950 196.950 67.050 199.050 ;
        RECT 65.400 178.050 66.600 196.950 ;
        RECT 64.950 175.950 67.050 178.050 ;
        RECT 65.400 169.050 66.600 175.950 ;
        RECT 74.400 172.050 75.600 199.950 ;
        RECT 80.100 198.600 84.000 199.050 ;
        RECT 80.100 196.950 84.600 198.600 ;
        RECT 83.400 190.050 84.600 196.950 ;
        RECT 82.950 187.950 85.050 190.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 73.950 169.950 76.050 172.050 ;
        RECT 64.950 166.950 67.050 169.050 ;
        RECT 83.400 163.050 84.600 178.950 ;
        RECT 82.950 160.950 85.050 163.050 ;
        RECT 56.400 152.400 60.600 153.600 ;
        RECT 56.400 142.050 57.600 152.400 ;
        RECT 55.950 139.950 58.050 142.050 ;
        RECT 49.950 136.950 52.050 139.050 ;
        RECT 50.400 130.050 51.600 136.950 ;
        RECT 49.950 127.950 52.050 130.050 ;
        RECT 55.950 127.950 58.050 130.050 ;
        RECT 50.400 106.050 51.600 127.950 ;
        RECT 52.950 109.950 55.050 112.050 ;
        RECT 49.950 103.950 52.050 106.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 53.400 94.200 54.600 109.950 ;
        RECT 56.400 97.050 57.600 127.950 ;
        RECT 61.950 126.600 66.000 127.050 ;
        RECT 61.950 124.950 66.600 126.600 ;
        RECT 68.100 124.950 70.200 127.050 ;
        RECT 65.400 121.050 66.600 124.950 ;
        RECT 64.950 118.950 67.050 121.050 ;
        RECT 68.400 115.050 69.600 124.950 ;
        RECT 86.400 124.050 87.600 205.950 ;
        RECT 95.400 202.050 96.600 208.950 ;
        RECT 94.950 199.950 97.050 202.050 ;
        RECT 95.400 193.050 96.600 199.950 ;
        RECT 100.800 193.950 102.900 196.050 ;
        RECT 94.950 190.950 97.050 193.050 ;
        RECT 101.400 184.050 102.600 193.950 ;
        RECT 100.950 181.950 103.050 184.050 ;
        RECT 101.400 175.050 102.600 181.950 ;
        RECT 100.950 172.950 103.050 175.050 ;
        RECT 91.950 169.950 94.050 172.050 ;
        RECT 92.400 166.050 93.600 169.950 ;
        RECT 88.950 164.400 93.600 166.050 ;
        RECT 88.950 163.950 93.000 164.400 ;
        RECT 100.950 163.950 103.050 166.050 ;
        RECT 101.400 160.050 102.600 163.950 ;
        RECT 100.950 157.950 103.050 160.050 ;
        RECT 104.400 139.050 105.600 211.950 ;
        RECT 88.950 136.950 91.050 139.050 ;
        RECT 103.950 136.950 106.050 139.050 ;
        RECT 89.400 127.050 90.600 136.950 ;
        RECT 107.400 136.050 108.600 242.400 ;
        RECT 109.950 241.950 112.050 242.400 ;
        RECT 125.400 241.050 126.600 244.950 ;
        RECT 116.100 238.950 118.200 241.050 ;
        RECT 125.100 238.950 127.200 241.050 ;
        RECT 116.400 235.050 117.600 238.950 ;
        RECT 131.400 237.600 132.600 262.950 ;
        RECT 134.400 262.050 135.600 265.950 ;
        RECT 139.950 262.950 142.050 268.050 ;
        RECT 133.950 259.950 136.050 262.050 ;
        RECT 146.400 253.050 147.600 271.950 ;
        RECT 155.400 271.050 156.600 274.950 ;
        RECT 151.950 269.400 156.600 271.050 ;
        RECT 151.950 268.950 156.000 269.400 ;
        RECT 172.950 268.950 175.050 271.050 ;
        RECT 148.950 265.950 151.050 268.050 ;
        RECT 161.100 267.000 163.200 268.050 ;
        RECT 160.950 265.950 163.200 267.000 ;
        RECT 169.950 265.950 172.050 268.050 ;
        RECT 149.400 262.050 150.600 265.950 ;
        RECT 160.950 262.950 163.050 265.950 ;
        RECT 148.800 259.950 150.900 262.050 ;
        RECT 152.100 259.950 154.200 262.050 ;
        RECT 145.950 250.950 148.050 253.050 ;
        RECT 139.950 240.600 142.050 244.050 ;
        RECT 152.400 241.050 153.600 259.950 ;
        RECT 157.950 253.950 160.050 256.050 ;
        RECT 158.400 247.050 159.600 253.950 ;
        RECT 157.950 244.950 160.050 247.050 ;
        RECT 158.400 241.050 159.600 244.950 ;
        RECT 170.400 244.050 171.600 265.950 ;
        RECT 169.950 241.950 172.050 244.050 ;
        RECT 173.400 241.050 174.600 268.950 ;
        RECT 175.950 262.950 178.050 265.050 ;
        RECT 176.400 259.050 177.600 262.950 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 137.400 240.000 142.050 240.600 ;
        RECT 137.400 239.400 141.600 240.000 ;
        RECT 137.400 237.600 138.600 239.400 ;
        RECT 151.800 238.950 153.900 241.050 ;
        RECT 155.100 239.400 159.600 241.050 ;
        RECT 155.100 238.950 159.000 239.400 ;
        RECT 172.950 238.950 175.050 241.050 ;
        RECT 128.400 236.400 132.600 237.600 ;
        RECT 134.400 237.000 138.600 237.600 ;
        RECT 133.950 236.400 138.600 237.000 ;
        RECT 115.950 232.950 118.050 235.050 ;
        RECT 128.400 217.050 129.600 236.400 ;
        RECT 133.950 235.050 136.050 236.400 ;
        RECT 133.800 234.000 136.050 235.050 ;
        RECT 133.800 232.950 135.900 234.000 ;
        RECT 137.100 232.950 139.200 235.050 ;
        RECT 127.950 214.950 130.050 217.050 ;
        RECT 137.400 214.050 138.600 232.950 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 208.950 142.050 211.050 ;
        RECT 118.950 202.950 121.050 205.050 ;
        RECT 119.400 199.050 120.600 202.950 ;
        RECT 140.400 199.050 141.600 208.950 ;
        RECT 152.400 208.050 153.600 238.950 ;
        RECT 160.950 232.950 163.050 235.050 ;
        RECT 161.400 229.050 162.600 232.950 ;
        RECT 160.950 226.950 163.050 229.050 ;
        RECT 151.950 205.950 154.050 208.050 ;
        RECT 148.950 199.950 151.050 202.050 ;
        RECT 118.800 196.950 120.900 199.050 ;
        RECT 124.950 196.950 127.050 199.050 ;
        RECT 130.950 198.600 135.000 199.050 ;
        RECT 130.950 196.950 135.600 198.600 ;
        RECT 139.950 196.950 142.050 199.050 ;
        RECT 112.950 193.950 115.050 196.050 ;
        RECT 113.400 178.050 114.600 193.950 ;
        RECT 112.950 175.950 115.050 178.050 ;
        RECT 113.400 169.050 114.600 175.950 ;
        RECT 119.400 175.050 120.600 196.950 ;
        RECT 125.400 184.050 126.600 196.950 ;
        RECT 127.950 193.950 130.050 196.050 ;
        RECT 128.400 184.050 129.600 193.950 ;
        RECT 134.400 187.050 135.600 196.950 ;
        RECT 133.950 184.950 136.050 187.050 ;
        RECT 124.800 181.950 126.900 184.050 ;
        RECT 128.100 181.950 130.200 184.050 ;
        RECT 118.950 172.950 121.050 175.050 ;
        RECT 109.950 167.400 114.600 169.050 ;
        RECT 109.950 166.950 114.000 167.400 ;
        RECT 119.400 163.050 120.600 172.950 ;
        RECT 128.400 166.050 129.600 181.950 ;
        RECT 127.950 163.950 130.050 166.050 ;
        RECT 134.400 163.050 135.600 184.950 ;
        RECT 149.400 175.050 150.600 199.950 ;
        RECT 161.400 193.050 162.600 226.950 ;
        RECT 166.950 217.950 169.050 220.050 ;
        RECT 167.400 196.050 168.600 217.950 ;
        RECT 176.400 205.050 177.600 256.950 ;
        RECT 185.400 256.050 186.600 322.950 ;
        RECT 191.400 319.050 192.600 322.950 ;
        RECT 190.950 316.950 193.050 319.050 ;
        RECT 191.400 310.050 192.600 316.950 ;
        RECT 190.950 307.950 193.050 310.050 ;
        RECT 190.950 265.950 193.050 268.050 ;
        RECT 178.950 253.950 181.050 256.050 ;
        RECT 184.950 253.950 187.050 256.050 ;
        RECT 179.400 217.050 180.600 253.950 ;
        RECT 191.400 244.050 192.600 265.950 ;
        RECT 194.400 265.050 195.600 466.950 ;
        RECT 196.950 460.950 199.050 463.050 ;
        RECT 197.400 385.050 198.600 460.950 ;
        RECT 203.400 454.050 204.600 478.950 ;
        RECT 206.400 457.050 207.600 526.950 ;
        RECT 218.400 526.050 219.600 538.950 ;
        RECT 217.950 523.950 220.050 526.050 ;
        RECT 214.800 520.950 216.900 523.050 ;
        RECT 215.400 508.050 216.600 520.950 ;
        RECT 214.950 505.950 217.050 508.050 ;
        RECT 208.950 487.950 211.050 490.050 ;
        RECT 209.400 472.050 210.600 487.950 ;
        RECT 208.950 469.950 211.050 472.050 ;
        RECT 218.400 463.050 219.600 523.950 ;
        RECT 221.400 511.050 222.600 541.950 ;
        RECT 230.400 529.050 231.600 592.950 ;
        RECT 239.400 577.050 240.600 592.950 ;
        RECT 238.950 574.950 241.050 577.050 ;
        RECT 232.950 571.950 235.050 574.050 ;
        RECT 233.400 559.050 234.600 571.950 ;
        RECT 238.950 565.950 241.050 568.050 ;
        RECT 233.400 557.400 238.050 559.050 ;
        RECT 234.000 556.950 238.050 557.400 ;
        RECT 239.400 553.050 240.600 565.950 ;
        RECT 238.950 550.950 241.050 553.050 ;
        RECT 232.950 538.950 235.050 541.050 ;
        RECT 233.400 535.050 234.600 538.950 ;
        RECT 242.400 535.050 243.600 619.800 ;
        RECT 245.400 607.200 246.600 682.950 ;
        RECT 248.400 676.050 249.600 688.950 ;
        RECT 253.950 685.950 256.050 688.050 ;
        RECT 247.950 673.950 250.050 676.050 ;
        RECT 248.400 670.050 249.600 673.950 ;
        RECT 254.400 670.050 255.600 685.950 ;
        RECT 263.400 685.050 264.600 691.950 ;
        RECT 262.950 682.950 265.050 685.050 ;
        RECT 259.950 679.950 262.050 682.050 ;
        RECT 260.400 673.050 261.600 679.950 ;
        RECT 269.400 673.050 270.600 703.950 ;
        RECT 285.000 702.600 288.900 703.050 ;
        RECT 284.400 700.950 288.900 702.600 ;
        RECT 277.950 694.950 280.050 697.050 ;
        RECT 278.400 673.050 279.600 694.950 ;
        RECT 284.400 691.050 285.600 700.950 ;
        RECT 283.950 688.950 286.050 691.050 ;
        RECT 286.950 679.950 289.050 682.050 ;
        RECT 260.400 671.400 265.050 673.050 ;
        RECT 261.000 670.950 265.050 671.400 ;
        RECT 268.950 670.950 271.050 673.050 ;
        RECT 277.800 670.950 279.900 673.050 ;
        RECT 248.100 667.950 250.200 670.050 ;
        RECT 253.950 667.950 256.050 670.050 ;
        RECT 254.400 646.050 255.600 667.950 ;
        RECT 253.950 643.950 256.050 646.050 ;
        RECT 263.400 640.050 264.600 670.950 ;
        RECT 287.400 670.050 288.600 679.950 ;
        RECT 286.950 669.600 289.050 670.050 ;
        RECT 286.950 668.400 291.600 669.600 ;
        RECT 286.950 667.950 289.050 668.400 ;
        RECT 290.400 664.050 291.600 668.400 ;
        RECT 293.400 667.050 294.600 709.950 ;
        RECT 301.800 703.950 303.900 706.050 ;
        RECT 305.100 705.000 307.200 706.050 ;
        RECT 304.950 703.950 307.200 705.000 ;
        RECT 302.400 700.050 303.600 703.950 ;
        RECT 304.950 702.600 307.050 703.950 ;
        RECT 316.950 702.600 319.050 703.050 ;
        RECT 304.950 702.000 319.050 702.600 ;
        RECT 305.400 701.400 319.050 702.000 ;
        RECT 316.950 700.950 319.050 701.400 ;
        RECT 302.100 697.950 304.200 700.050 ;
        RECT 311.100 697.950 313.200 700.050 ;
        RECT 311.400 691.050 312.600 697.950 ;
        RECT 316.950 694.950 319.050 697.050 ;
        RECT 310.950 688.950 313.050 691.050 ;
        RECT 307.950 676.950 310.050 679.050 ;
        RECT 299.400 669.000 303.600 669.600 ;
        RECT 298.950 668.400 303.600 669.000 ;
        RECT 298.950 667.050 301.050 668.400 ;
        RECT 292.950 664.950 295.050 667.050 ;
        RECT 298.800 666.000 301.050 667.050 ;
        RECT 298.800 664.950 300.900 666.000 ;
        RECT 289.950 661.950 292.050 664.050 ;
        RECT 286.950 658.950 289.050 661.050 ;
        RECT 287.400 655.050 288.600 658.950 ;
        RECT 302.400 658.050 303.600 668.400 ;
        RECT 308.400 661.050 309.600 676.950 ;
        RECT 317.400 673.050 318.600 694.950 ;
        RECT 316.950 669.000 319.050 673.050 ;
        RECT 317.400 668.400 318.600 669.000 ;
        RECT 307.950 658.950 310.050 661.050 ;
        RECT 301.950 655.950 304.050 658.050 ;
        RECT 286.950 652.950 289.050 655.050 ;
        RECT 262.950 637.950 265.050 640.050 ;
        RECT 274.950 637.950 277.050 640.050 ;
        RECT 275.400 634.050 276.600 637.950 ;
        RECT 259.950 631.950 262.050 634.050 ;
        RECT 268.800 633.600 273.000 634.050 ;
        RECT 268.800 633.000 273.600 633.600 ;
        RECT 268.800 631.950 274.050 633.000 ;
        RECT 274.950 631.950 277.050 634.050 ;
        RECT 252.000 630.600 255.900 631.050 ;
        RECT 251.400 628.950 255.900 630.600 ;
        RECT 251.400 622.050 252.600 628.950 ;
        RECT 260.400 628.050 261.600 631.950 ;
        RECT 271.950 631.050 274.050 631.950 ;
        RECT 265.950 628.950 268.050 631.050 ;
        RECT 271.950 630.000 274.200 631.050 ;
        RECT 272.100 628.950 274.200 630.000 ;
        RECT 283.950 628.950 286.050 631.050 ;
        RECT 259.950 625.950 262.050 628.050 ;
        RECT 250.950 619.950 253.050 622.050 ;
        RECT 266.400 619.050 267.600 628.950 ;
        RECT 271.950 622.950 274.050 625.050 ;
        RECT 265.950 616.950 268.050 619.050 ;
        RECT 244.950 605.100 247.050 607.200 ;
        RECT 246.000 603.900 249.000 604.050 ;
        RECT 244.950 603.450 249.000 603.900 ;
        RECT 244.950 601.950 249.600 603.450 ;
        RECT 244.950 601.800 247.050 601.950 ;
        RECT 248.400 592.050 249.600 601.950 ;
        RECT 266.100 592.950 268.200 595.050 ;
        RECT 247.950 589.950 250.050 592.050 ;
        RECT 266.400 583.050 267.600 592.950 ;
        RECT 268.950 589.950 271.050 592.050 ;
        RECT 265.950 580.950 268.050 583.050 ;
        RECT 244.950 574.950 247.050 577.050 ;
        RECT 259.950 574.950 262.050 577.050 ;
        RECT 245.400 552.600 246.600 574.950 ;
        RECT 247.950 568.950 250.050 571.050 ;
        RECT 248.400 562.050 249.600 568.950 ;
        RECT 260.400 565.050 261.600 574.950 ;
        RECT 262.950 571.950 265.050 574.050 ;
        RECT 259.950 562.950 262.050 565.050 ;
        RECT 247.950 559.950 250.050 562.050 ;
        RECT 248.400 556.050 249.600 559.950 ;
        RECT 263.400 556.050 264.600 571.950 ;
        RECT 265.950 562.950 268.050 565.050 ;
        RECT 266.400 559.050 267.600 562.950 ;
        RECT 265.950 556.950 268.050 559.050 ;
        RECT 247.800 553.950 249.900 556.050 ;
        RECT 262.950 553.950 265.050 556.050 ;
        RECT 245.400 551.400 249.600 552.600 ;
        RECT 232.950 532.950 235.050 535.050 ;
        RECT 241.950 532.950 244.050 535.050 ;
        RECT 229.950 526.950 232.050 529.050 ;
        RECT 236.100 526.950 238.200 529.050 ;
        RECT 236.400 517.050 237.600 526.950 ;
        RECT 248.400 526.050 249.600 551.400 ;
        RECT 265.950 550.950 268.050 553.050 ;
        RECT 259.950 535.950 262.050 538.050 ;
        RECT 260.400 532.050 261.600 535.950 ;
        RECT 259.950 528.000 262.050 532.050 ;
        RECT 266.400 529.050 267.600 550.950 ;
        RECT 260.400 527.400 261.600 528.000 ;
        RECT 265.950 526.950 268.050 529.050 ;
        RECT 241.950 523.950 244.050 526.050 ;
        RECT 247.950 523.950 250.050 526.050 ;
        RECT 226.800 514.950 228.900 517.050 ;
        RECT 235.950 514.950 238.050 517.050 ;
        RECT 220.950 508.950 223.050 511.050 ;
        RECT 220.950 493.950 223.050 496.050 ;
        RECT 217.950 460.950 220.050 463.050 ;
        RECT 205.950 454.950 208.050 457.050 ;
        RECT 221.400 454.050 222.600 493.950 ;
        RECT 227.400 454.050 228.600 514.950 ;
        RECT 232.950 499.950 235.050 502.050 ;
        RECT 202.950 451.950 205.050 454.050 ;
        RECT 220.950 451.950 223.050 454.050 ;
        RECT 227.100 451.950 229.200 454.050 ;
        RECT 217.950 448.950 220.050 451.050 ;
        RECT 202.950 442.950 205.050 448.050 ;
        RECT 203.400 412.050 204.600 442.950 ;
        RECT 218.400 415.050 219.600 448.950 ;
        RECT 221.400 442.050 222.600 451.950 ;
        RECT 233.400 448.050 234.600 499.950 ;
        RECT 236.400 484.050 237.600 514.950 ;
        RECT 242.400 496.050 243.600 523.950 ;
        RECT 253.950 511.950 256.050 514.050 ;
        RECT 241.950 493.950 244.050 496.050 ;
        RECT 254.400 493.050 255.600 511.950 ;
        RECT 259.950 499.950 262.050 502.050 ;
        RECT 260.400 496.050 261.600 499.950 ;
        RECT 259.950 493.950 262.050 496.050 ;
        RECT 253.800 490.950 255.900 493.050 ;
        RECT 257.100 492.000 259.200 493.050 ;
        RECT 256.950 490.950 259.200 492.000 ;
        RECT 256.950 489.600 259.050 490.950 ;
        RECT 266.400 490.050 267.600 526.950 ;
        RECT 269.400 493.050 270.600 589.950 ;
        RECT 272.400 585.600 273.600 622.950 ;
        RECT 284.400 601.050 285.600 628.950 ;
        RECT 280.950 599.400 285.600 601.050 ;
        RECT 280.950 598.950 285.000 599.400 ;
        RECT 287.400 595.050 288.600 652.950 ;
        RECT 289.950 649.950 292.050 652.050 ;
        RECT 290.400 639.600 291.600 649.950 ;
        RECT 290.400 638.400 294.600 639.600 ;
        RECT 293.400 631.050 294.600 638.400 ;
        RECT 304.950 633.600 307.050 637.050 ;
        RECT 308.400 633.600 309.600 658.950 ;
        RECT 310.950 643.950 313.050 646.050 ;
        RECT 304.950 633.000 309.600 633.600 ;
        RECT 305.400 632.400 309.600 633.000 ;
        RECT 290.100 628.950 294.600 631.050 ;
        RECT 298.950 628.950 301.050 631.050 ;
        RECT 286.950 589.950 289.050 595.050 ;
        RECT 272.400 584.400 276.600 585.600 ;
        RECT 271.950 580.950 274.050 583.050 ;
        RECT 272.400 553.050 273.600 580.950 ;
        RECT 271.950 550.950 274.050 553.050 ;
        RECT 275.400 541.050 276.600 584.400 ;
        RECT 293.400 577.050 294.600 628.950 ;
        RECT 295.950 625.950 298.050 628.050 ;
        RECT 296.400 610.050 297.600 625.950 ;
        RECT 299.400 616.050 300.600 628.950 ;
        RECT 298.950 613.950 301.050 616.050 ;
        RECT 308.400 613.050 309.600 632.400 ;
        RECT 311.400 631.050 312.600 643.950 ;
        RECT 322.950 637.950 325.050 640.050 ;
        RECT 316.950 631.950 319.050 634.050 ;
        RECT 311.100 628.950 313.200 631.050 ;
        RECT 311.400 616.050 312.600 628.950 ;
        RECT 317.400 628.050 318.600 631.950 ;
        RECT 323.400 631.050 324.600 637.950 ;
        RECT 322.950 628.950 325.050 631.050 ;
        RECT 316.800 625.950 318.900 628.050 ;
        RECT 319.950 616.950 322.050 619.050 ;
        RECT 310.950 613.950 313.050 616.050 ;
        RECT 316.950 613.950 319.050 616.050 ;
        RECT 307.950 610.950 310.050 613.050 ;
        RECT 295.950 607.950 298.050 610.050 ;
        RECT 313.950 607.950 316.050 610.050 ;
        RECT 314.400 601.050 315.600 607.950 ;
        RECT 313.950 598.950 316.050 601.050 ;
        RECT 317.400 598.050 318.600 613.950 ;
        RECT 316.950 595.950 319.050 598.050 ;
        RECT 317.400 589.050 318.600 595.950 ;
        RECT 298.950 586.950 301.050 589.050 ;
        RECT 316.950 586.950 319.050 589.050 ;
        RECT 292.950 574.950 295.050 577.050 ;
        RECT 277.950 565.950 280.050 568.050 ;
        RECT 295.950 565.950 298.050 568.050 ;
        RECT 278.400 550.050 279.600 565.950 ;
        RECT 283.950 559.950 286.050 562.050 ;
        RECT 284.400 556.050 285.600 559.950 ;
        RECT 296.400 556.050 297.600 565.950 ;
        RECT 283.950 553.950 286.050 556.050 ;
        RECT 295.950 553.950 298.050 556.050 ;
        RECT 277.950 547.950 280.050 550.050 ;
        RECT 286.950 544.950 289.050 547.050 ;
        RECT 274.950 538.950 277.050 541.050 ;
        RECT 271.950 532.950 274.050 535.050 ;
        RECT 268.950 490.950 271.050 493.050 ;
        RECT 254.400 489.000 259.050 489.600 ;
        RECT 254.400 488.400 258.600 489.000 ;
        RECT 235.800 481.950 237.900 484.050 ;
        RECT 247.950 481.950 250.050 484.050 ;
        RECT 236.400 457.050 237.600 481.950 ;
        RECT 235.950 454.950 238.050 457.050 ;
        RECT 232.950 445.950 235.050 448.050 ;
        RECT 220.950 439.950 223.050 442.050 ;
        RECT 248.400 436.050 249.600 481.950 ;
        RECT 247.950 433.950 250.050 436.050 ;
        RECT 248.400 415.050 249.600 433.950 ;
        RECT 254.400 430.050 255.600 488.400 ;
        RECT 259.950 487.950 262.050 490.050 ;
        RECT 265.950 487.950 268.050 490.050 ;
        RECT 253.950 427.950 256.050 430.050 ;
        RECT 260.400 424.050 261.600 487.950 ;
        RECT 262.950 466.950 265.050 469.050 ;
        RECT 263.400 454.050 264.600 466.950 ;
        RECT 265.950 454.950 268.050 457.050 ;
        RECT 262.950 451.950 265.050 454.050 ;
        RECT 259.950 421.950 262.050 424.050 ;
        RECT 250.950 415.950 253.050 418.050 ;
        RECT 217.950 412.950 220.050 415.050 ;
        RECT 247.950 412.950 250.050 415.050 ;
        RECT 202.950 409.950 205.050 412.050 ;
        RECT 227.100 409.950 229.200 412.050 ;
        RECT 217.950 394.950 220.050 397.050 ;
        RECT 208.950 391.950 211.050 394.050 ;
        RECT 205.950 385.950 208.050 388.050 ;
        RECT 196.950 382.950 199.050 385.050 ;
        RECT 196.950 373.950 199.050 376.050 ;
        RECT 197.400 349.050 198.600 373.950 ;
        RECT 196.950 346.950 199.050 349.050 ;
        RECT 206.400 346.050 207.600 385.950 ;
        RECT 209.400 355.050 210.600 391.950 ;
        RECT 214.950 379.950 217.050 382.050 ;
        RECT 215.400 370.050 216.600 379.950 ;
        RECT 214.950 367.950 217.050 370.050 ;
        RECT 211.950 364.950 214.050 367.050 ;
        RECT 208.950 352.950 211.050 355.050 ;
        RECT 205.950 343.950 208.050 346.050 ;
        RECT 201.000 342.600 205.050 343.050 ;
        RECT 200.400 340.950 205.050 342.600 ;
        RECT 200.400 318.600 201.600 340.950 ;
        RECT 202.950 334.950 205.050 337.050 ;
        RECT 203.400 325.050 204.600 334.950 ;
        RECT 212.400 334.050 213.600 364.950 ;
        RECT 215.400 343.050 216.600 367.950 ;
        RECT 214.950 340.950 217.050 343.050 ;
        RECT 211.950 331.950 214.050 334.050 ;
        RECT 214.950 325.950 217.050 328.050 ;
        RECT 202.950 322.950 205.050 325.050 ;
        RECT 197.400 317.400 201.600 318.600 ;
        RECT 197.400 307.050 198.600 317.400 ;
        RECT 215.400 316.050 216.600 325.950 ;
        RECT 218.400 324.600 219.600 394.950 ;
        RECT 227.400 394.050 228.600 409.950 ;
        RECT 247.950 397.950 250.050 400.050 ;
        RECT 226.950 391.950 229.050 394.050 ;
        RECT 241.950 391.950 244.050 394.050 ;
        RECT 229.950 385.950 232.050 388.050 ;
        RECT 225.000 381.600 229.050 382.050 ;
        RECT 224.400 379.950 229.050 381.600 ;
        RECT 224.400 346.050 225.600 379.950 ;
        RECT 230.400 376.050 231.600 385.950 ;
        RECT 242.400 385.050 243.600 391.950 ;
        RECT 241.950 382.950 244.050 385.050 ;
        RECT 235.950 376.950 238.050 379.050 ;
        RECT 229.950 373.950 232.050 376.050 ;
        RECT 226.950 346.950 229.050 349.050 ;
        RECT 232.950 346.950 235.050 349.050 ;
        RECT 223.950 343.950 226.050 346.050 ;
        RECT 227.400 337.050 228.600 346.950 ;
        RECT 233.400 340.050 234.600 346.950 ;
        RECT 232.950 337.950 235.050 340.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 236.400 331.050 237.600 376.950 ;
        RECT 238.950 358.950 241.050 361.050 ;
        RECT 239.400 336.600 240.600 358.950 ;
        RECT 241.950 340.950 244.050 346.050 ;
        RECT 239.400 335.400 243.600 336.600 ;
        RECT 235.950 328.950 238.050 331.050 ;
        RECT 218.400 323.400 222.600 324.600 ;
        RECT 199.950 313.950 202.050 316.050 ;
        RECT 215.400 314.400 220.050 316.050 ;
        RECT 216.000 313.950 220.050 314.400 ;
        RECT 200.400 310.050 201.600 313.950 ;
        RECT 221.400 310.050 222.600 323.400 ;
        RECT 223.950 316.950 226.050 319.050 ;
        RECT 242.400 318.600 243.600 335.400 ;
        RECT 248.400 322.050 249.600 397.950 ;
        RECT 251.400 361.200 252.600 415.950 ;
        RECT 253.950 412.950 256.050 415.050 ;
        RECT 254.400 397.050 255.600 412.950 ;
        RECT 266.400 409.050 267.600 454.950 ;
        RECT 268.950 442.950 271.050 445.050 ;
        RECT 256.950 406.950 259.050 409.050 ;
        RECT 265.950 406.950 268.050 409.050 ;
        RECT 253.950 394.950 256.050 397.050 ;
        RECT 253.950 388.950 256.050 391.050 ;
        RECT 250.950 359.100 253.050 361.200 ;
        RECT 250.950 355.800 253.050 357.900 ;
        RECT 247.950 319.950 250.050 322.050 ;
        RECT 242.400 317.400 246.600 318.600 ;
        RECT 224.400 313.050 225.600 316.950 ;
        RECT 232.950 313.950 235.050 316.050 ;
        RECT 223.950 310.950 226.050 313.050 ;
        RECT 200.400 308.400 205.050 310.050 ;
        RECT 201.000 307.950 205.050 308.400 ;
        RECT 220.950 307.950 223.050 310.050 ;
        RECT 226.950 307.950 229.050 310.050 ;
        RECT 197.400 306.900 201.000 307.050 ;
        RECT 197.400 305.250 202.050 306.900 ;
        RECT 198.000 304.950 202.050 305.250 ;
        RECT 199.950 304.800 202.050 304.950 ;
        RECT 227.400 298.050 228.600 307.950 ;
        RECT 226.950 295.950 229.050 298.050 ;
        RECT 233.400 289.050 234.600 313.950 ;
        RECT 245.400 307.050 246.600 317.400 ;
        RECT 248.400 316.050 249.600 319.950 ;
        RECT 247.950 313.950 250.050 316.050 ;
        RECT 251.400 310.050 252.600 355.800 ;
        RECT 254.400 343.050 255.600 388.950 ;
        RECT 253.950 340.950 256.050 343.050 ;
        RECT 257.400 319.050 258.600 406.950 ;
        RECT 266.400 397.050 267.600 406.950 ;
        RECT 265.950 394.950 268.050 397.050 ;
        RECT 265.950 388.950 268.050 391.050 ;
        RECT 266.400 388.050 267.600 388.950 ;
        RECT 262.800 382.950 264.900 385.050 ;
        RECT 265.950 384.000 268.050 388.050 ;
        RECT 266.400 383.400 267.600 384.000 ;
        RECT 259.950 379.950 262.050 382.050 ;
        RECT 260.400 370.050 261.600 379.950 ;
        RECT 259.950 367.950 262.050 370.050 ;
        RECT 263.400 358.050 264.600 382.950 ;
        RECT 269.400 382.050 270.600 442.950 ;
        RECT 272.400 442.050 273.600 532.950 ;
        RECT 280.950 529.950 283.050 532.050 ;
        RECT 277.950 520.950 280.050 523.050 ;
        RECT 278.400 508.050 279.600 520.950 ;
        RECT 277.950 505.950 280.050 508.050 ;
        RECT 281.400 505.050 282.600 529.950 ;
        RECT 287.400 523.050 288.600 544.950 ;
        RECT 295.950 529.950 298.050 532.050 ;
        RECT 287.400 521.400 292.050 523.050 ;
        RECT 288.000 520.950 292.050 521.400 ;
        RECT 283.950 514.950 286.050 517.050 ;
        RECT 280.950 502.950 283.050 505.050 ;
        RECT 284.400 490.050 285.600 514.950 ;
        RECT 296.400 508.050 297.600 529.950 ;
        RECT 299.400 517.050 300.600 586.950 ;
        RECT 313.950 583.950 316.050 586.050 ;
        RECT 302.100 571.950 304.200 574.050 ;
        RECT 302.400 565.050 303.600 571.950 ;
        RECT 314.400 568.050 315.600 583.950 ;
        RECT 314.100 565.950 316.200 568.050 ;
        RECT 301.950 562.950 304.050 565.050 ;
        RECT 307.800 559.950 309.900 562.050 ;
        RECT 316.950 559.950 319.050 562.050 ;
        RECT 304.950 556.950 307.050 559.050 ;
        RECT 305.400 553.050 306.600 556.950 ;
        RECT 304.950 550.950 307.050 553.050 ;
        RECT 308.400 550.050 309.600 559.950 ;
        RECT 317.400 556.050 318.600 559.950 ;
        RECT 316.950 553.950 319.050 556.050 ;
        RECT 307.950 547.950 310.050 550.050 ;
        RECT 313.950 544.950 316.050 547.050 ;
        RECT 314.400 540.600 315.600 544.950 ;
        RECT 311.400 539.400 315.600 540.600 ;
        RECT 301.950 535.950 304.050 538.050 ;
        RECT 302.400 532.050 303.600 535.950 ;
        RECT 302.100 529.950 304.200 532.050 ;
        RECT 311.400 526.050 312.600 539.400 ;
        RECT 317.400 529.050 318.600 553.950 ;
        RECT 316.950 526.950 319.050 529.050 ;
        RECT 310.950 523.950 313.050 526.050 ;
        RECT 316.950 520.950 319.050 523.050 ;
        RECT 298.950 514.950 301.050 517.050 ;
        RECT 304.950 514.950 307.050 517.050 ;
        RECT 295.950 505.950 298.050 508.050 ;
        RECT 298.950 502.950 301.050 505.050 ;
        RECT 295.950 496.950 298.050 499.050 ;
        RECT 283.950 487.950 286.050 490.050 ;
        RECT 292.950 487.950 295.050 490.050 ;
        RECT 289.950 484.950 292.050 487.050 ;
        RECT 274.950 475.950 277.050 478.050 ;
        RECT 275.400 457.050 276.600 475.950 ;
        RECT 286.950 472.950 289.050 475.050 ;
        RECT 277.950 463.950 280.050 466.050 ;
        RECT 274.950 454.950 277.050 457.050 ;
        RECT 271.950 439.950 274.050 442.050 ;
        RECT 278.400 418.050 279.600 463.950 ;
        RECT 280.950 454.950 283.050 457.050 ;
        RECT 281.400 448.050 282.600 454.950 ;
        RECT 287.400 454.050 288.600 472.950 ;
        RECT 283.950 452.400 288.600 454.050 ;
        RECT 283.950 451.950 288.000 452.400 ;
        RECT 280.950 445.950 283.050 448.050 ;
        RECT 277.950 415.950 280.050 418.050 ;
        RECT 273.000 411.600 277.050 412.050 ;
        RECT 272.400 409.950 277.050 411.600 ;
        RECT 272.400 400.050 273.600 409.950 ;
        RECT 281.400 409.050 282.600 445.950 ;
        RECT 290.400 433.050 291.600 484.950 ;
        RECT 293.400 454.050 294.600 487.950 ;
        RECT 296.400 484.050 297.600 496.950 ;
        RECT 295.950 481.950 298.050 484.050 ;
        RECT 299.400 466.050 300.600 502.950 ;
        RECT 305.400 501.600 306.600 514.950 ;
        RECT 317.400 502.050 318.600 520.950 ;
        RECT 302.400 500.400 306.600 501.600 ;
        RECT 302.400 466.050 303.600 500.400 ;
        RECT 316.950 499.950 319.050 502.050 ;
        RECT 309.000 489.600 313.050 490.050 ;
        RECT 308.400 487.950 313.050 489.600 ;
        RECT 316.950 487.950 319.050 490.050 ;
        RECT 308.400 466.050 309.600 487.950 ;
        RECT 317.400 472.050 318.600 487.950 ;
        RECT 320.400 475.050 321.600 616.950 ;
        RECT 329.400 607.050 330.600 718.950 ;
        RECT 356.400 700.050 357.600 733.950 ;
        RECT 370.950 727.950 373.050 730.050 ;
        RECT 367.950 709.950 370.050 712.050 ;
        RECT 361.950 700.950 364.050 703.050 ;
        RECT 352.800 697.950 354.900 700.050 ;
        RECT 356.400 698.400 361.050 700.050 ;
        RECT 357.000 697.950 361.050 698.400 ;
        RECT 343.950 685.950 346.050 688.050 ;
        RECT 344.400 673.050 345.600 685.950 ;
        RECT 353.400 685.050 354.600 697.950 ;
        RECT 362.400 691.050 363.600 700.950 ;
        RECT 364.950 697.950 367.050 700.050 ;
        RECT 361.950 688.950 364.050 691.050 ;
        RECT 352.950 682.950 355.050 685.050 ;
        RECT 344.400 671.400 349.050 673.050 ;
        RECT 345.000 670.950 349.050 671.400 ;
        RECT 362.400 670.050 363.600 688.950 ;
        RECT 365.400 682.050 366.600 697.950 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 364.950 673.950 367.050 676.050 ;
        RECT 338.100 667.950 340.200 670.050 ;
        RECT 361.950 667.950 364.050 670.050 ;
        RECT 334.800 664.950 336.900 667.050 ;
        RECT 335.400 661.200 336.600 664.950 ;
        RECT 334.950 659.100 337.050 661.200 ;
        RECT 334.950 655.800 337.050 657.900 ;
        RECT 335.400 637.050 336.600 655.800 ;
        RECT 338.400 652.050 339.600 667.950 ;
        RECT 355.950 661.950 358.050 664.050 ;
        RECT 343.950 655.950 346.050 658.050 ;
        RECT 337.950 649.950 340.050 652.050 ;
        RECT 334.950 634.950 337.050 637.050 ;
        RECT 344.400 631.050 345.600 655.950 ;
        RECT 356.400 646.050 357.600 661.950 ;
        RECT 361.950 649.950 364.050 652.050 ;
        RECT 355.950 643.950 358.050 646.050 ;
        RECT 355.950 637.950 358.050 640.050 ;
        RECT 347.100 631.950 349.200 634.050 ;
        RECT 334.950 628.950 337.050 631.050 ;
        RECT 343.800 628.950 345.900 631.050 ;
        RECT 335.400 619.050 336.600 628.950 ;
        RECT 337.950 625.950 340.050 628.050 ;
        RECT 334.950 616.950 337.050 619.050 ;
        RECT 329.400 605.400 334.050 607.050 ;
        RECT 330.000 604.950 334.050 605.400 ;
        RECT 338.400 604.050 339.600 625.950 ;
        RECT 347.400 625.050 348.600 631.950 ;
        RECT 356.400 628.050 357.600 637.950 ;
        RECT 355.950 625.950 358.050 628.050 ;
        RECT 346.950 622.950 349.050 625.050 ;
        RECT 352.950 619.950 355.050 622.050 ;
        RECT 343.950 610.950 346.050 613.050 ;
        RECT 325.950 601.950 328.050 604.050 ;
        RECT 337.950 601.950 340.050 604.050 ;
        RECT 326.400 582.600 327.600 601.950 ;
        RECT 344.400 595.050 345.600 610.950 ;
        RECT 331.950 592.950 334.050 595.050 ;
        RECT 343.950 592.950 346.050 595.050 ;
        RECT 326.400 581.400 330.600 582.600 ;
        RECT 322.950 574.950 325.050 577.050 ;
        RECT 323.400 520.050 324.600 574.950 ;
        RECT 329.400 562.050 330.600 581.400 ;
        RECT 328.950 559.950 331.050 562.050 ;
        RECT 328.950 550.950 331.050 556.050 ;
        RECT 332.400 523.050 333.600 592.950 ;
        RECT 334.950 577.950 337.050 580.050 ;
        RECT 335.400 556.050 336.600 577.950 ;
        RECT 353.400 562.050 354.600 619.950 ;
        RECT 362.400 601.050 363.600 649.950 ;
        RECT 365.400 613.050 366.600 673.950 ;
        RECT 364.950 610.950 367.050 613.050 ;
        RECT 361.950 598.950 364.050 601.050 ;
        RECT 368.400 586.050 369.600 709.950 ;
        RECT 371.400 619.050 372.600 727.950 ;
        RECT 373.950 724.950 376.050 727.050 ;
        RECT 374.400 622.050 375.600 724.950 ;
        RECT 389.400 718.050 390.600 736.950 ;
        RECT 388.950 715.950 391.050 718.050 ;
        RECT 398.400 703.050 399.600 742.950 ;
        RECT 400.950 736.950 403.050 739.050 ;
        RECT 401.400 715.050 402.600 736.950 ;
        RECT 404.400 718.050 405.600 742.950 ;
        RECT 413.400 721.050 414.600 743.400 ;
        RECT 415.950 742.950 418.050 743.400 ;
        RECT 419.400 730.050 420.600 745.950 ;
        RECT 434.400 745.050 435.600 751.950 ;
        RECT 433.950 742.950 436.050 745.050 ;
        RECT 436.950 739.950 439.050 742.050 ;
        RECT 426.000 738.600 430.050 739.050 ;
        RECT 425.400 736.950 430.050 738.600 ;
        RECT 418.950 727.950 421.050 730.050 ;
        RECT 425.400 727.050 426.600 736.950 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 430.950 724.950 433.050 727.050 ;
        RECT 412.950 718.950 415.050 721.050 ;
        RECT 425.400 718.050 426.600 724.950 ;
        RECT 403.950 715.950 406.050 718.050 ;
        RECT 415.800 715.950 417.900 718.050 ;
        RECT 419.100 715.950 421.200 718.050 ;
        RECT 424.950 715.950 427.050 718.050 ;
        RECT 400.950 712.950 403.050 715.050 ;
        RECT 378.000 702.600 382.050 703.050 ;
        RECT 377.400 700.950 382.050 702.600 ;
        RECT 392.100 700.950 394.200 703.050 ;
        RECT 397.950 700.950 400.050 703.050 ;
        RECT 377.400 673.200 378.600 700.950 ;
        RECT 392.400 679.050 393.600 700.950 ;
        RECT 391.950 676.950 394.050 679.050 ;
        RECT 376.950 671.100 379.050 673.200 ;
        RECT 388.950 670.950 391.050 673.050 ;
        RECT 378.000 669.600 382.050 670.050 ;
        RECT 377.400 667.950 382.050 669.600 ;
        RECT 377.400 658.050 378.600 667.950 ;
        RECT 389.400 664.050 390.600 670.950 ;
        RECT 394.800 667.950 396.900 670.050 ;
        RECT 395.400 664.050 396.600 667.950 ;
        RECT 382.950 661.950 385.050 664.050 ;
        RECT 388.950 661.950 391.050 664.050 ;
        RECT 394.950 661.950 397.050 664.050 ;
        RECT 376.950 655.950 379.050 658.050 ;
        RECT 376.950 646.950 379.050 649.050 ;
        RECT 377.400 625.050 378.600 646.950 ;
        RECT 383.400 637.050 384.600 661.950 ;
        RECT 401.400 655.050 402.600 712.950 ;
        RECT 406.950 700.950 409.050 703.050 ;
        RECT 403.950 691.950 406.050 694.050 ;
        RECT 404.400 679.050 405.600 691.950 ;
        RECT 403.950 676.950 406.050 679.050 ;
        RECT 407.400 675.600 408.600 700.950 ;
        RECT 416.400 699.600 417.600 715.950 ;
        RECT 419.400 703.200 420.600 715.950 ;
        RECT 418.950 701.100 421.050 703.200 ;
        RECT 420.000 699.600 424.050 700.050 ;
        RECT 416.400 698.400 424.050 699.600 ;
        RECT 419.400 697.950 424.050 698.400 ;
        RECT 412.950 682.950 415.050 685.050 ;
        RECT 409.950 676.950 412.050 679.050 ;
        RECT 404.400 675.000 408.600 675.600 ;
        RECT 403.950 674.400 408.600 675.000 ;
        RECT 403.950 673.050 406.050 674.400 ;
        RECT 410.400 673.050 411.600 676.950 ;
        RECT 403.800 672.000 406.050 673.050 ;
        RECT 403.800 670.950 405.900 672.000 ;
        RECT 409.950 670.950 412.050 673.050 ;
        RECT 403.950 664.950 406.050 667.050 ;
        RECT 409.950 664.950 412.050 667.050 ;
        RECT 404.400 661.050 405.600 664.950 ;
        RECT 403.950 658.950 406.050 661.050 ;
        RECT 394.950 652.950 397.050 655.050 ;
        RECT 400.950 652.950 403.050 655.050 ;
        RECT 382.950 634.950 385.050 637.050 ;
        RECT 383.400 628.050 384.600 634.950 ;
        RECT 395.400 634.050 396.600 652.950 ;
        RECT 410.400 646.050 411.600 664.950 ;
        RECT 409.950 643.950 412.050 646.050 ;
        RECT 395.100 631.950 397.200 634.050 ;
        RECT 385.950 630.600 390.000 631.050 ;
        RECT 385.950 629.400 393.600 630.600 ;
        RECT 385.950 628.950 390.600 629.400 ;
        RECT 382.950 625.950 385.050 628.050 ;
        RECT 376.950 622.950 379.050 625.050 ;
        RECT 373.950 619.950 376.050 622.050 ;
        RECT 382.950 619.950 385.050 622.050 ;
        RECT 370.950 616.950 373.050 619.050 ;
        RECT 379.950 613.950 382.050 616.050 ;
        RECT 370.950 601.950 373.050 604.050 ;
        RECT 371.400 594.600 372.600 601.950 ;
        RECT 380.400 601.050 381.600 613.950 ;
        RECT 379.950 598.950 382.050 601.050 ;
        RECT 383.400 597.600 384.600 619.950 ;
        RECT 389.400 616.050 390.600 628.950 ;
        RECT 392.400 625.050 393.600 629.400 ;
        RECT 406.950 628.950 409.050 631.050 ;
        RECT 399.000 627.600 402.900 628.050 ;
        RECT 398.400 625.950 402.900 627.600 ;
        RECT 391.950 622.950 394.050 625.050 ;
        RECT 388.950 613.950 391.050 616.050 ;
        RECT 391.950 610.950 394.050 613.050 ;
        RECT 380.400 596.400 384.600 597.600 ;
        RECT 371.400 593.400 375.600 594.600 ;
        RECT 370.950 586.950 373.050 589.050 ;
        RECT 367.950 583.950 370.050 586.050 ;
        RECT 364.950 568.950 367.050 571.050 ;
        RECT 337.950 559.950 340.050 562.050 ;
        RECT 352.950 559.950 355.050 562.050 ;
        RECT 358.950 559.950 361.050 562.050 ;
        RECT 334.950 553.950 337.050 556.050 ;
        RECT 335.400 550.050 336.600 553.950 ;
        RECT 334.950 547.950 337.050 550.050 ;
        RECT 338.400 532.050 339.600 559.950 ;
        RECT 352.950 553.950 355.050 556.050 ;
        RECT 349.950 541.950 352.050 544.050 ;
        RECT 350.400 532.050 351.600 541.950 ;
        RECT 337.950 529.950 340.050 532.050 ;
        RECT 349.950 529.950 352.050 532.050 ;
        RECT 353.400 529.200 354.600 553.950 ;
        RECT 359.400 553.050 360.600 559.950 ;
        RECT 365.400 559.050 366.600 568.950 ;
        RECT 361.950 557.400 366.600 559.050 ;
        RECT 361.950 556.950 366.000 557.400 ;
        RECT 371.400 555.600 372.600 586.950 ;
        RECT 368.400 554.400 372.600 555.600 ;
        RECT 358.950 550.950 361.050 553.050 ;
        RECT 355.950 547.950 358.050 550.050 ;
        RECT 340.950 526.950 343.050 529.050 ;
        RECT 352.950 527.100 355.050 529.200 ;
        RECT 331.950 520.950 334.050 523.050 ;
        RECT 337.950 520.950 340.050 523.050 ;
        RECT 322.950 517.950 325.050 520.050 ;
        RECT 338.400 517.050 339.600 520.950 ;
        RECT 337.950 514.950 340.050 517.050 ;
        RECT 335.100 511.950 337.200 514.050 ;
        RECT 328.950 490.950 331.050 496.050 ;
        RECT 326.400 486.000 327.600 486.600 ;
        RECT 325.950 481.950 328.050 486.000 ;
        RECT 322.950 478.950 325.050 481.050 ;
        RECT 319.950 472.950 322.050 475.050 ;
        RECT 316.950 469.950 319.050 472.050 ;
        RECT 313.950 466.950 316.050 469.050 ;
        RECT 298.800 463.950 300.900 466.050 ;
        RECT 302.100 463.950 304.200 466.050 ;
        RECT 307.950 463.950 310.050 466.050 ;
        RECT 308.400 457.050 309.600 463.950 ;
        RECT 314.400 457.200 315.600 466.950 ;
        RECT 316.950 460.050 319.050 463.050 ;
        RECT 316.950 459.000 319.200 460.050 ;
        RECT 317.100 457.950 319.200 459.000 ;
        RECT 307.800 454.950 309.900 457.050 ;
        RECT 313.800 455.100 315.900 457.200 ;
        RECT 293.400 452.400 298.050 454.050 ;
        RECT 294.000 451.950 298.050 452.400 ;
        RECT 311.100 453.600 315.000 454.050 ;
        RECT 311.100 451.950 315.600 453.600 ;
        RECT 304.950 442.950 307.050 445.050 ;
        RECT 289.950 430.950 292.050 433.050 ;
        RECT 295.950 424.950 298.050 427.050 ;
        RECT 286.950 421.950 289.050 424.050 ;
        RECT 283.950 415.950 286.050 418.050 ;
        RECT 280.950 406.950 283.050 409.050 ;
        RECT 271.950 397.950 274.050 400.050 ;
        RECT 277.950 397.950 280.050 400.050 ;
        RECT 274.950 382.950 277.050 385.050 ;
        RECT 269.400 380.400 274.050 382.050 ;
        RECT 270.000 379.950 274.050 380.400 ;
        RECT 265.950 376.950 268.050 379.050 ;
        RECT 275.400 378.600 276.600 382.950 ;
        RECT 272.400 377.400 276.600 378.600 ;
        RECT 262.950 355.950 265.050 358.050 ;
        RECT 266.400 349.050 267.600 376.950 ;
        RECT 265.950 346.950 268.050 349.050 ;
        RECT 266.400 337.050 267.600 346.950 ;
        RECT 272.400 343.050 273.600 377.400 ;
        RECT 278.400 375.600 279.600 397.950 ;
        RECT 280.950 388.950 283.050 391.050 ;
        RECT 281.400 379.050 282.600 388.950 ;
        RECT 280.950 376.950 283.050 379.050 ;
        RECT 284.400 376.050 285.600 415.950 ;
        RECT 287.400 379.050 288.600 421.950 ;
        RECT 290.400 414.000 291.600 414.600 ;
        RECT 289.950 409.950 292.050 414.000 ;
        RECT 290.400 388.050 291.600 409.950 ;
        RECT 292.950 406.950 295.050 409.050 ;
        RECT 289.950 385.950 292.050 388.050 ;
        RECT 286.950 376.950 289.050 379.050 ;
        RECT 293.400 376.050 294.600 406.950 ;
        RECT 296.400 391.050 297.600 424.950 ;
        RECT 305.400 421.050 306.600 442.950 ;
        RECT 314.400 442.050 315.600 451.950 ;
        RECT 313.950 439.950 316.050 442.050 ;
        RECT 317.400 426.600 318.600 457.950 ;
        RECT 319.950 451.950 322.050 454.050 ;
        RECT 320.400 430.050 321.600 451.950 ;
        RECT 319.950 427.950 322.050 430.050 ;
        RECT 323.400 427.050 324.600 478.950 ;
        RECT 326.400 469.050 327.600 481.950 ;
        RECT 325.950 466.950 328.050 469.050 ;
        RECT 335.400 463.050 336.600 511.950 ;
        RECT 337.950 505.950 340.050 508.050 ;
        RECT 338.400 490.050 339.600 505.950 ;
        RECT 337.950 487.950 340.050 490.050 ;
        RECT 334.950 460.950 337.050 463.050 ;
        RECT 327.000 456.600 331.050 457.050 ;
        RECT 326.400 454.950 331.050 456.600 ;
        RECT 326.400 430.050 327.600 454.950 ;
        RECT 334.950 439.950 337.050 442.050 ;
        RECT 325.950 427.950 328.050 430.050 ;
        RECT 314.400 425.400 318.600 426.600 ;
        RECT 314.400 424.050 315.600 425.400 ;
        RECT 322.950 424.950 325.050 427.050 ;
        RECT 313.800 421.950 315.900 424.050 ;
        RECT 304.950 418.950 307.050 421.050 ;
        RECT 314.400 412.050 315.600 421.950 ;
        RECT 325.800 415.950 327.900 418.050 ;
        RECT 329.100 415.950 331.200 418.050 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 298.950 409.950 301.050 412.050 ;
        RECT 314.400 410.400 319.050 412.050 ;
        RECT 315.000 409.950 319.050 410.400 ;
        RECT 295.950 388.950 298.050 391.050 ;
        RECT 299.400 382.050 300.600 409.950 ;
        RECT 323.400 394.050 324.600 412.950 ;
        RECT 322.950 391.950 325.050 394.050 ;
        RECT 319.950 388.950 322.050 391.050 ;
        RECT 313.950 382.950 316.050 385.050 ;
        RECT 298.950 379.950 301.050 382.050 ;
        RECT 295.950 376.950 298.050 379.050 ;
        RECT 306.000 378.600 310.050 379.050 ;
        RECT 305.400 376.950 310.050 378.600 ;
        RECT 275.400 374.400 279.600 375.600 ;
        RECT 271.950 340.950 274.050 343.050 ;
        RECT 265.950 334.950 268.050 337.050 ;
        RECT 256.950 316.950 259.050 319.050 ;
        RECT 253.950 313.950 256.050 316.050 ;
        RECT 250.950 307.950 253.050 310.050 ;
        RECT 244.950 304.950 247.050 307.050 ;
        RECT 251.400 301.050 252.600 307.950 ;
        RECT 254.400 307.050 255.600 313.950 ;
        RECT 257.400 313.050 258.600 316.950 ;
        RECT 256.950 310.950 259.050 313.050 ;
        RECT 266.400 312.600 267.600 334.950 ;
        RECT 271.950 313.950 274.050 316.050 ;
        RECT 266.400 311.400 270.600 312.600 ;
        RECT 262.950 307.950 265.050 310.050 ;
        RECT 254.100 306.600 256.200 307.050 ;
        RECT 254.100 305.400 258.600 306.600 ;
        RECT 254.100 304.950 256.200 305.400 ;
        RECT 235.950 298.950 238.050 301.050 ;
        RECT 250.950 298.950 253.050 301.050 ;
        RECT 232.950 286.950 235.050 289.050 ;
        RECT 226.950 277.950 229.050 280.050 ;
        RECT 196.950 268.950 199.050 271.050 ;
        RECT 217.950 268.950 220.050 271.050 ;
        RECT 193.950 262.950 196.050 265.050 ;
        RECT 197.400 250.050 198.600 268.950 ;
        RECT 202.950 265.950 205.050 268.050 ;
        RECT 203.400 253.050 204.600 265.950 ;
        RECT 205.950 253.950 208.050 256.050 ;
        RECT 202.950 250.950 205.050 253.050 ;
        RECT 196.950 247.950 199.050 250.050 ;
        RECT 190.950 241.950 193.050 244.050 ;
        RECT 183.000 237.600 187.050 238.050 ;
        RECT 182.400 235.950 187.050 237.600 ;
        RECT 199.950 235.950 202.050 238.050 ;
        RECT 182.400 229.050 183.600 235.950 ;
        RECT 200.400 232.050 201.600 235.950 ;
        RECT 199.950 229.950 202.050 232.050 ;
        RECT 181.950 226.950 184.050 229.050 ;
        RECT 181.950 217.950 184.050 220.050 ;
        RECT 178.950 214.950 181.050 217.050 ;
        RECT 182.400 205.050 183.600 217.950 ;
        RECT 184.800 211.950 186.900 214.050 ;
        RECT 175.950 202.950 178.050 205.050 ;
        RECT 181.950 202.950 184.050 205.050 ;
        RECT 176.400 199.050 177.600 202.950 ;
        RECT 185.400 199.050 186.600 211.950 ;
        RECT 190.950 208.950 193.050 211.050 ;
        RECT 191.400 202.050 192.600 208.950 ;
        RECT 190.950 199.950 193.050 202.050 ;
        RECT 175.800 196.950 177.900 199.050 ;
        RECT 181.800 196.950 183.900 199.050 ;
        RECT 185.100 196.950 187.200 199.050 ;
        RECT 167.400 194.400 172.050 196.050 ;
        RECT 168.000 193.950 172.050 194.400 ;
        RECT 160.950 190.950 163.050 193.050 ;
        RECT 154.950 187.950 157.050 190.050 ;
        RECT 139.950 172.950 142.050 175.050 ;
        RECT 148.950 172.950 151.050 175.050 ;
        RECT 140.400 169.050 141.600 172.950 ;
        RECT 151.950 169.950 154.050 172.050 ;
        RECT 139.950 166.950 142.050 169.050 ;
        RECT 118.950 160.950 121.050 163.050 ;
        RECT 133.950 160.950 136.050 163.050 ;
        RECT 152.400 160.050 153.600 169.950 ;
        RECT 155.400 169.050 156.600 187.950 ;
        RECT 160.950 184.950 163.050 187.050 ;
        RECT 161.400 169.050 162.600 184.950 ;
        RECT 182.400 184.050 183.600 196.950 ;
        RECT 184.950 187.950 187.050 190.050 ;
        RECT 181.950 181.950 184.050 184.050 ;
        RECT 169.950 175.950 172.050 178.050 ;
        RECT 154.950 166.950 157.050 169.050 ;
        RECT 161.100 166.950 163.200 169.050 ;
        RECT 167.100 166.950 169.200 169.050 ;
        RECT 145.950 157.950 148.050 160.050 ;
        RECT 151.950 157.950 154.050 160.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 111.000 129.600 115.050 130.050 ;
        RECT 110.400 127.950 115.050 129.600 ;
        RECT 127.950 127.950 130.050 130.050 ;
        RECT 91.800 127.050 93.900 127.200 ;
        RECT 89.400 125.400 93.900 127.050 ;
        RECT 90.000 125.100 93.900 125.400 ;
        RECT 90.000 124.950 93.000 125.100 ;
        RECT 103.800 124.950 105.900 127.050 ;
        RECT 85.950 121.950 88.050 124.050 ;
        RECT 93.000 123.600 96.900 124.050 ;
        RECT 92.400 121.950 96.900 123.600 ;
        RECT 92.400 115.050 93.600 121.950 ;
        RECT 104.400 118.050 105.600 124.950 ;
        RECT 103.950 115.950 106.050 118.050 ;
        RECT 110.400 115.050 111.600 127.950 ;
        RECT 121.950 124.950 124.050 127.050 ;
        RECT 122.400 115.050 123.600 124.950 ;
        RECT 128.400 115.050 129.600 127.950 ;
        RECT 139.950 124.950 142.050 127.050 ;
        RECT 140.400 115.050 141.600 124.950 ;
        RECT 146.400 124.050 147.600 157.950 ;
        RECT 167.400 157.050 168.600 166.950 ;
        RECT 166.950 154.950 169.050 157.050 ;
        RECT 167.400 150.600 168.600 154.950 ;
        RECT 164.400 149.400 168.600 150.600 ;
        RECT 151.950 139.950 154.050 142.050 ;
        RECT 145.950 121.950 148.050 124.050 ;
        RECT 67.950 112.950 70.050 115.050 ;
        RECT 91.950 112.950 94.050 115.050 ;
        RECT 109.950 112.950 112.050 115.050 ;
        RECT 121.950 112.950 124.050 115.050 ;
        RECT 127.950 112.950 130.050 115.050 ;
        RECT 139.800 112.950 141.900 115.050 ;
        RECT 73.950 109.950 76.050 112.050 ;
        RECT 55.950 94.950 58.050 97.050 ;
        RECT 52.800 92.100 54.900 94.200 ;
        RECT 74.400 94.050 75.600 109.950 ;
        RECT 112.950 103.950 115.050 106.050 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 89.400 97.050 90.600 100.950 ;
        RECT 113.400 100.050 114.600 103.950 ;
        RECT 112.950 97.950 115.050 100.050 ;
        RECT 88.950 94.950 91.050 97.050 ;
        RECT 100.950 94.950 103.050 97.050 ;
        RECT 73.950 91.950 76.050 94.050 ;
        RECT 95.100 91.950 97.200 94.050 ;
        RECT 55.950 90.600 58.050 91.050 ;
        RECT 47.400 90.000 58.050 90.600 ;
        RECT 46.950 89.400 58.050 90.000 ;
        RECT 46.950 85.950 49.050 89.400 ;
        RECT 55.950 88.950 58.050 89.400 ;
        RECT 95.400 88.050 96.600 91.950 ;
        RECT 94.950 85.950 97.050 88.050 ;
        RECT 40.950 82.950 43.050 85.050 ;
        RECT 52.950 82.950 55.050 85.050 ;
        RECT 82.950 82.950 85.050 85.050 ;
        RECT 25.950 76.950 28.050 79.050 ;
        RECT 26.400 58.050 27.600 76.950 ;
        RECT 31.950 64.950 34.050 67.050 ;
        RECT 25.950 55.950 28.050 58.050 ;
        RECT 32.400 55.050 33.600 64.950 ;
        RECT 37.950 61.950 40.050 64.050 ;
        RECT 32.100 52.950 34.200 55.050 ;
        RECT 13.950 46.950 16.050 52.050 ;
        RECT 32.400 49.050 33.600 52.950 ;
        RECT 38.400 52.050 39.600 61.950 ;
        RECT 46.950 52.950 49.050 55.050 ;
        RECT 37.950 49.950 40.050 52.050 ;
        RECT 31.950 46.950 34.050 49.050 ;
        RECT 25.950 40.950 28.050 43.050 ;
        RECT 19.950 25.950 22.050 28.050 ;
        RECT 20.400 22.050 21.600 25.950 ;
        RECT 26.400 22.050 27.600 40.950 ;
        RECT 47.400 31.050 48.600 52.950 ;
        RECT 53.400 52.050 54.600 82.950 ;
        RECT 79.950 58.950 82.050 61.050 ;
        RECT 70.950 57.600 75.000 58.050 ;
        RECT 70.950 55.950 75.600 57.600 ;
        RECT 60.000 54.600 64.050 55.050 ;
        RECT 59.400 52.950 64.050 54.600 ;
        RECT 52.950 49.950 55.050 52.050 ;
        RECT 59.400 43.050 60.600 52.950 ;
        RECT 67.950 43.950 70.050 46.050 ;
        RECT 58.950 40.950 61.050 43.050 ;
        RECT 46.950 28.950 49.050 31.050 ;
        RECT 43.950 25.950 46.050 28.050 ;
        RECT 49.950 25.950 52.050 28.050 ;
        RECT 44.400 22.050 45.600 25.950 ;
        RECT 19.950 19.950 22.050 22.050 ;
        RECT 26.100 19.950 28.200 22.050 ;
        RECT 43.950 19.950 46.050 22.050 ;
        RECT 50.400 13.050 51.600 25.950 ;
        RECT 68.400 22.050 69.600 43.950 ;
        RECT 64.950 20.400 69.600 22.050 ;
        RECT 64.950 19.950 69.000 20.400 ;
        RECT 74.400 19.050 75.600 55.950 ;
        RECT 80.400 49.050 81.600 58.950 ;
        RECT 83.400 55.050 84.600 82.950 ;
        RECT 91.950 79.950 94.050 82.050 ;
        RECT 83.400 53.400 88.050 55.050 ;
        RECT 84.000 52.950 88.050 53.400 ;
        RECT 79.950 46.950 82.050 49.050 ;
        RECT 92.400 43.050 93.600 79.950 ;
        RECT 101.400 70.050 102.600 94.950 ;
        RECT 113.400 94.050 114.600 97.950 ;
        RECT 128.400 94.050 129.600 112.950 ;
        RECT 152.400 109.050 153.600 139.950 ;
        RECT 157.800 121.950 159.900 124.050 ;
        RECT 158.400 115.050 159.600 121.950 ;
        RECT 157.950 112.950 160.050 115.050 ;
        RECT 136.950 106.950 139.050 109.050 ;
        RECT 151.950 106.950 154.050 109.050 ;
        RECT 109.950 92.400 114.600 94.050 ;
        RECT 109.950 91.950 114.000 92.400 ;
        RECT 127.950 91.950 130.050 94.050 ;
        RECT 103.950 88.950 106.050 91.050 ;
        RECT 94.950 67.950 97.050 70.050 ;
        RECT 100.950 67.950 103.050 70.050 ;
        RECT 95.400 49.050 96.600 67.950 ;
        RECT 104.400 64.050 105.600 88.950 ;
        RECT 128.400 88.050 129.600 91.950 ;
        RECT 127.950 85.950 130.050 88.050 ;
        RECT 118.950 73.950 121.050 76.050 ;
        RECT 109.800 64.950 111.900 67.050 ;
        RECT 103.950 61.950 106.050 64.050 ;
        RECT 101.100 54.600 105.000 55.050 ;
        RECT 101.100 52.950 105.600 54.600 ;
        RECT 98.100 49.950 100.200 52.050 ;
        RECT 94.800 46.950 96.900 49.050 ;
        RECT 91.950 40.950 94.050 43.050 ;
        RECT 76.950 37.950 79.050 40.050 ;
        RECT 77.400 31.050 78.600 37.950 ;
        RECT 76.950 28.950 79.050 31.050 ;
        RECT 77.400 22.050 78.600 28.950 ;
        RECT 82.950 22.950 85.050 25.050 ;
        RECT 76.950 19.950 79.050 22.050 ;
        RECT 73.950 16.950 76.050 19.050 ;
        RECT 49.950 10.950 52.050 13.050 ;
        RECT 83.400 10.050 84.600 22.950 ;
        RECT 92.400 22.050 93.600 40.950 ;
        RECT 98.400 28.050 99.600 49.950 ;
        RECT 104.400 43.050 105.600 52.950 ;
        RECT 110.400 52.050 111.600 64.950 ;
        RECT 119.400 58.050 120.600 73.950 ;
        RECT 133.950 70.950 136.050 73.050 ;
        RECT 124.950 61.950 127.050 64.050 ;
        RECT 118.950 55.950 121.050 58.050 ;
        RECT 125.400 55.050 126.600 61.950 ;
        RECT 125.400 53.400 130.050 55.050 ;
        RECT 126.000 52.950 130.050 53.400 ;
        RECT 134.400 52.050 135.600 70.950 ;
        RECT 110.100 49.950 112.200 52.050 ;
        RECT 133.950 49.950 136.050 52.050 ;
        RECT 118.950 43.950 121.050 46.050 ;
        RECT 103.950 40.950 106.050 43.050 ;
        RECT 97.950 25.950 100.050 28.050 ;
        RECT 106.950 22.950 109.050 28.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 92.400 20.400 97.050 22.050 ;
        RECT 93.000 19.950 97.050 20.400 ;
        RECT 113.400 13.050 114.600 22.950 ;
        RECT 119.400 19.050 120.600 43.950 ;
        RECT 137.400 37.050 138.600 106.950 ;
        RECT 148.950 103.950 151.050 106.050 ;
        RECT 149.400 94.050 150.600 103.950 ;
        RECT 160.950 97.950 163.050 103.050 ;
        RECT 149.100 91.950 151.200 94.050 ;
        RECT 157.950 82.950 160.050 85.050 ;
        RECT 158.400 58.050 159.600 82.950 ;
        RECT 164.400 82.050 165.600 149.400 ;
        RECT 170.400 124.050 171.600 175.950 ;
        RECT 178.950 172.950 181.050 175.050 ;
        RECT 179.400 166.050 180.600 172.950 ;
        RECT 175.950 164.400 180.600 166.050 ;
        RECT 175.950 163.950 180.000 164.400 ;
        RECT 182.100 163.950 184.200 166.050 ;
        RECT 172.950 160.950 175.050 163.050 ;
        RECT 173.400 142.050 174.600 160.950 ;
        RECT 182.400 154.050 183.600 163.950 ;
        RECT 181.950 151.950 184.050 154.050 ;
        RECT 172.950 139.950 175.050 142.050 ;
        RECT 178.950 130.950 181.050 133.050 ;
        RECT 179.400 124.050 180.600 130.950 ;
        RECT 169.800 121.950 171.900 124.050 ;
        RECT 179.400 122.400 184.050 124.050 ;
        RECT 180.000 121.950 184.050 122.400 ;
        RECT 170.400 103.050 171.600 121.950 ;
        RECT 172.950 112.950 175.050 115.050 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 173.400 94.050 174.600 112.950 ;
        RECT 185.400 106.050 186.600 187.950 ;
        RECT 193.950 181.950 196.050 184.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 188.400 127.050 189.600 178.950 ;
        RECT 194.400 163.050 195.600 181.950 ;
        RECT 206.400 178.050 207.600 253.950 ;
        RECT 218.400 244.050 219.600 268.950 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 217.950 241.950 220.050 244.050 ;
        RECT 211.950 238.950 214.050 241.050 ;
        RECT 221.100 238.950 223.200 241.050 ;
        RECT 212.400 229.050 213.600 238.950 ;
        RECT 217.950 235.950 220.050 238.050 ;
        RECT 218.400 232.050 219.600 235.950 ;
        RECT 217.950 229.950 220.050 232.050 ;
        RECT 211.950 226.950 214.050 229.050 ;
        RECT 221.400 223.050 222.600 238.950 ;
        RECT 224.400 235.050 225.600 256.950 ;
        RECT 223.950 232.950 226.050 235.050 ;
        RECT 220.950 220.950 223.050 223.050 ;
        RECT 211.950 214.950 214.050 217.050 ;
        RECT 212.400 202.050 213.600 214.950 ;
        RECT 227.400 211.050 228.600 277.950 ;
        RECT 229.950 265.950 232.050 268.050 ;
        RECT 230.400 214.050 231.600 265.950 ;
        RECT 236.400 247.200 237.600 298.950 ;
        RECT 253.950 292.950 256.050 295.050 ;
        RECT 254.400 277.050 255.600 292.950 ;
        RECT 253.950 274.950 256.050 277.050 ;
        RECT 244.950 268.950 247.050 271.050 ;
        RECT 245.400 256.050 246.600 268.950 ;
        RECT 257.400 258.600 258.600 305.400 ;
        RECT 259.950 280.950 262.050 283.050 ;
        RECT 260.400 277.050 261.600 280.950 ;
        RECT 263.400 280.050 264.600 307.950 ;
        RECT 269.400 292.050 270.600 311.400 ;
        RECT 268.950 289.950 271.050 292.050 ;
        RECT 272.400 280.050 273.600 313.950 ;
        RECT 275.400 310.050 276.600 374.400 ;
        RECT 283.950 373.950 286.050 376.050 ;
        RECT 292.950 373.950 295.050 376.050 ;
        RECT 284.400 361.050 285.600 373.950 ;
        RECT 283.950 358.950 286.050 361.050 ;
        RECT 296.400 346.050 297.600 376.950 ;
        RECT 305.400 370.050 306.600 376.950 ;
        RECT 314.400 376.050 315.600 382.950 ;
        RECT 320.400 382.050 321.600 388.950 ;
        RECT 326.400 385.050 327.600 415.950 ;
        RECT 329.400 406.050 330.600 415.950 ;
        RECT 328.950 403.950 331.050 406.050 ;
        RECT 335.400 391.050 336.600 439.950 ;
        RECT 338.400 424.050 339.600 487.950 ;
        RECT 341.400 427.050 342.600 526.950 ;
        RECT 352.950 523.800 355.050 525.900 ;
        RECT 343.950 514.950 346.050 517.050 ;
        RECT 344.400 511.050 345.600 514.950 ;
        RECT 343.950 508.950 346.050 511.050 ;
        RECT 343.950 499.950 346.050 502.050 ;
        RECT 344.400 490.050 345.600 499.950 ;
        RECT 343.800 489.000 345.900 490.050 ;
        RECT 343.800 487.950 346.050 489.000 ;
        RECT 343.950 486.000 346.050 487.950 ;
        RECT 344.400 485.400 345.600 486.000 ;
        RECT 349.950 484.950 352.050 487.050 ;
        RECT 350.400 475.050 351.600 484.950 ;
        RECT 353.400 478.050 354.600 523.800 ;
        RECT 356.400 481.050 357.600 547.950 ;
        RECT 361.950 535.950 364.050 538.050 ;
        RECT 362.400 523.050 363.600 535.950 ;
        RECT 364.950 523.950 367.050 526.050 ;
        RECT 361.950 520.950 364.050 523.050 ;
        RECT 365.400 496.050 366.600 523.950 ;
        RECT 368.400 499.050 369.600 554.400 ;
        RECT 370.950 550.950 373.050 553.050 ;
        RECT 367.950 496.950 370.050 499.050 ;
        RECT 364.950 493.950 367.050 496.050 ;
        RECT 361.950 481.950 364.050 484.050 ;
        RECT 355.950 478.950 358.050 481.050 ;
        RECT 362.400 478.050 363.600 481.950 ;
        RECT 352.950 475.950 355.050 478.050 ;
        RECT 361.950 475.950 364.050 478.050 ;
        RECT 349.950 472.950 352.050 475.050 ;
        RECT 355.950 472.950 358.050 475.050 ;
        RECT 346.950 469.950 349.050 472.050 ;
        RECT 347.400 457.050 348.600 469.950 ;
        RECT 352.950 460.950 355.050 463.050 ;
        RECT 353.400 457.050 354.600 460.950 ;
        RECT 356.400 457.050 357.600 472.950 ;
        RECT 361.950 466.950 364.050 469.050 ;
        RECT 343.950 455.400 348.600 457.050 ;
        RECT 343.950 454.950 348.000 455.400 ;
        RECT 352.800 454.950 354.900 457.050 ;
        RECT 356.400 454.950 361.050 457.050 ;
        RECT 343.950 448.950 346.050 451.050 ;
        RECT 344.400 442.050 345.600 448.950 ;
        RECT 343.950 439.950 346.050 442.050 ;
        RECT 340.950 424.950 343.050 427.050 ;
        RECT 337.950 421.950 340.050 424.050 ;
        RECT 341.400 408.600 342.600 424.950 ;
        RECT 338.400 407.400 342.600 408.600 ;
        RECT 334.950 388.950 337.050 391.050 ;
        RECT 328.950 385.950 331.050 388.050 ;
        RECT 326.100 382.950 328.200 385.050 ;
        RECT 320.400 379.950 324.900 382.050 ;
        RECT 313.950 373.950 316.050 376.050 ;
        RECT 304.950 367.950 307.050 370.050 ;
        RECT 298.950 349.950 301.050 352.050 ;
        RECT 299.400 346.050 300.600 349.950 ;
        RECT 295.800 343.950 297.900 346.050 ;
        RECT 299.100 343.950 301.200 346.050 ;
        RECT 307.950 343.950 310.050 346.050 ;
        RECT 289.950 340.950 292.050 343.050 ;
        RECT 277.800 337.950 279.900 340.050 ;
        RECT 282.000 339.600 285.900 340.050 ;
        RECT 281.400 337.950 285.900 339.600 ;
        RECT 278.400 331.050 279.600 337.950 ;
        RECT 277.950 328.950 280.050 331.050 ;
        RECT 281.400 316.050 282.600 337.950 ;
        RECT 283.950 319.950 286.050 322.050 ;
        RECT 280.950 313.950 283.050 316.050 ;
        RECT 284.400 313.050 285.600 319.950 ;
        RECT 283.950 310.950 286.050 313.050 ;
        RECT 274.800 307.950 276.900 310.050 ;
        RECT 290.400 286.050 291.600 340.950 ;
        RECT 308.400 340.050 309.600 343.950 ;
        RECT 292.950 339.600 297.000 340.050 ;
        RECT 292.950 337.950 297.600 339.600 ;
        RECT 307.950 337.950 310.050 340.050 ;
        RECT 296.400 325.050 297.600 337.950 ;
        RECT 295.950 322.950 298.050 325.050 ;
        RECT 301.950 319.950 304.050 322.050 ;
        RECT 302.400 310.050 303.600 319.950 ;
        RECT 302.400 308.400 307.050 310.050 ;
        RECT 303.000 307.950 307.050 308.400 ;
        RECT 294.000 306.600 297.900 307.050 ;
        RECT 293.400 304.950 297.900 306.600 ;
        RECT 289.950 283.950 292.050 286.050 ;
        RECT 293.400 283.050 294.600 304.950 ;
        RECT 298.950 298.950 301.050 301.050 ;
        RECT 299.400 283.050 300.600 298.950 ;
        RECT 308.400 289.050 309.600 337.950 ;
        RECT 314.400 336.600 315.600 373.950 ;
        RECT 320.400 352.050 321.600 379.950 ;
        RECT 322.950 373.950 325.050 376.050 ;
        RECT 319.950 349.950 322.050 352.050 ;
        RECT 311.400 335.400 315.600 336.600 ;
        RECT 311.400 325.050 312.600 335.400 ;
        RECT 310.950 322.950 313.050 325.050 ;
        RECT 311.400 316.050 312.600 322.950 ;
        RECT 313.950 316.950 316.050 319.050 ;
        RECT 310.950 313.950 313.050 316.050 ;
        RECT 314.400 307.050 315.600 316.950 ;
        RECT 316.950 313.950 319.050 316.050 ;
        RECT 313.950 304.950 316.050 307.050 ;
        RECT 317.400 304.050 318.600 313.950 ;
        RECT 319.950 304.050 322.050 307.050 ;
        RECT 316.800 301.950 318.900 304.050 ;
        RECT 319.950 303.000 322.200 304.050 ;
        RECT 320.100 301.950 322.200 303.000 ;
        RECT 310.950 292.950 313.050 295.050 ;
        RECT 307.950 286.950 310.050 289.050 ;
        RECT 292.950 280.950 295.050 283.050 ;
        RECT 298.950 280.950 301.050 283.050 ;
        RECT 262.800 277.950 264.900 280.050 ;
        RECT 271.950 277.950 274.050 280.050 ;
        RECT 259.950 274.950 262.050 277.050 ;
        RECT 260.400 268.050 261.600 274.950 ;
        RECT 280.950 271.950 283.050 274.050 ;
        RECT 268.950 268.950 271.050 271.050 ;
        RECT 259.950 265.950 262.050 268.050 ;
        RECT 259.950 259.950 262.050 262.050 ;
        RECT 254.400 257.400 258.600 258.600 ;
        RECT 244.950 253.950 247.050 256.050 ;
        RECT 241.950 250.950 244.050 253.050 ;
        RECT 235.950 245.100 238.050 247.200 ;
        RECT 235.950 241.800 238.050 243.900 ;
        RECT 236.400 238.050 237.600 241.800 ;
        RECT 242.400 238.050 243.600 250.950 ;
        RECT 247.950 247.950 250.050 250.050 ;
        RECT 248.400 238.050 249.600 247.950 ;
        RECT 254.400 247.050 255.600 257.400 ;
        RECT 253.950 244.950 256.050 247.050 ;
        RECT 235.950 235.950 238.050 238.050 ;
        RECT 241.800 235.950 243.900 238.050 ;
        RECT 247.950 235.950 250.050 238.050 ;
        RECT 256.950 235.950 259.050 238.050 ;
        RECT 257.400 229.050 258.600 235.950 ;
        RECT 256.950 226.950 259.050 229.050 ;
        RECT 235.950 223.950 238.050 226.050 ;
        RECT 229.950 211.950 232.050 214.050 ;
        RECT 226.950 208.950 229.050 211.050 ;
        RECT 227.400 207.600 228.600 208.950 ;
        RECT 227.400 206.400 231.600 207.600 ;
        RECT 230.400 202.050 231.600 206.400 ;
        RECT 211.950 199.950 214.050 202.050 ;
        RECT 229.950 199.950 232.050 202.050 ;
        RECT 226.950 196.950 229.050 199.050 ;
        RECT 205.950 175.950 208.050 178.050 ;
        RECT 202.950 169.950 205.050 175.050 ;
        RECT 217.950 169.950 220.050 172.050 ;
        RECT 196.950 163.950 199.050 166.050 ;
        RECT 193.950 160.950 196.050 163.050 ;
        RECT 197.400 160.050 198.600 163.950 ;
        RECT 218.400 163.050 219.600 169.950 ;
        RECT 205.950 160.950 208.050 163.050 ;
        RECT 217.950 160.950 220.050 163.050 ;
        RECT 196.950 157.950 199.050 160.050 ;
        RECT 206.400 154.050 207.600 160.950 ;
        RECT 205.950 151.950 208.050 154.050 ;
        RECT 196.950 136.950 199.050 139.050 ;
        RECT 197.400 130.050 198.600 136.950 ;
        RECT 196.950 127.950 199.050 130.050 ;
        RECT 202.950 127.950 205.050 130.050 ;
        RECT 187.800 124.950 189.900 127.050 ;
        RECT 190.800 121.950 192.900 124.050 ;
        RECT 191.400 118.050 192.600 121.950 ;
        RECT 196.950 118.950 199.050 121.050 ;
        RECT 190.950 115.950 193.050 118.050 ;
        RECT 197.400 109.050 198.600 118.950 ;
        RECT 196.950 106.950 199.050 109.050 ;
        RECT 184.950 103.950 187.050 106.050 ;
        RECT 181.950 100.950 184.050 103.050 ;
        RECT 182.400 94.050 183.600 100.950 ;
        RECT 187.950 94.950 190.050 97.050 ;
        RECT 173.400 92.400 177.900 94.050 ;
        RECT 174.000 91.950 177.900 92.400 ;
        RECT 181.950 91.950 184.050 94.050 ;
        RECT 163.950 79.950 166.050 82.050 ;
        RECT 169.950 79.950 172.050 82.050 ;
        RECT 170.400 61.050 171.600 79.950 ;
        RECT 178.950 70.950 181.050 73.050 ;
        RECT 157.950 55.950 160.050 58.050 ;
        RECT 163.950 55.950 166.050 61.050 ;
        RECT 169.800 58.950 171.900 61.050 ;
        RECT 179.400 55.050 180.600 70.950 ;
        RECT 188.400 70.050 189.600 94.950 ;
        RECT 197.400 93.600 198.600 106.950 ;
        RECT 203.400 100.050 204.600 127.950 ;
        RECT 217.800 124.950 219.900 127.050 ;
        RECT 223.950 124.950 226.050 127.050 ;
        RECT 218.400 106.050 219.600 124.950 ;
        RECT 224.400 115.050 225.600 124.950 ;
        RECT 227.400 121.050 228.600 196.950 ;
        RECT 236.400 181.200 237.600 223.950 ;
        RECT 260.400 208.050 261.600 259.950 ;
        RECT 262.950 244.950 265.050 247.050 ;
        RECT 259.950 205.950 262.050 208.050 ;
        RECT 263.400 202.050 264.600 244.950 ;
        RECT 265.950 232.950 268.050 235.050 ;
        RECT 262.950 199.950 265.050 202.050 ;
        RECT 244.950 196.950 247.050 199.050 ;
        RECT 235.950 179.100 238.050 181.200 ;
        RECT 235.950 175.800 238.050 177.900 ;
        RECT 232.950 157.950 235.050 160.050 ;
        RECT 233.400 142.050 234.600 157.950 ;
        RECT 232.950 139.950 235.050 142.050 ;
        RECT 236.400 133.050 237.600 175.800 ;
        RECT 238.800 160.950 240.900 163.050 ;
        RECT 239.400 157.050 240.600 160.950 ;
        RECT 238.950 154.950 241.050 157.050 ;
        RECT 235.950 130.950 238.050 133.050 ;
        RECT 236.400 124.050 237.600 130.950 ;
        RECT 245.400 130.050 246.600 196.950 ;
        RECT 253.950 193.800 256.050 195.900 ;
        RECT 250.950 187.950 253.050 190.050 ;
        RECT 251.400 175.050 252.600 187.950 ;
        RECT 250.950 172.950 253.050 175.050 ;
        RECT 254.400 172.050 255.600 193.800 ;
        RECT 263.400 193.050 264.600 199.950 ;
        RECT 266.400 198.600 267.600 232.950 ;
        RECT 269.400 220.050 270.600 268.950 ;
        RECT 281.400 265.050 282.600 271.950 ;
        RECT 311.400 271.050 312.600 292.950 ;
        RECT 316.950 286.950 319.050 289.050 ;
        RECT 289.950 268.950 292.050 271.050 ;
        RECT 299.100 270.000 301.200 271.050 ;
        RECT 298.950 268.950 301.200 270.000 ;
        RECT 310.950 268.950 313.050 271.050 ;
        RECT 280.800 264.000 282.900 265.050 ;
        RECT 280.800 262.950 283.050 264.000 ;
        RECT 280.950 259.950 283.050 262.950 ;
        RECT 290.400 259.050 291.600 268.950 ;
        RECT 298.950 265.950 301.050 268.950 ;
        RECT 289.950 256.950 292.050 259.050 ;
        RECT 310.950 256.950 313.050 259.050 ;
        RECT 283.950 250.950 286.050 253.050 ;
        RECT 280.950 238.950 283.050 244.050 ;
        RECT 284.400 232.050 285.600 250.950 ;
        RECT 286.950 247.950 289.050 250.050 ;
        RECT 287.400 241.050 288.600 247.950 ;
        RECT 290.400 244.050 291.600 256.950 ;
        RECT 307.950 250.950 310.050 253.050 ;
        RECT 289.950 241.950 292.050 244.050 ;
        RECT 286.950 238.950 289.050 241.050 ;
        RECT 301.950 240.600 306.000 241.050 ;
        RECT 301.950 238.950 306.600 240.600 ;
        RECT 295.950 235.950 298.050 238.050 ;
        RECT 283.950 229.950 286.050 232.050 ;
        RECT 277.950 223.950 280.050 226.050 ;
        RECT 268.950 217.950 271.050 220.050 ;
        RECT 274.950 205.950 277.050 208.050 ;
        RECT 268.950 198.600 271.050 199.050 ;
        RECT 266.400 197.400 271.050 198.600 ;
        RECT 268.950 196.950 271.050 197.400 ;
        RECT 263.100 190.950 265.200 193.050 ;
        RECT 269.400 187.050 270.600 196.950 ;
        RECT 259.950 184.950 262.050 187.050 ;
        RECT 268.800 184.950 270.900 187.050 ;
        RECT 253.950 169.950 256.050 172.050 ;
        RECT 260.400 169.050 261.600 184.950 ;
        RECT 275.400 175.050 276.600 205.950 ;
        RECT 278.400 178.050 279.600 223.950 ;
        RECT 296.400 223.050 297.600 235.950 ;
        RECT 305.400 235.050 306.600 238.950 ;
        RECT 304.950 232.950 307.050 235.050 ;
        RECT 308.400 226.050 309.600 250.950 ;
        RECT 307.950 223.950 310.050 226.050 ;
        RECT 295.950 220.950 298.050 223.050 ;
        RECT 311.400 202.050 312.600 256.950 ;
        RECT 317.400 205.050 318.600 286.950 ;
        RECT 320.400 244.050 321.600 301.950 ;
        RECT 323.400 286.050 324.600 373.950 ;
        RECT 329.400 370.050 330.600 385.950 ;
        RECT 328.950 367.950 331.050 370.050 ;
        RECT 325.950 349.950 328.050 352.050 ;
        RECT 326.400 346.050 327.600 349.950 ;
        RECT 328.950 346.050 331.050 346.200 ;
        RECT 326.400 344.550 331.050 346.050 ;
        RECT 327.000 344.100 331.050 344.550 ;
        RECT 327.000 343.950 330.000 344.100 ;
        RECT 328.950 340.800 331.050 342.900 ;
        RECT 322.950 283.950 325.050 286.050 ;
        RECT 322.950 277.950 325.050 280.050 ;
        RECT 323.400 268.050 324.600 277.950 ;
        RECT 329.400 271.050 330.600 340.800 ;
        RECT 334.950 328.950 337.050 331.050 ;
        RECT 335.400 307.050 336.600 328.950 ;
        RECT 338.400 319.050 339.600 407.400 ;
        RECT 340.950 403.950 343.050 406.050 ;
        RECT 341.400 388.050 342.600 403.950 ;
        RECT 340.950 385.950 343.050 388.050 ;
        RECT 344.400 376.050 345.600 439.950 ;
        RECT 346.950 436.950 349.050 439.050 ;
        RECT 347.400 433.050 348.600 436.950 ;
        RECT 346.950 430.950 349.050 433.050 ;
        RECT 347.400 412.050 348.600 430.950 ;
        RECT 352.950 427.950 355.050 430.050 ;
        RECT 353.400 412.050 354.600 427.950 ;
        RECT 356.400 418.050 357.600 454.950 ;
        RECT 358.950 445.950 361.050 448.050 ;
        RECT 355.950 415.950 358.050 418.050 ;
        RECT 346.950 409.950 349.050 412.050 ;
        RECT 353.400 409.950 358.050 412.050 ;
        RECT 347.400 400.050 348.600 409.950 ;
        RECT 346.950 397.950 349.050 400.050 ;
        RECT 353.400 394.050 354.600 409.950 ;
        RECT 359.400 406.050 360.600 445.950 ;
        RECT 358.950 403.950 361.050 406.050 ;
        RECT 352.950 393.600 355.050 394.050 ;
        RECT 350.400 392.400 355.050 393.600 ;
        RECT 346.950 385.950 349.050 388.050 ;
        RECT 347.400 382.050 348.600 385.950 ;
        RECT 346.950 379.950 349.050 382.050 ;
        RECT 343.950 373.950 346.050 376.050 ;
        RECT 347.400 363.600 348.600 379.950 ;
        RECT 344.400 362.400 348.600 363.600 ;
        RECT 344.400 340.050 345.600 362.400 ;
        RECT 350.400 340.050 351.600 392.400 ;
        RECT 352.950 391.950 355.050 392.400 ;
        RECT 362.400 385.050 363.600 466.950 ;
        RECT 365.400 463.050 366.600 493.950 ;
        RECT 368.400 469.050 369.600 496.950 ;
        RECT 367.950 466.950 370.050 469.050 ;
        RECT 371.400 466.050 372.600 550.950 ;
        RECT 374.400 535.050 375.600 593.400 ;
        RECT 380.400 577.050 381.600 596.400 ;
        RECT 385.950 595.950 388.050 598.050 ;
        RECT 386.400 577.050 387.600 595.950 ;
        RECT 379.950 574.950 382.050 577.050 ;
        RECT 385.950 574.950 388.050 577.050 ;
        RECT 376.950 568.950 379.050 571.050 ;
        RECT 377.400 562.050 378.600 568.950 ;
        RECT 392.400 562.050 393.600 610.950 ;
        RECT 398.400 610.050 399.600 625.950 ;
        RECT 407.400 625.050 408.600 628.950 ;
        RECT 413.400 628.050 414.600 682.950 ;
        RECT 419.400 670.050 420.600 697.950 ;
        RECT 431.400 691.050 432.600 724.950 ;
        RECT 437.400 721.050 438.600 739.950 ;
        RECT 443.400 727.050 444.600 769.950 ;
        RECT 446.100 744.600 450.000 745.050 ;
        RECT 446.100 742.950 450.600 744.600 ;
        RECT 449.400 730.050 450.600 742.950 ;
        RECT 457.950 733.950 460.050 736.050 ;
        RECT 454.950 730.950 457.050 733.050 ;
        RECT 448.950 727.950 451.050 730.050 ;
        RECT 442.950 724.950 445.050 727.050 ;
        RECT 439.950 721.950 442.050 724.050 ;
        RECT 436.950 718.950 439.050 721.050 ;
        RECT 437.400 703.050 438.600 718.950 ;
        RECT 440.400 712.050 441.600 721.950 ;
        RECT 439.950 709.950 442.050 712.050 ;
        RECT 451.950 706.950 454.050 709.050 ;
        RECT 445.950 703.950 448.050 706.050 ;
        RECT 436.950 700.950 439.050 703.050 ;
        RECT 446.400 700.050 447.600 703.950 ;
        RECT 445.950 699.600 450.000 700.050 ;
        RECT 445.950 697.950 450.600 699.600 ;
        RECT 436.950 694.950 439.050 697.050 ;
        RECT 430.950 688.950 433.050 691.050 ;
        RECT 437.400 682.050 438.600 694.950 ;
        RECT 439.950 688.950 442.050 691.050 ;
        RECT 436.950 679.950 439.050 682.050 ;
        RECT 437.400 676.050 438.600 679.950 ;
        RECT 436.800 673.950 438.900 676.050 ;
        RECT 415.950 668.400 420.600 670.050 ;
        RECT 415.950 667.950 420.000 668.400 ;
        RECT 424.950 664.950 427.050 667.050 ;
        RECT 425.400 661.050 426.600 664.950 ;
        RECT 424.950 658.950 427.050 661.050 ;
        RECT 425.400 640.050 426.600 658.950 ;
        RECT 430.950 652.950 433.050 655.050 ;
        RECT 424.950 637.950 427.050 640.050 ;
        RECT 413.100 625.950 415.200 628.050 ;
        RECT 418.800 625.950 420.900 628.050 ;
        RECT 406.950 622.950 409.050 625.050 ;
        RECT 419.400 610.050 420.600 625.950 ;
        RECT 431.400 625.050 432.600 652.950 ;
        RECT 440.400 634.050 441.600 688.950 ;
        RECT 445.950 682.950 448.050 685.050 ;
        RECT 446.400 679.050 447.600 682.950 ;
        RECT 445.950 676.950 448.050 679.050 ;
        RECT 449.400 676.050 450.600 697.950 ;
        RECT 452.400 697.050 453.600 706.950 ;
        RECT 451.950 694.950 454.050 697.050 ;
        RECT 455.400 676.050 456.600 730.950 ;
        RECT 458.400 721.050 459.600 733.950 ;
        RECT 457.950 718.950 460.050 721.050 ;
        RECT 461.400 679.050 462.600 802.950 ;
        RECT 467.400 772.050 468.600 811.950 ;
        RECT 470.400 802.050 471.600 841.950 ;
        RECT 476.400 817.050 477.600 844.950 ;
        RECT 485.400 835.050 486.600 850.950 ;
        RECT 511.950 847.950 514.050 850.050 ;
        RECT 512.400 844.050 513.600 847.950 ;
        RECT 575.400 847.050 576.600 850.950 ;
        RECT 526.950 844.950 529.050 847.050 ;
        RECT 562.950 844.950 565.050 847.050 ;
        RECT 574.950 844.950 577.050 847.050 ;
        RECT 511.950 841.950 514.050 844.050 ;
        RECT 484.950 832.950 487.050 835.050 ;
        RECT 512.400 829.050 513.600 841.950 ;
        RECT 517.950 835.950 520.050 838.050 ;
        RECT 508.800 826.950 510.900 829.050 ;
        RECT 512.100 826.950 514.200 829.050 ;
        RECT 502.950 820.950 505.050 823.050 ;
        RECT 484.950 817.950 487.050 820.050 ;
        RECT 475.950 814.950 478.050 817.050 ;
        RECT 485.400 811.050 486.600 817.950 ;
        RECT 503.400 817.050 504.600 820.950 ;
        RECT 505.950 817.950 508.050 820.050 ;
        RECT 502.800 814.950 504.900 817.050 ;
        RECT 478.950 808.950 481.050 811.050 ;
        RECT 485.100 808.950 487.200 811.050 ;
        RECT 469.950 799.950 472.050 802.050 ;
        RECT 479.400 799.050 480.600 808.950 ;
        RECT 478.950 796.950 481.050 799.050 ;
        RECT 506.400 784.050 507.600 817.950 ;
        RECT 505.950 781.950 508.050 784.050 ;
        RECT 478.950 775.950 481.050 778.050 ;
        RECT 493.950 775.950 496.050 778.050 ;
        RECT 466.950 769.950 469.050 772.050 ;
        RECT 469.950 757.950 472.050 760.050 ;
        RECT 463.950 733.950 466.050 736.050 ;
        RECT 464.400 703.050 465.600 733.950 ;
        RECT 470.400 732.600 471.600 757.950 ;
        RECT 467.400 731.400 471.600 732.600 ;
        RECT 467.400 706.050 468.600 731.400 ;
        RECT 472.950 727.950 475.050 730.050 ;
        RECT 466.950 703.950 469.050 706.050 ;
        RECT 463.950 700.950 466.050 703.050 ;
        RECT 473.400 697.050 474.600 727.950 ;
        RECT 479.400 709.050 480.600 775.950 ;
        RECT 484.950 772.950 487.050 775.050 ;
        RECT 485.400 769.050 486.600 772.950 ;
        RECT 494.400 772.050 495.600 775.950 ;
        RECT 499.950 774.600 504.000 775.050 ;
        RECT 499.950 772.950 504.600 774.600 ;
        RECT 493.950 769.950 496.050 772.050 ;
        RECT 484.950 766.950 487.050 769.050 ;
        RECT 485.400 745.050 486.600 766.950 ;
        RECT 484.800 742.950 486.900 745.050 ;
        RECT 481.950 724.950 484.050 727.050 ;
        RECT 482.400 718.050 483.600 724.950 ;
        RECT 484.950 718.950 487.050 721.050 ;
        RECT 481.950 715.950 484.050 718.050 ;
        RECT 478.950 706.950 481.050 709.050 ;
        RECT 485.400 706.050 486.600 718.950 ;
        RECT 494.400 709.050 495.600 769.950 ;
        RECT 503.400 769.050 504.600 772.950 ;
        RECT 509.400 772.050 510.600 826.950 ;
        RECT 514.950 820.950 517.050 823.050 ;
        RECT 511.950 817.950 514.050 820.050 ;
        RECT 512.400 799.050 513.600 817.950 ;
        RECT 515.400 811.050 516.600 820.950 ;
        RECT 514.950 808.950 517.050 811.050 ;
        RECT 511.950 796.950 514.050 799.050 ;
        RECT 518.400 772.050 519.600 835.950 ;
        RECT 527.400 805.050 528.600 844.950 ;
        RECT 563.400 838.050 564.600 844.950 ;
        RECT 568.950 838.950 571.050 841.050 ;
        RECT 553.950 835.950 556.050 838.050 ;
        RECT 562.950 835.950 565.050 838.050 ;
        RECT 532.950 811.950 535.050 814.050 ;
        RECT 545.100 813.600 549.000 814.050 ;
        RECT 545.100 811.950 549.600 813.600 ;
        RECT 526.950 802.950 529.050 805.050 ;
        RECT 527.400 778.050 528.600 802.950 ;
        RECT 533.400 802.050 534.600 811.950 ;
        RECT 548.400 805.050 549.600 811.950 ;
        RECT 547.950 802.950 550.050 805.050 ;
        RECT 532.950 799.950 535.050 802.050 ;
        RECT 526.950 775.950 529.050 778.050 ;
        RECT 509.100 769.950 511.200 772.050 ;
        RECT 517.950 769.950 520.050 772.050 ;
        RECT 502.950 766.950 505.050 769.050 ;
        RECT 514.950 766.950 517.050 769.050 ;
        RECT 502.950 760.950 505.050 763.050 ;
        RECT 503.400 751.050 504.600 760.950 ;
        RECT 515.400 757.050 516.600 766.950 ;
        RECT 514.950 754.950 517.050 757.050 ;
        RECT 502.950 748.950 505.050 751.050 ;
        RECT 508.950 748.950 511.050 751.050 ;
        RECT 509.400 745.050 510.600 748.950 ;
        RECT 508.950 742.950 511.050 745.050 ;
        RECT 502.950 739.950 505.050 742.050 ;
        RECT 487.950 706.950 490.050 709.050 ;
        RECT 493.950 706.950 496.050 709.050 ;
        RECT 475.950 703.950 478.050 706.050 ;
        RECT 481.950 704.400 486.600 706.050 ;
        RECT 481.950 703.950 486.000 704.400 ;
        RECT 469.950 695.400 474.600 697.050 ;
        RECT 469.950 694.950 474.000 695.400 ;
        RECT 460.950 676.950 463.050 679.050 ;
        RECT 469.950 676.950 472.050 679.050 ;
        RECT 448.950 673.950 451.050 676.050 ;
        RECT 454.950 673.950 457.050 676.050 ;
        RECT 442.950 646.950 445.050 649.050 ;
        RECT 439.950 631.950 442.050 634.050 ;
        RECT 443.400 631.050 444.600 646.950 ;
        RECT 451.950 634.950 454.050 637.050 ;
        RECT 442.950 628.950 445.050 631.050 ;
        RECT 448.950 628.950 451.050 631.050 ;
        RECT 430.950 622.950 433.050 625.050 ;
        RECT 397.950 607.950 400.050 610.050 ;
        RECT 418.950 607.950 421.050 610.050 ;
        RECT 418.950 600.600 423.000 601.050 ;
        RECT 418.950 598.950 423.600 600.600 ;
        RECT 409.950 595.950 412.050 598.050 ;
        RECT 397.800 592.950 399.900 595.050 ;
        RECT 401.100 594.600 405.000 595.050 ;
        RECT 401.100 592.950 405.600 594.600 ;
        RECT 398.400 568.050 399.600 592.950 ;
        RECT 404.400 586.050 405.600 592.950 ;
        RECT 403.950 585.600 406.050 586.050 ;
        RECT 403.950 584.400 408.600 585.600 ;
        RECT 403.950 583.950 406.050 584.400 ;
        RECT 397.950 565.950 400.050 568.050 ;
        RECT 407.400 562.200 408.600 584.400 ;
        RECT 410.400 574.050 411.600 595.950 ;
        RECT 422.400 595.050 423.600 598.950 ;
        RECT 430.950 595.950 433.050 598.050 ;
        RECT 443.400 597.600 444.600 628.950 ;
        RECT 445.950 610.950 448.050 613.050 ;
        RECT 446.400 601.050 447.600 610.950 ;
        RECT 449.400 604.050 450.600 628.950 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 445.950 598.950 448.050 601.050 ;
        RECT 443.400 596.400 447.600 597.600 ;
        RECT 421.950 592.950 424.050 595.050 ;
        RECT 431.400 586.050 432.600 595.950 ;
        RECT 430.950 583.950 433.050 586.050 ;
        RECT 439.950 574.950 442.050 577.050 ;
        RECT 409.950 571.950 412.050 574.050 ;
        RECT 427.950 565.950 430.050 568.050 ;
        RECT 376.950 559.950 379.050 562.050 ;
        RECT 391.950 559.950 394.050 562.050 ;
        RECT 406.950 560.100 409.050 562.200 ;
        RECT 388.950 550.950 391.050 553.050 ;
        RECT 382.950 538.950 385.050 541.050 ;
        RECT 373.950 532.950 376.050 535.050 ;
        RECT 373.950 517.950 376.050 520.050 ;
        RECT 374.400 469.050 375.600 517.950 ;
        RECT 376.950 505.950 379.050 508.050 ;
        RECT 377.400 472.200 378.600 505.950 ;
        RECT 383.400 487.050 384.600 538.950 ;
        RECT 389.400 520.050 390.600 550.950 ;
        RECT 392.400 547.050 393.600 559.950 ;
        RECT 428.400 559.050 429.600 565.950 ;
        RECT 433.950 561.600 438.000 562.050 ;
        RECT 433.950 559.950 438.600 561.600 ;
        RECT 406.950 556.800 409.050 558.900 ;
        RECT 421.800 556.950 423.900 559.050 ;
        RECT 427.950 556.950 430.050 559.050 ;
        RECT 397.950 553.950 400.050 556.050 ;
        RECT 391.950 544.950 394.050 547.050 ;
        RECT 398.400 532.050 399.600 553.950 ;
        RECT 407.400 553.050 408.600 556.800 ;
        RECT 412.950 555.600 417.000 556.050 ;
        RECT 412.950 553.950 417.600 555.600 ;
        RECT 406.950 550.950 409.050 553.050 ;
        RECT 409.950 547.950 412.050 550.050 ;
        RECT 397.950 529.950 400.050 532.050 ;
        RECT 410.400 529.050 411.600 547.950 ;
        RECT 416.400 538.050 417.600 553.950 ;
        RECT 422.400 550.050 423.600 556.950 ;
        RECT 437.400 553.050 438.600 559.950 ;
        RECT 436.950 550.950 439.050 553.050 ;
        RECT 421.950 547.950 424.050 550.050 ;
        RECT 440.400 549.600 441.600 574.950 ;
        RECT 442.950 562.950 445.050 565.050 ;
        RECT 443.400 559.050 444.600 562.950 ;
        RECT 442.950 556.950 445.050 559.050 ;
        RECT 440.400 548.400 444.600 549.600 ;
        RECT 439.950 544.950 442.050 547.050 ;
        RECT 415.950 535.950 418.050 538.050 ;
        RECT 427.950 535.950 430.050 538.050 ;
        RECT 436.950 535.950 439.050 538.050 ;
        RECT 391.950 526.950 394.050 529.050 ;
        RECT 407.100 527.400 411.600 529.050 ;
        RECT 407.100 526.950 411.000 527.400 ;
        RECT 388.950 517.950 391.050 520.050 ;
        RECT 383.400 485.400 388.050 487.050 ;
        RECT 384.000 484.950 388.050 485.400 ;
        RECT 376.950 470.100 379.050 472.200 ;
        RECT 386.400 472.050 387.600 484.950 ;
        RECT 385.950 469.950 388.050 472.050 ;
        RECT 374.400 468.900 378.000 469.050 ;
        RECT 374.400 466.950 379.050 468.900 ;
        RECT 370.950 463.950 373.050 466.050 ;
        RECT 364.950 460.950 367.050 463.050 ;
        RECT 370.950 451.950 373.050 454.050 ;
        RECT 371.400 427.050 372.600 451.950 ;
        RECT 374.400 448.050 375.600 466.950 ;
        RECT 376.950 466.800 379.050 466.950 ;
        RECT 388.950 460.950 391.050 463.050 ;
        RECT 389.400 454.050 390.600 460.950 ;
        RECT 379.950 451.950 382.050 454.050 ;
        RECT 385.950 452.400 390.600 454.050 ;
        RECT 385.950 451.950 390.000 452.400 ;
        RECT 373.950 445.950 376.050 448.050 ;
        RECT 370.950 424.950 373.050 427.050 ;
        RECT 376.950 424.950 379.050 427.050 ;
        RECT 370.950 418.950 373.050 421.050 ;
        RECT 365.100 417.600 369.000 418.050 ;
        RECT 365.100 415.950 369.600 417.600 ;
        RECT 368.400 394.050 369.600 415.950 ;
        RECT 367.950 391.950 370.050 394.050 ;
        RECT 364.950 388.950 367.050 391.050 ;
        RECT 352.950 382.950 355.050 385.050 ;
        RECT 361.950 382.950 364.050 385.050 ;
        RECT 353.400 352.200 354.600 382.950 ;
        RECT 352.950 350.100 355.050 352.200 ;
        RECT 365.400 349.050 366.600 388.950 ;
        RECT 367.950 379.950 370.050 382.050 ;
        RECT 368.400 373.050 369.600 379.950 ;
        RECT 367.950 370.950 370.050 373.050 ;
        RECT 371.400 367.050 372.600 418.950 ;
        RECT 373.950 394.950 376.050 397.050 ;
        RECT 370.950 364.950 373.050 367.050 ;
        RECT 374.400 364.050 375.600 394.950 ;
        RECT 377.400 388.050 378.600 424.950 ;
        RECT 380.400 412.050 381.600 451.950 ;
        RECT 392.400 450.600 393.600 526.950 ;
        RECT 400.950 523.950 403.050 526.050 ;
        RECT 401.400 487.050 402.600 523.950 ;
        RECT 407.400 508.050 408.600 526.950 ;
        RECT 421.950 523.950 424.050 526.050 ;
        RECT 428.400 525.600 429.600 535.950 ;
        RECT 437.400 529.050 438.600 535.950 ;
        RECT 440.400 532.200 441.600 544.950 ;
        RECT 439.950 530.100 442.050 532.200 ;
        RECT 436.800 526.950 438.900 529.050 ;
        RECT 440.100 526.800 442.200 528.900 ;
        RECT 433.950 525.600 436.050 526.050 ;
        RECT 428.400 524.400 436.050 525.600 ;
        RECT 433.950 523.950 436.050 524.400 ;
        RECT 406.950 505.950 409.050 508.050 ;
        RECT 406.950 499.950 409.050 502.050 ;
        RECT 407.400 490.050 408.600 499.950 ;
        RECT 422.400 499.050 423.600 523.950 ;
        RECT 424.950 514.950 427.050 517.050 ;
        RECT 421.950 496.950 424.050 499.050 ;
        RECT 425.400 496.050 426.600 514.950 ;
        RECT 440.400 502.050 441.600 526.800 ;
        RECT 439.950 499.950 442.050 502.050 ;
        RECT 409.950 493.950 412.050 496.050 ;
        RECT 424.950 493.950 427.050 496.050 ;
        RECT 406.950 487.950 409.050 490.050 ;
        RECT 397.950 485.400 402.600 487.050 ;
        RECT 397.950 484.950 402.000 485.400 ;
        RECT 398.400 481.050 399.600 484.950 ;
        RECT 410.400 481.050 411.600 493.950 ;
        RECT 418.950 490.950 421.050 493.050 ;
        RECT 419.400 484.050 420.600 490.950 ;
        RECT 418.950 481.950 421.050 484.050 ;
        RECT 397.950 478.950 400.050 481.050 ;
        RECT 409.950 478.950 412.050 481.050 ;
        RECT 415.950 478.950 418.050 481.050 ;
        RECT 433.950 478.950 436.050 481.050 ;
        RECT 410.400 466.050 411.600 478.950 ;
        RECT 397.950 463.950 400.050 466.050 ;
        RECT 409.950 463.950 412.050 466.050 ;
        RECT 395.100 454.950 397.200 457.050 ;
        RECT 395.400 451.050 396.600 454.950 ;
        RECT 398.400 454.050 399.600 463.950 ;
        RECT 416.400 463.050 417.600 478.950 ;
        RECT 418.950 475.950 421.050 478.050 ;
        RECT 415.950 460.950 418.050 463.050 ;
        RECT 403.950 457.950 406.050 460.050 ;
        RECT 412.950 457.950 415.050 460.050 ;
        RECT 404.400 454.050 405.600 457.950 ;
        RECT 397.950 451.950 400.050 454.050 ;
        RECT 403.950 451.950 406.050 454.050 ;
        RECT 394.950 450.600 397.050 451.050 ;
        RECT 392.400 449.400 397.050 450.600 ;
        RECT 394.950 448.950 397.050 449.400 ;
        RECT 382.950 442.950 385.050 445.050 ;
        RECT 379.950 409.950 382.050 412.050 ;
        RECT 383.400 391.050 384.600 442.950 ;
        RECT 398.400 442.050 399.600 451.950 ;
        RECT 397.950 439.950 400.050 442.050 ;
        RECT 391.950 433.950 394.050 436.050 ;
        RECT 385.950 421.950 388.050 424.050 ;
        RECT 386.400 412.050 387.600 421.950 ;
        RECT 388.950 415.950 391.050 418.050 ;
        RECT 386.100 409.950 388.200 412.050 ;
        RECT 385.950 397.950 388.050 400.050 ;
        RECT 382.950 388.950 385.050 391.050 ;
        RECT 386.400 388.050 387.600 397.950 ;
        RECT 376.950 385.950 379.050 388.050 ;
        RECT 385.950 384.000 388.050 388.050 ;
        RECT 386.400 383.400 387.600 384.000 ;
        RECT 389.400 382.050 390.600 415.950 ;
        RECT 388.950 379.950 391.050 382.050 ;
        RECT 373.950 361.950 376.050 364.050 ;
        RECT 392.400 363.600 393.600 433.950 ;
        RECT 406.950 430.950 409.050 433.050 ;
        RECT 400.950 424.950 403.050 427.050 ;
        RECT 401.400 379.050 402.600 424.950 ;
        RECT 400.950 376.950 403.050 379.050 ;
        RECT 389.400 362.400 393.600 363.600 ;
        RECT 389.400 355.050 390.600 362.400 ;
        RECT 376.950 352.950 379.050 355.050 ;
        RECT 388.950 352.950 391.050 355.050 ;
        RECT 377.400 349.050 378.600 352.950 ;
        RECT 352.950 346.800 355.050 348.900 ;
        RECT 364.950 346.950 367.050 349.050 ;
        RECT 376.950 346.950 379.050 349.050 ;
        RECT 343.800 337.950 345.900 340.050 ;
        RECT 349.950 337.950 352.050 340.050 ;
        RECT 337.950 316.950 340.050 319.050 ;
        RECT 331.950 305.400 336.600 307.050 ;
        RECT 331.950 304.950 336.000 305.400 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 335.400 271.050 336.600 289.950 ;
        RECT 337.950 283.950 340.050 286.050 ;
        RECT 343.950 283.950 346.050 286.050 ;
        RECT 328.950 268.950 331.050 271.050 ;
        RECT 334.950 268.950 337.050 271.050 ;
        RECT 323.400 266.400 328.050 268.050 ;
        RECT 324.000 265.950 328.050 266.400 ;
        RECT 319.950 241.950 322.050 244.050 ;
        RECT 328.950 241.950 331.050 244.050 ;
        RECT 319.950 235.950 322.050 238.050 ;
        RECT 316.950 202.950 319.050 205.050 ;
        RECT 310.950 199.950 313.050 202.050 ;
        RECT 302.100 196.950 304.200 199.050 ;
        RECT 289.950 187.950 292.050 190.050 ;
        RECT 277.950 175.950 280.050 178.050 ;
        RECT 271.950 173.400 276.600 175.050 ;
        RECT 271.950 172.950 276.000 173.400 ;
        RECT 268.950 169.950 271.050 172.050 ;
        RECT 277.950 169.950 280.050 172.050 ;
        RECT 256.950 167.400 261.600 169.050 ;
        RECT 256.950 166.950 261.000 167.400 ;
        RECT 269.400 163.050 270.600 169.950 ;
        RECT 268.950 160.950 271.050 163.050 ;
        RECT 274.950 148.950 277.050 151.050 ;
        RECT 275.400 139.050 276.600 148.950 ;
        RECT 274.950 136.950 277.050 139.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 253.950 130.950 256.050 133.050 ;
        RECT 244.950 127.950 247.050 130.050 ;
        RECT 245.400 124.050 246.600 127.950 ;
        RECT 254.400 124.050 255.600 130.950 ;
        RECT 265.950 127.950 268.050 130.050 ;
        RECT 266.400 124.050 267.600 127.950 ;
        RECT 235.950 121.950 238.050 124.050 ;
        RECT 244.950 121.950 247.050 124.050 ;
        RECT 253.950 121.950 256.050 124.050 ;
        RECT 262.950 122.400 267.600 124.050 ;
        RECT 262.950 121.950 267.000 122.400 ;
        RECT 272.400 121.050 273.600 133.950 ;
        RECT 226.950 118.950 229.050 121.050 ;
        RECT 271.950 118.950 274.050 121.050 ;
        RECT 238.950 115.950 241.050 118.050 ;
        RECT 268.950 115.950 271.050 118.050 ;
        RECT 223.950 112.950 226.050 115.050 ;
        RECT 217.950 103.950 220.050 106.050 ;
        RECT 202.950 97.950 205.050 100.050 ;
        RECT 194.400 93.000 198.600 93.600 ;
        RECT 193.950 92.400 198.600 93.000 ;
        RECT 193.950 88.950 196.050 92.400 ;
        RECT 218.400 90.600 219.600 103.950 ;
        RECT 224.400 97.050 225.600 112.950 ;
        RECT 232.950 109.950 235.050 112.050 ;
        RECT 229.950 97.950 232.050 100.050 ;
        RECT 223.950 94.950 226.050 97.050 ;
        RECT 230.400 94.050 231.600 97.950 ;
        RECT 233.400 97.050 234.600 109.950 ;
        RECT 239.400 103.050 240.600 115.950 ;
        RECT 244.950 103.950 247.050 106.050 ;
        RECT 262.950 103.950 265.050 106.050 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 239.400 97.050 240.600 100.950 ;
        RECT 232.950 94.950 235.050 97.050 ;
        RECT 238.800 94.950 240.900 97.050 ;
        RECT 245.400 94.050 246.600 103.950 ;
        RECT 263.400 97.050 264.600 103.950 ;
        RECT 262.800 94.950 264.900 97.050 ;
        RECT 269.400 94.050 270.600 115.950 ;
        RECT 275.400 103.050 276.600 136.950 ;
        RECT 274.950 100.950 277.050 103.050 ;
        RECT 275.400 97.050 276.600 100.950 ;
        RECT 274.950 94.950 277.050 97.050 ;
        RECT 229.950 91.950 232.050 94.050 ;
        RECT 245.400 92.400 250.050 94.050 ;
        RECT 246.000 91.950 250.050 92.400 ;
        RECT 268.950 91.950 271.050 94.050 ;
        RECT 223.950 90.600 226.050 91.050 ;
        RECT 218.400 89.400 226.050 90.600 ;
        RECT 223.950 88.950 226.050 89.400 ;
        RECT 247.950 82.950 250.050 85.050 ;
        RECT 220.950 79.950 223.050 82.050 ;
        RECT 193.950 73.950 196.050 76.050 ;
        RECT 187.950 67.950 190.050 70.050 ;
        RECT 187.950 58.950 190.050 61.050 ;
        RECT 188.400 55.050 189.600 58.950 ;
        RECT 194.400 58.050 195.600 73.950 ;
        RECT 221.400 61.050 222.600 79.950 ;
        RECT 226.950 67.950 229.050 70.050 ;
        RECT 220.950 58.950 223.050 61.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 201.000 57.600 205.050 58.050 ;
        RECT 200.400 55.950 205.050 57.600 ;
        RECT 150.000 54.600 154.050 55.050 ;
        RECT 149.400 52.950 154.050 54.600 ;
        RECT 178.950 52.950 181.050 55.050 ;
        RECT 188.400 53.400 193.050 55.050 ;
        RECT 189.000 52.950 193.050 53.400 ;
        RECT 149.400 49.050 150.600 52.950 ;
        RECT 181.950 49.950 184.050 52.050 ;
        RECT 148.950 46.950 151.050 49.050 ;
        RECT 127.950 34.950 130.050 37.050 ;
        RECT 136.950 34.950 139.050 37.050 ;
        RECT 128.400 22.050 129.600 34.950 ;
        RECT 182.400 34.050 183.600 49.950 ;
        RECT 200.400 43.050 201.600 55.950 ;
        RECT 221.400 52.050 222.600 58.950 ;
        RECT 227.400 55.050 228.600 67.950 ;
        RECT 244.950 58.950 247.050 61.050 ;
        RECT 227.400 53.400 231.900 55.050 ;
        RECT 228.000 52.950 231.900 53.400 ;
        RECT 211.950 46.950 214.050 52.050 ;
        RECT 220.950 49.950 223.050 52.050 ;
        RECT 199.950 40.950 202.050 43.050 ;
        RECT 172.950 31.950 175.050 34.050 ;
        RECT 181.950 31.950 184.050 34.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 124.950 19.950 129.600 22.050 ;
        RECT 118.950 16.950 121.050 19.050 ;
        RECT 112.950 10.950 115.050 13.050 ;
        RECT 82.950 7.950 85.050 10.050 ;
        RECT 128.400 7.050 129.600 19.950 ;
        RECT 131.400 19.050 132.600 22.950 ;
        RECT 173.400 22.200 174.600 31.950 ;
        RECT 200.400 28.050 201.600 40.950 ;
        RECT 214.950 31.950 217.050 34.050 ;
        RECT 211.950 28.950 214.050 31.050 ;
        RECT 181.950 24.600 184.050 28.050 ;
        RECT 199.950 25.950 202.050 28.050 ;
        RECT 181.950 24.000 186.600 24.600 ;
        RECT 182.400 23.400 186.600 24.000 ;
        RECT 136.950 19.950 139.050 22.050 ;
        RECT 166.950 19.950 169.050 22.050 ;
        RECT 172.800 20.100 174.900 22.200 ;
        RECT 181.950 19.950 184.050 22.050 ;
        RECT 131.400 17.400 136.050 19.050 ;
        RECT 132.000 16.950 136.050 17.400 ;
        RECT 137.400 10.050 138.600 19.950 ;
        RECT 167.400 16.050 168.600 19.950 ;
        RECT 174.000 18.600 178.050 19.050 ;
        RECT 173.400 16.950 178.050 18.600 ;
        RECT 166.950 13.950 169.050 16.050 ;
        RECT 173.400 10.050 174.600 16.950 ;
        RECT 182.400 16.050 183.600 19.950 ;
        RECT 185.400 18.600 186.600 23.400 ;
        RECT 205.950 22.950 208.050 25.050 ;
        RECT 196.950 19.950 199.050 22.050 ;
        RECT 193.950 18.600 196.050 19.050 ;
        RECT 185.400 17.400 196.050 18.600 ;
        RECT 193.950 16.950 196.050 17.400 ;
        RECT 197.400 16.050 198.600 19.950 ;
        RECT 181.950 13.950 184.050 16.050 ;
        RECT 196.950 13.950 199.050 16.050 ;
        RECT 197.400 10.050 198.600 13.950 ;
        RECT 206.400 10.050 207.600 22.950 ;
        RECT 212.400 19.050 213.600 28.950 ;
        RECT 215.400 22.050 216.600 31.950 ;
        RECT 217.950 28.950 223.050 31.050 ;
        RECT 245.400 28.050 246.600 58.950 ;
        RECT 248.400 55.050 249.600 82.950 ;
        RECT 274.950 73.950 277.050 76.050 ;
        RECT 271.950 57.600 274.050 58.050 ;
        RECT 266.400 56.400 274.050 57.600 ;
        RECT 248.400 53.400 253.050 55.050 ;
        RECT 249.000 52.950 253.050 53.400 ;
        RECT 253.950 46.950 256.050 49.050 ;
        RECT 254.400 40.050 255.600 46.950 ;
        RECT 253.950 37.950 256.050 40.050 ;
        RECT 247.950 31.950 250.050 34.050 ;
        RECT 235.950 24.600 240.000 25.050 ;
        RECT 235.950 22.950 240.600 24.600 ;
        RECT 244.950 24.000 247.050 28.050 ;
        RECT 245.400 23.400 246.600 24.000 ;
        RECT 215.400 20.400 220.050 22.050 ;
        RECT 216.000 19.950 220.050 20.400 ;
        RECT 211.950 16.950 214.050 19.050 ;
        RECT 239.400 10.050 240.600 22.950 ;
        RECT 248.400 22.050 249.600 31.950 ;
        RECT 266.400 22.050 267.600 56.400 ;
        RECT 271.950 55.950 274.050 56.400 ;
        RECT 275.400 55.050 276.600 73.950 ;
        RECT 278.400 58.050 279.600 169.950 ;
        RECT 290.400 169.050 291.600 187.950 ;
        RECT 295.950 181.950 298.050 184.050 ;
        RECT 296.400 169.050 297.600 181.950 ;
        RECT 289.950 166.950 292.050 169.050 ;
        RECT 295.950 166.950 298.050 169.050 ;
        RECT 298.950 136.950 301.050 139.050 ;
        RECT 280.950 130.950 283.050 133.050 ;
        RECT 281.400 124.050 282.600 130.950 ;
        RECT 299.400 130.050 300.600 136.950 ;
        RECT 302.400 133.050 303.600 196.950 ;
        RECT 310.950 190.950 313.050 193.050 ;
        RECT 304.950 163.950 307.050 166.050 ;
        RECT 305.400 160.050 306.600 163.950 ;
        RECT 304.950 157.950 307.050 160.050 ;
        RECT 307.950 133.950 310.050 136.050 ;
        RECT 301.950 130.950 304.050 133.050 ;
        RECT 286.950 127.950 289.050 130.050 ;
        RECT 298.950 127.950 301.050 130.050 ;
        RECT 287.400 124.050 288.600 127.950 ;
        RECT 308.400 127.050 309.600 133.950 ;
        RECT 292.950 124.950 295.050 127.050 ;
        RECT 304.950 124.950 309.600 127.050 ;
        RECT 280.800 121.950 282.900 124.050 ;
        RECT 286.950 121.950 289.050 124.050 ;
        RECT 293.400 118.050 294.600 124.950 ;
        RECT 292.950 115.950 295.050 118.050 ;
        RECT 295.950 112.950 298.050 115.050 ;
        RECT 304.950 112.950 307.050 115.050 ;
        RECT 289.950 109.950 292.050 112.050 ;
        RECT 290.400 97.050 291.600 109.950 ;
        RECT 296.400 97.050 297.600 112.950 ;
        RECT 289.950 94.950 292.050 97.050 ;
        RECT 295.950 94.950 298.050 97.050 ;
        RECT 305.400 67.050 306.600 112.950 ;
        RECT 308.400 112.050 309.600 124.950 ;
        RECT 311.400 124.050 312.600 190.950 ;
        RECT 320.400 169.050 321.600 235.950 ;
        RECT 325.950 190.950 328.050 193.050 ;
        RECT 319.950 166.950 322.050 169.050 ;
        RECT 326.400 163.050 327.600 190.950 ;
        RECT 325.950 160.950 328.050 163.050 ;
        RECT 311.400 122.400 316.050 124.050 ;
        RECT 312.000 121.950 316.050 122.400 ;
        RECT 319.950 118.950 322.050 121.050 ;
        RECT 307.950 109.950 310.050 112.050 ;
        RECT 320.400 91.050 321.600 118.950 ;
        RECT 322.950 103.950 325.050 106.050 ;
        RECT 323.400 100.050 324.600 103.950 ;
        RECT 322.950 97.950 325.050 100.050 ;
        RECT 323.400 94.050 324.600 97.950 ;
        RECT 323.400 92.400 328.050 94.050 ;
        RECT 324.000 91.950 328.050 92.400 ;
        RECT 316.950 89.400 321.600 91.050 ;
        RECT 316.950 88.950 321.000 89.400 ;
        RECT 325.950 85.950 328.050 88.050 ;
        RECT 326.400 73.050 327.600 85.950 ;
        RECT 325.950 70.950 328.050 73.050 ;
        RECT 329.400 67.050 330.600 241.950 ;
        RECT 338.400 241.050 339.600 283.950 ;
        RECT 344.400 271.050 345.600 283.950 ;
        RECT 350.400 277.050 351.600 337.950 ;
        RECT 353.400 286.050 354.600 346.800 ;
        RECT 373.950 343.950 376.050 346.050 ;
        RECT 385.950 343.950 388.050 346.050 ;
        RECT 397.950 343.950 400.050 346.050 ;
        RECT 355.950 340.950 358.050 343.050 ;
        RECT 356.400 328.050 357.600 340.950 ;
        RECT 355.950 325.950 358.050 328.050 ;
        RECT 370.950 325.950 373.050 328.050 ;
        RECT 364.950 316.950 367.050 319.050 ;
        RECT 365.400 310.050 366.600 316.950 ;
        RECT 371.400 313.050 372.600 325.950 ;
        RECT 367.950 310.950 372.600 313.050 ;
        RECT 364.950 307.950 367.050 310.050 ;
        RECT 371.400 298.050 372.600 310.950 ;
        RECT 370.950 295.950 373.050 298.050 ;
        RECT 374.400 295.050 375.600 343.950 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 377.400 328.050 378.600 334.950 ;
        RECT 382.950 328.950 385.050 331.050 ;
        RECT 376.950 325.950 379.050 328.050 ;
        RECT 376.950 316.950 379.050 319.050 ;
        RECT 377.400 313.050 378.600 316.950 ;
        RECT 377.400 311.400 382.050 313.050 ;
        RECT 378.000 310.950 382.050 311.400 ;
        RECT 376.950 295.950 379.050 298.050 ;
        RECT 373.950 292.950 376.050 295.050 ;
        RECT 352.950 283.950 355.050 286.050 ;
        RECT 361.950 277.950 364.050 280.050 ;
        RECT 349.950 274.950 352.050 277.050 ;
        RECT 362.400 271.050 363.600 277.950 ;
        RECT 370.950 271.950 373.050 274.050 ;
        RECT 343.950 268.950 346.050 271.050 ;
        RECT 361.950 268.950 364.050 271.050 ;
        RECT 371.400 268.050 372.600 271.950 ;
        RECT 377.400 271.050 378.600 295.950 ;
        RECT 376.950 268.950 379.050 271.050 ;
        RECT 352.800 267.600 354.900 268.050 ;
        RECT 359.100 267.600 361.200 268.050 ;
        RECT 352.800 266.400 361.200 267.600 ;
        RECT 352.800 265.950 354.900 266.400 ;
        RECT 359.100 265.950 361.200 266.400 ;
        RECT 370.950 265.950 373.050 268.050 ;
        RECT 355.950 262.950 358.050 265.050 ;
        RECT 343.950 244.950 346.050 247.050 ;
        RECT 337.950 238.950 340.050 241.050 ;
        RECT 344.400 238.050 345.600 244.950 ;
        RECT 331.950 235.950 334.050 238.050 ;
        RECT 343.950 235.950 346.050 238.050 ;
        RECT 332.400 223.050 333.600 235.950 ;
        RECT 346.950 223.950 349.050 226.050 ;
        RECT 331.950 220.950 334.050 223.050 ;
        RECT 331.950 202.950 334.050 205.050 ;
        RECT 332.400 154.050 333.600 202.950 ;
        RECT 339.000 201.600 343.050 202.050 ;
        RECT 338.400 199.950 343.050 201.600 ;
        RECT 334.950 187.950 337.050 193.050 ;
        RECT 338.400 187.050 339.600 199.950 ;
        RECT 347.400 196.050 348.600 223.950 ;
        RECT 349.800 214.950 351.900 217.050 ;
        RECT 353.100 214.950 355.200 217.050 ;
        RECT 350.400 211.050 351.600 214.950 ;
        RECT 349.950 208.950 352.050 211.050 ;
        RECT 353.400 202.200 354.600 214.950 ;
        RECT 352.950 200.100 355.050 202.200 ;
        RECT 352.950 196.800 355.050 198.900 ;
        RECT 346.950 193.950 349.050 196.050 ;
        RECT 337.950 184.950 340.050 187.050 ;
        RECT 343.950 184.950 346.050 187.050 ;
        RECT 338.400 169.050 339.600 184.950 ;
        RECT 344.400 178.050 345.600 184.950 ;
        RECT 353.400 184.050 354.600 196.800 ;
        RECT 356.400 187.050 357.600 262.950 ;
        RECT 364.950 253.950 367.050 256.050 ;
        RECT 358.950 235.950 361.050 238.050 ;
        RECT 359.400 214.050 360.600 235.950 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 365.400 211.050 366.600 253.950 ;
        RECT 367.950 247.950 370.050 250.050 ;
        RECT 364.950 208.950 367.050 211.050 ;
        RECT 358.950 205.950 361.050 208.050 ;
        RECT 359.400 199.050 360.600 205.950 ;
        RECT 365.400 202.050 366.600 208.950 ;
        RECT 368.400 205.050 369.600 247.950 ;
        RECT 370.950 238.950 373.050 241.050 ;
        RECT 371.400 214.050 372.600 238.950 ;
        RECT 383.400 220.050 384.600 328.950 ;
        RECT 386.400 313.200 387.600 343.950 ;
        RECT 388.950 340.950 391.050 343.050 ;
        RECT 385.950 311.100 388.050 313.200 ;
        RECT 389.400 310.050 390.600 340.950 ;
        RECT 398.400 310.050 399.600 343.950 ;
        RECT 407.400 343.050 408.600 430.950 ;
        RECT 413.400 415.050 414.600 457.950 ;
        RECT 412.950 412.950 415.050 415.050 ;
        RECT 415.950 409.950 418.050 412.050 ;
        RECT 409.950 406.950 412.050 409.050 ;
        RECT 410.400 403.050 411.600 406.950 ;
        RECT 416.400 406.050 417.600 409.950 ;
        RECT 415.950 403.950 418.050 406.050 ;
        RECT 409.950 400.950 412.050 403.050 ;
        RECT 419.400 394.050 420.600 475.950 ;
        RECT 427.950 472.950 430.050 475.050 ;
        RECT 428.400 457.050 429.600 472.950 ;
        RECT 434.400 472.050 435.600 478.950 ;
        RECT 443.400 474.600 444.600 548.400 ;
        RECT 446.400 505.050 447.600 596.400 ;
        RECT 452.400 595.050 453.600 634.950 ;
        RECT 451.950 592.950 454.050 595.050 ;
        RECT 455.400 580.050 456.600 673.950 ;
        RECT 457.950 670.950 460.050 673.050 ;
        RECT 463.950 670.950 466.050 673.050 ;
        RECT 458.400 652.050 459.600 670.950 ;
        RECT 464.400 658.050 465.600 670.950 ;
        RECT 463.950 655.950 466.050 658.050 ;
        RECT 457.950 649.950 460.050 652.050 ;
        RECT 458.400 646.050 459.600 649.950 ;
        RECT 457.950 643.950 460.050 646.050 ;
        RECT 470.400 634.050 471.600 676.950 ;
        RECT 476.400 672.600 477.600 703.950 ;
        RECT 481.950 694.950 484.050 697.050 ;
        RECT 482.400 673.050 483.600 694.950 ;
        RECT 488.400 673.050 489.600 706.950 ;
        RECT 497.100 703.950 499.200 706.050 ;
        RECT 497.400 685.050 498.600 703.950 ;
        RECT 496.950 682.950 499.050 685.050 ;
        RECT 503.400 679.050 504.600 739.950 ;
        RECT 509.400 738.600 510.600 742.950 ;
        RECT 506.400 737.400 510.600 738.600 ;
        RECT 506.400 709.050 507.600 737.400 ;
        RECT 508.950 718.950 511.050 721.050 ;
        RECT 505.950 706.950 508.050 709.050 ;
        RECT 506.400 688.050 507.600 706.950 ;
        RECT 505.950 685.950 508.050 688.050 ;
        RECT 502.950 676.950 505.050 679.050 ;
        RECT 499.950 673.950 502.050 676.050 ;
        RECT 473.400 672.000 477.600 672.600 ;
        RECT 472.950 671.400 477.600 672.000 ;
        RECT 472.950 670.050 475.050 671.400 ;
        RECT 481.800 670.950 483.900 673.050 ;
        RECT 487.950 670.950 490.050 673.050 ;
        RECT 500.400 670.050 501.600 673.950 ;
        RECT 506.400 673.050 507.600 685.950 ;
        RECT 505.950 670.950 508.050 673.050 ;
        RECT 472.800 669.000 475.050 670.050 ;
        RECT 472.800 667.950 474.900 669.000 ;
        RECT 478.950 667.950 481.050 670.050 ;
        RECT 484.950 667.950 487.050 670.050 ;
        RECT 499.950 667.950 502.050 670.050 ;
        RECT 472.950 637.950 475.050 640.050 ;
        RECT 469.950 631.950 472.050 634.050 ;
        RECT 473.400 631.050 474.600 637.950 ;
        RECT 479.400 634.050 480.600 667.950 ;
        RECT 485.400 664.050 486.600 667.950 ;
        RECT 484.950 661.950 487.050 664.050 ;
        RECT 478.950 631.950 481.050 634.050 ;
        RECT 473.400 629.400 478.050 631.050 ;
        RECT 474.000 628.950 478.050 629.400 ;
        RECT 457.950 622.950 460.050 625.050 ;
        RECT 458.400 604.050 459.600 622.950 ;
        RECT 479.400 613.050 480.600 631.950 ;
        RECT 485.400 628.050 486.600 661.950 ;
        RECT 490.950 658.950 493.050 661.050 ;
        RECT 491.400 631.050 492.600 658.950 ;
        RECT 499.950 634.950 502.050 637.050 ;
        RECT 487.950 629.400 492.600 631.050 ;
        RECT 487.950 628.950 492.000 629.400 ;
        RECT 494.100 628.950 496.200 631.050 ;
        RECT 484.950 625.950 487.050 628.050 ;
        RECT 494.400 622.050 495.600 628.950 ;
        RECT 500.400 625.050 501.600 634.950 ;
        RECT 505.950 625.950 508.050 628.050 ;
        RECT 499.950 622.950 502.050 625.050 ;
        RECT 493.950 619.950 496.050 622.050 ;
        RECT 484.950 613.950 487.050 616.050 ;
        RECT 478.950 610.950 481.050 613.050 ;
        RECT 457.950 600.000 460.050 604.050 ;
        RECT 458.400 599.400 459.600 600.000 ;
        RECT 463.800 595.950 465.900 598.050 ;
        RECT 481.950 597.600 484.050 601.050 ;
        RECT 485.400 597.600 486.600 613.950 ;
        RECT 500.400 610.050 501.600 622.950 ;
        RECT 506.400 622.050 507.600 625.950 ;
        RECT 505.950 619.950 508.050 622.050 ;
        RECT 499.950 607.950 502.050 610.050 ;
        RECT 490.950 604.950 493.050 607.050 ;
        RECT 481.950 597.000 486.600 597.600 ;
        RECT 482.400 596.400 486.600 597.000 ;
        RECT 460.950 592.950 463.050 595.050 ;
        RECT 457.950 586.950 460.050 589.050 ;
        RECT 458.400 583.050 459.600 586.950 ;
        RECT 457.950 580.950 460.050 583.050 ;
        RECT 454.950 577.950 457.050 580.050 ;
        RECT 461.400 571.050 462.600 592.950 ;
        RECT 460.950 568.950 463.050 571.050 ;
        RECT 464.400 568.050 465.600 595.950 ;
        RECT 475.950 594.600 480.000 595.050 ;
        RECT 475.950 592.950 480.600 594.600 ;
        RECT 488.100 592.950 490.200 595.050 ;
        RECT 479.400 580.050 480.600 592.950 ;
        RECT 478.950 577.950 481.050 580.050 ;
        RECT 488.400 577.050 489.600 592.950 ;
        RECT 466.950 574.950 469.050 577.050 ;
        RECT 487.950 574.950 490.050 577.050 ;
        RECT 467.400 571.050 468.600 574.950 ;
        RECT 469.950 571.950 472.050 574.050 ;
        RECT 466.950 568.950 469.050 571.050 ;
        RECT 451.950 565.950 454.050 568.050 ;
        RECT 457.950 565.950 460.050 568.050 ;
        RECT 463.950 565.950 466.050 568.050 ;
        RECT 452.400 556.050 453.600 565.950 ;
        RECT 458.400 559.050 459.600 565.950 ;
        RECT 470.400 562.050 471.600 571.950 ;
        RECT 487.950 565.950 490.050 568.050 ;
        RECT 469.950 559.950 472.050 562.050 ;
        RECT 457.800 556.950 459.900 559.050 ;
        RECT 448.950 554.400 453.600 556.050 ;
        RECT 448.950 553.950 453.000 554.400 ;
        RECT 458.400 541.050 459.600 556.950 ;
        RECT 470.400 556.050 471.600 559.950 ;
        RECT 461.100 553.950 463.200 556.050 ;
        RECT 469.950 553.950 472.050 556.050 ;
        RECT 479.100 555.600 483.000 556.050 ;
        RECT 479.100 553.950 483.600 555.600 ;
        RECT 461.400 550.050 462.600 553.950 ;
        RECT 463.950 550.950 466.050 553.050 ;
        RECT 460.950 547.950 463.050 550.050 ;
        RECT 457.950 538.950 460.050 541.050 ;
        RECT 454.800 523.950 456.900 526.050 ;
        RECT 445.950 502.950 448.050 505.050 ;
        RECT 455.400 495.600 456.600 523.950 ;
        RECT 464.400 523.050 465.600 550.950 ;
        RECT 466.950 532.950 469.050 535.050 ;
        RECT 467.400 526.050 468.600 532.950 ;
        RECT 470.400 528.600 471.600 553.950 ;
        RECT 482.400 544.050 483.600 553.950 ;
        RECT 481.950 541.950 484.050 544.050 ;
        RECT 478.950 538.950 481.050 541.050 ;
        RECT 479.400 529.050 480.600 538.950 ;
        RECT 488.400 535.050 489.600 565.950 ;
        RECT 491.400 553.050 492.600 604.950 ;
        RECT 506.400 604.050 507.600 619.950 ;
        RECT 505.950 601.950 508.050 604.050 ;
        RECT 505.950 577.950 508.050 580.050 ;
        RECT 502.950 559.950 505.050 565.050 ;
        RECT 490.950 550.950 493.050 553.050 ;
        RECT 487.950 532.950 490.050 535.050 ;
        RECT 491.400 532.050 492.600 550.950 ;
        RECT 502.950 538.950 505.050 541.050 ;
        RECT 484.950 529.050 487.050 532.050 ;
        RECT 490.950 529.950 493.050 532.050 ;
        RECT 503.400 529.050 504.600 538.950 ;
        RECT 470.400 527.400 474.600 528.600 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 463.950 520.950 466.050 523.050 ;
        RECT 473.400 514.050 474.600 527.400 ;
        RECT 478.800 526.950 480.900 529.050 ;
        RECT 484.950 528.000 487.200 529.050 ;
        RECT 485.100 526.950 487.200 528.000 ;
        RECT 502.950 526.950 505.050 529.050 ;
        RECT 472.950 511.950 475.050 514.050 ;
        RECT 484.950 511.950 487.050 514.050 ;
        RECT 460.950 508.950 463.050 511.050 ;
        RECT 455.400 494.400 459.600 495.600 ;
        RECT 448.950 490.950 451.050 493.050 ;
        RECT 453.000 492.600 457.050 493.050 ;
        RECT 452.400 490.950 457.050 492.600 ;
        RECT 449.400 487.050 450.600 490.950 ;
        RECT 448.950 484.950 451.050 487.050 ;
        RECT 443.400 473.400 447.600 474.600 ;
        RECT 433.950 469.950 436.050 472.050 ;
        RECT 442.950 469.950 445.050 472.050 ;
        RECT 436.950 463.950 439.050 466.050 ;
        RECT 433.950 457.950 436.050 460.050 ;
        RECT 424.950 455.400 429.600 457.050 ;
        RECT 424.950 454.950 429.000 455.400 ;
        RECT 424.950 445.950 427.050 448.050 ;
        RECT 421.950 442.950 424.050 445.050 ;
        RECT 418.950 391.950 421.050 394.050 ;
        RECT 409.950 364.950 412.050 367.050 ;
        RECT 410.400 349.050 411.600 364.950 ;
        RECT 409.950 346.950 412.050 349.050 ;
        RECT 406.950 340.950 409.050 343.050 ;
        RECT 412.950 328.950 415.050 331.050 ;
        RECT 402.000 312.600 406.050 313.050 ;
        RECT 388.950 309.600 391.050 310.050 ;
        RECT 386.400 308.400 391.050 309.600 ;
        RECT 382.950 217.950 385.050 220.050 ;
        RECT 370.950 211.950 373.050 214.050 ;
        RECT 367.950 202.950 370.050 205.050 ;
        RECT 365.100 199.950 367.200 202.050 ;
        RECT 359.400 196.950 364.050 199.050 ;
        RECT 370.950 196.950 373.050 199.050 ;
        RECT 377.400 198.000 378.600 198.600 ;
        RECT 359.400 187.050 360.600 196.950 ;
        RECT 355.800 184.950 357.900 187.050 ;
        RECT 359.100 184.950 361.200 187.050 ;
        RECT 352.950 181.950 355.050 184.050 ;
        RECT 349.950 178.950 352.050 181.050 ;
        RECT 343.950 175.950 346.050 178.050 ;
        RECT 343.950 169.950 346.050 172.050 ;
        RECT 334.950 167.400 339.600 169.050 ;
        RECT 334.950 166.950 339.000 167.400 ;
        RECT 344.400 166.050 345.600 169.950 ;
        RECT 350.400 169.050 351.600 178.950 ;
        RECT 352.950 175.950 355.050 178.050 ;
        RECT 349.950 166.950 352.050 169.050 ;
        RECT 343.800 163.950 345.900 166.050 ;
        RECT 334.950 160.950 337.050 163.050 ;
        RECT 331.950 151.950 334.050 154.050 ;
        RECT 331.950 124.950 334.050 127.050 ;
        RECT 332.400 118.050 333.600 124.950 ;
        RECT 331.950 115.950 334.050 118.050 ;
        RECT 332.400 106.050 333.600 115.950 ;
        RECT 331.950 103.950 334.050 106.050 ;
        RECT 335.400 67.050 336.600 160.950 ;
        RECT 346.950 136.950 349.050 139.050 ;
        RECT 340.950 130.950 343.050 133.050 ;
        RECT 341.400 124.050 342.600 130.950 ;
        RECT 347.400 127.050 348.600 136.950 ;
        RECT 346.950 124.950 349.050 127.050 ;
        RECT 340.950 121.950 343.050 124.050 ;
        RECT 353.400 97.050 354.600 175.950 ;
        RECT 361.950 169.950 364.050 172.050 ;
        RECT 362.400 166.050 363.600 169.950 ;
        RECT 371.400 169.050 372.600 196.950 ;
        RECT 376.950 193.950 379.050 198.000 ;
        RECT 373.950 187.950 376.050 190.050 ;
        RECT 370.950 166.950 373.050 169.050 ;
        RECT 374.400 166.050 375.600 187.950 ;
        RECT 377.400 175.050 378.600 193.950 ;
        RECT 382.950 181.950 385.050 184.050 ;
        RECT 376.950 172.950 379.050 175.050 ;
        RECT 383.400 166.050 384.600 181.950 ;
        RECT 358.950 164.400 363.600 166.050 ;
        RECT 358.950 163.950 363.000 164.400 ;
        RECT 373.950 163.950 376.050 166.050 ;
        RECT 383.100 163.950 385.200 166.050 ;
        RECT 364.950 148.950 367.050 151.050 ;
        RECT 365.400 126.600 366.600 148.950 ;
        RECT 383.400 135.600 384.600 163.950 ;
        RECT 380.400 134.400 384.600 135.600 ;
        RECT 370.950 127.950 373.050 130.050 ;
        RECT 365.400 125.400 369.600 126.600 ;
        RECT 361.950 121.950 364.050 124.050 ;
        RECT 355.950 97.950 358.050 100.050 ;
        RECT 342.000 96.600 346.050 97.050 ;
        RECT 341.400 94.950 346.050 96.600 ;
        RECT 352.950 94.950 355.050 97.050 ;
        RECT 341.400 70.050 342.600 94.950 ;
        RECT 340.950 67.950 343.050 70.050 ;
        RECT 304.950 64.950 307.050 67.050 ;
        RECT 316.950 64.950 319.050 67.050 ;
        RECT 328.950 64.950 331.050 67.050 ;
        RECT 334.950 64.950 337.050 67.050 ;
        RECT 304.950 58.950 307.050 61.050 ;
        RECT 277.950 55.950 280.050 58.050 ;
        RECT 274.950 52.950 277.050 55.050 ;
        RECT 292.950 52.950 295.050 55.050 ;
        RECT 271.950 49.950 274.050 52.050 ;
        RECT 268.950 25.950 271.050 28.050 ;
        RECT 248.400 20.400 253.050 22.050 ;
        RECT 249.000 19.950 253.050 20.400 ;
        RECT 265.950 19.950 268.050 22.050 ;
        RECT 269.400 16.050 270.600 25.950 ;
        RECT 268.950 13.950 271.050 16.050 ;
        RECT 272.400 13.050 273.600 49.950 ;
        RECT 286.950 43.950 289.050 46.050 ;
        RECT 277.950 34.950 280.050 37.050 ;
        RECT 278.400 22.050 279.600 34.950 ;
        RECT 287.400 22.050 288.600 43.950 ;
        RECT 293.400 31.050 294.600 52.950 ;
        RECT 305.400 49.050 306.600 58.950 ;
        RECT 317.400 58.050 318.600 64.950 ;
        RECT 334.950 58.950 337.050 61.050 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 304.950 46.950 307.050 49.050 ;
        RECT 310.950 43.950 313.050 46.050 ;
        RECT 295.950 34.950 298.050 37.050 ;
        RECT 296.400 31.050 297.600 34.950 ;
        RECT 292.800 28.950 294.900 31.050 ;
        RECT 296.100 28.950 298.200 31.050 ;
        RECT 301.950 28.950 304.050 31.050 ;
        RECT 302.400 25.050 303.600 28.950 ;
        RECT 311.400 28.050 312.600 43.950 ;
        RECT 317.100 40.950 319.200 43.050 ;
        RECT 317.400 28.050 318.600 40.950 ;
        RECT 322.950 37.950 325.050 40.050 ;
        RECT 323.400 31.050 324.600 37.950 ;
        RECT 335.400 37.050 336.600 58.950 ;
        RECT 356.400 58.050 357.600 97.950 ;
        RECT 359.400 96.000 360.600 96.600 ;
        RECT 358.950 94.050 361.050 96.000 ;
        RECT 358.800 93.000 361.050 94.050 ;
        RECT 358.800 91.950 360.900 93.000 ;
        RECT 359.400 88.050 360.600 91.950 ;
        RECT 362.400 91.050 363.600 121.950 ;
        RECT 364.950 115.950 367.050 118.050 ;
        RECT 365.400 103.050 366.600 115.950 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 368.400 100.050 369.600 125.400 ;
        RECT 367.950 97.950 370.050 100.050 ;
        RECT 371.400 97.200 372.600 127.950 ;
        RECT 380.400 127.200 381.600 134.400 ;
        RECT 386.400 130.050 387.600 308.400 ;
        RECT 388.950 307.950 391.050 308.400 ;
        RECT 394.950 308.400 399.600 310.050 ;
        RECT 401.400 310.950 406.050 312.600 ;
        RECT 394.950 307.950 399.000 308.400 ;
        RECT 388.950 277.950 391.050 280.050 ;
        RECT 389.400 271.050 390.600 277.950 ;
        RECT 395.400 274.050 396.600 307.950 ;
        RECT 401.400 301.050 402.600 310.950 ;
        RECT 406.950 307.950 409.050 310.050 ;
        RECT 400.950 298.950 403.050 301.050 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 395.400 272.400 400.050 274.050 ;
        RECT 396.000 271.950 400.050 272.400 ;
        RECT 388.950 268.950 391.050 271.050 ;
        RECT 388.950 262.950 391.050 265.050 ;
        RECT 389.400 151.050 390.600 262.950 ;
        RECT 404.400 253.050 405.600 289.950 ;
        RECT 403.950 250.950 406.050 253.050 ;
        RECT 407.400 241.050 408.600 307.950 ;
        RECT 409.950 259.950 412.050 262.050 ;
        RECT 403.950 239.400 408.600 241.050 ;
        RECT 403.950 238.950 408.000 239.400 ;
        RECT 406.950 232.950 409.050 235.050 ;
        RECT 407.400 226.050 408.600 232.950 ;
        RECT 406.950 223.950 409.050 226.050 ;
        RECT 391.950 205.950 394.050 208.050 ;
        RECT 392.400 199.050 393.600 205.950 ;
        RECT 391.950 196.950 394.050 199.050 ;
        RECT 397.950 196.950 400.050 199.050 ;
        RECT 398.400 187.050 399.600 196.950 ;
        RECT 397.950 184.950 400.050 187.050 ;
        RECT 406.950 181.950 409.050 184.050 ;
        RECT 407.400 169.050 408.600 181.950 ;
        RECT 406.950 166.950 409.050 169.050 ;
        RECT 391.950 163.950 394.050 166.050 ;
        RECT 388.950 148.950 391.050 151.050 ;
        RECT 385.950 127.950 388.050 130.050 ;
        RECT 379.950 125.100 382.050 127.200 ;
        RECT 392.400 127.050 393.600 163.950 ;
        RECT 410.400 157.050 411.600 259.950 ;
        RECT 413.400 253.050 414.600 328.950 ;
        RECT 419.400 310.050 420.600 391.950 ;
        RECT 422.400 373.200 423.600 442.950 ;
        RECT 421.950 371.100 424.050 373.200 ;
        RECT 421.950 367.800 424.050 369.900 ;
        RECT 422.400 343.050 423.600 367.800 ;
        RECT 421.950 340.950 424.050 343.050 ;
        RECT 425.400 331.050 426.600 445.950 ;
        RECT 427.950 415.950 430.050 421.050 ;
        RECT 434.400 414.600 435.600 457.950 ;
        RECT 437.400 427.050 438.600 463.950 ;
        RECT 443.400 436.050 444.600 469.950 ;
        RECT 446.400 445.050 447.600 473.400 ;
        RECT 445.950 442.950 448.050 445.050 ;
        RECT 442.950 433.950 445.050 436.050 ;
        RECT 452.400 433.050 453.600 490.950 ;
        RECT 458.400 490.050 459.600 494.400 ;
        RECT 457.950 487.950 460.050 490.050 ;
        RECT 457.950 442.950 460.050 445.050 ;
        RECT 454.950 433.950 457.050 436.050 ;
        RECT 451.950 430.950 454.050 433.050 ;
        RECT 436.950 424.950 439.050 427.050 ;
        RECT 448.950 418.950 451.050 421.050 ;
        RECT 434.400 413.400 438.600 414.600 ;
        RECT 433.950 409.950 436.050 412.050 ;
        RECT 427.950 406.950 430.050 409.050 ;
        RECT 428.400 403.050 429.600 406.950 ;
        RECT 427.950 400.950 430.050 403.050 ;
        RECT 434.400 399.600 435.600 409.950 ;
        RECT 431.400 398.400 435.600 399.600 ;
        RECT 431.400 394.050 432.600 398.400 ;
        RECT 437.400 397.050 438.600 413.400 ;
        RECT 439.950 412.950 442.050 415.050 ;
        RECT 440.400 403.050 441.600 412.950 ;
        RECT 449.400 412.050 450.600 418.950 ;
        RECT 455.400 415.050 456.600 433.950 ;
        RECT 454.950 412.950 457.050 415.050 ;
        RECT 448.950 409.950 451.050 412.050 ;
        RECT 442.950 403.950 445.050 406.050 ;
        RECT 439.950 400.950 442.050 403.050 ;
        RECT 436.950 394.950 439.050 397.050 ;
        RECT 430.950 391.950 433.050 394.050 ;
        RECT 443.400 385.050 444.600 403.950 ;
        RECT 458.400 403.050 459.600 442.950 ;
        RECT 457.950 400.950 460.050 403.050 ;
        RECT 454.950 394.950 457.050 397.050 ;
        RECT 437.400 384.000 438.600 384.600 ;
        RECT 436.950 382.050 439.050 384.000 ;
        RECT 443.400 383.400 448.050 385.050 ;
        RECT 444.000 382.950 448.050 383.400 ;
        RECT 436.800 381.000 439.050 382.050 ;
        RECT 436.800 379.950 438.900 381.000 ;
        RECT 448.950 379.950 451.050 382.050 ;
        RECT 430.950 376.950 433.050 379.050 ;
        RECT 431.400 361.050 432.600 376.950 ;
        RECT 437.400 370.050 438.600 379.950 ;
        RECT 436.950 367.950 439.050 370.050 ;
        RECT 430.950 358.950 433.050 361.050 ;
        RECT 436.950 358.950 439.050 361.050 ;
        RECT 430.950 352.950 433.050 355.050 ;
        RECT 427.950 337.950 430.050 340.050 ;
        RECT 424.950 328.950 427.050 331.050 ;
        RECT 421.950 319.950 424.050 322.050 ;
        RECT 422.400 316.050 423.600 319.950 ;
        RECT 421.950 313.950 424.050 316.050 ;
        RECT 422.400 310.050 423.600 313.950 ;
        RECT 418.800 307.950 420.900 310.050 ;
        RECT 422.100 307.950 424.200 310.050 ;
        RECT 428.400 307.050 429.600 337.950 ;
        RECT 427.950 304.950 430.050 307.050 ;
        RECT 415.950 301.950 418.050 304.050 ;
        RECT 416.400 283.050 417.600 301.950 ;
        RECT 431.400 301.050 432.600 352.950 ;
        RECT 437.400 328.050 438.600 358.950 ;
        RECT 439.950 346.950 442.050 349.050 ;
        RECT 436.950 325.950 439.050 328.050 ;
        RECT 440.400 322.050 441.600 346.950 ;
        RECT 445.950 340.950 448.050 343.050 ;
        RECT 446.400 337.050 447.600 340.950 ;
        RECT 442.950 335.400 447.600 337.050 ;
        RECT 442.950 334.950 447.000 335.400 ;
        RECT 449.400 333.600 450.600 379.950 ;
        RECT 455.400 340.050 456.600 394.950 ;
        RECT 458.400 352.050 459.600 400.950 ;
        RECT 461.400 397.050 462.600 508.950 ;
        RECT 472.950 502.950 475.050 505.050 ;
        RECT 463.950 487.950 466.050 490.050 ;
        RECT 464.400 460.050 465.600 487.950 ;
        RECT 469.950 481.950 472.050 484.050 ;
        RECT 463.800 457.950 465.900 460.050 ;
        RECT 467.100 457.950 469.200 460.050 ;
        RECT 467.400 448.050 468.600 457.950 ;
        RECT 470.400 454.050 471.600 481.950 ;
        RECT 473.400 472.050 474.600 502.950 ;
        RECT 485.400 490.050 486.600 511.950 ;
        RECT 506.400 505.200 507.600 577.950 ;
        RECT 505.950 503.100 508.050 505.200 ;
        RECT 505.950 499.800 508.050 501.900 ;
        RECT 484.950 487.950 487.050 490.050 ;
        RECT 487.950 484.950 490.050 487.050 ;
        RECT 484.950 472.950 487.050 478.050 ;
        RECT 472.950 469.950 475.050 472.050 ;
        RECT 484.950 466.950 487.050 469.050 ;
        RECT 469.800 451.950 471.900 454.050 ;
        RECT 485.400 448.050 486.600 466.950 ;
        RECT 488.400 457.050 489.600 484.950 ;
        RECT 506.400 478.050 507.600 499.800 ;
        RECT 505.950 475.950 508.050 478.050 ;
        RECT 505.950 466.950 508.050 469.050 ;
        RECT 506.400 463.050 507.600 466.950 ;
        RECT 505.950 460.950 508.050 463.050 ;
        RECT 493.950 457.050 496.050 460.050 ;
        RECT 487.800 454.950 489.900 457.050 ;
        RECT 493.950 456.000 496.200 457.050 ;
        RECT 494.100 454.950 496.200 456.000 ;
        RECT 499.950 454.950 502.050 457.050 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 466.950 430.950 469.050 433.050 ;
        RECT 463.950 427.950 466.050 430.050 ;
        RECT 464.400 418.050 465.600 427.950 ;
        RECT 463.950 415.950 466.050 418.050 ;
        RECT 460.950 394.950 463.050 397.050 ;
        RECT 461.400 385.050 462.600 394.950 ;
        RECT 460.950 382.950 463.050 385.050 ;
        RECT 463.950 358.950 466.050 361.050 ;
        RECT 457.950 349.950 460.050 352.050 ;
        RECT 464.400 340.050 465.600 358.950 ;
        RECT 467.400 348.600 468.600 430.950 ;
        RECT 500.400 430.050 501.600 454.950 ;
        RECT 509.400 454.050 510.600 718.950 ;
        RECT 511.950 703.950 514.050 706.050 ;
        RECT 512.400 697.050 513.600 703.950 ;
        RECT 515.400 703.050 516.600 754.950 ;
        RECT 520.950 745.950 523.050 748.050 ;
        RECT 517.950 736.950 520.050 739.050 ;
        RECT 518.400 712.050 519.600 736.950 ;
        RECT 521.400 736.050 522.600 745.950 ;
        RECT 533.400 742.050 534.600 799.950 ;
        RECT 535.950 790.950 538.050 793.050 ;
        RECT 526.950 739.950 529.050 742.050 ;
        RECT 532.950 739.950 535.050 742.050 ;
        RECT 520.950 733.950 523.050 736.050 ;
        RECT 523.950 724.950 526.050 727.050 ;
        RECT 517.950 709.950 520.050 712.050 ;
        RECT 514.950 700.950 517.050 703.050 ;
        RECT 518.400 700.050 519.600 709.950 ;
        RECT 524.400 703.050 525.600 724.950 ;
        RECT 523.950 702.600 526.050 703.050 ;
        RECT 521.400 701.400 526.050 702.600 ;
        RECT 517.950 697.950 520.050 700.050 ;
        RECT 511.950 694.950 514.050 697.050 ;
        RECT 512.400 661.050 513.600 694.950 ;
        RECT 514.950 691.950 517.050 694.050 ;
        RECT 515.400 670.050 516.600 691.950 ;
        RECT 515.400 668.400 520.050 670.050 ;
        RECT 516.000 667.950 520.050 668.400 ;
        RECT 511.950 658.950 514.050 661.050 ;
        RECT 521.400 645.600 522.600 701.400 ;
        RECT 523.950 700.950 526.050 701.400 ;
        RECT 527.400 667.050 528.600 739.950 ;
        RECT 536.400 721.050 537.600 790.950 ;
        RECT 554.400 784.050 555.600 835.950 ;
        RECT 565.950 826.950 568.050 829.050 ;
        RECT 566.400 811.050 567.600 826.950 ;
        RECT 569.400 817.050 570.600 838.950 ;
        RECT 575.400 837.600 576.600 844.950 ;
        RECT 602.400 841.050 603.600 862.950 ;
        RECT 635.400 847.050 636.600 862.950 ;
        RECT 641.400 853.050 642.600 865.950 ;
        RECT 640.800 850.950 642.900 853.050 ;
        RECT 644.100 847.950 646.200 850.050 ;
        RECT 715.950 847.950 718.050 850.050 ;
        RECT 634.950 844.950 637.050 847.050 ;
        RECT 601.950 838.950 604.050 841.050 ;
        RECT 631.950 838.950 634.050 841.050 ;
        RECT 572.400 836.400 576.600 837.600 ;
        RECT 572.400 829.050 573.600 836.400 ;
        RECT 577.950 832.950 580.050 835.050 ;
        RECT 616.950 832.950 619.050 835.050 ;
        RECT 571.950 826.950 574.050 829.050 ;
        RECT 568.800 814.950 570.900 817.050 ;
        RECT 572.100 814.950 574.200 817.050 ;
        RECT 565.800 808.950 567.900 811.050 ;
        RECT 562.800 805.950 564.900 808.050 ;
        RECT 563.400 787.050 564.600 805.950 ;
        RECT 562.950 784.950 565.050 787.050 ;
        RECT 553.950 781.950 556.050 784.050 ;
        RECT 555.000 774.600 559.200 775.050 ;
        RECT 554.400 774.000 559.200 774.600 ;
        RECT 553.950 772.950 559.200 774.000 ;
        RECT 553.950 772.200 556.050 772.950 ;
        RECT 538.950 769.950 541.050 772.050 ;
        RECT 553.800 771.000 556.050 772.200 ;
        RECT 553.800 770.100 555.900 771.000 ;
        RECT 562.950 769.950 565.050 772.050 ;
        RECT 539.400 748.050 540.600 769.950 ;
        RECT 553.950 766.800 556.050 768.900 ;
        RECT 544.950 763.950 547.050 766.050 ;
        RECT 538.950 745.950 541.050 748.050 ;
        RECT 535.950 718.950 538.050 721.050 ;
        RECT 539.400 703.050 540.600 745.950 ;
        RECT 545.400 724.050 546.600 763.950 ;
        RECT 550.950 760.950 553.050 763.050 ;
        RECT 547.950 736.950 550.050 739.050 ;
        RECT 544.950 721.950 547.050 724.050 ;
        RECT 541.950 718.950 544.050 721.050 ;
        RECT 538.950 700.950 541.050 703.050 ;
        RECT 532.950 696.600 537.000 697.050 ;
        RECT 532.950 694.950 537.600 696.600 ;
        RECT 536.400 685.050 537.600 694.950 ;
        RECT 535.950 682.950 538.050 685.050 ;
        RECT 542.400 681.600 543.600 718.950 ;
        RECT 548.400 694.050 549.600 736.950 ;
        RECT 547.950 691.950 550.050 694.050 ;
        RECT 539.400 680.400 543.600 681.600 ;
        RECT 532.950 669.600 537.000 670.050 ;
        RECT 532.950 667.950 537.600 669.600 ;
        RECT 526.950 664.950 529.050 667.050 ;
        RECT 521.400 645.000 525.600 645.600 ;
        RECT 521.400 644.400 526.050 645.000 ;
        RECT 511.950 640.950 514.050 643.050 ;
        RECT 523.950 640.950 526.050 644.400 ;
        RECT 512.400 634.050 513.600 640.950 ;
        RECT 514.950 634.950 517.050 637.050 ;
        RECT 511.950 631.950 514.050 634.050 ;
        RECT 512.100 625.950 514.200 628.050 ;
        RECT 512.400 616.050 513.600 625.950 ;
        RECT 511.950 613.950 514.050 616.050 ;
        RECT 511.950 607.950 514.050 610.050 ;
        RECT 512.400 568.050 513.600 607.950 ;
        RECT 511.950 565.950 514.050 568.050 ;
        RECT 511.950 559.950 514.050 562.050 ;
        RECT 512.400 556.050 513.600 559.950 ;
        RECT 511.950 553.950 514.050 556.050 ;
        RECT 512.400 532.050 513.600 553.950 ;
        RECT 511.950 529.950 514.050 532.050 ;
        RECT 515.400 528.600 516.600 634.950 ;
        RECT 536.400 634.200 537.600 667.950 ;
        RECT 539.400 637.050 540.600 680.400 ;
        RECT 551.400 679.050 552.600 760.950 ;
        RECT 554.400 721.050 555.600 766.800 ;
        RECT 563.400 751.050 564.600 769.950 ;
        RECT 562.950 748.950 565.050 751.050 ;
        RECT 562.950 741.600 567.000 742.050 ;
        RECT 562.950 739.950 567.600 741.600 ;
        RECT 566.400 736.050 567.600 739.950 ;
        RECT 565.950 733.950 568.050 736.050 ;
        RECT 562.950 730.950 565.050 733.050 ;
        RECT 553.950 718.950 556.050 721.050 ;
        RECT 559.950 711.600 562.050 712.050 ;
        RECT 563.400 711.600 564.600 730.950 ;
        RECT 569.400 718.050 570.600 814.950 ;
        RECT 572.400 811.200 573.600 814.950 ;
        RECT 571.950 809.100 574.050 811.200 ;
        RECT 571.950 805.800 574.050 807.900 ;
        RECT 572.400 760.050 573.600 805.800 ;
        RECT 578.400 799.050 579.600 832.950 ;
        RECT 617.400 829.050 618.600 832.950 ;
        RECT 632.400 829.050 633.600 838.950 ;
        RECT 616.950 826.950 619.050 829.050 ;
        RECT 631.950 826.950 634.050 829.050 ;
        RECT 580.950 817.950 583.050 820.050 ;
        RECT 578.100 796.950 580.200 799.050 ;
        RECT 581.400 793.050 582.600 817.950 ;
        RECT 634.950 817.050 637.050 820.050 ;
        RECT 634.950 816.000 637.200 817.050 ;
        RECT 635.100 814.950 637.200 816.000 ;
        RECT 595.950 811.950 598.050 814.050 ;
        RECT 631.800 811.950 633.900 814.050 ;
        RECT 583.950 805.950 586.050 811.050 ;
        RECT 589.950 808.950 592.050 811.050 ;
        RECT 583.950 793.950 586.050 796.050 ;
        RECT 580.950 790.950 583.050 793.050 ;
        RECT 577.950 787.950 580.050 790.050 ;
        RECT 578.400 772.050 579.600 787.950 ;
        RECT 574.950 769.950 579.600 772.050 ;
        RECT 571.950 757.950 574.050 760.050 ;
        RECT 578.400 745.050 579.600 769.950 ;
        RECT 584.400 769.050 585.600 793.950 ;
        RECT 590.400 787.200 591.600 808.950 ;
        RECT 596.400 805.050 597.600 811.950 ;
        RECT 604.950 805.950 607.050 808.050 ;
        RECT 595.950 802.950 598.050 805.050 ;
        RECT 596.400 796.050 597.600 802.950 ;
        RECT 595.950 793.950 598.050 796.050 ;
        RECT 589.950 785.100 592.050 787.200 ;
        RECT 589.950 781.800 592.050 783.900 ;
        RECT 583.950 766.950 586.050 769.050 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 584.400 748.050 585.600 757.950 ;
        RECT 590.400 757.050 591.600 781.800 ;
        RECT 592.950 778.950 595.050 781.050 ;
        RECT 589.950 754.950 592.050 757.050 ;
        RECT 593.400 751.050 594.600 778.950 ;
        RECT 598.950 769.950 601.050 772.050 ;
        RECT 599.400 763.050 600.600 769.950 ;
        RECT 605.400 769.050 606.600 805.950 ;
        RECT 622.950 796.950 625.050 799.050 ;
        RECT 623.400 772.050 624.600 796.950 ;
        RECT 632.400 796.050 633.600 811.950 ;
        RECT 631.950 793.950 634.050 796.050 ;
        RECT 644.400 787.050 645.600 847.950 ;
        RECT 649.950 844.950 652.050 847.050 ;
        RECT 664.950 844.950 667.050 847.050 ;
        RECT 644.100 784.950 646.200 787.050 ;
        RECT 650.400 781.050 651.600 844.950 ;
        RECT 665.400 835.050 666.600 844.950 ;
        RECT 691.950 838.950 694.050 841.050 ;
        RECT 655.950 832.950 658.050 835.050 ;
        RECT 664.950 832.950 667.050 835.050 ;
        RECT 656.400 793.050 657.600 832.950 ;
        RECT 673.950 823.950 676.050 826.050 ;
        RECT 674.400 811.050 675.600 823.950 ;
        RECT 692.400 820.050 693.600 838.950 ;
        RECT 716.400 829.050 717.600 847.950 ;
        RECT 719.400 844.050 720.600 865.950 ;
        RECT 740.400 847.050 741.600 865.950 ;
        RECT 760.950 847.950 763.050 850.050 ;
        RECT 740.100 844.950 742.200 847.050 ;
        RECT 718.950 841.950 721.050 844.050 ;
        RECT 761.400 841.050 762.600 847.950 ;
        RECT 772.950 844.950 775.050 847.050 ;
        RECT 781.950 846.600 786.000 847.050 ;
        RECT 781.950 844.950 786.600 846.600 ;
        RECT 727.950 838.950 730.050 841.050 ;
        RECT 760.950 838.950 763.050 841.050 ;
        RECT 715.950 826.950 718.050 829.050 ;
        RECT 709.950 823.950 712.050 826.050 ;
        RECT 682.950 817.950 685.050 820.050 ;
        RECT 692.400 818.400 697.050 820.050 ;
        RECT 693.000 817.950 697.050 818.400 ;
        RECT 673.950 808.950 676.050 811.050 ;
        RECT 683.400 799.050 684.600 817.950 ;
        RECT 710.400 817.050 711.600 823.950 ;
        RECT 709.800 814.950 711.900 817.050 ;
        RECT 691.800 811.950 693.900 814.050 ;
        RECT 682.950 796.950 685.050 799.050 ;
        RECT 692.400 796.050 693.600 811.950 ;
        RECT 710.400 808.050 711.600 814.950 ;
        RECT 728.400 810.600 729.600 838.950 ;
        RECT 757.950 829.950 760.050 832.050 ;
        RECT 758.400 820.050 759.600 829.950 ;
        RECT 766.950 826.950 769.050 829.050 ;
        RECT 757.950 817.950 760.050 820.050 ;
        RECT 730.950 814.050 733.050 814.200 ;
        RECT 730.950 813.750 735.000 814.050 ;
        RECT 730.950 812.100 735.600 813.750 ;
        RECT 732.000 811.950 735.600 812.100 ;
        RECT 739.950 811.950 742.050 814.050 ;
        RECT 754.950 811.950 757.050 814.050 ;
        RECT 730.950 810.600 733.050 810.900 ;
        RECT 728.400 809.400 733.050 810.600 ;
        RECT 730.950 808.800 733.050 809.400 ;
        RECT 697.950 805.950 700.050 808.050 ;
        RECT 709.950 805.950 712.050 808.050 ;
        RECT 688.800 793.950 690.900 796.050 ;
        RECT 692.100 793.950 694.200 796.050 ;
        RECT 655.950 790.950 658.050 793.050 ;
        RECT 634.800 778.950 636.900 781.050 ;
        RECT 649.950 778.950 652.050 781.050 ;
        RECT 629.100 775.950 631.200 778.050 ;
        RECT 625.800 772.950 627.900 775.050 ;
        RECT 613.950 769.950 616.050 772.050 ;
        RECT 623.100 769.950 625.200 772.050 ;
        RECT 605.400 767.400 610.050 769.050 ;
        RECT 606.000 766.950 610.050 767.400 ;
        RECT 614.400 766.050 615.600 769.950 ;
        RECT 613.950 763.950 616.050 766.050 ;
        RECT 622.950 765.600 625.050 766.050 ;
        RECT 626.400 765.600 627.600 772.950 ;
        RECT 622.950 764.400 627.600 765.600 ;
        RECT 622.950 763.950 625.050 764.400 ;
        RECT 598.800 760.950 600.900 763.050 ;
        RECT 602.100 760.950 604.200 763.050 ;
        RECT 583.950 745.950 586.050 748.050 ;
        RECT 592.950 747.000 595.050 751.050 ;
        RECT 593.400 746.400 594.600 747.000 ;
        RECT 578.400 743.400 583.050 745.050 ;
        RECT 579.000 742.950 583.050 743.400 ;
        RECT 589.950 739.950 592.050 742.050 ;
        RECT 568.950 715.950 571.050 718.050 ;
        RECT 559.950 710.400 564.600 711.600 ;
        RECT 559.950 709.950 562.050 710.400 ;
        RECT 560.400 700.050 561.600 709.950 ;
        RECT 590.400 709.050 591.600 739.950 ;
        RECT 595.950 736.950 598.050 739.050 ;
        RECT 592.950 721.950 595.050 724.050 ;
        RECT 593.400 712.050 594.600 721.950 ;
        RECT 592.950 709.950 595.050 712.050 ;
        RECT 589.950 706.950 592.050 709.050 ;
        RECT 565.950 703.950 568.050 706.050 ;
        RECT 559.950 697.950 562.050 700.050 ;
        RECT 566.400 697.050 567.600 703.950 ;
        RECT 571.950 700.950 574.050 703.050 ;
        RECT 565.950 694.950 568.050 697.050 ;
        RECT 568.950 693.600 571.050 694.050 ;
        RECT 572.400 693.600 573.600 700.950 ;
        RECT 590.400 700.050 591.600 706.950 ;
        RECT 596.400 703.050 597.600 736.950 ;
        RECT 598.950 733.950 601.050 736.050 ;
        RECT 599.400 724.050 600.600 733.950 ;
        RECT 598.950 721.950 601.050 724.050 ;
        RECT 595.950 700.950 598.050 703.050 ;
        RECT 589.800 699.000 591.900 700.050 ;
        RECT 589.800 697.950 592.050 699.000 ;
        RECT 589.950 696.000 592.050 697.950 ;
        RECT 590.400 695.400 591.600 696.000 ;
        RECT 568.950 692.400 573.600 693.600 ;
        RECT 568.950 691.950 571.050 692.400 ;
        RECT 550.950 676.950 553.050 679.050 ;
        RECT 547.950 673.950 550.050 676.050 ;
        RECT 548.400 670.050 549.600 673.950 ;
        RECT 550.800 670.950 552.900 673.050 ;
        RECT 556.950 670.950 559.050 673.050 ;
        RECT 547.950 667.950 550.050 670.050 ;
        RECT 548.400 655.050 549.600 667.950 ;
        RECT 547.950 652.950 550.050 655.050 ;
        RECT 551.400 649.050 552.600 670.950 ;
        RECT 550.950 646.950 553.050 649.050 ;
        RECT 538.950 634.950 541.050 637.050 ;
        RECT 535.950 632.100 538.050 634.200 ;
        RECT 535.950 625.950 538.050 630.900 ;
        RECT 523.950 622.950 526.050 625.050 ;
        RECT 541.950 622.950 544.050 625.050 ;
        RECT 524.400 598.050 525.600 622.950 ;
        RECT 535.950 601.950 538.050 604.050 ;
        RECT 519.000 597.600 522.900 598.050 ;
        RECT 518.400 595.950 522.900 597.600 ;
        RECT 524.400 596.400 529.050 598.050 ;
        RECT 525.000 595.950 529.050 596.400 ;
        RECT 518.400 580.050 519.600 595.950 ;
        RECT 532.950 592.950 535.050 595.050 ;
        RECT 533.400 580.050 534.600 592.950 ;
        RECT 536.400 592.050 537.600 601.950 ;
        RECT 542.400 598.050 543.600 622.950 ;
        RECT 557.400 618.600 558.600 670.950 ;
        RECT 569.400 670.050 570.600 691.950 ;
        RECT 583.950 688.950 586.050 691.050 ;
        RECT 584.400 673.050 585.600 688.950 ;
        RECT 592.950 676.950 595.050 679.050 ;
        RECT 593.400 673.050 594.600 676.950 ;
        RECT 595.950 673.950 598.050 676.050 ;
        RECT 583.950 670.950 586.050 673.050 ;
        RECT 592.800 670.950 594.900 673.050 ;
        RECT 568.950 667.950 571.050 670.050 ;
        RECT 574.800 664.950 576.900 667.050 ;
        RECT 575.400 661.050 576.600 664.950 ;
        RECT 589.950 661.950 592.050 664.050 ;
        RECT 574.950 658.950 577.050 661.050 ;
        RECT 568.950 652.950 571.050 655.050 ;
        RECT 562.950 646.950 565.050 649.050 ;
        RECT 563.400 637.050 564.600 646.950 ;
        RECT 562.950 634.950 565.050 637.050 ;
        RECT 569.400 634.050 570.600 652.950 ;
        RECT 569.400 632.400 574.050 634.050 ;
        RECT 570.000 631.950 574.050 632.400 ;
        RECT 577.950 631.950 580.050 634.050 ;
        RECT 554.400 617.400 558.600 618.600 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 541.950 595.950 544.050 598.050 ;
        RECT 535.950 589.950 538.050 592.050 ;
        RECT 517.950 577.950 520.050 580.050 ;
        RECT 532.950 577.950 535.050 580.050 ;
        RECT 541.950 577.950 544.050 580.050 ;
        RECT 532.950 562.950 535.050 565.050 ;
        RECT 533.400 553.050 534.600 562.950 ;
        RECT 542.400 562.200 543.600 577.950 ;
        RECT 547.950 565.950 550.050 568.050 ;
        RECT 541.950 560.100 544.050 562.200 ;
        RECT 548.400 559.050 549.600 565.950 ;
        RECT 541.950 556.800 544.050 558.900 ;
        RECT 547.950 556.950 550.050 559.050 ;
        RECT 532.950 550.950 535.050 553.050 ;
        RECT 520.950 547.950 523.050 550.050 ;
        RECT 515.400 527.400 519.600 528.600 ;
        RECT 514.950 514.950 517.050 517.050 ;
        RECT 511.950 505.950 514.050 508.050 ;
        RECT 512.400 487.050 513.600 505.950 ;
        RECT 511.950 484.950 514.050 487.050 ;
        RECT 515.400 484.050 516.600 514.950 ;
        RECT 518.400 502.050 519.600 527.400 ;
        RECT 517.950 499.950 520.050 502.050 ;
        RECT 521.400 487.050 522.600 547.950 ;
        RECT 542.400 538.050 543.600 556.800 ;
        RECT 541.950 535.950 544.050 538.050 ;
        RECT 523.950 529.950 526.050 532.050 ;
        RECT 524.400 523.050 525.600 529.950 ;
        RECT 542.400 526.050 543.600 535.950 ;
        RECT 544.950 529.950 547.050 532.050 ;
        RECT 539.100 524.400 543.600 526.050 ;
        RECT 539.100 523.950 543.000 524.400 ;
        RECT 523.950 520.950 526.050 523.050 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 520.950 484.950 523.050 487.050 ;
        RECT 514.950 481.950 517.050 484.050 ;
        RECT 511.950 475.950 514.050 478.050 ;
        RECT 505.950 451.950 510.600 454.050 ;
        RECT 509.400 445.050 510.600 451.950 ;
        RECT 512.400 451.050 513.600 475.950 ;
        RECT 511.950 448.950 514.050 451.050 ;
        RECT 508.950 442.950 511.050 445.050 ;
        RECT 496.800 427.950 498.900 430.050 ;
        RECT 500.100 427.950 502.200 430.050 ;
        RECT 497.400 421.050 498.600 427.950 ;
        RECT 515.400 427.050 516.600 481.950 ;
        RECT 517.950 478.950 520.050 481.050 ;
        RECT 518.400 454.050 519.600 478.950 ;
        RECT 521.400 466.050 522.600 484.950 ;
        RECT 536.400 484.050 537.600 490.950 ;
        RECT 535.950 483.600 538.050 484.050 ;
        RECT 535.950 482.400 540.600 483.600 ;
        RECT 535.950 481.950 538.050 482.400 ;
        RECT 526.950 469.950 529.050 472.050 ;
        RECT 520.950 463.950 523.050 466.050 ;
        RECT 517.950 451.950 520.050 454.050 ;
        RECT 518.400 436.050 519.600 451.950 ;
        RECT 517.950 433.950 520.050 436.050 ;
        RECT 517.950 427.950 520.050 430.050 ;
        RECT 514.950 424.950 517.050 427.050 ;
        RECT 497.400 419.400 502.050 421.050 ;
        RECT 498.000 418.950 502.050 419.400 ;
        RECT 499.950 409.950 502.050 412.050 ;
        RECT 484.950 406.950 487.050 409.050 ;
        RECT 490.950 406.950 493.050 409.050 ;
        RECT 485.400 397.050 486.600 406.950 ;
        RECT 491.400 397.050 492.600 406.950 ;
        RECT 493.950 397.950 496.050 400.050 ;
        RECT 484.950 394.950 487.050 397.050 ;
        RECT 490.950 394.950 493.050 397.050 ;
        RECT 481.950 393.600 484.050 394.050 ;
        RECT 476.400 392.400 484.050 393.600 ;
        RECT 469.950 379.950 472.050 382.050 ;
        RECT 470.400 367.050 471.600 379.950 ;
        RECT 469.950 364.950 472.050 367.050 ;
        RECT 476.400 355.050 477.600 392.400 ;
        RECT 481.950 391.950 484.050 392.400 ;
        RECT 494.400 385.050 495.600 397.950 ;
        RECT 500.400 397.050 501.600 409.950 ;
        RECT 511.950 403.950 514.050 406.050 ;
        RECT 508.950 400.950 511.050 403.050 ;
        RECT 499.950 394.950 502.050 397.050 ;
        RECT 502.950 388.950 505.050 391.050 ;
        RECT 493.800 382.950 495.900 385.050 ;
        RECT 503.400 379.050 504.600 388.950 ;
        RECT 487.950 376.950 490.050 379.050 ;
        RECT 502.950 376.950 505.050 379.050 ;
        RECT 488.400 373.050 489.600 376.950 ;
        RECT 487.950 370.950 490.050 373.050 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 481.950 364.950 484.050 367.050 ;
        RECT 475.950 352.950 478.050 355.050 ;
        RECT 467.400 347.400 471.600 348.600 ;
        RECT 454.950 337.950 457.050 340.050 ;
        RECT 464.100 337.950 466.200 340.050 ;
        RECT 457.950 334.950 460.050 337.050 ;
        RECT 446.400 332.400 450.600 333.600 ;
        RECT 442.950 325.950 445.050 328.050 ;
        RECT 439.950 319.950 442.050 322.050 ;
        RECT 439.950 307.950 442.050 310.050 ;
        RECT 421.950 298.950 424.050 301.050 ;
        RECT 430.950 298.950 433.050 301.050 ;
        RECT 422.400 295.050 423.600 298.950 ;
        RECT 427.950 295.950 430.050 298.050 ;
        RECT 421.950 292.950 424.050 295.050 ;
        RECT 415.950 280.950 418.050 283.050 ;
        RECT 422.400 279.600 423.600 292.950 ;
        RECT 419.400 278.400 423.600 279.600 ;
        RECT 419.400 265.050 420.600 278.400 ;
        RECT 428.400 265.050 429.600 295.950 ;
        RECT 440.400 294.600 441.600 307.950 ;
        RECT 437.400 294.000 441.600 294.600 ;
        RECT 436.950 293.400 441.600 294.000 ;
        RECT 436.950 289.950 439.050 293.400 ;
        RECT 439.950 286.950 442.050 289.050 ;
        RECT 440.400 277.050 441.600 286.950 ;
        RECT 439.950 274.950 442.050 277.050 ;
        RECT 443.400 271.050 444.600 325.950 ;
        RECT 431.100 268.950 433.200 271.050 ;
        RECT 442.950 268.950 445.050 271.050 ;
        RECT 418.950 264.600 421.050 265.050 ;
        RECT 416.400 263.400 421.050 264.600 ;
        RECT 412.950 250.950 415.050 253.050 ;
        RECT 416.400 250.050 417.600 263.400 ;
        RECT 418.950 262.950 421.050 263.400 ;
        RECT 427.950 262.950 430.050 265.050 ;
        RECT 415.950 247.950 418.050 250.050 ;
        RECT 427.950 241.950 430.050 244.050 ;
        RECT 414.000 240.600 418.050 241.050 ;
        RECT 413.400 238.950 418.050 240.600 ;
        RECT 413.400 229.050 414.600 238.950 ;
        RECT 428.400 232.050 429.600 241.950 ;
        RECT 431.400 241.050 432.600 268.950 ;
        RECT 446.400 268.050 447.600 332.400 ;
        RECT 451.950 313.950 454.050 316.050 ;
        RECT 448.950 304.950 451.050 307.050 ;
        RECT 449.400 292.050 450.600 304.950 ;
        RECT 448.950 289.950 451.050 292.050 ;
        RECT 449.400 274.050 450.600 289.950 ;
        RECT 448.950 271.950 451.050 274.050 ;
        RECT 433.950 267.600 438.000 268.050 ;
        RECT 433.950 265.950 438.600 267.600 ;
        RECT 445.950 265.950 448.050 268.050 ;
        RECT 434.400 247.200 435.600 265.950 ;
        RECT 437.400 256.200 438.600 265.950 ;
        RECT 452.400 265.050 453.600 313.950 ;
        RECT 454.950 310.950 457.050 313.050 ;
        RECT 455.400 289.050 456.600 310.950 ;
        RECT 454.950 286.950 457.050 289.050 ;
        RECT 458.400 286.050 459.600 334.950 ;
        RECT 463.950 319.950 466.050 322.050 ;
        RECT 464.400 313.050 465.600 319.950 ;
        RECT 470.400 316.050 471.600 347.400 ;
        RECT 474.000 339.600 478.050 340.050 ;
        RECT 473.400 337.950 478.050 339.600 ;
        RECT 469.950 313.950 472.050 316.050 ;
        RECT 466.800 313.050 468.900 313.200 ;
        RECT 464.400 311.400 468.900 313.050 ;
        RECT 465.000 311.100 468.900 311.400 ;
        RECT 465.000 310.950 468.000 311.100 ;
        RECT 465.000 309.900 468.000 310.050 ;
        RECT 463.950 309.450 468.000 309.900 ;
        RECT 463.950 307.950 468.600 309.450 ;
        RECT 463.950 307.800 466.050 307.950 ;
        RECT 467.400 298.050 468.600 307.950 ;
        RECT 473.400 298.050 474.600 337.950 ;
        RECT 482.400 319.050 483.600 364.950 ;
        RECT 484.950 343.950 487.050 346.050 ;
        RECT 490.950 343.950 493.050 346.050 ;
        RECT 485.400 337.200 486.600 343.950 ;
        RECT 484.950 335.100 487.050 337.200 ;
        RECT 484.950 331.800 487.050 333.900 ;
        RECT 481.950 316.950 484.050 319.050 ;
        RECT 485.400 307.050 486.600 331.800 ;
        RECT 491.400 322.050 492.600 343.950 ;
        RECT 497.400 325.050 498.600 367.950 ;
        RECT 509.400 364.050 510.600 400.950 ;
        RECT 512.400 397.050 513.600 403.950 ;
        RECT 514.950 397.950 517.050 400.050 ;
        RECT 511.950 394.950 514.050 397.050 ;
        RECT 512.400 385.050 513.600 394.950 ;
        RECT 515.400 394.050 516.600 397.950 ;
        RECT 514.950 391.950 517.050 394.050 ;
        RECT 518.400 391.050 519.600 427.950 ;
        RECT 517.950 388.950 520.050 391.050 ;
        RECT 511.950 382.950 514.050 385.050 ;
        RECT 515.100 379.950 517.200 382.050 ;
        RECT 515.400 376.050 516.600 379.950 ;
        RECT 517.800 376.950 519.900 379.050 ;
        RECT 521.100 376.950 523.200 379.050 ;
        RECT 514.950 373.950 517.050 376.050 ;
        RECT 511.950 370.950 514.050 373.050 ;
        RECT 508.950 361.950 511.050 364.050 ;
        RECT 505.800 337.950 507.900 340.050 ;
        RECT 506.400 325.050 507.600 337.950 ;
        RECT 512.400 337.050 513.600 370.950 ;
        RECT 515.400 346.050 516.600 373.950 ;
        RECT 514.950 343.950 517.050 346.050 ;
        RECT 514.950 337.950 517.050 340.050 ;
        RECT 511.950 334.950 514.050 337.050 ;
        RECT 511.950 325.950 514.050 328.050 ;
        RECT 496.950 322.950 499.050 325.050 ;
        RECT 505.950 322.950 508.050 325.050 ;
        RECT 490.950 319.950 493.050 322.050 ;
        RECT 491.400 310.050 492.600 319.950 ;
        RECT 499.950 316.950 502.050 319.050 ;
        RECT 491.100 307.950 493.200 310.050 ;
        RECT 481.950 305.400 486.600 307.050 ;
        RECT 481.950 304.950 486.000 305.400 ;
        RECT 466.950 295.950 469.050 298.050 ;
        RECT 472.950 295.950 475.050 298.050 ;
        RECT 496.950 295.950 499.050 298.050 ;
        RECT 469.950 292.950 472.050 295.050 ;
        RECT 475.950 292.950 478.050 295.050 ;
        RECT 457.950 283.950 460.050 286.050 ;
        RECT 470.400 283.050 471.600 292.950 ;
        RECT 469.950 280.950 472.050 283.050 ;
        RECT 466.950 277.950 469.050 280.050 ;
        RECT 463.950 271.050 466.050 271.200 ;
        RECT 467.400 271.050 468.600 277.950 ;
        RECT 472.950 271.950 475.050 277.050 ;
        RECT 454.950 270.600 459.000 271.050 ;
        RECT 454.950 268.950 459.600 270.600 ;
        RECT 463.950 269.550 468.600 271.050 ;
        RECT 463.950 269.100 468.000 269.550 ;
        RECT 465.000 268.950 468.000 269.100 ;
        RECT 439.950 262.950 442.050 265.050 ;
        RECT 451.800 262.950 453.900 265.050 ;
        RECT 455.100 262.950 457.200 265.050 ;
        RECT 436.950 254.100 439.050 256.200 ;
        RECT 436.950 250.800 439.050 252.900 ;
        RECT 433.950 245.100 436.050 247.200 ;
        RECT 433.950 241.800 436.050 243.900 ;
        RECT 431.100 238.950 433.200 241.050 ;
        RECT 430.950 232.950 433.050 235.050 ;
        RECT 427.950 229.950 430.050 232.050 ;
        RECT 412.950 226.950 415.050 229.050 ;
        RECT 418.950 226.950 421.050 229.050 ;
        RECT 419.400 217.050 420.600 226.950 ;
        RECT 431.400 226.050 432.600 232.950 ;
        RECT 430.950 223.950 433.050 226.050 ;
        RECT 418.950 214.950 421.050 217.050 ;
        RECT 434.400 202.050 435.600 241.800 ;
        RECT 433.950 199.950 436.050 202.050 ;
        RECT 412.800 196.950 414.900 199.050 ;
        RECT 413.400 187.050 414.600 196.950 ;
        RECT 418.950 190.950 421.050 193.050 ;
        RECT 412.950 184.950 415.050 187.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 413.400 166.050 414.600 178.950 ;
        RECT 419.400 175.050 420.600 190.950 ;
        RECT 427.950 187.950 430.050 190.050 ;
        RECT 418.950 172.950 421.050 175.050 ;
        RECT 424.950 169.950 427.050 172.050 ;
        RECT 412.950 163.950 415.050 166.050 ;
        RECT 403.950 154.950 406.050 157.050 ;
        RECT 409.950 154.950 412.050 157.050 ;
        RECT 397.950 142.950 400.050 145.050 ;
        RECT 392.100 124.950 394.200 127.050 ;
        RECT 398.400 124.050 399.600 142.950 ;
        RECT 376.950 123.600 381.000 124.050 ;
        RECT 376.950 121.950 381.600 123.600 ;
        RECT 386.400 123.000 387.600 123.600 ;
        RECT 380.400 115.050 381.600 121.950 ;
        RECT 385.950 118.950 388.050 123.000 ;
        RECT 397.950 121.950 400.050 124.050 ;
        RECT 379.950 112.950 382.050 115.050 ;
        RECT 386.400 112.050 387.600 118.950 ;
        RECT 385.950 109.950 388.050 112.050 ;
        RECT 398.400 106.050 399.600 121.950 ;
        RECT 400.950 117.600 403.050 118.050 ;
        RECT 404.400 117.600 405.600 154.950 ;
        RECT 409.950 148.950 412.050 151.050 ;
        RECT 410.400 118.050 411.600 148.950 ;
        RECT 425.400 130.050 426.600 169.950 ;
        RECT 428.400 169.050 429.600 187.950 ;
        RECT 434.400 181.050 435.600 199.950 ;
        RECT 433.950 178.950 436.050 181.050 ;
        RECT 427.950 166.950 430.050 169.050 ;
        RECT 428.400 157.050 429.600 166.950 ;
        RECT 430.950 163.950 433.050 166.050 ;
        RECT 427.950 154.950 430.050 157.050 ;
        RECT 427.950 133.950 430.050 136.050 ;
        RECT 421.950 128.400 426.600 130.050 ;
        RECT 421.950 127.950 426.000 128.400 ;
        RECT 428.400 127.050 429.600 133.950 ;
        RECT 431.400 133.050 432.600 163.950 ;
        RECT 437.400 133.200 438.600 250.800 ;
        RECT 440.400 238.050 441.600 262.950 ;
        RECT 442.950 250.950 445.050 253.050 ;
        RECT 439.950 235.950 442.050 238.050 ;
        RECT 439.950 211.950 442.050 214.050 ;
        RECT 440.400 202.050 441.600 211.950 ;
        RECT 443.400 208.050 444.600 250.950 ;
        RECT 446.100 234.600 450.000 235.050 ;
        RECT 446.100 232.950 450.600 234.600 ;
        RECT 449.400 223.050 450.600 232.950 ;
        RECT 448.950 220.950 451.050 223.050 ;
        RECT 442.950 205.950 445.050 208.050 ;
        RECT 439.950 199.950 442.050 202.050 ;
        RECT 443.400 196.050 444.600 205.950 ;
        RECT 452.400 199.050 453.600 262.950 ;
        RECT 455.400 244.200 456.600 262.950 ;
        RECT 458.400 259.050 459.600 268.950 ;
        RECT 476.400 268.050 477.600 292.950 ;
        RECT 484.950 289.950 487.050 292.050 ;
        RECT 490.950 289.950 493.050 292.050 ;
        RECT 485.400 286.050 486.600 289.950 ;
        RECT 484.950 283.950 487.050 286.050 ;
        RECT 491.400 280.050 492.600 289.950 ;
        RECT 490.950 274.950 493.050 280.050 ;
        RECT 482.100 271.950 484.200 274.050 ;
        RECT 463.950 265.800 466.050 267.900 ;
        RECT 476.400 267.600 481.050 268.050 ;
        RECT 482.400 267.600 483.600 271.950 ;
        RECT 484.950 268.950 487.050 271.050 ;
        RECT 476.400 266.400 483.600 267.600 ;
        RECT 477.000 265.950 481.050 266.400 ;
        RECT 457.950 256.950 460.050 259.050 ;
        RECT 454.950 242.100 457.050 244.200 ;
        RECT 454.950 238.800 457.050 240.900 ;
        RECT 455.400 205.050 456.600 238.800 ;
        RECT 464.400 238.050 465.600 265.800 ;
        RECT 485.400 253.050 486.600 268.950 ;
        RECT 484.950 250.950 487.050 253.050 ;
        RECT 497.400 252.600 498.600 295.950 ;
        RECT 500.400 274.050 501.600 316.950 ;
        RECT 512.400 310.050 513.600 325.950 ;
        RECT 515.400 324.600 516.600 337.950 ;
        RECT 518.400 327.600 519.600 376.950 ;
        RECT 521.400 331.050 522.600 376.950 ;
        RECT 527.400 367.050 528.600 469.950 ;
        RECT 539.400 457.050 540.600 482.400 ;
        RECT 531.000 456.600 534.900 457.050 ;
        RECT 530.400 454.950 534.900 456.600 ;
        RECT 538.950 454.950 541.050 457.050 ;
        RECT 530.400 442.050 531.600 454.950 ;
        RECT 532.800 448.950 534.900 451.050 ;
        RECT 536.100 448.950 538.200 451.050 ;
        RECT 529.950 439.950 532.050 442.050 ;
        RECT 530.400 397.050 531.600 439.950 ;
        RECT 529.950 394.950 532.050 397.050 ;
        RECT 526.950 364.950 529.050 367.050 ;
        RECT 530.400 346.050 531.600 394.950 ;
        RECT 533.400 379.050 534.600 448.950 ;
        RECT 536.400 424.050 537.600 448.950 ;
        RECT 542.100 445.950 544.200 448.050 ;
        RECT 535.950 421.950 538.050 424.050 ;
        RECT 542.400 421.050 543.600 445.950 ;
        RECT 541.950 418.950 544.050 421.050 ;
        RECT 539.100 412.950 541.200 415.050 ;
        RECT 535.950 391.950 538.050 394.050 ;
        RECT 532.950 376.950 535.050 379.050 ;
        RECT 529.950 343.950 532.050 346.050 ;
        RECT 523.800 339.000 525.900 340.050 ;
        RECT 523.800 337.950 526.050 339.000 ;
        RECT 523.950 334.950 526.050 337.950 ;
        RECT 529.950 334.950 532.050 337.050 ;
        RECT 520.950 328.950 523.050 331.050 ;
        RECT 518.400 326.400 522.600 327.600 ;
        RECT 515.400 323.400 519.600 324.600 ;
        RECT 511.950 309.600 514.050 310.050 ;
        RECT 509.400 308.400 514.050 309.600 ;
        RECT 505.950 301.950 508.050 304.050 ;
        RECT 502.950 286.950 505.050 289.050 ;
        RECT 499.950 271.950 502.050 274.050 ;
        RECT 503.400 256.050 504.600 286.950 ;
        RECT 502.950 253.950 505.050 256.050 ;
        RECT 497.400 251.400 501.600 252.600 ;
        RECT 469.950 247.950 472.050 250.050 ;
        RECT 470.400 238.050 471.600 247.950 ;
        RECT 485.400 244.050 486.600 250.950 ;
        RECT 484.950 241.950 487.050 244.050 ;
        RECT 457.950 235.950 460.050 238.050 ;
        RECT 463.800 235.950 465.900 238.050 ;
        RECT 470.100 235.950 472.200 238.050 ;
        RECT 454.950 202.950 457.050 205.050 ;
        RECT 451.950 198.600 454.050 199.050 ;
        RECT 449.400 197.400 454.050 198.600 ;
        RECT 442.950 193.950 445.050 196.050 ;
        RECT 442.950 184.950 445.050 187.050 ;
        RECT 430.950 130.950 433.050 133.050 ;
        RECT 436.950 131.100 439.050 133.200 ;
        RECT 436.950 127.800 439.050 129.900 ;
        RECT 415.950 124.950 418.050 127.050 ;
        RECT 428.400 125.400 433.050 127.050 ;
        RECT 429.000 124.950 433.050 125.400 ;
        RECT 400.950 116.400 405.600 117.600 ;
        RECT 400.950 115.950 403.050 116.400 ;
        RECT 409.950 115.950 412.050 118.050 ;
        RECT 391.950 103.950 394.050 106.050 ;
        RECT 397.950 103.950 400.050 106.050 ;
        RECT 370.950 95.100 373.050 97.200 ;
        RECT 392.400 94.050 393.600 103.950 ;
        RECT 401.400 100.050 402.600 115.950 ;
        RECT 416.400 109.050 417.600 124.950 ;
        RECT 421.950 118.950 424.050 121.050 ;
        RECT 418.950 112.950 421.050 115.050 ;
        RECT 409.950 106.950 412.050 109.050 ;
        RECT 415.950 106.950 418.050 109.050 ;
        RECT 403.950 103.950 406.050 106.050 ;
        RECT 400.950 97.950 403.050 100.050 ;
        RECT 370.950 91.800 373.050 93.900 ;
        RECT 388.950 92.400 393.600 94.050 ;
        RECT 388.950 91.950 393.000 92.400 ;
        RECT 361.950 88.950 364.050 91.050 ;
        RECT 358.950 85.950 361.050 88.050 ;
        RECT 358.950 79.950 361.050 82.050 ;
        RECT 359.400 61.050 360.600 79.950 ;
        RECT 364.800 61.950 366.900 64.050 ;
        RECT 368.100 61.950 370.200 64.050 ;
        RECT 359.100 58.950 361.200 61.050 ;
        RECT 355.800 55.950 357.900 58.050 ;
        RECT 365.400 55.050 366.600 61.950 ;
        RECT 364.950 52.950 367.050 55.050 ;
        RECT 334.950 34.950 337.050 37.050 ;
        RECT 340.950 34.950 343.050 37.050 ;
        RECT 322.950 28.950 325.050 31.050 ;
        RECT 331.950 28.950 334.050 31.050 ;
        RECT 310.950 25.950 313.050 28.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 316.950 24.000 319.050 28.050 ;
        RECT 317.400 23.400 318.600 24.000 ;
        RECT 323.400 22.050 324.600 28.950 ;
        RECT 278.400 20.400 282.900 22.050 ;
        RECT 279.000 19.950 282.900 20.400 ;
        RECT 286.950 19.950 289.050 22.050 ;
        RECT 322.950 19.950 325.050 22.050 ;
        RECT 332.400 19.050 333.600 28.950 ;
        RECT 341.400 19.050 342.600 34.950 ;
        RECT 358.950 31.950 361.050 34.050 ;
        RECT 359.400 28.050 360.600 31.950 ;
        RECT 358.950 25.950 361.050 28.050 ;
        RECT 368.400 25.050 369.600 61.950 ;
        RECT 371.400 40.050 372.600 91.800 ;
        RECT 401.400 91.050 402.600 97.950 ;
        RECT 397.800 90.000 399.900 91.050 ;
        RECT 397.800 88.950 400.050 90.000 ;
        RECT 401.100 88.950 403.200 91.050 ;
        RECT 397.950 85.950 400.050 88.950 ;
        RECT 391.950 82.950 394.050 85.050 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 382.950 57.600 387.000 58.050 ;
        RECT 382.950 55.950 387.600 57.600 ;
        RECT 370.950 37.950 373.050 40.050 ;
        RECT 374.400 31.050 375.600 55.950 ;
        RECT 386.400 43.050 387.600 55.950 ;
        RECT 392.400 55.050 393.600 82.950 ;
        RECT 404.400 64.050 405.600 103.950 ;
        RECT 406.950 97.050 409.050 97.200 ;
        RECT 410.400 97.050 411.600 106.950 ;
        RECT 406.950 95.550 411.600 97.050 ;
        RECT 406.950 95.100 411.000 95.550 ;
        RECT 408.000 94.950 411.000 95.100 ;
        RECT 406.950 91.800 409.050 93.900 ;
        RECT 407.400 88.050 408.600 91.800 ;
        RECT 406.950 85.950 409.050 88.050 ;
        RECT 403.950 61.950 406.050 64.050 ;
        RECT 419.400 58.050 420.600 112.950 ;
        RECT 406.950 55.950 409.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 391.950 52.950 394.050 55.050 ;
        RECT 407.400 52.050 408.600 55.950 ;
        RECT 413.100 54.600 417.000 55.050 ;
        RECT 413.100 52.950 417.600 54.600 ;
        RECT 406.950 49.950 409.050 52.050 ;
        RECT 403.950 46.950 406.050 49.050 ;
        RECT 385.950 40.950 388.050 43.050 ;
        RECT 373.950 28.950 376.050 31.050 ;
        RECT 367.950 22.950 370.050 25.050 ;
        RECT 349.800 21.600 351.900 22.050 ;
        RECT 356.100 21.600 358.200 22.050 ;
        RECT 349.800 20.400 358.200 21.600 ;
        RECT 349.800 19.950 351.900 20.400 ;
        RECT 356.100 19.950 358.200 20.400 ;
        RECT 368.400 19.050 369.600 22.950 ;
        RECT 404.400 22.050 405.600 46.950 ;
        RECT 416.400 34.050 417.600 52.950 ;
        RECT 422.400 52.050 423.600 118.950 ;
        RECT 424.950 115.950 427.050 118.050 ;
        RECT 425.400 85.050 426.600 115.950 ;
        RECT 437.400 115.050 438.600 127.800 ;
        RECT 436.950 112.950 439.050 115.050 ;
        RECT 436.950 97.950 439.050 100.050 ;
        RECT 437.400 91.050 438.600 97.950 ;
        RECT 443.400 97.050 444.600 184.950 ;
        RECT 445.950 130.950 448.050 133.050 ;
        RECT 446.400 103.050 447.600 130.950 ;
        RECT 449.400 124.050 450.600 197.400 ;
        RECT 451.950 196.950 454.050 197.400 ;
        RECT 458.400 196.050 459.600 235.950 ;
        RECT 470.400 223.050 471.600 235.950 ;
        RECT 500.400 226.050 501.600 251.400 ;
        RECT 506.400 235.050 507.600 301.950 ;
        RECT 509.400 280.050 510.600 308.400 ;
        RECT 511.950 307.950 514.050 308.400 ;
        RECT 511.950 286.950 514.050 289.050 ;
        RECT 512.400 283.050 513.600 286.950 ;
        RECT 511.950 280.950 514.050 283.050 ;
        RECT 508.950 277.950 511.050 280.050 ;
        RECT 511.950 268.050 514.050 268.200 ;
        RECT 510.000 267.600 514.050 268.050 ;
        RECT 509.400 266.100 514.050 267.600 ;
        RECT 509.400 265.950 513.000 266.100 ;
        RECT 509.400 247.050 510.600 265.950 ;
        RECT 518.400 265.200 519.600 323.400 ;
        RECT 521.400 283.050 522.600 326.400 ;
        RECT 526.950 325.950 529.050 328.050 ;
        RECT 527.400 313.050 528.600 325.950 ;
        RECT 530.400 313.050 531.600 334.950 ;
        RECT 526.800 310.950 528.900 313.050 ;
        RECT 530.400 311.400 535.050 313.050 ;
        RECT 531.000 310.950 535.050 311.400 ;
        RECT 536.400 310.050 537.600 391.950 ;
        RECT 539.400 388.050 540.600 412.950 ;
        RECT 545.400 394.200 546.600 529.950 ;
        RECT 551.400 520.050 552.600 601.950 ;
        RECT 554.400 601.050 555.600 617.400 ;
        RECT 556.950 610.950 559.050 613.050 ;
        RECT 553.950 598.950 556.050 601.050 ;
        RECT 557.400 562.050 558.600 610.950 ;
        RECT 578.400 604.050 579.600 631.950 ;
        RECT 587.400 630.000 588.600 630.600 ;
        RECT 586.950 625.950 589.050 630.000 ;
        RECT 587.400 625.050 588.600 625.950 ;
        RECT 586.950 622.950 589.050 625.050 ;
        RECT 580.950 619.950 583.050 622.050 ;
        RECT 574.950 601.950 579.600 604.050 ;
        RECT 562.950 592.950 565.050 595.050 ;
        RECT 563.400 580.050 564.600 592.950 ;
        RECT 578.400 583.050 579.600 601.950 ;
        RECT 577.950 580.950 580.050 583.050 ;
        RECT 562.950 577.950 565.050 580.050 ;
        RECT 563.400 574.050 564.600 577.950 ;
        RECT 562.950 571.950 565.050 574.050 ;
        RECT 568.950 562.950 571.050 565.050 ;
        RECT 557.400 559.950 562.050 562.050 ;
        RECT 557.400 556.050 558.600 559.950 ;
        RECT 569.400 559.050 570.600 562.950 ;
        RECT 562.950 556.950 565.050 559.050 ;
        RECT 568.950 556.950 571.050 559.050 ;
        RECT 577.800 556.950 579.900 559.050 ;
        RECT 556.950 553.950 559.050 556.050 ;
        RECT 559.950 538.950 562.050 541.050 ;
        RECT 560.400 526.050 561.600 538.950 ;
        RECT 563.400 538.050 564.600 556.950 ;
        RECT 578.400 550.050 579.600 556.950 ;
        RECT 577.950 547.950 580.050 550.050 ;
        RECT 571.950 544.950 574.050 547.050 ;
        RECT 562.950 535.950 565.050 538.050 ;
        RECT 556.950 524.400 561.600 526.050 ;
        RECT 556.950 523.950 561.000 524.400 ;
        RECT 550.950 517.950 553.050 520.050 ;
        RECT 550.950 508.950 553.050 511.050 ;
        RECT 551.400 484.050 552.600 508.950 ;
        RECT 556.950 499.950 559.050 502.050 ;
        RECT 557.400 484.050 558.600 499.950 ;
        RECT 551.400 482.400 555.900 484.050 ;
        RECT 552.000 481.950 555.900 482.400 ;
        RECT 557.100 481.950 559.200 484.050 ;
        RECT 565.950 481.950 568.050 484.050 ;
        RECT 550.800 466.950 552.900 469.050 ;
        RECT 554.100 466.950 556.200 469.050 ;
        RECT 547.950 463.950 550.050 466.050 ;
        RECT 548.400 451.050 549.600 463.950 ;
        RECT 547.950 448.950 550.050 451.050 ;
        RECT 551.400 445.050 552.600 466.950 ;
        RECT 550.950 442.950 553.050 445.050 ;
        RECT 547.950 421.950 550.050 424.050 ;
        RECT 548.400 412.200 549.600 421.950 ;
        RECT 550.950 418.950 553.050 421.050 ;
        RECT 547.950 410.100 550.050 412.200 ;
        RECT 547.950 406.800 550.050 408.900 ;
        RECT 544.950 392.100 547.050 394.200 ;
        RECT 538.950 384.000 541.050 388.050 ;
        RECT 544.950 385.950 547.050 390.900 ;
        RECT 539.400 383.400 540.600 384.000 ;
        RECT 548.400 382.050 549.600 406.800 ;
        RECT 547.950 379.950 550.050 382.050 ;
        RECT 548.400 358.050 549.600 379.950 ;
        RECT 547.950 355.950 550.050 358.050 ;
        RECT 551.400 355.050 552.600 418.950 ;
        RECT 554.400 376.050 555.600 466.950 ;
        RECT 566.400 457.050 567.600 481.950 ;
        RECT 565.950 454.950 568.050 457.050 ;
        RECT 559.950 451.950 562.050 454.050 ;
        RECT 556.950 448.950 559.050 451.050 ;
        RECT 557.400 433.050 558.600 448.950 ;
        RECT 560.400 448.050 561.600 451.950 ;
        RECT 559.950 445.950 562.050 448.050 ;
        RECT 566.400 433.050 567.600 454.950 ;
        RECT 556.950 430.950 559.050 433.050 ;
        RECT 565.950 430.950 568.050 433.050 ;
        RECT 559.950 424.950 562.050 427.050 ;
        RECT 565.950 424.950 568.050 427.050 ;
        RECT 556.950 421.950 559.050 424.050 ;
        RECT 553.950 373.950 556.050 376.050 ;
        RECT 557.400 361.050 558.600 421.950 ;
        RECT 560.400 415.050 561.600 424.950 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 560.400 367.050 561.600 412.950 ;
        RECT 566.400 412.050 567.600 424.950 ;
        RECT 572.400 424.050 573.600 544.950 ;
        RECT 574.950 541.950 577.050 544.050 ;
        RECT 575.400 535.050 576.600 541.950 ;
        RECT 574.950 532.950 577.050 535.050 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 575.400 472.050 576.600 523.950 ;
        RECT 581.400 523.200 582.600 619.950 ;
        RECT 583.950 613.950 586.050 616.050 ;
        RECT 584.400 601.050 585.600 613.950 ;
        RECT 583.950 598.950 586.050 601.050 ;
        RECT 584.400 595.200 585.600 598.950 ;
        RECT 583.950 593.100 586.050 595.200 ;
        RECT 583.950 589.800 586.050 591.900 ;
        RECT 580.950 521.100 583.050 523.200 ;
        RECT 580.950 517.800 583.050 519.900 ;
        RECT 577.950 502.950 580.050 505.050 ;
        RECT 574.950 469.950 577.050 472.050 ;
        RECT 578.400 439.050 579.600 502.950 ;
        RECT 577.950 436.950 580.050 439.050 ;
        RECT 577.950 430.950 580.050 433.050 ;
        RECT 571.950 421.950 574.050 424.050 ;
        RECT 578.400 412.050 579.600 430.950 ;
        RECT 581.400 421.050 582.600 517.800 ;
        RECT 584.400 517.050 585.600 589.800 ;
        RECT 590.400 586.050 591.600 661.950 ;
        RECT 592.950 631.950 595.050 634.050 ;
        RECT 593.400 592.050 594.600 631.950 ;
        RECT 596.400 601.050 597.600 673.950 ;
        RECT 599.400 664.050 600.600 721.950 ;
        RECT 602.400 715.050 603.600 760.950 ;
        RECT 613.950 748.950 616.050 751.050 ;
        RECT 614.400 745.050 615.600 748.950 ;
        RECT 614.400 743.400 618.900 745.050 ;
        RECT 615.000 742.950 618.900 743.400 ;
        RECT 610.950 736.950 613.050 739.050 ;
        RECT 604.800 727.950 606.900 730.050 ;
        RECT 608.100 727.950 610.200 730.050 ;
        RECT 601.950 712.950 604.050 715.050 ;
        RECT 605.400 697.050 606.600 727.950 ;
        RECT 608.400 712.050 609.600 727.950 ;
        RECT 611.400 721.050 612.600 736.950 ;
        RECT 616.950 733.950 619.050 736.050 ;
        RECT 617.400 727.050 618.600 733.950 ;
        RECT 623.400 733.050 624.600 763.950 ;
        RECT 629.400 760.050 630.600 775.950 ;
        RECT 635.400 772.050 636.600 778.950 ;
        RECT 673.950 775.950 676.050 778.050 ;
        RECT 651.000 774.600 655.200 775.050 ;
        RECT 650.400 772.950 655.200 774.600 ;
        RECT 634.950 769.950 637.050 772.050 ;
        RECT 643.950 769.950 646.050 772.050 ;
        RECT 628.950 757.950 631.050 760.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 634.950 754.950 637.050 757.050 ;
        RECT 635.400 748.050 636.600 754.950 ;
        RECT 625.800 745.950 627.900 748.050 ;
        RECT 634.950 745.950 637.050 748.050 ;
        RECT 626.400 736.050 627.600 745.950 ;
        RECT 635.400 739.050 636.600 745.950 ;
        RECT 634.950 736.950 637.050 739.050 ;
        RECT 625.950 733.950 628.050 736.050 ;
        RECT 622.950 730.950 625.050 733.050 ;
        RECT 616.950 724.950 619.050 727.050 ;
        RECT 610.950 718.950 613.050 721.050 ;
        RECT 607.950 709.950 610.050 712.050 ;
        RECT 604.950 694.950 607.050 697.050 ;
        RECT 604.950 682.950 607.050 685.050 ;
        RECT 605.400 673.050 606.600 682.950 ;
        RECT 605.400 671.400 610.050 673.050 ;
        RECT 606.000 670.950 610.050 671.400 ;
        RECT 598.950 661.950 601.050 664.050 ;
        RECT 601.950 649.950 604.050 652.050 ;
        RECT 602.400 631.050 603.600 649.950 ;
        RECT 598.950 628.950 603.600 631.050 ;
        RECT 602.400 622.050 603.600 628.950 ;
        RECT 601.950 619.950 604.050 622.050 ;
        RECT 611.400 616.050 612.600 718.950 ;
        RECT 613.950 715.950 616.050 718.050 ;
        RECT 614.400 703.050 615.600 715.950 ;
        RECT 613.950 700.950 616.050 703.050 ;
        RECT 617.400 634.050 618.600 724.950 ;
        RECT 622.950 715.950 625.050 718.050 ;
        RECT 619.950 703.950 622.050 706.050 ;
        RECT 620.400 682.050 621.600 703.950 ;
        RECT 619.950 679.950 622.050 682.050 ;
        RECT 616.950 631.950 619.050 634.050 ;
        RECT 616.950 625.950 619.050 628.050 ;
        RECT 613.950 619.950 616.050 622.050 ;
        RECT 617.400 621.600 618.600 625.950 ;
        RECT 617.400 620.400 621.600 621.600 ;
        RECT 610.950 613.950 613.050 616.050 ;
        RECT 595.800 598.950 597.900 601.050 ;
        RECT 592.950 589.950 595.050 592.050 ;
        RECT 586.800 583.950 588.900 586.050 ;
        RECT 590.100 583.950 592.200 586.050 ;
        RECT 587.400 556.050 588.600 583.950 ;
        RECT 595.950 580.950 598.050 583.050 ;
        RECT 589.950 559.950 592.050 562.050 ;
        RECT 586.950 553.950 589.050 556.050 ;
        RECT 586.950 538.950 589.050 541.050 ;
        RECT 583.950 514.950 586.050 517.050 ;
        RECT 583.950 508.950 586.050 511.050 ;
        RECT 584.400 484.050 585.600 508.950 ;
        RECT 583.950 481.950 586.050 484.050 ;
        RECT 587.400 460.050 588.600 538.950 ;
        RECT 586.950 457.950 589.050 460.050 ;
        RECT 583.950 454.950 586.050 457.050 ;
        RECT 580.950 418.950 583.050 421.050 ;
        RECT 584.400 418.050 585.600 454.950 ;
        RECT 587.400 436.050 588.600 457.950 ;
        RECT 586.950 433.950 589.050 436.050 ;
        RECT 590.400 420.600 591.600 559.950 ;
        RECT 592.950 514.950 595.050 517.050 ;
        RECT 593.400 484.050 594.600 514.950 ;
        RECT 592.950 481.950 595.050 484.050 ;
        RECT 596.400 448.050 597.600 580.950 ;
        RECT 614.400 580.050 615.600 619.950 ;
        RECT 598.950 577.950 601.050 580.050 ;
        RECT 613.950 577.950 616.050 580.050 ;
        RECT 599.400 559.050 600.600 577.950 ;
        RECT 620.400 577.050 621.600 620.400 ;
        RECT 623.400 616.050 624.600 715.950 ;
        RECT 635.400 700.050 636.600 736.950 ;
        RECT 641.400 718.050 642.600 757.950 ;
        RECT 644.400 754.050 645.600 769.950 ;
        RECT 643.950 751.950 646.050 754.050 ;
        RECT 643.950 739.950 646.050 742.050 ;
        RECT 644.400 721.050 645.600 739.950 ;
        RECT 650.400 724.050 651.600 772.950 ;
        RECT 667.950 768.600 670.050 772.050 ;
        RECT 665.400 768.000 670.050 768.600 ;
        RECT 665.400 767.400 669.600 768.000 ;
        RECT 658.950 763.950 661.050 766.050 ;
        RECT 659.400 754.050 660.600 763.950 ;
        RECT 665.400 760.050 666.600 767.400 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 658.950 751.950 661.050 754.050 ;
        RECT 659.400 748.050 660.600 751.950 ;
        RECT 658.800 745.950 660.900 748.050 ;
        RECT 670.950 745.950 673.050 748.050 ;
        RECT 664.950 739.950 667.050 742.050 ;
        RECT 665.400 736.050 666.600 739.950 ;
        RECT 658.950 733.950 661.050 736.050 ;
        RECT 664.950 733.950 667.050 736.050 ;
        RECT 649.950 721.950 652.050 724.050 ;
        RECT 643.950 718.950 646.050 721.050 ;
        RECT 640.950 715.950 643.050 718.050 ;
        RECT 646.950 700.950 649.050 703.050 ;
        RECT 625.950 697.950 628.050 700.050 ;
        RECT 634.950 697.950 637.050 700.050 ;
        RECT 626.400 676.050 627.600 697.950 ;
        RECT 637.950 676.950 640.050 679.050 ;
        RECT 625.950 673.950 628.050 676.050 ;
        RECT 631.950 673.950 634.050 676.050 ;
        RECT 632.400 667.050 633.600 673.950 ;
        RECT 631.950 664.950 634.050 667.050 ;
        RECT 638.400 637.050 639.600 676.950 ;
        RECT 647.400 676.050 648.600 700.950 ;
        RECT 652.950 694.950 655.050 697.050 ;
        RECT 653.400 688.050 654.600 694.950 ;
        RECT 652.950 685.950 655.050 688.050 ;
        RECT 647.100 673.950 649.200 676.050 ;
        RECT 643.800 672.000 645.900 673.050 ;
        RECT 643.800 670.950 646.050 672.000 ;
        RECT 643.950 670.050 646.050 670.950 ;
        RECT 643.950 669.000 649.200 670.050 ;
        RECT 644.400 667.950 649.200 669.000 ;
        RECT 637.950 634.950 640.050 637.050 ;
        RECT 622.950 613.950 625.050 616.050 ;
        RECT 628.950 613.800 631.050 615.900 ;
        RECT 625.950 598.950 628.050 601.050 ;
        RECT 619.950 574.950 622.050 577.050 ;
        RECT 613.950 571.950 616.050 574.050 ;
        RECT 598.950 556.950 601.050 559.050 ;
        RECT 599.400 508.050 600.600 556.950 ;
        RECT 606.000 555.600 610.050 556.050 ;
        RECT 605.400 553.950 610.050 555.600 ;
        RECT 605.400 550.050 606.600 553.950 ;
        RECT 604.950 547.950 607.050 550.050 ;
        RECT 605.100 523.950 607.200 526.050 ;
        RECT 605.400 511.050 606.600 523.950 ;
        RECT 604.950 508.950 607.050 511.050 ;
        RECT 598.950 505.950 601.050 508.050 ;
        RECT 610.950 499.950 613.050 502.050 ;
        RECT 603.000 498.600 607.050 499.050 ;
        RECT 602.400 496.950 607.050 498.600 ;
        RECT 602.400 451.050 603.600 496.950 ;
        RECT 611.400 469.050 612.600 499.950 ;
        RECT 614.400 498.600 615.600 571.950 ;
        RECT 620.400 571.050 621.600 574.950 ;
        RECT 619.950 568.950 622.050 571.050 ;
        RECT 626.400 562.050 627.600 598.950 ;
        RECT 625.950 559.950 628.050 562.050 ;
        RECT 616.950 558.600 621.000 559.050 ;
        RECT 616.950 556.950 621.600 558.600 ;
        RECT 620.400 547.050 621.600 556.950 ;
        RECT 623.400 555.000 624.600 555.600 ;
        RECT 622.950 550.950 625.050 555.000 ;
        RECT 619.950 544.950 622.050 547.050 ;
        RECT 623.400 544.050 624.600 550.950 ;
        RECT 629.400 550.050 630.600 613.800 ;
        RECT 634.950 586.950 637.050 589.050 ;
        RECT 635.400 556.050 636.600 586.950 ;
        RECT 631.950 554.400 636.600 556.050 ;
        RECT 631.950 553.950 636.000 554.400 ;
        RECT 628.950 547.950 631.050 550.050 ;
        RECT 622.950 541.950 625.050 544.050 ;
        RECT 625.950 535.950 628.050 538.050 ;
        RECT 616.950 529.950 619.050 532.050 ;
        RECT 617.400 508.050 618.600 529.950 ;
        RECT 626.400 526.050 627.600 535.950 ;
        RECT 638.400 529.050 639.600 634.950 ;
        RECT 644.400 634.050 645.600 667.950 ;
        RECT 659.400 658.050 660.600 733.950 ;
        RECT 671.400 724.050 672.600 745.950 ;
        RECT 674.400 745.050 675.600 775.950 ;
        RECT 689.400 775.050 690.600 793.950 ;
        RECT 694.950 775.950 697.050 778.050 ;
        RECT 686.100 773.400 690.600 775.050 ;
        RECT 686.100 772.950 690.000 773.400 ;
        RECT 688.950 763.950 691.050 766.050 ;
        RECT 676.950 751.950 679.050 754.050 ;
        RECT 677.400 748.050 678.600 751.950 ;
        RECT 676.800 745.950 678.900 748.050 ;
        RECT 685.950 745.950 688.050 748.050 ;
        RECT 673.800 742.950 675.900 745.050 ;
        RECT 682.950 739.950 685.050 742.050 ;
        RECT 683.400 733.050 684.600 739.950 ;
        RECT 682.950 730.950 685.050 733.050 ;
        RECT 673.950 724.950 676.050 727.050 ;
        RECT 670.950 721.950 673.050 724.050 ;
        RECT 674.400 721.050 675.600 724.950 ;
        RECT 673.950 718.950 676.050 721.050 ;
        RECT 674.400 706.050 675.600 718.950 ;
        RECT 686.400 718.050 687.600 745.950 ;
        RECT 685.950 715.950 688.050 718.050 ;
        RECT 686.400 706.050 687.600 715.950 ;
        RECT 673.950 703.950 676.050 706.050 ;
        RECT 685.950 703.950 688.050 706.050 ;
        RECT 681.000 702.600 685.050 703.050 ;
        RECT 680.400 700.950 685.050 702.600 ;
        RECT 666.000 699.600 670.050 700.050 ;
        RECT 665.400 697.950 670.050 699.600 ;
        RECT 665.400 679.050 666.600 697.950 ;
        RECT 673.950 691.950 676.050 694.050 ;
        RECT 664.950 676.950 667.050 679.050 ;
        RECT 665.400 664.050 666.600 676.950 ;
        RECT 664.950 661.950 667.050 664.050 ;
        RECT 649.950 655.950 652.050 658.050 ;
        RECT 658.950 655.950 661.050 658.050 ;
        RECT 643.950 631.950 646.050 634.050 ;
        RECT 644.400 595.050 645.600 631.950 ;
        RECT 650.400 619.050 651.600 655.950 ;
        RECT 674.400 655.050 675.600 691.950 ;
        RECT 680.400 691.050 681.600 700.950 ;
        RECT 679.950 688.950 682.050 691.050 ;
        RECT 680.400 685.200 681.600 688.950 ;
        RECT 689.400 688.050 690.600 763.950 ;
        RECT 695.400 754.050 696.600 775.950 ;
        RECT 698.400 772.050 699.600 805.950 ;
        RECT 703.950 802.950 706.050 805.050 ;
        RECT 727.950 802.950 730.050 805.050 ;
        RECT 704.400 775.050 705.600 802.950 ;
        RECT 728.400 799.050 729.600 802.950 ;
        RECT 727.950 796.950 730.050 799.050 ;
        RECT 731.400 796.050 732.600 808.800 ;
        RECT 734.400 802.050 735.600 811.950 ;
        RECT 740.400 802.050 741.600 811.950 ;
        RECT 755.400 808.050 756.600 811.950 ;
        RECT 754.950 805.950 757.050 808.050 ;
        RECT 733.950 799.950 736.050 802.050 ;
        RECT 739.950 799.950 742.050 802.050 ;
        RECT 730.950 793.950 733.050 796.050 ;
        RECT 709.950 790.950 712.050 793.050 ;
        RECT 703.950 772.950 706.050 775.050 ;
        RECT 697.950 769.950 700.050 772.050 ;
        RECT 710.400 766.050 711.600 790.950 ;
        RECT 731.400 783.600 732.600 793.950 ;
        RECT 731.400 782.400 735.600 783.600 ;
        RECT 718.950 772.950 721.050 775.050 ;
        RECT 709.950 763.950 712.050 766.050 ;
        RECT 715.950 763.950 718.050 766.050 ;
        RECT 694.950 751.950 697.050 754.050 ;
        RECT 716.400 745.050 717.600 763.950 ;
        RECT 719.400 763.200 720.600 772.950 ;
        RECT 734.400 772.050 735.600 782.400 ;
        RECT 755.400 778.050 756.600 805.950 ;
        RECT 763.950 796.950 766.050 799.050 ;
        RECT 764.400 778.050 765.600 796.950 ;
        RECT 754.950 775.950 757.050 778.050 ;
        RECT 763.950 775.950 766.050 778.050 ;
        RECT 745.950 774.600 750.000 775.050 ;
        RECT 745.950 772.950 750.600 774.600 ;
        RECT 734.400 770.400 739.050 772.050 ;
        RECT 735.000 769.950 739.050 770.400 ;
        RECT 730.950 766.950 733.050 769.050 ;
        RECT 718.950 761.100 721.050 763.200 ;
        RECT 718.950 757.800 721.050 759.900 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 719.400 754.050 720.600 757.800 ;
        RECT 718.950 751.950 721.050 754.050 ;
        RECT 716.400 743.400 721.050 745.050 ;
        RECT 717.000 742.950 721.050 743.400 ;
        RECT 728.400 742.050 729.600 757.950 ;
        RECT 694.950 738.600 699.000 739.050 ;
        RECT 703.950 738.600 706.050 742.050 ;
        RECT 709.950 739.950 712.050 742.050 ;
        RECT 727.950 739.950 730.050 742.050 ;
        RECT 694.950 736.950 699.600 738.600 ;
        RECT 703.950 738.000 708.600 738.600 ;
        RECT 704.400 737.400 708.600 738.000 ;
        RECT 698.400 724.050 699.600 736.950 ;
        RECT 697.950 721.950 700.050 724.050 ;
        RECT 694.950 700.950 697.050 703.050 ;
        RECT 688.950 685.950 691.050 688.050 ;
        RECT 679.950 683.100 682.050 685.200 ;
        RECT 695.400 684.600 696.600 700.950 ;
        RECT 703.950 697.950 706.050 700.050 ;
        RECT 704.400 694.050 705.600 697.950 ;
        RECT 703.950 691.950 706.050 694.050 ;
        RECT 692.400 683.400 696.600 684.600 ;
        RECT 679.950 679.800 682.050 681.900 ;
        RECT 680.400 667.050 681.600 679.800 ;
        RECT 692.400 673.050 693.600 683.400 ;
        RECT 700.950 682.950 703.050 685.050 ;
        RECT 691.800 670.950 693.900 673.050 ;
        RECT 687.000 669.600 691.050 670.050 ;
        RECT 686.400 667.950 691.050 669.600 ;
        RECT 679.950 664.950 682.050 667.050 ;
        RECT 686.400 655.050 687.600 667.950 ;
        RECT 688.950 661.950 691.050 664.050 ;
        RECT 673.950 652.950 676.050 655.050 ;
        RECT 685.950 652.950 688.050 655.050 ;
        RECT 655.950 646.950 658.050 649.050 ;
        RECT 682.950 646.950 685.050 649.050 ;
        RECT 656.400 631.050 657.600 646.950 ;
        RECT 683.400 631.050 684.600 646.950 ;
        RECT 655.800 628.950 657.900 631.050 ;
        RECT 662.100 628.950 664.200 631.050 ;
        RECT 682.950 628.950 685.050 631.050 ;
        RECT 662.400 622.050 663.600 628.950 ;
        RECT 676.950 627.600 681.000 628.050 ;
        RECT 689.400 627.600 690.600 661.950 ;
        RECT 692.400 645.600 693.600 670.950 ;
        RECT 694.950 667.950 697.050 670.050 ;
        RECT 695.400 649.050 696.600 667.950 ;
        RECT 701.400 652.050 702.600 682.950 ;
        RECT 704.400 682.050 705.600 691.950 ;
        RECT 703.950 679.950 706.050 682.050 ;
        RECT 703.950 670.950 706.050 673.050 ;
        RECT 704.400 655.050 705.600 670.950 ;
        RECT 707.400 667.050 708.600 737.400 ;
        RECT 710.400 727.050 711.600 739.950 ;
        RECT 709.950 724.950 712.050 727.050 ;
        RECT 731.400 721.050 732.600 766.950 ;
        RECT 749.400 766.050 750.600 772.950 ;
        RECT 752.400 771.000 753.600 771.600 ;
        RECT 751.950 766.950 754.050 771.000 ;
        RECT 748.950 763.950 751.050 766.050 ;
        RECT 752.400 763.050 753.600 766.950 ;
        RECT 757.950 763.950 760.050 766.050 ;
        RECT 751.950 760.950 754.050 763.050 ;
        RECT 758.400 736.050 759.600 763.950 ;
        RECT 763.950 754.950 766.050 757.050 ;
        RECT 757.950 733.950 760.050 736.050 ;
        RECT 764.400 733.050 765.600 754.950 ;
        RECT 754.950 730.950 757.050 733.050 ;
        RECT 763.950 730.950 766.050 733.050 ;
        RECT 730.950 718.950 733.050 721.050 ;
        RECT 755.400 718.050 756.600 730.950 ;
        RECT 709.950 715.950 712.050 718.050 ;
        RECT 754.950 715.950 757.050 718.050 ;
        RECT 710.400 685.050 711.600 715.950 ;
        RECT 742.950 705.600 747.000 706.050 ;
        RECT 742.950 703.950 747.600 705.600 ;
        RECT 760.950 703.950 763.050 706.050 ;
        RECT 724.950 699.600 727.050 703.050 ;
        RECT 733.950 699.600 736.050 700.050 ;
        RECT 724.950 699.000 736.050 699.600 ;
        RECT 725.400 698.400 736.050 699.000 ;
        RECT 733.950 697.950 736.050 698.400 ;
        RECT 718.950 694.950 721.050 697.050 ;
        RECT 714.000 690.600 718.050 691.050 ;
        RECT 713.400 688.950 718.050 690.600 ;
        RECT 709.950 682.950 712.050 685.050 ;
        RECT 713.400 682.050 714.600 688.950 ;
        RECT 719.400 685.050 720.600 694.950 ;
        RECT 724.950 688.950 727.050 691.050 ;
        RECT 718.950 682.950 721.050 685.050 ;
        RECT 712.950 679.950 715.050 682.050 ;
        RECT 710.100 670.950 712.200 673.050 ;
        RECT 706.950 664.950 709.050 667.050 ;
        RECT 703.950 652.950 706.050 655.050 ;
        RECT 700.950 649.950 703.050 652.050 ;
        RECT 710.400 649.050 711.600 670.950 ;
        RECT 712.950 664.950 715.050 667.050 ;
        RECT 694.950 646.950 697.050 649.050 ;
        RECT 709.950 646.950 712.050 649.050 ;
        RECT 692.400 644.400 696.600 645.600 ;
        RECT 695.400 637.050 696.600 644.400 ;
        RECT 694.950 634.950 697.050 637.050 ;
        RECT 676.950 625.950 681.600 627.600 ;
        RECT 689.400 626.400 693.600 627.600 ;
        RECT 661.950 619.950 664.050 622.050 ;
        RECT 649.950 616.950 652.050 619.050 ;
        RECT 658.950 616.950 661.050 619.050 ;
        RECT 643.950 592.950 646.050 595.050 ;
        RECT 655.950 583.950 658.050 586.050 ;
        RECT 640.950 580.950 643.050 583.050 ;
        RECT 641.400 532.050 642.600 580.950 ;
        RECT 643.950 555.600 648.000 556.050 ;
        RECT 643.950 553.950 648.600 555.600 ;
        RECT 647.400 538.050 648.600 553.950 ;
        RECT 652.950 550.950 655.050 553.050 ;
        RECT 653.400 544.050 654.600 550.950 ;
        RECT 652.950 541.950 655.050 544.050 ;
        RECT 646.950 535.950 649.050 538.050 ;
        RECT 640.950 529.950 643.050 532.050 ;
        RECT 637.950 526.950 640.050 529.050 ;
        RECT 646.950 528.600 651.000 529.050 ;
        RECT 646.950 526.950 651.600 528.600 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 622.950 520.950 625.050 523.050 ;
        RECT 619.950 508.950 622.050 511.050 ;
        RECT 616.950 505.950 619.050 508.050 ;
        RECT 614.400 497.400 618.600 498.600 ;
        RECT 613.950 493.950 616.050 496.050 ;
        RECT 614.400 490.050 615.600 493.950 ;
        RECT 613.950 487.950 616.050 490.050 ;
        RECT 610.950 466.950 613.050 469.050 ;
        RECT 613.950 454.950 616.050 457.050 ;
        RECT 614.400 451.050 615.600 454.950 ;
        RECT 601.950 448.950 604.050 451.050 ;
        RECT 613.950 448.950 616.050 451.050 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 613.950 442.950 616.050 445.050 ;
        RECT 611.100 439.950 613.200 442.050 ;
        RECT 601.950 436.950 604.050 439.050 ;
        RECT 602.400 424.050 603.600 436.950 ;
        RECT 601.950 421.950 604.050 424.050 ;
        RECT 611.400 423.600 612.600 439.950 ;
        RECT 614.400 427.050 615.600 442.950 ;
        RECT 617.400 442.200 618.600 497.400 ;
        RECT 616.950 440.100 619.050 442.200 ;
        RECT 616.950 436.800 619.050 438.900 ;
        RECT 613.950 424.950 616.050 427.050 ;
        RECT 605.400 422.400 612.600 423.600 ;
        RECT 590.400 419.400 594.600 420.600 ;
        RECT 583.950 415.950 586.050 418.050 ;
        RECT 589.950 412.950 592.050 415.050 ;
        RECT 565.950 409.950 568.050 412.050 ;
        RECT 574.950 410.400 579.600 412.050 ;
        RECT 574.950 409.950 579.000 410.400 ;
        RECT 566.400 400.050 567.600 409.950 ;
        RECT 575.400 403.050 576.600 409.950 ;
        RECT 590.400 406.050 591.600 412.950 ;
        RECT 589.950 403.950 592.050 406.050 ;
        RECT 574.950 400.950 577.050 403.050 ;
        RECT 565.950 397.950 568.050 400.050 ;
        RECT 589.950 391.950 592.050 394.050 ;
        RECT 574.950 384.600 579.000 385.050 ;
        RECT 583.950 384.600 588.000 385.050 ;
        RECT 574.950 382.950 579.600 384.600 ;
        RECT 583.950 382.950 588.600 384.600 ;
        RECT 559.950 364.950 562.050 367.050 ;
        RECT 571.950 364.950 574.050 367.050 ;
        RECT 556.800 358.950 558.900 361.050 ;
        RECT 560.100 358.950 562.200 361.050 ;
        RECT 550.950 352.950 553.050 355.050 ;
        RECT 560.400 349.050 561.600 358.950 ;
        RECT 565.950 352.950 568.050 355.050 ;
        RECT 559.950 346.950 562.050 349.050 ;
        RECT 560.400 343.050 561.600 346.950 ;
        RECT 538.950 340.950 541.050 343.050 ;
        RECT 560.100 340.950 562.200 343.050 ;
        RECT 539.400 322.050 540.600 340.950 ;
        RECT 553.950 334.950 556.050 337.050 ;
        RECT 544.950 331.950 547.050 334.050 ;
        RECT 538.950 319.950 541.050 322.050 ;
        RECT 536.400 308.400 541.050 310.050 ;
        RECT 537.000 307.950 541.050 308.400 ;
        RECT 526.950 304.950 529.050 307.050 ;
        RECT 527.400 286.050 528.600 304.950 ;
        RECT 545.400 304.050 546.600 331.950 ;
        RECT 554.400 325.050 555.600 334.950 ;
        RECT 547.950 322.950 550.050 325.050 ;
        RECT 553.950 322.950 556.050 325.050 ;
        RECT 548.400 316.050 549.600 322.950 ;
        RECT 556.950 316.950 559.050 319.050 ;
        RECT 548.400 314.400 553.050 316.050 ;
        RECT 549.000 313.950 553.050 314.400 ;
        RECT 536.100 301.950 538.200 304.050 ;
        RECT 544.950 301.950 547.050 304.050 ;
        RECT 532.950 298.950 535.050 301.050 ;
        RECT 533.400 286.050 534.600 298.950 ;
        RECT 526.950 283.950 529.050 286.050 ;
        RECT 532.950 283.950 535.050 286.050 ;
        RECT 520.950 280.950 523.050 283.050 ;
        RECT 529.950 280.950 532.050 283.050 ;
        RECT 523.950 271.950 526.050 274.050 ;
        RECT 517.950 263.100 520.050 265.200 ;
        RECT 517.950 259.800 520.050 261.900 ;
        RECT 508.950 244.950 511.050 247.050 ;
        RECT 505.950 232.950 508.050 235.050 ;
        RECT 481.950 223.950 484.050 226.050 ;
        RECT 499.950 223.950 502.050 226.050 ;
        RECT 469.950 220.950 472.050 223.050 ;
        RECT 466.950 217.950 469.050 220.050 ;
        RECT 472.950 217.950 475.050 220.050 ;
        RECT 467.400 196.050 468.600 217.950 ;
        RECT 473.400 199.050 474.600 217.950 ;
        RECT 478.950 202.950 481.050 205.050 ;
        RECT 479.400 199.050 480.600 202.950 ;
        RECT 472.800 198.000 474.900 199.050 ;
        RECT 472.800 196.950 475.050 198.000 ;
        RECT 478.950 196.950 481.050 199.050 ;
        RECT 457.950 193.950 460.050 196.050 ;
        RECT 463.950 194.400 468.600 196.050 ;
        RECT 472.950 195.000 475.050 196.950 ;
        RECT 473.400 194.400 474.600 195.000 ;
        RECT 463.950 193.950 468.000 194.400 ;
        RECT 457.950 187.950 460.050 190.050 ;
        RECT 454.950 172.950 457.050 175.050 ;
        RECT 451.950 169.950 454.050 172.050 ;
        RECT 452.400 166.050 453.600 169.950 ;
        RECT 451.950 163.950 454.050 166.050 ;
        RECT 455.400 147.600 456.600 172.950 ;
        RECT 458.400 160.050 459.600 187.950 ;
        RECT 466.950 178.950 469.050 181.050 ;
        RECT 463.950 169.950 466.050 172.050 ;
        RECT 460.950 160.950 463.050 163.050 ;
        RECT 457.950 157.950 460.050 160.050 ;
        RECT 452.400 146.400 456.600 147.600 ;
        RECT 452.400 127.050 453.600 146.400 ;
        RECT 458.400 127.050 459.600 157.950 ;
        RECT 461.400 157.050 462.600 160.950 ;
        RECT 460.950 154.950 463.050 157.050 ;
        RECT 464.400 133.050 465.600 169.950 ;
        RECT 467.400 169.050 468.600 178.950 ;
        RECT 482.400 178.050 483.600 223.950 ;
        RECT 508.950 217.950 511.050 220.050 ;
        RECT 490.950 202.950 493.050 205.050 ;
        RECT 484.950 190.950 487.050 193.050 ;
        RECT 481.950 175.950 484.050 178.050 ;
        RECT 466.950 166.950 469.050 169.050 ;
        RECT 472.950 160.950 475.050 163.050 ;
        RECT 473.400 136.050 474.600 160.950 ;
        RECT 478.950 157.950 481.050 163.050 ;
        RECT 475.950 142.950 478.050 145.050 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 463.800 130.950 465.900 133.050 ;
        RECT 467.400 130.050 468.600 133.950 ;
        RECT 467.100 127.950 469.200 130.050 ;
        RECT 476.400 127.050 477.600 142.950 ;
        RECT 485.400 142.050 486.600 190.950 ;
        RECT 491.400 175.050 492.600 202.950 ;
        RECT 509.400 193.050 510.600 217.950 ;
        RECT 518.400 217.050 519.600 259.800 ;
        RECT 524.400 250.050 525.600 271.950 ;
        RECT 526.950 256.950 529.050 259.050 ;
        RECT 523.950 247.950 526.050 250.050 ;
        RECT 527.400 244.050 528.600 256.950 ;
        RECT 526.950 240.000 529.050 244.050 ;
        RECT 527.400 239.400 528.600 240.000 ;
        RECT 520.950 237.600 525.000 238.050 ;
        RECT 530.400 237.600 531.600 280.950 ;
        RECT 536.400 274.050 537.600 301.950 ;
        RECT 550.950 292.950 553.050 295.050 ;
        RECT 551.400 283.050 552.600 292.950 ;
        RECT 557.400 285.600 558.600 316.950 ;
        RECT 559.950 304.950 562.050 307.050 ;
        RECT 560.400 286.050 561.600 304.950 ;
        RECT 554.400 284.400 558.600 285.600 ;
        RECT 550.950 280.950 553.050 283.050 ;
        RECT 554.400 277.050 555.600 284.400 ;
        RECT 559.950 283.950 562.050 286.050 ;
        RECT 556.950 280.950 559.050 283.050 ;
        RECT 566.400 282.600 567.600 352.950 ;
        RECT 572.400 319.050 573.600 364.950 ;
        RECT 578.400 358.050 579.600 382.950 ;
        RECT 587.400 361.050 588.600 382.950 ;
        RECT 586.950 358.950 589.050 361.050 ;
        RECT 577.950 355.950 580.050 358.050 ;
        RECT 583.950 352.950 586.050 355.050 ;
        RECT 584.400 349.050 585.600 352.950 ;
        RECT 583.800 346.950 585.900 349.050 ;
        RECT 587.100 346.950 589.200 349.050 ;
        RECT 577.800 340.950 579.900 343.050 ;
        RECT 583.950 340.950 586.050 343.050 ;
        RECT 578.400 337.050 579.600 340.950 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 574.950 328.950 577.050 331.050 ;
        RECT 571.950 316.950 574.050 319.050 ;
        RECT 572.100 310.950 574.200 313.050 ;
        RECT 563.400 281.400 567.600 282.600 ;
        RECT 544.950 274.950 547.050 277.050 ;
        RECT 553.950 274.950 556.050 277.050 ;
        RECT 535.950 271.950 538.050 274.050 ;
        RECT 535.950 259.950 538.050 262.050 ;
        RECT 520.950 235.950 525.600 237.600 ;
        RECT 524.400 232.050 525.600 235.950 ;
        RECT 527.400 236.400 531.600 237.600 ;
        RECT 523.950 229.950 526.050 232.050 ;
        RECT 517.950 214.950 520.050 217.050 ;
        RECT 511.950 211.800 514.050 213.900 ;
        RECT 496.950 190.950 499.050 193.050 ;
        RECT 508.950 190.950 511.050 193.050 ;
        RECT 497.400 181.050 498.600 190.950 ;
        RECT 505.950 181.950 508.050 184.050 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 499.950 175.950 502.050 178.050 ;
        RECT 490.950 172.950 493.050 175.050 ;
        RECT 500.400 172.050 501.600 175.950 ;
        RECT 496.800 171.000 498.900 172.050 ;
        RECT 500.100 171.000 502.200 172.050 ;
        RECT 496.800 169.950 499.050 171.000 ;
        RECT 496.950 169.050 499.050 169.950 ;
        RECT 496.800 168.000 499.050 169.050 ;
        RECT 499.950 169.950 502.200 171.000 ;
        RECT 499.950 168.000 502.050 169.950 ;
        RECT 496.800 166.950 498.900 168.000 ;
        RECT 500.400 167.400 501.600 168.000 ;
        RECT 499.950 151.950 502.050 154.050 ;
        RECT 484.950 139.950 487.050 142.050 ;
        RECT 497.100 127.950 499.200 130.050 ;
        RECT 451.950 124.950 454.050 127.050 ;
        RECT 457.950 124.950 460.050 127.050 ;
        RECT 475.950 124.950 478.050 127.050 ;
        RECT 487.800 126.000 489.900 127.050 ;
        RECT 487.800 124.950 490.050 126.000 ;
        RECT 448.950 121.950 451.050 124.050 ;
        RECT 472.950 121.950 475.050 124.050 ;
        RECT 487.950 123.600 490.050 124.950 ;
        RECT 487.950 123.000 492.600 123.600 ;
        RECT 488.400 122.400 492.600 123.000 ;
        RECT 449.400 118.050 450.600 121.950 ;
        RECT 448.950 115.950 451.050 118.050 ;
        RECT 473.400 112.050 474.600 121.950 ;
        RECT 481.950 112.950 484.050 115.050 ;
        RECT 472.950 109.950 475.050 112.050 ;
        RECT 451.950 103.950 454.050 106.050 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 442.950 94.950 445.050 97.050 ;
        RECT 443.400 91.050 444.600 94.950 ;
        RECT 452.400 94.050 453.600 103.950 ;
        RECT 482.400 100.050 483.600 112.950 ;
        RECT 484.950 109.950 487.050 112.050 ;
        RECT 481.950 97.950 484.050 100.050 ;
        RECT 458.100 94.950 460.200 97.050 ;
        RECT 448.950 92.400 453.600 94.050 ;
        RECT 448.950 91.950 453.000 92.400 ;
        RECT 436.950 88.950 439.050 91.050 ;
        RECT 443.100 88.950 445.200 91.050 ;
        RECT 424.950 82.950 427.050 85.050 ;
        RECT 451.950 76.950 454.050 79.050 ;
        RECT 430.950 70.950 433.050 73.050 ;
        RECT 421.950 49.950 424.050 52.050 ;
        RECT 421.950 40.950 424.050 43.050 ;
        RECT 415.950 31.950 418.050 34.050 ;
        RECT 422.400 28.050 423.600 40.950 ;
        RECT 431.400 28.050 432.600 70.950 ;
        RECT 436.950 58.950 439.050 61.050 ;
        RECT 437.400 55.050 438.600 58.950 ;
        RECT 436.950 52.950 439.050 55.050 ;
        RECT 442.800 52.950 444.900 55.050 ;
        RECT 443.400 40.050 444.600 52.950 ;
        RECT 452.400 52.050 453.600 76.950 ;
        RECT 451.800 49.950 453.900 52.050 ;
        RECT 455.100 49.950 457.200 52.050 ;
        RECT 455.400 43.050 456.600 49.950 ;
        RECT 458.400 49.050 459.600 94.950 ;
        RECT 482.400 94.050 483.600 97.950 ;
        RECT 469.950 91.950 472.050 94.050 ;
        RECT 482.100 91.950 484.200 94.050 ;
        RECT 460.950 88.950 463.050 91.050 ;
        RECT 461.400 70.050 462.600 88.950 ;
        RECT 463.800 73.950 465.900 76.050 ;
        RECT 467.100 73.950 469.200 76.050 ;
        RECT 464.400 70.050 465.600 73.950 ;
        RECT 460.800 67.950 462.900 70.050 ;
        RECT 464.100 67.950 466.200 70.050 ;
        RECT 467.400 52.050 468.600 73.950 ;
        RECT 466.950 49.950 469.050 52.050 ;
        RECT 457.950 46.950 460.050 49.050 ;
        RECT 454.950 40.950 457.050 43.050 ;
        RECT 442.950 37.950 445.050 40.050 ;
        RECT 421.950 25.950 424.050 28.050 ;
        RECT 430.950 25.950 433.050 28.050 ;
        RECT 403.950 19.950 406.050 22.050 ;
        RECT 442.950 19.950 445.050 22.050 ;
        RECT 448.950 19.950 451.050 22.050 ;
        RECT 332.400 17.400 336.900 19.050 ;
        RECT 333.000 16.950 336.900 17.400 ;
        RECT 340.950 16.950 343.050 19.050 ;
        RECT 367.950 16.950 370.050 19.050 ;
        RECT 271.950 10.950 274.050 13.050 ;
        RECT 136.950 7.950 139.050 10.050 ;
        RECT 172.950 7.950 175.050 10.050 ;
        RECT 196.950 7.950 199.050 10.050 ;
        RECT 205.950 7.950 208.050 10.050 ;
        RECT 238.950 7.950 241.050 10.050 ;
        RECT 443.400 7.050 444.600 19.950 ;
        RECT 127.950 4.950 130.050 7.050 ;
        RECT 442.950 4.950 445.050 7.050 ;
        RECT 449.400 4.050 450.600 19.950 ;
        RECT 467.400 6.600 468.600 49.950 ;
        RECT 470.400 37.050 471.600 91.950 ;
        RECT 485.400 76.050 486.600 109.950 ;
        RECT 491.400 103.050 492.600 122.400 ;
        RECT 497.400 112.050 498.600 127.950 ;
        RECT 496.950 109.950 499.050 112.050 ;
        RECT 500.400 106.050 501.600 151.950 ;
        RECT 506.400 130.050 507.600 181.950 ;
        RECT 512.400 130.050 513.600 211.800 ;
        RECT 518.400 196.050 519.600 214.950 ;
        RECT 514.800 193.950 519.600 196.050 ;
        RECT 518.400 184.200 519.600 193.950 ;
        RECT 517.950 182.100 520.050 184.200 ;
        RECT 527.400 181.050 528.600 236.400 ;
        RECT 532.950 232.950 535.050 235.050 ;
        RECT 529.950 223.950 532.050 226.050 ;
        RECT 517.950 178.800 520.050 180.900 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 514.950 163.950 517.050 166.050 ;
        RECT 505.950 127.950 508.050 130.050 ;
        RECT 511.950 127.950 514.050 130.050 ;
        RECT 515.400 124.050 516.600 163.950 ;
        RECT 514.950 121.950 517.050 124.050 ;
        RECT 518.400 121.050 519.600 178.800 ;
        RECT 520.950 175.950 523.050 178.050 ;
        RECT 502.800 118.950 504.900 121.050 ;
        RECT 506.100 118.950 508.200 121.050 ;
        RECT 517.950 118.950 520.050 121.050 ;
        RECT 503.400 112.050 504.600 118.950 ;
        RECT 502.950 109.950 505.050 112.050 ;
        RECT 499.950 103.950 502.050 106.050 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 499.950 97.950 502.050 100.050 ;
        RECT 484.950 73.950 487.050 76.050 ;
        RECT 473.100 51.600 477.000 52.050 ;
        RECT 473.100 49.950 477.600 51.600 ;
        RECT 476.400 40.050 477.600 49.950 ;
        RECT 484.950 46.950 487.050 49.050 ;
        RECT 475.950 37.950 478.050 40.050 ;
        RECT 469.950 34.950 472.050 37.050 ;
        RECT 485.400 25.050 486.600 46.950 ;
        RECT 500.400 28.050 501.600 97.950 ;
        RECT 499.950 25.950 502.050 28.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 506.400 22.050 507.600 118.950 ;
        RECT 517.950 112.950 520.050 115.050 ;
        RECT 511.950 106.950 514.050 109.050 ;
        RECT 508.950 103.950 511.050 106.050 ;
        RECT 509.400 31.050 510.600 103.950 ;
        RECT 512.400 94.050 513.600 106.950 ;
        RECT 518.400 94.050 519.600 112.950 ;
        RECT 521.400 100.050 522.600 175.950 ;
        RECT 526.950 172.950 529.050 175.050 ;
        RECT 527.400 166.050 528.600 172.950 ;
        RECT 524.100 164.400 528.600 166.050 ;
        RECT 524.100 163.950 528.000 164.400 ;
        RECT 524.400 127.200 525.600 163.950 ;
        RECT 530.400 139.050 531.600 223.950 ;
        RECT 533.400 142.050 534.600 232.950 ;
        RECT 532.950 139.950 535.050 142.050 ;
        RECT 529.950 136.950 532.050 139.050 ;
        RECT 536.400 130.050 537.600 259.950 ;
        RECT 538.950 232.950 541.050 235.050 ;
        RECT 535.950 127.950 538.050 130.050 ;
        RECT 523.800 125.100 525.900 127.200 ;
        RECT 539.400 127.050 540.600 232.950 ;
        RECT 545.400 214.050 546.600 274.950 ;
        RECT 550.950 271.050 553.050 274.050 ;
        RECT 557.400 271.050 558.600 280.950 ;
        RECT 550.950 270.000 553.200 271.050 ;
        RECT 551.100 268.950 553.200 270.000 ;
        RECT 556.950 268.950 559.050 271.050 ;
        RECT 563.400 270.600 564.600 281.400 ;
        RECT 565.950 277.950 568.050 280.050 ;
        RECT 560.400 270.000 564.600 270.600 ;
        RECT 559.950 269.400 564.600 270.000 ;
        RECT 566.400 271.050 567.600 277.950 ;
        RECT 572.400 274.050 573.600 310.950 ;
        RECT 575.400 310.050 576.600 328.950 ;
        RECT 584.400 310.050 585.600 340.950 ;
        RECT 587.400 340.050 588.600 346.950 ;
        RECT 586.950 337.950 589.050 340.050 ;
        RECT 590.400 334.050 591.600 391.950 ;
        RECT 589.950 331.950 592.050 334.050 ;
        RECT 586.950 322.950 589.050 325.050 ;
        RECT 575.400 308.400 580.050 310.050 ;
        RECT 576.000 307.950 580.050 308.400 ;
        RECT 583.800 307.950 585.900 310.050 ;
        RECT 574.950 304.800 577.050 306.900 ;
        RECT 575.400 295.050 576.600 304.800 ;
        RECT 574.950 292.950 577.050 295.050 ;
        RECT 583.950 285.600 586.050 286.050 ;
        RECT 587.400 285.600 588.600 322.950 ;
        RECT 593.400 313.050 594.600 419.400 ;
        RECT 602.400 415.050 603.600 421.950 ;
        RECT 601.950 412.950 604.050 415.050 ;
        RECT 598.950 379.950 601.050 382.050 ;
        RECT 599.400 358.200 600.600 379.950 ;
        RECT 601.950 367.950 604.050 370.050 ;
        RECT 598.950 356.100 601.050 358.200 ;
        RECT 598.950 352.800 601.050 354.900 ;
        RECT 595.950 349.950 598.050 352.050 ;
        RECT 596.400 346.050 597.600 349.950 ;
        RECT 595.950 343.950 598.050 346.050 ;
        RECT 595.950 322.950 598.050 325.050 ;
        RECT 596.400 319.050 597.600 322.950 ;
        RECT 599.400 319.050 600.600 352.800 ;
        RECT 602.400 325.050 603.600 367.950 ;
        RECT 605.400 337.050 606.600 422.400 ;
        RECT 607.950 415.950 610.050 421.050 ;
        RECT 613.950 418.950 616.050 421.050 ;
        RECT 608.100 411.600 612.000 412.050 ;
        RECT 608.100 409.950 612.600 411.600 ;
        RECT 607.950 400.950 610.050 403.050 ;
        RECT 608.400 394.050 609.600 400.950 ;
        RECT 607.800 391.950 609.900 394.050 ;
        RECT 611.400 388.050 612.600 409.950 ;
        RECT 610.950 385.950 613.050 388.050 ;
        RECT 614.400 385.050 615.600 418.950 ;
        RECT 617.400 415.050 618.600 436.800 ;
        RECT 620.400 433.050 621.600 508.950 ;
        RECT 623.400 433.050 624.600 520.950 ;
        RECT 638.400 520.050 639.600 526.950 ;
        RECT 637.950 517.950 640.050 520.050 ;
        RECT 634.950 502.950 637.050 505.050 ;
        RECT 625.950 487.950 628.050 490.050 ;
        RECT 626.400 451.050 627.600 487.950 ;
        RECT 635.400 484.050 636.600 502.950 ;
        RECT 638.400 496.050 639.600 517.950 ;
        RECT 650.400 496.050 651.600 526.950 ;
        RECT 656.400 505.050 657.600 583.950 ;
        RECT 655.950 502.950 658.050 505.050 ;
        RECT 659.400 499.050 660.600 616.950 ;
        RECT 680.400 610.050 681.600 625.950 ;
        RECT 679.950 607.950 682.050 610.050 ;
        RECT 692.400 607.050 693.600 626.400 ;
        RECT 700.950 625.950 703.050 628.050 ;
        RECT 710.100 627.600 712.200 628.050 ;
        RECT 713.400 627.600 714.600 664.950 ;
        RECT 719.400 655.050 720.600 682.950 ;
        RECT 725.400 679.050 726.600 688.950 ;
        RECT 746.400 679.050 747.600 703.950 ;
        RECT 724.950 676.950 727.050 679.050 ;
        RECT 745.950 676.950 748.050 679.050 ;
        RECT 757.950 676.950 760.050 679.050 ;
        RECT 730.950 670.950 733.050 673.050 ;
        RECT 718.950 652.950 721.050 655.050 ;
        RECT 731.400 649.050 732.600 670.950 ;
        RECT 736.950 661.950 739.050 667.050 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 718.950 634.950 721.050 637.050 ;
        RECT 710.100 626.400 714.600 627.600 ;
        RECT 710.100 625.950 712.200 626.400 ;
        RECT 673.950 601.950 676.050 607.050 ;
        RECT 682.950 603.600 685.050 607.050 ;
        RECT 691.950 604.950 694.050 607.050 ;
        RECT 682.950 603.000 687.600 603.600 ;
        RECT 683.400 602.400 687.600 603.000 ;
        RECT 667.950 592.950 670.050 595.050 ;
        RECT 676.950 592.950 679.050 595.050 ;
        RECT 668.400 556.050 669.600 592.950 ;
        RECT 670.950 589.950 673.050 592.050 ;
        RECT 671.400 583.050 672.600 589.950 ;
        RECT 677.400 589.050 678.600 592.950 ;
        RECT 676.950 586.950 679.050 589.050 ;
        RECT 670.800 580.950 672.900 583.050 ;
        RECT 674.100 580.950 676.200 583.050 ;
        RECT 667.950 555.600 672.000 556.050 ;
        RECT 667.950 553.950 672.600 555.600 ;
        RECT 664.950 541.950 667.050 544.050 ;
        RECT 665.400 535.050 666.600 541.950 ;
        RECT 671.400 541.050 672.600 553.950 ;
        RECT 670.950 538.950 673.050 541.050 ;
        RECT 664.950 532.950 667.050 535.050 ;
        RECT 658.800 496.950 660.900 499.050 ;
        RECT 637.950 493.950 640.050 496.050 ;
        RECT 649.950 493.950 652.050 496.050 ;
        RECT 655.950 493.950 658.050 496.050 ;
        RECT 638.400 487.050 639.600 493.950 ;
        RECT 643.950 490.950 646.050 493.050 ;
        RECT 638.100 484.950 640.200 487.050 ;
        RECT 644.400 484.050 645.600 490.950 ;
        RECT 656.400 487.050 657.600 493.950 ;
        RECT 656.400 485.400 661.050 487.050 ;
        RECT 657.000 484.950 661.050 485.400 ;
        RECT 634.950 481.950 637.050 484.050 ;
        RECT 644.400 482.400 649.050 484.050 ;
        RECT 645.000 481.950 649.050 482.400 ;
        RECT 665.400 478.050 666.600 532.950 ;
        RECT 667.950 522.600 672.000 523.050 ;
        RECT 667.950 520.950 672.600 522.600 ;
        RECT 671.400 517.200 672.600 520.950 ;
        RECT 670.950 515.100 673.050 517.200 ;
        RECT 670.950 511.800 673.050 513.900 ;
        RECT 671.400 490.050 672.600 511.800 ;
        RECT 670.950 487.950 673.050 490.050 ;
        RECT 646.950 475.950 649.050 478.050 ;
        RECT 664.950 475.950 667.050 478.050 ;
        RECT 643.950 472.950 646.050 475.050 ;
        RECT 634.800 460.950 636.900 463.050 ;
        RECT 635.400 451.050 636.600 460.950 ;
        RECT 625.950 448.950 628.050 451.050 ;
        RECT 634.950 448.950 637.050 451.050 ;
        RECT 625.950 442.950 628.050 445.050 ;
        RECT 619.800 430.950 621.900 433.050 ;
        RECT 623.100 430.950 625.200 433.050 ;
        RECT 626.400 417.600 627.600 442.950 ;
        RECT 644.400 439.050 645.600 472.950 ;
        RECT 647.400 454.050 648.600 475.950 ;
        RECT 674.400 475.050 675.600 580.950 ;
        RECT 676.950 574.950 679.050 577.050 ;
        RECT 677.400 478.050 678.600 574.950 ;
        RECT 686.400 559.050 687.600 602.400 ;
        RECT 701.400 595.050 702.600 625.950 ;
        RECT 710.400 613.050 711.600 625.950 ;
        RECT 709.950 610.950 712.050 613.050 ;
        RECT 712.950 607.950 715.050 610.050 ;
        RECT 709.950 604.950 712.050 607.050 ;
        RECT 706.950 598.950 709.050 601.050 ;
        RECT 692.100 592.950 694.200 595.050 ;
        RECT 700.950 592.950 703.050 595.050 ;
        RECT 692.400 577.050 693.600 592.950 ;
        RECT 691.950 574.950 694.050 577.050 ;
        RECT 685.950 556.950 688.050 559.050 ;
        RECT 679.950 555.600 684.000 556.050 ;
        RECT 679.950 553.950 684.600 555.600 ;
        RECT 683.400 538.050 684.600 553.950 ;
        RECT 682.950 535.950 685.050 538.050 ;
        RECT 679.950 526.950 682.050 529.050 ;
        RECT 680.400 496.050 681.600 526.950 ;
        RECT 692.400 526.050 693.600 574.950 ;
        RECT 707.400 574.050 708.600 598.950 ;
        RECT 710.400 586.050 711.600 604.950 ;
        RECT 710.100 583.950 712.200 586.050 ;
        RECT 706.950 571.950 709.050 574.050 ;
        RECT 713.400 556.050 714.600 607.950 ;
        RECT 719.400 607.050 720.600 634.950 ;
        RECT 730.950 622.950 733.050 625.050 ;
        RECT 736.950 622.950 739.050 625.050 ;
        RECT 727.950 613.950 730.050 616.050 ;
        RECT 718.950 604.950 721.050 607.050 ;
        RECT 728.400 604.050 729.600 613.950 ;
        RECT 727.950 601.950 730.050 604.050 ;
        RECT 731.400 601.050 732.600 622.950 ;
        RECT 737.400 610.050 738.600 622.950 ;
        RECT 746.400 610.050 747.600 676.950 ;
        RECT 754.950 667.950 757.050 670.050 ;
        RECT 751.950 664.950 754.050 667.050 ;
        RECT 752.400 652.050 753.600 664.950 ;
        RECT 755.400 664.050 756.600 667.950 ;
        RECT 754.950 661.950 757.050 664.050 ;
        RECT 751.950 649.950 754.050 652.050 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 755.400 628.050 756.600 646.950 ;
        RECT 751.800 625.950 753.900 628.050 ;
        RECT 755.100 625.950 757.200 628.050 ;
        RECT 736.950 607.950 739.050 610.050 ;
        RECT 745.950 607.950 748.050 610.050 ;
        RECT 721.950 598.950 724.050 601.050 ;
        RECT 731.100 598.950 733.200 601.050 ;
        RECT 722.400 574.050 723.600 598.950 ;
        RECT 724.950 595.950 727.050 598.050 ;
        RECT 725.400 589.050 726.600 595.950 ;
        RECT 724.950 586.950 727.050 589.050 ;
        RECT 727.950 583.950 730.050 586.050 ;
        RECT 721.950 571.950 724.050 574.050 ;
        RECT 703.950 555.600 708.000 556.050 ;
        RECT 703.950 553.950 708.600 555.600 ;
        RECT 713.400 554.400 718.050 556.050 ;
        RECT 714.000 553.950 718.050 554.400 ;
        RECT 722.100 553.950 724.200 556.050 ;
        RECT 707.400 544.050 708.600 553.950 ;
        RECT 716.400 547.050 717.600 553.950 ;
        RECT 715.950 544.950 718.050 547.050 ;
        RECT 706.950 541.950 709.050 544.050 ;
        RECT 712.950 541.950 715.050 544.050 ;
        RECT 718.950 541.950 721.050 544.050 ;
        RECT 709.950 529.950 712.050 532.050 ;
        RECT 688.950 523.950 693.600 526.050 ;
        RECT 692.400 520.050 693.600 523.950 ;
        RECT 710.400 523.050 711.600 529.950 ;
        RECT 706.950 520.950 711.600 523.050 ;
        RECT 691.950 517.950 694.050 520.050 ;
        RECT 685.950 514.950 688.050 517.050 ;
        RECT 686.400 508.050 687.600 514.950 ;
        RECT 710.400 511.050 711.600 520.950 ;
        RECT 709.950 508.950 712.050 511.050 ;
        RECT 685.950 505.950 688.050 508.050 ;
        RECT 679.950 493.950 682.050 496.050 ;
        RECT 682.950 484.950 685.050 487.050 ;
        RECT 676.950 475.950 679.050 478.050 ;
        RECT 673.950 472.950 676.050 475.050 ;
        RECT 661.950 469.950 664.050 472.050 ;
        RECT 652.950 457.950 655.050 460.050 ;
        RECT 646.800 451.950 648.900 454.050 ;
        RECT 644.100 436.950 646.200 439.050 ;
        RECT 647.400 436.050 648.600 451.950 ;
        RECT 653.400 441.600 654.600 457.950 ;
        RECT 662.400 454.050 663.600 469.950 ;
        RECT 664.950 463.950 667.050 466.050 ;
        RECT 665.400 457.050 666.600 463.950 ;
        RECT 676.950 460.950 679.050 463.050 ;
        RECT 664.950 454.950 667.050 457.050 ;
        RECT 661.950 451.950 664.050 454.050 ;
        RECT 665.400 448.050 666.600 454.950 ;
        RECT 672.000 450.600 675.900 451.050 ;
        RECT 671.400 448.950 675.900 450.600 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 671.400 442.050 672.600 448.950 ;
        RECT 650.400 440.400 654.600 441.600 ;
        RECT 637.950 433.950 640.050 436.050 ;
        RECT 646.950 433.950 649.050 436.050 ;
        RECT 638.400 418.050 639.600 433.950 ;
        RECT 623.400 416.400 627.600 417.600 ;
        RECT 616.950 412.950 619.050 415.050 ;
        RECT 619.950 406.950 622.050 409.050 ;
        RECT 620.400 385.050 621.600 406.950 ;
        RECT 607.950 382.950 610.050 385.050 ;
        RECT 613.800 382.950 615.900 385.050 ;
        RECT 619.800 382.950 621.900 385.050 ;
        RECT 608.400 363.600 609.600 382.950 ;
        RECT 623.400 373.050 624.600 416.400 ;
        RECT 637.950 415.950 640.050 418.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 625.950 409.950 628.050 412.050 ;
        RECT 626.400 406.050 627.600 409.950 ;
        RECT 625.950 403.950 628.050 406.050 ;
        RECT 629.400 400.050 630.600 412.950 ;
        RECT 638.400 403.050 639.600 415.950 ;
        RECT 650.400 415.050 651.600 440.400 ;
        RECT 670.950 439.950 673.050 442.050 ;
        RECT 652.800 436.950 654.900 439.050 ;
        RECT 677.400 438.600 678.600 460.950 ;
        RECT 683.400 454.050 684.600 484.950 ;
        RECT 686.400 457.200 687.600 505.950 ;
        RECT 691.950 502.950 694.050 505.050 ;
        RECT 688.950 496.950 691.050 499.050 ;
        RECT 689.400 463.050 690.600 496.950 ;
        RECT 692.400 463.050 693.600 502.950 ;
        RECT 710.400 496.050 711.600 508.950 ;
        RECT 713.400 505.050 714.600 541.950 ;
        RECT 719.400 529.050 720.600 541.950 ;
        RECT 722.400 541.050 723.600 553.950 ;
        RECT 724.950 544.950 727.050 547.050 ;
        RECT 721.950 538.950 724.050 541.050 ;
        RECT 718.950 526.950 721.050 529.050 ;
        RECT 712.950 502.950 715.050 505.050 ;
        RECT 709.950 493.950 712.050 496.050 ;
        RECT 713.400 490.050 714.600 502.950 ;
        RECT 721.950 493.950 724.050 496.050 ;
        RECT 718.950 490.950 721.050 493.050 ;
        RECT 712.950 487.950 715.050 490.050 ;
        RECT 719.400 487.050 720.600 490.950 ;
        RECT 709.950 484.950 712.050 487.050 ;
        RECT 718.950 484.950 721.050 487.050 ;
        RECT 697.950 478.950 700.050 481.050 ;
        RECT 688.800 460.950 690.900 463.050 ;
        RECT 692.100 460.950 694.200 463.050 ;
        RECT 685.950 455.100 688.050 457.200 ;
        RECT 683.400 453.900 687.000 454.050 ;
        RECT 683.400 452.250 688.050 453.900 ;
        RECT 684.000 451.950 688.050 452.250 ;
        RECT 685.950 451.800 688.050 451.950 ;
        RECT 698.400 445.050 699.600 478.950 ;
        RECT 710.400 472.050 711.600 484.950 ;
        RECT 715.950 481.950 718.050 484.050 ;
        RECT 709.950 469.950 712.050 472.050 ;
        RECT 706.950 460.950 709.050 463.050 ;
        RECT 703.950 451.950 706.050 454.050 ;
        RECT 697.950 442.950 700.050 445.050 ;
        RECT 682.950 439.950 685.050 442.050 ;
        RECT 674.400 437.400 678.600 438.600 ;
        RECT 649.950 412.950 652.050 415.050 ;
        RECT 640.950 406.950 643.050 409.050 ;
        RECT 641.400 403.050 642.600 406.950 ;
        RECT 637.800 400.950 639.900 403.050 ;
        RECT 641.100 400.950 643.200 403.050 ;
        RECT 628.950 397.950 631.050 400.050 ;
        RECT 625.950 388.950 628.050 391.050 ;
        RECT 641.400 390.600 642.600 400.950 ;
        RECT 646.950 397.950 649.050 400.050 ;
        RECT 643.950 394.950 646.050 397.050 ;
        RECT 638.400 389.400 642.600 390.600 ;
        RECT 626.400 382.050 627.600 388.950 ;
        RECT 638.400 385.050 639.600 389.400 ;
        RECT 635.100 382.950 639.600 385.050 ;
        RECT 626.400 380.400 631.050 382.050 ;
        RECT 627.000 379.950 631.050 380.400 ;
        RECT 613.950 370.950 616.050 373.050 ;
        RECT 622.950 370.950 625.050 373.050 ;
        RECT 608.400 362.400 612.600 363.600 ;
        RECT 611.400 349.050 612.600 362.400 ;
        RECT 614.400 355.050 615.600 370.950 ;
        RECT 625.950 364.950 628.050 367.050 ;
        RECT 613.950 352.950 616.050 355.050 ;
        RECT 626.400 354.600 627.600 364.950 ;
        RECT 638.400 364.050 639.600 382.950 ;
        RECT 644.400 382.050 645.600 394.950 ;
        RECT 643.800 381.600 645.900 382.050 ;
        RECT 641.400 380.400 645.900 381.600 ;
        RECT 641.400 376.050 642.600 380.400 ;
        RECT 643.800 379.950 645.900 380.400 ;
        RECT 647.400 379.050 648.600 397.950 ;
        RECT 647.100 376.950 649.200 379.050 ;
        RECT 640.950 373.950 643.050 376.050 ;
        RECT 647.400 367.050 648.600 376.950 ;
        RECT 646.950 364.950 649.050 367.050 ;
        RECT 637.950 361.950 640.050 364.050 ;
        RECT 640.950 358.950 643.050 361.050 ;
        RECT 626.400 353.400 630.600 354.600 ;
        RECT 622.950 349.950 625.050 352.050 ;
        RECT 610.950 346.950 613.050 349.050 ;
        RECT 616.950 343.950 619.050 349.050 ;
        RECT 623.400 343.050 624.600 349.950 ;
        RECT 629.400 349.050 630.600 353.400 ;
        RECT 631.950 349.950 634.050 352.050 ;
        RECT 628.950 346.950 631.050 349.050 ;
        RECT 623.400 341.400 628.050 343.050 ;
        RECT 624.000 340.950 628.050 341.400 ;
        RECT 604.950 334.950 607.050 337.050 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 610.950 331.950 613.050 334.050 ;
        RECT 604.950 328.950 607.050 331.050 ;
        RECT 601.950 322.950 604.050 325.050 ;
        RECT 595.800 316.950 597.900 319.050 ;
        RECT 599.100 316.950 601.200 319.050 ;
        RECT 601.950 313.950 604.050 316.050 ;
        RECT 592.950 310.950 595.050 313.050 ;
        RECT 589.950 306.600 592.050 310.050 ;
        RECT 589.950 306.000 594.600 306.600 ;
        RECT 590.400 305.400 594.600 306.000 ;
        RECT 583.950 284.400 588.600 285.600 ;
        RECT 583.950 283.950 586.050 284.400 ;
        RECT 584.400 277.050 585.600 283.950 ;
        RECT 583.800 274.950 585.900 277.050 ;
        RECT 571.950 271.950 574.050 274.050 ;
        RECT 580.950 271.950 583.050 274.050 ;
        RECT 566.400 269.400 571.200 271.050 ;
        RECT 559.950 265.950 562.050 269.400 ;
        RECT 567.000 268.950 571.200 269.400 ;
        RECT 566.100 265.950 568.200 268.050 ;
        RECT 566.400 256.050 567.600 265.950 ;
        RECT 574.950 262.950 577.050 265.050 ;
        RECT 565.950 253.950 568.050 256.050 ;
        RECT 547.950 250.950 550.050 253.050 ;
        RECT 568.950 250.950 571.050 253.050 ;
        RECT 548.400 235.050 549.600 250.950 ;
        RECT 569.400 244.050 570.600 250.950 ;
        RECT 562.950 241.950 565.050 244.050 ;
        RECT 568.950 241.950 571.050 244.050 ;
        RECT 548.400 233.400 553.050 235.050 ;
        RECT 549.000 232.950 553.050 233.400 ;
        RECT 544.950 211.950 547.050 214.050 ;
        RECT 541.950 202.950 544.050 205.050 ;
        RECT 542.400 175.050 543.600 202.950 ;
        RECT 553.950 195.600 558.000 196.050 ;
        RECT 553.950 193.950 558.600 195.600 ;
        RECT 557.400 184.050 558.600 193.950 ;
        RECT 563.400 193.050 564.600 241.950 ;
        RECT 575.400 238.050 576.600 262.950 ;
        RECT 581.400 246.600 582.600 271.950 ;
        RECT 587.100 270.600 591.000 271.050 ;
        RECT 587.100 268.950 591.600 270.600 ;
        RECT 583.950 265.950 586.050 268.050 ;
        RECT 584.400 250.050 585.600 265.950 ;
        RECT 590.400 262.200 591.600 268.950 ;
        RECT 589.950 260.100 592.050 262.200 ;
        RECT 589.950 256.800 592.050 258.900 ;
        RECT 583.950 247.950 586.050 250.050 ;
        RECT 581.400 245.400 585.600 246.600 ;
        RECT 580.950 241.950 583.050 244.050 ;
        RECT 574.950 235.950 577.050 238.050 ;
        RECT 568.950 220.950 571.050 223.050 ;
        RECT 569.400 199.050 570.600 220.950 ;
        RECT 568.800 196.950 570.900 199.050 ;
        RECT 577.950 193.950 580.050 196.050 ;
        RECT 562.950 190.950 565.050 193.050 ;
        RECT 556.950 181.950 559.050 184.050 ;
        RECT 562.950 178.950 565.050 181.050 ;
        RECT 541.950 172.950 544.050 175.050 ;
        RECT 563.400 169.050 564.600 178.950 ;
        RECT 578.400 169.050 579.600 193.950 ;
        RECT 581.400 171.600 582.600 241.950 ;
        RECT 584.400 205.050 585.600 245.400 ;
        RECT 583.950 202.950 586.050 205.050 ;
        RECT 586.950 196.950 589.050 199.050 ;
        RECT 587.400 187.050 588.600 196.950 ;
        RECT 586.950 184.950 589.050 187.050 ;
        RECT 581.400 170.400 585.600 171.600 ;
        RECT 541.950 166.950 544.050 169.050 ;
        RECT 559.950 167.400 564.600 169.050 ;
        RECT 577.950 168.600 580.050 169.050 ;
        RECT 577.950 167.400 582.600 168.600 ;
        RECT 559.950 166.950 564.000 167.400 ;
        RECT 577.950 166.950 580.050 167.400 ;
        RECT 542.400 151.050 543.600 166.950 ;
        RECT 562.950 163.800 565.050 165.900 ;
        RECT 541.950 148.950 544.050 151.050 ;
        RECT 547.800 148.950 549.900 151.050 ;
        RECT 538.800 124.950 540.900 127.050 ;
        RECT 525.000 123.600 528.900 124.050 ;
        RECT 524.400 121.950 528.900 123.600 ;
        RECT 524.400 112.050 525.600 121.950 ;
        RECT 532.950 115.950 535.050 118.050 ;
        RECT 526.950 112.950 529.050 115.050 ;
        RECT 523.950 109.950 526.050 112.050 ;
        RECT 520.950 97.950 523.050 100.050 ;
        RECT 523.950 94.950 526.050 97.050 ;
        RECT 512.400 92.400 516.900 94.050 ;
        RECT 513.000 91.950 516.900 92.400 ;
        RECT 518.100 91.950 520.200 94.050 ;
        RECT 518.400 61.050 519.600 91.950 ;
        RECT 511.950 58.950 514.050 61.050 ;
        RECT 517.950 58.950 520.050 61.050 ;
        RECT 512.400 55.050 513.600 58.950 ;
        RECT 511.950 52.950 514.050 55.050 ;
        RECT 520.950 54.600 523.050 58.050 ;
        RECT 524.400 54.600 525.600 94.950 ;
        RECT 520.950 54.000 525.600 54.600 ;
        RECT 521.400 53.400 525.600 54.000 ;
        RECT 527.400 52.050 528.600 112.950 ;
        RECT 533.400 100.050 534.600 115.950 ;
        RECT 539.400 103.050 540.600 124.950 ;
        RECT 538.950 100.950 541.050 103.050 ;
        RECT 532.950 97.950 535.050 100.050 ;
        RECT 539.400 97.050 540.600 100.950 ;
        RECT 538.950 94.950 541.050 97.050 ;
        RECT 544.950 91.950 547.050 94.050 ;
        RECT 535.800 90.000 537.900 91.050 ;
        RECT 535.800 88.950 538.050 90.000 ;
        RECT 539.100 88.950 541.200 91.050 ;
        RECT 535.950 85.950 538.050 88.950 ;
        RECT 539.400 52.050 540.600 88.950 ;
        RECT 545.400 70.050 546.600 91.950 ;
        RECT 548.400 91.050 549.600 148.950 ;
        RECT 563.400 148.050 564.600 163.800 ;
        RECT 562.950 145.950 565.050 148.050 ;
        RECT 568.950 142.950 571.050 145.050 ;
        RECT 559.950 136.950 562.050 139.050 ;
        RECT 560.400 100.050 561.600 136.950 ;
        RECT 569.400 124.050 570.600 142.950 ;
        RECT 574.950 139.950 577.050 142.050 ;
        RECT 568.950 121.950 571.050 124.050 ;
        RECT 550.950 97.950 553.050 100.050 ;
        RECT 559.950 97.950 562.050 100.050 ;
        RECT 547.950 88.950 550.050 91.050 ;
        RECT 551.400 88.050 552.600 97.950 ;
        RECT 550.950 85.950 553.050 88.050 ;
        RECT 569.400 73.050 570.600 121.950 ;
        RECT 575.400 106.050 576.600 139.950 ;
        RECT 581.400 130.050 582.600 167.400 ;
        RECT 580.950 127.950 583.050 130.050 ;
        RECT 580.950 112.950 583.050 115.050 ;
        RECT 574.950 103.950 577.050 106.050 ;
        RECT 568.950 70.950 571.050 73.050 ;
        RECT 544.950 67.950 547.050 70.050 ;
        RECT 562.950 67.950 565.050 70.050 ;
        RECT 518.400 51.000 519.600 51.600 ;
        RECT 517.950 46.950 520.050 51.000 ;
        RECT 526.950 49.950 529.050 52.050 ;
        RECT 538.950 49.950 541.050 52.050 ;
        RECT 563.400 49.050 564.600 67.950 ;
        RECT 568.950 55.950 571.050 58.050 ;
        RECT 562.950 46.950 565.050 49.050 ;
        RECT 508.950 28.950 511.050 31.050 ;
        RECT 505.950 19.950 508.050 22.050 ;
        RECT 518.400 7.050 519.600 46.950 ;
        RECT 569.400 22.050 570.600 55.950 ;
        RECT 575.400 55.050 576.600 103.950 ;
        RECT 574.950 52.950 577.050 55.050 ;
        RECT 581.400 22.050 582.600 112.950 ;
        RECT 584.400 70.050 585.600 170.400 ;
        RECT 590.400 165.600 591.600 256.800 ;
        RECT 593.400 253.050 594.600 305.400 ;
        RECT 595.950 301.950 598.050 304.050 ;
        RECT 596.400 255.600 597.600 301.950 ;
        RECT 598.950 295.950 601.050 298.050 ;
        RECT 599.400 259.050 600.600 295.950 ;
        RECT 602.400 292.050 603.600 313.950 ;
        RECT 605.400 310.050 606.600 328.950 ;
        RECT 607.950 322.950 610.050 325.050 ;
        RECT 608.400 316.050 609.600 322.950 ;
        RECT 607.950 313.950 610.050 316.050 ;
        RECT 611.400 310.050 612.600 331.950 ;
        RECT 604.950 307.950 607.050 310.050 ;
        RECT 611.100 307.950 613.200 310.050 ;
        RECT 605.400 301.050 606.600 307.950 ;
        RECT 604.950 298.950 607.050 301.050 ;
        RECT 601.950 289.950 604.050 292.050 ;
        RECT 604.950 280.950 607.050 283.050 ;
        RECT 605.400 268.050 606.600 280.950 ;
        RECT 614.400 277.050 615.600 334.950 ;
        RECT 628.950 331.950 631.050 334.050 ;
        RECT 622.950 325.950 625.050 328.050 ;
        RECT 623.400 322.050 624.600 325.950 ;
        RECT 622.950 319.950 625.050 322.050 ;
        RECT 625.950 310.950 628.050 313.050 ;
        RECT 622.950 304.950 625.050 307.050 ;
        RECT 616.950 292.800 619.050 294.900 ;
        RECT 613.950 274.950 616.050 277.050 ;
        RECT 604.950 265.950 607.050 268.050 ;
        RECT 613.800 267.000 615.900 268.050 ;
        RECT 613.800 265.950 616.050 267.000 ;
        RECT 613.950 262.950 616.050 265.950 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 596.400 254.400 600.600 255.600 ;
        RECT 592.950 250.950 595.050 253.050 ;
        RECT 599.400 246.600 600.600 254.400 ;
        RECT 604.950 253.950 607.050 256.050 ;
        RECT 593.400 245.400 600.600 246.600 ;
        RECT 593.400 208.050 594.600 245.400 ;
        RECT 605.400 244.050 606.600 253.950 ;
        RECT 604.950 241.950 607.050 244.050 ;
        RECT 595.950 240.600 600.000 241.050 ;
        RECT 595.950 238.950 600.600 240.600 ;
        RECT 599.400 217.050 600.600 238.950 ;
        RECT 613.950 229.950 616.050 232.050 ;
        RECT 598.950 214.950 601.050 217.050 ;
        RECT 614.400 214.050 615.600 229.950 ;
        RECT 613.950 211.950 616.050 214.050 ;
        RECT 592.950 205.950 595.050 208.050 ;
        RECT 601.950 205.950 604.050 208.050 ;
        RECT 595.950 202.950 598.050 205.050 ;
        RECT 596.400 196.050 597.600 202.950 ;
        RECT 595.950 193.950 598.050 196.050 ;
        RECT 602.400 192.600 603.600 205.950 ;
        RECT 599.400 191.400 603.600 192.600 ;
        RECT 599.400 180.600 600.600 191.400 ;
        RECT 596.400 179.400 600.600 180.600 ;
        RECT 596.400 169.050 597.600 179.400 ;
        RECT 598.950 169.950 601.050 172.050 ;
        RECT 596.100 166.950 598.200 169.050 ;
        RECT 590.400 164.400 594.600 165.600 ;
        RECT 586.950 133.950 589.050 136.050 ;
        RECT 587.400 127.050 588.600 133.950 ;
        RECT 586.950 124.950 589.050 127.050 ;
        RECT 593.400 124.050 594.600 164.400 ;
        RECT 595.950 160.950 598.050 163.050 ;
        RECT 596.400 126.600 597.600 160.950 ;
        RECT 599.400 133.050 600.600 169.950 ;
        RECT 612.000 168.600 616.050 169.050 ;
        RECT 611.400 166.950 616.050 168.600 ;
        RECT 611.400 163.050 612.600 166.950 ;
        RECT 617.400 166.050 618.600 292.800 ;
        RECT 623.400 283.050 624.600 304.950 ;
        RECT 626.400 301.200 627.600 310.950 ;
        RECT 629.400 307.050 630.600 331.950 ;
        RECT 628.950 304.950 631.050 307.050 ;
        RECT 625.950 299.100 628.050 301.200 ;
        RECT 622.950 280.950 625.050 283.050 ;
        RECT 619.950 271.950 622.050 274.050 ;
        RECT 620.400 268.050 621.600 271.950 ;
        RECT 628.950 268.950 631.050 271.050 ;
        RECT 620.100 267.600 622.200 268.050 ;
        RECT 620.100 266.400 624.600 267.600 ;
        RECT 620.100 265.950 622.200 266.400 ;
        RECT 619.950 256.950 622.050 259.050 ;
        RECT 620.400 238.050 621.600 256.950 ;
        RECT 619.950 235.950 622.050 238.050 ;
        RECT 623.400 232.050 624.600 266.400 ;
        RECT 629.400 241.050 630.600 268.950 ;
        RECT 632.400 247.200 633.600 349.950 ;
        RECT 634.950 346.950 637.050 349.050 ;
        RECT 635.400 274.050 636.600 346.950 ;
        RECT 637.800 337.950 639.900 340.050 ;
        RECT 638.400 313.050 639.600 337.950 ;
        RECT 637.950 310.950 640.050 313.050 ;
        RECT 637.950 301.950 640.050 304.050 ;
        RECT 634.950 271.950 637.050 274.050 ;
        RECT 634.800 267.000 636.900 268.050 ;
        RECT 634.800 265.950 637.050 267.000 ;
        RECT 634.950 262.950 637.050 265.950 ;
        RECT 631.950 245.100 634.050 247.200 ;
        RECT 638.400 244.050 639.600 301.950 ;
        RECT 641.400 295.050 642.600 358.950 ;
        RECT 643.950 355.950 646.050 358.050 ;
        RECT 644.400 322.050 645.600 355.950 ;
        RECT 653.400 352.050 654.600 436.950 ;
        RECT 670.950 433.950 673.050 436.050 ;
        RECT 655.950 430.950 658.050 433.050 ;
        RECT 661.950 430.950 664.050 433.050 ;
        RECT 656.400 358.050 657.600 430.950 ;
        RECT 662.400 411.600 663.600 430.950 ;
        RECT 667.950 418.950 670.050 421.050 ;
        RECT 659.400 410.400 663.600 411.600 ;
        RECT 659.400 394.050 660.600 410.400 ;
        RECT 661.950 406.950 664.050 409.050 ;
        RECT 658.950 391.950 661.050 394.050 ;
        RECT 662.400 388.050 663.600 406.950 ;
        RECT 668.400 388.200 669.600 418.950 ;
        RECT 661.950 385.950 664.050 388.050 ;
        RECT 667.950 386.100 670.050 388.200 ;
        RECT 667.950 384.600 670.050 384.900 ;
        RECT 671.400 384.600 672.600 433.950 ;
        RECT 667.950 383.400 672.600 384.600 ;
        RECT 667.950 382.800 670.050 383.400 ;
        RECT 661.950 379.950 664.050 382.050 ;
        RECT 662.400 376.050 663.600 379.950 ;
        RECT 661.950 373.950 664.050 376.050 ;
        RECT 655.950 355.950 658.050 358.050 ;
        RECT 661.950 352.950 664.050 355.050 ;
        RECT 652.950 349.950 655.050 352.050 ;
        RECT 662.400 349.050 663.600 352.950 ;
        RECT 664.950 349.950 667.050 352.050 ;
        RECT 661.950 346.950 664.050 349.050 ;
        RECT 646.950 343.950 649.050 346.050 ;
        RECT 652.950 343.950 655.050 346.050 ;
        RECT 647.400 340.050 648.600 343.950 ;
        RECT 646.950 337.950 649.050 340.050 ;
        RECT 643.950 319.950 646.050 322.050 ;
        RECT 646.950 312.600 651.000 313.050 ;
        RECT 646.950 310.950 651.600 312.600 ;
        RECT 650.400 304.050 651.600 310.950 ;
        RECT 653.400 310.050 654.600 343.950 ;
        RECT 662.400 313.050 663.600 346.950 ;
        RECT 665.400 319.200 666.600 349.950 ;
        RECT 668.400 325.200 669.600 382.800 ;
        RECT 670.950 373.950 673.050 376.050 ;
        RECT 667.950 323.100 670.050 325.200 ;
        RECT 667.950 319.800 670.050 321.900 ;
        RECT 664.950 317.100 667.050 319.200 ;
        RECT 664.950 313.800 667.050 315.900 ;
        RECT 661.950 310.950 664.050 313.050 ;
        RECT 652.950 307.950 655.050 310.050 ;
        RECT 655.950 304.950 658.050 307.050 ;
        RECT 649.950 301.950 652.050 304.050 ;
        RECT 646.950 298.950 649.050 301.050 ;
        RECT 643.950 295.950 646.050 298.050 ;
        RECT 640.950 292.950 643.050 295.050 ;
        RECT 640.950 274.950 643.050 277.050 ;
        RECT 631.950 241.800 634.050 243.900 ;
        RECT 637.950 241.950 640.050 244.050 ;
        RECT 628.950 238.950 631.050 241.050 ;
        RECT 632.400 238.050 633.600 241.800 ;
        RECT 632.100 235.950 634.200 238.050 ;
        RECT 622.950 229.950 625.050 232.050 ;
        RECT 631.950 229.950 634.050 232.050 ;
        RECT 622.950 223.950 625.050 226.050 ;
        RECT 619.950 208.950 622.050 211.050 ;
        RECT 620.400 202.050 621.600 208.950 ;
        RECT 619.950 199.950 622.050 202.050 ;
        RECT 620.400 196.050 621.600 199.950 ;
        RECT 619.950 193.950 622.050 196.050 ;
        RECT 617.400 164.400 622.050 166.050 ;
        RECT 618.000 163.950 622.050 164.400 ;
        RECT 610.950 160.950 613.050 163.050 ;
        RECT 623.400 148.050 624.600 223.950 ;
        RECT 632.400 199.050 633.600 229.950 ;
        RECT 641.400 226.050 642.600 274.950 ;
        RECT 640.950 223.950 643.050 226.050 ;
        RECT 640.950 214.950 643.050 217.050 ;
        RECT 641.400 205.050 642.600 214.950 ;
        RECT 640.950 202.950 643.050 205.050 ;
        RECT 634.950 199.950 637.050 202.050 ;
        RECT 631.950 196.950 634.050 199.050 ;
        RECT 631.950 181.950 634.050 184.050 ;
        RECT 632.400 166.050 633.600 181.950 ;
        RECT 631.950 163.950 634.050 166.050 ;
        RECT 635.400 163.050 636.600 199.950 ;
        RECT 641.400 196.050 642.600 202.950 ;
        RECT 640.950 193.950 643.050 196.050 ;
        RECT 644.400 175.050 645.600 295.950 ;
        RECT 647.400 246.600 648.600 298.950 ;
        RECT 651.000 270.600 655.050 271.050 ;
        RECT 650.400 268.950 655.050 270.600 ;
        RECT 650.400 250.050 651.600 268.950 ;
        RECT 656.400 268.050 657.600 304.950 ;
        RECT 665.400 298.050 666.600 313.800 ;
        RECT 664.950 295.950 667.050 298.050 ;
        RECT 658.950 292.950 661.050 295.050 ;
        RECT 659.400 270.600 660.600 292.950 ;
        RECT 661.950 289.950 664.050 292.050 ;
        RECT 662.400 283.050 663.600 289.950 ;
        RECT 661.950 280.950 664.050 283.050 ;
        RECT 661.950 270.600 664.050 271.050 ;
        RECT 659.400 269.400 664.050 270.600 ;
        RECT 661.950 268.950 664.050 269.400 ;
        RECT 655.950 265.950 658.050 268.050 ;
        RECT 652.950 262.950 655.050 265.050 ;
        RECT 649.950 247.950 652.050 250.050 ;
        RECT 647.400 245.400 651.600 246.600 ;
        RECT 646.950 241.950 649.050 244.050 ;
        RECT 647.400 238.050 648.600 241.950 ;
        RECT 647.100 235.950 649.200 238.050 ;
        RECT 650.400 235.050 651.600 245.400 ;
        RECT 650.100 232.950 652.200 235.050 ;
        RECT 646.950 220.950 649.050 223.050 ;
        RECT 647.400 193.050 648.600 220.950 ;
        RECT 650.400 217.050 651.600 232.950 ;
        RECT 653.400 220.050 654.600 262.950 ;
        RECT 656.400 256.050 657.600 265.950 ;
        RECT 655.950 253.950 658.050 256.050 ;
        RECT 658.950 241.950 661.050 244.050 ;
        RECT 659.400 223.050 660.600 241.950 ;
        RECT 658.950 220.950 661.050 223.050 ;
        RECT 652.950 217.950 655.050 220.050 ;
        RECT 649.950 214.950 652.050 217.050 ;
        RECT 655.950 211.950 658.050 214.050 ;
        RECT 656.400 202.050 657.600 211.950 ;
        RECT 652.950 200.400 657.600 202.050 ;
        RECT 652.950 199.950 657.000 200.400 ;
        RECT 646.950 190.950 649.050 193.050 ;
        RECT 643.950 172.950 646.050 175.050 ;
        RECT 653.400 172.050 654.600 199.950 ;
        RECT 662.400 196.050 663.600 268.950 ;
        RECT 664.950 265.950 667.050 268.050 ;
        RECT 665.400 226.050 666.600 265.950 ;
        RECT 668.400 244.050 669.600 319.800 ;
        RECT 671.400 313.050 672.600 373.950 ;
        RECT 674.400 373.050 675.600 437.400 ;
        RECT 676.950 433.950 679.050 436.050 ;
        RECT 677.400 421.050 678.600 433.950 ;
        RECT 676.950 418.950 679.050 421.050 ;
        RECT 679.950 409.950 682.050 412.050 ;
        RECT 673.950 370.950 676.050 373.050 ;
        RECT 676.950 364.950 679.050 367.050 ;
        RECT 677.400 346.050 678.600 364.950 ;
        RECT 680.400 361.050 681.600 409.950 ;
        RECT 683.400 376.050 684.600 439.950 ;
        RECT 697.950 427.950 700.050 430.050 ;
        RECT 698.400 415.050 699.600 427.950 ;
        RECT 700.950 418.950 703.050 421.050 ;
        RECT 695.100 413.400 699.600 415.050 ;
        RECT 695.100 412.950 699.000 413.400 ;
        RECT 691.800 409.950 693.900 412.050 ;
        RECT 692.400 405.600 693.600 409.950 ;
        RECT 689.400 405.000 693.600 405.600 ;
        RECT 688.950 404.400 693.600 405.000 ;
        RECT 688.950 400.950 691.050 404.400 ;
        RECT 695.400 403.050 696.600 412.950 ;
        RECT 701.400 412.050 702.600 418.950 ;
        RECT 700.950 409.950 703.050 412.050 ;
        RECT 694.950 400.950 697.050 403.050 ;
        RECT 704.400 400.050 705.600 451.950 ;
        RECT 703.950 397.950 706.050 400.050 ;
        RECT 688.950 391.950 691.050 394.050 ;
        RECT 685.950 388.950 688.050 391.050 ;
        RECT 686.400 382.050 687.600 388.950 ;
        RECT 685.950 379.950 688.050 382.050 ;
        RECT 682.950 373.950 685.050 376.050 ;
        RECT 679.950 358.950 682.050 361.050 ;
        RECT 682.950 349.950 685.050 352.050 ;
        RECT 683.400 346.050 684.600 349.950 ;
        RECT 676.950 342.600 679.050 346.050 ;
        RECT 682.950 343.950 685.050 346.050 ;
        RECT 674.400 342.000 679.050 342.600 ;
        RECT 674.400 341.400 678.600 342.000 ;
        RECT 674.400 331.050 675.600 341.400 ;
        RECT 678.000 339.900 681.000 340.050 ;
        RECT 677.100 339.600 681.000 339.900 ;
        RECT 677.100 337.950 681.600 339.600 ;
        RECT 677.100 337.800 679.200 337.950 ;
        RECT 673.950 328.950 676.050 331.050 ;
        RECT 673.950 316.950 676.050 319.050 ;
        RECT 670.950 310.950 673.050 313.050 ;
        RECT 674.400 310.050 675.600 316.950 ;
        RECT 680.400 310.050 681.600 337.950 ;
        RECT 685.950 334.950 688.050 337.050 ;
        RECT 686.400 319.050 687.600 334.950 ;
        RECT 685.950 316.950 688.050 319.050 ;
        RECT 682.950 312.600 687.000 313.050 ;
        RECT 682.950 310.950 687.600 312.600 ;
        RECT 673.950 307.950 676.050 310.050 ;
        RECT 679.950 307.950 682.050 310.050 ;
        RECT 670.950 298.950 673.050 301.050 ;
        RECT 671.400 268.050 672.600 298.950 ;
        RECT 674.400 274.050 675.600 307.950 ;
        RECT 686.400 304.050 687.600 310.950 ;
        RECT 685.950 301.950 688.050 304.050 ;
        RECT 689.400 301.050 690.600 391.950 ;
        RECT 703.950 382.950 706.050 385.050 ;
        RECT 704.400 379.050 705.600 382.950 ;
        RECT 691.950 376.950 694.050 379.050 ;
        RECT 703.950 376.950 706.050 379.050 ;
        RECT 692.400 355.050 693.600 376.950 ;
        RECT 707.400 376.050 708.600 460.950 ;
        RECT 716.400 460.050 717.600 481.950 ;
        RECT 718.950 475.950 721.050 478.050 ;
        RECT 715.950 456.000 718.050 460.050 ;
        RECT 716.400 455.400 717.600 456.000 ;
        RECT 716.100 451.800 718.200 453.900 ;
        RECT 712.800 448.950 714.900 451.050 ;
        RECT 713.400 445.200 714.600 448.950 ;
        RECT 716.400 448.050 717.600 451.800 ;
        RECT 715.950 445.950 718.050 448.050 ;
        RECT 712.950 443.100 715.050 445.200 ;
        RECT 712.950 439.800 715.050 441.900 ;
        RECT 709.950 427.950 712.050 430.050 ;
        RECT 710.400 412.050 711.600 427.950 ;
        RECT 709.950 409.950 712.050 412.050 ;
        RECT 709.950 403.950 712.050 406.050 ;
        RECT 710.400 385.050 711.600 403.950 ;
        RECT 713.400 400.050 714.600 439.800 ;
        RECT 719.400 436.050 720.600 475.950 ;
        RECT 718.950 433.950 721.050 436.050 ;
        RECT 722.400 424.050 723.600 493.950 ;
        RECT 721.950 421.950 724.050 424.050 ;
        RECT 720.000 414.600 724.050 415.050 ;
        RECT 719.400 412.950 724.050 414.600 ;
        RECT 719.400 409.050 720.600 412.950 ;
        RECT 718.950 408.600 721.050 409.050 ;
        RECT 716.400 407.400 721.050 408.600 ;
        RECT 712.950 397.950 715.050 400.050 ;
        RECT 709.950 382.950 712.050 385.050 ;
        RECT 716.400 382.050 717.600 407.400 ;
        RECT 718.950 406.950 721.050 407.400 ;
        RECT 718.950 400.950 721.050 403.050 ;
        RECT 719.400 388.050 720.600 400.950 ;
        RECT 719.400 386.400 724.050 388.050 ;
        RECT 720.000 385.950 724.050 386.400 ;
        RECT 715.950 379.950 718.050 382.050 ;
        RECT 706.950 373.950 709.050 376.050 ;
        RECT 712.950 373.950 715.050 376.050 ;
        RECT 694.950 370.950 697.050 373.050 ;
        RECT 709.950 370.950 712.050 373.050 ;
        RECT 691.950 352.950 694.050 355.050 ;
        RECT 691.950 343.950 694.050 346.050 ;
        RECT 692.400 322.050 693.600 343.950 ;
        RECT 691.950 319.950 694.050 322.050 ;
        RECT 688.950 298.950 691.050 301.050 ;
        RECT 679.950 295.950 682.050 298.050 ;
        RECT 673.950 271.950 676.050 274.050 ;
        RECT 676.950 268.950 679.050 271.050 ;
        RECT 670.800 265.950 672.900 268.050 ;
        RECT 674.100 265.950 676.200 268.050 ;
        RECT 674.400 253.050 675.600 265.950 ;
        RECT 677.400 262.050 678.600 268.950 ;
        RECT 676.950 259.950 679.050 262.050 ;
        RECT 680.400 259.050 681.600 295.950 ;
        RECT 682.950 286.950 685.050 289.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 673.950 250.950 676.050 253.050 ;
        RECT 679.950 247.950 682.050 250.050 ;
        RECT 680.400 244.050 681.600 247.950 ;
        RECT 667.950 241.950 670.050 244.050 ;
        RECT 679.950 241.950 682.050 244.050 ;
        RECT 667.950 235.950 670.050 238.050 ;
        RECT 664.950 223.950 667.050 226.050 ;
        RECT 668.400 202.050 669.600 235.950 ;
        RECT 670.950 232.950 673.050 235.050 ;
        RECT 671.400 211.050 672.600 232.950 ;
        RECT 673.950 229.950 676.050 232.050 ;
        RECT 670.950 208.950 673.050 211.050 ;
        RECT 667.950 199.950 670.050 202.050 ;
        RECT 670.950 196.950 673.050 199.050 ;
        RECT 661.950 193.950 664.050 196.050 ;
        RECT 655.950 190.950 658.050 193.050 ;
        RECT 652.950 169.950 655.050 172.050 ;
        RECT 649.950 163.950 652.050 166.050 ;
        RECT 628.950 160.950 631.050 163.050 ;
        RECT 634.950 160.950 637.050 163.050 ;
        RECT 641.100 162.000 643.200 163.050 ;
        RECT 640.950 160.950 643.200 162.000 ;
        RECT 646.950 160.950 649.050 163.050 ;
        RECT 625.950 154.950 628.050 157.050 ;
        RECT 610.950 145.950 613.050 148.050 ;
        RECT 622.950 145.950 625.050 148.050 ;
        RECT 604.950 142.950 607.050 145.050 ;
        RECT 605.400 133.050 606.600 142.950 ;
        RECT 598.950 130.950 601.050 133.050 ;
        RECT 604.950 130.950 607.050 133.050 ;
        RECT 596.400 125.400 600.600 126.600 ;
        RECT 592.950 121.950 595.050 124.050 ;
        RECT 593.400 112.050 594.600 121.950 ;
        RECT 592.950 109.950 595.050 112.050 ;
        RECT 599.400 109.050 600.600 125.400 ;
        RECT 607.950 124.950 610.050 127.050 ;
        RECT 604.950 118.950 607.050 121.050 ;
        RECT 589.950 106.950 592.050 109.050 ;
        RECT 598.950 106.950 601.050 109.050 ;
        RECT 583.950 67.950 586.050 70.050 ;
        RECT 590.400 25.050 591.600 106.950 ;
        RECT 595.950 100.950 598.050 103.050 ;
        RECT 592.950 97.950 595.050 100.050 ;
        RECT 593.400 94.050 594.600 97.950 ;
        RECT 596.400 97.050 597.600 100.950 ;
        RECT 596.400 95.400 601.050 97.050 ;
        RECT 597.000 94.950 601.050 95.400 ;
        RECT 592.950 91.950 595.050 94.050 ;
        RECT 601.950 82.950 604.050 85.050 ;
        RECT 602.400 58.050 603.600 82.950 ;
        RECT 601.950 55.950 604.050 58.050 ;
        RECT 592.950 49.950 595.050 52.050 ;
        RECT 589.800 22.950 591.900 25.050 ;
        RECT 593.400 22.050 594.600 49.950 ;
        RECT 605.400 49.050 606.600 118.950 ;
        RECT 608.400 94.050 609.600 124.950 ;
        RECT 607.950 91.950 610.050 94.050 ;
        RECT 604.950 46.950 607.050 49.050 ;
        RECT 568.800 19.950 570.900 22.050 ;
        RECT 580.950 19.950 583.050 22.050 ;
        RECT 592.950 19.950 595.050 22.050 ;
        RECT 541.950 18.600 546.000 19.050 ;
        RECT 541.950 16.950 546.600 18.600 ;
        RECT 565.800 18.000 567.900 19.050 ;
        RECT 565.800 16.950 568.050 18.000 ;
        RECT 526.950 10.950 529.050 16.050 ;
        RECT 545.400 13.200 546.600 16.950 ;
        RECT 565.950 13.950 568.050 16.950 ;
        RECT 544.950 11.100 547.050 13.200 ;
        RECT 611.400 7.050 612.600 145.950 ;
        RECT 616.950 139.950 619.050 142.050 ;
        RECT 613.950 136.950 616.050 139.050 ;
        RECT 614.400 25.050 615.600 136.950 ;
        RECT 617.400 133.050 618.600 139.950 ;
        RECT 626.400 139.050 627.600 154.950 ;
        RECT 625.950 136.950 628.050 139.050 ;
        RECT 616.950 130.950 619.050 133.050 ;
        RECT 624.000 129.600 628.050 130.050 ;
        RECT 623.400 127.950 628.050 129.600 ;
        RECT 623.400 121.050 624.600 127.950 ;
        RECT 629.400 127.050 630.600 160.950 ;
        RECT 635.400 157.050 636.600 160.950 ;
        RECT 640.950 157.950 643.050 160.950 ;
        RECT 647.400 157.050 648.600 160.950 ;
        RECT 634.950 154.950 637.050 157.050 ;
        RECT 646.950 154.950 649.050 157.050 ;
        RECT 646.950 145.950 649.050 148.050 ;
        RECT 634.950 130.950 637.050 133.050 ;
        RECT 635.400 127.050 636.600 130.950 ;
        RECT 628.950 124.950 631.050 127.050 ;
        RECT 634.800 124.950 636.900 127.050 ;
        RECT 642.000 123.600 646.050 124.050 ;
        RECT 641.400 121.950 646.050 123.600 ;
        RECT 622.950 118.950 625.050 121.050 ;
        RECT 641.400 106.050 642.600 121.950 ;
        RECT 625.950 103.950 628.050 106.050 ;
        RECT 640.950 103.950 643.050 106.050 ;
        RECT 626.400 97.050 627.600 103.950 ;
        RECT 641.400 100.050 642.600 103.950 ;
        RECT 647.400 103.200 648.600 145.950 ;
        RECT 650.400 145.050 651.600 163.950 ;
        RECT 656.400 148.050 657.600 190.950 ;
        RECT 671.400 157.050 672.600 196.950 ;
        RECT 670.950 154.950 673.050 157.050 ;
        RECT 674.400 151.050 675.600 229.950 ;
        RECT 683.400 193.050 684.600 286.950 ;
        RECT 695.400 280.050 696.600 370.950 ;
        RECT 700.950 364.950 703.050 367.050 ;
        RECT 701.400 352.050 702.600 364.950 ;
        RECT 706.950 361.950 709.050 364.050 ;
        RECT 703.950 358.950 706.050 361.050 ;
        RECT 700.950 349.950 703.050 352.050 ;
        RECT 700.800 343.050 702.900 343.200 ;
        RECT 699.000 342.600 702.900 343.050 ;
        RECT 698.400 341.100 702.900 342.600 ;
        RECT 698.400 340.950 702.000 341.100 ;
        RECT 698.400 334.050 699.600 340.950 ;
        RECT 704.400 339.600 705.600 358.950 ;
        RECT 707.400 352.050 708.600 361.950 ;
        RECT 706.950 349.950 709.050 352.050 ;
        RECT 707.400 346.050 708.600 349.950 ;
        RECT 706.950 343.950 709.050 346.050 ;
        RECT 701.400 339.000 705.600 339.600 ;
        RECT 700.950 338.400 705.600 339.000 ;
        RECT 700.950 334.950 703.050 338.400 ;
        RECT 697.950 331.950 700.050 334.050 ;
        RECT 698.400 322.050 699.600 331.950 ;
        RECT 697.950 319.950 700.050 322.050 ;
        RECT 707.400 319.050 708.600 343.950 ;
        RECT 706.950 316.950 709.050 319.050 ;
        RECT 706.950 310.950 709.050 313.050 ;
        RECT 710.400 312.600 711.600 370.950 ;
        RECT 713.400 316.050 714.600 373.950 ;
        RECT 715.950 361.950 718.050 364.050 ;
        RECT 712.950 313.950 715.050 316.050 ;
        RECT 710.400 311.400 714.600 312.600 ;
        RECT 697.950 301.950 700.050 304.050 ;
        RECT 694.950 277.950 697.050 280.050 ;
        RECT 685.950 274.950 688.050 277.050 ;
        RECT 678.000 192.600 681.900 193.050 ;
        RECT 677.400 190.950 681.900 192.600 ;
        RECT 683.100 190.950 685.200 193.050 ;
        RECT 673.950 148.950 676.050 151.050 ;
        RECT 655.950 145.950 658.050 148.050 ;
        RECT 649.950 142.950 652.050 145.050 ;
        RECT 661.950 142.950 664.050 145.050 ;
        RECT 655.950 139.950 658.050 142.050 ;
        RECT 652.950 124.950 655.050 127.050 ;
        RECT 653.400 121.050 654.600 124.950 ;
        RECT 652.950 118.950 655.050 121.050 ;
        RECT 656.400 109.050 657.600 139.950 ;
        RECT 658.950 124.950 661.050 127.050 ;
        RECT 655.950 106.950 658.050 109.050 ;
        RECT 646.950 101.100 649.050 103.200 ;
        RECT 640.800 97.950 642.900 100.050 ;
        RECT 646.950 97.800 649.050 99.900 ;
        RECT 622.950 94.950 627.600 97.050 ;
        RECT 626.400 67.050 627.600 94.950 ;
        RECT 631.950 91.950 634.050 94.050 ;
        RECT 625.950 64.950 628.050 67.050 ;
        RECT 632.400 61.050 633.600 91.950 ;
        RECT 647.400 91.050 648.600 97.800 ;
        RECT 659.400 97.050 660.600 124.950 ;
        RECT 662.400 121.050 663.600 142.950 ;
        RECT 677.400 139.050 678.600 190.950 ;
        RECT 686.400 190.200 687.600 274.950 ;
        RECT 688.950 271.950 691.050 274.050 ;
        RECT 689.400 268.050 690.600 271.950 ;
        RECT 689.400 266.400 694.050 268.050 ;
        RECT 690.000 265.950 694.050 266.400 ;
        RECT 694.950 262.950 697.050 265.050 ;
        RECT 688.950 256.950 691.050 259.050 ;
        RECT 689.400 217.200 690.600 256.950 ;
        RECT 691.950 253.950 694.050 256.050 ;
        RECT 688.950 215.100 691.050 217.200 ;
        RECT 688.950 213.600 691.050 213.900 ;
        RECT 692.400 213.600 693.600 253.950 ;
        RECT 695.400 253.200 696.600 262.950 ;
        RECT 694.950 251.100 697.050 253.200 ;
        RECT 694.800 247.800 696.900 249.900 ;
        RECT 695.400 238.050 696.600 247.800 ;
        RECT 694.950 235.950 697.050 238.050 ;
        RECT 698.400 220.050 699.600 301.950 ;
        RECT 700.950 298.950 703.050 301.050 ;
        RECT 701.400 283.050 702.600 298.950 ;
        RECT 700.950 280.950 703.050 283.050 ;
        RECT 703.950 277.950 706.050 280.050 ;
        RECT 701.100 268.950 703.200 271.050 ;
        RECT 701.400 265.050 702.600 268.950 ;
        RECT 700.950 262.950 703.050 265.050 ;
        RECT 704.400 255.600 705.600 277.950 ;
        RECT 707.400 259.200 708.600 310.950 ;
        RECT 709.950 265.950 712.050 268.050 ;
        RECT 706.950 257.100 709.050 259.200 ;
        RECT 701.400 254.400 705.600 255.600 ;
        RECT 701.400 235.050 702.600 254.400 ;
        RECT 706.950 253.800 709.050 255.900 ;
        RECT 707.400 250.050 708.600 253.800 ;
        RECT 706.950 247.950 709.050 250.050 ;
        RECT 710.400 235.050 711.600 265.950 ;
        RECT 700.950 232.950 703.050 235.050 ;
        RECT 709.950 232.950 712.050 235.050 ;
        RECT 700.950 223.950 703.050 226.050 ;
        RECT 697.950 217.950 700.050 220.050 ;
        RECT 688.950 212.400 693.600 213.600 ;
        RECT 688.950 211.800 691.050 212.400 ;
        RECT 689.400 196.050 690.600 211.800 ;
        RECT 694.950 205.950 697.050 208.050 ;
        RECT 695.400 202.050 696.600 205.950 ;
        RECT 694.950 199.950 697.050 202.050 ;
        RECT 688.950 193.950 691.050 196.050 ;
        RECT 695.100 195.600 699.000 196.050 ;
        RECT 695.100 193.950 699.600 195.600 ;
        RECT 698.400 193.050 699.600 193.950 ;
        RECT 691.950 190.950 694.050 193.050 ;
        RECT 697.950 190.950 700.050 193.050 ;
        RECT 685.950 188.100 688.050 190.200 ;
        RECT 685.950 184.800 688.050 186.900 ;
        RECT 679.950 172.950 682.050 175.050 ;
        RECT 676.950 136.950 679.050 139.050 ;
        RECT 667.950 124.950 670.050 127.050 ;
        RECT 674.100 126.600 678.000 127.050 ;
        RECT 674.100 124.950 678.600 126.600 ;
        RECT 661.800 118.950 663.900 121.050 ;
        RECT 668.400 118.050 669.600 124.950 ;
        RECT 667.950 115.950 670.050 118.050 ;
        RECT 664.950 109.950 667.050 112.050 ;
        RECT 670.950 109.950 673.050 112.050 ;
        RECT 665.400 100.050 666.600 109.950 ;
        RECT 665.100 97.950 667.200 100.050 ;
        RECT 659.400 95.400 663.900 97.050 ;
        RECT 660.000 94.950 663.900 95.400 ;
        RECT 646.950 88.950 649.050 91.050 ;
        RECT 671.400 70.050 672.600 109.950 ;
        RECT 677.400 106.050 678.600 124.950 ;
        RECT 680.400 112.050 681.600 172.950 ;
        RECT 686.400 166.050 687.600 184.800 ;
        RECT 692.400 184.050 693.600 190.950 ;
        RECT 691.950 181.950 694.050 184.050 ;
        RECT 698.400 172.050 699.600 190.950 ;
        RECT 701.400 178.050 702.600 223.950 ;
        RECT 706.950 220.950 709.050 223.050 ;
        RECT 703.950 214.950 706.050 217.050 ;
        RECT 700.950 175.950 703.050 178.050 ;
        RECT 688.950 169.950 691.050 172.050 ;
        RECT 697.950 169.950 700.050 172.050 ;
        RECT 682.950 164.400 687.600 166.050 ;
        RECT 682.950 163.950 687.000 164.400 ;
        RECT 689.400 163.050 690.600 169.950 ;
        RECT 695.100 163.950 697.200 166.050 ;
        RECT 688.950 160.950 691.050 163.050 ;
        RECT 695.400 121.050 696.600 163.950 ;
        RECT 704.400 163.050 705.600 214.950 ;
        RECT 707.400 199.050 708.600 220.950 ;
        RECT 706.950 196.950 709.050 199.050 ;
        RECT 713.400 187.050 714.600 311.400 ;
        RECT 716.400 289.050 717.600 361.950 ;
        RECT 725.400 355.050 726.600 544.950 ;
        RECT 728.400 496.050 729.600 583.950 ;
        RECT 732.000 552.600 736.050 553.050 ;
        RECT 731.400 550.950 736.050 552.600 ;
        RECT 731.400 505.050 732.600 550.950 ;
        RECT 737.400 547.050 738.600 607.950 ;
        RECT 752.400 595.050 753.600 625.950 ;
        RECT 755.400 613.050 756.600 625.950 ;
        RECT 754.950 610.950 757.050 613.050 ;
        RECT 739.950 592.950 742.050 595.050 ;
        RECT 751.800 592.950 753.900 595.050 ;
        RECT 740.400 552.600 741.600 592.950 ;
        RECT 745.950 574.950 748.050 577.050 ;
        RECT 746.400 565.050 747.600 574.950 ;
        RECT 745.950 562.950 748.050 565.050 ;
        RECT 746.400 559.200 747.600 562.950 ;
        RECT 745.950 557.100 748.050 559.200 ;
        RECT 742.950 555.600 747.000 556.050 ;
        RECT 742.950 553.950 747.600 555.600 ;
        RECT 749.100 553.950 751.200 556.050 ;
        RECT 740.400 551.400 744.600 552.600 ;
        RECT 736.950 544.950 739.050 547.050 ;
        RECT 737.400 529.050 738.600 544.950 ;
        RECT 739.950 541.950 742.050 544.050 ;
        RECT 740.400 532.050 741.600 541.950 ;
        RECT 739.950 529.950 742.050 532.050 ;
        RECT 733.950 527.400 738.600 529.050 ;
        RECT 733.950 526.950 738.000 527.400 ;
        RECT 730.950 502.950 733.050 505.050 ;
        RECT 739.950 502.950 742.050 505.050 ;
        RECT 740.400 499.050 741.600 502.950 ;
        RECT 739.950 496.950 742.050 499.050 ;
        RECT 727.950 493.950 730.050 496.050 ;
        RECT 740.400 487.050 741.600 496.950 ;
        RECT 739.950 484.950 742.050 487.050 ;
        RECT 727.950 472.950 730.050 475.050 ;
        RECT 728.400 451.050 729.600 472.950 ;
        RECT 730.950 463.950 733.050 466.050 ;
        RECT 731.400 454.050 732.600 463.950 ;
        RECT 730.800 451.950 732.900 454.050 ;
        RECT 727.800 448.950 729.900 451.050 ;
        RECT 739.950 448.950 742.050 451.050 ;
        RECT 736.950 436.800 739.050 438.900 ;
        RECT 737.400 427.050 738.600 436.800 ;
        RECT 740.400 430.050 741.600 448.950 ;
        RECT 743.400 439.050 744.600 551.400 ;
        RECT 746.400 511.050 747.600 553.950 ;
        RECT 749.400 541.050 750.600 553.950 ;
        RECT 755.400 550.050 756.600 610.950 ;
        RECT 754.950 547.950 757.050 550.050 ;
        RECT 758.400 541.050 759.600 676.950 ;
        RECT 761.400 670.050 762.600 703.950 ;
        RECT 763.950 694.950 766.050 697.050 ;
        RECT 761.100 667.950 763.200 670.050 ;
        RECT 760.950 649.950 763.050 652.050 ;
        RECT 748.950 538.950 751.050 541.050 ;
        RECT 757.950 538.950 760.050 541.050 ;
        RECT 761.400 538.050 762.600 649.950 ;
        RECT 764.400 580.050 765.600 694.950 ;
        RECT 767.400 685.050 768.600 826.950 ;
        RECT 769.950 820.950 772.050 823.050 ;
        RECT 770.400 808.050 771.600 820.950 ;
        RECT 773.400 817.050 774.600 844.950 ;
        RECT 785.400 826.050 786.600 844.950 ;
        RECT 791.100 841.950 793.200 844.050 ;
        RECT 809.100 841.950 811.200 844.050 ;
        RECT 784.950 823.950 787.050 826.050 ;
        RECT 787.950 820.050 790.050 823.050 ;
        RECT 781.950 817.950 784.050 820.050 ;
        RECT 787.950 819.000 790.200 820.050 ;
        RECT 788.100 817.950 790.200 819.000 ;
        RECT 773.400 815.400 778.050 817.050 ;
        RECT 774.000 814.950 778.050 815.400 ;
        RECT 769.950 805.950 772.050 808.050 ;
        RECT 782.400 805.050 783.600 817.950 ;
        RECT 787.950 811.950 790.050 814.050 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 788.400 769.050 789.600 811.950 ;
        RECT 787.950 766.950 790.050 769.050 ;
        RECT 791.400 765.600 792.600 841.950 ;
        RECT 805.800 838.950 807.900 841.050 ;
        RECT 802.950 829.950 805.050 832.050 ;
        RECT 793.950 823.950 796.050 826.050 ;
        RECT 788.400 764.400 792.600 765.600 ;
        RECT 772.950 757.950 775.050 760.050 ;
        RECT 773.400 748.050 774.600 757.950 ;
        RECT 781.950 751.950 784.050 754.050 ;
        RECT 772.950 745.950 775.050 748.050 ;
        RECT 779.100 739.950 781.200 742.050 ;
        RECT 769.950 727.950 772.050 730.050 ;
        RECT 766.950 682.950 769.050 685.050 ;
        RECT 770.400 637.050 771.600 727.950 ;
        RECT 779.400 700.050 780.600 739.950 ;
        RECT 775.950 698.400 780.600 700.050 ;
        RECT 775.950 697.950 780.000 698.400 ;
        RECT 775.950 691.950 778.050 694.050 ;
        RECT 776.400 688.050 777.600 691.950 ;
        RECT 775.950 685.950 778.050 688.050 ;
        RECT 772.950 673.950 775.050 676.050 ;
        RECT 773.400 669.600 774.600 673.950 ;
        RECT 776.400 673.050 777.600 685.950 ;
        RECT 782.400 679.050 783.600 751.950 ;
        RECT 788.400 697.050 789.600 764.400 ;
        RECT 794.400 754.050 795.600 823.950 ;
        RECT 803.400 817.050 804.600 829.950 ;
        RECT 806.400 829.050 807.600 838.950 ;
        RECT 805.950 826.950 808.050 829.050 ;
        RECT 802.950 814.950 805.050 817.050 ;
        RECT 793.950 751.950 796.050 754.050 ;
        RECT 809.400 747.600 810.600 841.950 ;
        RECT 811.950 820.950 814.050 823.050 ;
        RECT 812.400 820.050 813.600 820.950 ;
        RECT 811.950 816.000 814.050 820.050 ;
        RECT 812.400 815.400 813.600 816.000 ;
        RECT 811.950 808.950 814.050 811.050 ;
        RECT 812.400 763.050 813.600 808.950 ;
        RECT 815.400 799.050 816.600 865.950 ;
        RECT 837.000 843.600 841.050 844.050 ;
        RECT 836.400 841.950 841.050 843.600 ;
        RECT 836.400 826.050 837.600 841.950 ;
        RECT 850.950 829.950 853.050 832.050 ;
        RECT 835.950 823.950 838.050 826.050 ;
        RECT 838.950 817.950 841.050 820.050 ;
        RECT 823.950 814.950 826.050 817.050 ;
        RECT 814.950 796.950 817.050 799.050 ;
        RECT 814.950 790.950 817.050 793.050 ;
        RECT 815.400 775.050 816.600 790.950 ;
        RECT 824.400 784.050 825.600 814.950 ;
        RECT 832.800 811.950 834.900 814.050 ;
        RECT 833.400 799.050 834.600 811.950 ;
        RECT 839.400 802.050 840.600 817.950 ;
        RECT 845.100 811.950 847.200 814.050 ;
        RECT 838.950 799.950 841.050 802.050 ;
        RECT 832.950 796.950 835.050 799.050 ;
        RECT 823.950 781.950 826.050 784.050 ;
        RECT 814.950 772.950 817.050 775.050 ;
        RECT 826.950 772.950 829.050 775.050 ;
        RECT 823.950 766.950 826.050 769.050 ;
        RECT 811.950 760.950 814.050 763.050 ;
        RECT 806.400 746.400 810.600 747.600 ;
        RECT 796.950 742.950 799.050 745.050 ;
        RECT 790.950 697.950 793.050 700.050 ;
        RECT 787.950 694.950 790.050 697.050 ;
        RECT 781.950 676.950 784.050 679.050 ;
        RECT 775.800 670.950 777.900 673.050 ;
        RECT 779.100 672.600 783.000 673.050 ;
        RECT 779.100 670.950 783.600 672.600 ;
        RECT 773.400 668.400 777.600 669.600 ;
        RECT 769.950 634.950 772.050 637.050 ;
        RECT 776.400 628.050 777.600 668.400 ;
        RECT 782.400 640.050 783.600 670.950 ;
        RECT 787.950 667.950 790.050 670.050 ;
        RECT 788.400 646.050 789.600 667.950 ;
        RECT 791.400 649.050 792.600 697.950 ;
        RECT 797.400 694.050 798.600 742.950 ;
        RECT 806.400 730.200 807.600 746.400 ;
        RECT 812.400 745.050 813.600 760.950 ;
        RECT 810.000 744.600 814.050 745.050 ;
        RECT 809.400 742.950 814.050 744.600 ;
        RECT 809.400 739.050 810.600 742.950 ;
        RECT 824.400 739.050 825.600 766.950 ;
        RECT 808.950 736.950 811.050 739.050 ;
        RECT 824.100 738.000 826.200 739.050 ;
        RECT 823.950 736.950 826.200 738.000 ;
        RECT 823.950 733.950 826.050 736.950 ;
        RECT 805.950 728.100 808.050 730.200 ;
        RECT 805.950 724.800 808.050 726.900 ;
        RECT 820.950 724.950 823.050 727.050 ;
        RECT 806.400 703.050 807.600 724.800 ;
        RECT 806.400 701.400 811.050 703.050 ;
        RECT 807.000 700.950 811.050 701.400 ;
        RECT 796.950 691.950 799.050 694.050 ;
        RECT 799.950 688.950 802.050 691.050 ;
        RECT 800.400 685.050 801.600 688.950 ;
        RECT 799.950 682.950 802.050 685.050 ;
        RECT 805.950 682.950 808.050 685.050 ;
        RECT 800.400 673.050 801.600 682.950 ;
        RECT 796.950 671.400 801.600 673.050 ;
        RECT 796.950 670.950 801.000 671.400 ;
        RECT 806.400 670.050 807.600 682.950 ;
        RECT 821.400 673.050 822.600 724.950 ;
        RECT 827.400 724.050 828.600 772.950 ;
        RECT 833.400 757.050 834.600 796.950 ;
        RECT 845.400 775.050 846.600 811.950 ;
        RECT 851.400 811.050 852.600 829.950 ;
        RECT 850.950 808.950 853.050 811.050 ;
        RECT 844.950 772.950 847.050 775.050 ;
        RECT 838.950 760.950 841.050 766.050 ;
        RECT 832.950 754.950 835.050 757.050 ;
        RECT 853.950 754.950 856.050 757.050 ;
        RECT 832.950 745.950 835.050 748.050 ;
        RECT 826.950 721.950 829.050 724.050 ;
        RECT 833.400 703.050 834.600 745.950 ;
        RECT 838.950 736.950 841.050 739.050 ;
        RECT 839.400 733.050 840.600 736.950 ;
        RECT 841.950 733.950 844.050 736.050 ;
        RECT 838.950 730.950 841.050 733.050 ;
        RECT 832.950 700.950 835.050 703.050 ;
        RECT 827.100 697.950 829.200 700.050 ;
        RECT 827.400 688.050 828.600 697.950 ;
        RECT 826.950 685.950 829.050 688.050 ;
        RECT 832.950 682.950 835.050 685.050 ;
        RECT 833.400 673.050 834.600 682.950 ;
        RECT 820.950 670.950 823.050 673.050 ;
        RECT 833.400 671.400 838.050 673.050 ;
        RECT 834.000 670.950 838.050 671.400 ;
        RECT 805.950 667.950 808.050 670.050 ;
        RECT 817.950 667.950 820.050 670.050 ;
        RECT 814.950 661.950 817.050 664.050 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 787.950 643.950 790.050 646.050 ;
        RECT 781.950 637.950 784.050 640.050 ;
        RECT 782.400 634.050 783.600 637.950 ;
        RECT 787.950 634.950 790.050 637.050 ;
        RECT 805.950 634.950 808.050 640.050 ;
        RECT 781.950 631.950 784.050 634.050 ;
        RECT 769.950 625.950 772.050 628.050 ;
        RECT 776.100 625.950 778.200 628.050 ;
        RECT 788.400 627.600 789.600 634.950 ;
        RECT 793.950 631.950 796.050 634.050 ;
        RECT 785.400 627.000 789.600 627.600 ;
        RECT 784.950 626.400 789.600 627.000 ;
        RECT 770.400 601.050 771.600 625.950 ;
        RECT 772.950 607.950 775.050 610.050 ;
        RECT 769.800 598.950 771.900 601.050 ;
        RECT 770.400 595.050 771.600 598.950 ;
        RECT 769.950 592.950 772.050 595.050 ;
        RECT 763.950 577.950 766.050 580.050 ;
        RECT 764.400 568.050 765.600 577.950 ;
        RECT 763.950 565.950 766.050 568.050 ;
        RECT 763.950 559.950 766.050 562.050 ;
        RECT 764.400 553.050 765.600 559.950 ;
        RECT 763.950 550.950 766.050 553.050 ;
        RECT 766.950 547.950 769.050 550.050 ;
        RECT 773.400 549.600 774.600 607.950 ;
        RECT 770.400 548.400 774.600 549.600 ;
        RECT 760.950 535.950 763.050 538.050 ;
        RECT 757.950 529.950 760.050 532.050 ;
        RECT 754.950 523.950 757.050 526.050 ;
        RECT 745.950 508.950 748.050 511.050 ;
        RECT 755.400 508.050 756.600 523.950 ;
        RECT 754.950 505.950 757.050 508.050 ;
        RECT 745.950 487.950 748.050 493.050 ;
        RECT 758.400 484.050 759.600 529.950 ;
        RECT 760.950 514.950 763.050 517.050 ;
        RECT 761.400 487.050 762.600 514.950 ;
        RECT 763.950 490.950 766.050 493.050 ;
        RECT 760.950 484.950 763.050 487.050 ;
        RECT 757.950 481.950 760.050 484.050 ;
        RECT 758.400 472.050 759.600 481.950 ;
        RECT 760.950 478.950 763.050 481.050 ;
        RECT 748.950 469.950 751.050 472.050 ;
        RECT 757.950 469.950 760.050 472.050 ;
        RECT 749.400 454.050 750.600 469.950 ;
        RECT 746.100 452.400 750.600 454.050 ;
        RECT 746.100 451.950 750.000 452.400 ;
        RECT 746.400 448.050 747.600 451.950 ;
        RECT 761.400 451.050 762.600 478.950 ;
        RECT 760.950 448.950 763.050 451.050 ;
        RECT 764.400 448.050 765.600 490.950 ;
        RECT 767.400 478.050 768.600 547.950 ;
        RECT 766.950 475.950 769.050 478.050 ;
        RECT 770.400 475.050 771.600 548.400 ;
        RECT 776.400 546.600 777.600 625.950 ;
        RECT 784.950 622.950 787.050 626.400 ;
        RECT 778.950 598.950 781.050 601.050 ;
        RECT 779.400 577.050 780.600 598.950 ;
        RECT 784.950 594.600 789.000 595.050 ;
        RECT 784.950 592.950 789.600 594.600 ;
        RECT 788.400 589.050 789.600 592.950 ;
        RECT 787.950 586.950 790.050 589.050 ;
        RECT 778.950 574.950 781.050 577.050 ;
        RECT 788.400 574.050 789.600 586.950 ;
        RECT 794.400 580.050 795.600 631.950 ;
        RECT 815.400 625.050 816.600 661.950 ;
        RECT 818.400 634.050 819.600 667.950 ;
        RECT 820.950 664.950 823.050 667.050 ;
        RECT 817.950 631.950 820.050 634.050 ;
        RECT 821.400 631.050 822.600 664.950 ;
        RECT 842.400 664.050 843.600 733.950 ;
        RECT 844.950 730.950 847.050 733.050 ;
        RECT 845.400 700.050 846.600 730.950 ;
        RECT 844.950 697.950 847.050 700.050 ;
        RECT 841.950 661.950 844.050 664.050 ;
        RECT 838.950 643.950 841.050 646.050 ;
        RECT 820.950 628.950 823.050 631.050 ;
        RECT 827.100 628.950 829.200 631.050 ;
        RECT 832.950 628.950 835.050 631.050 ;
        RECT 814.950 622.950 817.050 625.050 ;
        RECT 823.950 622.950 826.050 625.050 ;
        RECT 817.950 616.950 820.050 619.050 ;
        RECT 805.950 601.950 808.050 604.050 ;
        RECT 806.400 598.050 807.600 601.950 ;
        RECT 805.950 595.950 808.050 598.050 ;
        RECT 793.950 577.950 796.050 580.050 ;
        RECT 814.950 574.950 817.050 577.050 ;
        RECT 781.950 571.950 784.050 574.050 ;
        RECT 787.950 571.950 790.050 574.050 ;
        RECT 796.950 571.950 799.050 574.050 ;
        RECT 778.950 565.950 781.050 568.050 ;
        RECT 773.400 545.400 777.600 546.600 ;
        RECT 773.400 502.050 774.600 545.400 ;
        RECT 779.400 531.600 780.600 565.950 ;
        RECT 782.400 559.050 783.600 571.950 ;
        RECT 781.950 556.950 784.050 559.050 ;
        RECT 797.400 556.050 798.600 571.950 ;
        RECT 815.400 556.050 816.600 574.950 ;
        RECT 793.950 554.400 798.600 556.050 ;
        RECT 793.950 553.950 798.000 554.400 ;
        RECT 805.950 553.950 808.050 556.050 ;
        RECT 812.100 554.400 816.600 556.050 ;
        RECT 812.100 553.950 816.000 554.400 ;
        RECT 784.950 547.950 787.050 550.050 ;
        RECT 781.950 538.950 784.050 541.050 ;
        RECT 776.400 530.400 780.600 531.600 ;
        RECT 772.950 499.950 775.050 502.050 ;
        RECT 772.950 487.950 775.050 490.050 ;
        RECT 773.400 481.050 774.600 487.950 ;
        RECT 772.950 478.950 775.050 481.050 ;
        RECT 769.950 472.950 772.050 475.050 ;
        RECT 772.950 469.950 775.050 472.050 ;
        RECT 766.950 463.950 769.050 466.050 ;
        RECT 767.400 454.050 768.600 463.950 ;
        RECT 766.950 451.950 769.050 454.050 ;
        RECT 769.950 448.950 772.050 451.050 ;
        RECT 745.950 445.950 748.050 448.050 ;
        RECT 763.800 445.950 765.900 448.050 ;
        RECT 767.100 445.950 769.200 448.050 ;
        RECT 742.950 436.950 745.050 439.050 ;
        RECT 748.950 436.950 751.050 439.050 ;
        RECT 749.400 433.050 750.600 436.950 ;
        RECT 748.950 430.950 751.050 433.050 ;
        RECT 760.950 430.950 763.050 433.050 ;
        RECT 739.950 427.950 742.050 430.050 ;
        RECT 736.950 424.950 739.050 427.050 ;
        RECT 733.950 421.950 736.050 424.050 ;
        RECT 730.950 397.950 733.050 400.050 ;
        RECT 731.400 367.050 732.600 397.950 ;
        RECT 734.400 376.050 735.600 421.950 ;
        RECT 758.100 417.000 760.200 418.050 ;
        RECT 757.950 415.950 760.200 417.000 ;
        RECT 757.950 415.050 760.050 415.950 ;
        RECT 754.800 414.000 760.050 415.050 ;
        RECT 754.800 413.400 759.600 414.000 ;
        RECT 754.800 412.950 759.000 413.400 ;
        RECT 751.950 409.950 754.050 412.050 ;
        RECT 748.950 400.950 751.050 403.050 ;
        RECT 742.950 397.950 745.050 400.050 ;
        RECT 733.950 373.950 736.050 376.050 ;
        RECT 730.950 364.950 733.050 367.050 ;
        RECT 724.950 352.950 727.050 355.050 ;
        RECT 724.950 346.950 727.050 349.050 ;
        RECT 725.400 343.050 726.600 346.950 ;
        RECT 731.400 346.050 732.600 364.950 ;
        RECT 739.950 352.950 742.050 355.050 ;
        RECT 730.950 343.950 733.050 346.050 ;
        RECT 721.800 342.000 723.900 343.050 ;
        RECT 721.800 340.950 724.050 342.000 ;
        RECT 725.400 341.400 730.050 343.050 ;
        RECT 726.000 340.950 730.050 341.400 ;
        RECT 721.950 337.950 724.050 340.950 ;
        RECT 722.400 322.050 723.600 337.950 ;
        RECT 724.950 334.950 727.050 337.050 ;
        RECT 721.950 319.950 724.050 322.050 ;
        RECT 721.950 313.950 724.050 316.050 ;
        RECT 722.400 307.050 723.600 313.950 ;
        RECT 725.400 313.050 726.600 334.950 ;
        RECT 731.400 325.050 732.600 343.950 ;
        RECT 736.950 340.950 739.050 343.050 ;
        RECT 737.400 334.050 738.600 340.950 ;
        RECT 736.950 331.950 739.050 334.050 ;
        RECT 731.100 322.950 733.200 325.050 ;
        RECT 736.950 322.950 739.050 325.050 ;
        RECT 724.950 310.950 727.050 313.050 ;
        RECT 737.400 307.050 738.600 322.950 ;
        RECT 722.100 304.950 724.200 307.050 ;
        RECT 737.100 304.950 739.200 307.050 ;
        RECT 727.950 295.950 730.050 298.050 ;
        RECT 715.800 286.950 717.900 289.050 ;
        RECT 719.100 286.950 721.200 289.050 ;
        RECT 719.400 277.200 720.600 286.950 ;
        RECT 721.950 283.950 724.050 286.050 ;
        RECT 718.950 275.100 721.050 277.200 ;
        RECT 718.950 271.800 721.050 273.900 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 716.400 244.050 717.600 256.950 ;
        RECT 719.400 253.050 720.600 271.800 ;
        RECT 722.400 268.050 723.600 283.950 ;
        RECT 722.100 265.950 724.200 268.050 ;
        RECT 718.950 250.950 721.050 253.050 ;
        RECT 715.950 241.950 718.050 244.050 ;
        RECT 719.400 241.050 720.600 250.950 ;
        RECT 728.400 250.050 729.600 295.950 ;
        RECT 733.950 289.950 736.050 292.050 ;
        RECT 734.400 286.050 735.600 289.950 ;
        RECT 733.950 283.950 736.050 286.050 ;
        RECT 740.400 283.050 741.600 352.950 ;
        RECT 743.400 337.050 744.600 397.950 ;
        RECT 745.950 373.950 748.050 376.050 ;
        RECT 746.400 346.050 747.600 373.950 ;
        RECT 745.950 343.950 748.050 346.050 ;
        RECT 745.950 337.950 748.050 340.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 746.400 319.050 747.600 337.950 ;
        RECT 749.400 328.050 750.600 400.950 ;
        RECT 752.400 340.050 753.600 409.950 ;
        RECT 761.400 394.050 762.600 430.950 ;
        RECT 760.950 391.950 763.050 394.050 ;
        RECT 767.400 385.050 768.600 445.950 ;
        RECT 770.400 430.050 771.600 448.950 ;
        RECT 773.400 448.200 774.600 469.950 ;
        RECT 772.950 446.100 775.050 448.200 ;
        RECT 772.950 442.800 775.050 444.900 ;
        RECT 769.950 427.950 772.050 430.050 ;
        RECT 773.400 400.050 774.600 442.800 ;
        RECT 776.400 430.050 777.600 530.400 ;
        RECT 778.950 526.950 781.050 529.050 ;
        RECT 779.400 508.050 780.600 526.950 ;
        RECT 778.950 505.950 781.050 508.050 ;
        RECT 782.400 499.050 783.600 538.950 ;
        RECT 785.400 532.050 786.600 547.950 ;
        RECT 806.400 544.050 807.600 553.950 ;
        RECT 805.950 541.950 808.050 544.050 ;
        RECT 784.950 529.950 787.050 532.050 ;
        RECT 785.400 526.050 786.600 529.950 ;
        RECT 788.100 526.950 790.200 529.050 ;
        RECT 784.950 523.950 787.050 526.050 ;
        RECT 788.400 523.050 789.600 526.950 ;
        RECT 787.950 520.950 790.050 523.050 ;
        RECT 805.950 520.950 808.050 523.050 ;
        RECT 793.950 508.950 796.050 511.050 ;
        RECT 781.950 496.950 784.050 499.050 ;
        RECT 787.950 496.950 790.050 499.050 ;
        RECT 784.950 493.950 787.050 496.050 ;
        RECT 778.950 481.950 781.050 484.050 ;
        RECT 779.400 460.050 780.600 481.950 ;
        RECT 778.950 457.950 781.050 460.050 ;
        RECT 778.950 451.950 781.050 454.050 ;
        RECT 775.950 427.950 778.050 430.050 ;
        RECT 779.400 426.600 780.600 451.950 ;
        RECT 785.400 445.050 786.600 493.950 ;
        RECT 788.400 466.050 789.600 496.950 ;
        RECT 794.400 490.050 795.600 508.950 ;
        RECT 793.950 487.950 796.050 490.050 ;
        RECT 799.950 484.950 802.050 487.050 ;
        RECT 793.950 481.950 796.050 484.050 ;
        RECT 787.950 463.950 790.050 466.050 ;
        RECT 788.400 450.600 789.600 463.950 ;
        RECT 794.400 460.050 795.600 481.950 ;
        RECT 793.800 457.950 795.900 460.050 ;
        RECT 797.100 457.950 799.200 460.050 ;
        RECT 794.400 454.050 795.600 457.950 ;
        RECT 790.950 452.400 795.600 454.050 ;
        RECT 790.950 451.950 795.000 452.400 ;
        RECT 797.400 451.050 798.600 457.950 ;
        RECT 800.400 457.050 801.600 484.950 ;
        RECT 802.950 478.950 805.050 481.050 ;
        RECT 803.400 460.050 804.600 478.950 ;
        RECT 802.950 457.950 805.050 460.050 ;
        RECT 800.100 454.950 802.200 457.050 ;
        RECT 803.100 451.950 805.200 454.050 ;
        RECT 788.400 450.000 792.600 450.600 ;
        RECT 788.400 449.400 793.050 450.000 ;
        RECT 790.950 445.950 793.050 449.400 ;
        RECT 796.950 448.950 799.050 451.050 ;
        RECT 784.950 442.950 787.050 445.050 ;
        RECT 793.950 439.950 796.050 442.050 ;
        RECT 787.950 430.950 790.050 433.050 ;
        RECT 776.400 425.400 780.600 426.600 ;
        RECT 776.400 415.050 777.600 425.400 ;
        RECT 778.950 418.950 781.050 421.050 ;
        RECT 775.800 412.950 777.900 415.050 ;
        RECT 779.400 412.050 780.600 418.950 ;
        RECT 778.950 409.950 781.050 412.050 ;
        RECT 778.950 403.950 781.050 406.050 ;
        RECT 772.800 397.950 774.900 400.050 ;
        RECT 776.100 397.950 778.200 400.050 ;
        RECT 766.950 382.950 769.050 385.050 ;
        RECT 773.100 376.950 775.200 379.050 ;
        RECT 773.400 370.050 774.600 376.950 ;
        RECT 772.950 367.950 775.050 370.050 ;
        RECT 757.950 358.950 760.050 361.050 ;
        RECT 754.950 346.950 757.050 349.050 ;
        RECT 755.400 340.050 756.600 346.950 ;
        RECT 751.800 337.950 753.900 340.050 ;
        RECT 755.100 337.950 757.200 340.050 ;
        RECT 754.950 331.950 757.050 334.050 ;
        RECT 748.950 325.950 751.050 328.050 ;
        RECT 745.950 316.950 748.050 319.050 ;
        RECT 742.950 310.950 745.050 313.050 ;
        RECT 736.800 280.950 738.900 283.050 ;
        RECT 740.100 280.950 742.200 283.050 ;
        RECT 737.400 277.050 738.600 280.950 ;
        RECT 736.950 274.950 739.050 277.050 ;
        RECT 743.400 276.600 744.600 310.950 ;
        RECT 749.400 300.600 750.600 325.950 ;
        RECT 746.400 299.400 750.600 300.600 ;
        RECT 746.400 292.050 747.600 299.400 ;
        RECT 755.400 298.050 756.600 331.950 ;
        RECT 758.400 310.050 759.600 358.950 ;
        RECT 772.950 355.950 775.050 358.050 ;
        RECT 773.400 343.050 774.600 355.950 ;
        RECT 772.950 342.600 775.050 343.050 ;
        RECT 770.400 341.400 775.050 342.600 ;
        RECT 761.100 340.050 763.200 340.200 ;
        RECT 761.100 339.600 765.000 340.050 ;
        RECT 761.100 338.100 765.600 339.600 ;
        RECT 762.000 337.950 765.600 338.100 ;
        RECT 760.950 334.800 763.050 336.900 ;
        RECT 757.950 307.950 760.050 310.050 ;
        RECT 754.950 295.950 757.050 298.050 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 740.400 276.000 744.600 276.600 ;
        RECT 739.950 275.400 744.600 276.000 ;
        RECT 737.400 271.050 738.600 274.950 ;
        RECT 739.950 271.950 742.050 275.400 ;
        RECT 746.400 271.050 747.600 289.950 ;
        RECT 761.400 289.050 762.600 334.800 ;
        RECT 764.400 319.050 765.600 337.950 ;
        RECT 770.400 331.050 771.600 341.400 ;
        RECT 772.950 340.950 775.050 341.400 ;
        RECT 776.400 334.050 777.600 397.950 ;
        RECT 779.400 352.050 780.600 403.950 ;
        RECT 788.400 400.050 789.600 430.950 ;
        RECT 787.950 397.950 790.050 400.050 ;
        RECT 781.950 382.950 784.050 385.050 ;
        RECT 782.400 361.050 783.600 382.950 ;
        RECT 781.950 358.950 784.050 361.050 ;
        RECT 778.950 349.950 781.050 352.050 ;
        RECT 781.950 343.950 784.050 346.050 ;
        RECT 775.950 331.950 778.050 334.050 ;
        RECT 769.950 328.950 772.050 331.050 ;
        RECT 769.950 322.950 772.050 325.050 ;
        RECT 763.950 316.950 766.050 319.050 ;
        RECT 770.400 310.050 771.600 322.950 ;
        RECT 775.950 310.950 778.050 313.050 ;
        RECT 769.800 307.950 771.900 310.050 ;
        RECT 776.400 304.200 777.600 310.950 ;
        RECT 775.950 303.600 778.050 304.200 ;
        RECT 773.400 302.400 778.050 303.600 ;
        RECT 769.950 298.950 772.050 301.050 ;
        RECT 760.950 286.950 763.050 289.050 ;
        RECT 770.400 286.050 771.600 298.950 ;
        RECT 769.950 283.950 772.050 286.050 ;
        RECT 766.950 280.950 769.050 283.050 ;
        RECT 751.950 271.950 754.050 274.050 ;
        RECT 757.950 271.950 760.050 274.050 ;
        RECT 736.950 268.950 739.050 271.050 ;
        RECT 746.400 269.400 751.050 271.050 ;
        RECT 747.000 268.950 751.050 269.400 ;
        RECT 736.950 262.950 739.050 265.050 ;
        RECT 727.950 247.950 730.050 250.050 ;
        RECT 724.950 241.950 727.050 244.050 ;
        RECT 718.800 238.950 720.900 241.050 ;
        RECT 715.950 235.950 718.050 238.050 ;
        RECT 721.800 235.950 723.900 238.050 ;
        RECT 716.400 229.050 717.600 235.950 ;
        RECT 722.400 232.050 723.600 235.950 ;
        RECT 721.950 229.950 724.050 232.050 ;
        RECT 715.800 226.950 717.900 229.050 ;
        RECT 719.100 226.950 721.200 229.050 ;
        RECT 719.400 208.050 720.600 226.950 ;
        RECT 718.950 205.950 721.050 208.050 ;
        RECT 719.400 199.200 720.600 205.950 ;
        RECT 725.400 205.050 726.600 241.950 ;
        RECT 728.400 214.050 729.600 247.950 ;
        RECT 737.400 217.050 738.600 262.950 ;
        RECT 742.950 256.950 745.050 259.050 ;
        RECT 743.400 250.050 744.600 256.950 ;
        RECT 749.400 256.050 750.600 268.950 ;
        RECT 748.950 253.950 751.050 256.050 ;
        RECT 742.950 247.950 745.050 250.050 ;
        RECT 743.400 244.050 744.600 247.950 ;
        RECT 742.800 241.950 744.900 244.050 ;
        RECT 746.100 240.000 748.200 241.050 ;
        RECT 745.950 238.950 748.200 240.000 ;
        RECT 745.950 238.050 748.050 238.950 ;
        RECT 742.800 237.000 748.050 238.050 ;
        RECT 742.800 235.950 747.600 237.000 ;
        RECT 739.950 220.950 742.050 223.050 ;
        RECT 736.950 214.950 739.050 217.050 ;
        RECT 740.400 214.050 741.600 220.950 ;
        RECT 742.950 217.950 745.050 220.050 ;
        RECT 727.800 211.950 729.900 214.050 ;
        RECT 739.950 211.950 742.050 214.050 ;
        RECT 733.950 205.950 736.050 208.050 ;
        RECT 724.950 202.950 727.050 205.050 ;
        RECT 730.950 202.950 733.050 205.050 ;
        RECT 718.800 197.100 720.900 199.200 ;
        RECT 724.950 196.950 727.050 199.050 ;
        RECT 720.000 195.600 724.050 196.050 ;
        RECT 719.400 193.950 724.050 195.600 ;
        RECT 712.950 184.950 715.050 187.050 ;
        RECT 703.950 160.950 706.050 163.050 ;
        RECT 706.950 157.950 709.050 160.050 ;
        RECT 700.950 139.950 703.050 142.050 ;
        RECT 701.400 124.050 702.600 139.950 ;
        RECT 707.400 136.050 708.600 157.950 ;
        RECT 719.400 145.050 720.600 193.950 ;
        RECT 725.400 193.050 726.600 196.950 ;
        RECT 724.950 190.950 727.050 193.050 ;
        RECT 727.950 175.950 730.050 178.050 ;
        RECT 724.950 160.950 727.050 163.050 ;
        RECT 725.400 145.050 726.600 160.950 ;
        RECT 718.950 142.950 721.050 145.050 ;
        RECT 724.950 142.950 727.050 145.050 ;
        RECT 728.400 139.050 729.600 175.950 ;
        RECT 731.400 172.050 732.600 202.950 ;
        RECT 734.400 196.050 735.600 205.950 ;
        RECT 740.400 196.050 741.600 211.950 ;
        RECT 743.400 211.050 744.600 217.950 ;
        RECT 742.950 208.950 745.050 211.050 ;
        RECT 746.400 205.050 747.600 235.950 ;
        RECT 752.400 214.050 753.600 271.950 ;
        RECT 758.400 262.050 759.600 271.950 ;
        RECT 763.950 270.600 766.050 274.050 ;
        RECT 761.400 270.000 766.050 270.600 ;
        RECT 761.400 269.400 765.600 270.000 ;
        RECT 761.400 265.050 762.600 269.400 ;
        RECT 764.100 265.800 766.200 267.900 ;
        RECT 760.950 262.950 763.050 265.050 ;
        RECT 757.950 261.600 760.050 262.050 ;
        RECT 755.400 260.400 760.050 261.600 ;
        RECT 755.400 253.050 756.600 260.400 ;
        RECT 757.950 259.950 760.050 260.400 ;
        RECT 754.950 250.950 757.050 253.050 ;
        RECT 755.400 241.050 756.600 250.950 ;
        RECT 754.950 238.950 757.050 241.050 ;
        RECT 764.400 237.600 765.600 265.800 ;
        RECT 761.400 236.400 765.600 237.600 ;
        RECT 757.950 220.950 760.050 223.050 ;
        RECT 751.950 211.950 754.050 214.050 ;
        RECT 758.400 207.600 759.600 220.950 ;
        RECT 755.400 206.400 759.600 207.600 ;
        RECT 745.950 202.950 748.050 205.050 ;
        RECT 751.950 199.950 754.050 202.050 ;
        RECT 742.950 196.950 745.050 199.050 ;
        RECT 733.950 193.950 736.050 196.050 ;
        RECT 739.950 193.950 742.050 196.050 ;
        RECT 736.950 187.950 739.050 190.050 ;
        RECT 733.950 184.950 736.050 187.050 ;
        RECT 730.950 169.950 733.050 172.050 ;
        RECT 730.950 163.950 733.050 166.050 ;
        RECT 731.400 157.050 732.600 163.950 ;
        RECT 730.950 154.950 733.050 157.050 ;
        RECT 734.400 153.600 735.600 184.950 ;
        RECT 731.400 152.400 735.600 153.600 ;
        RECT 721.950 136.950 724.050 139.050 ;
        RECT 727.950 136.950 730.050 139.050 ;
        RECT 707.400 134.400 712.050 136.050 ;
        RECT 708.000 133.950 712.050 134.400 ;
        RECT 718.950 133.950 721.050 136.050 ;
        RECT 719.400 130.050 720.600 133.950 ;
        RECT 715.950 128.400 720.600 130.050 ;
        RECT 715.950 127.950 720.000 128.400 ;
        RECT 722.400 127.050 723.600 136.950 ;
        RECT 731.400 136.050 732.600 152.400 ;
        RECT 731.100 133.950 733.200 136.050 ;
        RECT 737.400 130.050 738.600 187.950 ;
        RECT 739.950 181.950 742.050 184.050 ;
        RECT 736.950 127.950 739.050 130.050 ;
        RECT 718.800 124.800 720.900 126.900 ;
        RECT 722.400 125.400 727.050 127.050 ;
        RECT 740.400 126.600 741.600 181.950 ;
        RECT 743.400 181.050 744.600 196.950 ;
        RECT 752.400 190.200 753.600 199.950 ;
        RECT 751.950 188.100 754.050 190.200 ;
        RECT 751.950 184.800 754.050 186.900 ;
        RECT 748.950 181.950 751.050 184.050 ;
        RECT 742.950 178.950 745.050 181.050 ;
        RECT 749.400 175.050 750.600 181.950 ;
        RECT 748.950 172.950 751.050 175.050 ;
        RECT 752.400 172.050 753.600 184.800 ;
        RECT 751.950 169.950 754.050 172.050 ;
        RECT 744.000 168.600 748.050 169.050 ;
        RECT 743.400 166.950 748.050 168.600 ;
        RECT 743.400 133.050 744.600 166.950 ;
        RECT 755.400 157.050 756.600 206.400 ;
        RECT 761.400 205.050 762.600 236.400 ;
        RECT 767.400 234.600 768.600 280.950 ;
        RECT 770.400 274.200 771.600 283.950 ;
        RECT 769.950 272.100 772.050 274.200 ;
        RECT 769.950 268.800 772.050 270.900 ;
        RECT 770.400 262.050 771.600 268.800 ;
        RECT 773.400 262.200 774.600 302.400 ;
        RECT 775.950 302.100 778.050 302.400 ;
        RECT 782.400 301.050 783.600 343.950 ;
        RECT 794.400 343.050 795.600 439.950 ;
        RECT 803.400 433.050 804.600 451.950 ;
        RECT 802.950 430.950 805.050 433.050 ;
        RECT 806.400 424.050 807.600 520.950 ;
        RECT 814.950 487.950 817.050 490.050 ;
        RECT 811.950 478.950 814.050 481.050 ;
        RECT 808.950 472.950 811.050 475.050 ;
        RECT 809.400 436.050 810.600 472.950 ;
        RECT 808.950 433.950 811.050 436.050 ;
        RECT 805.950 421.950 808.050 424.050 ;
        RECT 812.400 421.050 813.600 478.950 ;
        RECT 815.400 454.050 816.600 487.950 ;
        RECT 818.400 469.050 819.600 616.950 ;
        RECT 820.950 580.950 823.050 583.050 ;
        RECT 821.400 523.050 822.600 580.950 ;
        RECT 824.400 553.050 825.600 622.950 ;
        RECT 827.400 604.050 828.600 628.950 ;
        RECT 826.950 601.950 829.050 604.050 ;
        RECT 823.950 550.950 826.050 553.050 ;
        RECT 826.950 529.950 829.050 532.050 ;
        RECT 820.950 520.950 823.050 523.050 ;
        RECT 827.400 490.050 828.600 529.950 ;
        RECT 833.400 514.050 834.600 628.950 ;
        RECT 835.950 622.950 838.050 625.050 ;
        RECT 832.950 511.950 835.050 514.050 ;
        RECT 829.950 502.950 832.050 505.050 ;
        RECT 826.950 487.950 829.050 490.050 ;
        RECT 820.950 484.950 823.050 487.050 ;
        RECT 821.400 472.050 822.600 484.950 ;
        RECT 830.400 481.050 831.600 502.950 ;
        RECT 836.400 496.050 837.600 622.950 ;
        RECT 839.400 598.050 840.600 643.950 ;
        RECT 845.400 627.600 846.600 697.950 ;
        RECT 847.950 628.950 850.050 631.050 ;
        RECT 842.400 626.400 846.600 627.600 ;
        RECT 842.400 619.050 843.600 626.400 ;
        RECT 844.950 622.950 847.050 625.050 ;
        RECT 841.950 616.950 844.050 619.050 ;
        RECT 845.400 610.050 846.600 622.950 ;
        RECT 848.400 610.050 849.600 628.950 ;
        RECT 844.800 607.950 846.900 610.050 ;
        RECT 848.100 607.950 850.200 610.050 ;
        RECT 847.950 598.950 850.050 601.050 ;
        RECT 838.950 595.950 841.050 598.050 ;
        RECT 844.950 511.950 847.050 514.050 ;
        RECT 841.950 508.950 844.050 511.050 ;
        RECT 835.950 493.950 838.050 496.050 ;
        RECT 829.950 478.950 832.050 481.050 ;
        RECT 842.400 475.050 843.600 508.950 ;
        RECT 826.950 472.950 829.050 475.050 ;
        RECT 841.950 472.950 844.050 475.050 ;
        RECT 820.950 469.950 823.050 472.050 ;
        RECT 817.950 466.950 820.050 469.050 ;
        RECT 820.950 457.950 823.050 460.050 ;
        RECT 814.950 451.950 817.050 454.050 ;
        RECT 821.400 451.050 822.600 457.950 ;
        RECT 827.400 456.600 828.600 472.950 ;
        RECT 832.950 469.950 835.050 472.050 ;
        RECT 833.400 460.050 834.600 469.950 ;
        RECT 841.950 466.950 844.050 469.050 ;
        RECT 829.950 458.400 834.600 460.050 ;
        RECT 829.950 457.950 834.000 458.400 ;
        RECT 827.400 455.400 831.600 456.600 ;
        RECT 826.950 451.950 829.050 454.050 ;
        RECT 820.950 448.950 823.050 451.050 ;
        RECT 827.400 421.050 828.600 451.950 ;
        RECT 830.400 442.050 831.600 455.400 ;
        RECT 838.950 454.950 841.050 457.050 ;
        RECT 832.950 442.950 835.050 445.050 ;
        RECT 829.950 439.950 832.050 442.050 ;
        RECT 811.950 418.950 814.050 421.050 ;
        RECT 826.950 418.950 829.050 421.050 ;
        RECT 802.950 415.950 805.050 418.050 ;
        RECT 803.400 412.050 804.600 415.950 ;
        RECT 810.000 414.600 814.050 415.050 ;
        RECT 809.400 412.950 814.050 414.600 ;
        RECT 817.950 412.950 820.050 415.050 ;
        RECT 827.100 412.950 829.200 415.050 ;
        RECT 802.950 409.950 805.050 412.050 ;
        RECT 803.400 405.600 804.600 409.950 ;
        RECT 800.400 404.400 804.600 405.600 ;
        RECT 800.400 388.200 801.600 404.400 ;
        RECT 803.100 400.950 805.200 403.050 ;
        RECT 803.400 391.050 804.600 400.950 ;
        RECT 809.400 397.050 810.600 412.950 ;
        RECT 818.400 403.050 819.600 412.950 ;
        RECT 817.950 400.950 820.050 403.050 ;
        RECT 808.950 394.950 811.050 397.050 ;
        RECT 820.950 394.950 823.050 397.050 ;
        RECT 802.950 388.950 805.050 391.050 ;
        RECT 817.950 388.950 820.050 391.050 ;
        RECT 799.950 386.100 802.050 388.200 ;
        RECT 814.950 385.950 817.050 388.050 ;
        RECT 801.000 384.600 805.050 385.050 ;
        RECT 800.400 382.950 805.050 384.600 ;
        RECT 796.950 367.950 799.050 370.050 ;
        RECT 797.400 358.050 798.600 367.950 ;
        RECT 800.400 367.050 801.600 382.950 ;
        RECT 815.400 381.600 816.600 385.950 ;
        RECT 812.400 380.400 816.600 381.600 ;
        RECT 812.400 379.050 813.600 380.400 ;
        RECT 808.950 377.400 813.600 379.050 ;
        RECT 808.950 376.950 813.000 377.400 ;
        RECT 799.950 364.950 802.050 367.050 ;
        RECT 818.400 358.050 819.600 388.950 ;
        RECT 821.400 382.050 822.600 394.950 ;
        RECT 827.400 385.050 828.600 412.950 ;
        RECT 833.400 391.200 834.600 442.950 ;
        RECT 839.400 441.600 840.600 454.950 ;
        RECT 836.400 440.400 840.600 441.600 ;
        RECT 832.950 389.100 835.050 391.200 ;
        RECT 832.950 385.800 835.050 387.900 ;
        RECT 826.950 382.950 829.050 385.050 ;
        RECT 820.950 379.950 823.050 382.050 ;
        RECT 821.400 370.050 822.600 379.950 ;
        RECT 827.400 379.050 828.600 382.950 ;
        RECT 826.950 376.950 829.050 379.050 ;
        RECT 820.950 367.950 823.050 370.050 ;
        RECT 829.950 367.950 832.050 370.050 ;
        RECT 823.950 358.950 826.050 361.050 ;
        RECT 796.950 355.950 799.050 358.050 ;
        RECT 805.950 355.950 808.050 358.050 ;
        RECT 817.950 355.950 820.050 358.050 ;
        RECT 797.400 346.050 798.600 355.950 ;
        RECT 806.400 349.050 807.600 355.950 ;
        RECT 817.950 349.950 820.050 352.050 ;
        RECT 805.950 346.950 808.050 349.050 ;
        RECT 814.950 346.950 817.050 349.050 ;
        RECT 796.950 343.950 799.050 346.050 ;
        RECT 811.950 343.950 814.050 346.050 ;
        RECT 787.800 340.950 789.900 343.050 ;
        RECT 794.100 340.950 796.200 343.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 785.400 328.050 786.600 334.950 ;
        RECT 788.400 331.050 789.600 340.950 ;
        RECT 796.950 337.950 799.050 340.050 ;
        RECT 802.950 337.950 805.050 340.050 ;
        RECT 787.950 328.950 790.050 331.050 ;
        RECT 784.950 325.950 787.050 328.050 ;
        RECT 797.400 322.050 798.600 337.950 ;
        RECT 799.950 334.950 802.050 337.050 ;
        RECT 796.950 319.950 799.050 322.050 ;
        RECT 784.950 316.950 787.050 319.050 ;
        RECT 800.400 318.600 801.600 334.950 ;
        RECT 803.400 319.050 804.600 337.950 ;
        RECT 808.950 328.950 811.050 331.050 ;
        RECT 805.950 319.950 808.050 322.050 ;
        RECT 797.400 317.400 801.600 318.600 ;
        RECT 776.100 298.800 778.200 300.900 ;
        RECT 781.950 298.950 784.050 301.050 ;
        RECT 769.800 259.950 771.900 262.050 ;
        RECT 773.100 260.100 775.200 262.200 ;
        RECT 772.950 256.800 775.050 258.900 ;
        RECT 773.400 247.050 774.600 256.800 ;
        RECT 772.950 244.950 775.050 247.050 ;
        RECT 769.950 241.950 772.050 244.050 ;
        RECT 764.400 233.400 768.600 234.600 ;
        RECT 760.950 202.950 763.050 205.050 ;
        RECT 764.400 192.600 765.600 233.400 ;
        RECT 766.950 229.950 769.050 232.050 ;
        RECT 767.400 217.050 768.600 229.950 ;
        RECT 770.400 226.050 771.600 241.950 ;
        RECT 776.400 241.050 777.600 298.800 ;
        RECT 785.400 274.050 786.600 316.950 ;
        RECT 788.100 312.600 792.000 313.050 ;
        RECT 788.100 310.950 792.600 312.600 ;
        RECT 794.100 310.950 796.200 313.050 ;
        RECT 791.400 283.050 792.600 310.950 ;
        RECT 794.400 304.050 795.600 310.950 ;
        RECT 793.950 301.950 796.050 304.050 ;
        RECT 793.950 289.950 796.050 292.050 ;
        RECT 790.950 280.950 793.050 283.050 ;
        RECT 794.400 274.050 795.600 289.950 ;
        RECT 784.950 271.950 787.050 274.050 ;
        RECT 794.100 271.950 796.200 274.050 ;
        RECT 794.400 268.050 795.600 271.950 ;
        RECT 793.950 265.950 796.050 268.050 ;
        RECT 790.950 259.950 793.050 262.050 ;
        RECT 781.950 256.950 784.050 259.050 ;
        RECT 776.400 238.950 781.050 241.050 ;
        RECT 776.400 235.050 777.600 238.950 ;
        RECT 775.950 232.950 778.050 235.050 ;
        RECT 769.950 223.950 772.050 226.050 ;
        RECT 782.400 225.600 783.600 256.950 ;
        RECT 791.400 253.050 792.600 259.950 ;
        RECT 790.950 250.950 793.050 253.050 ;
        RECT 794.400 247.050 795.600 265.950 ;
        RECT 797.400 261.600 798.600 317.400 ;
        RECT 803.100 316.950 805.200 319.050 ;
        RECT 802.950 307.950 805.050 310.050 ;
        RECT 799.950 304.950 802.050 307.050 ;
        RECT 800.400 286.050 801.600 304.950 ;
        RECT 803.400 301.050 804.600 307.950 ;
        RECT 802.950 298.950 805.050 301.050 ;
        RECT 799.950 283.950 802.050 286.050 ;
        RECT 797.400 260.400 801.600 261.600 ;
        RECT 796.950 256.950 799.050 259.050 ;
        RECT 793.950 244.950 796.050 247.050 ;
        RECT 790.950 232.950 793.050 235.050 ;
        RECT 791.400 226.050 792.600 232.950 ;
        RECT 779.400 224.400 783.600 225.600 ;
        RECT 772.950 220.950 775.050 223.050 ;
        RECT 766.950 214.950 769.050 217.050 ;
        RECT 766.950 208.950 769.050 211.050 ;
        RECT 761.400 191.400 765.600 192.600 ;
        RECT 767.400 192.600 768.600 208.950 ;
        RECT 773.400 196.050 774.600 220.950 ;
        RECT 779.400 219.600 780.600 224.400 ;
        RECT 790.950 223.950 793.050 226.050 ;
        RECT 797.400 223.050 798.600 256.950 ;
        RECT 800.400 244.050 801.600 260.400 ;
        RECT 802.950 259.950 805.050 262.050 ;
        RECT 803.400 256.050 804.600 259.950 ;
        RECT 802.950 253.950 805.050 256.050 ;
        RECT 806.400 252.600 807.600 319.950 ;
        RECT 809.400 273.600 810.600 328.950 ;
        RECT 812.400 328.050 813.600 343.950 ;
        RECT 811.950 325.950 814.050 328.050 ;
        RECT 815.400 289.050 816.600 346.950 ;
        RECT 818.400 337.050 819.600 349.950 ;
        RECT 824.400 343.050 825.600 358.950 ;
        RECT 830.400 346.050 831.600 367.950 ;
        RECT 833.400 352.050 834.600 385.800 ;
        RECT 836.400 352.050 837.600 440.400 ;
        RECT 838.950 436.950 841.050 439.050 ;
        RECT 832.800 349.950 834.900 352.050 ;
        RECT 836.100 349.950 838.200 352.050 ;
        RECT 829.950 343.950 832.050 346.050 ;
        RECT 823.950 340.950 826.050 343.050 ;
        RECT 820.950 337.950 823.050 340.050 ;
        RECT 829.800 339.000 831.900 340.050 ;
        RECT 834.000 339.600 838.050 340.050 ;
        RECT 829.800 337.950 832.050 339.000 ;
        RECT 817.950 334.950 820.050 337.050 ;
        RECT 821.400 334.050 822.600 337.950 ;
        RECT 829.950 336.600 832.050 337.950 ;
        RECT 824.400 336.000 832.050 336.600 ;
        RECT 833.400 337.950 838.050 339.600 ;
        RECT 824.400 335.400 831.600 336.000 ;
        RECT 820.950 331.950 823.050 334.050 ;
        RECT 824.400 330.600 825.600 335.400 ;
        RECT 833.400 334.050 834.600 337.950 ;
        RECT 829.950 332.400 834.600 334.050 ;
        RECT 829.950 331.950 834.000 332.400 ;
        RECT 821.400 329.400 825.600 330.600 ;
        RECT 821.400 325.050 822.600 329.400 ;
        RECT 820.950 322.950 823.050 325.050 ;
        RECT 839.400 319.050 840.600 436.950 ;
        RECT 842.400 376.050 843.600 466.950 ;
        RECT 845.400 439.050 846.600 511.950 ;
        RECT 844.950 436.950 847.050 439.050 ;
        RECT 848.400 415.050 849.600 598.950 ;
        RECT 850.950 592.950 853.050 595.050 ;
        RECT 851.400 555.600 852.600 592.950 ;
        RECT 854.400 559.050 855.600 754.950 ;
        RECT 853.950 556.950 856.050 559.050 ;
        RECT 851.400 554.400 855.600 555.600 ;
        RECT 850.950 550.950 853.050 553.050 ;
        RECT 847.950 412.950 850.050 415.050 ;
        RECT 851.400 409.050 852.600 550.950 ;
        RECT 844.950 406.950 847.050 409.050 ;
        RECT 850.950 406.950 853.050 409.050 ;
        RECT 841.950 373.950 844.050 376.050 ;
        RECT 845.400 373.050 846.600 406.950 ;
        RECT 850.950 400.950 853.050 403.050 ;
        RECT 851.400 391.050 852.600 400.950 ;
        RECT 850.950 388.950 853.050 391.050 ;
        RECT 854.400 388.050 855.600 554.400 ;
        RECT 856.950 532.950 859.050 535.050 ;
        RECT 857.400 424.050 858.600 532.950 ;
        RECT 856.950 421.950 859.050 424.050 ;
        RECT 853.950 385.950 856.050 388.050 ;
        RECT 847.950 382.950 850.050 385.050 ;
        RECT 844.950 370.950 847.050 373.050 ;
        RECT 841.950 325.950 844.050 328.050 ;
        RECT 817.950 316.950 820.050 319.050 ;
        RECT 826.950 316.950 829.050 319.050 ;
        RECT 838.950 316.950 841.050 319.050 ;
        RECT 818.400 294.600 819.600 316.950 ;
        RECT 818.400 293.400 822.600 294.600 ;
        RECT 814.950 286.950 817.050 289.050 ;
        RECT 821.400 285.600 822.600 293.400 ;
        RECT 821.400 284.400 825.600 285.600 ;
        RECT 820.950 280.950 823.050 283.050 ;
        RECT 809.400 272.400 813.600 273.600 ;
        RECT 812.400 262.050 813.600 272.400 ;
        RECT 814.950 265.950 817.050 268.050 ;
        RECT 811.950 259.950 814.050 262.050 ;
        RECT 815.400 256.200 816.600 265.950 ;
        RECT 817.950 259.950 820.050 262.050 ;
        RECT 811.800 253.950 813.900 256.050 ;
        RECT 815.100 254.100 817.200 256.200 ;
        RECT 803.400 251.400 807.600 252.600 ;
        RECT 799.950 241.950 802.050 244.050 ;
        RECT 796.800 220.950 798.900 223.050 ;
        RECT 800.100 220.950 802.200 223.050 ;
        RECT 776.400 218.400 780.600 219.600 ;
        RECT 776.400 208.050 777.600 218.400 ;
        RECT 784.950 217.950 787.050 220.050 ;
        RECT 775.950 205.950 778.050 208.050 ;
        RECT 772.800 193.950 774.900 196.050 ;
        RECT 779.100 193.950 781.200 196.050 ;
        RECT 769.950 192.600 772.050 193.050 ;
        RECT 767.400 191.400 772.050 192.600 ;
        RECT 748.950 154.950 751.050 157.050 ;
        RECT 754.950 154.950 757.050 157.050 ;
        RECT 749.400 148.050 750.600 154.950 ;
        RECT 761.400 154.050 762.600 191.400 ;
        RECT 769.950 190.950 772.050 191.400 ;
        RECT 763.950 187.950 766.050 190.050 ;
        RECT 764.400 175.050 765.600 187.950 ;
        RECT 770.400 178.050 771.600 190.950 ;
        RECT 779.400 190.050 780.600 193.950 ;
        RECT 778.950 187.950 781.050 190.050 ;
        RECT 785.400 184.050 786.600 217.950 ;
        RECT 796.950 214.950 799.050 217.050 ;
        RECT 790.950 211.950 793.050 214.050 ;
        RECT 787.950 202.950 790.050 205.050 ;
        RECT 784.950 181.950 787.050 184.050 ;
        RECT 769.950 175.950 772.050 178.050 ;
        RECT 788.400 175.050 789.600 202.950 ;
        RECT 763.950 172.950 766.050 175.050 ;
        RECT 772.950 172.950 775.050 175.050 ;
        RECT 787.950 172.950 790.050 175.050 ;
        RECT 766.950 166.950 769.050 169.050 ;
        RECT 767.400 163.050 768.600 166.950 ;
        RECT 773.400 166.050 774.600 172.950 ;
        RECT 775.950 169.950 778.050 172.050 ;
        RECT 769.950 164.400 774.600 166.050 ;
        RECT 769.950 163.950 774.000 164.400 ;
        RECT 766.950 160.950 769.050 163.050 ;
        RECT 751.950 151.950 754.050 154.050 ;
        RECT 760.950 151.950 763.050 154.050 ;
        RECT 748.950 145.950 751.050 148.050 ;
        RECT 745.950 136.950 748.050 139.050 ;
        RECT 742.950 130.950 745.050 133.050 ;
        RECT 723.000 124.950 727.050 125.400 ;
        RECT 737.400 125.400 741.600 126.600 ;
        RECT 701.400 122.400 706.050 124.050 ;
        RECT 702.000 121.950 706.050 122.400 ;
        RECT 694.950 118.950 697.050 121.050 ;
        RECT 688.950 115.950 691.050 118.050 ;
        RECT 679.950 109.950 682.050 112.050 ;
        RECT 676.950 103.950 679.050 106.050 ;
        RECT 689.400 103.050 690.600 115.950 ;
        RECT 688.950 100.950 691.050 103.050 ;
        RECT 676.950 97.950 679.050 100.050 ;
        RECT 677.400 91.050 678.600 97.950 ;
        RECT 695.400 97.050 696.600 118.950 ;
        RECT 712.950 106.950 715.050 109.050 ;
        RECT 700.950 103.950 703.050 106.050 ;
        RECT 694.950 94.950 697.050 97.050 ;
        RECT 701.400 94.050 702.600 103.950 ;
        RECT 706.950 94.950 709.050 97.050 ;
        RECT 697.950 92.400 702.600 94.050 ;
        RECT 697.950 91.950 702.000 92.400 ;
        RECT 676.950 88.950 679.050 91.050 ;
        RECT 682.950 76.950 685.050 79.050 ;
        RECT 670.950 67.950 673.050 70.050 ;
        RECT 683.400 67.050 684.600 76.950 ;
        RECT 688.950 73.950 691.050 76.050 ;
        RECT 682.950 64.950 685.050 67.050 ;
        RECT 689.400 61.050 690.600 73.950 ;
        RECT 700.950 70.950 703.050 73.050 ;
        RECT 697.950 67.950 700.050 70.050 ;
        RECT 694.950 64.950 697.050 67.050 ;
        RECT 631.950 58.950 634.050 61.050 ;
        RECT 688.800 58.950 690.900 61.050 ;
        RECT 695.400 58.050 696.600 64.950 ;
        RECT 625.950 55.950 628.050 58.050 ;
        RECT 646.800 57.600 648.900 58.050 ;
        RECT 653.100 57.600 655.200 58.050 ;
        RECT 646.800 56.400 655.200 57.600 ;
        RECT 646.800 55.950 648.900 56.400 ;
        RECT 653.100 55.950 655.200 56.400 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 692.100 56.400 696.600 58.050 ;
        RECT 692.100 55.950 696.000 56.400 ;
        RECT 626.400 52.050 627.600 55.950 ;
        RECT 625.950 49.950 628.050 52.050 ;
        RECT 665.400 40.050 666.600 55.950 ;
        RECT 670.800 54.600 672.900 55.050 ;
        RECT 679.950 54.600 682.050 55.050 ;
        RECT 670.800 53.400 682.050 54.600 ;
        RECT 670.800 52.950 672.900 53.400 ;
        RECT 679.950 52.950 682.050 53.400 ;
        RECT 683.400 43.050 684.600 55.950 ;
        RECT 691.950 43.950 694.050 46.050 ;
        RECT 682.950 40.950 685.050 43.050 ;
        RECT 664.950 37.950 667.050 40.050 ;
        RECT 692.400 28.050 693.600 43.950 ;
        RECT 698.400 37.050 699.600 67.950 ;
        RECT 701.400 46.050 702.600 70.950 ;
        RECT 707.400 70.050 708.600 94.950 ;
        RECT 713.400 94.050 714.600 106.950 ;
        RECT 719.400 106.050 720.600 124.800 ;
        RECT 733.950 112.950 736.050 115.050 ;
        RECT 730.950 106.950 733.050 109.050 ;
        RECT 718.950 103.950 721.050 106.050 ;
        RECT 727.950 103.950 730.050 106.050 ;
        RECT 712.950 91.950 715.050 94.050 ;
        RECT 725.100 93.000 727.200 94.050 ;
        RECT 724.950 91.950 727.200 93.000 ;
        RECT 724.950 91.050 727.050 91.950 ;
        RECT 721.800 90.000 727.050 91.050 ;
        RECT 721.800 89.400 726.600 90.000 ;
        RECT 721.800 88.950 726.000 89.400 ;
        RECT 728.400 88.050 729.600 103.950 ;
        RECT 727.950 85.950 730.050 88.050 ;
        RECT 721.950 79.950 724.050 82.050 ;
        RECT 722.400 70.050 723.600 79.950 ;
        RECT 706.950 67.950 709.050 70.050 ;
        RECT 721.950 67.950 724.050 70.050 ;
        RECT 707.400 60.600 708.600 67.950 ;
        RECT 704.400 59.400 708.600 60.600 ;
        RECT 704.400 55.050 705.600 59.400 ;
        RECT 712.950 58.950 715.050 64.050 ;
        RECT 722.400 55.050 723.600 67.950 ;
        RECT 703.950 52.950 706.050 55.050 ;
        RECT 721.950 52.950 724.050 55.050 ;
        RECT 724.950 51.600 727.050 52.050 ;
        RECT 731.400 51.600 732.600 106.950 ;
        RECT 724.950 50.400 732.600 51.600 ;
        RECT 724.950 49.950 727.050 50.400 ;
        RECT 700.950 43.950 703.050 46.050 ;
        RECT 724.950 40.950 727.050 43.050 ;
        RECT 718.950 37.950 721.050 40.050 ;
        RECT 697.950 34.950 700.050 37.050 ;
        RECT 658.950 25.950 661.050 28.050 ;
        RECT 691.950 25.950 694.050 28.050 ;
        RECT 715.950 25.950 718.050 28.050 ;
        RECT 614.400 23.400 619.050 25.050 ;
        RECT 615.000 22.950 619.050 23.400 ;
        RECT 637.950 22.950 640.050 25.050 ;
        RECT 625.950 16.950 628.050 19.050 ;
        RECT 631.950 16.950 634.050 22.050 ;
        RECT 626.400 10.050 627.600 16.950 ;
        RECT 638.400 16.050 639.600 22.950 ;
        RECT 659.400 19.050 660.600 25.950 ;
        RECT 685.950 22.050 688.050 25.050 ;
        RECT 692.400 22.050 693.600 25.950 ;
        RECT 679.950 19.950 682.050 22.050 ;
        RECT 685.800 21.000 688.050 22.050 ;
        RECT 685.800 19.950 687.900 21.000 ;
        RECT 691.950 19.950 694.050 22.050 ;
        RECT 655.950 17.400 660.600 19.050 ;
        RECT 655.950 16.950 660.000 17.400 ;
        RECT 637.800 13.950 639.900 16.050 ;
        RECT 641.100 15.000 643.200 16.050 ;
        RECT 640.950 13.950 643.200 15.000 ;
        RECT 646.950 13.950 649.050 16.050 ;
        RECT 640.950 10.950 643.050 13.950 ;
        RECT 647.400 10.050 648.600 13.950 ;
        RECT 625.950 7.950 628.050 10.050 ;
        RECT 646.950 7.950 649.050 10.050 ;
        RECT 464.400 6.000 468.600 6.600 ;
        RECT 463.950 5.400 468.600 6.000 ;
        RECT 448.950 1.950 451.050 4.050 ;
        RECT 463.950 1.950 466.050 5.400 ;
        RECT 517.950 4.950 520.050 7.050 ;
        RECT 610.950 4.950 613.050 7.050 ;
        RECT 680.400 4.050 681.600 19.950 ;
        RECT 716.400 19.050 717.600 25.950 ;
        RECT 719.400 25.050 720.600 37.950 ;
        RECT 718.950 22.950 721.050 25.050 ;
        RECT 725.400 22.050 726.600 40.950 ;
        RECT 725.400 20.400 730.050 22.050 ;
        RECT 726.000 19.950 730.050 20.400 ;
        RECT 734.400 19.050 735.600 112.950 ;
        RECT 737.400 79.050 738.600 125.400 ;
        RECT 739.950 109.950 742.050 112.050 ;
        RECT 736.950 76.950 739.050 79.050 ;
        RECT 736.950 58.950 739.050 61.050 ;
        RECT 737.400 22.050 738.600 58.950 ;
        RECT 740.400 28.050 741.600 109.950 ;
        RECT 742.950 91.950 745.050 94.050 ;
        RECT 743.400 61.050 744.600 91.950 ;
        RECT 746.400 67.050 747.600 136.950 ;
        RECT 748.800 124.950 750.900 127.050 ;
        RECT 749.400 121.050 750.600 124.950 ;
        RECT 748.950 118.950 751.050 121.050 ;
        RECT 748.950 112.950 751.050 115.050 ;
        RECT 749.400 94.050 750.600 112.950 ;
        RECT 748.950 91.950 751.050 94.050 ;
        RECT 748.950 73.950 751.050 76.050 ;
        RECT 745.950 64.950 748.050 67.050 ;
        RECT 749.400 61.050 750.600 73.950 ;
        RECT 742.950 58.950 745.050 61.050 ;
        RECT 748.950 58.950 751.050 61.050 ;
        RECT 752.400 49.050 753.600 151.950 ;
        RECT 766.950 148.950 769.050 151.050 ;
        RECT 763.950 145.950 766.050 148.050 ;
        RECT 757.950 136.950 760.050 139.050 ;
        RECT 754.950 133.950 757.050 136.050 ;
        RECT 755.400 106.050 756.600 133.950 ;
        RECT 754.950 103.950 757.050 106.050 ;
        RECT 758.400 97.050 759.600 136.950 ;
        RECT 754.800 95.400 759.600 97.050 ;
        RECT 754.800 94.950 759.000 95.400 ;
        RECT 760.950 94.950 763.050 97.050 ;
        RECT 754.950 82.950 757.050 85.050 ;
        RECT 755.400 64.050 756.600 82.950 ;
        RECT 761.400 76.050 762.600 94.950 ;
        RECT 760.950 73.950 763.050 76.050 ;
        RECT 764.400 64.050 765.600 145.950 ;
        RECT 754.950 61.950 757.050 64.050 ;
        RECT 763.950 61.950 766.050 64.050 ;
        RECT 755.400 58.050 756.600 61.950 ;
        RECT 755.400 56.400 760.050 58.050 ;
        RECT 756.000 55.950 760.050 56.400 ;
        RECT 751.950 46.950 754.050 49.050 ;
        RECT 757.950 46.950 760.050 49.050 ;
        RECT 763.950 46.950 766.050 49.050 ;
        RECT 742.950 28.950 745.050 31.050 ;
        RECT 739.950 25.950 742.050 28.050 ;
        RECT 743.400 25.050 744.600 28.950 ;
        RECT 758.400 25.050 759.600 46.950 ;
        RECT 764.400 40.050 765.600 46.950 ;
        RECT 767.400 43.050 768.600 148.950 ;
        RECT 769.950 142.950 772.050 145.050 ;
        RECT 770.400 103.050 771.600 142.950 ;
        RECT 776.400 139.050 777.600 169.950 ;
        RECT 788.400 166.050 789.600 172.950 ;
        RECT 780.000 165.600 784.050 166.050 ;
        RECT 779.400 163.950 784.050 165.600 ;
        RECT 787.950 163.950 790.050 166.050 ;
        RECT 779.400 160.050 780.600 163.950 ;
        RECT 791.400 163.050 792.600 211.950 ;
        RECT 797.400 198.600 798.600 214.950 ;
        RECT 794.400 197.400 798.600 198.600 ;
        RECT 794.400 190.050 795.600 197.400 ;
        RECT 796.950 193.950 799.050 196.050 ;
        RECT 793.950 187.950 796.050 190.050 ;
        RECT 797.400 181.050 798.600 193.950 ;
        RECT 800.400 184.050 801.600 220.950 ;
        RECT 799.950 181.950 802.050 184.050 ;
        RECT 796.950 178.950 799.050 181.050 ;
        RECT 803.400 180.600 804.600 251.400 ;
        RECT 808.950 241.950 811.050 244.050 ;
        RECT 809.400 214.200 810.600 241.950 ;
        RECT 812.400 217.050 813.600 253.950 ;
        RECT 814.950 250.800 817.050 252.900 ;
        RECT 811.950 214.950 814.050 217.050 ;
        RECT 808.950 212.100 811.050 214.200 ;
        RECT 815.400 211.050 816.600 250.800 ;
        RECT 818.400 220.050 819.600 259.950 ;
        RECT 821.400 250.050 822.600 280.950 ;
        RECT 820.950 247.950 823.050 250.050 ;
        RECT 824.400 243.600 825.600 284.400 ;
        RECT 827.400 283.050 828.600 316.950 ;
        RECT 832.950 310.950 835.050 316.050 ;
        RECT 835.950 307.950 838.050 310.050 ;
        RECT 832.950 295.950 835.050 298.050 ;
        RECT 833.400 283.050 834.600 295.950 ;
        RECT 836.400 285.600 837.600 307.950 ;
        RECT 842.400 304.050 843.600 325.950 ;
        RECT 848.400 304.050 849.600 382.950 ;
        RECT 850.950 376.950 853.050 379.050 ;
        RECT 851.400 358.050 852.600 376.950 ;
        RECT 853.950 373.950 856.050 376.050 ;
        RECT 850.950 355.950 853.050 358.050 ;
        RECT 850.950 349.950 853.050 352.050 ;
        RECT 851.400 310.050 852.600 349.950 ;
        RECT 850.950 307.950 853.050 310.050 ;
        RECT 841.950 301.950 844.050 304.050 ;
        RECT 847.950 301.950 850.050 304.050 ;
        RECT 854.400 301.050 855.600 373.950 ;
        RECT 856.950 367.950 859.050 370.050 ;
        RECT 857.400 361.050 858.600 367.950 ;
        RECT 856.950 358.950 859.050 361.050 ;
        RECT 856.950 352.950 859.050 355.050 ;
        RECT 857.400 316.050 858.600 352.950 ;
        RECT 856.950 313.950 859.050 316.050 ;
        RECT 844.950 298.950 847.050 301.050 ;
        RECT 853.950 298.950 856.050 301.050 ;
        RECT 845.400 295.050 846.600 298.950 ;
        RECT 847.950 295.950 850.050 298.050 ;
        RECT 844.950 292.950 847.050 295.050 ;
        RECT 841.950 286.950 844.050 289.050 ;
        RECT 836.400 284.400 840.600 285.600 ;
        RECT 826.800 280.950 828.900 283.050 ;
        RECT 832.950 280.950 835.050 283.050 ;
        RECT 839.400 274.050 840.600 284.400 ;
        RECT 838.950 271.950 841.050 274.050 ;
        RECT 835.950 268.950 838.050 271.050 ;
        RECT 829.950 259.950 832.050 262.050 ;
        RECT 826.950 253.950 829.050 256.050 ;
        RECT 821.400 242.400 825.600 243.600 ;
        RECT 817.950 217.950 820.050 220.050 ;
        RECT 821.400 213.600 822.600 242.400 ;
        RECT 827.400 241.050 828.600 253.950 ;
        RECT 823.950 239.400 828.600 241.050 ;
        RECT 823.950 238.950 828.000 239.400 ;
        RECT 824.400 235.050 825.600 238.950 ;
        RECT 830.400 238.050 831.600 259.950 ;
        RECT 832.950 256.950 835.050 259.050 ;
        RECT 833.400 253.050 834.600 256.950 ;
        RECT 832.950 250.950 835.050 253.050 ;
        RECT 836.400 238.050 837.600 268.950 ;
        RECT 839.400 267.000 840.600 267.600 ;
        RECT 838.950 262.950 841.050 267.000 ;
        RECT 839.400 250.050 840.600 262.950 ;
        RECT 838.950 247.950 841.050 250.050 ;
        RECT 842.400 247.050 843.600 286.950 ;
        RECT 844.950 262.950 847.050 265.050 ;
        RECT 845.400 256.050 846.600 262.950 ;
        RECT 844.950 253.950 847.050 256.050 ;
        RECT 841.950 244.950 844.050 247.050 ;
        RECT 844.950 241.950 847.050 244.050 ;
        RECT 841.950 238.950 844.050 241.050 ;
        RECT 828.000 237.900 831.600 238.050 ;
        RECT 826.950 236.250 831.600 237.900 ;
        RECT 833.100 236.400 837.600 238.050 ;
        RECT 826.950 235.950 831.000 236.250 ;
        RECT 833.100 235.950 837.000 236.400 ;
        RECT 826.950 235.800 829.050 235.950 ;
        RECT 823.950 232.950 826.050 235.050 ;
        RECT 838.950 232.950 841.050 235.050 ;
        RECT 824.400 229.050 825.600 232.950 ;
        RECT 823.950 228.600 826.050 229.050 ;
        RECT 823.950 227.400 828.600 228.600 ;
        RECT 823.950 226.950 826.050 227.400 ;
        RECT 821.400 212.400 825.600 213.600 ;
        RECT 808.950 208.800 811.050 210.900 ;
        RECT 814.950 208.950 817.050 211.050 ;
        RECT 805.950 193.950 808.050 196.050 ;
        RECT 800.400 179.400 804.600 180.600 ;
        RECT 796.950 169.950 799.050 172.050 ;
        RECT 790.950 160.950 793.050 163.050 ;
        RECT 797.400 160.050 798.600 169.950 ;
        RECT 778.950 157.950 781.050 160.050 ;
        RECT 796.950 157.950 799.050 160.050 ;
        RECT 775.950 136.950 778.050 139.050 ;
        RECT 779.400 136.050 780.600 157.950 ;
        RECT 793.950 139.950 796.050 142.050 ;
        RECT 784.950 136.950 787.050 139.050 ;
        RECT 778.950 133.950 781.050 136.050 ;
        RECT 785.400 133.050 786.600 136.950 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 775.950 130.950 778.050 133.050 ;
        RECT 784.950 130.950 787.050 133.050 ;
        RECT 776.400 127.050 777.600 130.950 ;
        RECT 775.950 124.950 778.050 127.050 ;
        RECT 772.950 121.950 775.050 124.050 ;
        RECT 773.400 118.050 774.600 121.950 ;
        RECT 772.950 115.950 775.050 118.050 ;
        RECT 791.400 109.050 792.600 133.950 ;
        RECT 794.400 130.050 795.600 139.950 ;
        RECT 800.400 136.050 801.600 179.400 ;
        RECT 806.400 169.050 807.600 193.950 ;
        RECT 805.950 166.950 808.050 169.050 ;
        RECT 809.400 142.050 810.600 208.800 ;
        RECT 824.400 208.050 825.600 212.400 ;
        RECT 827.400 211.050 828.600 227.400 ;
        RECT 830.100 226.950 832.200 229.050 ;
        RECT 826.950 208.950 829.050 211.050 ;
        RECT 823.950 205.950 826.050 208.050 ;
        RECT 817.950 202.950 820.050 205.050 ;
        RECT 811.950 199.950 814.050 202.050 ;
        RECT 812.400 196.050 813.600 199.950 ;
        RECT 818.400 199.050 819.600 202.950 ;
        RECT 818.100 196.950 820.200 199.050 ;
        RECT 812.100 193.950 814.200 196.050 ;
        RECT 820.950 187.950 823.050 190.050 ;
        RECT 811.950 169.950 814.050 172.050 ;
        RECT 808.950 139.950 811.050 142.050 ;
        RECT 799.950 133.950 802.050 136.050 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 793.950 127.950 796.050 130.050 ;
        RECT 802.950 127.950 805.050 133.050 ;
        RECT 809.400 124.050 810.600 133.950 ;
        RECT 809.100 121.950 811.200 124.050 ;
        RECT 802.950 118.950 805.050 121.050 ;
        RECT 790.950 106.950 793.050 109.050 ;
        RECT 799.950 106.950 802.050 109.050 ;
        RECT 769.950 100.950 772.050 103.050 ;
        RECT 778.950 97.950 781.050 100.050 ;
        RECT 779.400 94.050 780.600 97.950 ;
        RECT 791.400 97.200 792.600 106.950 ;
        RECT 796.950 103.950 799.050 106.050 ;
        RECT 790.950 95.100 793.050 97.200 ;
        RECT 769.950 91.950 772.050 94.050 ;
        RECT 775.950 92.400 780.600 94.050 ;
        RECT 792.000 93.900 795.000 94.050 ;
        RECT 790.950 93.450 795.000 93.900 ;
        RECT 775.950 91.950 780.000 92.400 ;
        RECT 790.950 91.950 795.600 93.450 ;
        RECT 770.400 48.600 771.600 91.950 ;
        RECT 790.950 91.800 793.050 91.950 ;
        RECT 785.100 90.000 787.200 91.050 ;
        RECT 784.950 88.950 787.200 90.000 ;
        RECT 784.950 88.050 787.050 88.950 ;
        RECT 781.800 85.950 783.900 88.050 ;
        RECT 784.950 87.000 787.200 88.050 ;
        RECT 785.100 85.950 787.200 87.000 ;
        RECT 782.400 76.050 783.600 85.950 ;
        RECT 794.400 82.050 795.600 91.950 ;
        RECT 793.950 79.950 796.050 82.050 ;
        RECT 772.950 73.950 775.050 76.050 ;
        RECT 781.950 73.950 784.050 76.050 ;
        RECT 773.400 61.050 774.600 73.950 ;
        RECT 784.950 70.950 787.050 73.050 ;
        RECT 772.950 58.950 775.050 61.050 ;
        RECT 785.400 58.050 786.600 70.950 ;
        RECT 797.400 61.050 798.600 103.950 ;
        RECT 796.950 58.950 799.050 61.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 797.400 55.050 798.600 58.950 ;
        RECT 772.800 54.600 774.900 55.050 ;
        RECT 779.100 54.600 781.200 55.050 ;
        RECT 772.800 53.400 781.200 54.600 ;
        RECT 772.800 52.950 774.900 53.400 ;
        RECT 779.100 52.950 781.200 53.400 ;
        RECT 794.100 53.400 798.600 55.050 ;
        RECT 794.100 52.950 798.000 53.400 ;
        RECT 770.400 47.400 786.600 48.600 ;
        RECT 766.950 40.950 769.050 43.050 ;
        RECT 763.950 37.950 766.050 40.050 ;
        RECT 775.950 37.950 778.050 40.050 ;
        RECT 742.950 22.950 745.050 25.050 ;
        RECT 757.950 22.950 760.050 25.050 ;
        RECT 776.400 22.050 777.600 37.950 ;
        RECT 737.400 20.400 742.050 22.050 ;
        RECT 738.000 19.950 742.050 20.400 ;
        RECT 766.950 19.950 769.050 22.050 ;
        RECT 775.950 19.950 778.050 22.050 ;
        RECT 715.950 16.950 718.050 19.050 ;
        RECT 730.950 17.400 735.600 19.050 ;
        RECT 730.950 16.950 735.000 17.400 ;
        RECT 745.950 15.600 748.050 16.050 ;
        RECT 745.950 14.400 762.600 15.600 ;
        RECT 745.950 13.950 748.050 14.400 ;
        RECT 679.950 1.950 682.050 4.050 ;
        RECT 761.400 3.600 762.600 14.400 ;
        RECT 767.400 7.050 768.600 19.950 ;
        RECT 785.400 13.050 786.600 47.400 ;
        RECT 790.950 34.950 793.050 37.050 ;
        RECT 791.400 28.050 792.600 34.950 ;
        RECT 796.950 28.950 799.050 31.050 ;
        RECT 790.950 25.950 793.050 28.050 ;
        RECT 797.400 25.050 798.600 28.950 ;
        RECT 796.950 22.950 799.050 25.050 ;
        RECT 800.400 22.050 801.600 106.950 ;
        RECT 803.400 97.050 804.600 118.950 ;
        RECT 809.400 106.050 810.600 121.950 ;
        RECT 812.400 112.050 813.600 169.950 ;
        RECT 821.400 169.050 822.600 187.950 ;
        RECT 820.950 166.950 823.050 169.050 ;
        RECT 814.950 157.950 817.050 160.050 ;
        RECT 815.400 136.050 816.600 157.950 ;
        RECT 817.950 154.950 820.050 157.050 ;
        RECT 818.400 142.050 819.600 154.950 ;
        RECT 824.400 148.050 825.600 205.950 ;
        RECT 826.950 181.950 829.050 184.050 ;
        RECT 827.400 166.050 828.600 181.950 ;
        RECT 830.400 172.050 831.600 226.950 ;
        RECT 835.950 223.950 838.050 226.050 ;
        RECT 832.950 214.950 835.050 217.050 ;
        RECT 833.400 205.050 834.600 214.950 ;
        RECT 832.950 202.950 835.050 205.050 ;
        RECT 833.400 175.050 834.600 202.950 ;
        RECT 836.400 178.050 837.600 223.950 ;
        RECT 839.400 181.050 840.600 232.950 ;
        RECT 842.400 232.050 843.600 238.950 ;
        RECT 841.950 229.950 844.050 232.050 ;
        RECT 845.400 223.050 846.600 241.950 ;
        RECT 848.400 229.050 849.600 295.950 ;
        RECT 853.950 292.950 856.050 295.050 ;
        RECT 850.950 262.950 853.050 265.050 ;
        RECT 851.400 253.050 852.600 262.950 ;
        RECT 854.400 262.200 855.600 292.950 ;
        RECT 853.950 260.100 856.050 262.200 ;
        RECT 853.950 256.800 856.050 258.900 ;
        RECT 850.950 250.950 853.050 253.050 ;
        RECT 850.950 244.950 853.050 247.050 ;
        RECT 847.950 226.950 850.050 229.050 ;
        RECT 844.950 220.950 847.050 223.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 838.950 178.950 841.050 181.050 ;
        RECT 835.950 175.950 838.050 178.050 ;
        RECT 832.950 172.950 835.050 175.050 ;
        RECT 829.950 169.950 832.050 172.050 ;
        RECT 835.950 169.950 838.050 172.050 ;
        RECT 826.950 163.950 829.050 166.050 ;
        RECT 832.950 151.950 835.050 154.050 ;
        RECT 823.950 145.950 826.050 148.050 ;
        RECT 829.950 145.950 832.050 148.050 ;
        RECT 818.400 140.400 823.050 142.050 ;
        RECT 819.000 139.950 823.050 140.400 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 830.400 133.050 831.600 145.950 ;
        RECT 833.400 142.050 834.600 151.950 ;
        RECT 832.950 139.950 835.050 142.050 ;
        RECT 820.950 130.950 823.050 133.050 ;
        RECT 829.950 130.950 832.050 133.050 ;
        RECT 814.950 127.950 817.050 130.050 ;
        RECT 815.400 124.050 816.600 127.950 ;
        RECT 821.400 127.050 822.600 130.950 ;
        RECT 820.950 126.600 825.000 127.050 ;
        RECT 820.950 124.950 825.600 126.600 ;
        RECT 815.100 121.950 817.200 124.050 ;
        RECT 811.950 109.950 814.050 112.050 ;
        RECT 808.950 103.950 811.050 106.050 ;
        RECT 815.400 100.050 816.600 121.950 ;
        RECT 824.400 121.050 825.600 124.950 ;
        RECT 830.400 124.050 831.600 130.950 ;
        RECT 830.100 121.950 832.200 124.050 ;
        RECT 823.950 118.950 826.050 121.050 ;
        RECT 832.950 100.950 835.050 103.050 ;
        RECT 808.950 97.950 811.050 100.050 ;
        RECT 815.400 98.400 819.900 100.050 ;
        RECT 816.000 97.950 819.900 98.400 ;
        RECT 821.100 97.950 823.200 100.050 ;
        RECT 803.400 95.400 808.050 97.050 ;
        RECT 804.000 94.950 808.050 95.400 ;
        RECT 805.950 82.950 808.050 85.050 ;
        RECT 802.950 76.950 805.050 79.050 ;
        RECT 803.400 28.050 804.600 76.950 ;
        RECT 806.400 34.050 807.600 82.950 ;
        RECT 809.400 58.050 810.600 97.950 ;
        RECT 821.400 70.050 822.600 97.950 ;
        RECT 829.950 88.950 832.050 91.050 ;
        RECT 830.400 76.050 831.600 88.950 ;
        RECT 829.950 73.950 832.050 76.050 ;
        RECT 820.950 67.950 823.050 70.050 ;
        RECT 811.950 64.950 814.050 67.050 ;
        RECT 808.950 55.950 811.050 58.050 ;
        RECT 808.950 46.950 811.050 49.050 ;
        RECT 809.400 37.050 810.600 46.950 ;
        RECT 808.950 34.950 811.050 37.050 ;
        RECT 805.950 31.950 808.050 34.050 ;
        RECT 812.400 31.050 813.600 64.950 ;
        RECT 830.400 58.050 831.600 73.950 ;
        RECT 814.950 54.600 817.050 58.050 ;
        RECT 829.950 55.950 832.050 58.050 ;
        RECT 814.950 54.000 819.600 54.600 ;
        RECT 815.400 53.400 819.600 54.000 ;
        RECT 814.950 46.950 817.050 49.050 ;
        RECT 811.950 28.950 814.050 31.050 ;
        RECT 802.950 25.950 805.050 28.050 ;
        RECT 799.950 19.950 802.050 22.050 ;
        RECT 793.950 13.950 796.050 19.050 ;
        RECT 784.950 10.950 787.050 13.050 ;
        RECT 766.950 4.950 769.050 7.050 ;
        RECT 772.950 3.600 775.050 7.050 ;
        RECT 815.400 4.050 816.600 46.950 ;
        RECT 818.400 46.050 819.600 53.400 ;
        RECT 817.950 43.950 820.050 46.050 ;
        RECT 817.950 34.950 820.050 37.050 ;
        RECT 818.400 19.050 819.600 34.950 ;
        RECT 833.400 34.050 834.600 100.950 ;
        RECT 832.950 31.950 835.050 34.050 ;
        RECT 836.400 30.600 837.600 169.950 ;
        RECT 842.400 169.050 843.600 211.950 ;
        RECT 847.950 190.950 850.050 193.050 ;
        RECT 844.950 184.950 847.050 187.050 ;
        RECT 841.950 166.950 844.050 169.050 ;
        RECT 838.950 160.950 841.050 163.050 ;
        RECT 839.400 151.200 840.600 160.950 ;
        RECT 838.950 149.100 841.050 151.200 ;
        RECT 838.950 145.800 841.050 147.900 ;
        RECT 839.400 130.050 840.600 145.800 ;
        RECT 845.400 144.600 846.600 184.950 ;
        RECT 848.400 178.050 849.600 190.950 ;
        RECT 851.400 187.050 852.600 244.950 ;
        RECT 854.400 235.050 855.600 256.800 ;
        RECT 856.950 250.950 859.050 253.050 ;
        RECT 857.400 244.050 858.600 250.950 ;
        RECT 856.950 241.950 859.050 244.050 ;
        RECT 853.950 232.950 856.050 235.050 ;
        RECT 853.950 220.950 856.050 223.050 ;
        RECT 850.950 184.950 853.050 187.050 ;
        RECT 854.400 183.600 855.600 220.950 ;
        RECT 856.950 208.950 859.050 211.050 ;
        RECT 851.400 182.400 855.600 183.600 ;
        RECT 847.950 175.950 850.050 178.050 ;
        RECT 845.400 143.400 849.600 144.600 ;
        RECT 844.950 139.950 847.050 142.050 ;
        RECT 838.950 127.950 841.050 130.050 ;
        RECT 845.400 124.050 846.600 139.950 ;
        RECT 844.800 121.950 846.900 124.050 ;
        RECT 841.950 112.950 844.050 115.050 ;
        RECT 838.950 55.950 841.050 58.050 ;
        RECT 839.400 46.200 840.600 55.950 ;
        RECT 838.950 44.100 841.050 46.200 ;
        RECT 838.950 40.800 841.050 42.900 ;
        RECT 839.400 31.050 840.600 40.800 ;
        RECT 833.400 29.400 837.600 30.600 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 817.950 16.950 820.050 19.050 ;
        RECT 827.400 13.050 828.600 22.950 ;
        RECT 833.400 22.050 834.600 29.400 ;
        RECT 838.950 28.950 841.050 31.050 ;
        RECT 832.950 19.950 835.050 22.050 ;
        RECT 842.400 16.050 843.600 112.950 ;
        RECT 848.400 109.050 849.600 143.400 ;
        RECT 851.400 129.600 852.600 182.400 ;
        RECT 853.950 178.950 856.050 181.050 ;
        RECT 854.400 139.050 855.600 178.950 ;
        RECT 853.950 136.950 856.050 139.050 ;
        RECT 851.400 128.400 855.600 129.600 ;
        RECT 850.950 124.950 853.050 127.050 ;
        RECT 847.950 106.950 850.050 109.050 ;
        RECT 851.400 85.050 852.600 124.950 ;
        RECT 850.950 82.950 853.050 85.050 ;
        RECT 844.950 61.950 847.050 64.050 ;
        RECT 845.400 55.050 846.600 61.950 ;
        RECT 850.950 58.950 853.050 61.050 ;
        RECT 844.950 52.950 847.050 55.050 ;
        RECT 851.400 49.050 852.600 58.950 ;
        RECT 850.950 46.950 853.050 49.050 ;
        RECT 841.950 13.950 844.050 16.050 ;
        RECT 826.950 10.950 829.050 13.050 ;
        RECT 854.400 7.050 855.600 128.400 ;
        RECT 857.400 40.050 858.600 208.950 ;
        RECT 856.950 37.950 859.050 40.050 ;
        RECT 853.950 4.950 856.050 7.050 ;
        RECT 761.400 3.000 775.050 3.600 ;
        RECT 761.400 2.400 774.600 3.000 ;
        RECT 814.950 1.950 817.050 4.050 ;
  END
END ALU_wrapper
END LIBRARY

