magic
tech scmos
magscale 1 30
timestamp 1727178187
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1555589239
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1555589239
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1555589239
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1555589239
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1555589239
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1555589239
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1555589239
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1555589239
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1555589239
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1555589239
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PIC  CIN_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_1
timestamp 1555589239
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_2
timestamp 1555589239
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_3
timestamp 1555589239
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_4
timestamp 1555589239
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  CIN_5
timestamp 1555589239
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use PIC  CLK
timestamp 1555589239
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use PIC  RDY_I
timestamp 1555589239
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use PIC  XIN_0
timestamp 1555589239
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC  XIN_1
timestamp 1555589239
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC  XIN_2
timestamp 1555589239
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  XIN_3
timestamp 1555589239
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC  YIN_0
timestamp 1555589239
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PIC  YIN_1
timestamp 1555589239
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_2
timestamp 1555589239
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN_3
timestamp 1555589239
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use POB8  VLD_O ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use POB8  XOUT_0
timestamp 1555589239
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use POB8  XOUT_1
timestamp 1555589239
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use POB8  XOUT_2
timestamp 1555589239
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use POB8  XOUT_3
timestamp 1555589239
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use POB8  YOUT_0
timestamp 1555589239
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_1
timestamp 1555589239
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_2
timestamp 1555589239
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use POB8  YOUT_3
timestamp 1555589239
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use PVSS  VSS_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use PVDD  VDD_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use PVDD  VDD_1
timestamp 1555589239
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use MY_LOGO  MY_LOGO_0
timestamp 1724157349
transform 1 0 149420 0 1 9675
box 180 225 21510 9045
<< end >>