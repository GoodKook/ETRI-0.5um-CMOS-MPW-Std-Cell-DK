VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fir_pe
  CLASS BLOCK ;
  FOREIGN fir_pe ;
  ORIGIN 6.000 6.000 ;
  SIZE 876.000 BY 834.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 819.300 873.450 821.700 ;
        RECT 864.450 743.700 873.450 819.300 ;
        RECT 0.600 741.300 873.450 743.700 ;
        RECT 658.800 735.300 660.600 741.300 ;
        RECT 667.800 735.300 669.600 741.300 ;
        RECT 626.400 665.700 628.200 671.700 ;
        RECT 635.100 665.700 636.900 671.700 ;
        RECT 674.400 665.700 676.200 671.700 ;
        RECT 683.400 665.700 685.200 671.700 ;
        RECT 864.450 665.700 873.450 741.300 ;
        RECT 0.600 663.300 873.450 665.700 ;
        RECT 864.450 587.700 873.450 663.300 ;
        RECT 0.600 585.300 873.450 587.700 ;
        RECT 743.400 509.700 745.200 515.700 ;
        RECT 752.400 509.700 754.200 515.700 ;
        RECT 818.400 509.700 820.200 515.700 ;
        RECT 827.400 509.700 829.200 515.700 ;
        RECT 864.450 509.700 873.450 585.300 ;
        RECT 0.600 507.300 873.450 509.700 ;
        RECT 218.100 501.300 219.900 507.300 ;
        RECT 226.800 501.300 228.600 507.300 ;
        RECT 671.400 501.300 673.200 507.300 ;
        RECT 680.100 501.300 681.900 507.300 ;
        RECT 755.400 501.300 757.200 507.300 ;
        RECT 764.400 501.300 766.200 507.300 ;
        RECT 155.400 431.700 157.200 437.700 ;
        RECT 164.100 431.700 165.900 437.700 ;
        RECT 260.400 431.700 262.200 437.700 ;
        RECT 269.400 431.700 271.200 437.700 ;
        RECT 835.800 431.700 837.600 437.700 ;
        RECT 844.800 431.700 846.600 437.700 ;
        RECT 864.450 431.700 873.450 507.300 ;
        RECT 0.600 429.300 873.450 431.700 ;
        RECT 152.100 353.700 153.900 359.700 ;
        RECT 160.800 353.700 162.600 359.700 ;
        RECT 864.450 353.700 873.450 429.300 ;
        RECT 0.600 351.300 873.450 353.700 ;
        RECT 236.400 275.700 238.200 281.700 ;
        RECT 245.400 275.700 247.200 281.700 ;
        RECT 676.800 275.700 678.600 281.700 ;
        RECT 685.800 275.700 687.600 281.700 ;
        RECT 864.450 275.700 873.450 351.300 ;
        RECT 0.600 273.300 873.450 275.700 ;
        RECT 269.100 197.700 270.900 203.700 ;
        RECT 277.800 197.700 279.600 203.700 ;
        RECT 722.400 197.700 724.200 203.700 ;
        RECT 731.400 197.700 733.200 203.700 ;
        RECT 864.450 197.700 873.450 273.300 ;
        RECT 0.600 195.300 873.450 197.700 ;
        RECT 101.400 119.700 103.200 125.700 ;
        RECT 110.400 119.700 112.200 125.700 ;
        RECT 864.450 119.700 873.450 195.300 ;
        RECT 0.600 117.300 873.450 119.700 ;
        RECT 13.800 111.300 15.600 117.300 ;
        RECT 22.800 111.300 24.600 117.300 ;
        RECT 95.100 111.300 96.900 117.300 ;
        RECT 103.800 111.300 105.600 117.300 ;
        RECT 864.450 41.700 873.450 117.300 ;
        RECT 0.600 39.300 873.450 41.700 ;
        RECT 864.450 0.300 873.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 782.700 -0.450 821.700 ;
        RECT -9.450 780.300 863.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT 658.800 704.700 660.600 715.500 ;
        RECT 667.800 704.700 669.600 715.500 ;
        RECT -9.450 702.300 863.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT 626.400 691.500 628.200 702.300 ;
        RECT 635.100 691.500 637.200 702.300 ;
        RECT 674.400 691.500 676.200 702.300 ;
        RECT 683.400 691.500 685.200 702.300 ;
        RECT -9.450 624.300 863.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT -9.450 546.300 863.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT 743.400 535.500 745.200 546.300 ;
        RECT 752.400 535.500 754.200 546.300 ;
        RECT 818.400 535.500 820.200 546.300 ;
        RECT 827.400 535.500 829.200 546.300 ;
        RECT 217.800 470.700 219.900 481.500 ;
        RECT 226.800 470.700 228.600 481.500 ;
        RECT 671.400 470.700 673.200 481.500 ;
        RECT 680.100 470.700 682.200 481.500 ;
        RECT 755.400 470.700 757.200 481.500 ;
        RECT 764.400 470.700 766.200 481.500 ;
        RECT -9.450 468.300 863.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT 155.400 457.500 157.200 468.300 ;
        RECT 164.100 457.500 166.200 468.300 ;
        RECT 260.400 457.500 262.200 468.300 ;
        RECT 269.400 457.500 271.200 468.300 ;
        RECT 835.800 457.500 837.600 468.300 ;
        RECT 844.800 457.500 846.600 468.300 ;
        RECT -9.450 390.300 863.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT 151.800 379.500 153.900 390.300 ;
        RECT 160.800 379.500 162.600 390.300 ;
        RECT -9.450 312.300 863.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT 236.400 301.500 238.200 312.300 ;
        RECT 245.400 301.500 247.200 312.300 ;
        RECT 676.800 301.500 678.600 312.300 ;
        RECT 685.800 301.500 687.600 312.300 ;
        RECT -9.450 234.300 863.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT 268.800 223.500 270.900 234.300 ;
        RECT 277.800 223.500 279.600 234.300 ;
        RECT 722.400 223.500 724.200 234.300 ;
        RECT 731.400 223.500 733.200 234.300 ;
        RECT -9.450 156.300 863.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT 101.400 145.500 103.200 156.300 ;
        RECT 110.400 145.500 112.200 156.300 ;
        RECT 13.800 80.700 15.600 91.500 ;
        RECT 22.800 80.700 24.600 91.500 ;
        RECT 94.800 80.700 96.900 91.500 ;
        RECT 103.800 80.700 105.600 91.500 ;
        RECT -9.450 78.300 863.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT -9.450 0.300 863.400 2.700 ;
    END
  END vdd
  PIN Cin[5]
    PORT
      LAYER metal1 ;
        RECT 508.950 651.450 513.000 652.050 ;
        RECT 508.950 649.950 513.450 651.450 ;
        RECT 512.550 642.900 513.450 649.950 ;
        RECT 511.950 640.800 514.050 642.900 ;
      LAYER metal2 ;
        RECT 581.400 814.050 582.450 828.450 ;
        RECT 568.950 811.950 571.050 814.050 ;
        RECT 580.950 811.950 583.050 814.050 ;
        RECT 569.400 801.450 570.450 811.950 ;
        RECT 569.400 800.400 573.450 801.450 ;
        RECT 572.400 754.050 573.450 800.400 ;
        RECT 541.950 751.950 544.050 754.050 ;
        RECT 571.950 751.950 574.050 754.050 ;
        RECT 542.400 739.050 543.450 751.950 ;
        RECT 526.950 736.950 529.050 739.050 ;
        RECT 541.950 736.950 544.050 739.050 ;
        RECT 527.400 730.050 528.450 736.950 ;
        RECT 526.950 727.950 529.050 730.050 ;
        RECT 523.950 721.950 526.050 724.050 ;
        RECT 524.400 688.050 525.450 721.950 ;
        RECT 523.950 685.950 526.050 688.050 ;
        RECT 508.950 676.950 511.050 679.050 ;
        RECT 509.400 652.050 510.450 676.950 ;
        RECT 508.950 649.950 511.050 652.050 ;
        RECT 461.400 644.400 462.600 646.800 ;
        RECT 461.400 625.050 462.450 644.400 ;
        RECT 511.950 640.800 514.050 642.900 ;
        RECT 512.400 625.050 513.450 640.800 ;
        RECT 461.400 622.950 466.050 625.050 ;
        RECT 511.950 622.950 514.050 625.050 ;
        RECT 461.400 610.200 462.450 622.950 ;
        RECT 541.950 622.800 544.050 624.900 ;
        RECT 419.400 606.450 420.600 606.600 ;
        RECT 421.950 606.450 424.050 610.050 ;
        RECT 448.950 607.950 451.050 610.050 ;
        RECT 460.950 608.100 463.050 610.200 ;
        RECT 542.400 610.050 543.450 622.800 ;
        RECT 541.950 607.950 544.050 610.050 ;
        RECT 419.400 606.000 424.050 606.450 ;
        RECT 419.400 605.400 423.450 606.000 ;
        RECT 419.400 604.200 420.600 605.400 ;
        RECT 449.400 573.450 450.450 607.950 ;
        RECT 568.950 604.800 571.050 606.900 ;
        RECT 569.400 604.200 570.600 604.800 ;
        RECT 449.400 572.400 453.450 573.450 ;
        RECT 407.400 567.000 408.600 568.800 ;
        RECT 406.950 562.950 409.050 567.000 ;
        RECT 430.950 562.950 433.050 565.050 ;
        RECT 431.400 559.050 432.450 562.950 ;
        RECT 452.400 559.050 453.450 572.400 ;
        RECT 430.950 556.950 433.050 559.050 ;
        RECT 451.800 556.950 453.900 559.050 ;
      LAYER metal3 ;
        RECT 568.950 813.600 571.050 814.050 ;
        RECT 580.950 813.600 583.050 814.050 ;
        RECT 568.950 812.400 583.050 813.600 ;
        RECT 568.950 811.950 571.050 812.400 ;
        RECT 580.950 811.950 583.050 812.400 ;
        RECT 541.950 753.600 544.050 754.050 ;
        RECT 571.950 753.600 574.050 754.050 ;
        RECT 541.950 752.400 574.050 753.600 ;
        RECT 541.950 751.950 544.050 752.400 ;
        RECT 571.950 751.950 574.050 752.400 ;
        RECT 526.950 738.600 529.050 739.050 ;
        RECT 541.950 738.600 544.050 739.050 ;
        RECT 526.950 737.400 544.050 738.600 ;
        RECT 526.950 736.950 529.050 737.400 ;
        RECT 541.950 736.950 544.050 737.400 ;
        RECT 526.950 727.950 529.050 730.050 ;
        RECT 527.400 724.050 528.600 727.950 ;
        RECT 523.950 722.400 528.600 724.050 ;
        RECT 523.950 721.950 528.000 722.400 ;
        RECT 523.950 687.600 526.050 688.050 ;
        RECT 509.400 686.400 526.050 687.600 ;
        RECT 509.400 679.050 510.600 686.400 ;
        RECT 523.950 685.950 526.050 686.400 ;
        RECT 508.950 676.950 511.050 679.050 ;
        RECT 463.950 624.600 466.050 625.050 ;
        RECT 511.950 624.600 514.050 625.050 ;
        RECT 541.950 624.600 544.050 624.900 ;
        RECT 463.950 623.400 544.050 624.600 ;
        RECT 463.950 622.950 466.050 623.400 ;
        RECT 511.950 622.950 514.050 623.400 ;
        RECT 541.950 622.800 544.050 623.400 ;
        RECT 421.950 609.600 424.050 610.050 ;
        RECT 448.950 609.600 451.050 610.050 ;
        RECT 460.950 609.600 463.050 610.200 ;
        RECT 421.950 608.400 463.050 609.600 ;
        RECT 421.950 607.950 424.050 608.400 ;
        RECT 448.950 607.950 451.050 608.400 ;
        RECT 460.950 608.100 463.050 608.400 ;
        RECT 541.950 609.600 544.050 610.050 ;
        RECT 541.950 608.400 564.600 609.600 ;
        RECT 541.950 607.950 544.050 608.400 ;
        RECT 563.400 606.600 564.600 608.400 ;
        RECT 568.950 606.600 571.050 606.900 ;
        RECT 563.400 605.400 571.050 606.600 ;
        RECT 568.950 604.800 571.050 605.400 ;
        RECT 406.950 564.600 409.050 565.050 ;
        RECT 430.950 564.600 433.050 565.050 ;
        RECT 406.950 563.400 433.050 564.600 ;
        RECT 406.950 562.950 409.050 563.400 ;
        RECT 430.950 562.950 433.050 563.400 ;
        RECT 430.950 558.600 433.050 559.050 ;
        RECT 451.800 558.600 453.900 559.050 ;
        RECT 430.950 557.400 453.900 558.600 ;
        RECT 430.950 556.950 433.050 557.400 ;
        RECT 451.800 556.950 453.900 557.400 ;
    END
  END Cin[5]
  PIN Cin[4]
    PORT
      LAYER metal1 ;
        RECT 646.950 762.450 651.000 763.050 ;
        RECT 646.950 760.950 651.450 762.450 ;
        RECT 643.950 753.450 646.050 754.050 ;
        RECT 650.550 753.450 651.450 760.950 ;
        RECT 643.950 752.550 651.450 753.450 ;
        RECT 643.950 751.950 646.050 752.550 ;
        RECT 432.000 651.450 436.050 652.050 ;
        RECT 431.550 649.950 436.050 651.450 ;
        RECT 431.550 646.050 432.450 649.950 ;
        RECT 431.550 644.550 436.050 646.050 ;
        RECT 432.000 643.950 436.050 644.550 ;
        RECT 298.950 606.450 303.000 607.050 ;
        RECT 601.950 606.450 604.050 607.050 ;
        RECT 298.950 604.950 303.450 606.450 ;
        RECT 302.550 601.050 303.450 604.950 ;
        RECT 298.950 599.550 303.450 601.050 ;
        RECT 596.550 605.550 604.050 606.450 ;
        RECT 596.550 601.050 597.450 605.550 ;
        RECT 601.950 604.950 604.050 605.550 ;
        RECT 596.550 599.550 601.050 601.050 ;
        RECT 298.950 598.950 303.000 599.550 ;
        RECT 597.000 598.950 601.050 599.550 ;
        RECT 598.950 574.950 601.050 577.050 ;
        RECT 282.000 573.450 286.050 574.050 ;
        RECT 281.550 571.950 286.050 573.450 ;
        RECT 281.550 568.050 282.450 571.950 ;
        RECT 281.550 566.550 286.050 568.050 ;
        RECT 282.000 565.950 286.050 566.550 ;
        RECT 592.950 567.450 595.050 568.050 ;
        RECT 599.550 567.450 600.450 574.950 ;
        RECT 592.950 566.550 600.450 567.450 ;
        RECT 592.950 565.950 595.050 566.550 ;
      LAYER metal2 ;
        RECT 575.400 820.050 576.450 828.450 ;
        RECT 584.400 824.400 627.450 825.450 ;
        RECT 584.400 820.050 585.450 824.400 ;
        RECT 574.950 817.950 577.050 820.050 ;
        RECT 583.950 817.950 586.050 820.050 ;
        RECT 626.400 808.050 627.450 824.400 ;
        RECT 625.950 805.950 628.050 808.050 ;
        RECT 634.950 799.950 637.050 802.050 ;
        RECT 635.400 795.450 636.450 799.950 ;
        RECT 635.400 794.400 639.450 795.450 ;
        RECT 638.400 772.050 639.450 794.400 ;
        RECT 637.950 769.950 640.050 772.050 ;
        RECT 646.950 769.950 649.050 772.050 ;
        RECT 647.400 763.050 648.450 769.950 ;
        RECT 646.950 760.950 649.050 763.050 ;
        RECT 643.950 751.950 646.050 754.050 ;
        RECT 644.400 730.050 645.450 751.950 ;
        RECT 643.950 727.950 646.050 730.050 ;
        RECT 643.950 721.950 646.050 724.050 ;
        RECT 644.400 670.050 645.450 721.950 ;
        RECT 559.950 667.950 562.050 670.050 ;
        RECT 277.950 650.250 280.050 652.350 ;
        RECT 286.950 650.250 289.050 652.350 ;
        RECT 278.400 649.500 279.600 650.250 ;
        RECT 287.400 646.050 288.450 650.250 ;
        RECT 433.950 649.950 436.050 655.050 ;
        RECT 442.950 650.250 445.050 652.350 ;
        RECT 560.400 651.600 561.450 667.950 ;
        RECT 587.400 667.050 588.450 669.450 ;
        RECT 643.950 667.950 646.050 670.050 ;
        RECT 586.950 664.950 589.050 667.050 ;
        RECT 595.950 664.950 598.050 667.050 ;
        RECT 587.400 651.600 588.450 664.950 ;
        RECT 443.400 649.500 444.600 650.250 ;
        RECT 560.400 649.500 561.600 651.600 ;
        RECT 587.400 649.500 588.600 651.600 ;
        RECT 296.400 646.050 297.600 646.800 ;
        RECT 286.950 643.950 289.050 646.050 ;
        RECT 295.950 643.950 298.050 646.050 ;
        RECT 433.950 643.950 436.050 646.050 ;
        RECT 296.400 610.050 297.450 643.950 ;
        RECT 434.400 640.050 435.450 643.950 ;
        RECT 596.400 643.050 597.450 664.950 ;
        RECT 595.950 640.950 598.050 643.050 ;
        RECT 601.950 640.800 604.050 642.900 ;
        RECT 322.950 637.950 325.050 640.050 ;
        RECT 433.950 637.950 436.050 640.050 ;
        RECT 323.400 621.450 324.450 637.950 ;
        RECT 320.400 620.400 324.450 621.450 ;
        RECT 320.400 610.050 321.450 620.400 ;
        RECT 295.950 609.450 298.050 610.050 ;
        RECT 295.950 609.000 300.450 609.450 ;
        RECT 295.950 608.400 301.050 609.000 ;
        RECT 295.950 607.950 298.050 608.400 ;
        RECT 298.950 604.950 301.050 608.400 ;
        RECT 319.800 607.950 321.900 610.050 ;
        RECT 602.400 607.050 603.450 640.800 ;
        RECT 601.950 604.950 604.050 607.050 ;
        RECT 602.400 604.200 603.600 604.950 ;
        RECT 298.950 598.950 301.050 601.050 ;
        RECT 598.950 598.950 601.050 601.050 ;
        RECT 299.400 580.050 300.450 598.950 ;
        RECT 289.950 577.950 292.050 580.050 ;
        RECT 298.950 577.950 301.050 580.050 ;
        RECT 283.950 571.950 286.050 577.050 ;
        RECT 290.400 574.350 291.450 577.950 ;
        RECT 599.400 577.050 600.450 598.950 ;
        RECT 598.950 574.950 601.050 577.050 ;
        RECT 289.950 572.250 292.050 574.350 ;
        RECT 290.400 571.500 291.600 572.250 ;
        RECT 521.400 568.050 522.600 568.800 ;
        RECT 593.400 568.050 594.600 568.800 ;
        RECT 283.950 565.950 286.050 568.050 ;
        RECT 508.950 565.950 511.050 568.050 ;
        RECT 520.950 565.950 523.050 568.050 ;
        RECT 592.950 565.950 595.050 568.050 ;
        RECT 284.400 541.050 285.450 565.950 ;
        RECT 509.400 553.050 510.450 565.950 ;
        RECT 430.950 550.950 433.050 553.050 ;
        RECT 508.950 550.950 511.050 553.050 ;
        RECT 532.950 550.950 535.050 553.050 ;
        RECT 431.400 547.050 432.450 550.950 ;
        RECT 533.400 547.050 534.450 550.950 ;
        RECT 593.400 547.050 594.450 565.950 ;
        RECT 430.950 544.950 433.050 547.050 ;
        RECT 532.950 544.950 535.050 547.050 ;
        RECT 592.950 544.950 595.050 547.050 ;
        RECT 394.950 541.950 397.050 544.050 ;
        RECT 283.950 538.950 286.050 541.050 ;
        RECT 355.950 538.950 358.050 541.050 ;
        RECT 356.400 528.600 357.450 538.950 ;
        RECT 395.400 535.050 396.450 541.950 ;
        RECT 406.950 541.800 409.050 543.900 ;
        RECT 407.400 535.050 408.450 541.800 ;
        RECT 394.950 532.950 397.050 535.050 ;
        RECT 406.950 532.950 409.050 535.050 ;
        RECT 593.400 532.050 594.450 544.950 ;
        RECT 592.950 529.950 595.050 532.050 ;
        RECT 356.400 526.200 357.600 528.600 ;
        RECT 604.950 528.000 607.050 532.050 ;
        RECT 605.400 526.200 606.600 528.000 ;
      LAYER metal3 ;
        RECT 574.950 819.600 577.050 820.050 ;
        RECT 583.950 819.600 586.050 820.050 ;
        RECT 574.950 818.400 586.050 819.600 ;
        RECT 574.950 817.950 577.050 818.400 ;
        RECT 583.950 817.950 586.050 818.400 ;
        RECT 625.950 807.600 630.000 808.050 ;
        RECT 625.950 805.950 630.600 807.600 ;
        RECT 629.400 804.600 630.600 805.950 ;
        RECT 629.400 803.400 633.600 804.600 ;
        RECT 632.400 802.050 633.600 803.400 ;
        RECT 632.400 800.400 637.050 802.050 ;
        RECT 633.000 799.950 637.050 800.400 ;
        RECT 637.950 771.600 640.050 772.050 ;
        RECT 646.950 771.600 649.050 772.050 ;
        RECT 637.950 770.400 649.050 771.600 ;
        RECT 637.950 769.950 640.050 770.400 ;
        RECT 646.950 769.950 649.050 770.400 ;
        RECT 643.950 727.950 646.050 730.050 ;
        RECT 644.400 724.050 645.600 727.950 ;
        RECT 643.950 721.950 646.050 724.050 ;
        RECT 559.950 669.600 562.050 670.050 ;
        RECT 643.950 669.600 646.050 670.050 ;
        RECT 559.950 668.400 646.050 669.600 ;
        RECT 559.950 667.950 562.050 668.400 ;
        RECT 587.400 667.050 588.600 668.400 ;
        RECT 643.950 667.950 646.050 668.400 ;
        RECT 586.950 666.600 589.050 667.050 ;
        RECT 595.950 666.600 598.050 667.050 ;
        RECT 586.950 665.400 598.050 666.600 ;
        RECT 586.950 664.950 589.050 665.400 ;
        RECT 595.950 664.950 598.050 665.400 ;
        RECT 277.950 651.900 280.050 652.350 ;
        RECT 286.950 651.900 289.050 652.350 ;
        RECT 277.950 650.700 289.050 651.900 ;
        RECT 433.950 651.600 436.050 655.050 ;
        RECT 442.950 651.600 445.050 652.350 ;
        RECT 433.950 651.000 445.050 651.600 ;
        RECT 277.950 650.250 280.050 650.700 ;
        RECT 286.950 650.250 289.050 650.700 ;
        RECT 434.400 650.400 445.050 651.000 ;
        RECT 442.950 650.250 445.050 650.400 ;
        RECT 286.950 645.600 289.050 646.050 ;
        RECT 295.950 645.600 298.050 646.050 ;
        RECT 286.950 644.400 298.050 645.600 ;
        RECT 286.950 643.950 289.050 644.400 ;
        RECT 295.950 643.950 298.050 644.400 ;
        RECT 595.950 642.600 598.050 643.050 ;
        RECT 601.950 642.600 604.050 642.900 ;
        RECT 595.950 641.400 604.050 642.600 ;
        RECT 595.950 640.950 598.050 641.400 ;
        RECT 601.950 640.800 604.050 641.400 ;
        RECT 322.950 639.600 325.050 640.050 ;
        RECT 433.950 639.600 436.050 640.050 ;
        RECT 322.950 638.400 396.600 639.600 ;
        RECT 322.950 637.950 325.050 638.400 ;
        RECT 395.400 636.600 396.600 638.400 ;
        RECT 407.400 638.400 436.050 639.600 ;
        RECT 407.400 636.600 408.600 638.400 ;
        RECT 433.950 637.950 436.050 638.400 ;
        RECT 395.400 635.400 408.600 636.600 ;
        RECT 295.950 609.600 298.050 610.050 ;
        RECT 319.800 609.600 321.900 610.050 ;
        RECT 295.950 608.400 321.900 609.600 ;
        RECT 295.950 607.950 298.050 608.400 ;
        RECT 319.800 607.950 321.900 608.400 ;
        RECT 289.950 579.600 292.050 580.050 ;
        RECT 298.950 579.600 301.050 580.050 ;
        RECT 289.950 578.400 301.050 579.600 ;
        RECT 289.950 577.950 292.050 578.400 ;
        RECT 298.950 577.950 301.050 578.400 ;
        RECT 283.950 573.600 286.050 577.050 ;
        RECT 289.950 573.600 292.050 574.350 ;
        RECT 283.950 573.000 292.050 573.600 ;
        RECT 284.400 572.400 292.050 573.000 ;
        RECT 289.950 572.250 292.050 572.400 ;
        RECT 508.950 567.600 511.050 568.050 ;
        RECT 520.950 567.600 523.050 568.050 ;
        RECT 508.950 566.400 523.050 567.600 ;
        RECT 508.950 565.950 511.050 566.400 ;
        RECT 520.950 565.950 523.050 566.400 ;
        RECT 430.950 552.600 433.050 553.050 ;
        RECT 508.950 552.600 511.050 553.050 ;
        RECT 532.950 552.600 535.050 553.050 ;
        RECT 430.950 551.400 535.050 552.600 ;
        RECT 430.950 550.950 433.050 551.400 ;
        RECT 508.950 550.950 511.050 551.400 ;
        RECT 532.950 550.950 535.050 551.400 ;
        RECT 430.950 546.600 433.050 547.050 ;
        RECT 425.400 545.400 433.050 546.600 ;
        RECT 393.000 543.600 397.050 544.050 ;
        RECT 356.400 542.400 366.600 543.600 ;
        RECT 356.400 541.050 357.600 542.400 ;
        RECT 283.950 540.600 286.050 541.050 ;
        RECT 355.950 540.600 358.050 541.050 ;
        RECT 283.950 539.400 358.050 540.600 ;
        RECT 365.400 540.600 366.600 542.400 ;
        RECT 392.400 541.950 397.050 543.600 ;
        RECT 406.950 543.600 409.050 543.900 ;
        RECT 425.400 543.600 426.600 545.400 ;
        RECT 430.950 544.950 433.050 545.400 ;
        RECT 532.950 546.600 535.050 547.050 ;
        RECT 592.950 546.600 595.050 547.050 ;
        RECT 532.950 545.400 595.050 546.600 ;
        RECT 532.950 544.950 535.050 545.400 ;
        RECT 592.950 544.950 595.050 545.400 ;
        RECT 406.950 542.400 426.600 543.600 ;
        RECT 392.400 540.600 393.600 541.950 ;
        RECT 406.950 541.800 409.050 542.400 ;
        RECT 365.400 539.400 393.600 540.600 ;
        RECT 283.950 538.950 286.050 539.400 ;
        RECT 355.950 538.950 358.050 539.400 ;
        RECT 394.950 534.600 397.050 535.050 ;
        RECT 406.950 534.600 409.050 535.050 ;
        RECT 394.950 533.400 409.050 534.600 ;
        RECT 394.950 532.950 397.050 533.400 ;
        RECT 406.950 532.950 409.050 533.400 ;
        RECT 592.950 531.600 595.050 532.050 ;
        RECT 604.950 531.600 607.050 532.050 ;
        RECT 592.950 530.400 607.050 531.600 ;
        RECT 592.950 529.950 595.050 530.400 ;
        RECT 604.950 529.950 607.050 530.400 ;
    END
  END Cin[4]
  PIN Cin[3]
    PORT
      LAYER metal1 ;
        RECT 559.950 573.450 564.000 574.050 ;
        RECT 559.950 571.950 564.450 573.450 ;
        RECT 556.950 567.450 559.050 568.050 ;
        RECT 563.550 567.450 564.450 571.950 ;
        RECT 556.950 566.550 564.450 567.450 ;
        RECT 556.950 565.950 559.050 566.550 ;
        RECT 301.950 528.450 304.050 529.050 ;
        RECT 310.950 528.450 313.050 529.050 ;
        RECT 301.950 527.550 313.050 528.450 ;
        RECT 301.950 526.950 304.050 527.550 ;
        RECT 310.950 526.950 313.050 527.550 ;
      LAYER metal2 ;
        RECT 569.400 823.050 570.450 828.450 ;
        RECT 568.950 820.950 571.050 823.050 ;
        RECT 586.950 820.950 589.050 823.050 ;
        RECT 587.400 811.050 588.450 820.950 ;
        RECT 586.950 808.950 589.050 811.050 ;
        RECT 607.950 808.950 610.050 811.050 ;
        RECT 608.400 790.050 609.450 808.950 ;
        RECT 607.950 787.950 610.050 790.050 ;
        RECT 628.950 787.800 631.050 789.900 ;
        RECT 629.400 742.050 630.450 787.800 ;
        RECT 628.950 739.950 631.050 742.050 ;
        RECT 646.950 739.950 649.050 742.050 ;
        RECT 647.400 715.050 648.450 739.950 ;
        RECT 580.950 712.950 583.050 715.050 ;
        RECT 646.950 712.950 649.050 715.050 ;
        RECT 581.400 673.050 582.450 712.950 ;
        RECT 562.950 670.950 565.050 673.050 ;
        RECT 580.950 670.950 583.050 673.050 ;
        RECT 563.400 661.050 564.450 670.950 ;
        RECT 541.950 658.950 544.050 661.050 ;
        RECT 553.950 658.950 556.050 661.050 ;
        RECT 562.950 658.950 565.050 661.050 ;
        RECT 542.400 651.600 543.450 658.950 ;
        RECT 554.400 652.050 555.450 658.950 ;
        RECT 563.400 654.450 564.450 658.950 ;
        RECT 563.400 653.400 567.450 654.450 ;
        RECT 542.400 649.500 543.600 651.600 ;
        RECT 553.950 649.950 556.050 652.050 ;
        RECT 566.400 651.600 567.450 653.400 ;
        RECT 566.400 649.500 567.600 651.600 ;
        RECT 457.950 643.950 460.050 646.050 ;
        RECT 484.800 643.950 486.900 646.050 ;
        RECT 547.950 643.950 550.050 646.050 ;
        RECT 458.400 637.050 459.450 643.950 ;
        RECT 485.400 637.050 486.450 643.950 ;
        RECT 548.400 637.050 549.450 643.950 ;
        RECT 583.950 640.950 586.050 643.050 ;
        RECT 424.950 634.950 427.050 637.050 ;
        RECT 457.950 634.950 460.050 637.050 ;
        RECT 484.950 634.950 487.050 637.050 ;
        RECT 547.950 634.950 550.050 637.050 ;
        RECT 425.400 600.750 426.450 634.950 ;
        RECT 548.400 607.050 549.450 634.950 ;
        RECT 584.400 619.050 585.450 640.950 ;
        RECT 583.950 616.950 586.050 619.050 ;
        RECT 610.950 616.950 613.050 619.050 ;
        RECT 547.950 604.950 550.050 607.050 ;
        RECT 584.400 606.600 585.450 616.950 ;
        RECT 611.400 610.050 612.450 616.950 ;
        RECT 610.950 607.950 613.050 610.050 ;
        RECT 584.400 604.200 585.600 606.600 ;
        RECT 622.950 606.000 625.050 610.050 ;
        RECT 623.400 604.200 624.600 606.000 ;
        RECT 437.400 600.750 438.600 601.500 ;
        RECT 424.950 598.650 427.050 600.750 ;
        RECT 436.950 598.650 439.050 600.750 ;
        RECT 559.950 598.950 562.050 601.050 ;
        RECT 425.400 586.050 426.450 598.650 ;
        RECT 361.950 583.950 364.050 586.050 ;
        RECT 424.950 583.950 427.050 586.050 ;
        RECT 310.950 572.250 313.050 574.350 ;
        RECT 311.400 571.500 312.600 572.250 ;
        RECT 310.950 565.950 313.050 568.050 ;
        RECT 311.400 532.050 312.450 565.950 ;
        RECT 362.400 552.450 363.450 583.950 ;
        RECT 560.400 574.050 561.450 598.950 ;
        RECT 559.950 571.950 562.050 574.050 ;
        RECT 557.400 568.050 558.600 568.800 ;
        RECT 556.950 565.950 559.050 568.050 ;
        RECT 557.400 553.050 558.450 565.950 ;
        RECT 586.950 556.950 589.050 559.050 ;
        RECT 628.800 556.950 630.900 559.050 ;
        RECT 587.400 553.050 588.450 556.950 ;
        RECT 359.400 551.400 363.450 552.450 ;
        RECT 301.950 526.950 304.050 529.050 ;
        RECT 310.950 526.950 313.050 532.050 ;
        RECT 359.400 529.050 360.450 551.400 ;
        RECT 556.950 550.950 559.050 553.050 ;
        RECT 586.950 550.950 589.050 553.050 ;
        RECT 629.400 544.050 630.450 556.950 ;
        RECT 628.950 541.950 631.050 544.050 ;
        RECT 661.950 541.950 664.050 544.050 ;
        RECT 337.950 526.950 340.050 529.050 ;
        RECT 358.950 526.950 361.050 529.050 ;
        RECT 662.400 528.600 663.450 541.950 ;
        RECT 302.400 526.200 303.600 526.950 ;
        RECT 338.400 526.200 339.600 526.950 ;
        RECT 662.400 526.200 663.600 528.600 ;
      LAYER metal3 ;
        RECT 568.950 822.600 571.050 823.050 ;
        RECT 586.950 822.600 589.050 823.050 ;
        RECT 568.950 821.400 589.050 822.600 ;
        RECT 568.950 820.950 571.050 821.400 ;
        RECT 586.950 820.950 589.050 821.400 ;
        RECT 586.950 810.600 589.050 811.050 ;
        RECT 607.950 810.600 610.050 811.050 ;
        RECT 586.950 809.400 610.050 810.600 ;
        RECT 586.950 808.950 589.050 809.400 ;
        RECT 607.950 808.950 610.050 809.400 ;
        RECT 607.950 789.600 610.050 790.050 ;
        RECT 628.950 789.600 631.050 789.900 ;
        RECT 607.950 788.400 631.050 789.600 ;
        RECT 607.950 787.950 610.050 788.400 ;
        RECT 628.950 787.800 631.050 788.400 ;
        RECT 628.950 741.600 631.050 742.050 ;
        RECT 646.950 741.600 649.050 742.050 ;
        RECT 628.950 740.400 649.050 741.600 ;
        RECT 628.950 739.950 631.050 740.400 ;
        RECT 646.950 739.950 649.050 740.400 ;
        RECT 580.950 714.600 583.050 715.050 ;
        RECT 646.950 714.600 649.050 715.050 ;
        RECT 580.950 713.400 649.050 714.600 ;
        RECT 580.950 712.950 583.050 713.400 ;
        RECT 646.950 712.950 649.050 713.400 ;
        RECT 562.950 672.600 565.050 673.050 ;
        RECT 580.950 672.600 583.050 673.050 ;
        RECT 562.950 671.400 583.050 672.600 ;
        RECT 562.950 670.950 565.050 671.400 ;
        RECT 580.950 670.950 583.050 671.400 ;
        RECT 541.950 660.600 544.050 661.050 ;
        RECT 553.950 660.600 556.050 661.050 ;
        RECT 562.950 660.600 565.050 661.050 ;
        RECT 541.950 659.400 565.050 660.600 ;
        RECT 541.950 658.950 544.050 659.400 ;
        RECT 553.950 658.950 556.050 659.400 ;
        RECT 562.950 658.950 565.050 659.400 ;
        RECT 553.950 651.600 558.000 652.050 ;
        RECT 553.950 649.950 558.600 651.600 ;
        RECT 457.950 645.600 460.050 646.050 ;
        RECT 484.800 645.600 486.900 646.050 ;
        RECT 457.950 644.400 486.900 645.600 ;
        RECT 457.950 643.950 460.050 644.400 ;
        RECT 484.800 643.950 486.900 644.400 ;
        RECT 547.950 645.600 550.050 646.050 ;
        RECT 557.400 645.600 558.600 649.950 ;
        RECT 547.950 644.400 561.600 645.600 ;
        RECT 547.950 643.950 550.050 644.400 ;
        RECT 560.400 642.600 561.600 644.400 ;
        RECT 583.950 642.600 586.050 643.050 ;
        RECT 560.400 641.400 586.050 642.600 ;
        RECT 583.950 640.950 586.050 641.400 ;
        RECT 424.950 636.600 427.050 637.050 ;
        RECT 457.950 636.600 460.050 637.050 ;
        RECT 424.950 635.400 460.050 636.600 ;
        RECT 424.950 634.950 427.050 635.400 ;
        RECT 457.950 634.950 460.050 635.400 ;
        RECT 484.950 636.600 487.050 637.050 ;
        RECT 547.950 636.600 550.050 637.050 ;
        RECT 484.950 635.400 550.050 636.600 ;
        RECT 484.950 634.950 487.050 635.400 ;
        RECT 547.950 634.950 550.050 635.400 ;
        RECT 583.950 618.600 586.050 619.050 ;
        RECT 610.950 618.600 613.050 619.050 ;
        RECT 583.950 617.400 613.050 618.600 ;
        RECT 583.950 616.950 586.050 617.400 ;
        RECT 610.950 616.950 613.050 617.400 ;
        RECT 610.950 609.600 613.050 610.050 ;
        RECT 622.950 609.600 625.050 610.050 ;
        RECT 610.950 608.400 625.050 609.600 ;
        RECT 610.950 607.950 613.050 608.400 ;
        RECT 622.950 607.950 625.050 608.400 ;
        RECT 547.950 606.600 550.050 607.050 ;
        RECT 547.950 605.400 561.600 606.600 ;
        RECT 547.950 604.950 550.050 605.400 ;
        RECT 560.400 601.050 561.600 605.400 ;
        RECT 424.950 600.300 427.050 600.750 ;
        RECT 436.950 600.300 439.050 600.750 ;
        RECT 424.950 599.100 439.050 600.300 ;
        RECT 424.950 598.650 427.050 599.100 ;
        RECT 436.950 598.650 439.050 599.100 ;
        RECT 559.950 598.950 562.050 601.050 ;
        RECT 361.950 585.600 364.050 586.050 ;
        RECT 424.950 585.600 427.050 586.050 ;
        RECT 361.950 584.400 427.050 585.600 ;
        RECT 361.950 583.950 364.050 584.400 ;
        RECT 424.950 583.950 427.050 584.400 ;
        RECT 310.950 572.250 313.050 574.350 ;
        RECT 311.400 568.050 312.600 572.250 ;
        RECT 310.950 565.950 313.050 568.050 ;
        RECT 586.950 558.600 589.050 559.050 ;
        RECT 628.800 558.600 630.900 559.050 ;
        RECT 586.950 557.400 630.900 558.600 ;
        RECT 586.950 556.950 589.050 557.400 ;
        RECT 628.800 556.950 630.900 557.400 ;
        RECT 556.950 552.600 559.050 553.050 ;
        RECT 586.950 552.600 589.050 553.050 ;
        RECT 556.950 551.400 589.050 552.600 ;
        RECT 556.950 550.950 559.050 551.400 ;
        RECT 586.950 550.950 589.050 551.400 ;
        RECT 628.950 543.600 631.050 544.050 ;
        RECT 661.950 543.600 664.050 544.050 ;
        RECT 628.950 542.400 664.050 543.600 ;
        RECT 628.950 541.950 631.050 542.400 ;
        RECT 661.950 541.950 664.050 542.400 ;
        RECT 310.950 528.600 313.050 532.050 ;
        RECT 337.950 528.600 340.050 529.050 ;
        RECT 358.950 528.600 361.050 529.050 ;
        RECT 310.950 528.000 361.050 528.600 ;
        RECT 311.400 527.400 361.050 528.000 ;
        RECT 337.950 526.950 340.050 527.400 ;
        RECT 358.950 526.950 361.050 527.400 ;
    END
  END Cin[3]
  PIN Cin[2]
    PORT
      LAYER metal1 ;
        RECT 589.950 801.450 592.050 802.050 ;
        RECT 595.950 801.450 598.050 802.050 ;
        RECT 589.950 800.550 598.050 801.450 ;
        RECT 589.950 799.950 592.050 800.550 ;
        RECT 595.950 799.950 598.050 800.550 ;
        RECT 703.950 765.450 706.050 766.050 ;
        RECT 703.950 765.000 711.450 765.450 ;
        RECT 703.950 764.550 712.050 765.000 ;
        RECT 703.950 763.950 706.050 764.550 ;
        RECT 709.950 760.800 712.050 764.550 ;
        RECT 696.000 729.450 700.050 730.050 ;
        RECT 695.550 727.950 700.050 729.450 ;
        RECT 695.550 724.050 696.450 727.950 ;
        RECT 691.950 722.550 696.450 724.050 ;
        RECT 691.950 721.950 696.000 722.550 ;
        RECT 166.950 645.450 169.050 646.050 ;
        RECT 172.950 645.450 175.050 646.050 ;
        RECT 166.950 644.550 175.050 645.450 ;
        RECT 166.950 643.950 169.050 644.550 ;
        RECT 172.950 643.950 175.050 644.550 ;
      LAYER metal2 ;
        RECT 512.400 825.450 513.450 828.450 ;
        RECT 512.400 824.400 519.450 825.450 ;
        RECT 232.950 820.950 235.050 823.050 ;
        RECT 304.950 820.950 307.050 823.050 ;
        RECT 463.950 820.950 466.050 823.050 ;
        RECT 233.400 814.050 234.450 820.950 ;
        RECT 208.950 811.950 211.050 814.050 ;
        RECT 232.950 811.950 235.050 814.050 ;
        RECT 209.400 766.050 210.450 811.950 ;
        RECT 233.400 807.600 234.450 811.950 ;
        RECT 305.400 811.050 306.450 820.950 ;
        RECT 304.950 808.950 307.050 811.050 ;
        RECT 310.950 808.950 313.050 811.050 ;
        RECT 233.400 805.500 234.600 807.600 ;
        RECT 311.400 781.050 312.450 808.950 ;
        RECT 464.400 808.050 465.450 820.950 ;
        RECT 475.950 819.450 478.050 823.050 ;
        RECT 512.400 820.050 513.450 824.400 ;
        RECT 518.400 820.050 519.450 824.400 ;
        RECT 631.950 820.950 634.050 823.050 ;
        RECT 685.950 820.950 688.050 823.050 ;
        RECT 481.950 819.450 484.050 820.050 ;
        RECT 475.950 819.000 484.050 819.450 ;
        RECT 476.400 818.400 484.050 819.000 ;
        RECT 481.950 817.950 484.050 818.400 ;
        RECT 511.950 817.950 514.050 820.050 ;
        RECT 517.950 817.950 520.050 820.050 ;
        RECT 559.950 817.950 562.050 820.050 ;
        RECT 560.400 811.050 561.450 817.950 ;
        RECT 632.400 817.050 633.450 820.950 ;
        RECT 589.950 814.950 592.050 817.050 ;
        RECT 607.950 816.450 610.050 817.050 ;
        RECT 613.950 816.450 616.050 817.050 ;
        RECT 607.950 815.400 616.050 816.450 ;
        RECT 607.950 814.950 610.050 815.400 ;
        RECT 613.950 814.950 616.050 815.400 ;
        RECT 631.950 814.950 634.050 817.050 ;
        RECT 559.950 808.950 562.050 811.050 ;
        RECT 463.950 805.950 466.050 808.050 ;
        RECT 590.400 805.050 591.450 814.950 ;
        RECT 686.400 814.050 687.450 820.950 ;
        RECT 685.950 811.950 688.050 814.050 ;
        RECT 697.950 811.950 700.050 814.050 ;
        RECT 338.400 800.400 339.600 802.800 ;
        RECT 338.400 781.050 339.450 800.400 ;
        RECT 463.950 799.950 466.050 802.050 ;
        RECT 589.950 799.950 592.050 805.050 ;
        RECT 596.400 802.050 597.600 802.800 ;
        RECT 595.950 799.950 598.050 802.050 ;
        RECT 310.950 778.950 313.050 781.050 ;
        RECT 337.950 778.950 340.050 781.050 ;
        RECT 464.400 778.050 465.450 799.950 ;
        RECT 463.950 775.950 466.050 778.050 ;
        RECT 698.400 775.050 699.450 811.950 ;
        RECT 697.950 772.950 700.050 775.050 ;
        RECT 703.950 772.950 706.050 775.050 ;
        RECT 704.400 766.050 705.450 772.950 ;
        RECT 199.950 763.950 202.050 766.050 ;
        RECT 208.950 763.950 211.050 766.050 ;
        RECT 703.950 763.950 706.050 766.050 ;
        RECT 200.400 733.050 201.450 763.950 ;
        RECT 709.950 760.800 712.050 762.900 ;
        RECT 710.400 745.050 711.450 760.800 ;
        RECT 697.950 742.800 700.050 744.900 ;
        RECT 709.950 742.950 712.050 745.050 ;
        RECT 184.950 730.950 187.050 733.050 ;
        RECT 199.950 730.950 202.050 733.050 ;
        RECT 161.400 724.050 162.600 724.800 ;
        RECT 185.400 724.050 186.450 730.950 ;
        RECT 698.400 730.050 699.450 742.800 ;
        RECT 697.950 727.950 700.050 730.050 ;
        RECT 160.950 723.450 163.050 724.050 ;
        RECT 158.400 722.400 163.050 723.450 ;
        RECT 158.400 658.050 159.450 722.400 ;
        RECT 160.950 721.950 163.050 722.400 ;
        RECT 184.800 721.950 186.900 724.050 ;
        RECT 691.950 721.950 694.050 724.050 ;
        RECT 692.400 718.050 693.450 721.950 ;
        RECT 661.950 715.950 664.050 718.050 ;
        RECT 691.950 715.950 694.050 718.050 ;
        RECT 589.950 700.950 592.050 703.050 ;
        RECT 598.950 700.950 601.050 703.050 ;
        RECT 590.400 684.600 591.450 700.950 ;
        RECT 599.400 691.050 600.450 700.950 ;
        RECT 662.400 694.050 663.450 715.950 ;
        RECT 661.950 691.950 664.050 694.050 ;
        RECT 598.950 688.950 601.050 691.050 ;
        RECT 607.950 688.950 610.050 691.050 ;
        RECT 608.400 684.600 609.450 688.950 ;
        RECT 590.400 682.200 591.600 684.600 ;
        RECT 608.400 682.200 609.600 684.600 ;
        RECT 157.950 655.950 160.050 658.050 ;
        RECT 172.950 655.950 175.050 658.050 ;
        RECT 167.400 646.050 168.600 646.800 ;
        RECT 173.400 646.050 174.450 655.950 ;
        RECT 166.950 643.950 169.050 646.050 ;
        RECT 172.950 643.950 175.050 646.050 ;
        RECT 167.400 622.050 168.450 643.950 ;
        RECT 157.950 619.950 160.050 622.050 ;
        RECT 166.800 619.950 168.900 622.050 ;
        RECT 158.400 607.050 159.450 619.950 ;
        RECT 157.950 604.950 160.050 607.050 ;
        RECT 154.950 598.950 157.050 601.050 ;
        RECT 155.400 585.450 156.450 598.950 ;
        RECT 155.400 584.400 159.450 585.450 ;
        RECT 145.950 577.800 148.050 579.900 ;
        RECT 151.950 579.600 154.050 580.050 ;
        RECT 158.400 579.600 159.450 584.400 ;
        RECT 151.950 578.550 159.450 579.600 ;
        RECT 151.950 577.950 154.050 578.550 ;
        RECT 146.400 574.050 147.450 577.800 ;
        RECT 145.950 571.950 148.050 574.050 ;
        RECT 145.950 565.950 148.050 568.050 ;
        RECT 146.400 529.050 147.450 565.950 ;
        RECT 145.950 526.950 148.050 529.050 ;
        RECT 163.950 523.800 166.050 525.900 ;
        RECT 164.400 508.050 165.450 523.800 ;
        RECT 163.950 505.950 166.050 508.050 ;
        RECT 187.950 505.950 190.050 508.050 ;
        RECT 188.400 490.050 189.450 505.950 ;
        RECT 197.400 490.050 198.600 490.800 ;
        RECT 187.950 487.950 190.050 490.050 ;
        RECT 196.950 487.950 199.050 490.050 ;
        RECT 188.400 463.050 189.450 487.950 ;
        RECT 181.950 460.950 184.050 463.050 ;
        RECT 187.950 460.950 190.050 463.050 ;
        RECT 182.400 450.600 183.450 460.950 ;
        RECT 182.400 448.200 183.600 450.600 ;
      LAYER metal3 ;
        RECT 232.950 822.600 235.050 823.050 ;
        RECT 304.950 822.600 307.050 823.050 ;
        RECT 232.950 821.400 307.050 822.600 ;
        RECT 232.950 820.950 235.050 821.400 ;
        RECT 304.950 820.950 307.050 821.400 ;
        RECT 463.950 822.600 466.050 823.050 ;
        RECT 475.950 822.600 478.050 823.050 ;
        RECT 463.950 821.400 478.050 822.600 ;
        RECT 463.950 820.950 466.050 821.400 ;
        RECT 475.950 820.950 478.050 821.400 ;
        RECT 631.950 822.600 634.050 823.050 ;
        RECT 685.950 822.600 688.050 823.050 ;
        RECT 631.950 821.400 688.050 822.600 ;
        RECT 631.950 820.950 634.050 821.400 ;
        RECT 685.950 820.950 688.050 821.400 ;
        RECT 481.950 819.600 484.050 820.050 ;
        RECT 511.950 819.600 514.050 820.050 ;
        RECT 481.950 818.400 514.050 819.600 ;
        RECT 481.950 817.950 484.050 818.400 ;
        RECT 511.950 817.950 514.050 818.400 ;
        RECT 517.950 819.600 520.050 820.050 ;
        RECT 559.950 819.600 562.050 820.050 ;
        RECT 517.950 818.400 562.050 819.600 ;
        RECT 517.950 817.950 520.050 818.400 ;
        RECT 559.950 817.950 562.050 818.400 ;
        RECT 589.950 816.600 592.050 817.050 ;
        RECT 607.950 816.600 610.050 817.050 ;
        RECT 589.950 815.400 610.050 816.600 ;
        RECT 589.950 814.950 592.050 815.400 ;
        RECT 607.950 814.950 610.050 815.400 ;
        RECT 613.950 816.600 616.050 817.050 ;
        RECT 631.950 816.600 634.050 817.050 ;
        RECT 613.950 815.400 634.050 816.600 ;
        RECT 613.950 814.950 616.050 815.400 ;
        RECT 631.950 814.950 634.050 815.400 ;
        RECT 208.950 813.600 211.050 814.050 ;
        RECT 232.950 813.600 235.050 814.050 ;
        RECT 208.950 812.400 235.050 813.600 ;
        RECT 208.950 811.950 211.050 812.400 ;
        RECT 232.950 811.950 235.050 812.400 ;
        RECT 685.950 813.600 688.050 814.050 ;
        RECT 697.950 813.600 700.050 814.050 ;
        RECT 685.950 812.400 700.050 813.600 ;
        RECT 685.950 811.950 688.050 812.400 ;
        RECT 697.950 811.950 700.050 812.400 ;
        RECT 304.950 810.600 307.050 811.050 ;
        RECT 310.950 810.600 313.050 811.050 ;
        RECT 304.950 809.400 313.050 810.600 ;
        RECT 304.950 808.950 307.050 809.400 ;
        RECT 310.950 808.950 313.050 809.400 ;
        RECT 559.950 808.950 562.050 811.050 ;
        RECT 463.950 805.950 466.050 808.050 ;
        RECT 464.400 802.050 465.600 805.950 ;
        RECT 560.400 804.600 561.600 808.950 ;
        RECT 589.950 804.600 592.050 805.050 ;
        RECT 560.400 803.400 592.050 804.600 ;
        RECT 589.950 802.950 592.050 803.400 ;
        RECT 463.950 799.950 466.050 802.050 ;
        RECT 310.950 780.600 313.050 781.050 ;
        RECT 337.950 780.600 340.050 781.050 ;
        RECT 310.950 779.400 408.600 780.600 ;
        RECT 310.950 778.950 313.050 779.400 ;
        RECT 337.950 778.950 340.050 779.400 ;
        RECT 407.400 777.600 408.600 779.400 ;
        RECT 463.950 777.600 466.050 778.050 ;
        RECT 407.400 776.400 466.050 777.600 ;
        RECT 463.950 775.950 466.050 776.400 ;
        RECT 697.950 774.600 700.050 775.050 ;
        RECT 703.950 774.600 706.050 775.050 ;
        RECT 697.950 773.400 706.050 774.600 ;
        RECT 697.950 772.950 700.050 773.400 ;
        RECT 703.950 772.950 706.050 773.400 ;
        RECT 199.950 765.600 202.050 766.050 ;
        RECT 208.950 765.600 211.050 766.050 ;
        RECT 199.950 764.400 211.050 765.600 ;
        RECT 199.950 763.950 202.050 764.400 ;
        RECT 208.950 763.950 211.050 764.400 ;
        RECT 697.950 744.600 700.050 744.900 ;
        RECT 709.950 744.600 712.050 745.050 ;
        RECT 697.950 743.400 712.050 744.600 ;
        RECT 697.950 742.800 700.050 743.400 ;
        RECT 709.950 742.950 712.050 743.400 ;
        RECT 184.950 732.600 187.050 733.050 ;
        RECT 199.950 732.600 202.050 733.050 ;
        RECT 184.950 731.400 202.050 732.600 ;
        RECT 184.950 730.950 187.050 731.400 ;
        RECT 199.950 730.950 202.050 731.400 ;
        RECT 160.950 723.600 163.050 724.050 ;
        RECT 184.800 723.600 186.900 724.050 ;
        RECT 160.950 722.400 186.900 723.600 ;
        RECT 160.950 721.950 163.050 722.400 ;
        RECT 184.800 721.950 186.900 722.400 ;
        RECT 661.950 717.600 664.050 718.050 ;
        RECT 691.950 717.600 694.050 718.050 ;
        RECT 661.950 716.400 694.050 717.600 ;
        RECT 661.950 715.950 664.050 716.400 ;
        RECT 691.950 715.950 694.050 716.400 ;
        RECT 589.950 702.600 592.050 703.050 ;
        RECT 598.950 702.600 601.050 703.050 ;
        RECT 589.950 701.400 601.050 702.600 ;
        RECT 589.950 700.950 592.050 701.400 ;
        RECT 598.950 700.950 601.050 701.400 ;
        RECT 660.000 693.600 664.050 694.050 ;
        RECT 659.400 691.950 664.050 693.600 ;
        RECT 598.950 690.600 601.050 691.050 ;
        RECT 607.950 690.600 610.050 691.050 ;
        RECT 659.400 690.600 660.600 691.950 ;
        RECT 598.950 689.400 660.600 690.600 ;
        RECT 598.950 688.950 601.050 689.400 ;
        RECT 607.950 688.950 610.050 689.400 ;
        RECT 157.950 657.600 160.050 658.050 ;
        RECT 172.950 657.600 175.050 658.050 ;
        RECT 157.950 656.400 175.050 657.600 ;
        RECT 157.950 655.950 160.050 656.400 ;
        RECT 172.950 655.950 175.050 656.400 ;
        RECT 157.950 621.600 160.050 622.050 ;
        RECT 166.800 621.600 168.900 622.050 ;
        RECT 157.950 620.400 168.900 621.600 ;
        RECT 157.950 619.950 160.050 620.400 ;
        RECT 166.800 619.950 168.900 620.400 ;
        RECT 157.950 603.600 160.050 607.050 ;
        RECT 155.400 603.000 160.050 603.600 ;
        RECT 154.950 602.400 159.600 603.000 ;
        RECT 154.950 598.950 157.050 602.400 ;
        RECT 145.950 579.600 148.050 579.900 ;
        RECT 151.950 579.600 154.050 580.050 ;
        RECT 145.950 578.400 154.050 579.600 ;
        RECT 145.950 577.800 148.050 578.400 ;
        RECT 151.950 577.950 154.050 578.400 ;
        RECT 145.950 571.950 148.050 574.050 ;
        RECT 146.400 568.050 147.600 571.950 ;
        RECT 145.950 565.950 148.050 568.050 ;
        RECT 145.950 528.600 148.050 529.050 ;
        RECT 145.950 528.000 165.600 528.600 ;
        RECT 145.950 527.400 166.050 528.000 ;
        RECT 145.950 526.950 148.050 527.400 ;
        RECT 163.950 523.800 166.050 527.400 ;
        RECT 163.950 507.600 166.050 508.050 ;
        RECT 187.950 507.600 190.050 508.050 ;
        RECT 163.950 506.400 190.050 507.600 ;
        RECT 163.950 505.950 166.050 506.400 ;
        RECT 187.950 505.950 190.050 506.400 ;
        RECT 187.950 489.600 190.050 490.050 ;
        RECT 196.950 489.600 199.050 490.050 ;
        RECT 187.950 488.400 199.050 489.600 ;
        RECT 187.950 487.950 190.050 488.400 ;
        RECT 196.950 487.950 199.050 488.400 ;
        RECT 181.950 462.600 184.050 463.050 ;
        RECT 187.950 462.600 190.050 463.050 ;
        RECT 181.950 461.400 190.050 462.600 ;
        RECT 181.950 460.950 184.050 461.400 ;
        RECT 187.950 460.950 190.050 461.400 ;
    END
  END Cin[2]
  PIN Cin[1]
    PORT
      LAYER metal1 ;
        RECT 508.950 763.950 511.050 766.050 ;
        RECT 509.550 757.050 510.450 763.950 ;
        RECT 505.950 755.550 510.450 757.050 ;
        RECT 505.950 754.950 510.000 755.550 ;
      LAYER metal2 ;
        RECT 503.400 823.050 504.450 828.450 ;
        RECT 484.950 820.950 487.050 823.050 ;
        RECT 502.950 820.950 505.050 823.050 ;
        RECT 358.950 817.950 361.050 820.050 ;
        RECT 427.950 817.950 430.050 820.050 ;
        RECT 359.400 811.050 360.450 817.950 ;
        RECT 346.950 808.950 349.050 811.050 ;
        RECT 145.950 805.950 148.050 808.050 ;
        RECT 157.950 806.100 160.050 808.200 ;
        RECT 146.400 784.050 147.450 805.950 ;
        RECT 158.400 805.350 159.600 806.100 ;
        RECT 347.400 787.050 348.450 808.950 ;
        RECT 358.950 807.000 361.050 811.050 ;
        RECT 359.400 805.350 360.600 807.000 ;
        RECT 428.400 787.050 429.450 817.950 ;
        RECT 485.400 816.450 486.450 820.950 ;
        RECT 482.400 815.400 486.450 816.450 ;
        RECT 482.400 801.450 483.450 815.400 ;
        RECT 479.400 800.400 483.450 801.450 ;
        RECT 479.400 787.050 480.450 800.400 ;
        RECT 328.950 784.950 331.050 787.050 ;
        RECT 346.950 784.950 349.050 787.050 ;
        RECT 427.950 784.950 430.050 787.050 ;
        RECT 478.950 784.950 481.050 787.050 ;
        RECT 508.950 784.950 511.050 787.050 ;
        RECT 145.950 781.950 148.050 784.050 ;
        RECT 157.950 781.950 160.050 784.050 ;
        RECT 158.400 775.050 159.450 781.950 ;
        RECT 329.400 775.050 330.450 784.950 ;
        RECT 157.950 772.950 160.050 775.050 ;
        RECT 328.950 772.950 331.050 775.050 ;
        RECT 158.400 745.050 159.450 772.950 ;
        RECT 509.400 766.050 510.450 784.950 ;
        RECT 508.950 763.950 511.050 766.050 ;
        RECT 505.950 754.950 508.050 757.050 ;
        RECT 157.950 742.950 160.050 745.050 ;
        RECT 172.950 742.950 175.050 745.050 ;
        RECT 173.400 729.600 174.450 742.950 ;
        RECT 506.400 733.050 507.450 754.950 ;
        RECT 173.400 727.350 174.600 729.600 ;
        RECT 496.950 729.000 499.050 733.050 ;
        RECT 505.950 730.950 508.050 733.050 ;
        RECT 497.400 727.350 498.600 729.000 ;
      LAYER metal3 ;
        RECT 484.950 822.600 487.050 823.050 ;
        RECT 502.950 822.600 505.050 823.050 ;
        RECT 484.950 821.400 505.050 822.600 ;
        RECT 484.950 820.950 487.050 821.400 ;
        RECT 502.950 820.950 505.050 821.400 ;
        RECT 358.950 819.600 361.050 820.050 ;
        RECT 427.950 819.600 430.050 820.050 ;
        RECT 358.950 818.400 430.050 819.600 ;
        RECT 358.950 817.950 361.050 818.400 ;
        RECT 427.950 817.950 430.050 818.400 ;
        RECT 346.950 810.600 349.050 811.050 ;
        RECT 358.950 810.600 361.050 811.050 ;
        RECT 346.950 809.400 361.050 810.600 ;
        RECT 346.950 808.950 349.050 809.400 ;
        RECT 358.950 808.950 361.050 809.400 ;
        RECT 145.950 807.600 148.050 808.050 ;
        RECT 157.950 807.600 160.050 808.200 ;
        RECT 145.950 806.400 160.050 807.600 ;
        RECT 145.950 805.950 148.050 806.400 ;
        RECT 157.950 806.100 160.050 806.400 ;
        RECT 328.950 786.600 331.050 787.050 ;
        RECT 346.950 786.600 349.050 787.050 ;
        RECT 328.950 785.400 349.050 786.600 ;
        RECT 328.950 784.950 331.050 785.400 ;
        RECT 346.950 784.950 349.050 785.400 ;
        RECT 427.950 786.600 430.050 787.050 ;
        RECT 478.950 786.600 481.050 787.050 ;
        RECT 508.950 786.600 511.050 787.050 ;
        RECT 427.950 785.400 511.050 786.600 ;
        RECT 427.950 784.950 430.050 785.400 ;
        RECT 478.950 784.950 481.050 785.400 ;
        RECT 508.950 784.950 511.050 785.400 ;
        RECT 145.950 783.600 148.050 784.050 ;
        RECT 157.950 783.600 160.050 784.050 ;
        RECT 145.950 782.400 160.050 783.600 ;
        RECT 145.950 781.950 148.050 782.400 ;
        RECT 157.950 781.950 160.050 782.400 ;
        RECT 157.950 774.600 160.050 775.050 ;
        RECT 328.950 774.600 331.050 775.050 ;
        RECT 157.950 773.400 331.050 774.600 ;
        RECT 157.950 772.950 160.050 773.400 ;
        RECT 328.950 772.950 331.050 773.400 ;
        RECT 157.950 744.600 160.050 745.050 ;
        RECT 172.950 744.600 175.050 745.050 ;
        RECT 157.950 743.400 175.050 744.600 ;
        RECT 157.950 742.950 160.050 743.400 ;
        RECT 172.950 742.950 175.050 743.400 ;
        RECT 496.950 732.600 499.050 733.050 ;
        RECT 505.950 732.600 508.050 733.050 ;
        RECT 496.950 731.400 508.050 732.600 ;
        RECT 496.950 730.950 499.050 731.400 ;
        RECT 505.950 730.950 508.050 731.400 ;
    END
  END Cin[1]
  PIN Cin[0]
    PORT
      LAYER metal2 ;
        RECT 494.400 827.400 498.450 828.450 ;
        RECT 494.400 825.450 495.450 827.400 ;
        RECT 491.400 824.400 495.450 825.450 ;
        RECT 433.950 820.950 436.050 823.050 ;
        RECT 220.950 817.950 223.050 820.050 ;
        RECT 221.400 808.200 222.450 817.950 ;
        RECT 434.400 811.050 435.450 820.950 ;
        RECT 491.400 817.050 492.450 824.400 ;
        RECT 442.950 814.950 445.050 817.050 ;
        RECT 490.800 814.950 492.900 817.050 ;
        RECT 443.400 811.050 444.450 814.950 ;
        RECT 433.950 808.950 436.050 811.050 ;
        RECT 442.950 808.950 445.050 811.050 ;
        RECT 220.950 806.100 223.050 808.200 ;
        RECT 443.400 807.600 444.450 808.950 ;
        RECT 221.400 805.350 222.600 806.100 ;
        RECT 443.400 805.350 444.600 807.600 ;
        RECT 238.800 799.950 240.900 802.050 ;
        RECT 239.400 762.450 240.450 799.950 ;
        RECT 239.400 761.400 243.450 762.450 ;
        RECT 242.400 745.050 243.450 761.400 ;
        RECT 241.950 742.950 244.050 745.050 ;
        RECT 271.950 742.950 274.050 745.050 ;
        RECT 160.950 715.950 163.050 718.050 ;
        RECT 161.400 685.050 162.450 715.950 ;
        RECT 232.950 715.800 235.050 717.900 ;
        RECT 233.400 703.050 234.450 715.800 ;
        RECT 272.400 703.050 273.450 742.950 ;
        RECT 232.950 700.950 235.050 703.050 ;
        RECT 271.950 700.950 274.050 703.050 ;
        RECT 272.400 697.050 273.450 700.950 ;
        RECT 271.950 694.950 274.050 697.050 ;
        RECT 280.950 694.950 283.050 697.050 ;
        RECT 160.950 682.950 163.050 685.050 ;
        RECT 152.400 679.050 153.600 679.650 ;
        RECT 152.400 677.400 157.050 679.050 ;
        RECT 266.400 678.000 267.600 679.650 ;
        RECT 153.000 676.950 157.050 677.400 ;
        RECT 265.950 673.950 268.050 678.000 ;
        RECT 281.400 676.050 282.450 694.950 ;
        RECT 280.950 673.950 283.050 676.050 ;
      LAYER metal3 ;
        RECT 433.950 822.600 436.050 823.050 ;
        RECT 314.400 821.400 436.050 822.600 ;
        RECT 220.950 819.600 223.050 820.050 ;
        RECT 314.400 819.600 315.600 821.400 ;
        RECT 433.950 820.950 436.050 821.400 ;
        RECT 220.950 818.400 315.600 819.600 ;
        RECT 220.950 817.950 223.050 818.400 ;
        RECT 442.950 816.600 445.050 817.050 ;
        RECT 490.800 816.600 492.900 817.050 ;
        RECT 442.950 815.400 492.900 816.600 ;
        RECT 442.950 814.950 445.050 815.400 ;
        RECT 490.800 814.950 492.900 815.400 ;
        RECT 433.950 810.600 436.050 811.050 ;
        RECT 442.950 810.600 445.050 811.050 ;
        RECT 433.950 809.400 445.050 810.600 ;
        RECT 433.950 808.950 436.050 809.400 ;
        RECT 442.950 808.950 445.050 809.400 ;
        RECT 220.950 807.600 223.050 808.200 ;
        RECT 220.950 806.400 237.600 807.600 ;
        RECT 220.950 806.100 223.050 806.400 ;
        RECT 236.400 804.600 237.600 806.400 ;
        RECT 236.400 804.000 240.450 804.600 ;
        RECT 236.400 803.400 241.050 804.000 ;
        RECT 238.950 802.050 241.050 803.400 ;
        RECT 238.800 801.000 241.050 802.050 ;
        RECT 238.800 799.950 240.900 801.000 ;
        RECT 241.950 744.600 244.050 745.050 ;
        RECT 271.950 744.600 274.050 745.050 ;
        RECT 241.950 743.400 274.050 744.600 ;
        RECT 241.950 742.950 244.050 743.400 ;
        RECT 271.950 742.950 274.050 743.400 ;
        RECT 160.950 717.600 163.050 718.050 ;
        RECT 232.950 717.600 235.050 717.900 ;
        RECT 160.950 716.400 235.050 717.600 ;
        RECT 160.950 715.950 163.050 716.400 ;
        RECT 232.950 715.800 235.050 716.400 ;
        RECT 232.950 702.600 235.050 703.050 ;
        RECT 271.950 702.600 274.050 703.050 ;
        RECT 232.950 701.400 274.050 702.600 ;
        RECT 232.950 700.950 235.050 701.400 ;
        RECT 271.950 700.950 274.050 701.400 ;
        RECT 271.950 696.600 274.050 697.050 ;
        RECT 280.950 696.600 283.050 697.050 ;
        RECT 271.950 695.400 283.050 696.600 ;
        RECT 271.950 694.950 274.050 695.400 ;
        RECT 280.950 694.950 283.050 695.400 ;
        RECT 160.950 684.600 163.050 685.050 ;
        RECT 155.400 683.400 163.050 684.600 ;
        RECT 155.400 679.050 156.600 683.400 ;
        RECT 160.950 682.950 163.050 683.400 ;
        RECT 154.950 676.950 157.050 679.050 ;
        RECT 265.950 675.600 268.050 676.050 ;
        RECT 280.950 675.600 283.050 676.050 ;
        RECT 265.950 674.400 283.050 675.600 ;
        RECT 265.950 673.950 268.050 674.400 ;
        RECT 280.950 673.950 283.050 674.400 ;
    END
  END Cin[0]
  PIN Rdy
    PORT
      LAYER metal2 ;
        RECT 1.950 298.950 4.050 301.050 ;
        RECT 55.950 298.950 58.050 301.050 ;
        RECT 2.400 295.050 3.450 298.950 ;
        RECT 1.950 292.950 4.050 295.050 ;
        RECT 56.400 294.600 57.450 298.950 ;
        RECT 56.400 292.350 57.600 294.600 ;
      LAYER metal3 ;
        RECT 1.950 300.600 4.050 301.050 ;
        RECT 55.950 300.600 58.050 301.050 ;
        RECT 1.950 299.400 58.050 300.600 ;
        RECT 1.950 298.950 4.050 299.400 ;
        RECT 55.950 298.950 58.050 299.400 ;
        RECT 1.950 294.600 4.050 295.050 ;
        RECT -3.600 293.400 4.050 294.600 ;
        RECT 1.950 292.950 4.050 293.400 ;
    END
  END Rdy
  PIN Vld
    PORT
      LAYER metal2 ;
        RECT 842.400 410.400 843.600 412.650 ;
        RECT 842.400 406.050 843.450 410.400 ;
        RECT 850.950 409.950 853.050 412.050 ;
        RECT 851.400 406.050 852.450 409.950 ;
        RECT 841.950 403.950 844.050 406.050 ;
        RECT 850.950 403.950 853.050 406.050 ;
      LAYER metal3 ;
        RECT 850.950 411.600 853.050 412.050 ;
        RECT 850.950 410.400 870.600 411.600 ;
        RECT 850.950 409.950 853.050 410.400 ;
        RECT 841.950 405.600 844.050 406.050 ;
        RECT 850.950 405.600 853.050 406.050 ;
        RECT 841.950 404.400 853.050 405.600 ;
        RECT 841.950 403.950 844.050 404.400 ;
        RECT 850.950 403.950 853.050 404.400 ;
    END
  END Vld
  PIN Xin[3]
    PORT
      LAYER metal1 ;
        RECT 6.000 528.450 10.050 529.050 ;
        RECT 5.550 526.950 10.050 528.450 ;
        RECT 5.550 523.050 6.450 526.950 ;
        RECT 5.550 521.550 10.050 523.050 ;
        RECT 6.000 520.950 10.050 521.550 ;
        RECT 424.950 486.450 427.050 487.050 ;
        RECT 439.950 486.450 442.050 487.050 ;
        RECT 424.950 485.550 442.050 486.450 ;
        RECT 424.950 484.950 427.050 485.550 ;
        RECT 439.950 484.950 442.050 485.550 ;
        RECT 55.950 456.450 58.050 457.050 ;
        RECT 67.950 456.450 70.050 457.050 ;
        RECT 55.950 455.550 70.050 456.450 ;
        RECT 55.950 454.950 58.050 455.550 ;
        RECT 67.950 454.950 70.050 455.550 ;
        RECT 216.000 450.450 220.050 451.050 ;
        RECT 215.550 448.950 220.050 450.450 ;
        RECT 215.550 445.050 216.450 448.950 ;
        RECT 215.550 443.550 220.050 445.050 ;
        RECT 216.000 442.950 220.050 443.550 ;
      LAYER metal2 ;
        RECT 7.950 532.950 10.050 535.050 ;
        RECT 8.400 529.050 9.450 532.950 ;
        RECT 7.950 526.950 10.050 529.050 ;
        RECT 481.950 526.950 484.050 529.050 ;
        RECT 490.950 526.950 493.050 529.050 ;
        RECT 7.950 520.950 10.050 523.050 ;
        RECT 8.400 517.050 9.450 520.950 ;
        RECT 7.950 514.950 10.050 517.050 ;
        RECT 19.950 514.950 22.050 517.050 ;
        RECT 20.400 460.050 21.450 514.950 ;
        RECT 482.400 511.050 483.450 526.950 ;
        RECT 491.400 526.200 492.600 526.950 ;
        RECT 481.950 508.950 484.050 511.050 ;
        RECT 490.950 508.950 493.050 511.050 ;
        RECT 491.400 496.050 492.450 508.950 ;
        RECT 490.950 493.950 493.050 496.050 ;
        RECT 494.400 490.050 495.600 490.800 ;
        RECT 493.950 487.950 496.050 490.050 ;
        RECT 424.950 484.950 427.050 487.050 ;
        RECT 439.950 484.950 442.050 487.050 ;
        RECT 148.950 475.950 151.050 478.050 ;
        RECT 217.950 475.950 220.050 478.050 ;
        RECT 67.950 460.950 70.050 463.050 ;
        RECT 88.950 460.950 91.050 463.050 ;
        RECT 19.950 457.950 22.050 460.050 ;
        RECT 55.950 454.950 58.050 460.050 ;
        RECT 68.400 457.050 69.450 460.950 ;
        RECT 89.400 457.050 90.450 460.950 ;
        RECT 149.400 460.050 150.450 475.950 ;
        RECT 148.950 457.950 151.050 460.050 ;
        RECT 67.950 454.950 70.050 457.050 ;
        RECT 88.950 454.950 91.050 457.050 ;
        RECT 218.400 451.050 219.450 475.950 ;
        RECT 425.400 469.050 426.450 484.950 ;
        RECT 440.400 481.050 441.450 484.950 ;
        RECT 439.950 478.950 442.050 481.050 ;
        RECT 469.950 478.950 472.050 481.050 ;
        RECT 391.950 466.950 394.050 469.050 ;
        RECT 424.950 466.950 427.050 469.050 ;
        RECT 217.950 448.950 220.050 451.050 ;
        RECT 392.400 450.450 393.450 466.950 ;
        RECT 470.400 466.050 471.450 478.950 ;
        RECT 494.400 466.050 495.450 487.950 ;
        RECT 469.950 463.950 472.050 466.050 ;
        RECT 493.950 463.950 496.050 466.050 ;
        RECT 389.400 449.400 393.450 450.450 ;
        RECT 217.950 442.950 220.050 445.050 ;
        RECT 218.400 427.050 219.450 442.950 ;
        RECT 244.950 439.950 247.050 442.050 ;
        RECT 286.950 439.950 289.050 442.050 ;
        RECT 245.400 427.050 246.450 439.950 ;
        RECT 287.400 427.050 288.450 439.950 ;
        RECT 389.400 436.050 390.450 449.400 ;
        RECT 346.950 433.950 349.050 436.050 ;
        RECT 388.950 433.950 391.050 436.050 ;
        RECT 217.950 424.950 220.050 427.050 ;
        RECT 244.950 424.950 247.050 427.050 ;
        RECT 286.950 424.950 289.050 427.050 ;
        RECT 316.950 426.450 321.000 427.050 ;
        RECT 316.950 426.000 321.450 426.450 ;
        RECT 316.950 424.950 322.050 426.000 ;
        RECT 319.950 421.950 322.050 424.950 ;
        RECT 347.400 424.050 348.450 433.950 ;
        RECT 346.950 421.950 349.050 424.050 ;
      LAYER metal3 ;
        RECT 7.950 534.600 10.050 535.050 ;
        RECT -3.600 533.400 10.050 534.600 ;
        RECT 7.950 532.950 10.050 533.400 ;
        RECT 481.950 528.600 484.050 529.050 ;
        RECT 490.950 528.600 493.050 529.050 ;
        RECT 481.950 527.400 493.050 528.600 ;
        RECT 481.950 526.950 484.050 527.400 ;
        RECT 490.950 526.950 493.050 527.400 ;
        RECT 7.950 516.600 10.050 517.050 ;
        RECT 19.950 516.600 22.050 517.050 ;
        RECT 7.950 515.400 22.050 516.600 ;
        RECT 7.950 514.950 10.050 515.400 ;
        RECT 19.950 514.950 22.050 515.400 ;
        RECT 481.950 510.600 484.050 511.050 ;
        RECT 490.950 510.600 493.050 511.050 ;
        RECT 481.950 509.400 493.050 510.600 ;
        RECT 481.950 508.950 484.050 509.400 ;
        RECT 490.950 508.950 493.050 509.400 ;
        RECT 490.950 492.600 493.050 496.050 ;
        RECT 490.950 492.000 495.600 492.600 ;
        RECT 491.400 491.400 496.050 492.000 ;
        RECT 493.950 487.950 496.050 491.400 ;
        RECT 439.950 480.600 442.050 481.050 ;
        RECT 469.950 480.600 472.050 481.050 ;
        RECT 439.950 479.400 472.050 480.600 ;
        RECT 439.950 478.950 442.050 479.400 ;
        RECT 469.950 478.950 472.050 479.400 ;
        RECT 148.950 477.600 151.050 478.050 ;
        RECT 217.950 477.600 220.050 478.050 ;
        RECT 148.950 476.400 220.050 477.600 ;
        RECT 148.950 475.950 151.050 476.400 ;
        RECT 217.950 475.950 220.050 476.400 ;
        RECT 391.950 468.600 394.050 469.050 ;
        RECT 424.950 468.600 427.050 469.050 ;
        RECT 391.950 467.400 427.050 468.600 ;
        RECT 391.950 466.950 394.050 467.400 ;
        RECT 424.950 466.950 427.050 467.400 ;
        RECT 469.950 465.600 472.050 466.050 ;
        RECT 493.950 465.600 496.050 466.050 ;
        RECT 469.950 464.400 496.050 465.600 ;
        RECT 469.950 463.950 472.050 464.400 ;
        RECT 493.950 463.950 496.050 464.400 ;
        RECT 67.950 462.600 70.050 463.050 ;
        RECT 88.950 462.600 91.050 463.050 ;
        RECT 67.950 461.400 91.050 462.600 ;
        RECT 67.950 460.950 70.050 461.400 ;
        RECT 88.950 460.950 91.050 461.400 ;
        RECT 19.950 459.600 22.050 460.050 ;
        RECT 55.950 459.600 58.050 460.050 ;
        RECT 148.950 459.600 151.050 460.050 ;
        RECT 19.950 458.400 58.050 459.600 ;
        RECT 19.950 457.950 22.050 458.400 ;
        RECT 55.950 457.950 58.050 458.400 ;
        RECT 113.400 458.400 151.050 459.600 ;
        RECT 88.950 456.600 91.050 457.050 ;
        RECT 113.400 456.600 114.600 458.400 ;
        RECT 148.950 457.950 151.050 458.400 ;
        RECT 88.950 455.400 114.600 456.600 ;
        RECT 88.950 454.950 91.050 455.400 ;
        RECT 244.950 441.600 247.050 442.050 ;
        RECT 286.950 441.600 289.050 442.050 ;
        RECT 244.950 440.400 289.050 441.600 ;
        RECT 244.950 439.950 247.050 440.400 ;
        RECT 286.950 439.950 289.050 440.400 ;
        RECT 346.950 435.600 349.050 436.050 ;
        RECT 388.950 435.600 391.050 436.050 ;
        RECT 346.950 434.400 391.050 435.600 ;
        RECT 346.950 433.950 349.050 434.400 ;
        RECT 388.950 433.950 391.050 434.400 ;
        RECT 217.950 426.600 220.050 427.050 ;
        RECT 244.950 426.600 247.050 427.050 ;
        RECT 217.950 425.400 247.050 426.600 ;
        RECT 217.950 424.950 220.050 425.400 ;
        RECT 244.950 424.950 247.050 425.400 ;
        RECT 286.950 426.600 289.050 427.050 ;
        RECT 316.950 426.600 319.050 427.050 ;
        RECT 286.950 425.400 319.050 426.600 ;
        RECT 286.950 424.950 289.050 425.400 ;
        RECT 316.950 424.950 319.050 425.400 ;
        RECT 319.950 423.600 322.050 424.050 ;
        RECT 346.950 423.600 349.050 424.050 ;
        RECT 319.950 422.400 349.050 423.600 ;
        RECT 319.950 421.950 322.050 422.400 ;
        RECT 346.950 421.950 349.050 422.400 ;
    END
  END Xin[3]
  PIN Xin[2]
    PORT
      LAYER metal1 ;
        RECT 292.950 483.450 295.050 483.900 ;
        RECT 301.950 483.450 304.050 484.050 ;
        RECT 292.950 482.550 304.050 483.450 ;
        RECT 292.950 481.800 295.050 482.550 ;
        RECT 301.950 481.950 304.050 482.550 ;
      LAYER metal2 ;
        RECT 466.950 562.950 469.050 565.050 ;
        RECT 493.950 562.950 496.050 565.050 ;
        RECT 467.400 559.050 468.450 562.950 ;
        RECT 454.950 556.800 457.050 558.900 ;
        RECT 466.950 556.950 469.050 559.050 ;
        RECT 455.400 547.050 456.450 556.800 ;
        RECT 439.950 544.950 442.050 547.050 ;
        RECT 454.950 544.950 457.050 547.050 ;
        RECT 440.400 529.050 441.450 544.950 ;
        RECT 494.400 538.050 495.450 562.950 ;
        RECT 493.950 535.950 496.050 538.050 ;
        RECT 526.950 535.950 529.050 538.050 ;
        RECT 4.950 526.950 7.050 529.050 ;
        RECT 437.400 528.450 438.600 528.600 ;
        RECT 439.950 528.450 442.050 529.050 ;
        RECT 437.400 527.400 442.050 528.450 ;
        RECT 5.400 505.050 6.450 526.950 ;
        RECT 437.400 526.200 438.600 527.400 ;
        RECT 439.950 526.950 442.050 527.400 ;
        RECT 527.400 528.600 528.450 535.950 ;
        RECT 527.400 526.200 528.600 528.600 ;
        RECT 439.950 520.950 442.050 523.050 ;
        RECT 440.400 508.050 441.450 520.950 ;
        RECT 433.950 505.950 436.050 508.050 ;
        RECT 439.950 505.950 442.050 508.050 ;
        RECT 4.950 502.950 7.050 505.050 ;
        RECT 55.950 502.950 58.050 505.050 ;
        RECT 56.400 469.050 57.450 502.950 ;
        RECT 434.400 496.050 435.450 505.950 ;
        RECT 433.950 493.950 436.050 496.050 ;
        RECT 433.950 487.950 436.050 490.050 ;
        RECT 106.950 478.950 109.050 481.050 ;
        RECT 145.950 478.950 148.050 481.050 ;
        RECT 253.950 478.950 256.050 481.050 ;
        RECT 292.950 478.950 295.050 483.900 ;
        RECT 301.950 481.950 304.050 484.050 ;
        RECT 107.400 469.050 108.450 478.950 ;
        RECT 146.400 469.050 147.450 478.950 ;
        RECT 254.400 469.050 255.450 478.950 ;
        RECT 302.400 469.050 303.450 481.950 ;
        RECT 55.950 466.950 58.050 469.050 ;
        RECT 106.950 466.950 109.050 469.050 ;
        RECT 145.950 466.950 148.050 469.050 ;
        RECT 253.950 466.950 256.050 469.050 ;
        RECT 301.950 466.950 304.050 469.050 ;
        RECT 310.950 466.950 313.050 469.050 ;
        RECT 311.400 460.050 312.450 466.950 ;
        RECT 310.950 457.950 313.050 460.050 ;
        RECT 434.400 457.050 435.450 487.950 ;
        RECT 433.950 454.950 436.050 457.050 ;
      LAYER metal3 ;
        RECT 466.950 564.600 469.050 565.050 ;
        RECT 493.950 564.600 496.050 565.050 ;
        RECT 466.950 563.400 496.050 564.600 ;
        RECT 466.950 562.950 469.050 563.400 ;
        RECT 493.950 562.950 496.050 563.400 ;
        RECT 454.950 558.600 457.050 558.900 ;
        RECT 466.950 558.600 469.050 559.050 ;
        RECT 454.950 557.400 469.050 558.600 ;
        RECT 454.950 556.800 457.050 557.400 ;
        RECT 466.950 556.950 469.050 557.400 ;
        RECT 439.950 546.600 442.050 547.050 ;
        RECT 454.950 546.600 457.050 547.050 ;
        RECT 439.950 545.400 457.050 546.600 ;
        RECT 439.950 544.950 442.050 545.400 ;
        RECT 454.950 544.950 457.050 545.400 ;
        RECT 493.950 537.600 496.050 538.050 ;
        RECT 526.950 537.600 529.050 538.050 ;
        RECT 493.950 536.400 529.050 537.600 ;
        RECT 493.950 535.950 496.050 536.400 ;
        RECT 526.950 535.950 529.050 536.400 ;
        RECT 4.950 528.600 7.050 529.050 ;
        RECT -3.600 527.400 7.050 528.600 ;
        RECT 4.950 526.950 7.050 527.400 ;
        RECT 439.950 526.950 442.050 529.050 ;
        RECT 440.400 523.050 441.600 526.950 ;
        RECT 439.950 520.950 442.050 523.050 ;
        RECT 433.950 507.600 436.050 508.050 ;
        RECT 439.950 507.600 442.050 508.050 ;
        RECT 433.950 506.400 442.050 507.600 ;
        RECT 433.950 505.950 436.050 506.400 ;
        RECT 439.950 505.950 442.050 506.400 ;
        RECT 4.950 504.600 7.050 505.050 ;
        RECT 55.950 504.600 58.050 505.050 ;
        RECT 4.950 503.400 58.050 504.600 ;
        RECT 4.950 502.950 7.050 503.400 ;
        RECT 55.950 502.950 58.050 503.400 ;
        RECT 433.950 493.950 436.050 496.050 ;
        RECT 434.400 490.050 435.600 493.950 ;
        RECT 433.950 487.950 436.050 490.050 ;
        RECT 106.950 480.600 109.050 481.050 ;
        RECT 145.950 480.600 148.050 481.050 ;
        RECT 106.950 479.400 148.050 480.600 ;
        RECT 106.950 478.950 109.050 479.400 ;
        RECT 145.950 478.950 148.050 479.400 ;
        RECT 253.950 480.600 256.050 481.050 ;
        RECT 292.950 480.600 295.050 481.050 ;
        RECT 253.950 479.400 295.050 480.600 ;
        RECT 253.950 478.950 256.050 479.400 ;
        RECT 292.950 478.950 295.050 479.400 ;
        RECT 55.950 468.600 58.050 469.050 ;
        RECT 106.950 468.600 109.050 469.050 ;
        RECT 55.950 467.400 109.050 468.600 ;
        RECT 55.950 466.950 58.050 467.400 ;
        RECT 106.950 466.950 109.050 467.400 ;
        RECT 145.950 468.600 148.050 469.050 ;
        RECT 253.950 468.600 256.050 469.050 ;
        RECT 145.950 467.400 256.050 468.600 ;
        RECT 145.950 466.950 148.050 467.400 ;
        RECT 253.950 466.950 256.050 467.400 ;
        RECT 301.950 468.600 304.050 469.050 ;
        RECT 310.950 468.600 313.050 469.050 ;
        RECT 301.950 467.400 313.050 468.600 ;
        RECT 301.950 466.950 304.050 467.400 ;
        RECT 310.950 466.950 313.050 467.400 ;
        RECT 310.950 459.600 313.050 460.050 ;
        RECT 310.950 458.400 393.600 459.600 ;
        RECT 310.950 457.950 313.050 458.400 ;
        RECT 392.400 456.600 393.600 458.400 ;
        RECT 433.950 456.600 436.050 457.050 ;
        RECT 392.400 455.400 436.050 456.600 ;
        RECT 433.950 454.950 436.050 455.400 ;
    END
  END Xin[2]
  PIN Xin[1]
    PORT
      LAYER metal1 ;
        RECT 91.950 486.450 94.050 487.050 ;
        RECT 103.950 486.450 106.050 487.050 ;
        RECT 91.950 485.550 106.050 486.450 ;
        RECT 91.950 484.950 94.050 485.550 ;
        RECT 103.950 484.950 106.050 485.550 ;
      LAYER metal2 ;
        RECT 391.950 528.000 394.050 531.900 ;
        RECT 392.400 526.200 393.600 528.000 ;
        RECT 400.950 520.950 403.050 523.050 ;
        RECT 401.400 511.050 402.450 520.950 ;
        RECT 334.950 508.800 337.050 510.900 ;
        RECT 400.950 508.950 403.050 511.050 ;
        RECT 335.400 496.050 336.450 508.800 ;
        RECT 334.950 493.950 337.050 496.050 ;
        RECT 91.950 484.950 94.050 487.050 ;
        RECT 92.400 472.050 93.450 484.950 ;
        RECT 103.950 481.950 106.050 487.050 ;
        RECT 325.950 484.950 328.050 487.050 ;
        RECT 193.950 481.950 196.050 484.050 ;
        RECT 43.950 469.950 46.050 472.050 ;
        RECT 91.950 469.950 94.050 472.050 ;
        RECT 44.400 466.050 45.450 469.950 ;
        RECT 1.950 463.950 4.050 466.050 ;
        RECT 43.950 463.950 46.050 466.050 ;
        RECT 2.400 457.050 3.450 463.950 ;
        RECT 194.400 457.050 195.450 481.950 ;
        RECT 326.400 463.050 327.450 484.950 ;
        RECT 295.950 460.050 298.050 463.050 ;
        RECT 325.950 460.950 328.050 463.050 ;
        RECT 346.950 460.950 349.050 463.050 ;
        RECT 292.950 459.000 298.050 460.050 ;
        RECT 292.950 458.400 297.450 459.000 ;
        RECT 292.950 457.950 297.000 458.400 ;
        RECT 1.950 454.950 4.050 457.050 ;
        RECT 193.950 454.950 196.050 457.050 ;
        RECT 347.400 450.600 348.450 460.950 ;
        RECT 347.400 448.200 348.600 450.600 ;
      LAYER metal3 ;
        RECT 391.950 531.600 394.050 531.900 ;
        RECT 391.950 530.400 405.600 531.600 ;
        RECT 391.950 529.800 394.050 530.400 ;
        RECT 404.400 523.050 405.600 530.400 ;
        RECT 400.950 521.400 405.600 523.050 ;
        RECT 400.950 520.950 405.000 521.400 ;
        RECT 334.950 510.600 337.050 510.900 ;
        RECT 400.950 510.600 403.050 511.050 ;
        RECT 334.950 509.400 403.050 510.600 ;
        RECT 334.950 508.800 337.050 509.400 ;
        RECT 400.950 508.950 403.050 509.400 ;
        RECT 334.950 493.950 337.050 496.050 ;
        RECT 335.400 489.600 336.600 493.950 ;
        RECT 326.400 489.000 336.600 489.600 ;
        RECT 325.950 488.400 336.600 489.000 ;
        RECT 325.950 484.950 328.050 488.400 ;
        RECT 103.950 483.600 106.050 484.050 ;
        RECT 193.950 483.600 196.050 484.050 ;
        RECT 103.950 482.400 196.050 483.600 ;
        RECT 103.950 481.950 106.050 482.400 ;
        RECT 193.950 481.950 196.050 482.400 ;
        RECT 43.950 471.600 46.050 472.050 ;
        RECT 91.950 471.600 94.050 472.050 ;
        RECT 43.950 470.400 94.050 471.600 ;
        RECT 43.950 469.950 46.050 470.400 ;
        RECT 91.950 469.950 94.050 470.400 ;
        RECT 1.950 465.600 4.050 466.050 ;
        RECT 43.950 465.600 46.050 466.050 ;
        RECT 1.950 464.400 46.050 465.600 ;
        RECT 1.950 463.950 4.050 464.400 ;
        RECT 43.950 463.950 46.050 464.400 ;
        RECT 295.950 462.600 298.050 463.050 ;
        RECT 325.950 462.600 328.050 463.050 ;
        RECT 346.950 462.600 349.050 463.050 ;
        RECT 295.950 461.400 349.050 462.600 ;
        RECT 295.950 460.950 298.050 461.400 ;
        RECT 325.950 460.950 328.050 461.400 ;
        RECT 346.950 460.950 349.050 461.400 ;
        RECT 292.950 459.600 295.050 460.050 ;
        RECT 224.400 458.400 295.050 459.600 ;
        RECT 1.950 456.600 4.050 457.050 ;
        RECT -3.600 455.400 4.050 456.600 ;
        RECT 1.950 454.950 4.050 455.400 ;
        RECT 193.950 456.600 196.050 457.050 ;
        RECT 224.400 456.600 225.600 458.400 ;
        RECT 292.950 457.950 295.050 458.400 ;
        RECT 193.950 455.400 225.600 456.600 ;
        RECT 193.950 454.950 196.050 455.400 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal2 ;
        RECT 1.950 448.950 4.050 451.050 ;
        RECT 418.950 448.950 421.050 451.050 ;
        RECT 424.950 448.950 427.050 451.050 ;
        RECT 430.950 448.950 433.050 451.050 ;
        RECT 2.400 397.050 3.450 448.950 ;
        RECT 419.400 448.200 420.600 448.950 ;
        RECT 425.400 430.050 426.450 448.950 ;
        RECT 431.400 448.200 432.600 448.950 ;
        RECT 424.950 427.950 427.050 430.050 ;
        RECT 436.950 427.950 439.050 430.050 ;
        RECT 143.400 401.400 150.450 402.450 ;
        RECT 143.400 397.050 144.450 401.400 ;
        RECT 1.950 394.950 4.050 397.050 ;
        RECT 139.950 395.400 144.450 397.050 ;
        RECT 139.950 394.950 144.000 395.400 ;
        RECT 149.400 385.050 150.450 401.400 ;
        RECT 437.400 400.050 438.450 427.950 ;
        RECT 379.950 397.950 382.050 400.050 ;
        RECT 436.950 397.950 439.050 400.050 ;
        RECT 166.950 394.950 169.050 397.050 ;
        RECT 181.950 394.950 184.050 397.050 ;
        RECT 167.400 385.050 168.450 394.950 ;
        RECT 182.400 385.050 183.450 394.950 ;
        RECT 380.400 385.050 381.450 397.950 ;
        RECT 148.950 382.950 151.050 385.050 ;
        RECT 166.950 382.950 169.050 385.050 ;
        RECT 181.950 382.950 184.050 385.050 ;
        RECT 379.950 382.950 382.050 385.050 ;
      LAYER metal3 ;
        RECT 1.950 450.600 4.050 451.050 ;
        RECT -3.600 449.400 4.050 450.600 ;
        RECT 1.950 448.950 4.050 449.400 ;
        RECT 418.950 450.600 421.050 451.050 ;
        RECT 424.950 450.600 427.050 451.050 ;
        RECT 430.950 450.600 433.050 451.050 ;
        RECT 418.950 449.400 433.050 450.600 ;
        RECT 418.950 448.950 421.050 449.400 ;
        RECT 424.950 448.950 427.050 449.400 ;
        RECT 430.950 448.950 433.050 449.400 ;
        RECT 424.950 429.600 427.050 430.050 ;
        RECT 436.950 429.600 439.050 430.050 ;
        RECT 424.950 428.400 439.050 429.600 ;
        RECT 424.950 427.950 427.050 428.400 ;
        RECT 436.950 427.950 439.050 428.400 ;
        RECT 379.950 399.600 382.050 400.050 ;
        RECT 436.950 399.600 439.050 400.050 ;
        RECT 379.950 398.400 439.050 399.600 ;
        RECT 379.950 397.950 382.050 398.400 ;
        RECT 436.950 397.950 439.050 398.400 ;
        RECT 1.950 396.600 4.050 397.050 ;
        RECT 139.950 396.600 142.050 397.050 ;
        RECT 1.950 395.400 142.050 396.600 ;
        RECT 1.950 394.950 4.050 395.400 ;
        RECT 139.950 394.950 142.050 395.400 ;
        RECT 166.950 396.600 169.050 397.050 ;
        RECT 181.950 396.600 184.050 397.050 ;
        RECT 166.950 395.400 184.050 396.600 ;
        RECT 166.950 394.950 169.050 395.400 ;
        RECT 181.950 394.950 184.050 395.400 ;
        RECT 148.950 384.600 151.050 385.050 ;
        RECT 166.950 384.600 169.050 385.050 ;
        RECT 148.950 383.400 169.050 384.600 ;
        RECT 148.950 382.950 151.050 383.400 ;
        RECT 166.950 382.950 169.050 383.400 ;
        RECT 181.950 384.600 184.050 385.050 ;
        RECT 379.950 384.600 382.050 385.050 ;
        RECT 181.950 383.400 382.050 384.600 ;
        RECT 181.950 382.950 184.050 383.400 ;
        RECT 379.950 382.950 382.050 383.400 ;
    END
  END Xin[0]
  PIN Xout[3]
    PORT
      LAYER metal2 ;
        RECT 817.950 606.000 820.050 610.050 ;
        RECT 818.400 604.350 819.600 606.000 ;
      LAYER metal3 ;
        RECT 830.400 611.400 870.600 612.600 ;
        RECT 817.950 609.600 820.050 610.050 ;
        RECT 830.400 609.600 831.600 611.400 ;
        RECT 817.950 608.400 831.600 609.600 ;
        RECT 817.950 607.950 820.050 608.400 ;
    END
  END Xout[3]
  PIN Xout[2]
    PORT
      LAYER metal2 ;
        RECT 853.950 605.100 856.050 607.200 ;
        RECT 854.400 604.350 855.600 605.100 ;
      LAYER metal3 ;
        RECT 853.950 606.600 856.050 607.200 ;
        RECT 853.950 605.400 870.600 606.600 ;
        RECT 853.950 605.100 856.050 605.400 ;
    END
  END Xout[2]
  PIN Xout[1]
    PORT
      LAYER metal2 ;
        RECT 824.400 568.050 825.600 568.650 ;
        RECT 824.400 566.400 829.050 568.050 ;
        RECT 825.000 565.950 829.050 566.400 ;
      LAYER metal3 ;
        RECT 826.950 567.600 829.050 568.050 ;
        RECT 826.950 566.400 870.600 567.600 ;
        RECT 826.950 565.950 829.050 566.400 ;
    END
  END Xout[1]
  PIN Xout[0]
    PORT
      LAYER metal2 ;
        RECT 817.950 449.100 820.050 451.200 ;
        RECT 818.400 448.350 819.600 449.100 ;
      LAYER metal3 ;
        RECT 817.950 450.600 820.050 451.200 ;
        RECT 817.950 449.400 870.600 450.600 ;
        RECT 817.950 449.100 820.050 449.400 ;
    END
  END Xout[0]
  PIN Yin[3]
    PORT
      LAYER metal1 ;
        RECT 487.950 27.450 492.000 28.050 ;
        RECT 487.950 25.950 492.450 27.450 ;
        RECT 491.550 22.050 492.450 25.950 ;
        RECT 491.550 20.550 496.050 22.050 ;
        RECT 492.000 19.950 496.050 20.550 ;
        RECT 505.950 6.450 508.050 7.050 ;
        RECT 511.950 6.450 514.050 7.050 ;
        RECT 505.950 5.550 514.050 6.450 ;
        RECT 505.950 4.950 508.050 5.550 ;
        RECT 511.950 4.950 514.050 5.550 ;
      LAYER metal2 ;
        RECT 486.000 27.600 490.050 28.050 ;
        RECT 485.400 25.950 490.050 27.600 ;
        RECT 485.400 25.350 486.600 25.950 ;
        RECT 493.950 19.950 496.050 22.050 ;
        RECT 494.400 0.450 495.450 19.950 ;
        RECT 504.000 6.450 508.050 7.050 ;
        RECT 503.400 4.950 508.050 6.450 ;
        RECT 511.950 4.950 514.050 7.050 ;
        RECT 503.400 0.450 504.450 4.950 ;
        RECT 494.400 -0.600 504.450 0.450 ;
        RECT 512.400 -2.550 513.450 4.950 ;
        RECT 512.400 -3.600 516.450 -2.550 ;
    END
  END Yin[3]
  PIN Yin[2]
    PORT
      LAYER metal2 ;
        RECT 515.400 53.400 516.600 55.650 ;
        RECT 515.400 43.050 516.450 53.400 ;
        RECT 493.950 40.950 496.050 43.050 ;
        RECT 514.950 40.950 517.050 43.050 ;
        RECT 494.400 28.050 495.450 40.950 ;
        RECT 493.950 25.950 496.050 28.050 ;
        RECT 499.950 19.950 502.050 22.050 ;
        RECT 500.400 4.050 501.450 19.950 ;
        RECT 499.950 1.950 502.050 4.050 ;
        RECT 508.950 1.950 511.050 4.050 ;
        RECT 509.400 -3.600 510.450 1.950 ;
      LAYER metal3 ;
        RECT 493.950 42.600 496.050 43.050 ;
        RECT 514.950 42.600 517.050 43.050 ;
        RECT 493.950 41.400 517.050 42.600 ;
        RECT 493.950 40.950 496.050 41.400 ;
        RECT 514.950 40.950 517.050 41.400 ;
        RECT 493.950 24.600 496.050 28.050 ;
        RECT 493.950 24.000 501.600 24.600 ;
        RECT 494.400 23.400 502.050 24.000 ;
        RECT 499.950 19.950 502.050 23.400 ;
        RECT 499.950 3.600 502.050 4.050 ;
        RECT 508.950 3.600 511.050 4.050 ;
        RECT 499.950 2.400 511.050 3.600 ;
        RECT 499.950 1.950 502.050 2.400 ;
        RECT 508.950 1.950 511.050 2.400 ;
    END
  END Yin[2]
  PIN Yin[1]
    PORT
      LAYER metal2 ;
        RECT 377.400 27.450 378.600 27.600 ;
        RECT 377.400 26.400 384.450 27.450 ;
        RECT 377.400 25.350 378.600 26.400 ;
        RECT 383.400 4.050 384.450 26.400 ;
        RECT 373.950 1.950 376.050 4.050 ;
        RECT 382.950 1.950 385.050 4.050 ;
        RECT 374.400 -3.600 375.450 1.950 ;
      LAYER metal3 ;
        RECT 373.950 3.600 376.050 4.050 ;
        RECT 382.950 3.600 385.050 4.050 ;
        RECT 373.950 2.400 385.050 3.600 ;
        RECT 373.950 1.950 376.050 2.400 ;
        RECT 382.950 1.950 385.050 2.400 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal2 ;
        RECT 355.950 26.100 358.050 28.200 ;
        RECT 356.400 25.350 357.600 26.100 ;
        RECT 352.950 19.950 355.050 22.050 ;
        RECT 353.400 4.050 354.450 19.950 ;
        RECT 352.950 1.950 355.050 4.050 ;
        RECT 358.950 1.950 361.050 4.050 ;
        RECT 359.400 -3.600 360.450 1.950 ;
      LAYER metal3 ;
        RECT 355.950 27.600 358.050 28.200 ;
        RECT 353.400 26.400 358.050 27.600 ;
        RECT 353.400 22.050 354.600 26.400 ;
        RECT 355.950 26.100 358.050 26.400 ;
        RECT 352.950 19.950 355.050 22.050 ;
        RECT 352.950 3.600 355.050 4.050 ;
        RECT 358.950 3.600 361.050 4.050 ;
        RECT 352.950 2.400 361.050 3.600 ;
        RECT 352.950 1.950 355.050 2.400 ;
        RECT 358.950 1.950 361.050 2.400 ;
    END
  END Yin[0]
  PIN Yout[3]
    PORT
      LAYER metal2 ;
        RECT 638.400 98.400 639.600 100.650 ;
        RECT 638.400 73.050 639.450 98.400 ;
        RECT 628.950 70.950 631.050 73.050 ;
        RECT 637.950 70.950 640.050 73.050 ;
        RECT 629.400 61.050 630.450 70.950 ;
        RECT 628.950 58.950 631.050 61.050 ;
        RECT 628.950 52.950 631.050 55.050 ;
        RECT 629.400 39.450 630.450 52.950 ;
        RECT 623.400 38.400 630.450 39.450 ;
        RECT 623.400 7.050 624.450 38.400 ;
        RECT 622.950 4.950 625.050 7.050 ;
        RECT 658.950 4.950 661.050 7.050 ;
        RECT 659.400 -3.600 660.450 4.950 ;
      LAYER metal3 ;
        RECT 628.950 72.600 631.050 73.050 ;
        RECT 637.950 72.600 640.050 73.050 ;
        RECT 628.950 71.400 640.050 72.600 ;
        RECT 628.950 70.950 631.050 71.400 ;
        RECT 637.950 70.950 640.050 71.400 ;
        RECT 628.950 58.950 631.050 61.050 ;
        RECT 629.400 55.050 630.600 58.950 ;
        RECT 628.950 52.950 631.050 55.050 ;
        RECT 622.950 6.600 625.050 7.050 ;
        RECT 658.950 6.600 661.050 7.050 ;
        RECT 622.950 5.400 661.050 6.600 ;
        RECT 622.950 4.950 625.050 5.400 ;
        RECT 658.950 4.950 661.050 5.400 ;
    END
  END Yout[3]
  PIN Yout[2]
    PORT
      LAYER metal1 ;
        RECT 637.950 63.450 640.050 64.050 ;
        RECT 632.550 62.550 640.050 63.450 ;
        RECT 632.550 54.450 633.450 62.550 ;
        RECT 637.950 61.950 640.050 62.550 ;
        RECT 632.550 53.550 636.450 54.450 ;
        RECT 635.550 51.450 636.450 53.550 ;
        RECT 635.550 51.000 639.450 51.450 ;
        RECT 635.550 50.550 640.050 51.000 ;
        RECT 637.950 46.800 640.050 50.550 ;
      LAYER metal2 ;
        RECT 637.950 61.950 640.050 67.050 ;
        RECT 658.950 64.950 661.050 67.050 ;
        RECT 659.400 60.600 660.450 64.950 ;
        RECT 659.400 58.350 660.600 60.600 ;
        RECT 637.950 46.800 640.050 48.900 ;
        RECT 638.400 4.050 639.450 46.800 ;
        RECT 637.950 1.950 640.050 4.050 ;
        RECT 652.950 1.950 655.050 4.050 ;
        RECT 653.400 -3.600 654.450 1.950 ;
      LAYER metal3 ;
        RECT 637.950 66.600 640.050 67.050 ;
        RECT 658.950 66.600 661.050 67.050 ;
        RECT 637.950 65.400 661.050 66.600 ;
        RECT 637.950 64.950 640.050 65.400 ;
        RECT 658.950 64.950 661.050 65.400 ;
        RECT 637.950 3.600 640.050 4.050 ;
        RECT 652.950 3.600 655.050 4.050 ;
        RECT 637.950 2.400 655.050 3.600 ;
        RECT 637.950 1.950 640.050 2.400 ;
        RECT 652.950 1.950 655.050 2.400 ;
    END
  END Yout[2]
  PIN Yout[1]
    PORT
      LAYER metal2 ;
        RECT 650.400 20.400 651.600 22.650 ;
        RECT 650.400 -2.550 651.450 20.400 ;
        RECT 647.400 -3.600 651.450 -2.550 ;
    END
  END Yout[1]
  PIN Yout[0]
    PORT
      LAYER metal1 ;
        RECT 619.950 63.450 622.050 64.050 ;
        RECT 614.550 62.550 622.050 63.450 ;
        RECT 614.550 55.050 615.450 62.550 ;
        RECT 619.950 61.950 622.050 62.550 ;
        RECT 614.550 53.550 619.050 55.050 ;
        RECT 615.000 52.950 619.050 53.550 ;
      LAYER metal2 ;
        RECT 620.400 98.400 621.600 100.650 ;
        RECT 620.400 64.050 621.450 98.400 ;
        RECT 619.950 61.950 622.050 64.050 ;
        RECT 616.950 52.950 619.050 55.050 ;
        RECT 617.400 27.450 618.450 52.950 ;
        RECT 617.400 26.400 621.450 27.450 ;
        RECT 620.400 -2.550 621.450 26.400 ;
        RECT 617.400 -3.600 621.450 -2.550 ;
    END
  END Yout[0]
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 478.950 816.450 481.050 817.050 ;
        RECT 487.950 816.450 490.050 817.050 ;
        RECT 478.950 815.550 490.050 816.450 ;
        RECT 478.950 814.950 481.050 815.550 ;
        RECT 487.950 814.950 490.050 815.550 ;
        RECT 457.950 810.450 460.050 811.050 ;
        RECT 472.950 810.450 475.050 811.050 ;
        RECT 457.950 809.550 475.050 810.450 ;
        RECT 457.950 808.950 460.050 809.550 ;
        RECT 472.950 808.950 475.050 809.550 ;
        RECT 517.950 528.450 522.000 529.050 ;
        RECT 517.950 526.950 522.450 528.450 ;
        RECT 521.550 519.450 522.450 526.950 ;
        RECT 526.950 519.450 529.050 520.050 ;
        RECT 521.550 518.550 529.050 519.450 ;
        RECT 526.950 517.950 529.050 518.550 ;
      LAYER metal2 ;
        RECT 488.400 827.400 492.450 828.450 ;
        RECT 488.400 817.050 489.450 827.400 ;
        RECT 478.950 816.450 481.050 817.050 ;
        RECT 473.400 815.400 481.050 816.450 ;
        RECT 473.400 811.050 474.450 815.400 ;
        RECT 478.950 814.950 481.050 815.400 ;
        RECT 487.950 814.950 490.050 817.050 ;
        RECT 457.950 805.950 460.050 811.050 ;
        RECT 472.950 808.950 475.050 811.050 ;
        RECT 442.950 796.950 445.050 799.050 ;
        RECT 443.400 733.050 444.450 796.950 ;
        RECT 442.950 730.950 445.050 733.050 ;
        RECT 439.950 721.950 442.050 724.050 ;
        RECT 440.400 685.050 441.450 721.950 ;
        RECT 439.950 682.950 442.050 685.050 ;
        RECT 430.950 673.950 433.050 676.050 ;
        RECT 431.400 645.450 432.450 673.950 ;
        RECT 428.400 644.400 432.450 645.450 ;
        RECT 428.400 577.050 429.450 644.400 ;
        RECT 427.950 574.950 430.050 577.050 ;
        RECT 481.950 565.950 484.050 568.050 ;
        RECT 482.400 544.050 483.450 565.950 ;
        RECT 481.950 541.950 484.050 544.050 ;
        RECT 517.950 541.950 520.050 544.050 ;
        RECT 518.400 529.050 519.450 541.950 ;
        RECT 517.950 526.950 520.050 529.050 ;
        RECT 526.950 517.950 529.050 520.050 ;
        RECT 527.400 496.050 528.450 517.950 ;
        RECT 526.950 493.950 529.050 496.050 ;
        RECT 526.800 487.950 528.900 490.050 ;
        RECT 527.400 484.050 528.450 487.950 ;
        RECT 526.950 481.950 529.050 484.050 ;
        RECT 538.950 481.950 541.050 484.050 ;
        RECT 539.400 442.050 540.450 481.950 ;
        RECT 532.950 439.950 535.050 442.050 ;
        RECT 538.950 439.950 541.050 442.050 ;
        RECT 503.400 412.050 504.600 412.800 ;
        RECT 518.400 412.050 519.600 412.800 ;
        RECT 533.400 412.050 534.450 439.950 ;
        RECT 502.950 409.950 505.050 412.050 ;
        RECT 517.950 411.450 520.050 412.050 ;
        RECT 517.950 410.400 522.450 411.450 ;
        RECT 517.950 409.950 520.050 410.400 ;
        RECT 521.400 361.050 522.450 410.400 ;
        RECT 532.950 409.950 535.050 412.050 ;
        RECT 478.950 358.950 481.050 361.050 ;
        RECT 520.950 358.950 523.050 361.050 ;
        RECT 479.400 301.050 480.450 358.950 ;
        RECT 427.950 298.950 430.050 301.050 ;
        RECT 478.950 298.950 481.050 301.050 ;
        RECT 508.950 298.950 511.050 301.050 ;
        RECT 428.400 286.050 429.450 298.950 ;
        RECT 509.400 294.600 510.450 298.950 ;
        RECT 509.400 292.200 510.600 294.600 ;
        RECT 421.950 283.650 424.050 285.750 ;
        RECT 427.950 283.950 430.050 286.050 ;
        RECT 143.400 254.400 144.600 256.800 ;
        RECT 143.400 229.050 144.450 254.400 ;
        RECT 422.400 253.050 423.450 283.650 ;
        RECT 166.950 250.950 169.050 253.050 ;
        RECT 421.950 250.950 424.050 253.050 ;
        RECT 430.950 250.950 433.050 253.050 ;
        RECT 167.400 229.050 168.450 250.950 ;
        RECT 142.950 226.950 145.050 229.050 ;
        RECT 166.950 226.950 169.050 229.050 ;
        RECT 167.400 178.050 168.450 226.950 ;
        RECT 431.400 220.050 432.450 250.950 ;
        RECT 430.950 217.950 433.050 220.050 ;
        RECT 469.950 217.950 472.050 220.050 ;
        RECT 176.400 178.050 177.600 178.800 ;
        RECT 464.400 178.050 465.600 178.800 ;
        RECT 470.400 178.050 471.450 217.950 ;
        RECT 478.950 216.000 481.050 220.050 ;
        RECT 479.400 214.200 480.600 216.000 ;
        RECT 166.950 175.950 169.050 178.050 ;
        RECT 175.950 175.950 178.050 178.050 ;
        RECT 463.950 175.950 466.050 178.050 ;
        RECT 469.950 175.950 472.050 178.050 ;
        RECT 575.400 176.400 576.600 178.800 ;
        RECT 470.400 169.050 471.450 175.950 ;
        RECT 575.400 169.050 576.450 176.400 ;
        RECT 469.950 166.950 472.050 169.050 ;
        RECT 574.950 166.950 577.050 169.050 ;
      LAYER metal3 ;
        RECT 457.950 805.950 460.050 808.050 ;
        RECT 442.950 798.600 445.050 799.050 ;
        RECT 458.400 798.600 459.600 805.950 ;
        RECT 442.950 797.400 459.600 798.600 ;
        RECT 442.950 796.950 445.050 797.400 ;
        RECT 442.950 730.950 445.050 733.050 ;
        RECT 443.400 726.600 444.600 730.950 ;
        RECT 440.400 726.000 444.600 726.600 ;
        RECT 439.950 725.400 444.600 726.000 ;
        RECT 439.950 721.950 442.050 725.400 ;
        RECT 439.950 681.600 442.050 685.050 ;
        RECT 439.950 681.000 453.600 681.600 ;
        RECT 440.400 680.400 453.600 681.000 ;
        RECT 430.950 675.600 433.050 676.050 ;
        RECT 452.400 675.600 453.600 680.400 ;
        RECT 430.950 674.400 453.600 675.600 ;
        RECT 430.950 673.950 433.050 674.400 ;
        RECT 427.950 576.600 432.000 577.050 ;
        RECT 427.950 574.950 432.600 576.600 ;
        RECT 431.400 570.600 432.600 574.950 ;
        RECT 431.400 569.400 471.600 570.600 ;
        RECT 470.400 567.600 471.600 569.400 ;
        RECT 481.950 567.600 484.050 568.050 ;
        RECT 470.400 566.400 484.050 567.600 ;
        RECT 481.950 565.950 484.050 566.400 ;
        RECT 481.950 543.600 484.050 544.050 ;
        RECT 517.950 543.600 520.050 544.050 ;
        RECT 481.950 542.400 520.050 543.600 ;
        RECT 481.950 541.950 484.050 542.400 ;
        RECT 517.950 541.950 520.050 542.400 ;
        RECT 526.950 493.950 529.050 496.050 ;
        RECT 527.400 490.050 528.600 493.950 ;
        RECT 526.800 487.950 528.900 490.050 ;
        RECT 526.950 483.600 529.050 484.050 ;
        RECT 538.950 483.600 541.050 484.050 ;
        RECT 526.950 482.400 541.050 483.600 ;
        RECT 526.950 481.950 529.050 482.400 ;
        RECT 538.950 481.950 541.050 482.400 ;
        RECT 532.950 441.600 535.050 442.050 ;
        RECT 538.950 441.600 541.050 442.050 ;
        RECT 532.950 440.400 541.050 441.600 ;
        RECT 532.950 439.950 535.050 440.400 ;
        RECT 538.950 439.950 541.050 440.400 ;
        RECT 502.950 411.600 505.050 412.050 ;
        RECT 517.950 411.600 520.050 412.050 ;
        RECT 532.950 411.600 535.050 412.050 ;
        RECT 502.950 410.400 535.050 411.600 ;
        RECT 502.950 409.950 505.050 410.400 ;
        RECT 517.950 409.950 520.050 410.400 ;
        RECT 532.950 409.950 535.050 410.400 ;
        RECT 478.950 360.600 481.050 361.050 ;
        RECT 520.950 360.600 523.050 361.050 ;
        RECT 478.950 359.400 523.050 360.600 ;
        RECT 478.950 358.950 481.050 359.400 ;
        RECT 520.950 358.950 523.050 359.400 ;
        RECT 427.950 300.600 430.050 301.050 ;
        RECT 478.950 300.600 481.050 301.050 ;
        RECT 508.950 300.600 511.050 301.050 ;
        RECT 427.950 299.400 511.050 300.600 ;
        RECT 427.950 298.950 430.050 299.400 ;
        RECT 478.950 298.950 481.050 299.400 ;
        RECT 508.950 298.950 511.050 299.400 ;
        RECT 421.950 285.600 424.050 285.750 ;
        RECT 427.950 285.600 430.050 286.050 ;
        RECT 421.950 284.400 430.050 285.600 ;
        RECT 421.950 283.650 424.050 284.400 ;
        RECT 427.950 283.950 430.050 284.400 ;
        RECT 166.950 252.600 169.050 253.050 ;
        RECT 421.950 252.600 424.050 253.050 ;
        RECT 430.950 252.600 433.050 253.050 ;
        RECT 166.950 251.400 433.050 252.600 ;
        RECT 166.950 250.950 169.050 251.400 ;
        RECT 421.950 250.950 424.050 251.400 ;
        RECT 430.950 250.950 433.050 251.400 ;
        RECT 142.950 228.600 145.050 229.050 ;
        RECT 166.950 228.600 169.050 229.050 ;
        RECT 142.950 227.400 169.050 228.600 ;
        RECT 142.950 226.950 145.050 227.400 ;
        RECT 166.950 226.950 169.050 227.400 ;
        RECT 430.950 219.600 433.050 220.050 ;
        RECT 469.950 219.600 472.050 220.050 ;
        RECT 478.950 219.600 481.050 220.050 ;
        RECT 430.950 218.400 481.050 219.600 ;
        RECT 430.950 217.950 433.050 218.400 ;
        RECT 469.950 217.950 472.050 218.400 ;
        RECT 478.950 217.950 481.050 218.400 ;
        RECT 166.950 177.600 169.050 178.050 ;
        RECT 175.950 177.600 178.050 178.050 ;
        RECT 166.950 176.400 178.050 177.600 ;
        RECT 166.950 175.950 169.050 176.400 ;
        RECT 175.950 175.950 178.050 176.400 ;
        RECT 463.950 177.600 466.050 178.050 ;
        RECT 469.950 177.600 472.050 178.050 ;
        RECT 463.950 176.400 472.050 177.600 ;
        RECT 463.950 175.950 466.050 176.400 ;
        RECT 469.950 175.950 472.050 176.400 ;
        RECT 469.950 168.600 472.050 169.050 ;
        RECT 574.950 168.600 577.050 169.050 ;
        RECT 469.950 167.400 577.050 168.600 ;
        RECT 469.950 166.950 472.050 167.400 ;
        RECT 574.950 166.950 577.050 167.400 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 11.700 815.400 13.500 819.000 ;
        RECT 14.700 813.600 16.500 818.400 ;
        RECT 11.400 812.400 16.500 813.600 ;
        RECT 19.200 812.400 21.000 819.000 ;
        RECT 11.400 805.200 12.300 812.400 ;
        RECT 29.400 809.400 31.200 819.000 ;
        RECT 36.000 810.000 37.800 818.400 ;
        RECT 55.200 810.000 57.000 818.400 ;
        RECT 36.000 808.800 39.300 810.000 ;
        RECT 14.100 805.200 15.900 807.000 ;
        RECT 20.100 805.200 21.900 807.000 ;
        RECT 29.100 805.200 30.900 807.000 ;
        RECT 35.100 805.200 36.900 807.000 ;
        RECT 38.400 805.200 39.300 808.800 ;
        RECT 53.700 808.800 57.000 810.000 ;
        RECT 61.800 809.400 63.600 819.000 ;
        RECT 71.700 812.400 73.500 819.000 ;
        RECT 76.800 811.200 78.600 818.400 ;
        RECT 74.400 810.300 78.600 811.200 ;
        RECT 49.950 807.450 52.050 808.050 ;
        RECT 44.550 806.550 52.050 807.450 ;
        RECT 10.950 803.100 13.050 805.200 ;
        RECT 13.950 803.100 16.050 805.200 ;
        RECT 16.950 803.100 19.050 805.200 ;
        RECT 19.950 803.100 22.050 805.200 ;
        RECT 28.950 803.100 31.050 805.200 ;
        RECT 31.950 803.100 34.050 805.200 ;
        RECT 34.950 803.100 37.050 805.200 ;
        RECT 37.950 803.100 40.050 805.200 ;
        RECT 11.400 795.600 12.300 803.100 ;
        RECT 17.100 801.300 18.900 803.100 ;
        RECT 32.100 801.300 33.900 803.100 ;
        RECT 16.950 798.450 19.050 799.050 ;
        RECT 34.950 798.450 37.050 799.050 ;
        RECT 16.950 797.550 37.050 798.450 ;
        RECT 16.950 796.950 19.050 797.550 ;
        RECT 34.950 796.950 37.050 797.550 ;
        RECT 10.800 783.600 12.600 795.600 ;
        RECT 13.800 794.700 21.600 795.600 ;
        RECT 13.800 783.600 15.600 794.700 ;
        RECT 16.800 783.000 18.600 793.800 ;
        RECT 19.800 783.600 21.600 794.700 ;
        RECT 38.400 790.800 39.300 803.100 ;
        RECT 44.550 801.450 45.450 806.550 ;
        RECT 49.950 805.950 52.050 806.550 ;
        RECT 53.700 805.200 54.600 808.800 ;
        RECT 56.100 805.200 57.900 807.000 ;
        RECT 62.100 805.200 63.900 807.000 ;
        RECT 71.100 805.200 72.900 807.000 ;
        RECT 74.400 805.200 75.600 810.300 ;
        RECT 94.200 810.000 96.000 818.400 ;
        RECT 92.700 808.800 96.000 810.000 ;
        RECT 100.800 809.400 102.600 819.000 ;
        RECT 110.700 812.400 112.500 819.000 ;
        RECT 115.800 811.200 117.600 818.400 ;
        RECT 128.400 815.400 130.200 819.000 ;
        RECT 131.400 815.400 133.200 818.400 ;
        RECT 134.400 815.400 136.200 819.000 ;
        RECT 113.400 810.300 117.600 811.200 ;
        RECT 77.100 805.200 78.900 807.000 ;
        RECT 92.700 805.200 93.600 808.800 ;
        RECT 95.100 805.200 96.900 807.000 ;
        RECT 101.100 805.200 102.900 807.000 ;
        RECT 110.100 805.200 111.900 807.000 ;
        RECT 113.400 805.200 114.600 810.300 ;
        RECT 116.100 805.200 117.900 807.000 ;
        RECT 52.950 803.100 55.050 805.200 ;
        RECT 55.950 803.100 58.050 805.200 ;
        RECT 58.950 803.100 61.050 805.200 ;
        RECT 61.950 803.100 64.050 805.200 ;
        RECT 70.950 803.100 73.050 805.200 ;
        RECT 73.950 803.100 76.050 805.200 ;
        RECT 76.950 803.100 79.050 805.200 ;
        RECT 91.950 803.100 94.050 805.200 ;
        RECT 94.950 803.100 97.050 805.200 ;
        RECT 97.950 803.100 100.050 805.200 ;
        RECT 100.950 803.100 103.050 805.200 ;
        RECT 109.950 803.100 112.050 805.200 ;
        RECT 112.950 803.100 115.050 805.200 ;
        RECT 115.950 803.100 118.050 805.200 ;
        RECT 131.700 805.050 132.600 815.400 ;
        RECT 151.800 812.400 153.600 818.400 ;
        RECT 154.800 815.400 156.600 819.000 ;
        RECT 157.800 815.400 159.600 818.400 ;
        RECT 151.800 805.050 153.000 812.400 ;
        RECT 158.400 811.500 159.600 815.400 ;
        RECT 153.900 810.600 159.600 811.500 ;
        RECT 167.400 810.600 169.200 818.400 ;
        RECT 171.900 812.400 173.700 819.000 ;
        RECT 174.900 814.200 176.700 818.400 ;
        RECT 174.900 812.400 177.600 814.200 ;
        RECT 193.500 812.400 195.300 819.000 ;
        RECT 198.000 812.400 199.800 818.400 ;
        RECT 202.500 812.400 204.300 819.000 ;
        RECT 214.800 812.400 216.600 818.400 ;
        RECT 217.800 815.400 219.600 819.000 ;
        RECT 220.800 815.400 222.600 818.400 ;
        RECT 173.100 810.600 174.900 811.500 ;
        RECT 153.900 809.700 155.850 810.600 ;
        RECT 167.400 809.700 174.900 810.600 ;
        RECT 41.550 801.000 45.450 801.450 ;
        RECT 40.950 800.550 45.450 801.000 ;
        RECT 40.950 796.950 43.050 800.550 ;
        RECT 32.700 789.900 39.300 790.800 ;
        RECT 32.700 789.600 34.200 789.900 ;
        RECT 29.400 783.000 31.200 789.600 ;
        RECT 32.400 783.600 34.200 789.600 ;
        RECT 38.400 789.600 39.300 789.900 ;
        RECT 53.700 790.800 54.600 803.100 ;
        RECT 59.100 801.300 60.900 803.100 ;
        RECT 53.700 789.900 60.300 790.800 ;
        RECT 53.700 789.600 54.600 789.900 ;
        RECT 35.400 783.000 37.200 789.000 ;
        RECT 38.400 783.600 40.200 789.600 ;
        RECT 52.800 783.600 54.600 789.600 ;
        RECT 58.800 789.600 60.300 789.900 ;
        RECT 74.400 789.600 75.600 803.100 ;
        RECT 92.700 790.800 93.600 803.100 ;
        RECT 98.100 801.300 99.900 803.100 ;
        RECT 100.950 801.450 103.050 802.050 ;
        RECT 109.950 801.450 112.050 802.050 ;
        RECT 100.950 800.550 112.050 801.450 ;
        RECT 100.950 799.950 103.050 800.550 ;
        RECT 109.950 799.950 112.050 800.550 ;
        RECT 92.700 789.900 99.300 790.800 ;
        RECT 92.700 789.600 93.600 789.900 ;
        RECT 55.800 783.000 57.600 789.000 ;
        RECT 58.800 783.600 60.600 789.600 ;
        RECT 61.800 783.000 63.600 789.600 ;
        RECT 71.400 783.000 73.200 789.600 ;
        RECT 74.400 783.600 76.200 789.600 ;
        RECT 77.400 783.000 79.200 789.600 ;
        RECT 91.800 783.600 93.600 789.600 ;
        RECT 97.800 789.600 99.300 789.900 ;
        RECT 113.400 789.600 114.600 803.100 ;
        RECT 127.950 802.950 130.050 805.050 ;
        RECT 130.950 802.950 133.050 805.050 ;
        RECT 133.950 802.950 136.050 805.050 ;
        RECT 151.800 802.950 154.050 805.050 ;
        RECT 128.100 801.150 129.900 802.950 ;
        RECT 131.700 795.600 132.600 802.950 ;
        RECT 134.100 801.150 135.900 802.950 ;
        RECT 151.800 795.600 153.000 802.950 ;
        RECT 154.950 798.300 155.850 809.700 ;
        RECT 167.100 805.200 168.900 807.000 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 166.950 803.100 169.050 805.200 ;
        RECT 158.100 801.150 159.900 802.950 ;
        RECT 153.900 797.400 155.850 798.300 ;
        RECT 153.900 796.500 159.600 797.400 ;
        RECT 94.800 783.000 96.600 789.000 ;
        RECT 97.800 783.600 99.600 789.600 ;
        RECT 100.800 783.000 102.600 789.600 ;
        RECT 110.400 783.000 112.200 789.600 ;
        RECT 113.400 783.600 115.200 789.600 ;
        RECT 116.400 783.000 118.200 789.600 ;
        RECT 128.400 783.000 130.200 795.600 ;
        RECT 131.700 794.400 135.300 795.600 ;
        RECT 133.500 783.600 135.300 794.400 ;
        RECT 151.800 783.600 153.600 795.600 ;
        RECT 158.400 789.600 159.600 796.500 ;
        RECT 170.400 789.600 171.300 809.700 ;
        RECT 176.700 805.200 177.600 812.400 ;
        RECT 191.100 805.200 192.900 807.000 ;
        RECT 198.000 805.200 199.050 812.400 ;
        RECT 203.100 805.200 204.900 807.000 ;
        RECT 172.950 803.100 175.050 805.200 ;
        RECT 175.950 803.100 178.050 805.200 ;
        RECT 190.950 803.100 193.050 805.200 ;
        RECT 193.950 803.100 196.050 805.200 ;
        RECT 196.950 803.100 199.050 805.200 ;
        RECT 199.950 803.100 202.050 805.200 ;
        RECT 202.950 803.100 205.050 805.200 ;
        RECT 214.800 805.050 216.000 812.400 ;
        RECT 221.400 811.500 222.600 815.400 ;
        RECT 230.700 812.400 232.500 819.000 ;
        RECT 235.200 812.400 237.000 818.400 ;
        RECT 239.700 812.400 241.500 819.000 ;
        RECT 216.900 810.600 222.600 811.500 ;
        RECT 216.900 809.700 218.850 810.600 ;
        RECT 173.100 801.300 174.900 803.100 ;
        RECT 176.700 795.600 177.600 803.100 ;
        RECT 194.100 801.300 195.900 803.100 ;
        RECT 198.000 797.400 198.900 803.100 ;
        RECT 200.100 801.300 201.900 803.100 ;
        RECT 214.800 802.950 217.050 805.050 ;
        RECT 193.800 796.500 198.900 797.400 ;
        RECT 154.800 783.000 156.600 789.600 ;
        RECT 157.800 783.600 159.600 789.600 ;
        RECT 167.400 783.000 169.200 789.600 ;
        RECT 170.400 783.600 172.200 789.600 ;
        RECT 173.400 783.000 175.200 789.600 ;
        RECT 176.400 783.600 178.200 795.600 ;
        RECT 190.800 784.500 192.600 795.600 ;
        RECT 193.800 785.400 195.600 796.500 ;
        RECT 214.800 795.600 216.000 802.950 ;
        RECT 217.950 798.300 218.850 809.700 ;
        RECT 230.100 805.200 231.900 807.000 ;
        RECT 235.950 805.200 237.000 812.400 ;
        RECT 259.200 810.000 261.000 818.400 ;
        RECT 257.700 808.800 261.000 810.000 ;
        RECT 265.800 809.400 267.600 819.000 ;
        RECT 275.700 812.400 277.500 819.000 ;
        RECT 280.800 811.200 282.600 818.400 ;
        RECT 293.700 812.400 295.500 819.000 ;
        RECT 298.200 812.400 300.000 818.400 ;
        RECT 302.700 812.400 304.500 819.000 ;
        RECT 319.800 815.400 321.600 818.400 ;
        RECT 322.800 815.400 324.600 819.000 ;
        RECT 278.400 810.300 282.600 811.200 ;
        RECT 242.100 805.200 243.900 807.000 ;
        RECT 257.700 805.200 258.600 808.800 ;
        RECT 260.100 805.200 261.900 807.000 ;
        RECT 266.100 805.200 267.900 807.000 ;
        RECT 275.100 805.200 276.900 807.000 ;
        RECT 278.400 805.200 279.600 810.300 ;
        RECT 281.100 805.200 282.900 807.000 ;
        RECT 293.100 805.200 294.900 807.000 ;
        RECT 298.950 805.200 300.000 812.400 ;
        RECT 305.100 805.200 306.900 807.000 ;
        RECT 220.950 802.950 223.050 805.050 ;
        RECT 229.950 803.100 232.050 805.200 ;
        RECT 232.950 803.100 235.050 805.200 ;
        RECT 235.950 803.100 238.050 805.200 ;
        RECT 238.950 803.100 241.050 805.200 ;
        RECT 241.950 803.100 244.050 805.200 ;
        RECT 256.950 803.100 259.050 805.200 ;
        RECT 259.950 803.100 262.050 805.200 ;
        RECT 262.950 803.100 265.050 805.200 ;
        RECT 265.950 803.100 268.050 805.200 ;
        RECT 274.950 803.100 277.050 805.200 ;
        RECT 277.950 803.100 280.050 805.200 ;
        RECT 280.950 803.100 283.050 805.200 ;
        RECT 292.950 803.100 295.050 805.200 ;
        RECT 295.950 803.100 298.050 805.200 ;
        RECT 298.950 803.100 301.050 805.200 ;
        RECT 301.950 803.100 304.050 805.200 ;
        RECT 304.950 803.100 307.050 805.200 ;
        RECT 320.400 805.050 321.600 815.400 ;
        RECT 332.700 812.400 334.500 819.000 ;
        RECT 337.800 811.200 339.600 818.400 ;
        RECT 335.400 810.300 339.600 811.200 ;
        RECT 352.800 812.400 354.600 818.400 ;
        RECT 355.800 815.400 357.600 819.000 ;
        RECT 358.800 815.400 360.600 818.400 ;
        RECT 332.100 805.200 333.900 807.000 ;
        RECT 335.400 805.200 336.600 810.300 ;
        RECT 338.100 805.200 339.900 807.000 ;
        RECT 221.100 801.150 222.900 802.950 ;
        RECT 233.100 801.300 234.900 803.100 ;
        RECT 216.900 797.400 218.850 798.300 ;
        RECT 236.100 797.400 237.000 803.100 ;
        RECT 239.100 801.300 240.900 803.100 ;
        RECT 216.900 796.500 222.600 797.400 ;
        RECT 236.100 796.500 241.200 797.400 ;
        RECT 196.800 794.400 204.600 795.300 ;
        RECT 196.800 784.500 198.600 794.400 ;
        RECT 190.800 783.600 198.600 784.500 ;
        RECT 199.800 783.000 201.600 793.500 ;
        RECT 202.800 783.600 204.600 794.400 ;
        RECT 214.800 783.600 216.600 795.600 ;
        RECT 221.400 789.600 222.600 796.500 ;
        RECT 217.800 783.000 219.600 789.600 ;
        RECT 220.800 783.600 222.600 789.600 ;
        RECT 230.400 794.400 238.200 795.300 ;
        RECT 230.400 783.600 232.200 794.400 ;
        RECT 233.400 783.000 235.200 793.500 ;
        RECT 236.400 784.500 238.200 794.400 ;
        RECT 239.400 785.400 241.200 796.500 ;
        RECT 242.400 784.500 244.200 795.600 ;
        RECT 257.700 790.800 258.600 803.100 ;
        RECT 263.100 801.300 264.900 803.100 ;
        RECT 257.700 789.900 264.300 790.800 ;
        RECT 257.700 789.600 258.600 789.900 ;
        RECT 236.400 783.600 244.200 784.500 ;
        RECT 256.800 783.600 258.600 789.600 ;
        RECT 262.800 789.600 264.300 789.900 ;
        RECT 278.400 789.600 279.600 803.100 ;
        RECT 296.100 801.300 297.900 803.100 ;
        RECT 299.100 797.400 300.000 803.100 ;
        RECT 302.100 801.300 303.900 803.100 ;
        RECT 319.950 802.950 322.050 805.050 ;
        RECT 322.950 802.950 325.050 805.050 ;
        RECT 331.950 803.100 334.050 805.200 ;
        RECT 334.950 803.100 337.050 805.200 ;
        RECT 337.950 803.100 340.050 805.200 ;
        RECT 352.800 805.050 354.000 812.400 ;
        RECT 359.400 811.500 360.600 815.400 ;
        RECT 372.300 814.200 374.100 818.400 ;
        RECT 354.900 810.600 360.600 811.500 ;
        RECT 371.400 812.400 374.100 814.200 ;
        RECT 375.300 812.400 377.100 819.000 ;
        RECT 354.900 809.700 356.850 810.600 ;
        RECT 299.100 796.500 304.200 797.400 ;
        RECT 293.400 794.400 301.200 795.300 ;
        RECT 259.800 783.000 261.600 789.000 ;
        RECT 262.800 783.600 264.600 789.600 ;
        RECT 265.800 783.000 267.600 789.600 ;
        RECT 275.400 783.000 277.200 789.600 ;
        RECT 278.400 783.600 280.200 789.600 ;
        RECT 281.400 783.000 283.200 789.600 ;
        RECT 293.400 783.600 295.200 794.400 ;
        RECT 296.400 783.000 298.200 793.500 ;
        RECT 299.400 784.500 301.200 794.400 ;
        RECT 302.400 785.400 304.200 796.500 ;
        RECT 305.400 784.500 307.200 795.600 ;
        RECT 320.400 789.600 321.600 802.950 ;
        RECT 323.100 801.150 324.900 802.950 ;
        RECT 335.400 789.600 336.600 803.100 ;
        RECT 352.800 802.950 355.050 805.050 ;
        RECT 352.800 795.600 354.000 802.950 ;
        RECT 355.950 798.300 356.850 809.700 ;
        RECT 371.400 805.200 372.300 812.400 ;
        RECT 374.100 810.600 375.900 811.500 ;
        RECT 379.800 810.600 381.600 818.400 ;
        RECT 389.400 813.300 391.200 818.400 ;
        RECT 392.400 814.200 394.200 819.000 ;
        RECT 395.400 813.300 397.200 818.400 ;
        RECT 389.400 811.950 397.200 813.300 ;
        RECT 398.400 812.400 400.200 818.400 ;
        RECT 410.700 812.400 412.500 819.000 ;
        RECT 415.200 812.400 417.000 818.400 ;
        RECT 419.700 812.400 421.500 819.000 ;
        RECT 436.800 812.400 438.600 818.400 ;
        RECT 439.800 815.400 441.600 819.000 ;
        RECT 442.800 815.400 444.600 818.400 ;
        RECT 452.400 815.400 454.200 819.000 ;
        RECT 455.400 815.400 457.200 818.400 ;
        RECT 374.100 809.700 381.600 810.600 ;
        RECT 398.400 810.300 399.600 812.400 ;
        RECT 358.950 802.950 361.050 805.050 ;
        RECT 370.950 803.100 373.050 805.200 ;
        RECT 373.950 803.100 376.050 805.200 ;
        RECT 359.100 801.150 360.900 802.950 ;
        RECT 354.900 797.400 356.850 798.300 ;
        RECT 354.900 796.500 360.600 797.400 ;
        RECT 299.400 783.600 307.200 784.500 ;
        RECT 319.800 783.600 321.600 789.600 ;
        RECT 322.800 783.000 324.600 789.600 ;
        RECT 332.400 783.000 334.200 789.600 ;
        RECT 335.400 783.600 337.200 789.600 ;
        RECT 338.400 783.000 340.200 789.600 ;
        RECT 352.800 783.600 354.600 795.600 ;
        RECT 359.400 789.600 360.600 796.500 ;
        RECT 371.400 795.600 372.300 803.100 ;
        RECT 374.100 801.300 375.900 803.100 ;
        RECT 355.800 783.000 357.600 789.600 ;
        RECT 358.800 783.600 360.600 789.600 ;
        RECT 370.800 783.600 372.600 795.600 ;
        RECT 377.700 789.600 378.600 809.700 ;
        RECT 395.850 809.250 399.600 810.300 ;
        RECT 380.100 805.200 381.900 807.000 ;
        RECT 379.950 803.100 382.050 805.200 ;
        RECT 392.100 805.050 393.900 806.850 ;
        RECT 395.850 805.050 397.050 809.250 ;
        RECT 398.100 805.050 399.900 806.850 ;
        RECT 410.100 805.200 411.900 807.000 ;
        RECT 415.950 805.200 417.000 812.400 ;
        RECT 418.950 810.450 421.050 811.050 ;
        RECT 430.950 810.450 433.050 811.050 ;
        RECT 418.950 809.550 433.050 810.450 ;
        RECT 418.950 808.950 421.050 809.550 ;
        RECT 430.950 808.950 433.050 809.550 ;
        RECT 422.100 805.200 423.900 807.000 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 391.950 802.950 394.050 805.050 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 409.950 803.100 412.050 805.200 ;
        RECT 412.950 803.100 415.050 805.200 ;
        RECT 415.950 803.100 418.050 805.200 ;
        RECT 418.950 803.100 421.050 805.200 ;
        RECT 421.950 803.100 424.050 805.200 ;
        RECT 436.800 805.050 438.000 812.400 ;
        RECT 443.400 811.500 444.600 815.400 ;
        RECT 438.900 810.600 444.600 811.500 ;
        RECT 438.900 809.700 440.850 810.600 ;
        RECT 389.100 801.150 390.900 802.950 ;
        RECT 373.800 783.000 375.600 789.600 ;
        RECT 376.800 783.600 378.600 789.600 ;
        RECT 379.800 783.000 381.600 789.600 ;
        RECT 389.700 783.000 391.500 795.600 ;
        RECT 394.950 789.600 396.150 802.950 ;
        RECT 413.100 801.300 414.900 803.100 ;
        RECT 416.100 797.400 417.000 803.100 ;
        RECT 419.100 801.300 420.900 803.100 ;
        RECT 436.800 802.950 439.050 805.050 ;
        RECT 416.100 796.500 421.200 797.400 ;
        RECT 410.400 794.400 418.200 795.300 ;
        RECT 394.800 783.600 396.600 789.600 ;
        RECT 397.800 783.000 399.600 789.600 ;
        RECT 410.400 783.600 412.200 794.400 ;
        RECT 413.400 783.000 415.200 793.500 ;
        RECT 416.400 784.500 418.200 794.400 ;
        RECT 419.400 785.400 421.200 796.500 ;
        RECT 436.800 795.600 438.000 802.950 ;
        RECT 439.950 798.300 440.850 809.700 ;
        RECT 455.400 805.050 456.600 815.400 ;
        RECT 468.000 812.400 469.800 819.000 ;
        RECT 472.500 813.600 474.300 818.400 ;
        RECT 475.500 815.400 477.300 819.000 ;
        RECT 472.500 812.400 477.600 813.600 ;
        RECT 467.100 805.200 468.900 807.000 ;
        RECT 473.100 805.200 474.900 807.000 ;
        RECT 476.700 805.200 477.600 812.400 ;
        RECT 493.200 810.000 495.000 818.400 ;
        RECT 491.700 808.800 495.000 810.000 ;
        RECT 499.800 809.400 501.600 819.000 ;
        RECT 509.400 809.400 511.200 819.000 ;
        RECT 516.000 810.000 517.800 818.400 ;
        RECT 531.000 812.400 532.800 819.000 ;
        RECT 535.500 813.600 537.300 818.400 ;
        RECT 538.500 815.400 540.300 819.000 ;
        RECT 535.500 812.400 540.600 813.600 ;
        RECT 553.800 812.400 555.600 818.400 ;
        RECT 516.000 808.800 519.300 810.000 ;
        RECT 491.700 805.200 492.600 808.800 ;
        RECT 494.100 805.200 495.900 807.000 ;
        RECT 500.100 805.200 501.900 807.000 ;
        RECT 509.100 805.200 510.900 807.000 ;
        RECT 515.100 805.200 516.900 807.000 ;
        RECT 518.400 805.200 519.300 808.800 ;
        RECT 530.100 805.200 531.900 807.000 ;
        RECT 536.100 805.200 537.900 807.000 ;
        RECT 539.700 805.200 540.600 812.400 ;
        RECT 554.400 810.300 555.600 812.400 ;
        RECT 556.800 813.300 558.600 818.400 ;
        RECT 559.800 814.200 561.600 819.000 ;
        RECT 562.800 813.300 564.600 818.400 ;
        RECT 556.800 811.950 564.600 813.300 ;
        RECT 574.800 812.400 576.600 818.400 ;
        RECT 565.950 810.450 568.050 811.050 ;
        RECT 571.950 810.450 574.050 811.050 ;
        RECT 554.400 809.250 558.150 810.300 ;
        RECT 541.950 807.450 546.000 808.050 ;
        RECT 541.950 805.950 546.450 807.450 ;
        RECT 442.950 802.950 445.050 805.050 ;
        RECT 451.950 802.950 454.050 805.050 ;
        RECT 454.950 802.950 457.050 805.050 ;
        RECT 466.950 803.100 469.050 805.200 ;
        RECT 469.950 803.100 472.050 805.200 ;
        RECT 472.950 803.100 475.050 805.200 ;
        RECT 475.950 803.100 478.050 805.200 ;
        RECT 490.950 803.100 493.050 805.200 ;
        RECT 493.950 803.100 496.050 805.200 ;
        RECT 496.950 803.100 499.050 805.200 ;
        RECT 499.950 803.100 502.050 805.200 ;
        RECT 508.950 803.100 511.050 805.200 ;
        RECT 511.950 803.100 514.050 805.200 ;
        RECT 514.950 803.100 517.050 805.200 ;
        RECT 517.950 803.100 520.050 805.200 ;
        RECT 529.950 803.100 532.050 805.200 ;
        RECT 532.950 803.100 535.050 805.200 ;
        RECT 535.950 803.100 538.050 805.200 ;
        RECT 538.950 803.100 541.050 805.200 ;
        RECT 443.100 801.150 444.900 802.950 ;
        RECT 452.100 801.150 453.900 802.950 ;
        RECT 438.900 797.400 440.850 798.300 ;
        RECT 438.900 796.500 444.600 797.400 ;
        RECT 422.400 784.500 424.200 795.600 ;
        RECT 416.400 783.600 424.200 784.500 ;
        RECT 436.800 783.600 438.600 795.600 ;
        RECT 443.400 789.600 444.600 796.500 ;
        RECT 455.400 789.600 456.600 802.950 ;
        RECT 470.100 801.300 471.900 803.100 ;
        RECT 457.950 798.450 460.050 799.050 ;
        RECT 472.950 798.450 475.050 799.050 ;
        RECT 457.950 797.550 475.050 798.450 ;
        RECT 457.950 796.950 460.050 797.550 ;
        RECT 472.950 796.950 475.050 797.550 ;
        RECT 476.700 795.600 477.600 803.100 ;
        RECT 467.400 794.700 475.200 795.600 ;
        RECT 439.800 783.000 441.600 789.600 ;
        RECT 442.800 783.600 444.600 789.600 ;
        RECT 452.400 783.000 454.200 789.600 ;
        RECT 455.400 783.600 457.200 789.600 ;
        RECT 467.400 783.600 469.200 794.700 ;
        RECT 470.400 783.000 472.200 793.800 ;
        RECT 473.400 783.600 475.200 794.700 ;
        RECT 476.400 783.600 478.200 795.600 ;
        RECT 491.700 790.800 492.600 803.100 ;
        RECT 497.100 801.300 498.900 803.100 ;
        RECT 512.100 801.300 513.900 803.100 ;
        RECT 493.950 798.450 496.050 799.050 ;
        RECT 514.950 798.450 517.050 799.050 ;
        RECT 493.950 797.550 517.050 798.450 ;
        RECT 493.950 796.950 496.050 797.550 ;
        RECT 514.950 796.950 517.050 797.550 ;
        RECT 493.950 795.450 496.050 795.900 ;
        RECT 499.950 795.450 502.050 796.050 ;
        RECT 493.950 794.550 502.050 795.450 ;
        RECT 493.950 793.800 496.050 794.550 ;
        RECT 499.950 793.950 502.050 794.550 ;
        RECT 518.400 790.800 519.300 803.100 ;
        RECT 533.100 801.300 534.900 803.100 ;
        RECT 539.700 795.600 540.600 803.100 ;
        RECT 545.550 802.050 546.450 805.950 ;
        RECT 554.100 805.050 555.900 806.850 ;
        RECT 556.950 805.050 558.150 809.250 ;
        RECT 565.950 809.550 574.050 810.450 ;
        RECT 565.950 808.950 568.050 809.550 ;
        RECT 571.950 808.950 574.050 809.550 ;
        RECT 575.400 810.300 576.600 812.400 ;
        RECT 577.800 813.300 579.600 818.400 ;
        RECT 580.800 814.200 582.600 819.000 ;
        RECT 583.800 813.300 585.600 818.400 ;
        RECT 577.800 811.950 585.600 813.300 ;
        RECT 596.400 811.200 598.200 818.400 ;
        RECT 601.500 812.400 603.300 819.000 ;
        RECT 613.800 812.400 615.600 818.400 ;
        RECT 596.400 810.300 600.600 811.200 ;
        RECT 575.400 809.250 579.150 810.300 ;
        RECT 560.100 805.050 561.900 806.850 ;
        RECT 575.100 805.050 576.900 806.850 ;
        RECT 577.950 805.050 579.150 809.250 ;
        RECT 581.100 805.050 582.900 806.850 ;
        RECT 596.100 805.200 597.900 807.000 ;
        RECT 599.400 805.200 600.600 810.300 ;
        RECT 614.400 810.300 615.600 812.400 ;
        RECT 616.800 813.300 618.600 818.400 ;
        RECT 619.800 814.200 621.600 819.000 ;
        RECT 622.800 813.300 624.600 818.400 ;
        RECT 635.700 815.400 637.500 819.000 ;
        RECT 638.700 813.600 640.500 818.400 ;
        RECT 616.800 811.950 624.600 813.300 ;
        RECT 635.400 812.400 640.500 813.600 ;
        RECT 643.200 812.400 645.000 819.000 ;
        RECT 614.400 809.250 618.150 810.300 ;
        RECT 602.100 805.200 603.900 807.000 ;
        RECT 553.950 802.950 556.050 805.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 562.950 802.950 565.050 805.050 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 583.950 802.950 586.050 805.050 ;
        RECT 595.950 803.100 598.050 805.200 ;
        RECT 598.950 803.100 601.050 805.200 ;
        RECT 601.950 803.100 604.050 805.200 ;
        RECT 614.100 805.050 615.900 806.850 ;
        RECT 616.950 805.050 618.150 809.250 ;
        RECT 620.100 805.050 621.900 806.850 ;
        RECT 635.400 805.200 636.300 812.400 ;
        RECT 658.200 810.000 660.000 818.400 ;
        RECT 656.700 808.800 660.000 810.000 ;
        RECT 664.800 809.400 666.600 819.000 ;
        RECT 674.400 815.400 676.200 819.000 ;
        RECT 677.400 815.400 679.200 818.400 ;
        RECT 689.400 815.400 691.200 819.000 ;
        RECT 692.400 815.400 694.200 818.400 ;
        RECT 638.100 805.200 639.900 807.000 ;
        RECT 644.100 805.200 645.900 807.000 ;
        RECT 656.700 805.200 657.600 808.800 ;
        RECT 659.100 805.200 660.900 807.000 ;
        RECT 665.100 805.200 666.900 807.000 ;
        RECT 541.950 800.550 546.450 802.050 ;
        RECT 541.950 799.950 546.000 800.550 ;
        RECT 491.700 789.900 498.300 790.800 ;
        RECT 491.700 789.600 492.600 789.900 ;
        RECT 490.800 783.600 492.600 789.600 ;
        RECT 496.800 789.600 498.300 789.900 ;
        RECT 512.700 789.900 519.300 790.800 ;
        RECT 512.700 789.600 514.200 789.900 ;
        RECT 493.800 783.000 495.600 789.000 ;
        RECT 496.800 783.600 498.600 789.600 ;
        RECT 499.800 783.000 501.600 789.600 ;
        RECT 509.400 783.000 511.200 789.600 ;
        RECT 512.400 783.600 514.200 789.600 ;
        RECT 518.400 789.600 519.300 789.900 ;
        RECT 530.400 794.700 538.200 795.600 ;
        RECT 515.400 783.000 517.200 789.000 ;
        RECT 518.400 783.600 520.200 789.600 ;
        RECT 530.400 783.600 532.200 794.700 ;
        RECT 533.400 783.000 535.200 793.800 ;
        RECT 536.400 783.600 538.200 794.700 ;
        RECT 539.400 783.600 541.200 795.600 ;
        RECT 557.850 789.600 559.050 802.950 ;
        RECT 563.100 801.150 564.900 802.950 ;
        RECT 565.950 798.450 568.050 799.050 ;
        RECT 574.950 798.450 577.050 799.050 ;
        RECT 565.950 797.550 577.050 798.450 ;
        RECT 565.950 796.950 568.050 797.550 ;
        RECT 574.950 796.950 577.050 797.550 ;
        RECT 554.400 783.000 556.200 789.600 ;
        RECT 557.400 783.600 559.200 789.600 ;
        RECT 562.500 783.000 564.300 795.600 ;
        RECT 578.850 789.600 580.050 802.950 ;
        RECT 584.100 801.150 585.900 802.950 ;
        RECT 575.400 783.000 577.200 789.600 ;
        RECT 578.400 783.600 580.200 789.600 ;
        RECT 583.500 783.000 585.300 795.600 ;
        RECT 599.400 789.600 600.600 803.100 ;
        RECT 613.950 802.950 616.050 805.050 ;
        RECT 616.950 802.950 619.050 805.050 ;
        RECT 619.950 802.950 622.050 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 634.950 803.100 637.050 805.200 ;
        RECT 637.950 803.100 640.050 805.200 ;
        RECT 640.950 803.100 643.050 805.200 ;
        RECT 643.950 803.100 646.050 805.200 ;
        RECT 655.950 803.100 658.050 805.200 ;
        RECT 658.950 803.100 661.050 805.200 ;
        RECT 661.950 803.100 664.050 805.200 ;
        RECT 664.950 803.100 667.050 805.200 ;
        RECT 677.400 805.050 678.600 815.400 ;
        RECT 692.400 805.050 693.600 815.400 ;
        RECT 705.000 812.400 706.800 819.000 ;
        RECT 709.500 813.600 711.300 818.400 ;
        RECT 712.500 815.400 714.300 819.000 ;
        RECT 709.500 812.400 714.600 813.600 ;
        RECT 704.100 805.200 705.900 807.000 ;
        RECT 710.100 805.200 711.900 807.000 ;
        RECT 713.700 805.200 714.600 812.400 ;
        RECT 725.400 813.300 727.200 818.400 ;
        RECT 728.400 814.200 730.200 819.000 ;
        RECT 731.400 813.300 733.200 818.400 ;
        RECT 725.400 811.950 733.200 813.300 ;
        RECT 734.400 812.400 736.200 818.400 ;
        RECT 747.000 812.400 748.800 819.000 ;
        RECT 751.500 813.600 753.300 818.400 ;
        RECT 754.500 815.400 756.300 819.000 ;
        RECT 751.500 812.400 756.600 813.600 ;
        RECT 767.700 812.400 769.500 819.000 ;
        RECT 734.400 810.300 735.600 812.400 ;
        RECT 731.850 809.250 735.600 810.300 ;
        RECT 617.850 789.600 619.050 802.950 ;
        RECT 623.100 801.150 624.900 802.950 ;
        RECT 635.400 795.600 636.300 803.100 ;
        RECT 641.100 801.300 642.900 803.100 ;
        RECT 595.800 783.000 597.600 789.600 ;
        RECT 598.800 783.600 600.600 789.600 ;
        RECT 601.800 783.000 603.600 789.600 ;
        RECT 614.400 783.000 616.200 789.600 ;
        RECT 617.400 783.600 619.200 789.600 ;
        RECT 622.500 783.000 624.300 795.600 ;
        RECT 634.800 783.600 636.600 795.600 ;
        RECT 637.800 794.700 645.600 795.600 ;
        RECT 637.800 783.600 639.600 794.700 ;
        RECT 640.800 783.000 642.600 793.800 ;
        RECT 643.800 783.600 645.600 794.700 ;
        RECT 656.700 790.800 657.600 803.100 ;
        RECT 662.100 801.300 663.900 803.100 ;
        RECT 673.950 802.950 676.050 805.050 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 688.950 802.950 691.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 703.950 803.100 706.050 805.200 ;
        RECT 706.950 803.100 709.050 805.200 ;
        RECT 709.950 803.100 712.050 805.200 ;
        RECT 712.950 803.100 715.050 805.200 ;
        RECT 728.100 805.050 729.900 806.850 ;
        RECT 731.850 805.050 733.050 809.250 ;
        RECT 734.100 805.050 735.900 806.850 ;
        RECT 746.100 805.200 747.900 807.000 ;
        RECT 752.100 805.200 753.900 807.000 ;
        RECT 755.700 805.200 756.600 812.400 ;
        RECT 772.800 811.200 774.600 818.400 ;
        RECT 786.000 812.400 787.800 819.000 ;
        RECT 790.500 813.600 792.300 818.400 ;
        RECT 793.500 815.400 795.300 819.000 ;
        RECT 790.500 812.400 795.600 813.600 ;
        RECT 808.800 812.400 810.600 818.400 ;
        RECT 770.400 810.300 774.600 811.200 ;
        RECT 767.100 805.200 768.900 807.000 ;
        RECT 770.400 805.200 771.600 810.300 ;
        RECT 773.100 805.200 774.900 807.000 ;
        RECT 785.100 805.200 786.900 807.000 ;
        RECT 791.100 805.200 792.900 807.000 ;
        RECT 794.700 805.200 795.600 812.400 ;
        RECT 809.400 810.300 810.600 812.400 ;
        RECT 811.800 813.300 813.600 818.400 ;
        RECT 814.800 814.200 816.600 819.000 ;
        RECT 817.800 813.300 819.600 818.400 ;
        RECT 811.800 811.950 819.600 813.300 ;
        RECT 827.400 813.300 829.200 818.400 ;
        RECT 830.400 814.200 832.200 819.000 ;
        RECT 833.400 813.300 835.200 818.400 ;
        RECT 827.400 811.950 835.200 813.300 ;
        RECT 836.400 812.400 838.200 818.400 ;
        RECT 836.400 810.300 837.600 812.400 ;
        RECT 809.400 809.250 813.150 810.300 ;
        RECT 674.100 801.150 675.900 802.950 ;
        RECT 664.950 798.450 667.050 799.050 ;
        RECT 673.950 798.450 676.050 799.050 ;
        RECT 664.950 797.550 676.050 798.450 ;
        RECT 664.950 796.950 667.050 797.550 ;
        RECT 673.950 796.950 676.050 797.550 ;
        RECT 656.700 789.900 663.300 790.800 ;
        RECT 656.700 789.600 657.600 789.900 ;
        RECT 655.800 783.600 657.600 789.600 ;
        RECT 661.800 789.600 663.300 789.900 ;
        RECT 677.400 789.600 678.600 802.950 ;
        RECT 689.100 801.150 690.900 802.950 ;
        RECT 692.400 789.600 693.600 802.950 ;
        RECT 707.100 801.300 708.900 803.100 ;
        RECT 713.700 795.600 714.600 803.100 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 727.950 802.950 730.050 805.050 ;
        RECT 730.950 802.950 733.050 805.050 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 745.950 803.100 748.050 805.200 ;
        RECT 748.950 803.100 751.050 805.200 ;
        RECT 751.950 803.100 754.050 805.200 ;
        RECT 754.950 803.100 757.050 805.200 ;
        RECT 766.950 803.100 769.050 805.200 ;
        RECT 769.950 803.100 772.050 805.200 ;
        RECT 772.950 803.100 775.050 805.200 ;
        RECT 784.950 803.100 787.050 805.200 ;
        RECT 787.950 803.100 790.050 805.200 ;
        RECT 790.950 803.100 793.050 805.200 ;
        RECT 793.950 803.100 796.050 805.200 ;
        RECT 809.100 805.050 810.900 806.850 ;
        RECT 811.950 805.050 813.150 809.250 ;
        RECT 833.850 809.250 837.600 810.300 ;
        RECT 815.100 805.050 816.900 806.850 ;
        RECT 830.100 805.050 831.900 806.850 ;
        RECT 833.850 805.050 835.050 809.250 ;
        RECT 836.100 805.050 837.900 806.850 ;
        RECT 725.100 801.150 726.900 802.950 ;
        RECT 704.400 794.700 712.200 795.600 ;
        RECT 658.800 783.000 660.600 789.000 ;
        RECT 661.800 783.600 663.600 789.600 ;
        RECT 664.800 783.000 666.600 789.600 ;
        RECT 674.400 783.000 676.200 789.600 ;
        RECT 677.400 783.600 679.200 789.600 ;
        RECT 689.400 783.000 691.200 789.600 ;
        RECT 692.400 783.600 694.200 789.600 ;
        RECT 704.400 783.600 706.200 794.700 ;
        RECT 707.400 783.000 709.200 793.800 ;
        RECT 710.400 783.600 712.200 794.700 ;
        RECT 713.400 783.600 715.200 795.600 ;
        RECT 725.700 783.000 727.500 795.600 ;
        RECT 730.950 789.600 732.150 802.950 ;
        RECT 749.100 801.300 750.900 803.100 ;
        RECT 742.950 798.450 745.050 799.050 ;
        RECT 751.950 798.450 754.050 799.050 ;
        RECT 742.950 797.550 754.050 798.450 ;
        RECT 742.950 796.950 745.050 797.550 ;
        RECT 751.950 796.950 754.050 797.550 ;
        RECT 755.700 795.600 756.600 803.100 ;
        RECT 746.400 794.700 754.200 795.600 ;
        RECT 730.800 783.600 732.600 789.600 ;
        RECT 733.800 783.000 735.600 789.600 ;
        RECT 746.400 783.600 748.200 794.700 ;
        RECT 749.400 783.000 751.200 793.800 ;
        RECT 752.400 783.600 754.200 794.700 ;
        RECT 755.400 783.600 757.200 795.600 ;
        RECT 770.400 789.600 771.600 803.100 ;
        RECT 788.100 801.300 789.900 803.100 ;
        RECT 794.700 795.600 795.600 803.100 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 811.950 802.950 814.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 817.950 802.950 820.050 805.050 ;
        RECT 826.950 802.950 829.050 805.050 ;
        RECT 829.950 802.950 832.050 805.050 ;
        RECT 832.950 802.950 835.050 805.050 ;
        RECT 835.950 802.950 838.050 805.050 ;
        RECT 785.400 794.700 793.200 795.600 ;
        RECT 767.400 783.000 769.200 789.600 ;
        RECT 770.400 783.600 772.200 789.600 ;
        RECT 773.400 783.000 775.200 789.600 ;
        RECT 785.400 783.600 787.200 794.700 ;
        RECT 788.400 783.000 790.200 793.800 ;
        RECT 791.400 783.600 793.200 794.700 ;
        RECT 794.400 783.600 796.200 795.600 ;
        RECT 812.850 789.600 814.050 802.950 ;
        RECT 818.100 801.150 819.900 802.950 ;
        RECT 827.100 801.150 828.900 802.950 ;
        RECT 809.400 783.000 811.200 789.600 ;
        RECT 812.400 783.600 814.200 789.600 ;
        RECT 817.500 783.000 819.300 795.600 ;
        RECT 827.700 783.000 829.500 795.600 ;
        RECT 832.950 789.600 834.150 802.950 ;
        RECT 832.800 783.600 834.600 789.600 ;
        RECT 835.800 783.000 837.600 789.600 ;
        RECT 11.400 773.400 13.200 780.000 ;
        RECT 14.400 773.400 16.200 779.400 ;
        RECT 14.850 760.050 16.050 773.400 ;
        RECT 19.500 767.400 21.300 780.000 ;
        RECT 29.700 767.400 31.500 780.000 ;
        RECT 34.800 773.400 36.600 779.400 ;
        RECT 37.800 773.400 39.600 780.000 ;
        RECT 52.800 773.400 54.600 779.400 ;
        RECT 55.800 773.400 57.600 780.000 ;
        RECT 20.100 760.050 21.900 761.850 ;
        RECT 29.100 760.050 30.900 761.850 ;
        RECT 34.950 760.050 36.150 773.400 ;
        RECT 53.400 760.050 54.600 773.400 ;
        RECT 67.800 767.400 69.600 779.400 ;
        RECT 70.800 768.300 72.600 779.400 ;
        RECT 73.800 769.200 75.600 780.000 ;
        RECT 76.800 768.300 78.600 779.400 ;
        RECT 88.800 773.400 90.600 779.400 ;
        RECT 91.800 774.000 93.600 780.000 ;
        RECT 70.800 767.400 78.600 768.300 ;
        RECT 89.700 773.100 90.600 773.400 ;
        RECT 94.800 773.400 96.600 779.400 ;
        RECT 97.800 773.400 99.600 780.000 ;
        RECT 107.400 773.400 109.200 780.000 ;
        RECT 110.400 773.400 112.200 779.400 ;
        RECT 94.800 773.100 96.300 773.400 ;
        RECT 89.700 772.200 96.300 773.100 ;
        RECT 56.100 760.050 57.900 761.850 ;
        RECT 10.950 757.950 13.050 760.050 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 28.950 757.950 31.050 760.050 ;
        RECT 31.950 757.950 34.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 52.950 757.950 55.050 760.050 ;
        RECT 55.950 757.950 58.050 760.050 ;
        RECT 68.400 759.900 69.300 767.400 ;
        RECT 79.950 762.450 84.000 763.050 ;
        RECT 74.100 759.900 75.900 761.700 ;
        RECT 79.950 760.950 84.450 762.450 ;
        RECT 11.100 756.150 12.900 757.950 ;
        RECT 13.950 753.750 15.150 757.950 ;
        RECT 17.100 756.150 18.900 757.950 ;
        RECT 32.100 756.150 33.900 757.950 ;
        RECT 11.400 752.700 15.150 753.750 ;
        RECT 35.850 753.750 37.050 757.950 ;
        RECT 38.100 756.150 39.900 757.950 ;
        RECT 35.850 752.700 39.600 753.750 ;
        RECT 11.400 750.600 12.600 752.700 ;
        RECT 10.800 744.600 12.600 750.600 ;
        RECT 13.800 749.700 21.600 751.050 ;
        RECT 13.800 744.600 15.600 749.700 ;
        RECT 16.800 744.000 18.600 748.800 ;
        RECT 19.800 744.600 21.600 749.700 ;
        RECT 29.400 749.700 37.200 751.050 ;
        RECT 29.400 744.600 31.200 749.700 ;
        RECT 32.400 744.000 34.200 748.800 ;
        RECT 35.400 744.600 37.200 749.700 ;
        RECT 38.400 750.600 39.600 752.700 ;
        RECT 38.400 744.600 40.200 750.600 ;
        RECT 53.400 747.600 54.600 757.950 ;
        RECT 67.950 757.800 70.050 759.900 ;
        RECT 70.950 757.800 73.050 759.900 ;
        RECT 73.950 757.800 76.050 759.900 ;
        RECT 76.950 757.800 79.050 759.900 ;
        RECT 68.400 750.600 69.300 757.800 ;
        RECT 71.100 756.000 72.900 757.800 ;
        RECT 77.100 756.000 78.900 757.800 ;
        RECT 83.550 757.050 84.450 760.950 ;
        RECT 89.700 759.900 90.600 772.200 ;
        RECT 97.950 768.450 100.050 769.050 ;
        RECT 106.950 768.450 109.050 769.050 ;
        RECT 97.950 767.550 109.050 768.450 ;
        RECT 97.950 766.950 100.050 767.550 ;
        RECT 106.950 766.950 109.050 767.550 ;
        RECT 91.950 765.450 94.050 766.050 ;
        RECT 100.950 765.450 103.050 766.050 ;
        RECT 91.950 764.550 103.050 765.450 ;
        RECT 91.950 763.950 94.050 764.550 ;
        RECT 100.950 763.950 103.050 764.550 ;
        RECT 95.100 759.900 96.900 761.700 ;
        RECT 107.100 760.050 108.900 761.850 ;
        RECT 110.400 760.050 111.600 773.400 ;
        RECT 122.400 768.300 124.200 779.400 ;
        RECT 125.400 769.200 127.200 780.000 ;
        RECT 128.400 768.300 130.200 779.400 ;
        RECT 122.400 767.400 130.200 768.300 ;
        RECT 131.400 767.400 133.200 779.400 ;
        RECT 143.400 773.400 145.200 780.000 ;
        RECT 146.400 773.400 148.200 779.400 ;
        RECT 149.400 773.400 151.200 780.000 ;
        RECT 88.950 757.800 91.050 759.900 ;
        RECT 91.950 757.800 94.050 759.900 ;
        RECT 94.950 757.800 97.050 759.900 ;
        RECT 97.950 757.800 100.050 759.900 ;
        RECT 106.950 757.950 109.050 760.050 ;
        RECT 109.950 757.950 112.050 760.050 ;
        RECT 125.100 759.900 126.900 761.700 ;
        RECT 131.700 759.900 132.600 767.400 ;
        RECT 138.000 762.450 142.050 763.050 ;
        RECT 137.550 760.950 142.050 762.450 ;
        RECT 79.950 755.550 84.450 757.050 ;
        RECT 79.950 754.950 84.000 755.550 ;
        RECT 89.700 754.200 90.600 757.800 ;
        RECT 92.100 756.000 93.900 757.800 ;
        RECT 98.100 756.000 99.900 757.800 ;
        RECT 89.700 753.000 93.000 754.200 ;
        RECT 68.400 749.400 73.500 750.600 ;
        RECT 52.800 744.600 54.600 747.600 ;
        RECT 55.800 744.000 57.600 747.600 ;
        RECT 68.700 744.000 70.500 747.600 ;
        RECT 71.700 744.600 73.500 749.400 ;
        RECT 76.200 744.000 78.000 750.600 ;
        RECT 91.200 744.600 93.000 753.000 ;
        RECT 97.800 744.000 99.600 753.600 ;
        RECT 110.400 747.600 111.600 757.950 ;
        RECT 121.950 757.800 124.050 759.900 ;
        RECT 124.950 757.800 127.050 759.900 ;
        RECT 127.950 757.800 130.050 759.900 ;
        RECT 130.950 757.800 133.050 759.900 ;
        RECT 122.100 756.000 123.900 757.800 ;
        RECT 128.100 756.000 129.900 757.800 ;
        RECT 131.700 750.600 132.600 757.800 ;
        RECT 137.550 757.050 138.450 760.950 ;
        RECT 142.950 757.800 145.050 759.900 ;
        RECT 133.950 755.550 138.450 757.050 ;
        RECT 143.100 756.000 144.900 757.800 ;
        RECT 133.950 754.950 138.000 755.550 ;
        RECT 146.400 753.300 147.300 773.400 ;
        RECT 152.400 767.400 154.200 779.400 ;
        RECT 164.400 773.400 166.200 780.000 ;
        RECT 167.400 773.400 169.200 779.400 ;
        RECT 170.400 773.400 172.200 780.000 ;
        RECT 149.100 759.900 150.900 761.700 ;
        RECT 152.700 759.900 153.600 767.400 ;
        RECT 167.400 759.900 168.600 773.400 ;
        RECT 182.700 767.400 184.500 780.000 ;
        RECT 187.800 773.400 189.600 779.400 ;
        RECT 190.800 773.400 192.600 780.000 ;
        RECT 206.400 773.400 208.200 780.000 ;
        RECT 209.400 773.400 211.200 779.400 ;
        RECT 182.100 760.050 183.900 761.850 ;
        RECT 187.950 760.050 189.150 773.400 ;
        RECT 209.850 760.050 211.050 773.400 ;
        RECT 214.500 767.400 216.300 780.000 ;
        RECT 227.400 773.400 229.200 780.000 ;
        RECT 230.400 773.400 232.200 779.400 ;
        RECT 215.100 760.050 216.900 761.850 ;
        RECT 230.850 760.050 232.050 773.400 ;
        RECT 235.500 767.400 237.300 780.000 ;
        RECT 247.800 773.400 249.600 779.400 ;
        RECT 250.800 774.000 252.600 780.000 ;
        RECT 248.700 773.100 249.600 773.400 ;
        RECT 253.800 773.400 255.600 779.400 ;
        RECT 256.800 773.400 258.600 780.000 ;
        RECT 266.400 773.400 268.200 780.000 ;
        RECT 269.400 773.400 271.200 779.400 ;
        RECT 272.400 774.000 274.200 780.000 ;
        RECT 253.800 773.100 255.300 773.400 ;
        RECT 248.700 772.200 255.300 773.100 ;
        RECT 269.700 773.100 271.200 773.400 ;
        RECT 275.400 773.400 277.200 779.400 ;
        RECT 275.400 773.100 276.300 773.400 ;
        RECT 269.700 772.200 276.300 773.100 ;
        RECT 236.100 760.050 237.900 761.850 ;
        RECT 148.950 757.800 151.050 759.900 ;
        RECT 151.950 757.800 154.050 759.900 ;
        RECT 163.950 757.800 166.050 759.900 ;
        RECT 166.950 757.800 169.050 759.900 ;
        RECT 169.950 757.800 172.050 759.900 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 205.950 757.950 208.050 760.050 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 226.950 757.950 229.050 760.050 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 248.700 759.900 249.600 772.200 ;
        RECT 254.100 759.900 255.900 761.700 ;
        RECT 269.100 759.900 270.900 761.700 ;
        RECT 275.400 759.900 276.300 772.200 ;
        RECT 287.400 768.300 289.200 779.400 ;
        RECT 290.400 769.200 292.200 780.000 ;
        RECT 293.400 768.300 295.200 779.400 ;
        RECT 287.400 767.400 295.200 768.300 ;
        RECT 296.400 767.400 298.200 779.400 ;
        RECT 310.800 773.400 312.600 779.400 ;
        RECT 313.800 774.000 315.600 780.000 ;
        RECT 311.700 773.100 312.600 773.400 ;
        RECT 316.800 773.400 318.600 779.400 ;
        RECT 319.800 773.400 321.600 780.000 ;
        RECT 316.800 773.100 318.300 773.400 ;
        RECT 311.700 772.200 318.300 773.100 ;
        RECT 292.950 765.450 295.050 766.050 ;
        RECT 287.550 764.550 295.050 765.450 ;
        RECT 287.550 762.450 288.450 764.550 ;
        RECT 292.950 763.950 295.050 764.550 ;
        RECT 281.550 761.550 288.450 762.450 ;
        RECT 107.400 744.000 109.200 747.600 ;
        RECT 110.400 744.600 112.200 747.600 ;
        RECT 123.000 744.000 124.800 750.600 ;
        RECT 127.500 749.400 132.600 750.600 ;
        RECT 143.400 752.400 150.900 753.300 ;
        RECT 127.500 744.600 129.300 749.400 ;
        RECT 130.500 744.000 132.300 747.600 ;
        RECT 143.400 744.600 145.200 752.400 ;
        RECT 149.100 751.500 150.900 752.400 ;
        RECT 152.700 750.600 153.600 757.800 ;
        RECT 164.100 756.000 165.900 757.800 ;
        RECT 167.400 752.700 168.600 757.800 ;
        RECT 170.100 756.000 171.900 757.800 ;
        RECT 185.100 756.150 186.900 757.950 ;
        RECT 188.850 753.750 190.050 757.950 ;
        RECT 191.100 756.150 192.900 757.950 ;
        RECT 206.100 756.150 207.900 757.950 ;
        RECT 208.950 753.750 210.150 757.950 ;
        RECT 212.100 756.150 213.900 757.950 ;
        RECT 227.100 756.150 228.900 757.950 ;
        RECT 229.950 753.750 231.150 757.950 ;
        RECT 233.100 756.150 234.900 757.950 ;
        RECT 247.950 757.800 250.050 759.900 ;
        RECT 250.950 757.800 253.050 759.900 ;
        RECT 253.950 757.800 256.050 759.900 ;
        RECT 256.950 757.800 259.050 759.900 ;
        RECT 265.950 757.800 268.050 759.900 ;
        RECT 268.950 757.800 271.050 759.900 ;
        RECT 271.950 757.800 274.050 759.900 ;
        RECT 274.950 757.800 277.050 759.900 ;
        RECT 188.850 752.700 192.600 753.750 ;
        RECT 167.400 751.800 171.600 752.700 ;
        RECT 147.900 744.000 149.700 750.600 ;
        RECT 150.900 748.800 153.600 750.600 ;
        RECT 150.900 744.600 152.700 748.800 ;
        RECT 164.700 744.000 166.500 750.600 ;
        RECT 169.800 744.600 171.600 751.800 ;
        RECT 182.400 749.700 190.200 751.050 ;
        RECT 182.400 744.600 184.200 749.700 ;
        RECT 185.400 744.000 187.200 748.800 ;
        RECT 188.400 744.600 190.200 749.700 ;
        RECT 191.400 750.600 192.600 752.700 ;
        RECT 206.400 752.700 210.150 753.750 ;
        RECT 227.400 752.700 231.150 753.750 ;
        RECT 248.700 754.200 249.600 757.800 ;
        RECT 251.100 756.000 252.900 757.800 ;
        RECT 257.100 756.000 258.900 757.800 ;
        RECT 266.100 756.000 267.900 757.800 ;
        RECT 272.100 756.000 273.900 757.800 ;
        RECT 275.400 754.200 276.300 757.800 ;
        RECT 281.550 757.050 282.450 761.550 ;
        RECT 290.100 759.900 291.900 761.700 ;
        RECT 296.700 759.900 297.600 767.400 ;
        RECT 311.700 759.900 312.600 772.200 ;
        RECT 331.800 767.400 333.600 779.400 ;
        RECT 334.800 768.300 336.600 779.400 ;
        RECT 337.800 769.200 339.600 780.000 ;
        RECT 340.800 768.300 342.600 779.400 ;
        RECT 352.800 773.400 354.600 779.400 ;
        RECT 355.800 774.000 357.600 780.000 ;
        RECT 334.800 767.400 342.600 768.300 ;
        RECT 353.700 773.100 354.600 773.400 ;
        RECT 358.800 773.400 360.600 779.400 ;
        RECT 361.800 773.400 363.600 780.000 ;
        RECT 373.800 773.400 375.600 780.000 ;
        RECT 376.800 773.400 378.600 779.400 ;
        RECT 379.800 773.400 381.600 780.000 ;
        RECT 391.800 773.400 393.600 779.400 ;
        RECT 394.800 774.000 396.600 780.000 ;
        RECT 358.800 773.100 360.300 773.400 ;
        RECT 353.700 772.200 360.300 773.100 ;
        RECT 313.950 765.450 316.050 766.050 ;
        RECT 325.950 765.450 328.050 766.050 ;
        RECT 313.950 764.550 328.050 765.450 ;
        RECT 313.950 763.950 316.050 764.550 ;
        RECT 325.950 763.950 328.050 764.550 ;
        RECT 317.100 759.900 318.900 761.700 ;
        RECT 332.400 759.900 333.300 767.400 ;
        RECT 338.100 759.900 339.900 761.700 ;
        RECT 353.700 759.900 354.600 772.200 ;
        RECT 358.950 768.450 361.050 769.050 ;
        RECT 373.950 768.450 376.050 769.050 ;
        RECT 358.950 767.550 376.050 768.450 ;
        RECT 358.950 766.950 361.050 767.550 ;
        RECT 373.950 766.950 376.050 767.550 ;
        RECT 355.950 765.450 358.050 766.050 ;
        RECT 355.950 764.550 363.450 765.450 ;
        RECT 355.950 763.950 358.050 764.550 ;
        RECT 362.550 762.450 363.450 764.550 ;
        RECT 359.100 759.900 360.900 761.700 ;
        RECT 362.550 761.550 369.450 762.450 ;
        RECT 286.950 757.800 289.050 759.900 ;
        RECT 289.950 757.800 292.050 759.900 ;
        RECT 292.950 757.800 295.050 759.900 ;
        RECT 295.950 757.800 298.050 759.900 ;
        RECT 310.950 757.800 313.050 759.900 ;
        RECT 313.950 757.800 316.050 759.900 ;
        RECT 316.950 757.800 319.050 759.900 ;
        RECT 319.950 757.800 322.050 759.900 ;
        RECT 331.950 757.800 334.050 759.900 ;
        RECT 334.950 757.800 337.050 759.900 ;
        RECT 337.950 757.800 340.050 759.900 ;
        RECT 340.950 757.800 343.050 759.900 ;
        RECT 352.950 757.800 355.050 759.900 ;
        RECT 355.950 757.800 358.050 759.900 ;
        RECT 358.950 757.800 361.050 759.900 ;
        RECT 361.950 757.800 364.050 759.900 ;
        RECT 277.950 755.550 282.450 757.050 ;
        RECT 287.100 756.000 288.900 757.800 ;
        RECT 293.100 756.000 294.900 757.800 ;
        RECT 277.950 754.950 282.000 755.550 ;
        RECT 248.700 753.000 252.000 754.200 ;
        RECT 206.400 750.600 207.600 752.700 ;
        RECT 191.400 744.600 193.200 750.600 ;
        RECT 205.800 744.600 207.600 750.600 ;
        RECT 208.800 749.700 216.600 751.050 ;
        RECT 227.400 750.600 228.600 752.700 ;
        RECT 208.800 744.600 210.600 749.700 ;
        RECT 211.800 744.000 213.600 748.800 ;
        RECT 214.800 744.600 216.600 749.700 ;
        RECT 226.800 744.600 228.600 750.600 ;
        RECT 229.800 749.700 237.600 751.050 ;
        RECT 229.800 744.600 231.600 749.700 ;
        RECT 232.800 744.000 234.600 748.800 ;
        RECT 235.800 744.600 237.600 749.700 ;
        RECT 250.200 744.600 252.000 753.000 ;
        RECT 256.800 744.000 258.600 753.600 ;
        RECT 266.400 744.000 268.200 753.600 ;
        RECT 273.000 753.000 276.300 754.200 ;
        RECT 273.000 744.600 274.800 753.000 ;
        RECT 296.700 750.600 297.600 757.800 ;
        RECT 311.700 754.200 312.600 757.800 ;
        RECT 314.100 756.000 315.900 757.800 ;
        RECT 320.100 756.000 321.900 757.800 ;
        RECT 311.700 753.000 315.000 754.200 ;
        RECT 288.000 744.000 289.800 750.600 ;
        RECT 292.500 749.400 297.600 750.600 ;
        RECT 292.500 744.600 294.300 749.400 ;
        RECT 295.500 744.000 297.300 747.600 ;
        RECT 313.200 744.600 315.000 753.000 ;
        RECT 319.800 744.000 321.600 753.600 ;
        RECT 332.400 750.600 333.300 757.800 ;
        RECT 335.100 756.000 336.900 757.800 ;
        RECT 341.100 756.000 342.900 757.800 ;
        RECT 353.700 754.200 354.600 757.800 ;
        RECT 356.100 756.000 357.900 757.800 ;
        RECT 362.100 756.000 363.900 757.800 ;
        RECT 368.550 757.050 369.450 761.550 ;
        RECT 377.400 759.900 378.600 773.400 ;
        RECT 392.700 773.100 393.600 773.400 ;
        RECT 397.800 773.400 399.600 779.400 ;
        RECT 400.800 773.400 402.600 780.000 ;
        RECT 410.400 773.400 412.200 780.000 ;
        RECT 413.400 773.400 415.200 779.400 ;
        RECT 416.400 773.400 418.200 780.000 ;
        RECT 428.400 773.400 430.200 780.000 ;
        RECT 431.400 773.400 433.200 779.400 ;
        RECT 434.400 774.000 436.200 780.000 ;
        RECT 397.800 773.100 399.300 773.400 ;
        RECT 392.700 772.200 399.300 773.100 ;
        RECT 379.950 762.450 382.050 763.050 ;
        RECT 385.950 762.450 388.050 763.050 ;
        RECT 379.950 761.550 388.050 762.450 ;
        RECT 379.950 760.950 382.050 761.550 ;
        RECT 385.950 760.950 388.050 761.550 ;
        RECT 392.700 759.900 393.600 772.200 ;
        RECT 394.950 765.450 397.050 766.050 ;
        RECT 403.950 765.450 406.050 766.050 ;
        RECT 394.950 764.550 406.050 765.450 ;
        RECT 394.950 763.950 397.050 764.550 ;
        RECT 403.950 763.950 406.050 764.550 ;
        RECT 398.100 759.900 399.900 761.700 ;
        RECT 413.400 759.900 414.600 773.400 ;
        RECT 431.700 773.100 433.200 773.400 ;
        RECT 437.400 773.400 439.200 779.400 ;
        RECT 437.400 773.100 438.300 773.400 ;
        RECT 431.700 772.200 438.300 773.100 ;
        RECT 415.950 771.450 418.050 772.050 ;
        RECT 427.950 771.450 430.050 772.050 ;
        RECT 415.950 770.550 430.050 771.450 ;
        RECT 415.950 769.950 418.050 770.550 ;
        RECT 427.950 769.950 430.050 770.550 ;
        RECT 427.950 762.450 430.050 763.050 ;
        RECT 422.550 761.550 430.050 762.450 ;
        RECT 373.950 757.800 376.050 759.900 ;
        RECT 376.950 757.800 379.050 759.900 ;
        RECT 379.950 757.800 382.050 759.900 ;
        RECT 391.950 757.800 394.050 759.900 ;
        RECT 394.950 757.800 397.050 759.900 ;
        RECT 397.950 757.800 400.050 759.900 ;
        RECT 400.950 757.800 403.050 759.900 ;
        RECT 409.950 757.800 412.050 759.900 ;
        RECT 412.950 757.800 415.050 759.900 ;
        RECT 415.950 757.800 418.050 759.900 ;
        RECT 368.550 755.550 373.050 757.050 ;
        RECT 374.100 756.000 375.900 757.800 ;
        RECT 369.000 754.950 373.050 755.550 ;
        RECT 353.700 753.000 357.000 754.200 ;
        RECT 332.400 749.400 337.500 750.600 ;
        RECT 332.700 744.000 334.500 747.600 ;
        RECT 335.700 744.600 337.500 749.400 ;
        RECT 340.200 744.000 342.000 750.600 ;
        RECT 355.200 744.600 357.000 753.000 ;
        RECT 361.800 744.000 363.600 753.600 ;
        RECT 377.400 752.700 378.600 757.800 ;
        RECT 380.100 756.000 381.900 757.800 ;
        RECT 392.700 754.200 393.600 757.800 ;
        RECT 395.100 756.000 396.900 757.800 ;
        RECT 401.100 756.000 402.900 757.800 ;
        RECT 410.100 756.000 411.900 757.800 ;
        RECT 392.700 753.000 396.000 754.200 ;
        RECT 374.400 751.800 378.600 752.700 ;
        RECT 374.400 744.600 376.200 751.800 ;
        RECT 379.500 744.000 381.300 750.600 ;
        RECT 394.200 744.600 396.000 753.000 ;
        RECT 400.800 744.000 402.600 753.600 ;
        RECT 413.400 752.700 414.600 757.800 ;
        RECT 416.100 756.000 417.900 757.800 ;
        RECT 422.550 757.050 423.450 761.550 ;
        RECT 427.950 760.950 430.050 761.550 ;
        RECT 431.100 759.900 432.900 761.700 ;
        RECT 437.400 759.900 438.300 772.200 ;
        RECT 451.800 767.400 453.600 779.400 ;
        RECT 454.800 768.300 456.600 779.400 ;
        RECT 457.800 769.200 459.600 780.000 ;
        RECT 460.800 768.300 462.600 779.400 ;
        RECT 472.800 773.400 474.600 779.400 ;
        RECT 475.800 774.000 477.600 780.000 ;
        RECT 454.800 767.400 462.600 768.300 ;
        RECT 473.700 773.100 474.600 773.400 ;
        RECT 478.800 773.400 480.600 779.400 ;
        RECT 481.800 773.400 483.600 780.000 ;
        RECT 478.800 773.100 480.300 773.400 ;
        RECT 473.700 772.200 480.300 773.100 ;
        RECT 452.400 759.900 453.300 767.400 ;
        RECT 454.950 765.450 457.050 766.050 ;
        RECT 466.950 765.450 469.050 766.050 ;
        RECT 454.950 764.550 469.050 765.450 ;
        RECT 454.950 763.950 457.050 764.550 ;
        RECT 466.950 763.950 469.050 764.550 ;
        RECT 458.100 759.900 459.900 761.700 ;
        RECT 473.700 759.900 474.600 772.200 ;
        RECT 481.950 771.450 484.050 772.050 ;
        RECT 487.950 771.450 490.050 772.050 ;
        RECT 481.950 770.550 490.050 771.450 ;
        RECT 481.950 769.950 484.050 770.550 ;
        RECT 487.950 769.950 490.050 770.550 ;
        RECT 493.800 767.400 495.600 779.400 ;
        RECT 496.800 768.300 498.600 779.400 ;
        RECT 499.800 769.200 501.600 780.000 ;
        RECT 502.800 768.300 504.600 779.400 ;
        RECT 514.800 773.400 516.600 779.400 ;
        RECT 517.800 774.000 519.600 780.000 ;
        RECT 496.800 767.400 504.600 768.300 ;
        RECT 515.700 773.100 516.600 773.400 ;
        RECT 520.800 773.400 522.600 779.400 ;
        RECT 523.800 773.400 525.600 780.000 ;
        RECT 520.800 773.100 522.300 773.400 ;
        RECT 515.700 772.200 522.300 773.100 ;
        RECT 479.100 759.900 480.900 761.700 ;
        RECT 494.400 759.900 495.300 767.400 ;
        RECT 500.100 759.900 501.900 761.700 ;
        RECT 515.700 759.900 516.600 772.200 ;
        RECT 533.700 767.400 535.500 780.000 ;
        RECT 538.800 773.400 540.600 779.400 ;
        RECT 541.800 773.400 543.600 780.000 ;
        RECT 521.100 759.900 522.900 761.700 ;
        RECT 533.100 760.050 534.900 761.850 ;
        RECT 538.950 760.050 540.150 773.400 ;
        RECT 556.800 767.400 558.600 779.400 ;
        RECT 559.800 773.400 561.600 780.000 ;
        RECT 562.800 773.400 564.600 779.400 ;
        RECT 565.800 773.400 567.600 780.000 ;
        RECT 577.800 778.500 585.600 779.400 ;
        RECT 550.950 763.950 553.050 766.050 ;
        RECT 427.950 757.800 430.050 759.900 ;
        RECT 430.950 757.800 433.050 759.900 ;
        RECT 433.950 757.800 436.050 759.900 ;
        RECT 436.950 757.800 439.050 759.900 ;
        RECT 451.950 757.800 454.050 759.900 ;
        RECT 454.950 757.800 457.050 759.900 ;
        RECT 457.950 757.800 460.050 759.900 ;
        RECT 460.950 757.800 463.050 759.900 ;
        RECT 472.950 757.800 475.050 759.900 ;
        RECT 475.950 757.800 478.050 759.900 ;
        RECT 478.950 757.800 481.050 759.900 ;
        RECT 481.950 757.800 484.050 759.900 ;
        RECT 493.950 757.800 496.050 759.900 ;
        RECT 496.950 757.800 499.050 759.900 ;
        RECT 499.950 757.800 502.050 759.900 ;
        RECT 502.950 757.800 505.050 759.900 ;
        RECT 514.950 757.800 517.050 759.900 ;
        RECT 517.950 757.800 520.050 759.900 ;
        RECT 520.950 757.800 523.050 759.900 ;
        RECT 523.950 757.800 526.050 759.900 ;
        RECT 532.950 757.950 535.050 760.050 ;
        RECT 535.950 757.950 538.050 760.050 ;
        RECT 538.950 757.950 541.050 760.050 ;
        RECT 541.950 757.950 544.050 760.050 ;
        RECT 422.550 755.550 427.050 757.050 ;
        RECT 428.100 756.000 429.900 757.800 ;
        RECT 434.100 756.000 435.900 757.800 ;
        RECT 423.000 754.950 427.050 755.550 ;
        RECT 437.400 754.200 438.300 757.800 ;
        RECT 413.400 751.800 417.600 752.700 ;
        RECT 410.700 744.000 412.500 750.600 ;
        RECT 415.800 744.600 417.600 751.800 ;
        RECT 428.400 744.000 430.200 753.600 ;
        RECT 435.000 753.000 438.300 754.200 ;
        RECT 435.000 744.600 436.800 753.000 ;
        RECT 452.400 750.600 453.300 757.800 ;
        RECT 455.100 756.000 456.900 757.800 ;
        RECT 461.100 756.000 462.900 757.800 ;
        RECT 473.700 754.200 474.600 757.800 ;
        RECT 476.100 756.000 477.900 757.800 ;
        RECT 482.100 756.000 483.900 757.800 ;
        RECT 473.700 753.000 477.000 754.200 ;
        RECT 452.400 749.400 457.500 750.600 ;
        RECT 452.700 744.000 454.500 747.600 ;
        RECT 455.700 744.600 457.500 749.400 ;
        RECT 460.200 744.000 462.000 750.600 ;
        RECT 475.200 744.600 477.000 753.000 ;
        RECT 481.800 744.000 483.600 753.600 ;
        RECT 494.400 750.600 495.300 757.800 ;
        RECT 497.100 756.000 498.900 757.800 ;
        RECT 503.100 756.000 504.900 757.800 ;
        RECT 515.700 754.200 516.600 757.800 ;
        RECT 518.100 756.000 519.900 757.800 ;
        RECT 524.100 756.000 525.900 757.800 ;
        RECT 536.100 756.150 537.900 757.950 ;
        RECT 499.950 753.450 502.050 753.600 ;
        RECT 511.950 753.450 514.050 754.050 ;
        RECT 499.950 752.550 514.050 753.450 ;
        RECT 515.700 753.000 519.000 754.200 ;
        RECT 539.850 753.750 541.050 757.950 ;
        RECT 542.100 756.150 543.900 757.950 ;
        RECT 544.950 756.450 547.050 757.050 ;
        RECT 551.550 756.450 552.450 763.950 ;
        RECT 557.400 759.900 558.300 767.400 ;
        RECT 560.100 759.900 561.900 761.700 ;
        RECT 556.950 757.800 559.050 759.900 ;
        RECT 559.950 757.800 562.050 759.900 ;
        RECT 544.950 755.550 552.450 756.450 ;
        RECT 544.950 754.950 547.050 755.550 ;
        RECT 499.950 751.500 502.050 752.550 ;
        RECT 511.950 751.950 514.050 752.550 ;
        RECT 494.400 749.400 499.500 750.600 ;
        RECT 494.700 744.000 496.500 747.600 ;
        RECT 497.700 744.600 499.500 749.400 ;
        RECT 502.200 744.000 504.000 750.600 ;
        RECT 517.200 744.600 519.000 753.000 ;
        RECT 523.800 744.000 525.600 753.600 ;
        RECT 539.850 752.700 543.600 753.750 ;
        RECT 533.400 749.700 541.200 751.050 ;
        RECT 533.400 744.600 535.200 749.700 ;
        RECT 536.400 744.000 538.200 748.800 ;
        RECT 539.400 744.600 541.200 749.700 ;
        RECT 542.400 750.600 543.600 752.700 ;
        RECT 557.400 750.600 558.300 757.800 ;
        RECT 563.700 753.300 564.600 773.400 ;
        RECT 577.800 767.400 579.600 778.500 ;
        RECT 580.800 766.500 582.600 777.600 ;
        RECT 583.800 768.600 585.600 778.500 ;
        RECT 586.800 769.500 588.600 780.000 ;
        RECT 589.800 768.600 591.600 779.400 ;
        RECT 601.800 773.400 603.600 780.000 ;
        RECT 604.800 773.400 606.600 779.400 ;
        RECT 607.800 773.400 609.600 780.000 ;
        RECT 583.800 767.700 591.600 768.600 ;
        RECT 580.800 765.600 585.900 766.500 ;
        RECT 577.950 762.450 580.050 763.050 ;
        RECT 572.550 761.550 580.050 762.450 ;
        RECT 565.950 757.800 568.050 759.900 ;
        RECT 566.100 756.000 567.900 757.800 ;
        RECT 572.550 757.050 573.450 761.550 ;
        RECT 577.950 760.950 580.050 761.550 ;
        RECT 581.100 759.900 582.900 761.700 ;
        RECT 585.000 759.900 585.900 765.600 ;
        RECT 589.950 765.450 592.050 766.050 ;
        RECT 598.950 765.450 601.050 766.050 ;
        RECT 589.950 764.550 601.050 765.450 ;
        RECT 589.950 763.950 592.050 764.550 ;
        RECT 598.950 763.950 601.050 764.550 ;
        RECT 589.950 762.450 592.050 762.900 ;
        RECT 595.950 762.450 598.050 763.050 ;
        RECT 587.100 759.900 588.900 761.700 ;
        RECT 589.950 761.550 598.050 762.450 ;
        RECT 589.950 760.800 592.050 761.550 ;
        RECT 595.950 760.950 598.050 761.550 ;
        RECT 605.400 759.900 606.600 773.400 ;
        RECT 617.400 767.400 619.200 780.000 ;
        RECT 622.500 768.600 624.300 779.400 ;
        RECT 637.800 773.400 639.600 780.000 ;
        RECT 640.800 773.400 642.600 779.400 ;
        RECT 643.800 773.400 645.600 780.000 ;
        RECT 656.400 773.400 658.200 780.000 ;
        RECT 659.400 773.400 661.200 779.400 ;
        RECT 620.700 767.400 624.300 768.600 ;
        RECT 617.100 760.050 618.900 761.850 ;
        RECT 620.700 760.050 621.600 767.400 ;
        RECT 631.950 762.450 634.050 763.050 ;
        RECT 637.950 762.450 640.050 763.050 ;
        RECT 623.100 760.050 624.900 761.850 ;
        RECT 631.950 761.550 640.050 762.450 ;
        RECT 631.950 760.950 634.050 761.550 ;
        RECT 637.950 760.950 640.050 761.550 ;
        RECT 577.950 757.800 580.050 759.900 ;
        RECT 580.950 757.800 583.050 759.900 ;
        RECT 583.950 757.800 586.050 759.900 ;
        RECT 586.950 757.800 589.050 759.900 ;
        RECT 589.950 757.800 592.050 759.900 ;
        RECT 601.950 757.800 604.050 759.900 ;
        RECT 604.950 757.800 607.050 759.900 ;
        RECT 607.950 757.800 610.050 759.900 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 622.950 757.950 625.050 760.050 ;
        RECT 641.400 759.900 642.600 773.400 ;
        RECT 659.850 760.050 661.050 773.400 ;
        RECT 664.500 767.400 666.300 780.000 ;
        RECT 674.400 767.400 676.200 780.000 ;
        RECT 679.500 768.600 681.300 779.400 ;
        RECT 695.400 773.400 697.200 780.000 ;
        RECT 698.400 773.400 700.200 779.400 ;
        RECT 677.700 767.400 681.300 768.600 ;
        RECT 665.100 760.050 666.900 761.850 ;
        RECT 674.100 760.050 675.900 761.850 ;
        RECT 677.700 760.050 678.600 767.400 ;
        RECT 682.950 762.450 685.050 763.050 ;
        RECT 680.100 760.050 681.900 761.850 ;
        RECT 682.950 761.550 690.450 762.450 ;
        RECT 682.950 760.950 685.050 761.550 ;
        RECT 568.950 755.550 573.450 757.050 ;
        RECT 578.100 756.000 579.900 757.800 ;
        RECT 568.950 754.950 573.000 755.550 ;
        RECT 560.100 752.400 567.600 753.300 ;
        RECT 560.100 751.500 561.900 752.400 ;
        RECT 542.400 744.600 544.200 750.600 ;
        RECT 557.400 748.800 560.100 750.600 ;
        RECT 558.300 744.600 560.100 748.800 ;
        RECT 561.300 744.000 563.100 750.600 ;
        RECT 565.800 744.600 567.600 752.400 ;
        RECT 585.000 750.600 586.050 757.800 ;
        RECT 590.100 756.000 591.900 757.800 ;
        RECT 602.100 756.000 603.900 757.800 ;
        RECT 605.400 752.700 606.600 757.800 ;
        RECT 608.100 756.000 609.900 757.800 ;
        RECT 602.400 751.800 606.600 752.700 ;
        RECT 580.500 744.000 582.300 750.600 ;
        RECT 585.000 744.600 586.800 750.600 ;
        RECT 589.500 744.000 591.300 750.600 ;
        RECT 602.400 744.600 604.200 751.800 ;
        RECT 607.500 744.000 609.300 750.600 ;
        RECT 620.700 747.600 621.600 757.950 ;
        RECT 637.950 757.800 640.050 759.900 ;
        RECT 640.950 757.800 643.050 759.900 ;
        RECT 643.950 757.800 646.050 759.900 ;
        RECT 655.950 757.950 658.050 760.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 673.950 757.950 676.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 679.950 757.950 682.050 760.050 ;
        RECT 638.100 756.000 639.900 757.800 ;
        RECT 641.400 752.700 642.600 757.800 ;
        RECT 644.100 756.000 645.900 757.800 ;
        RECT 656.100 756.150 657.900 757.950 ;
        RECT 658.950 753.750 660.150 757.950 ;
        RECT 662.100 756.150 663.900 757.950 ;
        RECT 638.400 751.800 642.600 752.700 ;
        RECT 656.400 752.700 660.150 753.750 ;
        RECT 617.400 744.000 619.200 747.600 ;
        RECT 620.400 744.600 622.200 747.600 ;
        RECT 623.400 744.000 625.200 747.600 ;
        RECT 638.400 744.600 640.200 751.800 ;
        RECT 656.400 750.600 657.600 752.700 ;
        RECT 643.500 744.000 645.300 750.600 ;
        RECT 655.800 744.600 657.600 750.600 ;
        RECT 658.800 749.700 666.600 751.050 ;
        RECT 658.800 744.600 660.600 749.700 ;
        RECT 661.800 744.000 663.600 748.800 ;
        RECT 664.800 744.600 666.600 749.700 ;
        RECT 677.700 747.600 678.600 757.950 ;
        RECT 689.550 757.050 690.450 761.550 ;
        RECT 698.850 760.050 700.050 773.400 ;
        RECT 703.500 767.400 705.300 780.000 ;
        RECT 716.700 768.600 718.500 779.400 ;
        RECT 716.700 767.400 720.300 768.600 ;
        RECT 721.800 767.400 723.600 780.000 ;
        RECT 731.400 773.400 733.200 780.000 ;
        RECT 734.400 773.400 736.200 779.400 ;
        RECT 737.400 773.400 739.200 780.000 ;
        RECT 749.400 773.400 751.200 780.000 ;
        RECT 752.400 773.400 754.200 779.400 ;
        RECT 755.400 774.000 757.200 780.000 ;
        RECT 704.100 760.050 705.900 761.850 ;
        RECT 716.100 760.050 717.900 761.850 ;
        RECT 719.400 760.050 720.300 767.400 ;
        RECT 722.100 760.050 723.900 761.850 ;
        RECT 694.950 757.950 697.050 760.050 ;
        RECT 697.950 757.950 700.050 760.050 ;
        RECT 700.950 757.950 703.050 760.050 ;
        RECT 703.950 757.950 706.050 760.050 ;
        RECT 715.950 757.950 718.050 760.050 ;
        RECT 718.950 757.950 721.050 760.050 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 734.400 759.900 735.600 773.400 ;
        RECT 752.700 773.100 754.200 773.400 ;
        RECT 758.400 773.400 760.200 779.400 ;
        RECT 770.400 773.400 772.200 780.000 ;
        RECT 773.400 773.400 775.200 779.400 ;
        RECT 776.400 774.000 778.200 780.000 ;
        RECT 758.400 773.100 759.300 773.400 ;
        RECT 752.700 772.200 759.300 773.100 ;
        RECT 773.700 773.100 775.200 773.400 ;
        RECT 779.400 773.400 781.200 779.400 ;
        RECT 779.400 773.100 780.300 773.400 ;
        RECT 773.700 772.200 780.300 773.100 ;
        RECT 744.000 762.450 748.050 763.050 ;
        RECT 743.550 760.950 748.050 762.450 ;
        RECT 689.550 755.550 694.050 757.050 ;
        RECT 695.100 756.150 696.900 757.950 ;
        RECT 690.000 754.950 694.050 755.550 ;
        RECT 697.950 753.750 699.150 757.950 ;
        RECT 701.100 756.150 702.900 757.950 ;
        RECT 695.400 752.700 699.150 753.750 ;
        RECT 695.400 750.600 696.600 752.700 ;
        RECT 674.400 744.000 676.200 747.600 ;
        RECT 677.400 744.600 679.200 747.600 ;
        RECT 680.400 744.000 682.200 747.600 ;
        RECT 694.800 744.600 696.600 750.600 ;
        RECT 697.800 749.700 705.600 751.050 ;
        RECT 697.800 744.600 699.600 749.700 ;
        RECT 700.800 744.000 702.600 748.800 ;
        RECT 703.800 744.600 705.600 749.700 ;
        RECT 719.400 747.600 720.300 757.950 ;
        RECT 730.950 757.800 733.050 759.900 ;
        RECT 733.950 757.800 736.050 759.900 ;
        RECT 736.950 757.800 739.050 759.900 ;
        RECT 731.100 756.000 732.900 757.800 ;
        RECT 721.950 753.450 724.050 754.050 ;
        RECT 727.950 753.450 730.050 754.050 ;
        RECT 721.950 752.550 730.050 753.450 ;
        RECT 721.950 751.950 724.050 752.550 ;
        RECT 727.950 751.950 730.050 752.550 ;
        RECT 734.400 752.700 735.600 757.800 ;
        RECT 737.100 756.000 738.900 757.800 ;
        RECT 743.550 757.050 744.450 760.950 ;
        RECT 752.100 759.900 753.900 761.700 ;
        RECT 758.400 759.900 759.300 772.200 ;
        RECT 773.100 759.900 774.900 761.700 ;
        RECT 779.400 759.900 780.300 772.200 ;
        RECT 793.800 767.400 795.600 779.400 ;
        RECT 796.800 768.300 798.600 779.400 ;
        RECT 799.800 769.200 801.600 780.000 ;
        RECT 802.800 768.300 804.600 779.400 ;
        RECT 812.400 773.400 814.200 780.000 ;
        RECT 815.400 773.400 817.200 779.400 ;
        RECT 818.400 773.400 820.200 780.000 ;
        RECT 830.400 773.400 832.200 780.000 ;
        RECT 833.400 773.400 835.200 779.400 ;
        RECT 836.400 774.000 838.200 780.000 ;
        RECT 796.800 767.400 804.600 768.300 ;
        RECT 794.400 759.900 795.300 767.400 ;
        RECT 796.950 765.450 799.050 766.050 ;
        RECT 802.950 765.450 805.050 766.050 ;
        RECT 796.950 764.550 805.050 765.450 ;
        RECT 796.950 763.950 799.050 764.550 ;
        RECT 802.950 763.950 805.050 764.550 ;
        RECT 800.100 759.900 801.900 761.700 ;
        RECT 815.400 759.900 816.600 773.400 ;
        RECT 833.700 773.100 835.200 773.400 ;
        RECT 839.400 773.400 841.200 779.400 ;
        RECT 851.400 773.400 853.200 780.000 ;
        RECT 854.400 773.400 856.200 779.400 ;
        RECT 839.400 773.100 840.300 773.400 ;
        RECT 833.700 772.200 840.300 773.100 ;
        RECT 820.950 765.450 823.050 766.050 ;
        RECT 835.950 765.450 838.050 766.050 ;
        RECT 820.950 764.550 838.050 765.450 ;
        RECT 820.950 763.950 823.050 764.550 ;
        RECT 835.950 763.950 838.050 764.550 ;
        RECT 825.000 762.450 829.050 763.050 ;
        RECT 824.550 760.950 829.050 762.450 ;
        RECT 748.950 757.800 751.050 759.900 ;
        RECT 751.950 757.800 754.050 759.900 ;
        RECT 754.950 757.800 757.050 759.900 ;
        RECT 757.950 757.800 760.050 759.900 ;
        RECT 769.950 757.800 772.050 759.900 ;
        RECT 772.950 757.800 775.050 759.900 ;
        RECT 775.950 757.800 778.050 759.900 ;
        RECT 778.950 757.800 781.050 759.900 ;
        RECT 793.950 757.800 796.050 759.900 ;
        RECT 796.950 757.800 799.050 759.900 ;
        RECT 799.950 757.800 802.050 759.900 ;
        RECT 802.950 757.800 805.050 759.900 ;
        RECT 811.950 757.800 814.050 759.900 ;
        RECT 814.950 757.800 817.050 759.900 ;
        RECT 817.950 757.800 820.050 759.900 ;
        RECT 739.950 755.550 744.450 757.050 ;
        RECT 749.100 756.000 750.900 757.800 ;
        RECT 755.100 756.000 756.900 757.800 ;
        RECT 739.950 754.950 744.000 755.550 ;
        RECT 758.400 754.200 759.300 757.800 ;
        RECT 770.100 756.000 771.900 757.800 ;
        RECT 776.100 756.000 777.900 757.800 ;
        RECT 779.400 754.200 780.300 757.800 ;
        RECT 781.950 756.450 784.050 757.050 ;
        RECT 787.950 756.450 790.050 757.050 ;
        RECT 781.950 755.550 790.050 756.450 ;
        RECT 781.950 754.950 784.050 755.550 ;
        RECT 787.950 754.950 790.050 755.550 ;
        RECT 734.400 751.800 738.600 752.700 ;
        RECT 715.800 744.000 717.600 747.600 ;
        RECT 718.800 744.600 720.600 747.600 ;
        RECT 721.800 744.000 723.600 747.600 ;
        RECT 731.700 744.000 733.500 750.600 ;
        RECT 736.800 744.600 738.600 751.800 ;
        RECT 749.400 744.000 751.200 753.600 ;
        RECT 756.000 753.000 759.300 754.200 ;
        RECT 756.000 744.600 757.800 753.000 ;
        RECT 770.400 744.000 772.200 753.600 ;
        RECT 777.000 753.000 780.300 754.200 ;
        RECT 777.000 744.600 778.800 753.000 ;
        RECT 794.400 750.600 795.300 757.800 ;
        RECT 797.100 756.000 798.900 757.800 ;
        RECT 803.100 756.000 804.900 757.800 ;
        RECT 812.100 756.000 813.900 757.800 ;
        RECT 815.400 752.700 816.600 757.800 ;
        RECT 818.100 756.000 819.900 757.800 ;
        RECT 824.550 757.050 825.450 760.950 ;
        RECT 833.100 759.900 834.900 761.700 ;
        RECT 839.400 759.900 840.300 772.200 ;
        RECT 851.100 760.050 852.900 761.850 ;
        RECT 854.400 760.050 855.600 773.400 ;
        RECT 829.950 757.800 832.050 759.900 ;
        RECT 832.950 757.800 835.050 759.900 ;
        RECT 835.950 757.800 838.050 759.900 ;
        RECT 838.950 757.800 841.050 759.900 ;
        RECT 850.950 757.950 853.050 760.050 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 824.550 755.550 829.050 757.050 ;
        RECT 830.100 756.000 831.900 757.800 ;
        RECT 836.100 756.000 837.900 757.800 ;
        RECT 825.000 754.950 829.050 755.550 ;
        RECT 839.400 754.200 840.300 757.800 ;
        RECT 815.400 751.800 819.600 752.700 ;
        RECT 794.400 749.400 799.500 750.600 ;
        RECT 794.700 744.000 796.500 747.600 ;
        RECT 797.700 744.600 799.500 749.400 ;
        RECT 802.200 744.000 804.000 750.600 ;
        RECT 812.700 744.000 814.500 750.600 ;
        RECT 817.800 744.600 819.600 751.800 ;
        RECT 830.400 744.000 832.200 753.600 ;
        RECT 837.000 753.000 840.300 754.200 ;
        RECT 837.000 744.600 838.800 753.000 ;
        RECT 854.400 747.600 855.600 757.950 ;
        RECT 851.400 744.000 853.200 747.600 ;
        RECT 854.400 744.600 856.200 747.600 ;
        RECT 13.200 732.000 15.000 740.400 ;
        RECT 11.700 730.800 15.000 732.000 ;
        RECT 19.800 731.400 21.600 741.000 ;
        RECT 30.000 734.400 31.800 741.000 ;
        RECT 34.500 735.600 36.300 740.400 ;
        RECT 37.500 737.400 39.300 741.000 ;
        RECT 34.500 734.400 39.600 735.600 ;
        RECT 11.700 727.200 12.600 730.800 ;
        RECT 14.100 727.200 15.900 729.000 ;
        RECT 20.100 727.200 21.900 729.000 ;
        RECT 29.100 727.200 30.900 729.000 ;
        RECT 35.100 727.200 36.900 729.000 ;
        RECT 38.700 727.200 39.600 734.400 ;
        RECT 55.200 732.000 57.000 740.400 ;
        RECT 53.700 730.800 57.000 732.000 ;
        RECT 61.800 731.400 63.600 741.000 ;
        RECT 76.200 732.000 78.000 740.400 ;
        RECT 74.700 730.800 78.000 732.000 ;
        RECT 82.800 731.400 84.600 741.000 ;
        RECT 93.000 734.400 94.800 741.000 ;
        RECT 97.500 735.600 99.300 740.400 ;
        RECT 100.500 737.400 102.300 741.000 ;
        RECT 97.500 734.400 102.600 735.600 ;
        RECT 115.800 734.400 117.600 740.400 ;
        RECT 53.700 727.200 54.600 730.800 ;
        RECT 69.000 729.450 73.050 730.050 ;
        RECT 56.100 727.200 57.900 729.000 ;
        RECT 62.100 727.200 63.900 729.000 ;
        RECT 68.550 727.950 73.050 729.450 ;
        RECT 10.950 725.100 13.050 727.200 ;
        RECT 13.950 725.100 16.050 727.200 ;
        RECT 16.950 725.100 19.050 727.200 ;
        RECT 19.950 725.100 22.050 727.200 ;
        RECT 28.950 725.100 31.050 727.200 ;
        RECT 31.950 725.100 34.050 727.200 ;
        RECT 34.950 725.100 37.050 727.200 ;
        RECT 37.950 725.100 40.050 727.200 ;
        RECT 52.950 725.100 55.050 727.200 ;
        RECT 55.950 725.100 58.050 727.200 ;
        RECT 58.950 725.100 61.050 727.200 ;
        RECT 61.950 725.100 64.050 727.200 ;
        RECT 11.700 712.800 12.600 725.100 ;
        RECT 17.100 723.300 18.900 725.100 ;
        RECT 32.100 723.300 33.900 725.100 ;
        RECT 38.700 717.600 39.600 725.100 ;
        RECT 29.400 716.700 37.200 717.600 ;
        RECT 11.700 711.900 18.300 712.800 ;
        RECT 11.700 711.600 12.600 711.900 ;
        RECT 10.800 705.600 12.600 711.600 ;
        RECT 16.800 711.600 18.300 711.900 ;
        RECT 13.800 705.000 15.600 711.000 ;
        RECT 16.800 705.600 18.600 711.600 ;
        RECT 19.800 705.000 21.600 711.600 ;
        RECT 29.400 705.600 31.200 716.700 ;
        RECT 32.400 705.000 34.200 715.800 ;
        RECT 35.400 705.600 37.200 716.700 ;
        RECT 38.400 705.600 40.200 717.600 ;
        RECT 53.700 712.800 54.600 725.100 ;
        RECT 59.100 723.300 60.900 725.100 ;
        RECT 61.950 723.450 64.050 724.050 ;
        RECT 68.550 723.450 69.450 727.950 ;
        RECT 74.700 727.200 75.600 730.800 ;
        RECT 77.100 727.200 78.900 729.000 ;
        RECT 83.100 727.200 84.900 729.000 ;
        RECT 92.100 727.200 93.900 729.000 ;
        RECT 98.100 727.200 99.900 729.000 ;
        RECT 101.700 727.200 102.600 734.400 ;
        RECT 116.400 732.300 117.600 734.400 ;
        RECT 118.800 735.300 120.600 740.400 ;
        RECT 121.800 736.200 123.600 741.000 ;
        RECT 124.800 735.300 126.600 740.400 ;
        RECT 118.800 733.950 126.600 735.300 ;
        RECT 136.800 734.400 138.600 740.400 ;
        RECT 137.400 732.300 138.600 734.400 ;
        RECT 139.800 735.300 141.600 740.400 ;
        RECT 142.800 736.200 144.600 741.000 ;
        RECT 145.800 735.300 147.600 740.400 ;
        RECT 139.800 733.950 147.600 735.300 ;
        RECT 155.700 734.400 157.500 741.000 ;
        RECT 160.800 733.200 162.600 740.400 ;
        RECT 158.400 732.300 162.600 733.200 ;
        RECT 173.400 737.400 175.200 740.400 ;
        RECT 176.400 737.400 178.200 741.000 ;
        RECT 173.400 733.500 174.600 737.400 ;
        RECT 179.400 734.400 181.200 740.400 ;
        RECT 192.000 734.400 193.800 741.000 ;
        RECT 196.500 735.600 198.300 740.400 ;
        RECT 199.500 737.400 201.300 741.000 ;
        RECT 196.500 734.400 201.600 735.600 ;
        RECT 173.400 732.600 179.100 733.500 ;
        RECT 116.400 731.250 120.150 732.300 ;
        RECT 137.400 731.250 141.150 732.300 ;
        RECT 103.950 729.450 106.050 730.050 ;
        RECT 103.950 728.550 111.450 729.450 ;
        RECT 103.950 727.950 106.050 728.550 ;
        RECT 73.950 725.100 76.050 727.200 ;
        RECT 76.950 725.100 79.050 727.200 ;
        RECT 79.950 725.100 82.050 727.200 ;
        RECT 82.950 725.100 85.050 727.200 ;
        RECT 91.950 725.100 94.050 727.200 ;
        RECT 94.950 725.100 97.050 727.200 ;
        RECT 97.950 725.100 100.050 727.200 ;
        RECT 100.950 725.100 103.050 727.200 ;
        RECT 61.950 722.550 69.450 723.450 ;
        RECT 61.950 721.950 64.050 722.550 ;
        RECT 74.700 712.800 75.600 725.100 ;
        RECT 80.100 723.300 81.900 725.100 ;
        RECT 95.100 723.300 96.900 725.100 ;
        RECT 82.950 720.450 85.050 721.050 ;
        RECT 97.950 720.450 100.050 721.050 ;
        RECT 82.950 719.550 100.050 720.450 ;
        RECT 82.950 718.950 85.050 719.550 ;
        RECT 97.950 718.950 100.050 719.550 ;
        RECT 101.700 717.600 102.600 725.100 ;
        RECT 110.550 724.050 111.450 728.550 ;
        RECT 116.100 727.050 117.900 728.850 ;
        RECT 118.950 727.050 120.150 731.250 ;
        RECT 122.100 727.050 123.900 728.850 ;
        RECT 137.100 727.050 138.900 728.850 ;
        RECT 139.950 727.050 141.150 731.250 ;
        RECT 143.100 727.050 144.900 728.850 ;
        RECT 155.100 727.200 156.900 729.000 ;
        RECT 158.400 727.200 159.600 732.300 ;
        RECT 177.150 731.700 179.100 732.600 ;
        RECT 163.950 729.450 168.000 730.050 ;
        RECT 161.100 727.200 162.900 729.000 ;
        RECT 163.950 727.950 168.450 729.450 ;
        RECT 115.950 724.950 118.050 727.050 ;
        RECT 118.950 724.950 121.050 727.050 ;
        RECT 121.950 724.950 124.050 727.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 136.950 724.950 139.050 727.050 ;
        RECT 139.950 724.950 142.050 727.050 ;
        RECT 142.950 724.950 145.050 727.050 ;
        RECT 145.950 724.950 148.050 727.050 ;
        RECT 154.950 725.100 157.050 727.200 ;
        RECT 157.950 725.100 160.050 727.200 ;
        RECT 160.950 725.100 163.050 727.200 ;
        RECT 110.550 722.550 115.050 724.050 ;
        RECT 111.000 721.950 115.050 722.550 ;
        RECT 92.400 716.700 100.200 717.600 ;
        RECT 53.700 711.900 60.300 712.800 ;
        RECT 53.700 711.600 54.600 711.900 ;
        RECT 52.800 705.600 54.600 711.600 ;
        RECT 58.800 711.600 60.300 711.900 ;
        RECT 74.700 711.900 81.300 712.800 ;
        RECT 74.700 711.600 75.600 711.900 ;
        RECT 55.800 705.000 57.600 711.000 ;
        RECT 58.800 705.600 60.600 711.600 ;
        RECT 61.800 705.000 63.600 711.600 ;
        RECT 73.800 705.600 75.600 711.600 ;
        RECT 79.800 711.600 81.300 711.900 ;
        RECT 76.800 705.000 78.600 711.000 ;
        RECT 79.800 705.600 81.600 711.600 ;
        RECT 82.800 705.000 84.600 711.600 ;
        RECT 92.400 705.600 94.200 716.700 ;
        RECT 95.400 705.000 97.200 715.800 ;
        RECT 98.400 705.600 100.200 716.700 ;
        RECT 101.400 705.600 103.200 717.600 ;
        RECT 119.850 711.600 121.050 724.950 ;
        RECT 125.100 723.150 126.900 724.950 ;
        RECT 116.400 705.000 118.200 711.600 ;
        RECT 119.400 705.600 121.200 711.600 ;
        RECT 124.500 705.000 126.300 717.600 ;
        RECT 140.850 711.600 142.050 724.950 ;
        RECT 146.100 723.150 147.900 724.950 ;
        RECT 137.400 705.000 139.200 711.600 ;
        RECT 140.400 705.600 142.200 711.600 ;
        RECT 145.500 705.000 147.300 717.600 ;
        RECT 158.400 711.600 159.600 725.100 ;
        RECT 167.550 724.050 168.450 727.950 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 167.550 722.550 172.050 724.050 ;
        RECT 173.100 723.150 174.900 724.950 ;
        RECT 168.000 721.950 172.050 722.550 ;
        RECT 177.150 720.300 178.050 731.700 ;
        RECT 180.000 727.050 181.200 734.400 ;
        RECT 191.100 727.200 192.900 729.000 ;
        RECT 197.100 727.200 198.900 729.000 ;
        RECT 200.700 727.200 201.600 734.400 ;
        RECT 217.200 732.000 219.000 740.400 ;
        RECT 215.700 730.800 219.000 732.000 ;
        RECT 223.800 731.400 225.600 741.000 ;
        RECT 234.000 734.400 235.800 741.000 ;
        RECT 238.500 735.600 240.300 740.400 ;
        RECT 241.500 737.400 243.300 741.000 ;
        RECT 238.500 734.400 243.600 735.600 ;
        RECT 226.950 732.450 229.050 733.050 ;
        RECT 235.950 732.450 238.050 733.050 ;
        RECT 226.950 731.550 238.050 732.450 ;
        RECT 226.950 730.950 229.050 731.550 ;
        RECT 235.950 730.950 238.050 731.550 ;
        RECT 215.700 727.200 216.600 730.800 ;
        RECT 218.100 727.200 219.900 729.000 ;
        RECT 224.100 727.200 225.900 729.000 ;
        RECT 233.100 727.200 234.900 729.000 ;
        RECT 239.100 727.200 240.900 729.000 ;
        RECT 242.700 727.200 243.600 734.400 ;
        RECT 259.200 732.000 261.000 740.400 ;
        RECT 257.700 730.800 261.000 732.000 ;
        RECT 265.800 731.400 267.600 741.000 ;
        RECT 278.700 737.400 280.500 741.000 ;
        RECT 281.700 735.600 283.500 740.400 ;
        RECT 278.400 734.400 283.500 735.600 ;
        RECT 286.200 734.400 288.000 741.000 ;
        RECT 296.400 735.300 298.200 740.400 ;
        RECT 299.400 736.200 301.200 741.000 ;
        RECT 302.400 735.300 304.200 740.400 ;
        RECT 257.700 727.200 258.600 730.800 ;
        RECT 260.100 727.200 261.900 729.000 ;
        RECT 266.100 727.200 267.900 729.000 ;
        RECT 278.400 727.200 279.300 734.400 ;
        RECT 296.400 733.950 304.200 735.300 ;
        RECT 305.400 734.400 307.200 740.400 ;
        RECT 317.400 737.400 319.200 741.000 ;
        RECT 320.400 737.400 322.200 740.400 ;
        RECT 305.400 732.300 306.600 734.400 ;
        RECT 302.850 731.250 306.600 732.300 ;
        RECT 281.100 727.200 282.900 729.000 ;
        RECT 287.100 727.200 288.900 729.000 ;
        RECT 178.950 724.950 181.200 727.050 ;
        RECT 190.950 725.100 193.050 727.200 ;
        RECT 193.950 725.100 196.050 727.200 ;
        RECT 196.950 725.100 199.050 727.200 ;
        RECT 199.950 725.100 202.050 727.200 ;
        RECT 214.950 725.100 217.050 727.200 ;
        RECT 217.950 725.100 220.050 727.200 ;
        RECT 220.950 725.100 223.050 727.200 ;
        RECT 223.950 725.100 226.050 727.200 ;
        RECT 232.950 725.100 235.050 727.200 ;
        RECT 235.950 725.100 238.050 727.200 ;
        RECT 238.950 725.100 241.050 727.200 ;
        RECT 241.950 725.100 244.050 727.200 ;
        RECT 247.950 726.450 252.000 727.050 ;
        RECT 177.150 719.400 179.100 720.300 ;
        RECT 173.400 718.500 179.100 719.400 ;
        RECT 173.400 711.600 174.600 718.500 ;
        RECT 180.000 717.600 181.200 724.950 ;
        RECT 194.100 723.300 195.900 725.100 ;
        RECT 200.700 717.600 201.600 725.100 ;
        RECT 155.400 705.000 157.200 711.600 ;
        RECT 158.400 705.600 160.200 711.600 ;
        RECT 161.400 705.000 163.200 711.600 ;
        RECT 173.400 705.600 175.200 711.600 ;
        RECT 176.400 705.000 178.200 711.600 ;
        RECT 179.400 705.600 181.200 717.600 ;
        RECT 191.400 716.700 199.200 717.600 ;
        RECT 191.400 705.600 193.200 716.700 ;
        RECT 194.400 705.000 196.200 715.800 ;
        RECT 197.400 705.600 199.200 716.700 ;
        RECT 200.400 705.600 202.200 717.600 ;
        RECT 215.700 712.800 216.600 725.100 ;
        RECT 221.100 723.300 222.900 725.100 ;
        RECT 236.100 723.300 237.900 725.100 ;
        RECT 217.950 720.450 220.050 721.050 ;
        RECT 232.950 720.450 235.050 721.050 ;
        RECT 217.950 719.550 235.050 720.450 ;
        RECT 217.950 718.950 220.050 719.550 ;
        RECT 232.950 718.950 235.050 719.550 ;
        RECT 242.700 717.600 243.600 725.100 ;
        RECT 247.950 724.950 252.450 726.450 ;
        RECT 256.950 725.100 259.050 727.200 ;
        RECT 259.950 725.100 262.050 727.200 ;
        RECT 262.950 725.100 265.050 727.200 ;
        RECT 265.950 725.100 268.050 727.200 ;
        RECT 277.950 725.100 280.050 727.200 ;
        RECT 280.950 725.100 283.050 727.200 ;
        RECT 283.950 725.100 286.050 727.200 ;
        RECT 286.950 725.100 289.050 727.200 ;
        RECT 299.100 727.050 300.900 728.850 ;
        RECT 302.850 727.050 304.050 731.250 ;
        RECT 305.100 727.050 306.900 728.850 ;
        RECT 320.400 727.050 321.600 737.400 ;
        RECT 333.000 734.400 334.800 741.000 ;
        RECT 337.500 735.600 339.300 740.400 ;
        RECT 340.500 737.400 342.300 741.000 ;
        RECT 337.500 734.400 342.600 735.600 ;
        RECT 355.800 734.400 357.600 740.400 ;
        RECT 332.100 727.200 333.900 729.000 ;
        RECT 338.100 727.200 339.900 729.000 ;
        RECT 341.700 727.200 342.600 734.400 ;
        RECT 356.400 732.300 357.600 734.400 ;
        RECT 358.800 735.300 360.600 740.400 ;
        RECT 361.800 736.200 363.600 741.000 ;
        RECT 364.800 735.300 366.600 740.400 ;
        RECT 358.800 733.950 366.600 735.300 ;
        RECT 376.800 734.400 378.600 740.400 ;
        RECT 377.400 732.300 378.600 734.400 ;
        RECT 379.800 735.300 381.600 740.400 ;
        RECT 382.800 736.200 384.600 741.000 ;
        RECT 385.800 735.300 387.600 740.400 ;
        RECT 379.800 733.950 387.600 735.300 ;
        RECT 395.400 735.300 397.200 740.400 ;
        RECT 398.400 736.200 400.200 741.000 ;
        RECT 401.400 735.300 403.200 740.400 ;
        RECT 395.400 733.950 403.200 735.300 ;
        RECT 404.400 734.400 406.200 740.400 ;
        RECT 404.400 732.300 405.600 734.400 ;
        RECT 356.400 731.250 360.150 732.300 ;
        RECT 377.400 731.250 381.150 732.300 ;
        RECT 251.550 724.050 252.450 724.950 ;
        RECT 251.550 722.550 256.050 724.050 ;
        RECT 252.000 721.950 256.050 722.550 ;
        RECT 233.400 716.700 241.200 717.600 ;
        RECT 215.700 711.900 222.300 712.800 ;
        RECT 215.700 711.600 216.600 711.900 ;
        RECT 214.800 705.600 216.600 711.600 ;
        RECT 220.800 711.600 222.300 711.900 ;
        RECT 217.800 705.000 219.600 711.000 ;
        RECT 220.800 705.600 222.600 711.600 ;
        RECT 223.800 705.000 225.600 711.600 ;
        RECT 233.400 705.600 235.200 716.700 ;
        RECT 236.400 705.000 238.200 715.800 ;
        RECT 239.400 705.600 241.200 716.700 ;
        RECT 242.400 705.600 244.200 717.600 ;
        RECT 257.700 712.800 258.600 725.100 ;
        RECT 263.100 723.300 264.900 725.100 ;
        RECT 278.400 717.600 279.300 725.100 ;
        RECT 284.100 723.300 285.900 725.100 ;
        RECT 295.950 724.950 298.050 727.050 ;
        RECT 298.950 724.950 301.050 727.050 ;
        RECT 301.950 724.950 304.050 727.050 ;
        RECT 304.950 724.950 307.050 727.050 ;
        RECT 316.950 724.950 319.050 727.050 ;
        RECT 319.950 724.950 322.050 727.050 ;
        RECT 331.950 725.100 334.050 727.200 ;
        RECT 334.950 725.100 337.050 727.200 ;
        RECT 337.950 725.100 340.050 727.200 ;
        RECT 340.950 725.100 343.050 727.200 ;
        RECT 356.100 727.050 357.900 728.850 ;
        RECT 358.950 727.050 360.150 731.250 ;
        RECT 362.100 727.050 363.900 728.850 ;
        RECT 377.100 727.050 378.900 728.850 ;
        RECT 379.950 727.050 381.150 731.250 ;
        RECT 401.850 731.250 405.600 732.300 ;
        RECT 421.200 732.000 423.000 740.400 ;
        RECT 383.100 727.050 384.900 728.850 ;
        RECT 398.100 727.050 399.900 728.850 ;
        RECT 401.850 727.050 403.050 731.250 ;
        RECT 419.700 730.800 423.000 732.000 ;
        RECT 427.800 731.400 429.600 741.000 ;
        RECT 438.000 734.400 439.800 741.000 ;
        RECT 442.500 735.600 444.300 740.400 ;
        RECT 445.500 737.400 447.300 741.000 ;
        RECT 462.300 736.200 464.100 740.400 ;
        RECT 442.500 734.400 447.600 735.600 ;
        RECT 406.950 729.450 411.000 730.050 ;
        RECT 404.100 727.050 405.900 728.850 ;
        RECT 406.950 727.950 411.450 729.450 ;
        RECT 296.100 723.150 297.900 724.950 ;
        RECT 289.950 720.450 292.050 721.050 ;
        RECT 295.950 720.450 298.050 721.050 ;
        RECT 289.950 719.550 298.050 720.450 ;
        RECT 289.950 718.950 292.050 719.550 ;
        RECT 295.950 718.950 298.050 719.550 ;
        RECT 257.700 711.900 264.300 712.800 ;
        RECT 257.700 711.600 258.600 711.900 ;
        RECT 256.800 705.600 258.600 711.600 ;
        RECT 262.800 711.600 264.300 711.900 ;
        RECT 259.800 705.000 261.600 711.000 ;
        RECT 262.800 705.600 264.600 711.600 ;
        RECT 265.800 705.000 267.600 711.600 ;
        RECT 277.800 705.600 279.600 717.600 ;
        RECT 280.800 716.700 288.600 717.600 ;
        RECT 280.800 705.600 282.600 716.700 ;
        RECT 283.800 705.000 285.600 715.800 ;
        RECT 286.800 705.600 288.600 716.700 ;
        RECT 296.700 705.000 298.500 717.600 ;
        RECT 301.950 711.600 303.150 724.950 ;
        RECT 317.100 723.150 318.900 724.950 ;
        RECT 320.400 711.600 321.600 724.950 ;
        RECT 335.100 723.300 336.900 725.100 ;
        RECT 341.700 717.600 342.600 725.100 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 358.950 724.950 361.050 727.050 ;
        RECT 361.950 724.950 364.050 727.050 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 379.950 724.950 382.050 727.050 ;
        RECT 382.950 724.950 385.050 727.050 ;
        RECT 385.950 724.950 388.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 400.950 724.950 403.050 727.050 ;
        RECT 403.950 724.950 406.050 727.050 ;
        RECT 332.400 716.700 340.200 717.600 ;
        RECT 301.800 705.600 303.600 711.600 ;
        RECT 304.800 705.000 306.600 711.600 ;
        RECT 317.400 705.000 319.200 711.600 ;
        RECT 320.400 705.600 322.200 711.600 ;
        RECT 332.400 705.600 334.200 716.700 ;
        RECT 335.400 705.000 337.200 715.800 ;
        RECT 338.400 705.600 340.200 716.700 ;
        RECT 341.400 705.600 343.200 717.600 ;
        RECT 359.850 711.600 361.050 724.950 ;
        RECT 365.100 723.150 366.900 724.950 ;
        RECT 364.950 720.450 369.000 721.050 ;
        RECT 364.950 718.950 369.450 720.450 ;
        RECT 356.400 705.000 358.200 711.600 ;
        RECT 359.400 705.600 361.200 711.600 ;
        RECT 364.500 705.000 366.300 717.600 ;
        RECT 368.550 717.450 369.450 718.950 ;
        RECT 376.950 717.450 379.050 718.050 ;
        RECT 368.550 716.550 379.050 717.450 ;
        RECT 376.950 715.950 379.050 716.550 ;
        RECT 380.850 711.600 382.050 724.950 ;
        RECT 386.100 723.150 387.900 724.950 ;
        RECT 395.100 723.150 396.900 724.950 ;
        RECT 377.400 705.000 379.200 711.600 ;
        RECT 380.400 705.600 382.200 711.600 ;
        RECT 385.500 705.000 387.300 717.600 ;
        RECT 395.700 705.000 397.500 717.600 ;
        RECT 400.950 711.600 402.150 724.950 ;
        RECT 410.550 723.450 411.450 727.950 ;
        RECT 419.700 727.200 420.600 730.800 ;
        RECT 422.100 727.200 423.900 729.000 ;
        RECT 428.100 727.200 429.900 729.000 ;
        RECT 437.100 727.200 438.900 729.000 ;
        RECT 443.100 727.200 444.900 729.000 ;
        RECT 446.700 727.200 447.600 734.400 ;
        RECT 461.400 734.400 464.100 736.200 ;
        RECT 465.300 734.400 467.100 741.000 ;
        RECT 461.400 727.200 462.300 734.400 ;
        RECT 464.100 732.600 465.900 733.500 ;
        RECT 469.800 732.600 471.600 740.400 ;
        RECT 464.100 731.700 471.600 732.600 ;
        RECT 482.400 733.200 484.200 740.400 ;
        RECT 487.500 734.400 489.300 741.000 ;
        RECT 497.400 737.400 499.200 740.400 ;
        RECT 500.400 737.400 502.200 741.000 ;
        RECT 497.400 733.500 498.600 737.400 ;
        RECT 503.400 734.400 505.200 740.400 ;
        RECT 517.800 737.400 519.600 740.400 ;
        RECT 520.800 737.400 522.600 741.000 ;
        RECT 482.400 732.300 486.600 733.200 ;
        RECT 497.400 732.600 503.100 733.500 ;
        RECT 418.950 725.100 421.050 727.200 ;
        RECT 421.950 725.100 424.050 727.200 ;
        RECT 424.950 725.100 427.050 727.200 ;
        RECT 427.950 725.100 430.050 727.200 ;
        RECT 436.950 725.100 439.050 727.200 ;
        RECT 439.950 725.100 442.050 727.200 ;
        RECT 442.950 725.100 445.050 727.200 ;
        RECT 445.950 725.100 448.050 727.200 ;
        RECT 460.950 725.100 463.050 727.200 ;
        RECT 463.950 725.100 466.050 727.200 ;
        RECT 415.950 723.450 418.050 724.050 ;
        RECT 410.550 722.550 418.050 723.450 ;
        RECT 415.950 721.950 418.050 722.550 ;
        RECT 419.700 712.800 420.600 725.100 ;
        RECT 425.100 723.300 426.900 725.100 ;
        RECT 440.100 723.300 441.900 725.100 ;
        RECT 446.700 717.600 447.600 725.100 ;
        RECT 461.400 717.600 462.300 725.100 ;
        RECT 464.100 723.300 465.900 725.100 ;
        RECT 437.400 716.700 445.200 717.600 ;
        RECT 419.700 711.900 426.300 712.800 ;
        RECT 419.700 711.600 420.600 711.900 ;
        RECT 400.800 705.600 402.600 711.600 ;
        RECT 403.800 705.000 405.600 711.600 ;
        RECT 418.800 705.600 420.600 711.600 ;
        RECT 424.800 711.600 426.300 711.900 ;
        RECT 421.800 705.000 423.600 711.000 ;
        RECT 424.800 705.600 426.600 711.600 ;
        RECT 427.800 705.000 429.600 711.600 ;
        RECT 437.400 705.600 439.200 716.700 ;
        RECT 440.400 705.000 442.200 715.800 ;
        RECT 443.400 705.600 445.200 716.700 ;
        RECT 446.400 705.600 448.200 717.600 ;
        RECT 460.800 705.600 462.600 717.600 ;
        RECT 467.700 711.600 468.600 731.700 ;
        RECT 470.100 727.200 471.900 729.000 ;
        RECT 482.100 727.200 483.900 729.000 ;
        RECT 485.400 727.200 486.600 732.300 ;
        RECT 501.150 731.700 503.100 732.600 ;
        RECT 488.100 727.200 489.900 729.000 ;
        RECT 469.950 725.100 472.050 727.200 ;
        RECT 481.950 725.100 484.050 727.200 ;
        RECT 484.950 725.100 487.050 727.200 ;
        RECT 487.950 725.100 490.050 727.200 ;
        RECT 469.950 723.450 472.050 724.050 ;
        RECT 481.950 723.450 484.050 724.050 ;
        RECT 469.950 722.550 484.050 723.450 ;
        RECT 469.950 721.950 472.050 722.550 ;
        RECT 481.950 721.950 484.050 722.550 ;
        RECT 485.400 711.600 486.600 725.100 ;
        RECT 496.950 724.950 499.050 727.050 ;
        RECT 497.100 723.150 498.900 724.950 ;
        RECT 501.150 720.300 502.050 731.700 ;
        RECT 504.000 727.050 505.200 734.400 ;
        RECT 508.950 729.450 511.050 730.050 ;
        RECT 514.950 729.450 517.050 730.050 ;
        RECT 508.950 728.550 517.050 729.450 ;
        RECT 508.950 727.950 511.050 728.550 ;
        RECT 514.950 727.950 517.050 728.550 ;
        RECT 518.400 727.050 519.600 737.400 ;
        RECT 530.400 735.300 532.200 740.400 ;
        RECT 533.400 736.200 535.200 741.000 ;
        RECT 536.400 735.300 538.200 740.400 ;
        RECT 530.400 733.950 538.200 735.300 ;
        RECT 539.400 734.400 541.200 740.400 ;
        RECT 551.400 735.300 553.200 740.400 ;
        RECT 554.400 736.200 556.200 741.000 ;
        RECT 557.400 735.300 559.200 740.400 ;
        RECT 539.400 732.300 540.600 734.400 ;
        RECT 551.400 733.950 559.200 735.300 ;
        RECT 560.400 734.400 562.200 740.400 ;
        RECT 573.000 734.400 574.800 741.000 ;
        RECT 577.500 735.600 579.300 740.400 ;
        RECT 580.500 737.400 582.300 741.000 ;
        RECT 577.500 734.400 582.600 735.600 ;
        RECT 560.400 732.300 561.600 734.400 ;
        RECT 536.850 731.250 540.600 732.300 ;
        RECT 557.850 731.250 561.600 732.300 ;
        RECT 533.100 727.050 534.900 728.850 ;
        RECT 536.850 727.050 538.050 731.250 ;
        RECT 539.100 727.050 540.900 728.850 ;
        RECT 554.100 727.050 555.900 728.850 ;
        RECT 557.850 727.050 559.050 731.250 ;
        RECT 562.950 729.450 567.000 730.050 ;
        RECT 560.100 727.050 561.900 728.850 ;
        RECT 562.950 727.950 567.450 729.450 ;
        RECT 502.950 724.950 505.200 727.050 ;
        RECT 517.950 724.950 520.050 727.050 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 556.950 724.950 559.050 727.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 501.150 719.400 503.100 720.300 ;
        RECT 497.400 718.500 503.100 719.400 ;
        RECT 497.400 711.600 498.600 718.500 ;
        RECT 504.000 717.600 505.200 724.950 ;
        RECT 463.800 705.000 465.600 711.600 ;
        RECT 466.800 705.600 468.600 711.600 ;
        RECT 469.800 705.000 471.600 711.600 ;
        RECT 481.800 705.000 483.600 711.600 ;
        RECT 484.800 705.600 486.600 711.600 ;
        RECT 487.800 705.000 489.600 711.600 ;
        RECT 497.400 705.600 499.200 711.600 ;
        RECT 500.400 705.000 502.200 711.600 ;
        RECT 503.400 705.600 505.200 717.600 ;
        RECT 518.400 711.600 519.600 724.950 ;
        RECT 521.100 723.150 522.900 724.950 ;
        RECT 530.100 723.150 531.900 724.950 ;
        RECT 517.800 705.600 519.600 711.600 ;
        RECT 520.800 705.000 522.600 711.600 ;
        RECT 530.700 705.000 532.500 717.600 ;
        RECT 535.950 711.600 537.150 724.950 ;
        RECT 551.100 723.150 552.900 724.950 ;
        RECT 535.800 705.600 537.600 711.600 ;
        RECT 538.800 705.000 540.600 711.600 ;
        RECT 551.700 705.000 553.500 717.600 ;
        RECT 556.950 711.600 558.150 724.950 ;
        RECT 566.550 724.050 567.450 727.950 ;
        RECT 572.100 727.200 573.900 729.000 ;
        RECT 578.100 727.200 579.900 729.000 ;
        RECT 581.700 727.200 582.600 734.400 ;
        RECT 596.400 733.200 598.200 740.400 ;
        RECT 601.500 734.400 603.300 741.000 ;
        RECT 611.400 735.300 613.200 740.400 ;
        RECT 614.400 736.200 616.200 741.000 ;
        RECT 617.400 735.300 619.200 740.400 ;
        RECT 611.400 733.950 619.200 735.300 ;
        RECT 620.400 734.400 622.200 740.400 ;
        RECT 632.400 735.300 634.200 740.400 ;
        RECT 635.400 736.200 637.200 741.000 ;
        RECT 680.400 740.400 681.600 741.000 ;
        RECT 638.400 735.300 640.200 740.400 ;
        RECT 596.400 732.300 600.600 733.200 ;
        RECT 620.400 732.300 621.600 734.400 ;
        RECT 632.400 733.950 640.200 735.300 ;
        RECT 641.400 734.400 643.200 740.400 ;
        RECT 655.800 734.400 657.600 740.400 ;
        RECT 663.300 734.400 665.100 740.400 ;
        RECT 670.800 734.400 672.600 740.400 ;
        RECT 680.400 737.400 682.200 740.400 ;
        RECT 683.400 737.400 685.200 740.400 ;
        RECT 686.400 737.400 688.200 741.000 ;
        RECT 641.400 732.300 642.600 734.400 ;
        RECT 655.800 733.500 660.600 734.400 ;
        RECT 658.500 732.300 660.600 733.500 ;
        RECT 663.600 732.900 664.800 734.400 ;
        RECT 596.100 727.200 597.900 729.000 ;
        RECT 599.400 727.200 600.600 732.300 ;
        RECT 617.850 731.250 621.600 732.300 ;
        RECT 638.850 731.250 642.600 732.300 ;
        RECT 602.100 727.200 603.900 729.000 ;
        RECT 571.950 725.100 574.050 727.200 ;
        RECT 574.950 725.100 577.050 727.200 ;
        RECT 577.950 725.100 580.050 727.200 ;
        RECT 580.950 725.100 583.050 727.200 ;
        RECT 595.950 725.100 598.050 727.200 ;
        RECT 598.950 725.100 601.050 727.200 ;
        RECT 601.950 725.100 604.050 727.200 ;
        RECT 614.100 727.050 615.900 728.850 ;
        RECT 617.850 727.050 619.050 731.250 ;
        RECT 620.100 727.050 621.900 728.850 ;
        RECT 635.100 727.050 636.900 728.850 ;
        RECT 638.850 727.050 640.050 731.250 ;
        RECT 661.950 730.800 664.800 732.900 ;
        RECT 670.800 732.600 672.000 734.400 ;
        RECT 641.100 727.050 642.900 728.850 ;
        RECT 660.750 727.800 662.850 729.900 ;
        RECT 566.550 722.550 571.050 724.050 ;
        RECT 575.100 723.300 576.900 725.100 ;
        RECT 567.000 721.950 571.050 722.550 ;
        RECT 562.950 720.450 565.050 721.050 ;
        RECT 577.950 720.450 580.050 720.900 ;
        RECT 562.950 719.550 580.050 720.450 ;
        RECT 562.950 718.950 565.050 719.550 ;
        RECT 577.950 718.800 580.050 719.550 ;
        RECT 581.700 717.600 582.600 725.100 ;
        RECT 589.950 723.450 592.050 724.050 ;
        RECT 595.950 723.450 598.050 724.050 ;
        RECT 589.950 722.550 598.050 723.450 ;
        RECT 589.950 721.950 592.050 722.550 ;
        RECT 595.950 721.950 598.050 722.550 ;
        RECT 572.400 716.700 580.200 717.600 ;
        RECT 556.800 705.600 558.600 711.600 ;
        RECT 559.800 705.000 561.600 711.600 ;
        RECT 572.400 705.600 574.200 716.700 ;
        RECT 575.400 705.000 577.200 715.800 ;
        RECT 578.400 705.600 580.200 716.700 ;
        RECT 581.400 705.600 583.200 717.600 ;
        RECT 599.400 711.600 600.600 725.100 ;
        RECT 610.950 724.950 613.050 727.050 ;
        RECT 613.950 724.950 616.050 727.050 ;
        RECT 616.950 724.950 619.050 727.050 ;
        RECT 619.950 724.950 622.050 727.050 ;
        RECT 631.950 724.950 634.050 727.050 ;
        RECT 634.950 724.950 637.050 727.050 ;
        RECT 637.950 724.950 640.050 727.050 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 655.950 725.100 658.050 727.200 ;
        RECT 660.600 726.000 662.400 727.800 ;
        RECT 663.750 725.100 664.800 730.800 ;
        RECT 665.700 731.700 672.000 732.600 ;
        RECT 684.300 733.200 685.200 737.400 ;
        RECT 689.400 734.400 691.200 740.400 ;
        RECT 701.400 735.300 703.200 740.400 ;
        RECT 704.400 736.200 706.200 741.000 ;
        RECT 707.400 735.300 709.200 740.400 ;
        RECT 684.300 732.300 687.600 733.200 ;
        RECT 665.700 729.600 667.800 731.700 ;
        RECT 685.800 731.400 687.600 732.300 ;
        RECT 665.700 727.800 667.500 729.600 ;
        RECT 670.950 727.200 672.750 729.000 ;
        RECT 670.950 726.300 673.050 727.200 ;
        RECT 680.100 727.050 681.900 728.850 ;
        RECT 611.100 723.150 612.900 724.950 ;
        RECT 595.800 705.000 597.600 711.600 ;
        RECT 598.800 705.600 600.600 711.600 ;
        RECT 601.800 705.000 603.600 711.600 ;
        RECT 611.700 705.000 613.500 717.600 ;
        RECT 616.950 711.600 618.150 724.950 ;
        RECT 632.100 723.150 633.900 724.950 ;
        RECT 616.800 705.600 618.600 711.600 ;
        RECT 619.800 705.000 621.600 711.600 ;
        RECT 632.700 705.000 634.500 717.600 ;
        RECT 637.950 711.600 639.150 724.950 ;
        RECT 649.950 723.450 652.050 724.050 ;
        RECT 656.100 723.450 657.900 725.100 ;
        RECT 662.400 724.200 664.800 725.100 ;
        RECT 665.700 725.100 673.050 726.300 ;
        RECT 665.700 724.500 667.500 725.100 ;
        RECT 679.950 724.950 682.050 727.050 ;
        RECT 682.950 724.950 685.050 727.050 ;
        RECT 649.950 723.300 657.900 723.450 ;
        RECT 649.950 722.550 657.450 723.300 ;
        RECT 649.950 721.950 652.050 722.550 ;
        RECT 661.950 722.100 664.050 724.200 ;
        RECT 640.950 720.450 643.050 720.750 ;
        RECT 652.950 720.450 655.050 721.050 ;
        RECT 640.950 719.550 655.050 720.450 ;
        RECT 640.950 718.650 643.050 719.550 ;
        RECT 652.950 718.950 655.050 719.550 ;
        RECT 663.000 720.000 663.900 722.100 ;
        RECT 664.950 721.500 668.700 723.300 ;
        RECT 683.100 723.150 684.900 724.950 ;
        RECT 664.950 721.200 667.050 721.500 ;
        RECT 686.700 720.900 687.600 731.400 ;
        RECT 690.000 727.050 691.050 734.400 ;
        RECT 701.400 733.950 709.200 735.300 ;
        RECT 710.400 734.400 712.200 740.400 ;
        RECT 725.700 737.400 727.500 741.000 ;
        RECT 728.700 735.600 730.500 740.400 ;
        RECT 725.400 734.400 730.500 735.600 ;
        RECT 733.200 734.400 735.000 741.000 ;
        RECT 743.400 735.300 745.200 740.400 ;
        RECT 746.400 736.200 748.200 741.000 ;
        RECT 749.400 735.300 751.200 740.400 ;
        RECT 710.400 732.300 711.600 734.400 ;
        RECT 707.850 731.250 711.600 732.300 ;
        RECT 704.100 727.050 705.900 728.850 ;
        RECT 707.850 727.050 709.050 731.250 ;
        RECT 710.100 727.050 711.900 728.850 ;
        RECT 725.400 727.200 726.300 734.400 ;
        RECT 743.400 733.950 751.200 735.300 ;
        RECT 752.400 734.400 754.200 740.400 ;
        RECT 765.000 734.400 766.800 741.000 ;
        RECT 769.500 735.600 771.300 740.400 ;
        RECT 772.500 737.400 774.300 741.000 ;
        RECT 769.500 734.400 774.600 735.600 ;
        RECT 752.400 732.300 753.600 734.400 ;
        RECT 749.850 731.250 753.600 732.300 ;
        RECT 728.100 727.200 729.900 729.000 ;
        RECT 734.100 727.200 735.900 729.000 ;
        RECT 685.800 720.300 687.600 720.900 ;
        RECT 663.000 719.100 664.500 720.000 ;
        RECT 658.500 717.600 660.600 718.500 ;
        RECT 655.800 716.400 660.600 717.600 ;
        RECT 663.300 717.600 664.500 719.100 ;
        RECT 668.100 717.600 670.200 719.700 ;
        RECT 680.400 719.100 687.600 720.300 ;
        RECT 688.950 724.950 691.050 727.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 706.950 724.950 709.050 727.050 ;
        RECT 709.950 724.950 712.050 727.050 ;
        RECT 724.950 725.100 727.050 727.200 ;
        RECT 727.950 725.100 730.050 727.200 ;
        RECT 730.950 725.100 733.050 727.200 ;
        RECT 733.950 725.100 736.050 727.200 ;
        RECT 746.100 727.050 747.900 728.850 ;
        RECT 749.850 727.050 751.050 731.250 ;
        RECT 752.100 727.050 753.900 728.850 ;
        RECT 764.100 727.200 765.900 729.000 ;
        RECT 770.100 727.200 771.900 729.000 ;
        RECT 773.700 727.200 774.600 734.400 ;
        RECT 785.400 731.400 787.200 741.000 ;
        RECT 792.000 732.000 793.800 740.400 ;
        RECT 808.800 734.400 810.600 740.400 ;
        RECT 809.400 732.300 810.600 734.400 ;
        RECT 811.800 735.300 813.600 740.400 ;
        RECT 814.800 736.200 816.600 741.000 ;
        RECT 817.800 735.300 819.600 740.400 ;
        RECT 830.700 737.400 832.500 741.000 ;
        RECT 833.700 735.600 835.500 740.400 ;
        RECT 811.800 733.950 819.600 735.300 ;
        RECT 830.400 734.400 835.500 735.600 ;
        RECT 838.200 734.400 840.000 741.000 ;
        RECT 848.400 735.300 850.200 740.400 ;
        RECT 851.400 736.200 853.200 741.000 ;
        RECT 854.400 735.300 856.200 740.400 ;
        RECT 792.000 730.800 795.300 732.000 ;
        RECT 809.400 731.250 813.150 732.300 ;
        RECT 785.100 727.200 786.900 729.000 ;
        RECT 791.100 727.200 792.900 729.000 ;
        RECT 794.400 727.200 795.300 730.800 ;
        RECT 680.400 717.600 681.600 719.100 ;
        RECT 688.950 717.600 690.300 724.950 ;
        RECT 701.100 723.150 702.900 724.950 ;
        RECT 637.800 705.600 639.600 711.600 ;
        RECT 640.800 705.000 642.600 711.600 ;
        RECT 655.800 705.600 657.600 716.400 ;
        RECT 663.300 705.600 665.100 717.600 ;
        RECT 668.100 716.700 672.600 717.600 ;
        RECT 670.800 705.600 672.600 716.700 ;
        RECT 680.400 705.600 682.200 717.600 ;
        RECT 684.900 705.000 686.700 717.600 ;
        RECT 687.900 716.100 690.300 717.600 ;
        RECT 687.900 705.600 689.700 716.100 ;
        RECT 701.700 705.000 703.500 717.600 ;
        RECT 706.950 711.600 708.150 724.950 ;
        RECT 725.400 717.600 726.300 725.100 ;
        RECT 731.100 723.300 732.900 725.100 ;
        RECT 742.950 724.950 745.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 763.950 725.100 766.050 727.200 ;
        RECT 766.950 725.100 769.050 727.200 ;
        RECT 769.950 725.100 772.050 727.200 ;
        RECT 772.950 725.100 775.050 727.200 ;
        RECT 784.950 725.100 787.050 727.200 ;
        RECT 787.950 725.100 790.050 727.200 ;
        RECT 790.950 725.100 793.050 727.200 ;
        RECT 793.950 725.100 796.050 727.200 ;
        RECT 809.100 727.050 810.900 728.850 ;
        RECT 811.950 727.050 813.150 731.250 ;
        RECT 815.100 727.050 816.900 728.850 ;
        RECT 830.400 727.200 831.300 734.400 ;
        RECT 848.400 733.950 856.200 735.300 ;
        RECT 857.400 734.400 859.200 740.400 ;
        RECT 857.400 732.300 858.600 734.400 ;
        RECT 854.850 731.250 858.600 732.300 ;
        RECT 833.100 727.200 834.900 729.000 ;
        RECT 839.100 727.200 840.900 729.000 ;
        RECT 743.100 723.150 744.900 724.950 ;
        RECT 706.800 705.600 708.600 711.600 ;
        RECT 709.800 705.000 711.600 711.600 ;
        RECT 724.800 705.600 726.600 717.600 ;
        RECT 727.800 716.700 735.600 717.600 ;
        RECT 727.800 705.600 729.600 716.700 ;
        RECT 730.800 705.000 732.600 715.800 ;
        RECT 733.800 705.600 735.600 716.700 ;
        RECT 743.700 705.000 745.500 717.600 ;
        RECT 748.950 711.600 750.150 724.950 ;
        RECT 767.100 723.300 768.900 725.100 ;
        RECT 773.700 717.600 774.600 725.100 ;
        RECT 778.950 723.450 781.050 724.050 ;
        RECT 784.950 723.450 787.050 724.050 ;
        RECT 778.950 722.550 787.050 723.450 ;
        RECT 788.100 723.300 789.900 725.100 ;
        RECT 778.950 721.950 781.050 722.550 ;
        RECT 784.950 721.950 787.050 722.550 ;
        RECT 764.400 716.700 772.200 717.600 ;
        RECT 748.800 705.600 750.600 711.600 ;
        RECT 751.800 705.000 753.600 711.600 ;
        RECT 764.400 705.600 766.200 716.700 ;
        RECT 767.400 705.000 769.200 715.800 ;
        RECT 770.400 705.600 772.200 716.700 ;
        RECT 773.400 705.600 775.200 717.600 ;
        RECT 794.400 712.800 795.300 725.100 ;
        RECT 808.950 724.950 811.050 727.050 ;
        RECT 811.950 724.950 814.050 727.050 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 829.950 725.100 832.050 727.200 ;
        RECT 832.950 725.100 835.050 727.200 ;
        RECT 835.950 725.100 838.050 727.200 ;
        RECT 838.950 725.100 841.050 727.200 ;
        RECT 851.100 727.050 852.900 728.850 ;
        RECT 854.850 727.050 856.050 731.250 ;
        RECT 857.100 727.050 858.900 728.850 ;
        RECT 788.700 711.900 795.300 712.800 ;
        RECT 788.700 711.600 790.200 711.900 ;
        RECT 785.400 705.000 787.200 711.600 ;
        RECT 788.400 705.600 790.200 711.600 ;
        RECT 794.400 711.600 795.300 711.900 ;
        RECT 812.850 711.600 814.050 724.950 ;
        RECT 818.100 723.150 819.900 724.950 ;
        RECT 830.400 717.600 831.300 725.100 ;
        RECT 836.100 723.300 837.900 725.100 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 853.950 724.950 856.050 727.050 ;
        RECT 856.950 724.950 859.050 727.050 ;
        RECT 848.100 723.150 849.900 724.950 ;
        RECT 832.950 720.450 835.050 721.050 ;
        RECT 844.950 720.450 847.050 721.050 ;
        RECT 832.950 719.550 847.050 720.450 ;
        RECT 832.950 718.950 835.050 719.550 ;
        RECT 844.950 718.950 847.050 719.550 ;
        RECT 791.400 705.000 793.200 711.000 ;
        RECT 794.400 705.600 796.200 711.600 ;
        RECT 809.400 705.000 811.200 711.600 ;
        RECT 812.400 705.600 814.200 711.600 ;
        RECT 817.500 705.000 819.300 717.600 ;
        RECT 829.800 705.600 831.600 717.600 ;
        RECT 832.800 716.700 840.600 717.600 ;
        RECT 832.800 705.600 834.600 716.700 ;
        RECT 835.800 705.000 837.600 715.800 ;
        RECT 838.800 705.600 840.600 716.700 ;
        RECT 848.700 705.000 850.500 717.600 ;
        RECT 853.950 711.600 855.150 724.950 ;
        RECT 853.800 705.600 855.600 711.600 ;
        RECT 856.800 705.000 858.600 711.600 ;
        RECT 10.800 695.400 12.600 701.400 ;
        RECT 13.800 695.400 15.600 702.000 ;
        RECT 11.400 682.050 12.600 695.400 ;
        RECT 27.300 689.400 29.100 702.000 ;
        RECT 31.800 689.400 35.100 701.400 ;
        RECT 37.800 689.400 39.600 702.000 ;
        RECT 47.400 689.400 49.200 702.000 ;
        RECT 52.500 690.600 54.300 701.400 ;
        RECT 65.400 695.400 67.200 702.000 ;
        RECT 68.400 695.400 70.200 701.400 ;
        RECT 50.700 689.400 54.300 690.600 ;
        RECT 14.100 682.050 15.900 683.850 ;
        RECT 10.950 679.950 13.050 682.050 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 26.100 681.900 27.900 683.700 ;
        RECT 32.700 681.900 33.900 689.400 ;
        RECT 38.100 681.900 39.900 683.700 ;
        RECT 47.100 682.050 48.900 683.850 ;
        RECT 50.700 682.050 51.600 689.400 ;
        RECT 53.100 682.050 54.900 683.850 ;
        RECT 65.100 682.050 66.900 683.850 ;
        RECT 68.400 682.050 69.600 695.400 ;
        RECT 80.400 690.300 82.200 701.400 ;
        RECT 83.400 691.200 85.200 702.000 ;
        RECT 86.400 690.300 88.200 701.400 ;
        RECT 80.400 689.400 88.200 690.300 ;
        RECT 89.400 689.400 91.200 701.400 ;
        RECT 103.800 695.400 105.600 702.000 ;
        RECT 106.800 695.400 108.600 701.400 ;
        RECT 109.800 695.400 111.600 702.000 ;
        RECT 11.400 669.600 12.600 679.950 ;
        RECT 25.950 679.800 28.050 681.900 ;
        RECT 28.950 679.800 31.050 681.900 ;
        RECT 31.950 679.800 34.050 681.900 ;
        RECT 34.950 679.800 37.050 681.900 ;
        RECT 37.950 679.800 40.050 681.900 ;
        RECT 46.950 679.950 49.050 682.050 ;
        RECT 49.950 679.950 52.050 682.050 ;
        RECT 52.950 679.950 55.050 682.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 67.950 679.950 70.050 682.050 ;
        RECT 83.100 681.900 84.900 683.700 ;
        RECT 89.700 681.900 90.600 689.400 ;
        RECT 94.950 687.450 97.050 688.050 ;
        RECT 103.950 687.450 106.050 688.050 ;
        RECT 94.950 686.550 106.050 687.450 ;
        RECT 94.950 685.950 97.050 686.550 ;
        RECT 103.950 685.950 106.050 686.550 ;
        RECT 91.950 684.450 96.000 685.050 ;
        RECT 91.950 682.950 96.450 684.450 ;
        RECT 29.100 678.000 30.900 679.800 ;
        RECT 33.000 677.400 34.050 679.800 ;
        RECT 35.100 678.000 36.900 679.800 ;
        RECT 32.700 675.300 33.900 677.400 ;
        RECT 29.400 674.100 33.900 675.300 ;
        RECT 29.400 672.600 30.300 674.100 ;
        RECT 10.800 666.600 12.600 669.600 ;
        RECT 13.800 666.000 15.600 669.600 ;
        RECT 25.800 667.500 27.600 672.600 ;
        RECT 28.800 668.400 30.600 672.600 ;
        RECT 31.800 672.000 39.600 672.900 ;
        RECT 31.800 667.500 33.600 672.000 ;
        RECT 25.800 666.600 33.600 667.500 ;
        RECT 34.800 666.000 36.600 671.100 ;
        RECT 37.800 666.600 39.600 672.000 ;
        RECT 50.700 669.600 51.600 679.950 ;
        RECT 52.950 675.450 55.050 676.050 ;
        RECT 58.950 675.450 61.050 676.050 ;
        RECT 52.950 674.550 61.050 675.450 ;
        RECT 52.950 673.950 55.050 674.550 ;
        RECT 58.950 673.950 61.050 674.550 ;
        RECT 68.400 669.600 69.600 679.950 ;
        RECT 79.950 679.800 82.050 681.900 ;
        RECT 82.950 679.800 85.050 681.900 ;
        RECT 85.950 679.800 88.050 681.900 ;
        RECT 88.950 679.800 91.050 681.900 ;
        RECT 95.550 681.450 96.450 682.950 ;
        RECT 107.400 681.900 108.600 695.400 ;
        RECT 119.400 690.600 121.200 701.400 ;
        RECT 122.400 691.500 124.200 702.000 ;
        RECT 125.400 700.500 133.200 701.400 ;
        RECT 125.400 690.600 127.200 700.500 ;
        RECT 119.400 689.700 127.200 690.600 ;
        RECT 128.400 688.500 130.200 699.600 ;
        RECT 131.400 689.400 133.200 700.500 ;
        RECT 145.800 689.400 147.600 701.400 ;
        RECT 148.800 695.400 150.600 702.000 ;
        RECT 151.800 695.400 153.600 701.400 ;
        RECT 163.800 695.400 165.600 701.400 ;
        RECT 166.800 696.000 168.600 702.000 ;
        RECT 125.100 687.600 130.200 688.500 ;
        RECT 122.100 681.900 123.900 683.700 ;
        RECT 125.100 681.900 126.000 687.600 ;
        RECT 130.950 684.450 133.050 684.900 ;
        RECT 139.950 684.450 142.050 685.050 ;
        RECT 128.100 681.900 129.900 683.700 ;
        RECT 130.950 683.550 142.050 684.450 ;
        RECT 130.950 682.800 133.050 683.550 ;
        RECT 139.950 682.950 142.050 683.550 ;
        RECT 145.800 682.050 147.000 689.400 ;
        RECT 152.400 688.500 153.600 695.400 ;
        RECT 147.900 687.600 153.600 688.500 ;
        RECT 164.700 695.100 165.600 695.400 ;
        RECT 169.800 695.400 171.600 701.400 ;
        RECT 172.800 695.400 174.600 702.000 ;
        RECT 182.400 695.400 184.200 702.000 ;
        RECT 185.400 695.400 187.200 701.400 ;
        RECT 188.400 696.000 190.200 702.000 ;
        RECT 169.800 695.100 171.300 695.400 ;
        RECT 164.700 694.200 171.300 695.100 ;
        RECT 185.700 695.100 187.200 695.400 ;
        RECT 191.400 695.400 193.200 701.400 ;
        RECT 191.400 695.100 192.300 695.400 ;
        RECT 185.700 694.200 192.300 695.100 ;
        RECT 147.900 686.700 149.850 687.600 ;
        RECT 95.550 680.550 99.450 681.450 ;
        RECT 80.100 678.000 81.900 679.800 ;
        RECT 86.100 678.000 87.900 679.800 ;
        RECT 89.700 672.600 90.600 679.800 ;
        RECT 98.550 679.050 99.450 680.550 ;
        RECT 103.950 679.800 106.050 681.900 ;
        RECT 106.950 679.800 109.050 681.900 ;
        RECT 109.950 679.800 112.050 681.900 ;
        RECT 118.950 679.800 121.050 681.900 ;
        RECT 121.950 679.800 124.050 681.900 ;
        RECT 124.950 679.800 127.050 681.900 ;
        RECT 127.950 679.800 130.050 681.900 ;
        RECT 130.950 679.800 133.050 681.900 ;
        RECT 145.800 679.950 148.050 682.050 ;
        RECT 98.550 677.550 103.050 679.050 ;
        RECT 104.100 678.000 105.900 679.800 ;
        RECT 99.000 676.950 103.050 677.550 ;
        RECT 107.400 674.700 108.600 679.800 ;
        RECT 110.100 678.000 111.900 679.800 ;
        RECT 119.100 678.000 120.900 679.800 ;
        RECT 47.400 666.000 49.200 669.600 ;
        RECT 50.400 666.600 52.200 669.600 ;
        RECT 53.400 666.000 55.200 669.600 ;
        RECT 65.400 666.000 67.200 669.600 ;
        RECT 68.400 666.600 70.200 669.600 ;
        RECT 81.000 666.000 82.800 672.600 ;
        RECT 85.500 671.400 90.600 672.600 ;
        RECT 104.400 673.800 108.600 674.700 ;
        RECT 85.500 666.600 87.300 671.400 ;
        RECT 88.500 666.000 90.300 669.600 ;
        RECT 104.400 666.600 106.200 673.800 ;
        RECT 124.950 672.600 126.000 679.800 ;
        RECT 131.100 678.000 132.900 679.800 ;
        RECT 145.800 672.600 147.000 679.950 ;
        RECT 148.950 675.300 149.850 686.700 ;
        RECT 152.100 682.050 153.900 683.850 ;
        RECT 151.950 679.950 154.050 682.050 ;
        RECT 164.700 681.900 165.600 694.200 ;
        RECT 172.950 684.450 175.050 685.050 ;
        RECT 181.950 684.450 184.050 685.050 ;
        RECT 170.100 681.900 171.900 683.700 ;
        RECT 172.950 683.550 184.050 684.450 ;
        RECT 172.950 682.950 175.050 683.550 ;
        RECT 181.950 682.950 184.050 683.550 ;
        RECT 185.100 681.900 186.900 683.700 ;
        RECT 191.400 681.900 192.300 694.200 ;
        RECT 203.700 689.400 205.500 702.000 ;
        RECT 208.800 695.400 210.600 701.400 ;
        RECT 211.800 695.400 213.600 702.000 ;
        RECT 227.400 695.400 229.200 702.000 ;
        RECT 230.400 695.400 232.200 701.400 ;
        RECT 203.100 682.050 204.900 683.850 ;
        RECT 208.950 682.050 210.150 695.400 ;
        RECT 230.850 682.050 232.050 695.400 ;
        RECT 235.500 689.400 237.300 702.000 ;
        RECT 248.400 695.400 250.200 702.000 ;
        RECT 251.400 695.400 253.200 701.400 ;
        RECT 236.100 682.050 237.900 683.850 ;
        RECT 251.850 682.050 253.050 695.400 ;
        RECT 256.500 689.400 258.300 702.000 ;
        RECT 266.400 695.400 268.200 701.400 ;
        RECT 269.400 695.400 271.200 702.000 ;
        RECT 266.400 688.500 267.600 695.400 ;
        RECT 272.400 689.400 274.200 701.400 ;
        RECT 286.800 695.400 288.600 702.000 ;
        RECT 289.800 695.400 291.600 701.400 ;
        RECT 292.800 695.400 294.600 702.000 ;
        RECT 266.400 687.600 272.100 688.500 ;
        RECT 270.150 686.700 272.100 687.600 ;
        RECT 257.100 682.050 258.900 683.850 ;
        RECT 266.100 682.050 267.900 683.850 ;
        RECT 163.950 679.800 166.050 681.900 ;
        RECT 166.950 679.800 169.050 681.900 ;
        RECT 169.950 679.800 172.050 681.900 ;
        RECT 172.950 679.800 175.050 681.900 ;
        RECT 181.950 679.800 184.050 681.900 ;
        RECT 184.950 679.800 187.050 681.900 ;
        RECT 187.950 679.800 190.050 681.900 ;
        RECT 190.950 679.800 193.050 681.900 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 211.950 679.950 214.050 682.050 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 235.950 679.950 238.050 682.050 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 256.950 679.950 259.050 682.050 ;
        RECT 265.950 679.950 268.050 682.050 ;
        RECT 147.900 674.400 149.850 675.300 ;
        RECT 164.700 676.200 165.600 679.800 ;
        RECT 167.100 678.000 168.900 679.800 ;
        RECT 173.100 678.000 174.900 679.800 ;
        RECT 182.100 678.000 183.900 679.800 ;
        RECT 188.100 678.000 189.900 679.800 ;
        RECT 191.400 676.200 192.300 679.800 ;
        RECT 206.100 678.150 207.900 679.950 ;
        RECT 164.700 675.000 168.000 676.200 ;
        RECT 147.900 673.500 153.600 674.400 ;
        RECT 109.500 666.000 111.300 672.600 ;
        RECT 119.700 666.000 121.500 672.600 ;
        RECT 124.200 666.600 126.000 672.600 ;
        RECT 128.700 666.000 130.500 672.600 ;
        RECT 145.800 666.600 147.600 672.600 ;
        RECT 152.400 669.600 153.600 673.500 ;
        RECT 148.800 666.000 150.600 669.600 ;
        RECT 151.800 666.600 153.600 669.600 ;
        RECT 166.200 666.600 168.000 675.000 ;
        RECT 172.800 666.000 174.600 675.600 ;
        RECT 182.400 666.000 184.200 675.600 ;
        RECT 189.000 675.000 192.300 676.200 ;
        RECT 209.850 675.750 211.050 679.950 ;
        RECT 212.100 678.150 213.900 679.950 ;
        RECT 227.100 678.150 228.900 679.950 ;
        RECT 229.950 675.750 231.150 679.950 ;
        RECT 233.100 678.150 234.900 679.950 ;
        RECT 248.100 678.150 249.900 679.950 ;
        RECT 250.950 675.750 252.150 679.950 ;
        RECT 254.100 678.150 255.900 679.950 ;
        RECT 189.000 666.600 190.800 675.000 ;
        RECT 209.850 674.700 213.600 675.750 ;
        RECT 203.400 671.700 211.200 673.050 ;
        RECT 203.400 666.600 205.200 671.700 ;
        RECT 206.400 666.000 208.200 670.800 ;
        RECT 209.400 666.600 211.200 671.700 ;
        RECT 212.400 672.600 213.600 674.700 ;
        RECT 227.400 674.700 231.150 675.750 ;
        RECT 248.400 674.700 252.150 675.750 ;
        RECT 270.150 675.300 271.050 686.700 ;
        RECT 273.000 682.050 274.200 689.400 ;
        RECT 271.950 679.950 274.200 682.050 ;
        RECT 290.400 681.900 291.600 695.400 ;
        RECT 304.800 689.400 306.600 701.400 ;
        RECT 307.800 695.400 309.600 702.000 ;
        RECT 310.800 695.400 312.600 701.400 ;
        RECT 313.800 695.400 315.600 702.000 ;
        RECT 323.400 695.400 325.200 702.000 ;
        RECT 326.400 695.400 328.200 701.400 ;
        RECT 329.400 696.000 331.200 702.000 ;
        RECT 305.400 681.900 306.300 689.400 ;
        RECT 308.100 681.900 309.900 683.700 ;
        RECT 227.400 672.600 228.600 674.700 ;
        RECT 212.400 666.600 214.200 672.600 ;
        RECT 226.800 666.600 228.600 672.600 ;
        RECT 229.800 671.700 237.600 673.050 ;
        RECT 248.400 672.600 249.600 674.700 ;
        RECT 270.150 674.400 272.100 675.300 ;
        RECT 266.400 673.500 272.100 674.400 ;
        RECT 229.800 666.600 231.600 671.700 ;
        RECT 232.800 666.000 234.600 670.800 ;
        RECT 235.800 666.600 237.600 671.700 ;
        RECT 247.800 666.600 249.600 672.600 ;
        RECT 250.800 671.700 258.600 673.050 ;
        RECT 250.800 666.600 252.600 671.700 ;
        RECT 253.800 666.000 255.600 670.800 ;
        RECT 256.800 666.600 258.600 671.700 ;
        RECT 266.400 669.600 267.600 673.500 ;
        RECT 273.000 672.600 274.200 679.950 ;
        RECT 286.950 679.800 289.050 681.900 ;
        RECT 289.950 679.800 292.050 681.900 ;
        RECT 292.950 679.800 295.050 681.900 ;
        RECT 304.950 679.800 307.050 681.900 ;
        RECT 307.950 679.800 310.050 681.900 ;
        RECT 287.100 678.000 288.900 679.800 ;
        RECT 290.400 674.700 291.600 679.800 ;
        RECT 293.100 678.000 294.900 679.800 ;
        RECT 266.400 666.600 268.200 669.600 ;
        RECT 269.400 666.000 271.200 669.600 ;
        RECT 272.400 666.600 274.200 672.600 ;
        RECT 287.400 673.800 291.600 674.700 ;
        RECT 287.400 666.600 289.200 673.800 ;
        RECT 305.400 672.600 306.300 679.800 ;
        RECT 311.700 675.300 312.600 695.400 ;
        RECT 326.700 695.100 328.200 695.400 ;
        RECT 332.400 695.400 334.200 701.400 ;
        RECT 346.800 695.400 348.600 702.000 ;
        RECT 349.800 695.400 351.600 701.400 ;
        RECT 352.800 695.400 354.600 702.000 ;
        RECT 362.400 695.400 364.200 702.000 ;
        RECT 365.400 695.400 367.200 701.400 ;
        RECT 368.400 696.000 370.200 702.000 ;
        RECT 332.400 695.100 333.300 695.400 ;
        RECT 326.700 694.200 333.300 695.100 ;
        RECT 326.100 681.900 327.900 683.700 ;
        RECT 332.400 681.900 333.300 694.200 ;
        RECT 342.000 684.450 346.050 685.050 ;
        RECT 341.550 682.950 346.050 684.450 ;
        RECT 313.950 679.800 316.050 681.900 ;
        RECT 322.950 679.800 325.050 681.900 ;
        RECT 325.950 679.800 328.050 681.900 ;
        RECT 328.950 679.800 331.050 681.900 ;
        RECT 331.950 679.800 334.050 681.900 ;
        RECT 314.100 678.000 315.900 679.800 ;
        RECT 323.100 678.000 324.900 679.800 ;
        RECT 329.100 678.000 330.900 679.800 ;
        RECT 332.400 676.200 333.300 679.800 ;
        RECT 341.550 679.050 342.450 682.950 ;
        RECT 350.400 681.900 351.600 695.400 ;
        RECT 365.700 695.100 367.200 695.400 ;
        RECT 371.400 695.400 373.200 701.400 ;
        RECT 385.800 695.400 387.600 701.400 ;
        RECT 388.800 696.000 390.600 702.000 ;
        RECT 371.400 695.100 372.300 695.400 ;
        RECT 365.700 694.200 372.300 695.100 ;
        RECT 365.100 681.900 366.900 683.700 ;
        RECT 371.400 681.900 372.300 694.200 ;
        RECT 386.700 695.100 387.600 695.400 ;
        RECT 391.800 695.400 393.600 701.400 ;
        RECT 394.800 695.400 396.600 702.000 ;
        RECT 391.800 695.100 393.300 695.400 ;
        RECT 386.700 694.200 393.300 695.100 ;
        RECT 386.700 681.900 387.600 694.200 ;
        RECT 404.400 690.300 406.200 701.400 ;
        RECT 407.400 691.200 409.200 702.000 ;
        RECT 410.400 690.300 412.200 701.400 ;
        RECT 404.400 689.400 412.200 690.300 ;
        RECT 413.400 689.400 415.200 701.400 ;
        RECT 427.800 689.400 429.600 701.400 ;
        RECT 430.800 690.300 432.600 701.400 ;
        RECT 433.800 691.200 435.600 702.000 ;
        RECT 436.800 690.300 438.600 701.400 ;
        RECT 446.400 695.400 448.200 702.000 ;
        RECT 449.400 695.400 451.200 701.400 ;
        RECT 452.400 696.000 454.200 702.000 ;
        RECT 449.700 695.100 451.200 695.400 ;
        RECT 455.400 695.400 457.200 701.400 ;
        RECT 467.400 695.400 469.200 702.000 ;
        RECT 470.400 695.400 472.200 701.400 ;
        RECT 455.400 695.100 456.300 695.400 ;
        RECT 449.700 694.200 456.300 695.100 ;
        RECT 430.800 689.400 438.600 690.300 ;
        RECT 388.950 687.450 391.050 688.050 ;
        RECT 403.950 687.450 406.050 688.050 ;
        RECT 388.950 686.550 406.050 687.450 ;
        RECT 388.950 685.950 391.050 686.550 ;
        RECT 403.950 685.950 406.050 686.550 ;
        RECT 392.100 681.900 393.900 683.700 ;
        RECT 407.100 681.900 408.900 683.700 ;
        RECT 413.700 681.900 414.600 689.400 ;
        RECT 415.950 684.450 420.000 685.050 ;
        RECT 415.950 682.950 420.450 684.450 ;
        RECT 346.950 679.800 349.050 681.900 ;
        RECT 349.950 679.800 352.050 681.900 ;
        RECT 352.950 679.800 355.050 681.900 ;
        RECT 361.950 679.800 364.050 681.900 ;
        RECT 364.950 679.800 367.050 681.900 ;
        RECT 367.950 679.800 370.050 681.900 ;
        RECT 370.950 679.800 373.050 681.900 ;
        RECT 385.950 679.800 388.050 681.900 ;
        RECT 388.950 679.800 391.050 681.900 ;
        RECT 391.950 679.800 394.050 681.900 ;
        RECT 394.950 679.800 397.050 681.900 ;
        RECT 403.950 679.800 406.050 681.900 ;
        RECT 406.950 679.800 409.050 681.900 ;
        RECT 409.950 679.800 412.050 681.900 ;
        RECT 412.950 679.800 415.050 681.900 ;
        RECT 341.550 677.550 346.050 679.050 ;
        RECT 347.100 678.000 348.900 679.800 ;
        RECT 342.000 676.950 346.050 677.550 ;
        RECT 308.100 674.400 315.600 675.300 ;
        RECT 308.100 673.500 309.900 674.400 ;
        RECT 292.500 666.000 294.300 672.600 ;
        RECT 305.400 670.800 308.100 672.600 ;
        RECT 306.300 666.600 308.100 670.800 ;
        RECT 309.300 666.000 311.100 672.600 ;
        RECT 313.800 666.600 315.600 674.400 ;
        RECT 323.400 666.000 325.200 675.600 ;
        RECT 330.000 675.000 333.300 676.200 ;
        RECT 330.000 666.600 331.800 675.000 ;
        RECT 350.400 674.700 351.600 679.800 ;
        RECT 353.100 678.000 354.900 679.800 ;
        RECT 362.100 678.000 363.900 679.800 ;
        RECT 368.100 678.000 369.900 679.800 ;
        RECT 371.400 676.200 372.300 679.800 ;
        RECT 347.400 673.800 351.600 674.700 ;
        RECT 347.400 666.600 349.200 673.800 ;
        RECT 352.500 666.000 354.300 672.600 ;
        RECT 362.400 666.000 364.200 675.600 ;
        RECT 369.000 675.000 372.300 676.200 ;
        RECT 386.700 676.200 387.600 679.800 ;
        RECT 389.100 678.000 390.900 679.800 ;
        RECT 395.100 678.000 396.900 679.800 ;
        RECT 404.100 678.000 405.900 679.800 ;
        RECT 410.100 678.000 411.900 679.800 ;
        RECT 386.700 675.000 390.000 676.200 ;
        RECT 369.000 666.600 370.800 675.000 ;
        RECT 388.200 666.600 390.000 675.000 ;
        RECT 394.800 666.000 396.600 675.600 ;
        RECT 413.700 672.600 414.600 679.800 ;
        RECT 419.550 679.050 420.450 682.950 ;
        RECT 428.400 681.900 429.300 689.400 ;
        RECT 434.100 681.900 435.900 683.700 ;
        RECT 449.100 681.900 450.900 683.700 ;
        RECT 455.400 681.900 456.300 694.200 ;
        RECT 467.100 682.050 468.900 683.850 ;
        RECT 470.400 682.050 471.600 695.400 ;
        RECT 482.700 689.400 484.500 702.000 ;
        RECT 487.800 695.400 489.600 701.400 ;
        RECT 490.800 695.400 492.600 702.000 ;
        RECT 503.400 695.400 505.200 702.000 ;
        RECT 506.400 695.400 508.200 701.400 ;
        RECT 520.800 695.400 522.600 701.400 ;
        RECT 523.800 696.000 525.600 702.000 ;
        RECT 472.950 684.450 477.000 685.050 ;
        RECT 472.950 682.950 477.450 684.450 ;
        RECT 427.950 679.800 430.050 681.900 ;
        RECT 430.950 679.800 433.050 681.900 ;
        RECT 433.950 679.800 436.050 681.900 ;
        RECT 436.950 679.800 439.050 681.900 ;
        RECT 445.950 679.800 448.050 681.900 ;
        RECT 448.950 679.800 451.050 681.900 ;
        RECT 451.950 679.800 454.050 681.900 ;
        RECT 454.950 679.800 457.050 681.900 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 415.950 677.550 420.450 679.050 ;
        RECT 415.950 676.950 420.000 677.550 ;
        RECT 405.000 666.000 406.800 672.600 ;
        RECT 409.500 671.400 414.600 672.600 ;
        RECT 428.400 672.600 429.300 679.800 ;
        RECT 431.100 678.000 432.900 679.800 ;
        RECT 437.100 678.000 438.900 679.800 ;
        RECT 446.100 678.000 447.900 679.800 ;
        RECT 452.100 678.000 453.900 679.800 ;
        RECT 455.400 676.200 456.300 679.800 ;
        RECT 428.400 671.400 433.500 672.600 ;
        RECT 409.500 666.600 411.300 671.400 ;
        RECT 412.500 666.000 414.300 669.600 ;
        RECT 428.700 666.000 430.500 669.600 ;
        RECT 431.700 666.600 433.500 671.400 ;
        RECT 436.200 666.000 438.000 672.600 ;
        RECT 446.400 666.000 448.200 675.600 ;
        RECT 453.000 675.000 456.300 676.200 ;
        RECT 453.000 666.600 454.800 675.000 ;
        RECT 470.400 669.600 471.600 679.950 ;
        RECT 476.550 679.050 477.450 682.950 ;
        RECT 482.100 682.050 483.900 683.850 ;
        RECT 487.950 682.050 489.150 695.400 ;
        RECT 498.000 684.450 502.050 685.050 ;
        RECT 497.550 682.950 502.050 684.450 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 484.950 679.950 487.050 682.050 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 490.950 679.950 493.050 682.050 ;
        RECT 476.550 677.550 481.050 679.050 ;
        RECT 485.100 678.150 486.900 679.950 ;
        RECT 477.000 676.950 481.050 677.550 ;
        RECT 488.850 675.750 490.050 679.950 ;
        RECT 491.100 678.150 492.900 679.950 ;
        RECT 497.550 679.050 498.450 682.950 ;
        RECT 503.100 682.050 504.900 683.850 ;
        RECT 506.400 682.050 507.600 695.400 ;
        RECT 521.700 695.100 522.600 695.400 ;
        RECT 526.800 695.400 528.600 701.400 ;
        RECT 529.800 695.400 531.600 702.000 ;
        RECT 539.400 695.400 541.200 702.000 ;
        RECT 542.400 695.400 544.200 701.400 ;
        RECT 545.400 695.400 547.200 702.000 ;
        RECT 557.400 695.400 559.200 702.000 ;
        RECT 560.400 695.400 562.200 701.400 ;
        RECT 526.800 695.100 528.300 695.400 ;
        RECT 521.700 694.200 528.300 695.100 ;
        RECT 508.950 684.450 511.050 685.050 ;
        RECT 508.950 683.550 516.450 684.450 ;
        RECT 508.950 682.950 511.050 683.550 ;
        RECT 502.950 679.950 505.050 682.050 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 493.950 677.550 498.450 679.050 ;
        RECT 493.950 676.950 498.000 677.550 ;
        RECT 488.850 674.700 492.600 675.750 ;
        RECT 482.400 671.700 490.200 673.050 ;
        RECT 467.400 666.000 469.200 669.600 ;
        RECT 470.400 666.600 472.200 669.600 ;
        RECT 482.400 666.600 484.200 671.700 ;
        RECT 485.400 666.000 487.200 670.800 ;
        RECT 488.400 666.600 490.200 671.700 ;
        RECT 491.400 672.600 492.600 674.700 ;
        RECT 491.400 666.600 493.200 672.600 ;
        RECT 506.400 669.600 507.600 679.950 ;
        RECT 515.550 679.050 516.450 683.550 ;
        RECT 521.700 681.900 522.600 694.200 ;
        RECT 529.950 687.450 532.050 688.050 ;
        RECT 535.950 687.450 538.050 688.050 ;
        RECT 529.950 686.550 538.050 687.450 ;
        RECT 529.950 685.950 532.050 686.550 ;
        RECT 535.950 685.950 538.050 686.550 ;
        RECT 532.950 684.450 535.050 685.050 ;
        RECT 538.950 684.450 541.050 684.900 ;
        RECT 527.100 681.900 528.900 683.700 ;
        RECT 532.950 683.550 541.050 684.450 ;
        RECT 532.950 682.950 535.050 683.550 ;
        RECT 538.950 682.800 541.050 683.550 ;
        RECT 542.400 681.900 543.600 695.400 ;
        RECT 557.100 682.050 558.900 683.850 ;
        RECT 560.400 682.050 561.600 695.400 ;
        RECT 572.400 689.400 574.200 702.000 ;
        RECT 575.400 689.400 577.200 701.400 ;
        RECT 589.800 695.400 591.600 702.000 ;
        RECT 592.800 695.400 594.600 701.400 ;
        RECT 595.800 695.400 597.600 702.000 ;
        RECT 607.800 695.400 609.600 702.000 ;
        RECT 610.800 695.400 612.600 701.400 ;
        RECT 613.800 695.400 615.600 702.000 ;
        RECT 520.950 679.800 523.050 681.900 ;
        RECT 523.950 679.800 526.050 681.900 ;
        RECT 526.950 679.800 529.050 681.900 ;
        RECT 529.950 679.800 532.050 681.900 ;
        RECT 538.950 679.800 541.050 681.900 ;
        RECT 541.950 679.800 544.050 681.900 ;
        RECT 544.950 679.800 547.050 681.900 ;
        RECT 556.950 679.950 559.050 682.050 ;
        RECT 559.950 679.950 562.050 682.050 ;
        RECT 575.400 681.900 576.600 689.400 ;
        RECT 593.400 681.900 594.600 695.400 ;
        RECT 611.400 681.900 612.600 695.400 ;
        RECT 623.400 690.300 625.200 701.400 ;
        RECT 630.900 690.300 632.700 701.400 ;
        RECT 638.400 690.600 640.200 701.400 ;
        RECT 623.400 689.100 628.200 690.300 ;
        RECT 630.900 689.400 634.200 690.300 ;
        RECT 626.100 688.200 628.200 689.100 ;
        RECT 626.100 687.300 631.350 688.200 ;
        RECT 629.550 685.200 631.350 687.300 ;
        RECT 633.000 684.900 634.200 689.400 ;
        RECT 635.100 689.400 640.200 690.600 ;
        RECT 650.700 689.400 652.500 702.000 ;
        RECT 655.800 695.400 657.600 701.400 ;
        RECT 658.800 695.400 660.600 702.000 ;
        RECT 635.100 688.500 637.200 689.400 ;
        RECT 632.250 684.300 634.350 684.900 ;
        RECT 628.200 682.200 630.000 684.000 ;
        RECT 631.350 682.800 634.350 684.300 ;
        RECT 638.550 683.700 645.450 684.450 ;
        RECT 638.100 683.550 645.450 683.700 ;
        RECT 515.550 677.550 520.050 679.050 ;
        RECT 516.000 676.950 520.050 677.550 ;
        RECT 521.700 676.200 522.600 679.800 ;
        RECT 524.100 678.000 525.900 679.800 ;
        RECT 530.100 678.000 531.900 679.800 ;
        RECT 539.100 678.000 540.900 679.800 ;
        RECT 521.700 675.000 525.000 676.200 ;
        RECT 503.400 666.000 505.200 669.600 ;
        RECT 506.400 666.600 508.200 669.600 ;
        RECT 523.200 666.600 525.000 675.000 ;
        RECT 529.800 666.000 531.600 675.600 ;
        RECT 542.400 674.700 543.600 679.800 ;
        RECT 545.100 678.000 546.900 679.800 ;
        RECT 547.950 675.450 550.050 676.050 ;
        RECT 556.950 675.450 559.050 676.050 ;
        RECT 542.400 673.800 546.600 674.700 ;
        RECT 547.950 674.550 559.050 675.450 ;
        RECT 547.950 673.950 550.050 674.550 ;
        RECT 556.950 673.950 559.050 674.550 ;
        RECT 539.700 666.000 541.500 672.600 ;
        RECT 544.800 666.600 546.600 673.800 ;
        RECT 560.400 669.600 561.600 679.950 ;
        RECT 571.950 679.800 574.050 681.900 ;
        RECT 574.950 679.800 577.050 681.900 ;
        RECT 589.950 679.800 592.050 681.900 ;
        RECT 592.950 679.800 595.050 681.900 ;
        RECT 595.950 679.800 598.050 681.900 ;
        RECT 607.950 679.800 610.050 681.900 ;
        RECT 610.950 679.800 613.050 681.900 ;
        RECT 613.950 679.800 616.050 681.900 ;
        RECT 622.950 679.800 625.050 681.900 ;
        RECT 628.200 680.100 630.300 682.200 ;
        RECT 572.100 678.000 573.900 679.800 ;
        RECT 575.400 672.600 576.600 679.800 ;
        RECT 590.100 678.000 591.900 679.800 ;
        RECT 593.400 674.700 594.600 679.800 ;
        RECT 596.100 678.000 597.900 679.800 ;
        RECT 608.100 678.000 609.900 679.800 ;
        RECT 611.400 674.700 612.600 679.800 ;
        RECT 614.100 678.000 615.900 679.800 ;
        RECT 623.250 679.200 625.050 679.800 ;
        RECT 623.250 678.000 630.300 679.200 ;
        RECT 628.200 677.100 630.300 678.000 ;
        RECT 625.650 675.000 627.750 675.600 ;
        RECT 628.650 675.300 630.450 677.100 ;
        RECT 631.350 676.200 632.250 682.800 ;
        RECT 638.100 681.900 639.900 683.550 ;
        RECT 633.300 680.100 635.100 681.900 ;
        RECT 633.150 678.000 635.250 680.100 ;
        RECT 637.950 679.800 640.050 681.900 ;
        RECT 644.550 679.050 645.450 683.550 ;
        RECT 650.100 682.050 651.900 683.850 ;
        RECT 655.950 682.050 657.150 695.400 ;
        RECT 671.400 690.300 673.200 701.400 ;
        RECT 678.900 697.050 680.700 701.400 ;
        RECT 678.900 694.950 682.050 697.050 ;
        RECT 671.400 689.400 675.900 690.300 ;
        RECT 678.900 689.400 680.700 694.950 ;
        RECT 686.400 690.600 688.200 701.400 ;
        RECT 698.400 695.400 700.200 702.000 ;
        RECT 701.400 695.400 703.200 701.400 ;
        RECT 704.400 696.000 706.200 702.000 ;
        RECT 701.700 695.100 703.200 695.400 ;
        RECT 707.400 695.400 709.200 701.400 ;
        RECT 719.400 695.400 721.200 702.000 ;
        RECT 722.400 695.400 724.200 701.400 ;
        RECT 725.400 696.000 727.200 702.000 ;
        RECT 707.400 695.100 708.300 695.400 ;
        RECT 701.700 694.200 708.300 695.100 ;
        RECT 722.700 695.100 724.200 695.400 ;
        RECT 728.400 695.400 730.200 701.400 ;
        RECT 743.400 695.400 745.200 702.000 ;
        RECT 746.400 695.400 748.200 701.400 ;
        RECT 728.400 695.100 729.300 695.400 ;
        RECT 722.700 694.200 729.300 695.100 ;
        RECT 673.800 687.300 675.900 689.400 ;
        RECT 679.500 687.900 680.700 689.400 ;
        RECT 683.400 689.400 688.200 690.600 ;
        RECT 683.400 688.500 685.500 689.400 ;
        RECT 679.500 687.000 681.000 687.900 ;
        RECT 676.950 685.500 679.050 685.800 ;
        RECT 675.300 683.700 679.050 685.500 ;
        RECT 680.100 684.900 681.000 687.000 ;
        RECT 679.950 682.800 682.050 684.900 ;
        RECT 691.950 684.450 694.050 685.050 ;
        RECT 686.550 683.700 694.050 684.450 ;
        RECT 686.100 683.550 694.050 683.700 ;
        RECT 649.950 679.950 652.050 682.050 ;
        RECT 652.950 679.950 655.050 682.050 ;
        RECT 655.950 679.950 658.050 682.050 ;
        RECT 658.950 679.950 661.050 682.050 ;
        RECT 676.500 681.900 678.300 682.500 ;
        RECT 670.950 680.700 678.300 681.900 ;
        RECT 679.200 681.900 681.600 682.800 ;
        RECT 686.100 681.900 687.900 683.550 ;
        RECT 691.950 682.950 694.050 683.550 ;
        RECT 701.100 681.900 702.900 683.700 ;
        RECT 707.400 681.900 708.300 694.200 ;
        RECT 722.100 681.900 723.900 683.700 ;
        RECT 728.400 681.900 729.300 694.200 ;
        RECT 746.850 682.050 748.050 695.400 ;
        RECT 751.500 689.400 753.300 702.000 ;
        RECT 761.700 689.400 763.500 702.000 ;
        RECT 766.800 695.400 768.600 701.400 ;
        RECT 769.800 695.400 771.600 702.000 ;
        RECT 782.400 695.400 784.200 702.000 ;
        RECT 785.400 695.400 787.200 701.400 ;
        RECT 799.800 695.400 801.600 701.400 ;
        RECT 802.800 695.400 804.600 702.000 ;
        RECT 812.400 695.400 814.200 702.000 ;
        RECT 815.400 695.400 817.200 701.400 ;
        RECT 818.400 696.000 820.200 702.000 ;
        RECT 752.100 682.050 753.900 683.850 ;
        RECT 761.100 682.050 762.900 683.850 ;
        RECT 766.950 682.050 768.150 695.400 ;
        RECT 782.100 682.050 783.900 683.850 ;
        RECT 785.400 682.050 786.600 695.400 ;
        RECT 800.400 682.050 801.600 695.400 ;
        RECT 815.700 695.100 817.200 695.400 ;
        RECT 821.400 695.400 823.200 701.400 ;
        RECT 833.400 695.400 835.200 702.000 ;
        RECT 836.400 695.400 838.200 701.400 ;
        RECT 839.400 696.000 841.200 702.000 ;
        RECT 821.400 695.100 822.300 695.400 ;
        RECT 815.700 694.200 822.300 695.100 ;
        RECT 836.700 695.100 838.200 695.400 ;
        RECT 842.400 695.400 844.200 701.400 ;
        RECT 842.400 695.100 843.300 695.400 ;
        RECT 836.700 694.200 843.300 695.100 ;
        RECT 803.100 682.050 804.900 683.850 ;
        RECT 644.550 677.550 649.050 679.050 ;
        RECT 653.100 678.150 654.900 679.950 ;
        RECT 645.000 676.950 649.050 677.550 ;
        RECT 590.400 673.800 594.600 674.700 ;
        RECT 608.400 673.800 612.600 674.700 ;
        RECT 557.400 666.000 559.200 669.600 ;
        RECT 560.400 666.600 562.200 669.600 ;
        RECT 572.400 666.000 574.200 672.600 ;
        RECT 575.400 666.600 577.200 672.600 ;
        RECT 590.400 666.600 592.200 673.800 ;
        RECT 595.500 666.000 597.300 672.600 ;
        RECT 608.400 666.600 610.200 673.800 ;
        RECT 623.400 673.500 627.750 675.000 ;
        RECT 631.350 674.100 634.350 676.200 ;
        RECT 623.400 672.600 624.900 673.500 ;
        RECT 613.500 666.000 615.300 672.600 ;
        RECT 623.400 666.600 625.200 672.600 ;
        RECT 631.350 672.000 632.250 674.100 ;
        RECT 635.700 673.500 637.800 675.900 ;
        RECT 656.850 675.750 658.050 679.950 ;
        RECT 659.100 678.150 660.900 679.950 ;
        RECT 670.950 679.800 673.050 680.700 ;
        RECT 671.250 678.000 673.050 679.800 ;
        RECT 676.500 677.400 678.300 679.200 ;
        RECT 656.850 674.700 660.600 675.750 ;
        RECT 676.200 675.300 678.300 677.400 ;
        RECT 635.700 672.600 640.200 673.500 ;
        RECT 630.600 666.600 632.400 672.000 ;
        RECT 638.400 666.600 640.200 672.600 ;
        RECT 650.400 671.700 658.200 673.050 ;
        RECT 650.400 666.600 652.200 671.700 ;
        RECT 653.400 666.000 655.200 670.800 ;
        RECT 656.400 666.600 658.200 671.700 ;
        RECT 659.400 672.600 660.600 674.700 ;
        RECT 672.000 674.400 678.300 675.300 ;
        RECT 679.200 676.200 680.250 681.900 ;
        RECT 681.600 679.200 683.400 681.000 ;
        RECT 685.950 679.800 688.050 681.900 ;
        RECT 697.950 679.800 700.050 681.900 ;
        RECT 700.950 679.800 703.050 681.900 ;
        RECT 703.950 679.800 706.050 681.900 ;
        RECT 706.950 679.800 709.050 681.900 ;
        RECT 718.950 679.800 721.050 681.900 ;
        RECT 721.950 679.800 724.050 681.900 ;
        RECT 724.950 679.800 727.050 681.900 ;
        RECT 727.950 679.800 730.050 681.900 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 748.950 679.950 751.050 682.050 ;
        RECT 751.950 679.950 754.050 682.050 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 769.950 679.950 772.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 784.950 679.950 787.050 682.050 ;
        RECT 799.950 679.950 802.050 682.050 ;
        RECT 802.950 679.950 805.050 682.050 ;
        RECT 815.100 681.900 816.900 683.700 ;
        RECT 821.400 681.900 822.300 694.200 ;
        RECT 836.100 681.900 837.900 683.700 ;
        RECT 842.400 681.900 843.300 694.200 ;
        RECT 681.150 677.100 683.250 679.200 ;
        RECT 698.100 678.000 699.900 679.800 ;
        RECT 704.100 678.000 705.900 679.800 ;
        RECT 707.400 676.200 708.300 679.800 ;
        RECT 719.100 678.000 720.900 679.800 ;
        RECT 725.100 678.000 726.900 679.800 ;
        RECT 728.400 676.200 729.300 679.800 ;
        RECT 743.100 678.150 744.900 679.950 ;
        RECT 672.000 672.600 673.200 674.400 ;
        RECT 679.200 674.100 682.050 676.200 ;
        RECT 679.200 672.600 680.400 674.100 ;
        RECT 683.400 673.500 685.500 674.700 ;
        RECT 683.400 672.600 688.200 673.500 ;
        RECT 659.400 666.600 661.200 672.600 ;
        RECT 671.400 666.600 673.200 672.600 ;
        RECT 678.900 666.600 680.700 672.600 ;
        RECT 686.400 666.600 688.200 672.600 ;
        RECT 698.400 666.000 700.200 675.600 ;
        RECT 705.000 675.000 708.300 676.200 ;
        RECT 705.000 666.600 706.800 675.000 ;
        RECT 719.400 666.000 721.200 675.600 ;
        RECT 726.000 675.000 729.300 676.200 ;
        RECT 745.950 675.750 747.150 679.950 ;
        RECT 749.100 678.150 750.900 679.950 ;
        RECT 764.100 678.150 765.900 679.950 ;
        RECT 726.000 666.600 727.800 675.000 ;
        RECT 743.400 674.700 747.150 675.750 ;
        RECT 767.850 675.750 769.050 679.950 ;
        RECT 770.100 678.150 771.900 679.950 ;
        RECT 767.850 674.700 771.600 675.750 ;
        RECT 743.400 672.600 744.600 674.700 ;
        RECT 742.800 666.600 744.600 672.600 ;
        RECT 745.800 671.700 753.600 673.050 ;
        RECT 745.800 666.600 747.600 671.700 ;
        RECT 748.800 666.000 750.600 670.800 ;
        RECT 751.800 666.600 753.600 671.700 ;
        RECT 761.400 671.700 769.200 673.050 ;
        RECT 761.400 666.600 763.200 671.700 ;
        RECT 764.400 666.000 766.200 670.800 ;
        RECT 767.400 666.600 769.200 671.700 ;
        RECT 770.400 672.600 771.600 674.700 ;
        RECT 770.400 666.600 772.200 672.600 ;
        RECT 785.400 669.600 786.600 679.950 ;
        RECT 800.400 669.600 801.600 679.950 ;
        RECT 811.950 679.800 814.050 681.900 ;
        RECT 814.950 679.800 817.050 681.900 ;
        RECT 817.950 679.800 820.050 681.900 ;
        RECT 820.950 679.800 823.050 681.900 ;
        RECT 832.950 679.800 835.050 681.900 ;
        RECT 835.950 679.800 838.050 681.900 ;
        RECT 838.950 679.800 841.050 681.900 ;
        RECT 841.950 679.800 844.050 681.900 ;
        RECT 812.100 678.000 813.900 679.800 ;
        RECT 818.100 678.000 819.900 679.800 ;
        RECT 821.400 676.200 822.300 679.800 ;
        RECT 833.100 678.000 834.900 679.800 ;
        RECT 839.100 678.000 840.900 679.800 ;
        RECT 842.400 676.200 843.300 679.800 ;
        RECT 782.400 666.000 784.200 669.600 ;
        RECT 785.400 666.600 787.200 669.600 ;
        RECT 799.800 666.600 801.600 669.600 ;
        RECT 802.800 666.000 804.600 669.600 ;
        RECT 812.400 666.000 814.200 675.600 ;
        RECT 819.000 675.000 822.300 676.200 ;
        RECT 819.000 666.600 820.800 675.000 ;
        RECT 833.400 666.000 835.200 675.600 ;
        RECT 840.000 675.000 843.300 676.200 ;
        RECT 840.000 666.600 841.800 675.000 ;
        RECT 10.800 659.400 12.600 662.400 ;
        RECT 13.800 659.400 15.600 663.000 ;
        RECT 11.400 649.050 12.600 659.400 ;
        RECT 25.800 656.400 27.600 662.400 ;
        RECT 13.950 654.450 16.050 654.900 ;
        RECT 22.950 654.450 25.050 655.050 ;
        RECT 13.950 653.550 25.050 654.450 ;
        RECT 13.950 652.800 16.050 653.550 ;
        RECT 22.950 652.950 25.050 653.550 ;
        RECT 26.400 654.300 27.600 656.400 ;
        RECT 28.800 657.300 30.600 662.400 ;
        RECT 31.800 658.200 33.600 663.000 ;
        RECT 34.800 657.300 36.600 662.400 ;
        RECT 28.800 655.950 36.600 657.300 ;
        RECT 44.400 657.300 46.200 662.400 ;
        RECT 47.400 658.200 49.200 663.000 ;
        RECT 50.400 657.300 52.200 662.400 ;
        RECT 44.400 655.950 52.200 657.300 ;
        RECT 53.400 656.400 55.200 662.400 ;
        RECT 53.400 654.300 54.600 656.400 ;
        RECT 26.400 653.250 30.150 654.300 ;
        RECT 26.100 649.050 27.900 650.850 ;
        RECT 28.950 649.050 30.150 653.250 ;
        RECT 50.850 653.250 54.600 654.300 ;
        RECT 65.400 653.400 67.200 663.000 ;
        RECT 72.000 654.000 73.800 662.400 ;
        RECT 87.000 656.400 88.800 663.000 ;
        RECT 91.500 657.600 93.300 662.400 ;
        RECT 94.500 659.400 96.300 663.000 ;
        RECT 111.300 658.200 113.100 662.400 ;
        RECT 91.500 656.400 96.600 657.600 ;
        RECT 32.100 649.050 33.900 650.850 ;
        RECT 47.100 649.050 48.900 650.850 ;
        RECT 50.850 649.050 52.050 653.250 ;
        RECT 72.000 652.800 75.300 654.000 ;
        RECT 53.100 649.050 54.900 650.850 ;
        RECT 65.100 649.200 66.900 651.000 ;
        RECT 71.100 649.200 72.900 651.000 ;
        RECT 74.400 649.200 75.300 652.800 ;
        RECT 76.950 651.450 81.000 652.050 ;
        RECT 76.950 649.950 81.450 651.450 ;
        RECT 10.950 646.950 13.050 649.050 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 25.950 646.950 28.050 649.050 ;
        RECT 28.950 646.950 31.050 649.050 ;
        RECT 31.950 646.950 34.050 649.050 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 43.950 646.950 46.050 649.050 ;
        RECT 46.950 646.950 49.050 649.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 52.950 646.950 55.050 649.050 ;
        RECT 64.950 647.100 67.050 649.200 ;
        RECT 67.950 647.100 70.050 649.200 ;
        RECT 70.950 647.100 73.050 649.200 ;
        RECT 73.950 647.100 76.050 649.200 ;
        RECT 11.400 633.600 12.600 646.950 ;
        RECT 14.100 645.150 15.900 646.950 ;
        RECT 29.850 633.600 31.050 646.950 ;
        RECT 35.100 645.150 36.900 646.950 ;
        RECT 44.100 645.150 45.900 646.950 ;
        RECT 10.800 627.600 12.600 633.600 ;
        RECT 13.800 627.000 15.600 633.600 ;
        RECT 26.400 627.000 28.200 633.600 ;
        RECT 29.400 627.600 31.200 633.600 ;
        RECT 34.500 627.000 36.300 639.600 ;
        RECT 44.700 627.000 46.500 639.600 ;
        RECT 49.950 633.600 51.150 646.950 ;
        RECT 68.100 645.300 69.900 647.100 ;
        RECT 74.400 634.800 75.300 647.100 ;
        RECT 80.550 646.050 81.450 649.950 ;
        RECT 86.100 649.200 87.900 651.000 ;
        RECT 92.100 649.200 93.900 651.000 ;
        RECT 95.700 649.200 96.600 656.400 ;
        RECT 110.400 656.400 113.100 658.200 ;
        RECT 114.300 656.400 116.100 663.000 ;
        RECT 100.950 654.450 103.050 655.050 ;
        RECT 106.950 654.450 109.050 655.050 ;
        RECT 100.950 653.550 109.050 654.450 ;
        RECT 100.950 652.950 103.050 653.550 ;
        RECT 106.950 652.950 109.050 653.550 ;
        RECT 97.950 651.450 100.050 652.050 ;
        RECT 103.950 651.450 106.050 652.050 ;
        RECT 97.950 650.550 106.050 651.450 ;
        RECT 97.950 649.950 100.050 650.550 ;
        RECT 103.950 649.950 106.050 650.550 ;
        RECT 110.400 649.200 111.300 656.400 ;
        RECT 113.100 654.600 114.900 655.500 ;
        RECT 118.800 654.600 120.600 662.400 ;
        RECT 128.700 656.400 130.500 663.000 ;
        RECT 133.800 655.200 135.600 662.400 ;
        RECT 146.400 659.400 148.200 663.000 ;
        RECT 149.400 659.400 151.200 662.400 ;
        RECT 113.100 653.700 120.600 654.600 ;
        RECT 131.400 654.300 135.600 655.200 ;
        RECT 85.950 647.100 88.050 649.200 ;
        RECT 88.950 647.100 91.050 649.200 ;
        RECT 91.950 647.100 94.050 649.200 ;
        RECT 94.950 647.100 97.050 649.200 ;
        RECT 109.950 647.100 112.050 649.200 ;
        RECT 112.950 647.100 115.050 649.200 ;
        RECT 76.950 644.550 81.450 646.050 ;
        RECT 89.100 645.300 90.900 647.100 ;
        RECT 76.950 643.950 81.000 644.550 ;
        RECT 95.700 639.600 96.600 647.100 ;
        RECT 110.400 639.600 111.300 647.100 ;
        RECT 113.100 645.300 114.900 647.100 ;
        RECT 68.700 633.900 75.300 634.800 ;
        RECT 68.700 633.600 70.200 633.900 ;
        RECT 49.800 627.600 51.600 633.600 ;
        RECT 52.800 627.000 54.600 633.600 ;
        RECT 65.400 627.000 67.200 633.600 ;
        RECT 68.400 627.600 70.200 633.600 ;
        RECT 74.400 633.600 75.300 633.900 ;
        RECT 86.400 638.700 94.200 639.600 ;
        RECT 71.400 627.000 73.200 633.000 ;
        RECT 74.400 627.600 76.200 633.600 ;
        RECT 86.400 627.600 88.200 638.700 ;
        RECT 89.400 627.000 91.200 637.800 ;
        RECT 92.400 627.600 94.200 638.700 ;
        RECT 95.400 627.600 97.200 639.600 ;
        RECT 109.800 627.600 111.600 639.600 ;
        RECT 116.700 633.600 117.600 653.700 ;
        RECT 119.100 649.200 120.900 651.000 ;
        RECT 128.100 649.200 129.900 651.000 ;
        RECT 131.400 649.200 132.600 654.300 ;
        RECT 134.100 649.200 135.900 651.000 ;
        RECT 118.950 647.100 121.050 649.200 ;
        RECT 127.950 647.100 130.050 649.200 ;
        RECT 130.950 647.100 133.050 649.200 ;
        RECT 133.950 647.100 136.050 649.200 ;
        RECT 149.400 649.050 150.600 659.400 ;
        RECT 161.700 656.400 163.500 663.000 ;
        RECT 166.800 655.200 168.600 662.400 ;
        RECT 181.800 659.400 183.600 662.400 ;
        RECT 184.800 659.400 186.600 663.000 ;
        RECT 164.400 654.300 168.600 655.200 ;
        RECT 161.100 649.200 162.900 651.000 ;
        RECT 164.400 649.200 165.600 654.300 ;
        RECT 167.100 649.200 168.900 651.000 ;
        RECT 131.400 633.600 132.600 647.100 ;
        RECT 145.950 646.950 148.050 649.050 ;
        RECT 148.950 646.950 151.050 649.050 ;
        RECT 160.950 647.100 163.050 649.200 ;
        RECT 163.950 647.100 166.050 649.200 ;
        RECT 166.950 647.100 169.050 649.200 ;
        RECT 182.400 649.050 183.600 659.400 ;
        RECT 199.200 654.000 201.000 662.400 ;
        RECT 197.700 652.800 201.000 654.000 ;
        RECT 205.800 653.400 207.600 663.000 ;
        RECT 216.000 656.400 217.800 663.000 ;
        RECT 220.500 657.600 222.300 662.400 ;
        RECT 223.500 659.400 225.300 663.000 ;
        RECT 236.400 659.400 238.200 663.000 ;
        RECT 239.400 659.400 241.200 662.400 ;
        RECT 220.500 656.400 225.600 657.600 ;
        RECT 192.000 651.450 196.050 652.050 ;
        RECT 191.550 649.950 196.050 651.450 ;
        RECT 146.100 645.150 147.900 646.950 ;
        RECT 149.400 633.600 150.600 646.950 ;
        RECT 164.400 633.600 165.600 647.100 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 182.400 633.600 183.600 646.950 ;
        RECT 185.100 645.150 186.900 646.950 ;
        RECT 191.550 646.050 192.450 649.950 ;
        RECT 197.700 649.200 198.600 652.800 ;
        RECT 200.100 649.200 201.900 651.000 ;
        RECT 206.100 649.200 207.900 651.000 ;
        RECT 215.100 649.200 216.900 651.000 ;
        RECT 221.100 649.200 222.900 651.000 ;
        RECT 224.700 649.200 225.600 656.400 ;
        RECT 196.950 647.100 199.050 649.200 ;
        RECT 199.950 647.100 202.050 649.200 ;
        RECT 202.950 647.100 205.050 649.200 ;
        RECT 205.950 647.100 208.050 649.200 ;
        RECT 214.950 647.100 217.050 649.200 ;
        RECT 217.950 647.100 220.050 649.200 ;
        RECT 220.950 647.100 223.050 649.200 ;
        RECT 223.950 647.100 226.050 649.200 ;
        RECT 239.400 649.050 240.600 659.400 ;
        RECT 252.000 656.400 253.800 663.000 ;
        RECT 256.500 657.600 258.300 662.400 ;
        RECT 259.500 659.400 261.300 663.000 ;
        RECT 256.500 656.400 261.600 657.600 ;
        RECT 251.100 649.200 252.900 651.000 ;
        RECT 257.100 649.200 258.900 651.000 ;
        RECT 260.700 649.200 261.600 656.400 ;
        RECT 272.400 654.600 274.200 662.400 ;
        RECT 276.900 656.400 278.700 663.000 ;
        RECT 279.900 658.200 281.700 662.400 ;
        RECT 279.900 656.400 282.600 658.200 ;
        RECT 278.100 654.600 279.900 655.500 ;
        RECT 272.400 653.700 279.900 654.600 ;
        RECT 272.100 649.200 273.900 651.000 ;
        RECT 187.950 644.550 192.450 646.050 ;
        RECT 187.950 643.950 192.000 644.550 ;
        RECT 197.700 634.800 198.600 647.100 ;
        RECT 203.100 645.300 204.900 647.100 ;
        RECT 218.100 645.300 219.900 647.100 ;
        RECT 199.950 642.450 202.050 643.050 ;
        RECT 214.950 642.450 217.050 643.050 ;
        RECT 199.950 641.550 217.050 642.450 ;
        RECT 199.950 640.950 202.050 641.550 ;
        RECT 214.950 640.950 217.050 641.550 ;
        RECT 202.950 639.450 205.050 640.050 ;
        RECT 208.950 639.450 211.050 640.050 ;
        RECT 224.700 639.600 225.600 647.100 ;
        RECT 235.950 646.950 238.050 649.050 ;
        RECT 238.950 646.950 241.050 649.050 ;
        RECT 250.950 647.100 253.050 649.200 ;
        RECT 253.950 647.100 256.050 649.200 ;
        RECT 256.950 647.100 259.050 649.200 ;
        RECT 259.950 647.100 262.050 649.200 ;
        RECT 271.950 647.100 274.050 649.200 ;
        RECT 236.100 645.150 237.900 646.950 ;
        RECT 202.950 638.550 211.050 639.450 ;
        RECT 202.950 637.950 205.050 638.550 ;
        RECT 208.950 637.950 211.050 638.550 ;
        RECT 215.400 638.700 223.200 639.600 ;
        RECT 197.700 633.900 204.300 634.800 ;
        RECT 197.700 633.600 198.600 633.900 ;
        RECT 112.800 627.000 114.600 633.600 ;
        RECT 115.800 627.600 117.600 633.600 ;
        RECT 118.800 627.000 120.600 633.600 ;
        RECT 128.400 627.000 130.200 633.600 ;
        RECT 131.400 627.600 133.200 633.600 ;
        RECT 134.400 627.000 136.200 633.600 ;
        RECT 146.400 627.000 148.200 633.600 ;
        RECT 149.400 627.600 151.200 633.600 ;
        RECT 161.400 627.000 163.200 633.600 ;
        RECT 164.400 627.600 166.200 633.600 ;
        RECT 167.400 627.000 169.200 633.600 ;
        RECT 181.800 627.600 183.600 633.600 ;
        RECT 184.800 627.000 186.600 633.600 ;
        RECT 196.800 627.600 198.600 633.600 ;
        RECT 202.800 633.600 204.300 633.900 ;
        RECT 199.800 627.000 201.600 633.000 ;
        RECT 202.800 627.600 204.600 633.600 ;
        RECT 205.800 627.000 207.600 633.600 ;
        RECT 215.400 627.600 217.200 638.700 ;
        RECT 218.400 627.000 220.200 637.800 ;
        RECT 221.400 627.600 223.200 638.700 ;
        RECT 224.400 627.600 226.200 639.600 ;
        RECT 239.400 633.600 240.600 646.950 ;
        RECT 254.100 645.300 255.900 647.100 ;
        RECT 241.950 642.450 244.050 643.050 ;
        RECT 256.950 642.450 259.050 643.050 ;
        RECT 241.950 641.550 259.050 642.450 ;
        RECT 241.950 640.950 244.050 641.550 ;
        RECT 256.950 640.950 259.050 641.550 ;
        RECT 260.700 639.600 261.600 647.100 ;
        RECT 251.400 638.700 259.200 639.600 ;
        RECT 236.400 627.000 238.200 633.600 ;
        RECT 239.400 627.600 241.200 633.600 ;
        RECT 251.400 627.600 253.200 638.700 ;
        RECT 254.400 627.000 256.200 637.800 ;
        RECT 257.400 627.600 259.200 638.700 ;
        RECT 260.400 627.600 262.200 639.600 ;
        RECT 275.400 633.600 276.300 653.700 ;
        RECT 281.700 649.200 282.600 656.400 ;
        RECT 296.400 655.200 298.200 662.400 ;
        RECT 301.500 656.400 303.300 663.000 ;
        RECT 313.800 656.400 315.600 662.400 ;
        RECT 296.400 654.300 300.600 655.200 ;
        RECT 296.100 649.200 297.900 651.000 ;
        RECT 299.400 649.200 300.600 654.300 ;
        RECT 314.400 654.300 315.600 656.400 ;
        RECT 316.800 657.300 318.600 662.400 ;
        RECT 319.800 658.200 321.600 663.000 ;
        RECT 322.800 657.300 324.600 662.400 ;
        RECT 334.800 659.400 336.600 662.400 ;
        RECT 337.800 659.400 339.600 663.000 ;
        RECT 316.800 655.950 324.600 657.300 ;
        RECT 314.400 653.250 318.150 654.300 ;
        RECT 302.100 649.200 303.900 651.000 ;
        RECT 277.950 647.100 280.050 649.200 ;
        RECT 280.950 647.100 283.050 649.200 ;
        RECT 295.950 647.100 298.050 649.200 ;
        RECT 298.950 647.100 301.050 649.200 ;
        RECT 301.950 647.100 304.050 649.200 ;
        RECT 314.100 649.050 315.900 650.850 ;
        RECT 316.950 649.050 318.150 653.250 ;
        RECT 330.000 651.450 334.050 652.050 ;
        RECT 320.100 649.050 321.900 650.850 ;
        RECT 329.550 649.950 334.050 651.450 ;
        RECT 278.100 645.300 279.900 647.100 ;
        RECT 281.700 639.600 282.600 647.100 ;
        RECT 272.400 627.000 274.200 633.600 ;
        RECT 275.400 627.600 277.200 633.600 ;
        RECT 278.400 627.000 280.200 633.600 ;
        RECT 281.400 627.600 283.200 639.600 ;
        RECT 299.400 633.600 300.600 647.100 ;
        RECT 313.950 646.950 316.050 649.050 ;
        RECT 316.950 646.950 319.050 649.050 ;
        RECT 319.950 646.950 322.050 649.050 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 317.850 633.600 319.050 646.950 ;
        RECT 323.100 645.150 324.900 646.950 ;
        RECT 329.550 646.050 330.450 649.950 ;
        RECT 335.400 649.050 336.600 659.400 ;
        RECT 347.700 656.400 349.500 663.000 ;
        RECT 352.800 655.200 354.600 662.400 ;
        RECT 365.400 657.300 367.200 662.400 ;
        RECT 368.400 658.200 370.200 663.000 ;
        RECT 371.400 657.300 373.200 662.400 ;
        RECT 365.400 655.950 373.200 657.300 ;
        RECT 374.400 656.400 376.200 662.400 ;
        RECT 388.800 656.400 390.600 662.400 ;
        RECT 391.800 656.400 393.600 663.000 ;
        RECT 403.800 656.400 405.600 662.400 ;
        RECT 350.400 654.300 354.600 655.200 ;
        RECT 374.400 654.300 375.600 656.400 ;
        RECT 347.100 649.200 348.900 651.000 ;
        RECT 350.400 649.200 351.600 654.300 ;
        RECT 371.850 653.250 375.600 654.300 ;
        RECT 360.000 651.450 364.050 652.050 ;
        RECT 353.100 649.200 354.900 651.000 ;
        RECT 359.550 649.950 364.050 651.450 ;
        RECT 334.950 646.950 337.050 649.050 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 346.950 647.100 349.050 649.200 ;
        RECT 349.950 647.100 352.050 649.200 ;
        RECT 352.950 647.100 355.050 649.200 ;
        RECT 329.550 644.550 334.050 646.050 ;
        RECT 330.000 643.950 334.050 644.550 ;
        RECT 295.800 627.000 297.600 633.600 ;
        RECT 298.800 627.600 300.600 633.600 ;
        RECT 301.800 627.000 303.600 633.600 ;
        RECT 314.400 627.000 316.200 633.600 ;
        RECT 317.400 627.600 319.200 633.600 ;
        RECT 322.500 627.000 324.300 639.600 ;
        RECT 335.400 633.600 336.600 646.950 ;
        RECT 338.100 645.150 339.900 646.950 ;
        RECT 350.400 633.600 351.600 647.100 ;
        RECT 359.550 646.050 360.450 649.950 ;
        RECT 368.100 649.050 369.900 650.850 ;
        RECT 371.850 649.050 373.050 653.250 ;
        RECT 374.100 649.050 375.900 650.850 ;
        RECT 389.400 649.200 390.600 656.400 ;
        RECT 404.400 654.300 405.600 656.400 ;
        RECT 406.800 657.300 408.600 662.400 ;
        RECT 409.800 658.200 411.600 663.000 ;
        RECT 412.800 657.300 414.600 662.400 ;
        RECT 406.800 655.950 414.600 657.300 ;
        RECT 422.400 656.400 424.200 663.000 ;
        RECT 425.400 656.400 427.200 662.400 ;
        RECT 404.400 653.250 408.150 654.300 ;
        RECT 392.100 649.200 393.900 651.000 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 367.950 646.950 370.050 649.050 ;
        RECT 370.950 646.950 373.050 649.050 ;
        RECT 373.950 646.950 376.050 649.050 ;
        RECT 388.950 647.100 391.050 649.200 ;
        RECT 391.950 647.100 394.050 649.200 ;
        RECT 404.100 649.050 405.900 650.850 ;
        RECT 406.950 649.050 408.150 653.250 ;
        RECT 410.100 649.050 411.900 650.850 ;
        RECT 422.100 649.200 423.900 651.000 ;
        RECT 425.400 649.200 426.600 656.400 ;
        RECT 437.400 654.600 439.200 662.400 ;
        RECT 441.900 656.400 443.700 663.000 ;
        RECT 444.900 658.200 446.700 662.400 ;
        RECT 444.900 656.400 447.600 658.200 ;
        RECT 443.100 654.600 444.900 655.500 ;
        RECT 437.400 653.700 444.900 654.600 ;
        RECT 437.100 649.200 438.900 651.000 ;
        RECT 355.950 644.550 360.450 646.050 ;
        RECT 365.100 645.150 366.900 646.950 ;
        RECT 355.950 643.950 360.000 644.550 ;
        RECT 334.800 627.600 336.600 633.600 ;
        RECT 337.800 627.000 339.600 633.600 ;
        RECT 347.400 627.000 349.200 633.600 ;
        RECT 350.400 627.600 352.200 633.600 ;
        RECT 353.400 627.000 355.200 633.600 ;
        RECT 365.700 627.000 367.500 639.600 ;
        RECT 370.950 633.600 372.150 646.950 ;
        RECT 389.400 639.600 390.600 647.100 ;
        RECT 403.950 646.950 406.050 649.050 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 421.950 647.100 424.050 649.200 ;
        RECT 424.950 647.100 427.050 649.200 ;
        RECT 436.950 647.100 439.050 649.200 ;
        RECT 370.800 627.600 372.600 633.600 ;
        RECT 373.800 627.000 375.600 633.600 ;
        RECT 388.800 627.600 390.600 639.600 ;
        RECT 391.800 627.000 393.600 639.600 ;
        RECT 407.850 633.600 409.050 646.950 ;
        RECT 413.100 645.150 414.900 646.950 ;
        RECT 425.400 639.600 426.600 647.100 ;
        RECT 404.400 627.000 406.200 633.600 ;
        RECT 407.400 627.600 409.200 633.600 ;
        RECT 412.500 627.000 414.300 639.600 ;
        RECT 422.400 627.000 424.200 639.600 ;
        RECT 425.400 627.600 427.200 639.600 ;
        RECT 440.400 633.600 441.300 653.700 ;
        RECT 446.700 649.200 447.600 656.400 ;
        RECT 461.400 655.200 463.200 662.400 ;
        RECT 466.500 656.400 468.300 663.000 ;
        RECT 461.400 654.300 465.600 655.200 ;
        RECT 461.100 649.200 462.900 651.000 ;
        RECT 464.400 649.200 465.600 654.300 ;
        RECT 481.200 654.000 483.000 662.400 ;
        RECT 479.700 652.800 483.000 654.000 ;
        RECT 487.800 653.400 489.600 663.000 ;
        RECT 497.400 657.300 499.200 662.400 ;
        RECT 500.400 658.200 502.200 663.000 ;
        RECT 503.400 657.300 505.200 662.400 ;
        RECT 497.400 655.950 505.200 657.300 ;
        RECT 506.400 656.400 508.200 662.400 ;
        RECT 518.700 656.400 520.500 663.000 ;
        RECT 506.400 654.300 507.600 656.400 ;
        RECT 523.800 655.200 525.600 662.400 ;
        RECT 503.850 653.250 507.600 654.300 ;
        RECT 521.400 654.300 525.600 655.200 ;
        RECT 536.400 654.600 538.200 662.400 ;
        RECT 540.900 656.400 542.700 663.000 ;
        RECT 543.900 658.200 545.700 662.400 ;
        RECT 543.900 656.400 546.600 658.200 ;
        RECT 557.700 656.400 559.500 663.000 ;
        RECT 562.200 656.400 564.000 662.400 ;
        RECT 566.700 656.400 568.500 663.000 ;
        RECT 542.100 654.600 543.900 655.500 ;
        RECT 467.100 649.200 468.900 651.000 ;
        RECT 479.700 649.200 480.600 652.800 ;
        RECT 482.100 649.200 483.900 651.000 ;
        RECT 488.100 649.200 489.900 651.000 ;
        RECT 442.950 647.100 445.050 649.200 ;
        RECT 445.950 647.100 448.050 649.200 ;
        RECT 460.950 647.100 463.050 649.200 ;
        RECT 463.950 647.100 466.050 649.200 ;
        RECT 466.950 647.100 469.050 649.200 ;
        RECT 478.950 647.100 481.050 649.200 ;
        RECT 481.950 647.100 484.050 649.200 ;
        RECT 484.950 647.100 487.050 649.200 ;
        RECT 487.950 647.100 490.050 649.200 ;
        RECT 500.100 649.050 501.900 650.850 ;
        RECT 503.850 649.050 505.050 653.250 ;
        RECT 506.100 649.050 507.900 650.850 ;
        RECT 518.100 649.200 519.900 651.000 ;
        RECT 521.400 649.200 522.600 654.300 ;
        RECT 536.400 653.700 543.900 654.600 ;
        RECT 524.100 649.200 525.900 651.000 ;
        RECT 536.100 649.200 537.900 651.000 ;
        RECT 443.100 645.300 444.900 647.100 ;
        RECT 446.700 639.600 447.600 647.100 ;
        RECT 437.400 627.000 439.200 633.600 ;
        RECT 440.400 627.600 442.200 633.600 ;
        RECT 443.400 627.000 445.200 633.600 ;
        RECT 446.400 627.600 448.200 639.600 ;
        RECT 464.400 633.600 465.600 647.100 ;
        RECT 479.700 634.800 480.600 647.100 ;
        RECT 485.100 645.300 486.900 647.100 ;
        RECT 496.950 646.950 499.050 649.050 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 517.950 647.100 520.050 649.200 ;
        RECT 520.950 647.100 523.050 649.200 ;
        RECT 523.950 647.100 526.050 649.200 ;
        RECT 535.950 647.100 538.050 649.200 ;
        RECT 497.100 645.150 498.900 646.950 ;
        RECT 479.700 633.900 486.300 634.800 ;
        RECT 479.700 633.600 480.600 633.900 ;
        RECT 460.800 627.000 462.600 633.600 ;
        RECT 463.800 627.600 465.600 633.600 ;
        RECT 466.800 627.000 468.600 633.600 ;
        RECT 478.800 627.600 480.600 633.600 ;
        RECT 484.800 633.600 486.300 633.900 ;
        RECT 481.800 627.000 483.600 633.000 ;
        RECT 484.800 627.600 486.600 633.600 ;
        RECT 487.800 627.000 489.600 633.600 ;
        RECT 497.700 627.000 499.500 639.600 ;
        RECT 502.950 633.600 504.150 646.950 ;
        RECT 521.400 633.600 522.600 647.100 ;
        RECT 535.950 645.450 538.050 646.050 ;
        RECT 527.550 645.000 538.050 645.450 ;
        RECT 526.950 644.550 538.050 645.000 ;
        RECT 526.950 640.950 529.050 644.550 ;
        RECT 535.950 643.950 538.050 644.550 ;
        RECT 539.400 633.600 540.300 653.700 ;
        RECT 545.700 649.200 546.600 656.400 ;
        RECT 557.100 649.200 558.900 651.000 ;
        RECT 562.950 649.200 564.000 656.400 ;
        RECT 581.400 654.600 583.200 662.400 ;
        RECT 585.900 656.400 587.700 663.000 ;
        RECT 588.900 658.200 590.700 662.400 ;
        RECT 588.900 656.400 591.600 658.200 ;
        RECT 603.000 656.400 604.800 663.000 ;
        RECT 607.500 657.600 609.300 662.400 ;
        RECT 610.500 659.400 612.300 663.000 ;
        RECT 607.500 656.400 612.600 657.600 ;
        RECT 623.700 656.400 625.500 663.000 ;
        RECT 628.200 656.400 630.000 662.400 ;
        RECT 632.700 656.400 634.500 663.000 ;
        RECT 649.800 659.400 651.600 663.000 ;
        RECT 652.800 659.400 654.600 662.400 ;
        RECT 655.800 659.400 657.600 663.000 ;
        RECT 587.100 654.600 588.900 655.500 ;
        RECT 581.400 653.700 588.900 654.600 ;
        RECT 571.950 651.450 576.000 652.050 ;
        RECT 569.100 649.200 570.900 651.000 ;
        RECT 571.950 649.950 576.450 651.450 ;
        RECT 541.950 647.100 544.050 649.200 ;
        RECT 544.950 647.100 547.050 649.200 ;
        RECT 556.950 647.100 559.050 649.200 ;
        RECT 559.950 647.100 562.050 649.200 ;
        RECT 562.950 647.100 565.050 649.200 ;
        RECT 565.950 647.100 568.050 649.200 ;
        RECT 568.950 647.100 571.050 649.200 ;
        RECT 542.100 645.300 543.900 647.100 ;
        RECT 545.700 639.600 546.600 647.100 ;
        RECT 560.100 645.300 561.900 647.100 ;
        RECT 563.100 641.400 564.000 647.100 ;
        RECT 566.100 645.300 567.900 647.100 ;
        RECT 568.950 645.450 571.050 646.050 ;
        RECT 575.550 645.450 576.450 649.950 ;
        RECT 581.100 649.200 582.900 651.000 ;
        RECT 580.950 647.100 583.050 649.200 ;
        RECT 580.950 645.450 583.050 646.050 ;
        RECT 568.950 644.550 583.050 645.450 ;
        RECT 568.950 643.950 571.050 644.550 ;
        RECT 580.950 643.950 583.050 644.550 ;
        RECT 563.100 640.500 568.200 641.400 ;
        RECT 502.800 627.600 504.600 633.600 ;
        RECT 505.800 627.000 507.600 633.600 ;
        RECT 518.400 627.000 520.200 633.600 ;
        RECT 521.400 627.600 523.200 633.600 ;
        RECT 524.400 627.000 526.200 633.600 ;
        RECT 536.400 627.000 538.200 633.600 ;
        RECT 539.400 627.600 541.200 633.600 ;
        RECT 542.400 627.000 544.200 633.600 ;
        RECT 545.400 627.600 547.200 639.600 ;
        RECT 557.400 638.400 565.200 639.300 ;
        RECT 557.400 627.600 559.200 638.400 ;
        RECT 560.400 627.000 562.200 637.500 ;
        RECT 563.400 628.500 565.200 638.400 ;
        RECT 566.400 629.400 568.200 640.500 ;
        RECT 569.400 628.500 571.200 639.600 ;
        RECT 584.400 633.600 585.300 653.700 ;
        RECT 590.700 649.200 591.600 656.400 ;
        RECT 604.950 654.450 607.050 655.050 ;
        RECT 599.550 653.550 607.050 654.450 ;
        RECT 599.550 651.450 600.450 653.550 ;
        RECT 604.950 652.950 607.050 653.550 ;
        RECT 596.550 650.550 600.450 651.450 ;
        RECT 586.950 647.100 589.050 649.200 ;
        RECT 589.950 647.100 592.050 649.200 ;
        RECT 587.100 645.300 588.900 647.100 ;
        RECT 590.700 639.600 591.600 647.100 ;
        RECT 596.550 646.050 597.450 650.550 ;
        RECT 602.100 649.200 603.900 651.000 ;
        RECT 608.100 649.200 609.900 651.000 ;
        RECT 611.700 649.200 612.600 656.400 ;
        RECT 615.000 654.450 619.050 655.050 ;
        RECT 622.950 654.450 625.050 655.050 ;
        RECT 614.550 653.550 625.050 654.450 ;
        RECT 615.000 652.950 619.050 653.550 ;
        RECT 622.950 652.950 625.050 653.550 ;
        RECT 623.100 649.200 624.900 651.000 ;
        RECT 628.950 649.200 630.000 656.400 ;
        RECT 635.100 649.200 636.900 651.000 ;
        RECT 601.950 647.100 604.050 649.200 ;
        RECT 604.950 647.100 607.050 649.200 ;
        RECT 607.950 647.100 610.050 649.200 ;
        RECT 610.950 647.100 613.050 649.200 ;
        RECT 622.950 647.100 625.050 649.200 ;
        RECT 625.950 647.100 628.050 649.200 ;
        RECT 628.950 647.100 631.050 649.200 ;
        RECT 631.950 647.100 634.050 649.200 ;
        RECT 634.950 647.100 637.050 649.200 ;
        RECT 653.400 649.050 654.300 659.400 ;
        RECT 668.400 655.200 670.200 662.400 ;
        RECT 673.500 656.400 675.300 663.000 ;
        RECT 668.400 654.300 672.600 655.200 ;
        RECT 668.100 649.200 669.900 651.000 ;
        RECT 671.400 649.200 672.600 654.300 ;
        RECT 683.400 653.400 685.200 663.000 ;
        RECT 690.000 654.000 691.800 662.400 ;
        RECT 705.000 656.400 706.800 663.000 ;
        RECT 709.500 657.600 711.300 662.400 ;
        RECT 712.500 659.400 714.300 663.000 ;
        RECT 727.800 659.400 729.600 662.400 ;
        RECT 730.800 659.400 732.600 663.000 ;
        RECT 709.500 656.400 714.600 657.600 ;
        RECT 690.000 652.800 693.300 654.000 ;
        RECT 674.100 649.200 675.900 651.000 ;
        RECT 683.100 649.200 684.900 651.000 ;
        RECT 689.100 649.200 690.900 651.000 ;
        RECT 692.400 649.200 693.300 652.800 ;
        RECT 704.100 649.200 705.900 651.000 ;
        RECT 710.100 649.200 711.900 651.000 ;
        RECT 713.700 649.200 714.600 656.400 ;
        RECT 592.950 644.550 597.450 646.050 ;
        RECT 605.100 645.300 606.900 647.100 ;
        RECT 592.950 643.950 597.000 644.550 ;
        RECT 611.700 639.600 612.600 647.100 ;
        RECT 613.950 645.450 616.050 646.050 ;
        RECT 622.950 645.450 625.050 646.050 ;
        RECT 613.950 644.550 625.050 645.450 ;
        RECT 626.100 645.300 627.900 647.100 ;
        RECT 613.950 643.950 616.050 644.550 ;
        RECT 622.950 643.950 625.050 644.550 ;
        RECT 629.100 641.400 630.000 647.100 ;
        RECT 632.100 645.300 633.900 647.100 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 652.950 646.950 655.050 649.050 ;
        RECT 655.950 646.950 658.050 649.050 ;
        RECT 667.950 647.100 670.050 649.200 ;
        RECT 670.950 647.100 673.050 649.200 ;
        RECT 673.950 647.100 676.050 649.200 ;
        RECT 682.950 647.100 685.050 649.200 ;
        RECT 685.950 647.100 688.050 649.200 ;
        RECT 688.950 647.100 691.050 649.200 ;
        RECT 691.950 647.100 694.050 649.200 ;
        RECT 703.950 647.100 706.050 649.200 ;
        RECT 706.950 647.100 709.050 649.200 ;
        RECT 709.950 647.100 712.050 649.200 ;
        RECT 712.950 647.100 715.050 649.200 ;
        RECT 728.400 649.050 729.600 659.400 ;
        RECT 740.400 653.400 742.200 663.000 ;
        RECT 747.000 654.000 748.800 662.400 ;
        RECT 747.000 652.800 750.300 654.000 ;
        RECT 761.400 653.400 763.200 663.000 ;
        RECT 768.000 654.000 769.800 662.400 ;
        RECT 782.700 656.400 784.500 663.000 ;
        RECT 787.800 655.200 789.600 662.400 ;
        RECT 785.400 654.300 789.600 655.200 ;
        RECT 803.400 655.200 805.200 662.400 ;
        RECT 808.500 656.400 810.300 663.000 ;
        RECT 803.400 654.300 807.600 655.200 ;
        RECT 768.000 652.800 771.300 654.000 ;
        RECT 740.100 649.200 741.900 651.000 ;
        RECT 746.100 649.200 747.900 651.000 ;
        RECT 749.400 649.200 750.300 652.800 ;
        RECT 751.950 651.450 756.000 652.050 ;
        RECT 751.950 649.950 756.450 651.450 ;
        RECT 634.950 645.450 637.050 646.050 ;
        RECT 640.950 645.450 643.050 646.050 ;
        RECT 634.950 644.550 643.050 645.450 ;
        RECT 650.100 645.150 651.900 646.950 ;
        RECT 634.950 643.950 637.050 644.550 ;
        RECT 640.950 643.950 643.050 644.550 ;
        RECT 629.100 640.500 634.200 641.400 ;
        RECT 563.400 627.600 571.200 628.500 ;
        RECT 581.400 627.000 583.200 633.600 ;
        RECT 584.400 627.600 586.200 633.600 ;
        RECT 587.400 627.000 589.200 633.600 ;
        RECT 590.400 627.600 592.200 639.600 ;
        RECT 602.400 638.700 610.200 639.600 ;
        RECT 602.400 627.600 604.200 638.700 ;
        RECT 605.400 627.000 607.200 637.800 ;
        RECT 608.400 627.600 610.200 638.700 ;
        RECT 611.400 627.600 613.200 639.600 ;
        RECT 623.400 638.400 631.200 639.300 ;
        RECT 623.400 627.600 625.200 638.400 ;
        RECT 626.400 627.000 628.200 637.500 ;
        RECT 629.400 628.500 631.200 638.400 ;
        RECT 632.400 629.400 634.200 640.500 ;
        RECT 653.400 639.600 654.300 646.950 ;
        RECT 656.100 645.150 657.900 646.950 ;
        RECT 635.400 628.500 637.200 639.600 ;
        RECT 629.400 627.600 637.200 628.500 ;
        RECT 650.700 638.400 654.300 639.600 ;
        RECT 650.700 627.600 652.500 638.400 ;
        RECT 655.800 627.000 657.600 639.600 ;
        RECT 671.400 633.600 672.600 647.100 ;
        RECT 673.950 645.450 676.050 646.050 ;
        RECT 682.950 645.450 685.050 646.050 ;
        RECT 673.950 644.550 685.050 645.450 ;
        RECT 686.100 645.300 687.900 647.100 ;
        RECT 673.950 643.950 676.050 644.550 ;
        RECT 682.950 643.950 685.050 644.550 ;
        RECT 692.400 634.800 693.300 647.100 ;
        RECT 707.100 645.300 708.900 647.100 ;
        RECT 713.700 639.600 714.600 647.100 ;
        RECT 727.950 646.950 730.050 649.050 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 739.950 647.100 742.050 649.200 ;
        RECT 742.950 647.100 745.050 649.200 ;
        RECT 745.950 647.100 748.050 649.200 ;
        RECT 748.950 647.100 751.050 649.200 ;
        RECT 686.700 633.900 693.300 634.800 ;
        RECT 686.700 633.600 688.200 633.900 ;
        RECT 667.800 627.000 669.600 633.600 ;
        RECT 670.800 627.600 672.600 633.600 ;
        RECT 673.800 627.000 675.600 633.600 ;
        RECT 683.400 627.000 685.200 633.600 ;
        RECT 686.400 627.600 688.200 633.600 ;
        RECT 692.400 633.600 693.300 633.900 ;
        RECT 704.400 638.700 712.200 639.600 ;
        RECT 689.400 627.000 691.200 633.000 ;
        RECT 692.400 627.600 694.200 633.600 ;
        RECT 704.400 627.600 706.200 638.700 ;
        RECT 707.400 627.000 709.200 637.800 ;
        RECT 710.400 627.600 712.200 638.700 ;
        RECT 713.400 627.600 715.200 639.600 ;
        RECT 728.400 633.600 729.600 646.950 ;
        RECT 731.100 645.150 732.900 646.950 ;
        RECT 743.100 645.300 744.900 647.100 ;
        RECT 749.400 634.800 750.300 647.100 ;
        RECT 755.550 645.450 756.450 649.950 ;
        RECT 761.100 649.200 762.900 651.000 ;
        RECT 767.100 649.200 768.900 651.000 ;
        RECT 770.400 649.200 771.300 652.800 ;
        RECT 772.950 651.450 777.000 652.050 ;
        RECT 772.950 649.950 777.450 651.450 ;
        RECT 760.950 647.100 763.050 649.200 ;
        RECT 763.950 647.100 766.050 649.200 ;
        RECT 766.950 647.100 769.050 649.200 ;
        RECT 769.950 647.100 772.050 649.200 ;
        RECT 752.550 645.000 756.450 645.450 ;
        RECT 764.100 645.300 765.900 647.100 ;
        RECT 751.950 644.550 756.450 645.000 ;
        RECT 751.950 640.950 754.050 644.550 ;
        RECT 757.950 642.450 760.050 643.050 ;
        RECT 766.950 642.450 769.050 643.050 ;
        RECT 757.950 641.550 769.050 642.450 ;
        RECT 757.950 640.950 760.050 641.550 ;
        RECT 766.950 640.950 769.050 641.550 ;
        RECT 770.400 634.800 771.300 647.100 ;
        RECT 776.550 645.450 777.450 649.950 ;
        RECT 782.100 649.200 783.900 651.000 ;
        RECT 785.400 649.200 786.600 654.300 ;
        RECT 788.100 649.200 789.900 651.000 ;
        RECT 803.100 649.200 804.900 651.000 ;
        RECT 806.400 649.200 807.600 654.300 ;
        RECT 818.400 653.400 820.200 663.000 ;
        RECT 825.000 654.000 826.800 662.400 ;
        RECT 825.000 652.800 828.300 654.000 ;
        RECT 839.400 653.400 841.200 663.000 ;
        RECT 846.000 654.000 847.800 662.400 ;
        RECT 846.000 652.800 849.300 654.000 ;
        RECT 809.100 649.200 810.900 651.000 ;
        RECT 818.100 649.200 819.900 651.000 ;
        RECT 824.100 649.200 825.900 651.000 ;
        RECT 827.400 649.200 828.300 652.800 ;
        RECT 839.100 649.200 840.900 651.000 ;
        RECT 845.100 649.200 846.900 651.000 ;
        RECT 848.400 649.200 849.300 652.800 ;
        RECT 781.950 647.100 784.050 649.200 ;
        RECT 784.950 647.100 787.050 649.200 ;
        RECT 787.950 647.100 790.050 649.200 ;
        RECT 802.950 647.100 805.050 649.200 ;
        RECT 805.950 647.100 808.050 649.200 ;
        RECT 808.950 647.100 811.050 649.200 ;
        RECT 817.950 647.100 820.050 649.200 ;
        RECT 820.950 647.100 823.050 649.200 ;
        RECT 823.950 647.100 826.050 649.200 ;
        RECT 826.950 647.100 829.050 649.200 ;
        RECT 838.950 647.100 841.050 649.200 ;
        RECT 841.950 647.100 844.050 649.200 ;
        RECT 844.950 647.100 847.050 649.200 ;
        RECT 847.950 647.100 850.050 649.200 ;
        RECT 781.950 645.450 784.050 646.050 ;
        RECT 776.550 644.550 784.050 645.450 ;
        RECT 781.950 643.950 784.050 644.550 ;
        RECT 743.700 633.900 750.300 634.800 ;
        RECT 743.700 633.600 745.200 633.900 ;
        RECT 727.800 627.600 729.600 633.600 ;
        RECT 730.800 627.000 732.600 633.600 ;
        RECT 740.400 627.000 742.200 633.600 ;
        RECT 743.400 627.600 745.200 633.600 ;
        RECT 749.400 633.600 750.300 633.900 ;
        RECT 764.700 633.900 771.300 634.800 ;
        RECT 764.700 633.600 766.200 633.900 ;
        RECT 746.400 627.000 748.200 633.000 ;
        RECT 749.400 627.600 751.200 633.600 ;
        RECT 761.400 627.000 763.200 633.600 ;
        RECT 764.400 627.600 766.200 633.600 ;
        RECT 770.400 633.600 771.300 633.900 ;
        RECT 785.400 633.600 786.600 647.100 ;
        RECT 793.950 639.450 796.050 640.050 ;
        RECT 799.950 639.450 802.050 640.050 ;
        RECT 793.950 638.550 802.050 639.450 ;
        RECT 793.950 637.950 796.050 638.550 ;
        RECT 799.950 637.950 802.050 638.550 ;
        RECT 787.950 636.450 790.050 636.900 ;
        RECT 796.950 636.450 799.050 637.050 ;
        RECT 802.950 636.450 805.050 637.050 ;
        RECT 787.950 635.550 805.050 636.450 ;
        RECT 787.950 634.800 790.050 635.550 ;
        RECT 796.950 634.950 799.050 635.550 ;
        RECT 802.950 634.950 805.050 635.550 ;
        RECT 806.400 633.600 807.600 647.100 ;
        RECT 821.100 645.300 822.900 647.100 ;
        RECT 827.400 634.800 828.300 647.100 ;
        RECT 842.100 645.300 843.900 647.100 ;
        RECT 848.400 634.800 849.300 647.100 ;
        RECT 821.700 633.900 828.300 634.800 ;
        RECT 821.700 633.600 823.200 633.900 ;
        RECT 767.400 627.000 769.200 633.000 ;
        RECT 770.400 627.600 772.200 633.600 ;
        RECT 782.400 627.000 784.200 633.600 ;
        RECT 785.400 627.600 787.200 633.600 ;
        RECT 788.400 627.000 790.200 633.600 ;
        RECT 802.800 627.000 804.600 633.600 ;
        RECT 805.800 627.600 807.600 633.600 ;
        RECT 808.800 627.000 810.600 633.600 ;
        RECT 818.400 627.000 820.200 633.600 ;
        RECT 821.400 627.600 823.200 633.600 ;
        RECT 827.400 633.600 828.300 633.900 ;
        RECT 842.700 633.900 849.300 634.800 ;
        RECT 842.700 633.600 844.200 633.900 ;
        RECT 824.400 627.000 826.200 633.000 ;
        RECT 827.400 627.600 829.200 633.600 ;
        RECT 839.400 627.000 841.200 633.600 ;
        RECT 842.400 627.600 844.200 633.600 ;
        RECT 848.400 633.600 849.300 633.900 ;
        RECT 845.400 627.000 847.200 633.000 ;
        RECT 848.400 627.600 850.200 633.600 ;
        RECT 10.800 617.400 12.600 623.400 ;
        RECT 13.800 618.000 15.600 624.000 ;
        RECT 11.700 617.100 12.600 617.400 ;
        RECT 16.800 617.400 18.600 623.400 ;
        RECT 19.800 617.400 21.600 624.000 ;
        RECT 16.800 617.100 18.300 617.400 ;
        RECT 11.700 616.200 18.300 617.100 ;
        RECT 11.700 603.900 12.600 616.200 ;
        RECT 29.400 612.300 31.200 623.400 ;
        RECT 32.400 613.200 34.200 624.000 ;
        RECT 35.400 612.300 37.200 623.400 ;
        RECT 29.400 611.400 37.200 612.300 ;
        RECT 38.400 611.400 40.200 623.400 ;
        RECT 52.800 617.400 54.600 623.400 ;
        RECT 55.800 618.000 57.600 624.000 ;
        RECT 53.700 617.100 54.600 617.400 ;
        RECT 58.800 617.400 60.600 623.400 ;
        RECT 61.800 617.400 63.600 624.000 ;
        RECT 71.400 617.400 73.200 624.000 ;
        RECT 74.400 617.400 76.200 623.400 ;
        RECT 77.400 618.000 79.200 624.000 ;
        RECT 58.800 617.100 60.300 617.400 ;
        RECT 53.700 616.200 60.300 617.100 ;
        RECT 74.700 617.100 76.200 617.400 ;
        RECT 80.400 617.400 82.200 623.400 ;
        RECT 92.400 617.400 94.200 624.000 ;
        RECT 95.400 617.400 97.200 623.400 ;
        RECT 98.400 618.000 100.200 624.000 ;
        RECT 80.400 617.100 81.300 617.400 ;
        RECT 74.700 616.200 81.300 617.100 ;
        RECT 95.700 617.100 97.200 617.400 ;
        RECT 101.400 617.400 103.200 623.400 ;
        RECT 116.400 617.400 118.200 624.000 ;
        RECT 119.400 617.400 121.200 623.400 ;
        RECT 101.400 617.100 102.300 617.400 ;
        RECT 95.700 616.200 102.300 617.100 ;
        RECT 13.950 609.450 16.050 610.050 ;
        RECT 34.950 609.450 37.050 610.050 ;
        RECT 13.950 608.550 37.050 609.450 ;
        RECT 13.950 607.950 16.050 608.550 ;
        RECT 34.950 607.950 37.050 608.550 ;
        RECT 17.100 603.900 18.900 605.700 ;
        RECT 32.100 603.900 33.900 605.700 ;
        RECT 38.700 603.900 39.600 611.400 ;
        RECT 53.700 603.900 54.600 616.200 ;
        RECT 59.100 603.900 60.900 605.700 ;
        RECT 74.100 603.900 75.900 605.700 ;
        RECT 80.400 603.900 81.300 616.200 ;
        RECT 85.950 612.450 88.050 613.050 ;
        RECT 94.950 612.450 97.050 613.050 ;
        RECT 85.950 611.550 97.050 612.450 ;
        RECT 85.950 610.950 88.050 611.550 ;
        RECT 94.950 610.950 97.050 611.550 ;
        RECT 97.950 609.450 100.050 610.050 ;
        RECT 92.550 608.550 100.050 609.450 ;
        RECT 92.550 606.450 93.450 608.550 ;
        RECT 97.950 607.950 100.050 608.550 ;
        RECT 86.550 605.550 93.450 606.450 ;
        RECT 10.950 601.800 13.050 603.900 ;
        RECT 13.950 601.800 16.050 603.900 ;
        RECT 16.950 601.800 19.050 603.900 ;
        RECT 19.950 601.800 22.050 603.900 ;
        RECT 28.950 601.800 31.050 603.900 ;
        RECT 31.950 601.800 34.050 603.900 ;
        RECT 34.950 601.800 37.050 603.900 ;
        RECT 37.950 601.800 40.050 603.900 ;
        RECT 52.950 601.800 55.050 603.900 ;
        RECT 55.950 601.800 58.050 603.900 ;
        RECT 58.950 601.800 61.050 603.900 ;
        RECT 61.950 601.800 64.050 603.900 ;
        RECT 70.950 601.800 73.050 603.900 ;
        RECT 73.950 601.800 76.050 603.900 ;
        RECT 76.950 601.800 79.050 603.900 ;
        RECT 79.950 601.800 82.050 603.900 ;
        RECT 11.700 598.200 12.600 601.800 ;
        RECT 14.100 600.000 15.900 601.800 ;
        RECT 20.100 600.000 21.900 601.800 ;
        RECT 29.100 600.000 30.900 601.800 ;
        RECT 35.100 600.000 36.900 601.800 ;
        RECT 11.700 597.000 15.000 598.200 ;
        RECT 13.200 588.600 15.000 597.000 ;
        RECT 19.800 588.000 21.600 597.600 ;
        RECT 38.700 594.600 39.600 601.800 ;
        RECT 53.700 598.200 54.600 601.800 ;
        RECT 56.100 600.000 57.900 601.800 ;
        RECT 62.100 600.000 63.900 601.800 ;
        RECT 71.100 600.000 72.900 601.800 ;
        RECT 77.100 600.000 78.900 601.800 ;
        RECT 80.400 598.200 81.300 601.800 ;
        RECT 86.550 601.050 87.450 605.550 ;
        RECT 95.100 603.900 96.900 605.700 ;
        RECT 101.400 603.900 102.300 616.200 ;
        RECT 111.000 606.450 115.050 607.050 ;
        RECT 110.550 604.950 115.050 606.450 ;
        RECT 91.950 601.800 94.050 603.900 ;
        RECT 94.950 601.800 97.050 603.900 ;
        RECT 97.950 601.800 100.050 603.900 ;
        RECT 100.950 601.800 103.050 603.900 ;
        RECT 82.950 599.550 87.450 601.050 ;
        RECT 92.100 600.000 93.900 601.800 ;
        RECT 98.100 600.000 99.900 601.800 ;
        RECT 82.950 598.950 87.000 599.550 ;
        RECT 101.400 598.200 102.300 601.800 ;
        RECT 110.550 600.900 111.450 604.950 ;
        RECT 119.850 604.050 121.050 617.400 ;
        RECT 124.500 611.400 126.300 624.000 ;
        RECT 134.700 611.400 136.500 624.000 ;
        RECT 139.800 617.400 141.600 623.400 ;
        RECT 142.800 617.400 144.600 624.000 ;
        RECT 157.800 617.400 159.600 623.400 ;
        RECT 160.800 618.000 162.600 624.000 ;
        RECT 125.100 604.050 126.900 605.850 ;
        RECT 134.100 604.050 135.900 605.850 ;
        RECT 139.950 604.050 141.150 617.400 ;
        RECT 158.700 617.100 159.600 617.400 ;
        RECT 163.800 617.400 165.600 623.400 ;
        RECT 166.800 617.400 168.600 624.000 ;
        RECT 178.800 617.400 180.600 624.000 ;
        RECT 181.800 617.400 183.600 623.400 ;
        RECT 184.800 617.400 186.600 624.000 ;
        RECT 194.400 617.400 196.200 624.000 ;
        RECT 197.400 617.400 199.200 623.400 ;
        RECT 163.800 617.100 165.300 617.400 ;
        RECT 158.700 616.200 165.300 617.100 ;
        RECT 142.950 609.450 145.050 610.200 ;
        RECT 151.950 609.450 154.050 610.050 ;
        RECT 142.950 608.550 154.050 609.450 ;
        RECT 142.950 608.100 145.050 608.550 ;
        RECT 151.950 607.950 154.050 608.550 ;
        RECT 115.950 601.950 118.050 604.050 ;
        RECT 118.950 601.950 121.050 604.050 ;
        RECT 121.950 601.950 124.050 604.050 ;
        RECT 124.950 601.950 127.050 604.050 ;
        RECT 133.950 601.950 136.050 604.050 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 158.700 603.900 159.600 616.200 ;
        RECT 164.100 603.900 165.900 605.700 ;
        RECT 182.400 603.900 183.600 617.400 ;
        RECT 194.100 604.050 195.900 605.850 ;
        RECT 197.400 604.050 198.600 617.400 ;
        RECT 209.400 612.300 211.200 623.400 ;
        RECT 212.400 613.200 214.200 624.000 ;
        RECT 215.400 612.300 217.200 623.400 ;
        RECT 209.400 611.400 217.200 612.300 ;
        RECT 218.400 611.400 220.200 623.400 ;
        RECT 230.400 617.400 232.200 624.000 ;
        RECT 233.400 617.400 235.200 623.400 ;
        RECT 247.800 617.400 249.600 623.400 ;
        RECT 250.800 618.000 252.600 624.000 ;
        RECT 109.950 598.800 112.050 600.900 ;
        RECT 116.100 600.150 117.900 601.950 ;
        RECT 53.700 597.000 57.000 598.200 ;
        RECT 30.000 588.000 31.800 594.600 ;
        RECT 34.500 593.400 39.600 594.600 ;
        RECT 34.500 588.600 36.300 593.400 ;
        RECT 37.500 588.000 39.300 591.600 ;
        RECT 55.200 588.600 57.000 597.000 ;
        RECT 61.800 588.000 63.600 597.600 ;
        RECT 71.400 588.000 73.200 597.600 ;
        RECT 78.000 597.000 81.300 598.200 ;
        RECT 78.000 588.600 79.800 597.000 ;
        RECT 92.400 588.000 94.200 597.600 ;
        RECT 99.000 597.000 102.300 598.200 ;
        RECT 118.950 597.750 120.150 601.950 ;
        RECT 122.100 600.150 123.900 601.950 ;
        RECT 137.100 600.150 138.900 601.950 ;
        RECT 99.000 588.600 100.800 597.000 ;
        RECT 116.400 596.700 120.150 597.750 ;
        RECT 140.850 597.750 142.050 601.950 ;
        RECT 143.100 600.150 144.900 601.950 ;
        RECT 157.950 601.800 160.050 603.900 ;
        RECT 160.950 601.800 163.050 603.900 ;
        RECT 163.950 601.800 166.050 603.900 ;
        RECT 166.950 601.800 169.050 603.900 ;
        RECT 178.950 601.800 181.050 603.900 ;
        RECT 181.950 601.800 184.050 603.900 ;
        RECT 184.950 601.800 187.050 603.900 ;
        RECT 193.950 601.950 196.050 604.050 ;
        RECT 196.950 601.950 199.050 604.050 ;
        RECT 212.100 603.900 213.900 605.700 ;
        RECT 218.700 603.900 219.600 611.400 ;
        RECT 230.100 604.050 231.900 605.850 ;
        RECT 233.400 604.050 234.600 617.400 ;
        RECT 248.700 617.100 249.600 617.400 ;
        RECT 253.800 617.400 255.600 623.400 ;
        RECT 256.800 617.400 258.600 624.000 ;
        RECT 269.400 617.400 271.200 624.000 ;
        RECT 272.400 617.400 274.200 623.400 ;
        RECT 253.800 617.100 255.300 617.400 ;
        RECT 248.700 616.200 255.300 617.100 ;
        RECT 158.700 598.200 159.600 601.800 ;
        RECT 161.100 600.000 162.900 601.800 ;
        RECT 167.100 600.000 168.900 601.800 ;
        RECT 179.100 600.000 180.900 601.800 ;
        RECT 140.850 596.700 144.600 597.750 ;
        RECT 158.700 597.000 162.000 598.200 ;
        RECT 116.400 594.600 117.600 596.700 ;
        RECT 115.800 588.600 117.600 594.600 ;
        RECT 118.800 593.700 126.600 595.050 ;
        RECT 118.800 588.600 120.600 593.700 ;
        RECT 121.800 588.000 123.600 592.800 ;
        RECT 124.800 588.600 126.600 593.700 ;
        RECT 134.400 593.700 142.200 595.050 ;
        RECT 134.400 588.600 136.200 593.700 ;
        RECT 137.400 588.000 139.200 592.800 ;
        RECT 140.400 588.600 142.200 593.700 ;
        RECT 143.400 594.600 144.600 596.700 ;
        RECT 143.400 588.600 145.200 594.600 ;
        RECT 160.200 588.600 162.000 597.000 ;
        RECT 166.800 588.000 168.600 597.600 ;
        RECT 182.400 596.700 183.600 601.800 ;
        RECT 185.100 600.000 186.900 601.800 ;
        RECT 179.400 595.800 183.600 596.700 ;
        RECT 179.400 588.600 181.200 595.800 ;
        RECT 184.500 588.000 186.300 594.600 ;
        RECT 197.400 591.600 198.600 601.950 ;
        RECT 208.950 601.800 211.050 603.900 ;
        RECT 211.950 601.800 214.050 603.900 ;
        RECT 214.950 601.800 217.050 603.900 ;
        RECT 217.950 601.800 220.050 603.900 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 232.950 601.950 235.050 604.050 ;
        RECT 248.700 603.900 249.600 616.200 ;
        RECT 254.100 603.900 255.900 605.700 ;
        RECT 272.850 604.050 274.050 617.400 ;
        RECT 277.500 611.400 279.300 624.000 ;
        RECT 287.400 612.300 289.200 623.400 ;
        RECT 290.400 613.200 292.200 624.000 ;
        RECT 293.400 612.300 295.200 623.400 ;
        RECT 287.400 611.400 295.200 612.300 ;
        RECT 296.400 611.400 298.200 623.400 ;
        RECT 311.400 617.400 313.200 624.000 ;
        RECT 314.400 617.400 316.200 623.400 ;
        RECT 277.950 609.450 280.050 610.050 ;
        RECT 292.950 609.450 295.050 610.050 ;
        RECT 277.950 608.550 295.050 609.450 ;
        RECT 277.950 607.950 280.050 608.550 ;
        RECT 292.950 607.950 295.050 608.550 ;
        RECT 278.100 604.050 279.900 605.850 ;
        RECT 209.100 600.000 210.900 601.800 ;
        RECT 215.100 600.000 216.900 601.800 ;
        RECT 218.700 594.600 219.600 601.800 ;
        RECT 194.400 588.000 196.200 591.600 ;
        RECT 197.400 588.600 199.200 591.600 ;
        RECT 210.000 588.000 211.800 594.600 ;
        RECT 214.500 593.400 219.600 594.600 ;
        RECT 214.500 588.600 216.300 593.400 ;
        RECT 233.400 591.600 234.600 601.950 ;
        RECT 247.950 601.800 250.050 603.900 ;
        RECT 250.950 601.800 253.050 603.900 ;
        RECT 253.950 601.800 256.050 603.900 ;
        RECT 256.950 601.800 259.050 603.900 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 274.950 601.950 277.050 604.050 ;
        RECT 277.950 601.950 280.050 604.050 ;
        RECT 290.100 603.900 291.900 605.700 ;
        RECT 296.700 603.900 297.600 611.400 ;
        RECT 306.000 606.450 310.050 607.050 ;
        RECT 305.550 604.950 310.050 606.450 ;
        RECT 248.700 598.200 249.600 601.800 ;
        RECT 251.100 600.000 252.900 601.800 ;
        RECT 257.100 600.000 258.900 601.800 ;
        RECT 269.100 600.150 270.900 601.950 ;
        RECT 248.700 597.000 252.000 598.200 ;
        RECT 271.950 597.750 273.150 601.950 ;
        RECT 275.100 600.150 276.900 601.950 ;
        RECT 286.950 601.800 289.050 603.900 ;
        RECT 289.950 601.800 292.050 603.900 ;
        RECT 292.950 601.800 295.050 603.900 ;
        RECT 295.950 601.800 298.050 603.900 ;
        RECT 287.100 600.000 288.900 601.800 ;
        RECT 293.100 600.000 294.900 601.800 ;
        RECT 217.500 588.000 219.300 591.600 ;
        RECT 230.400 588.000 232.200 591.600 ;
        RECT 233.400 588.600 235.200 591.600 ;
        RECT 250.200 588.600 252.000 597.000 ;
        RECT 256.800 588.000 258.600 597.600 ;
        RECT 269.400 596.700 273.150 597.750 ;
        RECT 269.400 594.600 270.600 596.700 ;
        RECT 268.800 588.600 270.600 594.600 ;
        RECT 271.800 593.700 279.600 595.050 ;
        RECT 296.700 594.600 297.600 601.800 ;
        RECT 305.550 601.050 306.450 604.950 ;
        RECT 314.850 604.050 316.050 617.400 ;
        RECT 319.500 611.400 321.300 624.000 ;
        RECT 331.800 617.400 333.600 623.400 ;
        RECT 334.800 618.000 336.600 624.000 ;
        RECT 332.700 617.100 333.600 617.400 ;
        RECT 337.800 617.400 339.600 623.400 ;
        RECT 340.800 617.400 342.600 624.000 ;
        RECT 353.400 617.400 355.200 624.000 ;
        RECT 356.400 617.400 358.200 623.400 ;
        RECT 337.800 617.100 339.300 617.400 ;
        RECT 332.700 616.200 339.300 617.100 ;
        RECT 327.000 606.450 331.050 607.050 ;
        RECT 320.100 604.050 321.900 605.850 ;
        RECT 326.550 604.950 331.050 606.450 ;
        RECT 310.950 601.950 313.050 604.050 ;
        RECT 313.950 601.950 316.050 604.050 ;
        RECT 316.950 601.950 319.050 604.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 305.550 599.550 310.050 601.050 ;
        RECT 311.100 600.150 312.900 601.950 ;
        RECT 306.000 598.950 310.050 599.550 ;
        RECT 313.950 597.750 315.150 601.950 ;
        RECT 317.100 600.150 318.900 601.950 ;
        RECT 326.550 601.050 327.450 604.950 ;
        RECT 332.700 603.900 333.600 616.200 ;
        RECT 338.100 603.900 339.900 605.700 ;
        RECT 356.850 604.050 358.050 617.400 ;
        RECT 361.500 611.400 363.300 624.000 ;
        RECT 373.800 617.400 375.600 623.400 ;
        RECT 376.800 618.000 378.600 624.000 ;
        RECT 374.700 617.100 375.600 617.400 ;
        RECT 379.800 617.400 381.600 623.400 ;
        RECT 382.800 617.400 384.600 624.000 ;
        RECT 395.400 617.400 397.200 624.000 ;
        RECT 398.400 617.400 400.200 623.400 ;
        RECT 379.800 617.100 381.300 617.400 ;
        RECT 374.700 616.200 381.300 617.100 ;
        RECT 369.000 606.450 373.050 607.050 ;
        RECT 362.100 604.050 363.900 605.850 ;
        RECT 368.550 604.950 373.050 606.450 ;
        RECT 331.950 601.800 334.050 603.900 ;
        RECT 334.950 601.800 337.050 603.900 ;
        RECT 337.950 601.800 340.050 603.900 ;
        RECT 340.950 601.800 343.050 603.900 ;
        RECT 352.950 601.950 355.050 604.050 ;
        RECT 355.950 601.950 358.050 604.050 ;
        RECT 358.950 601.950 361.050 604.050 ;
        RECT 361.950 601.950 364.050 604.050 ;
        RECT 326.550 599.550 331.050 601.050 ;
        RECT 327.000 598.950 331.050 599.550 ;
        RECT 311.400 596.700 315.150 597.750 ;
        RECT 332.700 598.200 333.600 601.800 ;
        RECT 335.100 600.000 336.900 601.800 ;
        RECT 341.100 600.000 342.900 601.800 ;
        RECT 353.100 600.150 354.900 601.950 ;
        RECT 332.700 597.000 336.000 598.200 ;
        RECT 355.950 597.750 357.150 601.950 ;
        RECT 359.100 600.150 360.900 601.950 ;
        RECT 368.550 598.050 369.450 604.950 ;
        RECT 374.700 603.900 375.600 616.200 ;
        RECT 385.950 606.450 388.050 607.050 ;
        RECT 391.950 606.450 394.050 607.050 ;
        RECT 380.100 603.900 381.900 605.700 ;
        RECT 385.950 605.550 394.050 606.450 ;
        RECT 385.950 604.950 388.050 605.550 ;
        RECT 391.950 604.950 394.050 605.550 ;
        RECT 398.850 604.050 400.050 617.400 ;
        RECT 403.500 611.400 405.300 624.000 ;
        RECT 413.400 617.400 415.200 624.000 ;
        RECT 416.400 617.400 418.200 623.400 ;
        RECT 419.400 617.400 421.200 624.000 ;
        RECT 404.100 604.050 405.900 605.850 ;
        RECT 373.950 601.800 376.050 603.900 ;
        RECT 376.950 601.800 379.050 603.900 ;
        RECT 379.950 601.800 382.050 603.900 ;
        RECT 382.950 601.800 385.050 603.900 ;
        RECT 394.950 601.950 397.050 604.050 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 400.950 601.950 403.050 604.050 ;
        RECT 403.950 601.950 406.050 604.050 ;
        RECT 416.400 603.900 417.600 617.400 ;
        RECT 433.800 611.400 435.600 623.400 ;
        RECT 436.800 617.400 438.600 624.000 ;
        RECT 439.800 617.400 441.600 623.400 ;
        RECT 442.800 617.400 444.600 624.000 ;
        RECT 455.400 617.400 457.200 624.000 ;
        RECT 458.400 617.400 460.200 623.400 ;
        RECT 434.400 603.900 435.300 611.400 ;
        RECT 437.100 603.900 438.900 605.700 ;
        RECT 374.700 598.200 375.600 601.800 ;
        RECT 377.100 600.000 378.900 601.800 ;
        RECT 383.100 600.000 384.900 601.800 ;
        RECT 395.100 600.150 396.900 601.950 ;
        RECT 311.400 594.600 312.600 596.700 ;
        RECT 271.800 588.600 273.600 593.700 ;
        RECT 274.800 588.000 276.600 592.800 ;
        RECT 277.800 588.600 279.600 593.700 ;
        RECT 288.000 588.000 289.800 594.600 ;
        RECT 292.500 593.400 297.600 594.600 ;
        RECT 292.500 588.600 294.300 593.400 ;
        RECT 295.500 588.000 297.300 591.600 ;
        RECT 310.800 588.600 312.600 594.600 ;
        RECT 313.800 593.700 321.600 595.050 ;
        RECT 313.800 588.600 315.600 593.700 ;
        RECT 316.800 588.000 318.600 592.800 ;
        RECT 319.800 588.600 321.600 593.700 ;
        RECT 334.200 588.600 336.000 597.000 ;
        RECT 340.800 588.000 342.600 597.600 ;
        RECT 353.400 596.700 357.150 597.750 ;
        RECT 353.400 594.600 354.600 596.700 ;
        RECT 367.950 595.950 370.050 598.050 ;
        RECT 374.700 597.000 378.000 598.200 ;
        RECT 397.950 597.750 399.150 601.950 ;
        RECT 401.100 600.150 402.900 601.950 ;
        RECT 412.950 601.800 415.050 603.900 ;
        RECT 415.950 601.800 418.050 603.900 ;
        RECT 418.950 601.800 421.050 603.900 ;
        RECT 433.950 601.800 436.050 603.900 ;
        RECT 436.950 601.800 439.050 603.900 ;
        RECT 413.100 600.000 414.900 601.800 ;
        RECT 352.800 588.600 354.600 594.600 ;
        RECT 355.800 593.700 363.600 595.050 ;
        RECT 355.800 588.600 357.600 593.700 ;
        RECT 358.800 588.000 360.600 592.800 ;
        RECT 361.800 588.600 363.600 593.700 ;
        RECT 376.200 588.600 378.000 597.000 ;
        RECT 382.800 588.000 384.600 597.600 ;
        RECT 395.400 596.700 399.150 597.750 ;
        RECT 416.400 596.700 417.600 601.800 ;
        RECT 419.100 600.000 420.900 601.800 ;
        RECT 395.400 594.600 396.600 596.700 ;
        RECT 416.400 595.800 420.600 596.700 ;
        RECT 394.800 588.600 396.600 594.600 ;
        RECT 397.800 593.700 405.600 595.050 ;
        RECT 397.800 588.600 399.600 593.700 ;
        RECT 400.800 588.000 402.600 592.800 ;
        RECT 403.800 588.600 405.600 593.700 ;
        RECT 413.700 588.000 415.500 594.600 ;
        RECT 418.800 588.600 420.600 595.800 ;
        RECT 434.400 594.600 435.300 601.800 ;
        RECT 440.700 597.300 441.600 617.400 ;
        RECT 445.950 609.450 448.050 610.050 ;
        RECT 454.950 609.450 457.050 610.050 ;
        RECT 445.950 608.550 457.050 609.450 ;
        RECT 445.950 607.950 448.050 608.550 ;
        RECT 454.950 607.950 457.050 608.550 ;
        RECT 458.850 604.050 460.050 617.400 ;
        RECT 463.500 611.400 465.300 624.000 ;
        RECT 475.800 617.400 477.600 624.000 ;
        RECT 478.800 617.400 480.600 623.400 ;
        RECT 481.800 617.400 483.600 624.000 ;
        RECT 493.800 617.400 495.600 624.000 ;
        RECT 496.800 617.400 498.600 623.400 ;
        RECT 499.800 617.400 501.600 624.000 ;
        RECT 512.400 617.400 514.200 624.000 ;
        RECT 515.400 617.400 517.200 623.400 ;
        RECT 471.000 606.450 475.050 607.050 ;
        RECT 464.100 604.050 465.900 605.850 ;
        RECT 470.550 604.950 475.050 606.450 ;
        RECT 442.950 601.800 445.050 603.900 ;
        RECT 454.950 601.950 457.050 604.050 ;
        RECT 457.950 601.950 460.050 604.050 ;
        RECT 460.950 601.950 463.050 604.050 ;
        RECT 463.950 601.950 466.050 604.050 ;
        RECT 443.100 600.000 444.900 601.800 ;
        RECT 455.100 600.150 456.900 601.950 ;
        RECT 457.950 597.750 459.150 601.950 ;
        RECT 461.100 600.150 462.900 601.950 ;
        RECT 470.550 601.050 471.450 604.950 ;
        RECT 479.400 603.900 480.600 617.400 ;
        RECT 493.950 606.450 496.050 607.050 ;
        RECT 488.550 605.550 496.050 606.450 ;
        RECT 475.950 601.800 478.050 603.900 ;
        RECT 478.950 601.800 481.050 603.900 ;
        RECT 481.950 601.800 484.050 603.900 ;
        RECT 470.550 599.550 475.050 601.050 ;
        RECT 476.100 600.000 477.900 601.800 ;
        RECT 471.000 598.950 475.050 599.550 ;
        RECT 437.100 596.400 444.600 597.300 ;
        RECT 437.100 595.500 438.900 596.400 ;
        RECT 434.400 592.800 437.100 594.600 ;
        RECT 435.300 588.600 437.100 592.800 ;
        RECT 438.300 588.000 440.100 594.600 ;
        RECT 442.800 588.600 444.600 596.400 ;
        RECT 455.400 596.700 459.150 597.750 ;
        RECT 479.400 596.700 480.600 601.800 ;
        RECT 482.100 600.000 483.900 601.800 ;
        RECT 488.550 601.050 489.450 605.550 ;
        RECT 493.950 604.950 496.050 605.550 ;
        RECT 497.400 603.900 498.600 617.400 ;
        RECT 508.950 610.950 511.050 613.050 ;
        RECT 499.950 609.450 502.050 610.050 ;
        RECT 505.950 609.450 508.050 610.050 ;
        RECT 499.950 608.550 508.050 609.450 ;
        RECT 499.950 607.950 502.050 608.550 ;
        RECT 505.950 607.950 508.050 608.550 ;
        RECT 509.550 606.450 510.450 610.950 ;
        RECT 506.550 605.550 510.450 606.450 ;
        RECT 493.950 601.800 496.050 603.900 ;
        RECT 496.950 601.800 499.050 603.900 ;
        RECT 499.950 601.800 502.050 603.900 ;
        RECT 488.550 599.550 493.050 601.050 ;
        RECT 494.100 600.000 495.900 601.800 ;
        RECT 489.000 598.950 493.050 599.550 ;
        RECT 497.400 596.700 498.600 601.800 ;
        RECT 500.100 600.000 501.900 601.800 ;
        RECT 506.550 601.050 507.450 605.550 ;
        RECT 515.850 604.050 517.050 617.400 ;
        RECT 520.500 611.400 522.300 624.000 ;
        RECT 530.700 611.400 532.500 624.000 ;
        RECT 535.800 617.400 537.600 623.400 ;
        RECT 538.800 617.400 540.600 624.000 ;
        RECT 521.100 604.050 522.900 605.850 ;
        RECT 530.100 604.050 531.900 605.850 ;
        RECT 535.950 604.050 537.150 617.400 ;
        RECT 551.400 611.400 553.200 624.000 ;
        RECT 556.500 612.600 558.300 623.400 ;
        RECT 554.700 611.400 558.300 612.600 ;
        RECT 569.400 611.400 571.200 624.000 ;
        RECT 572.400 611.400 574.200 623.400 ;
        RECT 584.400 611.400 586.200 624.000 ;
        RECT 587.400 611.400 589.200 623.400 ;
        RECT 601.800 617.400 603.600 624.000 ;
        RECT 604.800 617.400 606.600 623.400 ;
        RECT 607.800 617.400 609.600 624.000 ;
        RECT 617.400 617.400 619.200 624.000 ;
        RECT 620.400 617.400 622.200 623.400 ;
        RECT 623.400 617.400 625.200 624.000 ;
        RECT 538.950 609.450 541.050 610.050 ;
        RECT 544.950 609.450 547.050 609.900 ;
        RECT 538.950 608.550 547.050 609.450 ;
        RECT 538.950 607.950 541.050 608.550 ;
        RECT 544.950 607.800 547.050 608.550 ;
        RECT 551.100 604.050 552.900 605.850 ;
        RECT 554.700 604.050 555.600 611.400 ;
        RECT 556.950 609.450 559.050 610.050 ;
        RECT 568.950 609.450 571.050 610.050 ;
        RECT 556.950 608.550 571.050 609.450 ;
        RECT 556.950 607.950 559.050 608.550 ;
        RECT 568.950 607.950 571.050 608.550 ;
        RECT 557.100 604.050 558.900 605.850 ;
        RECT 511.950 601.950 514.050 604.050 ;
        RECT 514.950 601.950 517.050 604.050 ;
        RECT 517.950 601.950 520.050 604.050 ;
        RECT 520.950 601.950 523.050 604.050 ;
        RECT 529.950 601.950 532.050 604.050 ;
        RECT 532.950 601.950 535.050 604.050 ;
        RECT 535.950 601.950 538.050 604.050 ;
        RECT 538.950 601.950 541.050 604.050 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 553.950 601.950 556.050 604.050 ;
        RECT 556.950 601.950 559.050 604.050 ;
        RECT 572.400 603.900 573.600 611.400 ;
        RECT 579.000 606.450 583.050 607.050 ;
        RECT 578.550 604.950 583.050 606.450 ;
        RECT 502.950 599.550 507.450 601.050 ;
        RECT 512.100 600.150 513.900 601.950 ;
        RECT 502.950 598.950 507.000 599.550 ;
        RECT 514.950 597.750 516.150 601.950 ;
        RECT 518.100 600.150 519.900 601.950 ;
        RECT 533.100 600.150 534.900 601.950 ;
        RECT 455.400 594.600 456.600 596.700 ;
        RECT 476.400 595.800 480.600 596.700 ;
        RECT 494.400 595.800 498.600 596.700 ;
        RECT 512.400 596.700 516.150 597.750 ;
        RECT 536.850 597.750 538.050 601.950 ;
        RECT 539.100 600.150 540.900 601.950 ;
        RECT 536.850 596.700 540.600 597.750 ;
        RECT 454.800 588.600 456.600 594.600 ;
        RECT 457.800 593.700 465.600 595.050 ;
        RECT 457.800 588.600 459.600 593.700 ;
        RECT 460.800 588.000 462.600 592.800 ;
        RECT 463.800 588.600 465.600 593.700 ;
        RECT 476.400 588.600 478.200 595.800 ;
        RECT 481.500 588.000 483.300 594.600 ;
        RECT 494.400 588.600 496.200 595.800 ;
        RECT 512.400 594.600 513.600 596.700 ;
        RECT 499.500 588.000 501.300 594.600 ;
        RECT 511.800 588.600 513.600 594.600 ;
        RECT 514.800 593.700 522.600 595.050 ;
        RECT 514.800 588.600 516.600 593.700 ;
        RECT 517.800 588.000 519.600 592.800 ;
        RECT 520.800 588.600 522.600 593.700 ;
        RECT 530.400 593.700 538.200 595.050 ;
        RECT 530.400 588.600 532.200 593.700 ;
        RECT 533.400 588.000 535.200 592.800 ;
        RECT 536.400 588.600 538.200 593.700 ;
        RECT 539.400 594.600 540.600 596.700 ;
        RECT 539.400 588.600 541.200 594.600 ;
        RECT 554.700 591.600 555.600 601.950 ;
        RECT 568.950 601.800 571.050 603.900 ;
        RECT 571.950 601.800 574.050 603.900 ;
        RECT 569.100 600.000 570.900 601.800 ;
        RECT 572.400 594.600 573.600 601.800 ;
        RECT 578.550 601.050 579.450 604.950 ;
        RECT 587.400 603.900 588.600 611.400 ;
        RECT 605.400 603.900 606.600 617.400 ;
        RECT 607.950 609.450 610.050 610.050 ;
        RECT 616.950 609.450 619.050 610.050 ;
        RECT 607.950 608.550 619.050 609.450 ;
        RECT 607.950 607.950 610.050 608.550 ;
        RECT 616.950 607.950 619.050 608.550 ;
        RECT 620.400 603.900 621.600 617.400 ;
        RECT 635.700 611.400 637.500 624.000 ;
        RECT 640.800 617.400 642.600 623.400 ;
        RECT 643.800 617.400 645.600 624.000 ;
        RECT 659.400 617.400 661.200 624.000 ;
        RECT 662.400 617.400 664.200 623.400 ;
        RECT 635.100 604.050 636.900 605.850 ;
        RECT 640.950 604.050 642.150 617.400 ;
        RECT 646.950 606.450 651.000 607.050 ;
        RECT 654.000 606.450 658.050 607.050 ;
        RECT 646.950 604.950 651.450 606.450 ;
        RECT 583.950 601.800 586.050 603.900 ;
        RECT 586.950 601.800 589.050 603.900 ;
        RECT 601.950 601.800 604.050 603.900 ;
        RECT 604.950 601.800 607.050 603.900 ;
        RECT 607.950 601.800 610.050 603.900 ;
        RECT 616.950 601.800 619.050 603.900 ;
        RECT 619.950 601.800 622.050 603.900 ;
        RECT 622.950 601.800 625.050 603.900 ;
        RECT 634.950 601.950 637.050 604.050 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 574.950 599.550 579.450 601.050 ;
        RECT 584.100 600.000 585.900 601.800 ;
        RECT 574.950 598.950 579.000 599.550 ;
        RECT 587.400 594.600 588.600 601.800 ;
        RECT 602.100 600.000 603.900 601.800 ;
        RECT 605.400 596.700 606.600 601.800 ;
        RECT 608.100 600.000 609.900 601.800 ;
        RECT 617.100 600.000 618.900 601.800 ;
        RECT 602.400 595.800 606.600 596.700 ;
        RECT 620.400 596.700 621.600 601.800 ;
        RECT 623.100 600.000 624.900 601.800 ;
        RECT 638.100 600.150 639.900 601.950 ;
        RECT 641.850 597.750 643.050 601.950 ;
        RECT 644.100 600.150 645.900 601.950 ;
        RECT 650.550 601.050 651.450 604.950 ;
        RECT 646.950 599.550 651.450 601.050 ;
        RECT 653.550 604.950 658.050 606.450 ;
        RECT 653.550 601.050 654.450 604.950 ;
        RECT 662.850 604.050 664.050 617.400 ;
        RECT 667.500 611.400 669.300 624.000 ;
        RECT 677.700 611.400 679.500 624.000 ;
        RECT 682.800 617.400 684.600 623.400 ;
        RECT 685.800 617.400 687.600 624.000 ;
        RECT 668.100 604.050 669.900 605.850 ;
        RECT 677.100 604.050 678.900 605.850 ;
        RECT 682.950 604.050 684.150 617.400 ;
        RECT 698.400 612.300 700.200 623.400 ;
        RECT 701.400 613.200 703.200 624.000 ;
        RECT 704.400 612.300 706.200 623.400 ;
        RECT 698.400 611.400 706.200 612.300 ;
        RECT 707.400 611.400 709.200 623.400 ;
        RECT 719.400 617.400 721.200 624.000 ;
        RECT 722.400 617.400 724.200 623.400 ;
        RECT 725.400 618.000 727.200 624.000 ;
        RECT 722.700 617.100 724.200 617.400 ;
        RECT 728.400 617.400 730.200 623.400 ;
        RECT 740.400 617.400 742.200 624.000 ;
        RECT 743.400 617.400 745.200 623.400 ;
        RECT 755.400 617.400 757.200 624.000 ;
        RECT 758.400 617.400 760.200 623.400 ;
        RECT 761.400 618.000 763.200 624.000 ;
        RECT 728.400 617.100 729.300 617.400 ;
        RECT 722.700 616.200 729.300 617.100 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 676.950 601.950 679.050 604.050 ;
        RECT 679.950 601.950 682.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 701.100 603.900 702.900 605.700 ;
        RECT 707.700 603.900 708.600 611.400 ;
        RECT 722.100 603.900 723.900 605.700 ;
        RECT 728.400 603.900 729.300 616.200 ;
        RECT 740.100 604.050 741.900 605.850 ;
        RECT 743.400 604.050 744.600 617.400 ;
        RECT 758.700 617.100 760.200 617.400 ;
        RECT 764.400 617.400 766.200 623.400 ;
        RECT 778.800 617.400 780.600 624.000 ;
        RECT 781.800 617.400 783.600 623.400 ;
        RECT 784.800 617.400 786.600 624.000 ;
        RECT 796.800 617.400 798.600 624.000 ;
        RECT 799.800 617.400 801.600 623.400 ;
        RECT 802.800 617.400 804.600 624.000 ;
        RECT 812.400 617.400 814.200 623.400 ;
        RECT 815.400 617.400 817.200 624.000 ;
        RECT 764.400 617.100 765.300 617.400 ;
        RECT 758.700 616.200 765.300 617.100 ;
        RECT 748.950 606.450 751.050 607.050 ;
        RECT 754.950 606.450 757.050 607.050 ;
        RECT 748.950 605.550 757.050 606.450 ;
        RECT 748.950 604.950 751.050 605.550 ;
        RECT 754.950 604.950 757.050 605.550 ;
        RECT 653.550 599.550 658.050 601.050 ;
        RECT 659.100 600.150 660.900 601.950 ;
        RECT 646.950 598.950 651.000 599.550 ;
        RECT 654.000 598.950 658.050 599.550 ;
        RECT 661.950 597.750 663.150 601.950 ;
        RECT 665.100 600.150 666.900 601.950 ;
        RECT 680.100 600.150 681.900 601.950 ;
        RECT 641.850 596.700 645.600 597.750 ;
        RECT 620.400 595.800 624.600 596.700 ;
        RECT 551.400 588.000 553.200 591.600 ;
        RECT 554.400 588.600 556.200 591.600 ;
        RECT 557.400 588.000 559.200 591.600 ;
        RECT 569.400 588.000 571.200 594.600 ;
        RECT 572.400 588.600 574.200 594.600 ;
        RECT 584.400 588.000 586.200 594.600 ;
        RECT 587.400 588.600 589.200 594.600 ;
        RECT 602.400 588.600 604.200 595.800 ;
        RECT 607.500 588.000 609.300 594.600 ;
        RECT 617.700 588.000 619.500 594.600 ;
        RECT 622.800 588.600 624.600 595.800 ;
        RECT 635.400 593.700 643.200 595.050 ;
        RECT 635.400 588.600 637.200 593.700 ;
        RECT 638.400 588.000 640.200 592.800 ;
        RECT 641.400 588.600 643.200 593.700 ;
        RECT 644.400 594.600 645.600 596.700 ;
        RECT 659.400 596.700 663.150 597.750 ;
        RECT 683.850 597.750 685.050 601.950 ;
        RECT 686.100 600.150 687.900 601.950 ;
        RECT 697.950 601.800 700.050 603.900 ;
        RECT 700.950 601.800 703.050 603.900 ;
        RECT 703.950 601.800 706.050 603.900 ;
        RECT 706.950 601.800 709.050 603.900 ;
        RECT 718.950 601.800 721.050 603.900 ;
        RECT 721.950 601.800 724.050 603.900 ;
        RECT 724.950 601.800 727.050 603.900 ;
        RECT 727.950 601.800 730.050 603.900 ;
        RECT 739.950 601.950 742.050 604.050 ;
        RECT 742.950 601.950 745.050 604.050 ;
        RECT 758.100 603.900 759.900 605.700 ;
        RECT 764.400 603.900 765.300 616.200 ;
        RECT 782.400 603.900 783.600 617.400 ;
        RECT 784.950 606.450 787.050 607.050 ;
        RECT 784.950 605.550 792.450 606.450 ;
        RECT 784.950 604.950 787.050 605.550 ;
        RECT 698.100 600.000 699.900 601.800 ;
        RECT 704.100 600.000 705.900 601.800 ;
        RECT 683.850 596.700 687.600 597.750 ;
        RECT 659.400 594.600 660.600 596.700 ;
        RECT 644.400 588.600 646.200 594.600 ;
        RECT 658.800 588.600 660.600 594.600 ;
        RECT 661.800 593.700 669.600 595.050 ;
        RECT 661.800 588.600 663.600 593.700 ;
        RECT 664.800 588.000 666.600 592.800 ;
        RECT 667.800 588.600 669.600 593.700 ;
        RECT 677.400 593.700 685.200 595.050 ;
        RECT 677.400 588.600 679.200 593.700 ;
        RECT 680.400 588.000 682.200 592.800 ;
        RECT 683.400 588.600 685.200 593.700 ;
        RECT 686.400 594.600 687.600 596.700 ;
        RECT 688.950 597.450 691.050 598.050 ;
        RECT 694.950 597.450 697.050 598.050 ;
        RECT 688.950 596.550 697.050 597.450 ;
        RECT 688.950 595.950 691.050 596.550 ;
        RECT 694.950 595.950 697.050 596.550 ;
        RECT 707.700 594.600 708.600 601.800 ;
        RECT 719.100 600.000 720.900 601.800 ;
        RECT 725.100 600.000 726.900 601.800 ;
        RECT 728.400 598.200 729.300 601.800 ;
        RECT 686.400 588.600 688.200 594.600 ;
        RECT 699.000 588.000 700.800 594.600 ;
        RECT 703.500 593.400 708.600 594.600 ;
        RECT 703.500 588.600 705.300 593.400 ;
        RECT 706.500 588.000 708.300 591.600 ;
        RECT 719.400 588.000 721.200 597.600 ;
        RECT 726.000 597.000 729.300 598.200 ;
        RECT 726.000 588.600 727.800 597.000 ;
        RECT 743.400 591.600 744.600 601.950 ;
        RECT 754.950 601.800 757.050 603.900 ;
        RECT 757.950 601.800 760.050 603.900 ;
        RECT 760.950 601.800 763.050 603.900 ;
        RECT 763.950 601.800 766.050 603.900 ;
        RECT 778.950 601.800 781.050 603.900 ;
        RECT 781.950 601.800 784.050 603.900 ;
        RECT 784.950 601.800 787.050 603.900 ;
        RECT 755.100 600.000 756.900 601.800 ;
        RECT 761.100 600.000 762.900 601.800 ;
        RECT 764.400 598.200 765.300 601.800 ;
        RECT 779.100 600.000 780.900 601.800 ;
        RECT 740.400 588.000 742.200 591.600 ;
        RECT 743.400 588.600 745.200 591.600 ;
        RECT 755.400 588.000 757.200 597.600 ;
        RECT 762.000 597.000 765.300 598.200 ;
        RECT 762.000 588.600 763.800 597.000 ;
        RECT 782.400 596.700 783.600 601.800 ;
        RECT 785.100 600.000 786.900 601.800 ;
        RECT 791.550 601.050 792.450 605.550 ;
        RECT 800.400 603.900 801.600 617.400 ;
        RECT 812.400 610.500 813.600 617.400 ;
        RECT 818.400 611.400 820.200 623.400 ;
        RECT 830.400 611.400 832.200 624.000 ;
        RECT 835.500 612.600 837.300 623.400 ;
        RECT 833.700 611.400 837.300 612.600 ;
        RECT 848.400 617.400 850.200 623.400 ;
        RECT 851.400 617.400 853.200 624.000 ;
        RECT 812.400 609.600 818.100 610.500 ;
        RECT 816.150 608.700 818.100 609.600 ;
        RECT 812.100 604.050 813.900 605.850 ;
        RECT 796.950 601.800 799.050 603.900 ;
        RECT 799.950 601.800 802.050 603.900 ;
        RECT 802.950 601.800 805.050 603.900 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 791.550 599.550 796.050 601.050 ;
        RECT 797.100 600.000 798.900 601.800 ;
        RECT 792.000 598.950 796.050 599.550 ;
        RECT 800.400 596.700 801.600 601.800 ;
        RECT 803.100 600.000 804.900 601.800 ;
        RECT 779.400 595.800 783.600 596.700 ;
        RECT 797.400 595.800 801.600 596.700 ;
        RECT 816.150 597.300 817.050 608.700 ;
        RECT 819.000 604.050 820.200 611.400 ;
        RECT 830.100 604.050 831.900 605.850 ;
        RECT 833.700 604.050 834.600 611.400 ;
        RECT 848.400 610.500 849.600 617.400 ;
        RECT 854.400 611.400 856.200 623.400 ;
        RECT 848.400 609.600 854.100 610.500 ;
        RECT 852.150 608.700 854.100 609.600 ;
        RECT 836.100 604.050 837.900 605.850 ;
        RECT 848.100 604.050 849.900 605.850 ;
        RECT 817.950 601.950 820.200 604.050 ;
        RECT 829.950 601.950 832.050 604.050 ;
        RECT 832.950 601.950 835.050 604.050 ;
        RECT 835.950 601.950 838.050 604.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 816.150 596.400 818.100 597.300 ;
        RECT 779.400 588.600 781.200 595.800 ;
        RECT 784.500 588.000 786.300 594.600 ;
        RECT 797.400 588.600 799.200 595.800 ;
        RECT 812.400 595.500 818.100 596.400 ;
        RECT 802.500 588.000 804.300 594.600 ;
        RECT 812.400 591.600 813.600 595.500 ;
        RECT 819.000 594.600 820.200 601.950 ;
        RECT 812.400 588.600 814.200 591.600 ;
        RECT 815.400 588.000 817.200 591.600 ;
        RECT 818.400 588.600 820.200 594.600 ;
        RECT 833.700 591.600 834.600 601.950 ;
        RECT 852.150 597.300 853.050 608.700 ;
        RECT 855.000 604.050 856.200 611.400 ;
        RECT 853.950 601.950 856.200 604.050 ;
        RECT 852.150 596.400 854.100 597.300 ;
        RECT 848.400 595.500 854.100 596.400 ;
        RECT 848.400 591.600 849.600 595.500 ;
        RECT 855.000 594.600 856.200 601.950 ;
        RECT 830.400 588.000 832.200 591.600 ;
        RECT 833.400 588.600 835.200 591.600 ;
        RECT 836.400 588.000 838.200 591.600 ;
        RECT 848.400 588.600 850.200 591.600 ;
        RECT 851.400 588.000 853.200 591.600 ;
        RECT 854.400 588.600 856.200 594.600 ;
        RECT 10.800 581.400 12.600 584.400 ;
        RECT 13.800 581.400 15.600 585.000 ;
        RECT 11.400 571.050 12.600 581.400 ;
        RECT 24.000 578.400 25.800 585.000 ;
        RECT 28.500 579.600 30.300 584.400 ;
        RECT 31.500 581.400 33.300 585.000 ;
        RECT 28.500 578.400 33.600 579.600 ;
        RECT 46.800 578.400 48.600 584.400 ;
        RECT 23.100 571.200 24.900 573.000 ;
        RECT 29.100 571.200 30.900 573.000 ;
        RECT 32.700 571.200 33.600 578.400 ;
        RECT 47.400 576.300 48.600 578.400 ;
        RECT 49.800 579.300 51.600 584.400 ;
        RECT 52.800 580.200 54.600 585.000 ;
        RECT 55.800 579.300 57.600 584.400 ;
        RECT 68.700 581.400 70.500 585.000 ;
        RECT 71.700 579.600 73.500 584.400 ;
        RECT 49.800 577.950 57.600 579.300 ;
        RECT 68.400 578.400 73.500 579.600 ;
        RECT 76.200 578.400 78.000 585.000 ;
        RECT 47.400 575.250 51.150 576.300 ;
        RECT 10.950 568.950 13.050 571.050 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 22.950 569.100 25.050 571.200 ;
        RECT 25.950 569.100 28.050 571.200 ;
        RECT 28.950 569.100 31.050 571.200 ;
        RECT 31.950 569.100 34.050 571.200 ;
        RECT 47.100 571.050 48.900 572.850 ;
        RECT 49.950 571.050 51.150 575.250 ;
        RECT 53.100 571.050 54.900 572.850 ;
        RECT 68.400 571.200 69.300 578.400 ;
        RECT 86.400 575.400 88.200 585.000 ;
        RECT 93.000 576.000 94.800 584.400 ;
        RECT 107.400 579.300 109.200 584.400 ;
        RECT 110.400 580.200 112.200 585.000 ;
        RECT 113.400 579.300 115.200 584.400 ;
        RECT 107.400 577.950 115.200 579.300 ;
        RECT 116.400 578.400 118.200 584.400 ;
        RECT 116.400 576.300 117.600 578.400 ;
        RECT 93.000 574.800 96.300 576.000 ;
        RECT 71.100 571.200 72.900 573.000 ;
        RECT 77.100 571.200 78.900 573.000 ;
        RECT 86.100 571.200 87.900 573.000 ;
        RECT 92.100 571.200 93.900 573.000 ;
        RECT 95.400 571.200 96.300 574.800 ;
        RECT 113.850 575.250 117.600 576.300 ;
        RECT 128.400 575.400 130.200 585.000 ;
        RECT 135.000 576.000 136.800 584.400 ;
        RECT 150.000 578.400 151.800 585.000 ;
        RECT 154.500 579.600 156.300 584.400 ;
        RECT 157.500 581.400 159.300 585.000 ;
        RECT 154.500 578.400 159.600 579.600 ;
        RECT 142.950 576.450 145.050 577.050 ;
        RECT 154.950 576.450 157.050 577.050 ;
        RECT 97.950 573.450 102.000 574.050 ;
        RECT 97.950 571.950 102.450 573.450 ;
        RECT 11.400 555.600 12.600 568.950 ;
        RECT 14.100 567.150 15.900 568.950 ;
        RECT 26.100 567.300 27.900 569.100 ;
        RECT 32.700 561.600 33.600 569.100 ;
        RECT 46.950 568.950 49.050 571.050 ;
        RECT 49.950 568.950 52.050 571.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 55.950 568.950 58.050 571.050 ;
        RECT 67.950 569.100 70.050 571.200 ;
        RECT 70.950 569.100 73.050 571.200 ;
        RECT 73.950 569.100 76.050 571.200 ;
        RECT 76.950 569.100 79.050 571.200 ;
        RECT 85.950 569.100 88.050 571.200 ;
        RECT 88.950 569.100 91.050 571.200 ;
        RECT 91.950 569.100 94.050 571.200 ;
        RECT 94.950 569.100 97.050 571.200 ;
        RECT 23.400 560.700 31.200 561.600 ;
        RECT 10.800 549.600 12.600 555.600 ;
        RECT 13.800 549.000 15.600 555.600 ;
        RECT 23.400 549.600 25.200 560.700 ;
        RECT 26.400 549.000 28.200 559.800 ;
        RECT 29.400 549.600 31.200 560.700 ;
        RECT 32.400 549.600 34.200 561.600 ;
        RECT 50.850 555.600 52.050 568.950 ;
        RECT 56.100 567.150 57.900 568.950 ;
        RECT 68.400 561.600 69.300 569.100 ;
        RECT 74.100 567.300 75.900 569.100 ;
        RECT 89.100 567.300 90.900 569.100 ;
        RECT 47.400 549.000 49.200 555.600 ;
        RECT 50.400 549.600 52.200 555.600 ;
        RECT 55.500 549.000 57.300 561.600 ;
        RECT 67.800 549.600 69.600 561.600 ;
        RECT 70.800 560.700 78.600 561.600 ;
        RECT 70.800 549.600 72.600 560.700 ;
        RECT 73.800 549.000 75.600 559.800 ;
        RECT 76.800 549.600 78.600 560.700 ;
        RECT 95.400 556.800 96.300 569.100 ;
        RECT 101.550 568.050 102.450 571.950 ;
        RECT 110.100 571.050 111.900 572.850 ;
        RECT 113.850 571.050 115.050 575.250 ;
        RECT 135.000 574.800 138.300 576.000 ;
        RECT 142.950 575.550 157.050 576.450 ;
        RECT 142.950 574.950 145.050 575.550 ;
        RECT 154.950 574.950 157.050 575.550 ;
        RECT 123.000 573.450 127.050 574.050 ;
        RECT 116.100 571.050 117.900 572.850 ;
        RECT 122.550 571.950 127.050 573.450 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 112.950 568.950 115.050 571.050 ;
        RECT 115.950 568.950 118.050 571.050 ;
        RECT 101.550 566.550 106.050 568.050 ;
        RECT 107.100 567.150 108.900 568.950 ;
        RECT 102.000 565.950 106.050 566.550 ;
        RECT 89.700 555.900 96.300 556.800 ;
        RECT 89.700 555.600 91.200 555.900 ;
        RECT 86.400 549.000 88.200 555.600 ;
        RECT 89.400 549.600 91.200 555.600 ;
        RECT 95.400 555.600 96.300 555.900 ;
        RECT 92.400 549.000 94.200 555.000 ;
        RECT 95.400 549.600 97.200 555.600 ;
        RECT 107.700 549.000 109.500 561.600 ;
        RECT 112.950 555.600 114.150 568.950 ;
        RECT 122.550 568.050 123.450 571.950 ;
        RECT 128.100 571.200 129.900 573.000 ;
        RECT 134.100 571.200 135.900 573.000 ;
        RECT 137.400 571.200 138.300 574.800 ;
        RECT 149.100 571.200 150.900 573.000 ;
        RECT 155.100 571.200 156.900 573.000 ;
        RECT 158.700 571.200 159.600 578.400 ;
        RECT 175.200 576.000 177.000 584.400 ;
        RECT 173.700 574.800 177.000 576.000 ;
        RECT 181.800 575.400 183.600 585.000 ;
        RECT 194.400 577.200 196.200 584.400 ;
        RECT 199.500 578.400 201.300 585.000 ;
        RECT 209.400 579.300 211.200 584.400 ;
        RECT 212.400 580.200 214.200 585.000 ;
        RECT 215.400 579.300 217.200 584.400 ;
        RECT 209.400 577.950 217.200 579.300 ;
        RECT 218.400 578.400 220.200 584.400 ;
        RECT 194.400 576.300 198.600 577.200 ;
        RECT 218.400 576.300 219.600 578.400 ;
        RECT 160.950 573.450 163.050 574.050 ;
        RECT 160.950 572.550 168.450 573.450 ;
        RECT 160.950 571.950 163.050 572.550 ;
        RECT 127.950 569.100 130.050 571.200 ;
        RECT 130.950 569.100 133.050 571.200 ;
        RECT 133.950 569.100 136.050 571.200 ;
        RECT 136.950 569.100 139.050 571.200 ;
        RECT 148.950 569.100 151.050 571.200 ;
        RECT 151.950 569.100 154.050 571.200 ;
        RECT 154.950 569.100 157.050 571.200 ;
        RECT 157.950 569.100 160.050 571.200 ;
        RECT 122.550 566.550 127.050 568.050 ;
        RECT 131.100 567.300 132.900 569.100 ;
        RECT 123.000 565.950 127.050 566.550 ;
        RECT 137.400 556.800 138.300 569.100 ;
        RECT 142.950 567.450 145.050 567.900 ;
        RECT 148.950 567.450 151.050 568.050 ;
        RECT 142.950 566.550 151.050 567.450 ;
        RECT 152.100 567.300 153.900 569.100 ;
        RECT 142.950 565.800 145.050 566.550 ;
        RECT 148.950 565.950 151.050 566.550 ;
        RECT 158.700 561.600 159.600 569.100 ;
        RECT 167.550 568.050 168.450 572.550 ;
        RECT 173.700 571.200 174.600 574.800 ;
        RECT 176.100 571.200 177.900 573.000 ;
        RECT 182.100 571.200 183.900 573.000 ;
        RECT 194.100 571.200 195.900 573.000 ;
        RECT 197.400 571.200 198.600 576.300 ;
        RECT 215.850 575.250 219.600 576.300 ;
        RECT 235.200 576.000 237.000 584.400 ;
        RECT 200.100 571.200 201.900 573.000 ;
        RECT 172.950 569.100 175.050 571.200 ;
        RECT 175.950 569.100 178.050 571.200 ;
        RECT 178.950 569.100 181.050 571.200 ;
        RECT 181.950 569.100 184.050 571.200 ;
        RECT 193.950 569.100 196.050 571.200 ;
        RECT 196.950 569.100 199.050 571.200 ;
        RECT 199.950 569.100 202.050 571.200 ;
        RECT 212.100 571.050 213.900 572.850 ;
        RECT 215.850 571.050 217.050 575.250 ;
        RECT 233.700 574.800 237.000 576.000 ;
        RECT 241.800 575.400 243.600 585.000 ;
        RECT 251.700 578.400 253.500 585.000 ;
        RECT 256.800 577.200 258.600 584.400 ;
        RECT 271.800 578.400 273.600 584.400 ;
        RECT 274.800 578.400 276.600 585.000 ;
        RECT 288.300 580.200 290.100 584.400 ;
        RECT 287.400 578.400 290.100 580.200 ;
        RECT 291.300 578.400 293.100 585.000 ;
        RECT 254.400 576.300 258.600 577.200 ;
        RECT 218.100 571.050 219.900 572.850 ;
        RECT 233.700 571.200 234.600 574.800 ;
        RECT 236.100 571.200 237.900 573.000 ;
        RECT 242.100 571.200 243.900 573.000 ;
        RECT 251.100 571.200 252.900 573.000 ;
        RECT 254.400 571.200 255.600 576.300 ;
        RECT 267.000 573.450 271.050 574.050 ;
        RECT 257.100 571.200 258.900 573.000 ;
        RECT 266.550 571.950 271.050 573.450 ;
        RECT 167.550 566.550 172.050 568.050 ;
        RECT 168.000 565.950 172.050 566.550 ;
        RECT 131.700 555.900 138.300 556.800 ;
        RECT 131.700 555.600 133.200 555.900 ;
        RECT 112.800 549.600 114.600 555.600 ;
        RECT 115.800 549.000 117.600 555.600 ;
        RECT 128.400 549.000 130.200 555.600 ;
        RECT 131.400 549.600 133.200 555.600 ;
        RECT 137.400 555.600 138.300 555.900 ;
        RECT 149.400 560.700 157.200 561.600 ;
        RECT 134.400 549.000 136.200 555.000 ;
        RECT 137.400 549.600 139.200 555.600 ;
        RECT 149.400 549.600 151.200 560.700 ;
        RECT 152.400 549.000 154.200 559.800 ;
        RECT 155.400 549.600 157.200 560.700 ;
        RECT 158.400 549.600 160.200 561.600 ;
        RECT 173.700 556.800 174.600 569.100 ;
        RECT 179.100 567.300 180.900 569.100 ;
        RECT 175.950 564.450 178.050 565.050 ;
        RECT 187.950 564.450 190.050 565.050 ;
        RECT 175.950 563.550 190.050 564.450 ;
        RECT 175.950 562.950 178.050 563.550 ;
        RECT 187.950 562.950 190.050 563.550 ;
        RECT 173.700 555.900 180.300 556.800 ;
        RECT 173.700 555.600 174.600 555.900 ;
        RECT 172.800 549.600 174.600 555.600 ;
        RECT 178.800 555.600 180.300 555.900 ;
        RECT 197.400 555.600 198.600 569.100 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 214.950 568.950 217.050 571.050 ;
        RECT 217.950 568.950 220.050 571.050 ;
        RECT 209.100 567.150 210.900 568.950 ;
        RECT 175.800 549.000 177.600 555.000 ;
        RECT 178.800 549.600 180.600 555.600 ;
        RECT 181.800 549.000 183.600 555.600 ;
        RECT 193.800 549.000 195.600 555.600 ;
        RECT 196.800 549.600 198.600 555.600 ;
        RECT 199.800 549.000 201.600 555.600 ;
        RECT 209.700 549.000 211.500 561.600 ;
        RECT 214.950 555.600 216.150 568.950 ;
        RECT 220.950 567.450 223.050 568.050 ;
        RECT 226.950 567.450 229.050 571.050 ;
        RECT 232.950 569.100 235.050 571.200 ;
        RECT 235.950 569.100 238.050 571.200 ;
        RECT 238.950 569.100 241.050 571.200 ;
        RECT 241.950 569.100 244.050 571.200 ;
        RECT 250.950 569.100 253.050 571.200 ;
        RECT 253.950 569.100 256.050 571.200 ;
        RECT 256.950 569.100 259.050 571.200 ;
        RECT 220.950 567.000 229.050 567.450 ;
        RECT 220.950 566.550 228.450 567.000 ;
        RECT 220.950 565.950 223.050 566.550 ;
        RECT 233.700 556.800 234.600 569.100 ;
        RECT 239.100 567.300 240.900 569.100 ;
        RECT 241.950 567.450 244.050 568.050 ;
        RECT 250.950 567.450 253.050 568.050 ;
        RECT 241.950 566.550 253.050 567.450 ;
        RECT 241.950 565.950 244.050 566.550 ;
        RECT 250.950 565.950 253.050 566.550 ;
        RECT 233.700 555.900 240.300 556.800 ;
        RECT 233.700 555.600 234.600 555.900 ;
        RECT 214.800 549.600 216.600 555.600 ;
        RECT 217.800 549.000 219.600 555.600 ;
        RECT 232.800 549.600 234.600 555.600 ;
        RECT 238.800 555.600 240.300 555.900 ;
        RECT 254.400 555.600 255.600 569.100 ;
        RECT 266.550 568.050 267.450 571.950 ;
        RECT 272.400 571.200 273.600 578.400 ;
        RECT 275.100 571.200 276.900 573.000 ;
        RECT 287.400 571.200 288.300 578.400 ;
        RECT 290.100 576.600 291.900 577.500 ;
        RECT 295.800 576.600 297.600 584.400 ;
        RECT 290.100 575.700 297.600 576.600 ;
        RECT 305.400 576.600 307.200 584.400 ;
        RECT 309.900 578.400 311.700 585.000 ;
        RECT 312.900 580.200 314.700 584.400 ;
        RECT 312.900 578.400 315.600 580.200 ;
        RECT 311.100 576.600 312.900 577.500 ;
        RECT 305.400 575.700 312.900 576.600 ;
        RECT 271.950 569.100 274.050 571.200 ;
        RECT 274.950 569.100 277.050 571.200 ;
        RECT 286.950 569.100 289.050 571.200 ;
        RECT 289.950 569.100 292.050 571.200 ;
        RECT 256.950 567.450 259.050 568.050 ;
        RECT 262.950 567.450 265.050 568.050 ;
        RECT 256.950 566.550 265.050 567.450 ;
        RECT 266.550 566.550 271.050 568.050 ;
        RECT 256.950 565.950 259.050 566.550 ;
        RECT 262.950 565.950 265.050 566.550 ;
        RECT 267.000 565.950 271.050 566.550 ;
        RECT 272.400 561.600 273.600 569.100 ;
        RECT 287.400 561.600 288.300 569.100 ;
        RECT 290.100 567.300 291.900 569.100 ;
        RECT 235.800 549.000 237.600 555.000 ;
        RECT 238.800 549.600 240.600 555.600 ;
        RECT 241.800 549.000 243.600 555.600 ;
        RECT 251.400 549.000 253.200 555.600 ;
        RECT 254.400 549.600 256.200 555.600 ;
        RECT 257.400 549.000 259.200 555.600 ;
        RECT 271.800 549.600 273.600 561.600 ;
        RECT 274.800 549.000 276.600 561.600 ;
        RECT 286.800 549.600 288.600 561.600 ;
        RECT 293.700 555.600 294.600 575.700 ;
        RECT 296.100 571.200 297.900 573.000 ;
        RECT 305.100 571.200 306.900 573.000 ;
        RECT 295.950 569.100 298.050 571.200 ;
        RECT 304.950 569.100 307.050 571.200 ;
        RECT 308.400 555.600 309.300 575.700 ;
        RECT 314.700 571.200 315.600 578.400 ;
        RECT 326.400 579.300 328.200 584.400 ;
        RECT 329.400 580.200 331.200 585.000 ;
        RECT 332.400 579.300 334.200 584.400 ;
        RECT 326.400 577.950 334.200 579.300 ;
        RECT 335.400 578.400 337.200 584.400 ;
        RECT 335.400 576.300 336.600 578.400 ;
        RECT 350.400 577.200 352.200 584.400 ;
        RECT 355.500 578.400 357.300 585.000 ;
        RECT 350.400 576.300 354.600 577.200 ;
        RECT 332.850 575.250 336.600 576.300 ;
        RECT 316.950 573.450 321.000 574.050 ;
        RECT 316.950 571.950 321.450 573.450 ;
        RECT 310.950 569.100 313.050 571.200 ;
        RECT 313.950 569.100 316.050 571.200 ;
        RECT 311.100 567.300 312.900 569.100 ;
        RECT 314.700 561.600 315.600 569.100 ;
        RECT 320.550 564.450 321.450 571.950 ;
        RECT 329.100 571.050 330.900 572.850 ;
        RECT 332.850 571.050 334.050 575.250 ;
        RECT 335.100 571.050 336.900 572.850 ;
        RECT 350.100 571.200 351.900 573.000 ;
        RECT 353.400 571.200 354.600 576.300 ;
        RECT 355.950 576.450 358.050 577.050 ;
        RECT 364.950 576.450 367.050 577.050 ;
        RECT 355.950 575.550 367.050 576.450 ;
        RECT 370.200 576.000 372.000 584.400 ;
        RECT 355.950 574.950 358.050 575.550 ;
        RECT 364.950 574.950 367.050 575.550 ;
        RECT 368.700 574.800 372.000 576.000 ;
        RECT 376.800 575.400 378.600 585.000 ;
        RECT 386.400 581.400 388.200 585.000 ;
        RECT 389.400 581.400 391.200 584.400 ;
        RECT 356.100 571.200 357.900 573.000 ;
        RECT 368.700 571.200 369.600 574.800 ;
        RECT 371.100 571.200 372.900 573.000 ;
        RECT 377.100 571.200 378.900 573.000 ;
        RECT 325.950 568.950 328.050 571.050 ;
        RECT 328.950 568.950 331.050 571.050 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 349.950 569.100 352.050 571.200 ;
        RECT 352.950 569.100 355.050 571.200 ;
        RECT 355.950 569.100 358.050 571.200 ;
        RECT 367.950 569.100 370.050 571.200 ;
        RECT 370.950 569.100 373.050 571.200 ;
        RECT 373.950 569.100 376.050 571.200 ;
        RECT 376.950 569.100 379.050 571.200 ;
        RECT 389.400 571.050 390.600 581.400 ;
        RECT 401.700 578.400 403.500 585.000 ;
        RECT 406.800 577.200 408.600 584.400 ;
        RECT 421.800 578.400 423.600 584.400 ;
        RECT 404.400 576.300 408.600 577.200 ;
        RECT 422.400 576.300 423.600 578.400 ;
        RECT 424.800 579.300 426.600 584.400 ;
        RECT 427.800 580.200 429.600 585.000 ;
        RECT 430.800 579.300 432.600 584.400 ;
        RECT 424.800 577.950 432.600 579.300 ;
        RECT 435.150 578.400 436.950 584.400 ;
        RECT 438.150 581.400 439.950 585.000 ;
        RECT 442.950 582.300 444.750 584.400 ;
        RECT 441.000 581.400 444.750 582.300 ;
        RECT 447.450 581.400 449.250 585.000 ;
        RECT 450.750 581.400 452.550 584.400 ;
        RECT 454.350 581.400 456.150 585.000 ;
        RECT 458.550 581.400 460.350 584.400 ;
        RECT 463.350 581.400 465.150 585.000 ;
        RECT 441.000 580.500 442.050 581.400 ;
        RECT 450.750 580.500 451.800 581.400 ;
        RECT 439.950 578.400 442.050 580.500 ;
        RECT 396.000 573.450 400.050 574.050 ;
        RECT 395.550 571.950 400.050 573.450 ;
        RECT 326.100 567.150 327.900 568.950 ;
        RECT 325.950 564.450 328.050 565.050 ;
        RECT 320.550 563.550 328.050 564.450 ;
        RECT 325.950 562.950 328.050 563.550 ;
        RECT 289.800 549.000 291.600 555.600 ;
        RECT 292.800 549.600 294.600 555.600 ;
        RECT 295.800 549.000 297.600 555.600 ;
        RECT 305.400 549.000 307.200 555.600 ;
        RECT 308.400 549.600 310.200 555.600 ;
        RECT 311.400 549.000 313.200 555.600 ;
        RECT 314.400 549.600 316.200 561.600 ;
        RECT 326.700 549.000 328.500 561.600 ;
        RECT 331.950 555.600 333.150 568.950 ;
        RECT 353.400 555.600 354.600 569.100 ;
        RECT 368.700 556.800 369.600 569.100 ;
        RECT 374.100 567.300 375.900 569.100 ;
        RECT 385.950 568.950 388.050 571.050 ;
        RECT 388.950 568.950 391.050 571.050 ;
        RECT 386.100 567.150 387.900 568.950 ;
        RECT 368.700 555.900 375.300 556.800 ;
        RECT 368.700 555.600 369.600 555.900 ;
        RECT 331.800 549.600 333.600 555.600 ;
        RECT 334.800 549.000 336.600 555.600 ;
        RECT 349.800 549.000 351.600 555.600 ;
        RECT 352.800 549.600 354.600 555.600 ;
        RECT 355.800 549.000 357.600 555.600 ;
        RECT 367.800 549.600 369.600 555.600 ;
        RECT 373.800 555.600 375.300 555.900 ;
        RECT 389.400 555.600 390.600 568.950 ;
        RECT 395.550 568.050 396.450 571.950 ;
        RECT 401.100 571.200 402.900 573.000 ;
        RECT 404.400 571.200 405.600 576.300 ;
        RECT 422.400 575.250 426.150 576.300 ;
        RECT 407.100 571.200 408.900 573.000 ;
        RECT 400.950 569.100 403.050 571.200 ;
        RECT 403.950 569.100 406.050 571.200 ;
        RECT 406.950 569.100 409.050 571.200 ;
        RECT 422.100 571.050 423.900 572.850 ;
        RECT 424.950 571.050 426.150 575.250 ;
        RECT 428.100 571.050 429.900 572.850 ;
        RECT 391.950 566.550 396.450 568.050 ;
        RECT 391.950 565.950 396.000 566.550 ;
        RECT 404.400 555.600 405.600 569.100 ;
        RECT 421.950 568.950 424.050 571.050 ;
        RECT 424.950 568.950 427.050 571.050 ;
        RECT 427.950 568.950 430.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 425.850 555.600 427.050 568.950 ;
        RECT 431.100 567.150 432.900 568.950 ;
        RECT 435.150 563.700 436.050 578.400 ;
        RECT 443.550 577.800 445.350 579.600 ;
        RECT 446.850 579.450 451.800 580.500 ;
        RECT 459.300 580.500 460.350 581.400 ;
        RECT 446.850 578.700 448.650 579.450 ;
        RECT 459.300 579.300 463.050 580.500 ;
        RECT 460.950 578.400 463.050 579.300 ;
        RECT 466.650 578.400 468.450 584.400 ;
        RECT 443.850 576.000 444.900 577.800 ;
        RECT 454.050 576.000 455.850 576.600 ;
        RECT 443.850 574.800 455.850 576.000 ;
        RECT 438.000 573.600 444.900 574.800 ;
        RECT 438.000 572.850 438.900 573.600 ;
        RECT 443.100 573.000 444.900 573.600 ;
        RECT 437.100 571.050 438.900 572.850 ;
        RECT 440.100 571.800 441.900 572.400 ;
        RECT 436.950 568.950 439.050 571.050 ;
        RECT 440.100 570.600 448.050 571.800 ;
        RECT 445.950 568.950 448.050 570.600 ;
        RECT 444.450 563.700 446.250 564.000 ;
        RECT 435.150 563.100 446.250 563.700 ;
        RECT 435.150 562.500 452.850 563.100 ;
        RECT 435.150 561.600 436.050 562.500 ;
        RECT 444.450 562.200 452.850 562.500 ;
        RECT 370.800 549.000 372.600 555.000 ;
        RECT 373.800 549.600 375.600 555.600 ;
        RECT 376.800 549.000 378.600 555.600 ;
        RECT 386.400 549.000 388.200 555.600 ;
        RECT 389.400 549.600 391.200 555.600 ;
        RECT 401.400 549.000 403.200 555.600 ;
        RECT 404.400 549.600 406.200 555.600 ;
        RECT 407.400 549.000 409.200 555.600 ;
        RECT 422.400 549.000 424.200 555.600 ;
        RECT 425.400 549.600 427.200 555.600 ;
        RECT 430.500 549.000 432.300 561.600 ;
        RECT 435.150 549.600 436.950 561.600 ;
        RECT 449.250 560.700 451.050 561.300 ;
        RECT 443.550 559.500 451.050 560.700 ;
        RECT 451.950 560.100 452.850 562.200 ;
        RECT 454.950 562.200 455.850 574.800 ;
        RECT 467.250 571.050 468.450 578.400 ;
        RECT 479.400 577.200 481.200 584.400 ;
        RECT 484.500 578.400 486.300 585.000 ;
        RECT 496.800 578.400 498.600 584.400 ;
        RECT 479.400 576.300 483.600 577.200 ;
        RECT 479.100 571.200 480.900 573.000 ;
        RECT 482.400 571.200 483.600 576.300 ;
        RECT 497.400 576.300 498.600 578.400 ;
        RECT 499.800 579.300 501.600 584.400 ;
        RECT 502.800 580.200 504.600 585.000 ;
        RECT 505.800 579.300 507.600 584.400 ;
        RECT 499.800 577.950 507.600 579.300 ;
        RECT 517.800 578.400 519.600 584.400 ;
        RECT 520.800 578.400 522.600 585.000 ;
        RECT 530.400 579.300 532.200 584.400 ;
        RECT 533.400 580.200 535.200 585.000 ;
        RECT 536.400 579.300 538.200 584.400 ;
        RECT 497.400 575.250 501.150 576.300 ;
        RECT 485.100 571.200 486.900 573.000 ;
        RECT 462.150 569.250 468.450 571.050 ;
        RECT 463.950 568.950 468.450 569.250 ;
        RECT 478.950 569.100 481.050 571.200 ;
        RECT 481.950 569.100 484.050 571.200 ;
        RECT 484.950 569.100 487.050 571.200 ;
        RECT 497.100 571.050 498.900 572.850 ;
        RECT 499.950 571.050 501.150 575.250 ;
        RECT 503.100 571.050 504.900 572.850 ;
        RECT 518.400 571.200 519.600 578.400 ;
        RECT 530.400 577.950 538.200 579.300 ;
        RECT 539.400 578.400 541.200 584.400 ;
        RECT 551.700 578.400 553.500 585.000 ;
        RECT 539.400 576.300 540.600 578.400 ;
        RECT 556.800 577.200 558.600 584.400 ;
        RECT 569.400 581.400 571.200 585.000 ;
        RECT 572.400 581.400 574.200 584.400 ;
        RECT 575.400 581.400 577.200 585.000 ;
        RECT 536.850 575.250 540.600 576.300 ;
        RECT 544.950 576.450 547.050 577.050 ;
        RECT 550.950 576.450 553.050 576.900 ;
        RECT 544.950 575.550 553.050 576.450 ;
        RECT 521.100 571.200 522.900 573.000 ;
        RECT 464.250 563.400 466.050 565.200 ;
        RECT 460.950 562.200 465.150 563.400 ;
        RECT 454.950 561.300 460.050 562.200 ;
        RECT 460.950 561.300 463.050 562.200 ;
        RECT 467.250 561.600 468.450 568.950 ;
        RECT 459.150 560.400 460.050 561.300 ;
        RECT 456.450 560.100 458.250 560.400 ;
        RECT 443.550 558.600 444.750 559.500 ;
        RECT 451.950 559.200 458.250 560.100 ;
        RECT 456.450 558.600 458.250 559.200 ;
        RECT 459.150 558.600 461.850 560.400 ;
        RECT 439.950 556.500 444.750 558.600 ;
        RECT 447.450 557.550 449.250 558.300 ;
        RECT 452.250 557.550 454.050 558.300 ;
        RECT 447.450 556.500 454.050 557.550 ;
        RECT 443.550 555.600 444.750 556.500 ;
        RECT 438.150 549.000 439.950 555.600 ;
        RECT 443.550 549.600 445.350 555.600 ;
        RECT 448.350 549.000 450.150 555.600 ;
        RECT 451.350 549.600 453.150 556.500 ;
        RECT 459.150 555.600 463.050 557.700 ;
        RECT 454.950 549.000 456.750 555.600 ;
        RECT 459.150 549.600 460.950 555.600 ;
        RECT 463.650 549.000 465.450 552.600 ;
        RECT 466.650 549.600 468.450 561.600 ;
        RECT 482.400 555.600 483.600 569.100 ;
        RECT 496.950 568.950 499.050 571.050 ;
        RECT 499.950 568.950 502.050 571.050 ;
        RECT 502.950 568.950 505.050 571.050 ;
        RECT 505.950 568.950 508.050 571.050 ;
        RECT 517.950 569.100 520.050 571.200 ;
        RECT 520.950 569.100 523.050 571.200 ;
        RECT 533.100 571.050 534.900 572.850 ;
        RECT 536.850 571.050 538.050 575.250 ;
        RECT 544.950 574.950 547.050 575.550 ;
        RECT 550.950 574.800 553.050 575.550 ;
        RECT 554.400 576.300 558.600 577.200 ;
        RECT 539.100 571.050 540.900 572.850 ;
        RECT 551.100 571.200 552.900 573.000 ;
        RECT 554.400 571.200 555.600 576.300 ;
        RECT 557.100 571.200 558.900 573.000 ;
        RECT 500.850 555.600 502.050 568.950 ;
        RECT 506.100 567.150 507.900 568.950 ;
        RECT 518.400 561.600 519.600 569.100 ;
        RECT 529.950 568.950 532.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 550.950 569.100 553.050 571.200 ;
        RECT 553.950 569.100 556.050 571.200 ;
        RECT 556.950 569.100 559.050 571.200 ;
        RECT 572.700 571.050 573.600 581.400 ;
        RECT 587.700 578.400 589.500 585.000 ;
        RECT 592.800 577.200 594.600 584.400 ;
        RECT 605.400 579.300 607.200 584.400 ;
        RECT 608.400 580.200 610.200 585.000 ;
        RECT 611.400 579.300 613.200 584.400 ;
        RECT 605.400 577.950 613.200 579.300 ;
        RECT 614.400 578.400 616.200 584.400 ;
        RECT 628.800 581.400 630.600 585.000 ;
        RECT 631.800 581.400 633.600 584.400 ;
        RECT 634.800 581.400 636.600 585.000 ;
        RECT 644.400 584.400 645.600 585.000 ;
        RECT 644.400 581.400 646.200 584.400 ;
        RECT 647.400 581.400 649.200 584.400 ;
        RECT 650.400 581.400 652.200 585.000 ;
        RECT 590.400 576.300 594.600 577.200 ;
        RECT 614.400 576.300 615.600 578.400 ;
        RECT 587.100 571.200 588.900 573.000 ;
        RECT 590.400 571.200 591.600 576.300 ;
        RECT 611.850 575.250 615.600 576.300 ;
        RECT 593.100 571.200 594.900 573.000 ;
        RECT 530.100 567.150 531.900 568.950 ;
        RECT 478.800 549.000 480.600 555.600 ;
        RECT 481.800 549.600 483.600 555.600 ;
        RECT 484.800 549.000 486.600 555.600 ;
        RECT 497.400 549.000 499.200 555.600 ;
        RECT 500.400 549.600 502.200 555.600 ;
        RECT 505.500 549.000 507.300 561.600 ;
        RECT 517.800 549.600 519.600 561.600 ;
        RECT 520.800 549.000 522.600 561.600 ;
        RECT 530.700 549.000 532.500 561.600 ;
        RECT 535.950 555.600 537.150 568.950 ;
        RECT 554.400 555.600 555.600 569.100 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 571.950 568.950 574.050 571.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 569.100 567.150 570.900 568.950 ;
        RECT 572.700 561.600 573.600 568.950 ;
        RECT 575.100 567.150 576.900 568.950 ;
        RECT 580.950 567.450 583.050 571.050 ;
        RECT 586.950 569.100 589.050 571.200 ;
        RECT 589.950 569.100 592.050 571.200 ;
        RECT 592.950 569.100 595.050 571.200 ;
        RECT 608.100 571.050 609.900 572.850 ;
        RECT 611.850 571.050 613.050 575.250 ;
        RECT 614.100 571.050 615.900 572.850 ;
        RECT 622.950 571.950 625.050 574.050 ;
        RECT 586.950 567.450 589.050 568.050 ;
        RECT 580.950 567.000 589.050 567.450 ;
        RECT 581.550 566.550 589.050 567.000 ;
        RECT 586.950 565.950 589.050 566.550 ;
        RECT 535.800 549.600 537.600 555.600 ;
        RECT 538.800 549.000 540.600 555.600 ;
        RECT 551.400 549.000 553.200 555.600 ;
        RECT 554.400 549.600 556.200 555.600 ;
        RECT 557.400 549.000 559.200 555.600 ;
        RECT 569.400 549.000 571.200 561.600 ;
        RECT 572.700 560.400 576.300 561.600 ;
        RECT 574.500 549.600 576.300 560.400 ;
        RECT 590.400 555.600 591.600 569.100 ;
        RECT 604.950 568.950 607.050 571.050 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 605.100 567.150 606.900 568.950 ;
        RECT 587.400 549.000 589.200 555.600 ;
        RECT 590.400 549.600 592.200 555.600 ;
        RECT 593.400 549.000 595.200 555.600 ;
        RECT 605.700 549.000 607.500 561.600 ;
        RECT 610.950 555.600 612.150 568.950 ;
        RECT 623.550 568.050 624.450 571.950 ;
        RECT 632.400 571.050 633.300 581.400 ;
        RECT 648.300 577.200 649.200 581.400 ;
        RECT 653.400 578.400 655.200 584.400 ;
        RECT 648.300 576.300 651.600 577.200 ;
        RECT 649.800 575.400 651.600 576.300 ;
        RECT 644.100 571.050 645.900 572.850 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 634.950 568.950 637.050 571.050 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 623.550 566.550 628.050 568.050 ;
        RECT 629.100 567.150 630.900 568.950 ;
        RECT 624.000 565.950 628.050 566.550 ;
        RECT 632.400 561.600 633.300 568.950 ;
        RECT 635.100 567.150 636.900 568.950 ;
        RECT 647.100 567.150 648.900 568.950 ;
        RECT 650.700 564.900 651.600 575.400 ;
        RECT 654.000 571.050 655.050 578.400 ;
        RECT 658.950 574.950 661.050 577.050 ;
        RECT 665.400 575.400 667.200 585.000 ;
        RECT 672.000 576.000 673.800 584.400 ;
        RECT 688.800 581.400 690.600 584.400 ;
        RECT 691.800 581.400 693.600 585.000 ;
        RECT 649.800 564.300 651.600 564.900 ;
        RECT 644.400 563.100 651.600 564.300 ;
        RECT 652.950 568.950 655.050 571.050 ;
        RECT 644.400 561.600 645.600 563.100 ;
        RECT 652.950 561.600 654.300 568.950 ;
        RECT 659.550 568.050 660.450 574.950 ;
        RECT 672.000 574.800 675.300 576.000 ;
        RECT 665.100 571.200 666.900 573.000 ;
        RECT 671.100 571.200 672.900 573.000 ;
        RECT 674.400 571.200 675.300 574.800 ;
        RECT 664.950 569.100 667.050 571.200 ;
        RECT 667.950 569.100 670.050 571.200 ;
        RECT 670.950 569.100 673.050 571.200 ;
        RECT 673.950 569.100 676.050 571.200 ;
        RECT 689.400 571.050 690.600 581.400 ;
        RECT 703.800 578.400 705.600 584.400 ;
        RECT 704.400 576.300 705.600 578.400 ;
        RECT 706.800 579.300 708.600 584.400 ;
        RECT 709.800 580.200 711.600 585.000 ;
        RECT 712.800 579.300 714.600 584.400 ;
        RECT 724.800 581.400 726.600 584.400 ;
        RECT 727.800 581.400 729.600 585.000 ;
        RECT 740.700 581.400 742.500 585.000 ;
        RECT 706.800 577.950 714.600 579.300 ;
        RECT 704.400 575.250 708.150 576.300 ;
        RECT 704.100 571.050 705.900 572.850 ;
        RECT 706.950 571.050 708.150 575.250 ;
        RECT 710.100 571.050 711.900 572.850 ;
        RECT 725.400 571.050 726.600 581.400 ;
        RECT 743.700 579.600 745.500 584.400 ;
        RECT 740.400 578.400 745.500 579.600 ;
        RECT 748.200 578.400 750.000 585.000 ;
        RECT 740.400 571.200 741.300 578.400 ;
        RECT 758.400 576.600 760.200 584.400 ;
        RECT 762.900 578.400 764.700 585.000 ;
        RECT 765.900 580.200 767.700 584.400 ;
        RECT 765.900 578.400 768.600 580.200 ;
        RECT 781.800 578.400 783.600 584.400 ;
        RECT 784.800 581.400 786.600 585.000 ;
        RECT 791.400 584.400 792.600 585.000 ;
        RECT 787.800 581.400 789.600 584.400 ;
        RECT 790.800 581.400 792.600 584.400 ;
        RECT 764.100 576.600 765.900 577.500 ;
        RECT 758.400 575.700 765.900 576.600 ;
        RECT 743.100 571.200 744.900 573.000 ;
        RECT 749.100 571.200 750.900 573.000 ;
        RECT 758.100 571.200 759.900 573.000 ;
        RECT 655.950 566.550 660.450 568.050 ;
        RECT 668.100 567.300 669.900 569.100 ;
        RECT 655.950 565.950 660.000 566.550 ;
        RECT 629.700 560.400 633.300 561.600 ;
        RECT 610.800 549.600 612.600 555.600 ;
        RECT 613.800 549.000 615.600 555.600 ;
        RECT 629.700 549.600 631.500 560.400 ;
        RECT 634.800 549.000 636.600 561.600 ;
        RECT 644.400 549.600 646.200 561.600 ;
        RECT 648.900 549.000 650.700 561.600 ;
        RECT 651.900 560.100 654.300 561.600 ;
        RECT 658.950 561.450 661.050 562.050 ;
        RECT 670.950 561.450 673.050 561.900 ;
        RECT 658.950 560.550 673.050 561.450 ;
        RECT 651.900 549.600 653.700 560.100 ;
        RECT 658.950 559.950 661.050 560.550 ;
        RECT 670.950 559.800 673.050 560.550 ;
        RECT 674.400 556.800 675.300 569.100 ;
        RECT 688.950 568.950 691.050 571.050 ;
        RECT 691.950 568.950 694.050 571.050 ;
        RECT 703.950 568.950 706.050 571.050 ;
        RECT 706.950 568.950 709.050 571.050 ;
        RECT 709.950 568.950 712.050 571.050 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 724.950 568.950 727.050 571.050 ;
        RECT 727.950 568.950 730.050 571.050 ;
        RECT 739.950 569.100 742.050 571.200 ;
        RECT 742.950 569.100 745.050 571.200 ;
        RECT 745.950 569.100 748.050 571.200 ;
        RECT 748.950 569.100 751.050 571.200 ;
        RECT 757.950 569.100 760.050 571.200 ;
        RECT 668.700 555.900 675.300 556.800 ;
        RECT 668.700 555.600 670.200 555.900 ;
        RECT 665.400 549.000 667.200 555.600 ;
        RECT 668.400 549.600 670.200 555.600 ;
        RECT 674.400 555.600 675.300 555.900 ;
        RECT 689.400 555.600 690.600 568.950 ;
        RECT 692.100 567.150 693.900 568.950 ;
        RECT 707.850 555.600 709.050 568.950 ;
        RECT 713.100 567.150 714.900 568.950 ;
        RECT 671.400 549.000 673.200 555.000 ;
        RECT 674.400 549.600 676.200 555.600 ;
        RECT 688.800 549.600 690.600 555.600 ;
        RECT 691.800 549.000 693.600 555.600 ;
        RECT 704.400 549.000 706.200 555.600 ;
        RECT 707.400 549.600 709.200 555.600 ;
        RECT 712.500 549.000 714.300 561.600 ;
        RECT 725.400 555.600 726.600 568.950 ;
        RECT 728.100 567.150 729.900 568.950 ;
        RECT 740.400 561.600 741.300 569.100 ;
        RECT 746.100 567.300 747.900 569.100 ;
        RECT 724.800 549.600 726.600 555.600 ;
        RECT 727.800 549.000 729.600 555.600 ;
        RECT 739.800 549.600 741.600 561.600 ;
        RECT 742.800 560.700 750.600 561.600 ;
        RECT 742.800 549.600 744.600 560.700 ;
        RECT 745.800 549.000 747.600 559.800 ;
        RECT 748.800 549.600 750.600 560.700 ;
        RECT 761.400 555.600 762.300 575.700 ;
        RECT 767.700 571.200 768.600 578.400 ;
        RECT 763.950 569.100 766.050 571.200 ;
        RECT 766.950 569.100 769.050 571.200 ;
        RECT 781.950 571.050 783.000 578.400 ;
        RECT 787.800 577.200 788.700 581.400 ;
        RECT 800.700 578.400 802.500 585.000 ;
        RECT 805.800 577.200 807.600 584.400 ;
        RECT 785.400 576.300 788.700 577.200 ;
        RECT 803.400 576.300 807.600 577.200 ;
        RECT 818.400 581.400 820.200 584.400 ;
        RECT 821.400 581.400 823.200 585.000 ;
        RECT 818.400 577.500 819.600 581.400 ;
        RECT 824.400 578.400 826.200 584.400 ;
        RECT 818.400 576.600 824.100 577.500 ;
        RECT 785.400 575.400 787.200 576.300 ;
        RECT 764.100 567.300 765.900 569.100 ;
        RECT 767.700 561.600 768.600 569.100 ;
        RECT 781.950 568.950 784.050 571.050 ;
        RECT 782.700 561.600 784.050 568.950 ;
        RECT 785.400 564.900 786.300 575.400 ;
        RECT 791.100 571.050 792.900 572.850 ;
        RECT 800.100 571.200 801.900 573.000 ;
        RECT 803.400 571.200 804.600 576.300 ;
        RECT 822.150 575.700 824.100 576.600 ;
        RECT 806.100 571.200 807.900 573.000 ;
        RECT 787.950 568.950 790.050 571.050 ;
        RECT 790.950 568.950 793.050 571.050 ;
        RECT 799.950 569.100 802.050 571.200 ;
        RECT 802.950 569.100 805.050 571.200 ;
        RECT 805.950 569.100 808.050 571.200 ;
        RECT 788.100 567.150 789.900 568.950 ;
        RECT 785.400 564.300 787.200 564.900 ;
        RECT 785.400 563.100 792.600 564.300 ;
        RECT 791.400 561.600 792.600 563.100 ;
        RECT 758.400 549.000 760.200 555.600 ;
        RECT 761.400 549.600 763.200 555.600 ;
        RECT 764.400 549.000 766.200 555.600 ;
        RECT 767.400 549.600 769.200 561.600 ;
        RECT 782.700 560.100 785.100 561.600 ;
        RECT 783.300 549.600 785.100 560.100 ;
        RECT 786.300 549.000 788.100 561.600 ;
        RECT 790.800 549.600 792.600 561.600 ;
        RECT 803.400 555.600 804.600 569.100 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 818.100 567.150 819.900 568.950 ;
        RECT 822.150 564.300 823.050 575.700 ;
        RECT 825.000 571.050 826.200 578.400 ;
        RECT 836.400 576.600 838.200 584.400 ;
        RECT 840.900 578.400 842.700 585.000 ;
        RECT 843.900 580.200 845.700 584.400 ;
        RECT 843.900 578.400 846.600 580.200 ;
        RECT 842.100 576.600 843.900 577.500 ;
        RECT 836.400 575.700 843.900 576.600 ;
        RECT 831.000 573.450 835.050 574.050 ;
        RECT 823.950 568.950 826.200 571.050 ;
        RECT 822.150 563.400 824.100 564.300 ;
        RECT 818.400 562.500 824.100 563.400 ;
        RECT 818.400 555.600 819.600 562.500 ;
        RECT 825.000 561.600 826.200 568.950 ;
        RECT 830.550 571.950 835.050 573.450 ;
        RECT 830.550 568.050 831.450 571.950 ;
        RECT 836.100 571.200 837.900 573.000 ;
        RECT 835.950 569.100 838.050 571.200 ;
        RECT 830.550 566.550 835.050 568.050 ;
        RECT 831.000 565.950 835.050 566.550 ;
        RECT 800.400 549.000 802.200 555.600 ;
        RECT 803.400 549.600 805.200 555.600 ;
        RECT 806.400 549.000 808.200 555.600 ;
        RECT 818.400 549.600 820.200 555.600 ;
        RECT 821.400 549.000 823.200 555.600 ;
        RECT 824.400 549.600 826.200 561.600 ;
        RECT 839.400 555.600 840.300 575.700 ;
        RECT 845.700 571.200 846.600 578.400 ;
        RECT 841.950 569.100 844.050 571.200 ;
        RECT 844.950 569.100 847.050 571.200 ;
        RECT 842.100 567.300 843.900 569.100 ;
        RECT 845.700 561.600 846.600 569.100 ;
        RECT 836.400 549.000 838.200 555.600 ;
        RECT 839.400 549.600 841.200 555.600 ;
        RECT 842.400 549.000 844.200 555.600 ;
        RECT 845.400 549.600 847.200 561.600 ;
        RECT 10.800 533.400 12.600 545.400 ;
        RECT 13.800 534.300 15.600 545.400 ;
        RECT 16.800 535.200 18.600 546.000 ;
        RECT 19.800 534.300 21.600 545.400 ;
        RECT 29.400 539.400 31.200 546.000 ;
        RECT 32.400 539.400 34.200 545.400 ;
        RECT 35.400 540.000 37.200 546.000 ;
        RECT 32.700 539.100 34.200 539.400 ;
        RECT 38.400 539.400 40.200 545.400 ;
        RECT 50.400 539.400 52.200 546.000 ;
        RECT 53.400 539.400 55.200 545.400 ;
        RECT 56.400 540.000 58.200 546.000 ;
        RECT 38.400 539.100 39.300 539.400 ;
        RECT 32.700 538.200 39.300 539.100 ;
        RECT 53.700 539.100 55.200 539.400 ;
        RECT 59.400 539.400 61.200 545.400 ;
        RECT 59.400 539.100 60.300 539.400 ;
        RECT 53.700 538.200 60.300 539.100 ;
        RECT 13.800 533.400 21.600 534.300 ;
        RECT 11.400 525.900 12.300 533.400 ;
        RECT 13.950 531.450 16.050 532.050 ;
        RECT 28.950 531.450 31.050 532.050 ;
        RECT 13.950 530.550 31.050 531.450 ;
        RECT 13.950 529.950 16.050 530.550 ;
        RECT 28.950 529.950 31.050 530.550 ;
        RECT 17.100 525.900 18.900 527.700 ;
        RECT 32.100 525.900 33.900 527.700 ;
        RECT 38.400 525.900 39.300 538.200 ;
        RECT 43.950 528.450 46.050 529.050 ;
        RECT 49.950 528.450 52.050 529.050 ;
        RECT 43.950 527.550 52.050 528.450 ;
        RECT 43.950 526.950 46.050 527.550 ;
        RECT 49.950 526.950 52.050 527.550 ;
        RECT 53.100 525.900 54.900 527.700 ;
        RECT 59.400 525.900 60.300 538.200 ;
        RECT 73.800 533.400 75.600 545.400 ;
        RECT 76.800 534.300 78.600 545.400 ;
        RECT 79.800 535.200 81.600 546.000 ;
        RECT 82.800 534.300 84.600 545.400 ;
        RECT 76.800 533.400 84.600 534.300 ;
        RECT 94.800 533.400 96.600 545.400 ;
        RECT 97.800 534.300 99.600 545.400 ;
        RECT 100.800 535.200 102.600 546.000 ;
        RECT 103.800 534.300 105.600 545.400 ;
        RECT 115.800 539.400 117.600 545.400 ;
        RECT 118.800 540.000 120.600 546.000 ;
        RECT 97.800 533.400 105.600 534.300 ;
        RECT 116.700 539.100 117.600 539.400 ;
        RECT 121.800 539.400 123.600 545.400 ;
        RECT 124.800 539.400 126.600 546.000 ;
        RECT 134.400 539.400 136.200 546.000 ;
        RECT 137.400 539.400 139.200 545.400 ;
        RECT 121.800 539.100 123.300 539.400 ;
        RECT 116.700 538.200 123.300 539.100 ;
        RECT 74.400 525.900 75.300 533.400 ;
        RECT 82.950 528.450 85.050 529.050 ;
        RECT 88.950 528.450 91.050 529.050 ;
        RECT 80.100 525.900 81.900 527.700 ;
        RECT 82.950 527.550 91.050 528.450 ;
        RECT 82.950 526.950 85.050 527.550 ;
        RECT 88.950 526.950 91.050 527.550 ;
        RECT 95.400 525.900 96.300 533.400 ;
        RECT 101.100 525.900 102.900 527.700 ;
        RECT 116.700 525.900 117.600 538.200 ;
        RECT 118.950 531.450 121.050 532.050 ;
        RECT 124.950 531.450 127.050 532.050 ;
        RECT 118.950 530.550 127.050 531.450 ;
        RECT 118.950 529.950 121.050 530.550 ;
        RECT 124.950 529.950 127.050 530.550 ;
        RECT 122.100 525.900 123.900 527.700 ;
        RECT 134.100 526.050 135.900 527.850 ;
        RECT 137.400 526.050 138.600 539.400 ;
        RECT 149.700 533.400 151.500 546.000 ;
        RECT 154.800 539.400 156.600 545.400 ;
        RECT 157.800 539.400 159.600 546.000 ;
        RECT 172.800 544.500 180.600 545.400 ;
        RECT 139.950 528.450 144.000 529.050 ;
        RECT 139.950 526.950 144.450 528.450 ;
        RECT 10.950 523.800 13.050 525.900 ;
        RECT 13.950 523.800 16.050 525.900 ;
        RECT 16.950 523.800 19.050 525.900 ;
        RECT 19.950 523.800 22.050 525.900 ;
        RECT 28.950 523.800 31.050 525.900 ;
        RECT 31.950 523.800 34.050 525.900 ;
        RECT 34.950 523.800 37.050 525.900 ;
        RECT 37.950 523.800 40.050 525.900 ;
        RECT 49.950 523.800 52.050 525.900 ;
        RECT 52.950 523.800 55.050 525.900 ;
        RECT 55.950 523.800 58.050 525.900 ;
        RECT 58.950 523.800 61.050 525.900 ;
        RECT 73.950 523.800 76.050 525.900 ;
        RECT 76.950 523.800 79.050 525.900 ;
        RECT 79.950 523.800 82.050 525.900 ;
        RECT 82.950 523.800 85.050 525.900 ;
        RECT 94.950 523.800 97.050 525.900 ;
        RECT 97.950 523.800 100.050 525.900 ;
        RECT 100.950 523.800 103.050 525.900 ;
        RECT 103.950 523.800 106.050 525.900 ;
        RECT 115.950 523.800 118.050 525.900 ;
        RECT 118.950 523.800 121.050 525.900 ;
        RECT 121.950 523.800 124.050 525.900 ;
        RECT 124.950 523.800 127.050 525.900 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 11.400 516.600 12.300 523.800 ;
        RECT 14.100 522.000 15.900 523.800 ;
        RECT 20.100 522.000 21.900 523.800 ;
        RECT 29.100 522.000 30.900 523.800 ;
        RECT 35.100 522.000 36.900 523.800 ;
        RECT 38.400 520.200 39.300 523.800 ;
        RECT 50.100 522.000 51.900 523.800 ;
        RECT 56.100 522.000 57.900 523.800 ;
        RECT 59.400 520.200 60.300 523.800 ;
        RECT 11.400 515.400 16.500 516.600 ;
        RECT 11.700 510.000 13.500 513.600 ;
        RECT 14.700 510.600 16.500 515.400 ;
        RECT 19.200 510.000 21.000 516.600 ;
        RECT 29.400 510.000 31.200 519.600 ;
        RECT 36.000 519.000 39.300 520.200 ;
        RECT 36.000 510.600 37.800 519.000 ;
        RECT 50.400 510.000 52.200 519.600 ;
        RECT 57.000 519.000 60.300 520.200 ;
        RECT 57.000 510.600 58.800 519.000 ;
        RECT 74.400 516.600 75.300 523.800 ;
        RECT 77.100 522.000 78.900 523.800 ;
        RECT 83.100 522.000 84.900 523.800 ;
        RECT 79.950 519.450 82.050 520.050 ;
        RECT 88.950 519.450 91.050 520.050 ;
        RECT 79.950 518.550 91.050 519.450 ;
        RECT 79.950 517.950 82.050 518.550 ;
        RECT 88.950 517.950 91.050 518.550 ;
        RECT 95.400 516.600 96.300 523.800 ;
        RECT 98.100 522.000 99.900 523.800 ;
        RECT 104.100 522.000 105.900 523.800 ;
        RECT 116.700 520.200 117.600 523.800 ;
        RECT 119.100 522.000 120.900 523.800 ;
        RECT 125.100 522.000 126.900 523.800 ;
        RECT 97.950 519.450 100.050 520.050 ;
        RECT 112.950 519.450 115.050 520.050 ;
        RECT 97.950 518.550 115.050 519.450 ;
        RECT 116.700 519.000 120.000 520.200 ;
        RECT 97.950 517.950 100.050 518.550 ;
        RECT 112.950 517.950 115.050 518.550 ;
        RECT 74.400 515.400 79.500 516.600 ;
        RECT 74.700 510.000 76.500 513.600 ;
        RECT 77.700 510.600 79.500 515.400 ;
        RECT 82.200 510.000 84.000 516.600 ;
        RECT 95.400 515.400 100.500 516.600 ;
        RECT 95.700 510.000 97.500 513.600 ;
        RECT 98.700 510.600 100.500 515.400 ;
        RECT 103.200 510.000 105.000 516.600 ;
        RECT 118.200 510.600 120.000 519.000 ;
        RECT 124.800 510.000 126.600 519.600 ;
        RECT 137.400 513.600 138.600 523.950 ;
        RECT 143.550 523.050 144.450 526.950 ;
        RECT 149.100 526.050 150.900 527.850 ;
        RECT 154.950 526.050 156.150 539.400 ;
        RECT 172.800 533.400 174.600 544.500 ;
        RECT 175.800 532.500 177.600 543.600 ;
        RECT 178.800 534.600 180.600 544.500 ;
        RECT 181.800 535.500 183.600 546.000 ;
        RECT 184.800 534.600 186.600 545.400 ;
        RECT 194.400 539.400 196.200 546.000 ;
        RECT 197.400 539.400 199.200 545.400 ;
        RECT 200.400 539.400 202.200 546.000 ;
        RECT 178.800 533.700 186.600 534.600 ;
        RECT 175.800 531.600 180.900 532.500 ;
        RECT 163.950 526.950 166.050 529.050 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 143.550 521.550 148.050 523.050 ;
        RECT 152.100 522.150 153.900 523.950 ;
        RECT 144.000 520.950 148.050 521.550 ;
        RECT 155.850 519.750 157.050 523.950 ;
        RECT 158.100 522.150 159.900 523.950 ;
        RECT 164.550 523.050 165.450 526.950 ;
        RECT 176.100 525.900 177.900 527.700 ;
        RECT 180.000 525.900 180.900 531.600 ;
        RECT 182.100 525.900 183.900 527.700 ;
        RECT 172.950 523.800 175.050 525.900 ;
        RECT 175.950 523.800 178.050 525.900 ;
        RECT 178.950 523.800 181.050 525.900 ;
        RECT 181.950 523.800 184.050 525.900 ;
        RECT 184.950 523.800 187.050 525.900 ;
        RECT 193.950 523.800 196.050 525.900 ;
        RECT 160.950 521.550 165.450 523.050 ;
        RECT 173.100 522.000 174.900 523.800 ;
        RECT 160.950 520.950 165.000 521.550 ;
        RECT 155.850 518.700 159.600 519.750 ;
        RECT 149.400 515.700 157.200 517.050 ;
        RECT 134.400 510.000 136.200 513.600 ;
        RECT 137.400 510.600 139.200 513.600 ;
        RECT 149.400 510.600 151.200 515.700 ;
        RECT 152.400 510.000 154.200 514.800 ;
        RECT 155.400 510.600 157.200 515.700 ;
        RECT 158.400 516.600 159.600 518.700 ;
        RECT 180.000 516.600 181.050 523.800 ;
        RECT 185.100 522.000 186.900 523.800 ;
        RECT 194.100 522.000 195.900 523.800 ;
        RECT 197.400 519.300 198.300 539.400 ;
        RECT 203.400 533.400 205.200 545.400 ;
        RECT 215.400 539.400 217.200 546.000 ;
        RECT 218.400 539.400 220.200 545.400 ;
        RECT 221.400 539.400 223.200 546.000 ;
        RECT 200.100 525.900 201.900 527.700 ;
        RECT 203.700 525.900 204.600 533.400 ;
        RECT 214.950 528.450 217.050 529.050 ;
        RECT 209.550 527.550 217.050 528.450 ;
        RECT 199.950 523.800 202.050 525.900 ;
        RECT 202.950 523.800 205.050 525.900 ;
        RECT 194.400 518.400 201.900 519.300 ;
        RECT 158.400 510.600 160.200 516.600 ;
        RECT 175.500 510.000 177.300 516.600 ;
        RECT 180.000 510.600 181.800 516.600 ;
        RECT 184.500 510.000 186.300 516.600 ;
        RECT 194.400 510.600 196.200 518.400 ;
        RECT 200.100 517.500 201.900 518.400 ;
        RECT 203.700 516.600 204.600 523.800 ;
        RECT 209.550 523.050 210.450 527.550 ;
        RECT 214.950 526.950 217.050 527.550 ;
        RECT 218.400 525.900 219.600 539.400 ;
        RECT 235.800 533.400 237.600 545.400 ;
        RECT 238.800 534.300 240.600 545.400 ;
        RECT 241.800 535.200 243.600 546.000 ;
        RECT 244.800 534.300 246.600 545.400 ;
        RECT 257.400 539.400 259.200 546.000 ;
        RECT 260.400 539.400 262.200 545.400 ;
        RECT 238.800 533.400 246.600 534.300 ;
        RECT 236.400 525.900 237.300 533.400 ;
        RECT 242.100 525.900 243.900 527.700 ;
        RECT 260.850 526.050 262.050 539.400 ;
        RECT 265.500 533.400 267.300 546.000 ;
        RECT 278.400 539.400 280.200 546.000 ;
        RECT 281.400 539.400 283.200 545.400 ;
        RECT 273.000 528.450 277.050 529.050 ;
        RECT 266.100 526.050 267.900 527.850 ;
        RECT 272.550 526.950 277.050 528.450 ;
        RECT 214.950 523.800 217.050 525.900 ;
        RECT 217.950 523.800 220.050 525.900 ;
        RECT 220.950 523.800 223.050 525.900 ;
        RECT 235.950 523.800 238.050 525.900 ;
        RECT 238.950 523.800 241.050 525.900 ;
        RECT 241.950 523.800 244.050 525.900 ;
        RECT 244.950 523.800 247.050 525.900 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 205.950 521.550 210.450 523.050 ;
        RECT 215.100 522.000 216.900 523.800 ;
        RECT 205.950 520.950 210.000 521.550 ;
        RECT 218.400 518.700 219.600 523.800 ;
        RECT 221.100 522.000 222.900 523.800 ;
        RECT 218.400 517.800 222.600 518.700 ;
        RECT 198.900 510.000 200.700 516.600 ;
        RECT 201.900 514.800 204.600 516.600 ;
        RECT 201.900 510.600 203.700 514.800 ;
        RECT 215.700 510.000 217.500 516.600 ;
        RECT 220.800 510.600 222.600 517.800 ;
        RECT 236.400 516.600 237.300 523.800 ;
        RECT 239.100 522.000 240.900 523.800 ;
        RECT 245.100 522.000 246.900 523.800 ;
        RECT 257.100 522.150 258.900 523.950 ;
        RECT 259.950 519.750 261.150 523.950 ;
        RECT 263.100 522.150 264.900 523.950 ;
        RECT 272.550 523.050 273.450 526.950 ;
        RECT 281.850 526.050 283.050 539.400 ;
        RECT 286.500 533.400 288.300 546.000 ;
        RECT 296.400 539.400 298.200 546.000 ;
        RECT 299.400 539.400 301.200 545.400 ;
        RECT 302.400 539.400 304.200 546.000 ;
        RECT 287.100 526.050 288.900 527.850 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 286.950 523.950 289.050 526.050 ;
        RECT 299.400 525.900 300.600 539.400 ;
        RECT 314.700 533.400 316.500 546.000 ;
        RECT 319.800 539.400 321.600 545.400 ;
        RECT 322.800 539.400 324.600 546.000 ;
        RECT 337.800 539.400 339.600 546.000 ;
        RECT 340.800 539.400 342.600 545.400 ;
        RECT 343.800 539.400 345.600 546.000 ;
        RECT 355.800 539.400 357.600 546.000 ;
        RECT 358.800 539.400 360.600 545.400 ;
        RECT 361.800 539.400 363.600 546.000 ;
        RECT 374.400 539.400 376.200 546.000 ;
        RECT 377.400 539.400 379.200 545.400 ;
        RECT 314.100 526.050 315.900 527.850 ;
        RECT 319.950 526.050 321.150 539.400 ;
        RECT 325.950 528.450 328.050 532.050 ;
        RECT 325.950 528.000 330.450 528.450 ;
        RECT 326.550 527.550 330.450 528.000 ;
        RECT 268.950 521.550 273.450 523.050 ;
        RECT 278.100 522.150 279.900 523.950 ;
        RECT 268.950 520.950 273.000 521.550 ;
        RECT 280.950 519.750 282.150 523.950 ;
        RECT 284.100 522.150 285.900 523.950 ;
        RECT 295.950 523.800 298.050 525.900 ;
        RECT 298.950 523.800 301.050 525.900 ;
        RECT 301.950 523.800 304.050 525.900 ;
        RECT 313.950 523.950 316.050 526.050 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 319.950 523.950 322.050 526.050 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 296.100 522.000 297.900 523.800 ;
        RECT 257.400 518.700 261.150 519.750 ;
        RECT 278.400 518.700 282.150 519.750 ;
        RECT 299.400 518.700 300.600 523.800 ;
        RECT 302.100 522.000 303.900 523.800 ;
        RECT 317.100 522.150 318.900 523.950 ;
        RECT 320.850 519.750 322.050 523.950 ;
        RECT 323.100 522.150 324.900 523.950 ;
        RECT 329.550 522.450 330.450 527.550 ;
        RECT 341.400 525.900 342.600 539.400 ;
        RECT 359.400 525.900 360.600 539.400 ;
        RECT 367.950 531.450 370.050 532.050 ;
        RECT 373.950 531.450 376.050 532.050 ;
        RECT 367.950 530.550 376.050 531.450 ;
        RECT 367.950 529.950 370.050 530.550 ;
        RECT 373.950 529.950 376.050 530.550 ;
        RECT 364.950 528.450 369.000 529.050 ;
        RECT 364.950 526.950 369.450 528.450 ;
        RECT 337.950 523.800 340.050 525.900 ;
        RECT 340.950 523.800 343.050 525.900 ;
        RECT 343.950 523.800 346.050 525.900 ;
        RECT 355.950 523.800 358.050 525.900 ;
        RECT 358.950 523.800 361.050 525.900 ;
        RECT 361.950 523.800 364.050 525.900 ;
        RECT 334.950 522.450 337.050 523.050 ;
        RECT 329.550 521.550 337.050 522.450 ;
        RECT 338.100 522.000 339.900 523.800 ;
        RECT 334.950 520.950 337.050 521.550 ;
        RECT 320.850 518.700 324.600 519.750 ;
        RECT 341.400 518.700 342.600 523.800 ;
        RECT 344.100 522.000 345.900 523.800 ;
        RECT 356.100 522.000 357.900 523.800 ;
        RECT 359.400 518.700 360.600 523.800 ;
        RECT 362.100 522.000 363.900 523.800 ;
        RECT 368.550 523.050 369.450 526.950 ;
        RECT 377.850 526.050 379.050 539.400 ;
        RECT 382.500 533.400 384.300 546.000 ;
        RECT 392.400 539.400 394.200 546.000 ;
        RECT 395.400 539.400 397.200 545.400 ;
        RECT 398.400 539.400 400.200 546.000 ;
        RECT 383.100 526.050 384.900 527.850 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 376.950 523.950 379.050 526.050 ;
        RECT 379.950 523.950 382.050 526.050 ;
        RECT 382.950 523.950 385.050 526.050 ;
        RECT 395.400 525.900 396.600 539.400 ;
        RECT 410.700 533.400 412.500 546.000 ;
        RECT 415.800 539.400 417.600 545.400 ;
        RECT 418.800 539.400 420.600 546.000 ;
        RECT 431.400 539.400 433.200 546.000 ;
        RECT 434.400 539.400 436.200 545.400 ;
        RECT 437.400 539.400 439.200 546.000 ;
        RECT 408.000 531.900 411.000 532.050 ;
        RECT 406.950 531.450 411.000 531.900 ;
        RECT 404.550 530.550 411.450 531.450 ;
        RECT 364.950 521.550 369.450 523.050 ;
        RECT 374.100 522.150 375.900 523.950 ;
        RECT 364.950 520.950 369.000 521.550 ;
        RECT 376.950 519.750 378.150 523.950 ;
        RECT 380.100 522.150 381.900 523.950 ;
        RECT 391.950 523.800 394.050 525.900 ;
        RECT 394.950 523.800 397.050 525.900 ;
        RECT 397.950 523.800 400.050 525.900 ;
        RECT 392.100 522.000 393.900 523.800 ;
        RECT 257.400 516.600 258.600 518.700 ;
        RECT 236.400 515.400 241.500 516.600 ;
        RECT 236.700 510.000 238.500 513.600 ;
        RECT 239.700 510.600 241.500 515.400 ;
        RECT 244.200 510.000 246.000 516.600 ;
        RECT 256.800 510.600 258.600 516.600 ;
        RECT 259.800 515.700 267.600 517.050 ;
        RECT 278.400 516.600 279.600 518.700 ;
        RECT 299.400 517.800 303.600 518.700 ;
        RECT 259.800 510.600 261.600 515.700 ;
        RECT 262.800 510.000 264.600 514.800 ;
        RECT 265.800 510.600 267.600 515.700 ;
        RECT 277.800 510.600 279.600 516.600 ;
        RECT 280.800 515.700 288.600 517.050 ;
        RECT 280.800 510.600 282.600 515.700 ;
        RECT 283.800 510.000 285.600 514.800 ;
        RECT 286.800 510.600 288.600 515.700 ;
        RECT 296.700 510.000 298.500 516.600 ;
        RECT 301.800 510.600 303.600 517.800 ;
        RECT 314.400 515.700 322.200 517.050 ;
        RECT 314.400 510.600 316.200 515.700 ;
        RECT 317.400 510.000 319.200 514.800 ;
        RECT 320.400 510.600 322.200 515.700 ;
        RECT 323.400 516.600 324.600 518.700 ;
        RECT 338.400 517.800 342.600 518.700 ;
        RECT 356.400 517.800 360.600 518.700 ;
        RECT 374.400 518.700 378.150 519.750 ;
        RECT 395.400 518.700 396.600 523.800 ;
        RECT 398.100 522.000 399.900 523.800 ;
        RECT 404.550 523.050 405.450 530.550 ;
        RECT 406.950 529.950 411.000 530.550 ;
        RECT 406.950 529.800 409.050 529.950 ;
        RECT 410.100 526.050 411.900 527.850 ;
        RECT 415.950 526.050 417.150 539.400 ;
        RECT 421.950 534.450 424.050 535.050 ;
        RECT 430.950 534.450 433.050 535.050 ;
        RECT 421.950 533.550 433.050 534.450 ;
        RECT 421.950 532.950 424.050 533.550 ;
        RECT 430.950 532.950 433.050 533.550 ;
        RECT 424.950 528.450 427.050 529.050 ;
        RECT 430.950 528.450 433.050 529.050 ;
        RECT 424.950 527.550 433.050 528.450 ;
        RECT 424.950 526.950 427.050 527.550 ;
        RECT 430.950 526.950 433.050 527.550 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 434.400 525.900 435.600 539.400 ;
        RECT 444.150 533.400 445.950 545.400 ;
        RECT 447.150 539.400 448.950 546.000 ;
        RECT 452.550 539.400 454.350 545.400 ;
        RECT 457.350 539.400 459.150 546.000 ;
        RECT 452.550 538.500 453.750 539.400 ;
        RECT 460.350 538.500 462.150 545.400 ;
        RECT 463.950 539.400 465.750 546.000 ;
        RECT 468.150 539.400 469.950 545.400 ;
        RECT 472.650 542.400 474.450 546.000 ;
        RECT 448.950 536.400 453.750 538.500 ;
        RECT 456.450 537.450 463.050 538.500 ;
        RECT 456.450 536.700 458.250 537.450 ;
        RECT 461.250 536.700 463.050 537.450 ;
        RECT 468.150 537.300 472.050 539.400 ;
        RECT 452.550 535.500 453.750 536.400 ;
        RECT 465.450 535.800 467.250 536.400 ;
        RECT 452.550 534.300 460.050 535.500 ;
        RECT 458.250 533.700 460.050 534.300 ;
        RECT 460.950 534.900 467.250 535.800 ;
        RECT 444.150 532.500 445.050 533.400 ;
        RECT 460.950 532.800 461.850 534.900 ;
        RECT 465.450 534.600 467.250 534.900 ;
        RECT 468.150 534.600 470.850 536.400 ;
        RECT 468.150 533.700 469.050 534.600 ;
        RECT 453.450 532.500 461.850 532.800 ;
        RECT 444.150 531.900 461.850 532.500 ;
        RECT 463.950 532.800 469.050 533.700 ;
        RECT 469.950 532.800 472.050 533.700 ;
        RECT 475.650 533.400 477.450 545.400 ;
        RECT 490.800 539.400 492.600 546.000 ;
        RECT 493.800 539.400 495.600 545.400 ;
        RECT 496.800 539.400 498.600 546.000 ;
        RECT 444.150 531.300 455.250 531.900 ;
        RECT 404.550 521.550 409.050 523.050 ;
        RECT 413.100 522.150 414.900 523.950 ;
        RECT 405.000 520.950 409.050 521.550 ;
        RECT 416.850 519.750 418.050 523.950 ;
        RECT 419.100 522.150 420.900 523.950 ;
        RECT 430.950 523.800 433.050 525.900 ;
        RECT 433.950 523.800 436.050 525.900 ;
        RECT 436.950 523.800 439.050 525.900 ;
        RECT 431.100 522.000 432.900 523.800 ;
        RECT 416.850 518.700 420.600 519.750 ;
        RECT 323.400 510.600 325.200 516.600 ;
        RECT 328.950 513.450 331.050 514.050 ;
        RECT 334.950 513.450 337.050 514.050 ;
        RECT 328.950 512.550 337.050 513.450 ;
        RECT 328.950 511.950 331.050 512.550 ;
        RECT 334.950 511.950 337.050 512.550 ;
        RECT 338.400 510.600 340.200 517.800 ;
        RECT 343.500 510.000 345.300 516.600 ;
        RECT 356.400 510.600 358.200 517.800 ;
        RECT 374.400 516.600 375.600 518.700 ;
        RECT 395.400 517.800 399.600 518.700 ;
        RECT 361.500 510.000 363.300 516.600 ;
        RECT 373.800 510.600 375.600 516.600 ;
        RECT 376.800 515.700 384.600 517.050 ;
        RECT 376.800 510.600 378.600 515.700 ;
        RECT 379.800 510.000 381.600 514.800 ;
        RECT 382.800 510.600 384.600 515.700 ;
        RECT 392.700 510.000 394.500 516.600 ;
        RECT 397.800 510.600 399.600 517.800 ;
        RECT 410.400 515.700 418.200 517.050 ;
        RECT 410.400 510.600 412.200 515.700 ;
        RECT 413.400 510.000 415.200 514.800 ;
        RECT 416.400 510.600 418.200 515.700 ;
        RECT 419.400 516.600 420.600 518.700 ;
        RECT 434.400 518.700 435.600 523.800 ;
        RECT 437.100 522.000 438.900 523.800 ;
        RECT 434.400 517.800 438.600 518.700 ;
        RECT 419.400 510.600 421.200 516.600 ;
        RECT 431.700 510.000 433.500 516.600 ;
        RECT 436.800 510.600 438.600 517.800 ;
        RECT 444.150 516.600 445.050 531.300 ;
        RECT 453.450 531.000 455.250 531.300 ;
        RECT 445.950 523.950 448.050 526.050 ;
        RECT 454.950 524.400 457.050 526.050 ;
        RECT 446.100 522.150 447.900 523.950 ;
        RECT 449.100 523.200 457.050 524.400 ;
        RECT 449.100 522.600 450.900 523.200 ;
        RECT 447.000 521.400 447.900 522.150 ;
        RECT 452.100 521.400 453.900 522.000 ;
        RECT 447.000 520.200 453.900 521.400 ;
        RECT 463.950 520.200 464.850 532.800 ;
        RECT 469.950 531.600 474.150 532.800 ;
        RECT 473.250 529.800 475.050 531.600 ;
        RECT 476.250 526.050 477.450 533.400 ;
        RECT 484.950 529.950 487.050 532.050 ;
        RECT 472.950 525.750 477.450 526.050 ;
        RECT 471.150 523.950 477.450 525.750 ;
        RECT 452.850 519.000 464.850 520.200 ;
        RECT 452.850 517.200 453.900 519.000 ;
        RECT 463.050 518.400 464.850 519.000 ;
        RECT 444.150 510.600 445.950 516.600 ;
        RECT 448.950 514.500 451.050 516.600 ;
        RECT 452.550 515.400 454.350 517.200 ;
        RECT 476.250 516.600 477.450 523.950 ;
        RECT 485.550 523.050 486.450 529.950 ;
        RECT 494.400 525.900 495.600 539.400 ;
        RECT 506.700 533.400 508.500 546.000 ;
        RECT 511.800 539.400 513.600 545.400 ;
        RECT 514.800 539.400 516.600 546.000 ;
        RECT 527.400 539.400 529.200 546.000 ;
        RECT 530.400 539.400 532.200 545.400 ;
        RECT 533.400 539.400 535.200 546.000 ;
        RECT 548.400 539.400 550.200 546.000 ;
        RECT 551.400 539.400 553.200 545.400 ;
        RECT 506.100 526.050 507.900 527.850 ;
        RECT 511.950 526.050 513.150 539.400 ;
        RECT 490.950 523.800 493.050 525.900 ;
        RECT 493.950 523.800 496.050 525.900 ;
        RECT 496.950 523.800 499.050 525.900 ;
        RECT 505.950 523.950 508.050 526.050 ;
        RECT 508.950 523.950 511.050 526.050 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 514.950 523.950 517.050 526.050 ;
        RECT 530.400 525.900 531.600 539.400 ;
        RECT 532.950 528.450 535.050 529.050 ;
        RECT 538.950 528.450 541.050 529.050 ;
        RECT 532.950 527.550 541.050 528.450 ;
        RECT 532.950 526.950 535.050 527.550 ;
        RECT 538.950 526.950 541.050 527.550 ;
        RECT 551.850 526.050 553.050 539.400 ;
        RECT 556.500 533.400 558.300 546.000 ;
        RECT 561.150 533.400 562.950 545.400 ;
        RECT 564.150 539.400 565.950 546.000 ;
        RECT 569.550 539.400 571.350 545.400 ;
        RECT 574.350 539.400 576.150 546.000 ;
        RECT 569.550 538.500 570.750 539.400 ;
        RECT 577.350 538.500 579.150 545.400 ;
        RECT 580.950 539.400 582.750 546.000 ;
        RECT 585.150 539.400 586.950 545.400 ;
        RECT 589.650 542.400 591.450 546.000 ;
        RECT 565.950 536.400 570.750 538.500 ;
        RECT 573.450 537.450 580.050 538.500 ;
        RECT 573.450 536.700 575.250 537.450 ;
        RECT 578.250 536.700 580.050 537.450 ;
        RECT 585.150 537.300 589.050 539.400 ;
        RECT 569.550 535.500 570.750 536.400 ;
        RECT 582.450 535.800 584.250 536.400 ;
        RECT 569.550 534.300 577.050 535.500 ;
        RECT 575.250 533.700 577.050 534.300 ;
        RECT 577.950 534.900 584.250 535.800 ;
        RECT 561.150 532.500 562.050 533.400 ;
        RECT 577.950 532.800 578.850 534.900 ;
        RECT 582.450 534.600 584.250 534.900 ;
        RECT 585.150 534.600 587.850 536.400 ;
        RECT 585.150 533.700 586.050 534.600 ;
        RECT 570.450 532.500 578.850 532.800 ;
        RECT 561.150 531.900 578.850 532.500 ;
        RECT 580.950 532.800 586.050 533.700 ;
        RECT 586.950 532.800 589.050 533.700 ;
        RECT 592.650 533.400 594.450 545.400 ;
        RECT 604.800 539.400 606.600 546.000 ;
        RECT 607.800 539.400 609.600 545.400 ;
        RECT 610.800 539.400 612.600 546.000 ;
        RECT 561.150 531.300 572.250 531.900 ;
        RECT 557.100 526.050 558.900 527.850 ;
        RECT 485.550 521.550 490.050 523.050 ;
        RECT 491.100 522.000 492.900 523.800 ;
        RECT 486.000 520.950 490.050 521.550 ;
        RECT 494.400 518.700 495.600 523.800 ;
        RECT 497.100 522.000 498.900 523.800 ;
        RECT 509.100 522.150 510.900 523.950 ;
        RECT 512.850 519.750 514.050 523.950 ;
        RECT 515.100 522.150 516.900 523.950 ;
        RECT 526.950 523.800 529.050 525.900 ;
        RECT 529.950 523.800 532.050 525.900 ;
        RECT 532.950 523.800 535.050 525.900 ;
        RECT 547.950 523.950 550.050 526.050 ;
        RECT 550.950 523.950 553.050 526.050 ;
        RECT 553.950 523.950 556.050 526.050 ;
        RECT 556.950 523.950 559.050 526.050 ;
        RECT 527.100 522.000 528.900 523.800 ;
        RECT 512.850 518.700 516.600 519.750 ;
        RECT 455.850 515.550 457.650 516.300 ;
        RECT 469.950 515.700 472.050 516.600 ;
        RECT 455.850 514.500 460.800 515.550 ;
        RECT 450.000 513.600 451.050 514.500 ;
        RECT 459.750 513.600 460.800 514.500 ;
        RECT 468.300 514.500 472.050 515.700 ;
        RECT 468.300 513.600 469.350 514.500 ;
        RECT 447.150 510.000 448.950 513.600 ;
        RECT 450.000 512.700 453.750 513.600 ;
        RECT 451.950 510.600 453.750 512.700 ;
        RECT 456.450 510.000 458.250 513.600 ;
        RECT 459.750 510.600 461.550 513.600 ;
        RECT 463.350 510.000 465.150 513.600 ;
        RECT 467.550 510.600 469.350 513.600 ;
        RECT 472.350 510.000 474.150 513.600 ;
        RECT 475.650 510.600 477.450 516.600 ;
        RECT 491.400 517.800 495.600 518.700 ;
        RECT 491.400 510.600 493.200 517.800 ;
        RECT 496.500 510.000 498.300 516.600 ;
        RECT 506.400 515.700 514.200 517.050 ;
        RECT 506.400 510.600 508.200 515.700 ;
        RECT 509.400 510.000 511.200 514.800 ;
        RECT 512.400 510.600 514.200 515.700 ;
        RECT 515.400 516.600 516.600 518.700 ;
        RECT 530.400 518.700 531.600 523.800 ;
        RECT 533.100 522.000 534.900 523.800 ;
        RECT 538.950 522.450 541.050 523.050 ;
        RECT 544.950 522.450 547.050 523.050 ;
        RECT 538.950 521.550 547.050 522.450 ;
        RECT 548.100 522.150 549.900 523.950 ;
        RECT 538.950 520.950 541.050 521.550 ;
        RECT 544.950 520.950 547.050 521.550 ;
        RECT 550.950 519.750 552.150 523.950 ;
        RECT 554.100 522.150 555.900 523.950 ;
        RECT 548.400 518.700 552.150 519.750 ;
        RECT 530.400 517.800 534.600 518.700 ;
        RECT 515.400 510.600 517.200 516.600 ;
        RECT 527.700 510.000 529.500 516.600 ;
        RECT 532.800 510.600 534.600 517.800 ;
        RECT 548.400 516.600 549.600 518.700 ;
        RECT 547.800 510.600 549.600 516.600 ;
        RECT 550.800 515.700 558.600 517.050 ;
        RECT 550.800 510.600 552.600 515.700 ;
        RECT 553.800 510.000 555.600 514.800 ;
        RECT 556.800 510.600 558.600 515.700 ;
        RECT 561.150 516.600 562.050 531.300 ;
        RECT 570.450 531.000 572.250 531.300 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 571.950 524.400 574.050 526.050 ;
        RECT 563.100 522.150 564.900 523.950 ;
        RECT 566.100 523.200 574.050 524.400 ;
        RECT 566.100 522.600 567.900 523.200 ;
        RECT 564.000 521.400 564.900 522.150 ;
        RECT 569.100 521.400 570.900 522.000 ;
        RECT 564.000 520.200 570.900 521.400 ;
        RECT 580.950 520.200 581.850 532.800 ;
        RECT 586.950 531.600 591.150 532.800 ;
        RECT 590.250 529.800 592.050 531.600 ;
        RECT 593.250 526.050 594.450 533.400 ;
        RECT 589.950 525.750 594.450 526.050 ;
        RECT 608.400 525.900 609.600 539.400 ;
        RECT 615.150 533.400 616.950 545.400 ;
        RECT 618.150 539.400 619.950 546.000 ;
        RECT 623.550 539.400 625.350 545.400 ;
        RECT 628.350 539.400 630.150 546.000 ;
        RECT 623.550 538.500 624.750 539.400 ;
        RECT 631.350 538.500 633.150 545.400 ;
        RECT 634.950 539.400 636.750 546.000 ;
        RECT 639.150 539.400 640.950 545.400 ;
        RECT 643.650 542.400 645.450 546.000 ;
        RECT 619.950 536.400 624.750 538.500 ;
        RECT 627.450 537.450 634.050 538.500 ;
        RECT 627.450 536.700 629.250 537.450 ;
        RECT 632.250 536.700 634.050 537.450 ;
        RECT 639.150 537.300 643.050 539.400 ;
        RECT 623.550 535.500 624.750 536.400 ;
        RECT 636.450 535.800 638.250 536.400 ;
        RECT 623.550 534.300 631.050 535.500 ;
        RECT 629.250 533.700 631.050 534.300 ;
        RECT 631.950 534.900 638.250 535.800 ;
        RECT 615.150 532.500 616.050 533.400 ;
        RECT 631.950 532.800 632.850 534.900 ;
        RECT 636.450 534.600 638.250 534.900 ;
        RECT 639.150 534.600 641.850 536.400 ;
        RECT 639.150 533.700 640.050 534.600 ;
        RECT 624.450 532.500 632.850 532.800 ;
        RECT 615.150 531.900 632.850 532.500 ;
        RECT 634.950 532.800 640.050 533.700 ;
        RECT 640.950 532.800 643.050 533.700 ;
        RECT 646.650 533.400 648.450 545.400 ;
        RECT 656.400 539.400 658.200 546.000 ;
        RECT 659.400 539.400 661.200 545.400 ;
        RECT 662.400 539.400 664.200 546.000 ;
        RECT 615.150 531.300 626.250 531.900 ;
        RECT 588.150 523.950 594.450 525.750 ;
        RECT 569.850 519.000 581.850 520.200 ;
        RECT 569.850 517.200 570.900 519.000 ;
        RECT 580.050 518.400 581.850 519.000 ;
        RECT 561.150 510.600 562.950 516.600 ;
        RECT 565.950 514.500 568.050 516.600 ;
        RECT 569.550 515.400 571.350 517.200 ;
        RECT 593.250 516.600 594.450 523.950 ;
        RECT 604.950 523.800 607.050 525.900 ;
        RECT 607.950 523.800 610.050 525.900 ;
        RECT 610.950 523.800 613.050 525.900 ;
        RECT 605.100 522.000 606.900 523.800 ;
        RECT 608.400 518.700 609.600 523.800 ;
        RECT 611.100 522.000 612.900 523.800 ;
        RECT 572.850 515.550 574.650 516.300 ;
        RECT 586.950 515.700 589.050 516.600 ;
        RECT 572.850 514.500 577.800 515.550 ;
        RECT 567.000 513.600 568.050 514.500 ;
        RECT 576.750 513.600 577.800 514.500 ;
        RECT 585.300 514.500 589.050 515.700 ;
        RECT 585.300 513.600 586.350 514.500 ;
        RECT 564.150 510.000 565.950 513.600 ;
        RECT 567.000 512.700 570.750 513.600 ;
        RECT 568.950 510.600 570.750 512.700 ;
        RECT 573.450 510.000 575.250 513.600 ;
        RECT 576.750 510.600 578.550 513.600 ;
        RECT 580.350 510.000 582.150 513.600 ;
        RECT 584.550 510.600 586.350 513.600 ;
        RECT 589.350 510.000 591.150 513.600 ;
        RECT 592.650 510.600 594.450 516.600 ;
        RECT 605.400 517.800 609.600 518.700 ;
        RECT 605.400 510.600 607.200 517.800 ;
        RECT 615.150 516.600 616.050 531.300 ;
        RECT 624.450 531.000 626.250 531.300 ;
        RECT 616.950 523.950 619.050 526.050 ;
        RECT 625.950 524.400 628.050 526.050 ;
        RECT 617.100 522.150 618.900 523.950 ;
        RECT 620.100 523.200 628.050 524.400 ;
        RECT 620.100 522.600 621.900 523.200 ;
        RECT 618.000 521.400 618.900 522.150 ;
        RECT 623.100 521.400 624.900 522.000 ;
        RECT 618.000 520.200 624.900 521.400 ;
        RECT 634.950 520.200 635.850 532.800 ;
        RECT 640.950 531.600 645.150 532.800 ;
        RECT 644.250 529.800 646.050 531.600 ;
        RECT 647.250 526.050 648.450 533.400 ;
        RECT 649.950 529.950 652.050 532.050 ;
        RECT 643.950 525.750 648.450 526.050 ;
        RECT 642.150 523.950 648.450 525.750 ;
        RECT 623.850 519.000 635.850 520.200 ;
        RECT 623.850 517.200 624.900 519.000 ;
        RECT 634.050 518.400 635.850 519.000 ;
        RECT 610.500 510.000 612.300 516.600 ;
        RECT 615.150 510.600 616.950 516.600 ;
        RECT 619.950 514.500 622.050 516.600 ;
        RECT 623.550 515.400 625.350 517.200 ;
        RECT 647.250 516.600 648.450 523.950 ;
        RECT 650.550 523.050 651.450 529.950 ;
        RECT 659.400 525.900 660.600 539.400 ;
        RECT 674.700 533.400 676.500 546.000 ;
        RECT 679.800 539.400 681.600 545.400 ;
        RECT 682.800 539.400 684.600 546.000 ;
        RECT 698.400 539.400 700.200 546.000 ;
        RECT 701.400 539.400 703.200 545.400 ;
        RECT 669.000 528.450 673.050 529.050 ;
        RECT 668.550 526.950 673.050 528.450 ;
        RECT 655.950 523.800 658.050 525.900 ;
        RECT 658.950 523.800 661.050 525.900 ;
        RECT 661.950 523.800 664.050 525.900 ;
        RECT 650.550 521.550 655.050 523.050 ;
        RECT 656.100 522.000 657.900 523.800 ;
        RECT 651.000 520.950 655.050 521.550 ;
        RECT 659.400 518.700 660.600 523.800 ;
        RECT 662.100 522.000 663.900 523.800 ;
        RECT 668.550 523.050 669.450 526.950 ;
        RECT 674.100 526.050 675.900 527.850 ;
        RECT 679.950 526.050 681.150 539.400 ;
        RECT 701.850 526.050 703.050 539.400 ;
        RECT 706.500 533.400 708.300 546.000 ;
        RECT 716.400 533.400 718.200 546.000 ;
        RECT 720.900 533.400 724.200 545.400 ;
        RECT 726.900 533.400 728.700 546.000 ;
        RECT 740.400 534.300 742.200 545.400 ;
        RECT 747.900 544.050 749.700 545.400 ;
        RECT 747.900 541.950 751.050 544.050 ;
        RECT 740.400 533.400 744.900 534.300 ;
        RECT 747.900 533.400 749.700 541.950 ;
        RECT 755.400 534.600 757.200 545.400 ;
        RECT 767.400 539.400 769.200 546.000 ;
        RECT 770.400 539.400 772.200 545.400 ;
        RECT 782.400 539.400 784.200 546.000 ;
        RECT 785.400 539.400 787.200 545.400 ;
        RECT 788.400 539.400 790.200 546.000 ;
        RECT 800.400 539.400 802.200 546.000 ;
        RECT 803.400 539.400 805.200 545.400 ;
        RECT 707.100 526.050 708.900 527.850 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 682.950 523.950 685.050 526.050 ;
        RECT 697.950 523.950 700.050 526.050 ;
        RECT 700.950 523.950 703.050 526.050 ;
        RECT 703.950 523.950 706.050 526.050 ;
        RECT 706.950 523.950 709.050 526.050 ;
        RECT 716.100 525.900 717.900 527.700 ;
        RECT 722.100 525.900 723.300 533.400 ;
        RECT 742.800 531.300 744.900 533.400 ;
        RECT 748.500 531.900 749.700 533.400 ;
        RECT 752.400 533.400 757.200 534.600 ;
        RECT 752.400 532.500 754.500 533.400 ;
        RECT 748.500 531.000 750.000 531.900 ;
        RECT 745.950 529.500 748.050 529.800 ;
        RECT 735.000 528.450 739.050 529.050 ;
        RECT 728.100 525.900 729.900 527.700 ;
        RECT 734.550 526.950 739.050 528.450 ;
        RECT 744.300 527.700 748.050 529.500 ;
        RECT 749.100 528.900 750.000 531.000 ;
        RECT 668.550 521.550 673.050 523.050 ;
        RECT 677.100 522.150 678.900 523.950 ;
        RECT 669.000 520.950 673.050 521.550 ;
        RECT 680.850 519.750 682.050 523.950 ;
        RECT 683.100 522.150 684.900 523.950 ;
        RECT 698.100 522.150 699.900 523.950 ;
        RECT 680.850 518.700 684.600 519.750 ;
        RECT 659.400 517.800 663.600 518.700 ;
        RECT 626.850 515.550 628.650 516.300 ;
        RECT 640.950 515.700 643.050 516.600 ;
        RECT 626.850 514.500 631.800 515.550 ;
        RECT 621.000 513.600 622.050 514.500 ;
        RECT 630.750 513.600 631.800 514.500 ;
        RECT 639.300 514.500 643.050 515.700 ;
        RECT 639.300 513.600 640.350 514.500 ;
        RECT 618.150 510.000 619.950 513.600 ;
        RECT 621.000 512.700 624.750 513.600 ;
        RECT 622.950 510.600 624.750 512.700 ;
        RECT 627.450 510.000 629.250 513.600 ;
        RECT 630.750 510.600 632.550 513.600 ;
        RECT 634.350 510.000 636.150 513.600 ;
        RECT 638.550 510.600 640.350 513.600 ;
        RECT 643.350 510.000 645.150 513.600 ;
        RECT 646.650 510.600 648.450 516.600 ;
        RECT 656.700 510.000 658.500 516.600 ;
        RECT 661.800 510.600 663.600 517.800 ;
        RECT 674.400 515.700 682.200 517.050 ;
        RECT 674.400 510.600 676.200 515.700 ;
        RECT 677.400 510.000 679.200 514.800 ;
        RECT 680.400 510.600 682.200 515.700 ;
        RECT 683.400 516.600 684.600 518.700 ;
        RECT 685.950 519.450 688.050 520.050 ;
        RECT 691.950 519.450 694.050 519.900 ;
        RECT 700.950 519.750 702.150 523.950 ;
        RECT 704.100 522.150 705.900 523.950 ;
        RECT 715.950 523.800 718.050 525.900 ;
        RECT 718.950 523.800 721.050 525.900 ;
        RECT 721.950 523.800 724.050 525.900 ;
        RECT 724.950 523.800 727.050 525.900 ;
        RECT 727.950 523.800 730.050 525.900 ;
        RECT 719.100 522.000 720.900 523.800 ;
        RECT 721.950 521.400 723.000 523.800 ;
        RECT 725.100 522.000 726.900 523.800 ;
        RECT 734.550 523.050 735.450 526.950 ;
        RECT 748.950 526.800 751.050 528.900 ;
        RECT 756.000 528.450 760.050 529.050 ;
        RECT 755.550 527.700 760.050 528.450 ;
        RECT 755.100 526.950 760.050 527.700 ;
        RECT 745.500 525.900 747.300 526.500 ;
        RECT 739.950 524.700 747.300 525.900 ;
        RECT 748.200 525.900 750.600 526.800 ;
        RECT 755.100 525.900 756.900 526.950 ;
        RECT 767.100 526.050 768.900 527.850 ;
        RECT 770.400 526.050 771.600 539.400 ;
        RECT 739.950 523.800 742.050 524.700 ;
        RECT 730.950 521.550 735.450 523.050 ;
        RECT 740.250 522.000 742.050 523.800 ;
        RECT 685.950 518.550 694.050 519.450 ;
        RECT 685.950 517.950 688.050 518.550 ;
        RECT 691.950 517.800 694.050 518.550 ;
        RECT 698.400 518.700 702.150 519.750 ;
        RECT 722.100 519.300 723.300 521.400 ;
        RECT 730.950 520.950 735.000 521.550 ;
        RECT 745.500 521.400 747.300 523.200 ;
        RECT 745.200 519.300 747.300 521.400 ;
        RECT 698.400 516.600 699.600 518.700 ;
        RECT 722.100 518.100 726.600 519.300 ;
        RECT 683.400 510.600 685.200 516.600 ;
        RECT 697.800 510.600 699.600 516.600 ;
        RECT 700.800 515.700 708.600 517.050 ;
        RECT 700.800 510.600 702.600 515.700 ;
        RECT 703.800 510.000 705.600 514.800 ;
        RECT 706.800 510.600 708.600 515.700 ;
        RECT 716.400 516.000 724.200 516.900 ;
        RECT 725.700 516.600 726.600 518.100 ;
        RECT 741.000 518.400 747.300 519.300 ;
        RECT 748.200 520.200 749.250 525.900 ;
        RECT 750.600 523.200 752.400 525.000 ;
        RECT 754.950 523.800 757.050 525.900 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 769.950 523.950 772.050 526.050 ;
        RECT 785.400 525.900 786.600 539.400 ;
        RECT 800.100 526.050 801.900 527.850 ;
        RECT 803.400 526.050 804.600 539.400 ;
        RECT 815.400 534.300 817.200 545.400 ;
        RECT 815.400 533.400 819.900 534.300 ;
        RECT 822.900 533.400 824.700 545.400 ;
        RECT 830.400 534.600 832.200 545.400 ;
        RECT 842.400 539.400 844.200 546.000 ;
        RECT 845.400 539.400 847.200 545.400 ;
        RECT 848.400 540.000 850.200 546.000 ;
        RECT 845.700 539.100 847.200 539.400 ;
        RECT 851.400 539.400 853.200 545.400 ;
        RECT 851.400 539.100 852.300 539.400 ;
        RECT 845.700 538.200 852.300 539.100 ;
        RECT 817.800 531.300 819.900 533.400 ;
        RECT 823.500 531.900 824.700 533.400 ;
        RECT 827.400 533.400 832.200 534.600 ;
        RECT 827.400 532.500 829.500 533.400 ;
        RECT 823.500 531.000 825.000 531.900 ;
        RECT 820.950 529.500 823.050 529.800 ;
        RECT 819.300 527.700 823.050 529.500 ;
        RECT 824.100 528.900 825.000 531.000 ;
        RECT 823.950 526.800 826.050 528.900 ;
        RECT 838.950 528.450 841.050 529.050 ;
        RECT 830.550 527.700 841.050 528.450 ;
        RECT 830.100 527.550 841.050 527.700 ;
        RECT 750.150 521.100 752.250 523.200 ;
        RECT 741.000 516.600 742.200 518.400 ;
        RECT 748.200 518.100 751.050 520.200 ;
        RECT 748.200 516.600 749.400 518.100 ;
        RECT 752.400 517.500 754.500 518.700 ;
        RECT 752.400 516.600 757.200 517.500 ;
        RECT 716.400 510.600 718.200 516.000 ;
        RECT 719.400 510.000 721.200 515.100 ;
        RECT 722.400 511.500 724.200 516.000 ;
        RECT 725.400 512.400 727.200 516.600 ;
        RECT 728.400 511.500 730.200 516.600 ;
        RECT 722.400 510.600 730.200 511.500 ;
        RECT 740.400 510.600 742.200 516.600 ;
        RECT 747.900 510.600 749.700 516.600 ;
        RECT 755.400 510.600 757.200 516.600 ;
        RECT 770.400 513.600 771.600 523.950 ;
        RECT 781.950 523.800 784.050 525.900 ;
        RECT 784.950 523.800 787.050 525.900 ;
        RECT 787.950 523.800 790.050 525.900 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 820.500 525.900 822.300 526.500 ;
        RECT 814.950 524.700 822.300 525.900 ;
        RECT 823.200 525.900 825.600 526.800 ;
        RECT 830.100 525.900 831.900 527.550 ;
        RECT 838.950 526.950 841.050 527.550 ;
        RECT 845.100 525.900 846.900 527.700 ;
        RECT 851.400 525.900 852.300 538.200 ;
        RECT 856.950 529.950 859.050 532.050 ;
        RECT 782.100 522.000 783.900 523.800 ;
        RECT 785.400 518.700 786.600 523.800 ;
        RECT 788.100 522.000 789.900 523.800 ;
        RECT 785.400 517.800 789.600 518.700 ;
        RECT 767.400 510.000 769.200 513.600 ;
        RECT 770.400 510.600 772.200 513.600 ;
        RECT 782.700 510.000 784.500 516.600 ;
        RECT 787.800 510.600 789.600 517.800 ;
        RECT 803.400 513.600 804.600 523.950 ;
        RECT 814.950 523.800 817.050 524.700 ;
        RECT 815.250 522.000 817.050 523.800 ;
        RECT 820.500 521.400 822.300 523.200 ;
        RECT 820.200 519.300 822.300 521.400 ;
        RECT 816.000 518.400 822.300 519.300 ;
        RECT 823.200 520.200 824.250 525.900 ;
        RECT 825.600 523.200 827.400 525.000 ;
        RECT 829.950 523.800 832.050 525.900 ;
        RECT 841.950 523.800 844.050 525.900 ;
        RECT 844.950 523.800 847.050 525.900 ;
        RECT 847.950 523.800 850.050 525.900 ;
        RECT 850.950 523.800 853.050 525.900 ;
        RECT 825.150 521.100 827.250 523.200 ;
        RECT 842.100 522.000 843.900 523.800 ;
        RECT 848.100 522.000 849.900 523.800 ;
        RECT 851.400 520.200 852.300 523.800 ;
        RECT 816.000 516.600 817.200 518.400 ;
        RECT 823.200 518.100 826.050 520.200 ;
        RECT 823.200 516.600 824.400 518.100 ;
        RECT 827.400 517.500 829.500 518.700 ;
        RECT 827.400 516.600 832.200 517.500 ;
        RECT 800.400 510.000 802.200 513.600 ;
        RECT 803.400 510.600 805.200 513.600 ;
        RECT 815.400 510.600 817.200 516.600 ;
        RECT 822.900 510.600 824.700 516.600 ;
        RECT 830.400 510.600 832.200 516.600 ;
        RECT 842.400 510.000 844.200 519.600 ;
        RECT 849.000 519.000 852.300 520.200 ;
        RECT 849.000 510.600 850.800 519.000 ;
        RECT 857.550 516.900 858.450 529.950 ;
        RECT 856.950 514.800 859.050 516.900 ;
        RECT 10.800 503.400 12.600 506.400 ;
        RECT 13.800 503.400 15.600 507.000 ;
        RECT 25.800 503.400 27.600 506.400 ;
        RECT 28.800 503.400 30.600 507.000 ;
        RECT 11.400 493.050 12.600 503.400 ;
        RECT 26.400 493.050 27.600 503.400 ;
        RECT 40.800 500.400 42.600 506.400 ;
        RECT 28.950 498.450 31.050 499.050 ;
        RECT 34.950 498.450 37.050 499.050 ;
        RECT 28.950 497.550 37.050 498.450 ;
        RECT 28.950 496.950 31.050 497.550 ;
        RECT 34.950 496.950 37.050 497.550 ;
        RECT 41.400 498.300 42.600 500.400 ;
        RECT 43.800 501.300 45.600 506.400 ;
        RECT 46.800 502.200 48.600 507.000 ;
        RECT 49.800 501.300 51.600 506.400 ;
        RECT 62.700 503.400 64.500 507.000 ;
        RECT 65.700 501.600 67.500 506.400 ;
        RECT 43.800 499.950 51.600 501.300 ;
        RECT 62.400 500.400 67.500 501.600 ;
        RECT 70.200 500.400 72.000 507.000 ;
        RECT 82.800 500.400 84.600 506.400 ;
        RECT 41.400 497.250 45.150 498.300 ;
        RECT 41.100 493.050 42.900 494.850 ;
        RECT 43.950 493.050 45.150 497.250 ;
        RECT 47.100 493.050 48.900 494.850 ;
        RECT 62.400 493.200 63.300 500.400 ;
        RECT 83.400 498.300 84.600 500.400 ;
        RECT 85.800 501.300 87.600 506.400 ;
        RECT 88.800 502.200 90.600 507.000 ;
        RECT 91.800 501.300 93.600 506.400 ;
        RECT 103.800 503.400 105.600 507.000 ;
        RECT 106.800 503.400 108.600 506.400 ;
        RECT 109.800 503.400 111.600 507.000 ;
        RECT 121.800 503.400 123.600 506.400 ;
        RECT 124.800 503.400 126.600 507.000 ;
        RECT 85.800 499.950 93.600 501.300 ;
        RECT 83.400 497.250 87.150 498.300 ;
        RECT 65.100 493.200 66.900 495.000 ;
        RECT 71.100 493.200 72.900 495.000 ;
        RECT 10.950 490.950 13.050 493.050 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 25.950 490.950 28.050 493.050 ;
        RECT 28.950 490.950 31.050 493.050 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 43.950 490.950 46.050 493.050 ;
        RECT 46.950 490.950 49.050 493.050 ;
        RECT 49.950 490.950 52.050 493.050 ;
        RECT 61.950 491.100 64.050 493.200 ;
        RECT 64.950 491.100 67.050 493.200 ;
        RECT 67.950 491.100 70.050 493.200 ;
        RECT 70.950 491.100 73.050 493.200 ;
        RECT 83.100 493.050 84.900 494.850 ;
        RECT 85.950 493.050 87.150 497.250 ;
        RECT 94.950 495.450 99.000 496.050 ;
        RECT 89.100 493.050 90.900 494.850 ;
        RECT 94.950 493.950 99.450 495.450 ;
        RECT 11.400 477.600 12.600 490.950 ;
        RECT 14.100 489.150 15.900 490.950 ;
        RECT 26.400 477.600 27.600 490.950 ;
        RECT 29.100 489.150 30.900 490.950 ;
        RECT 44.850 477.600 46.050 490.950 ;
        RECT 50.100 489.150 51.900 490.950 ;
        RECT 62.400 483.600 63.300 491.100 ;
        RECT 68.100 489.300 69.900 491.100 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 85.950 490.950 88.050 493.050 ;
        RECT 88.950 490.950 91.050 493.050 ;
        RECT 91.950 490.950 94.050 493.050 ;
        RECT 10.800 471.600 12.600 477.600 ;
        RECT 13.800 471.000 15.600 477.600 ;
        RECT 25.800 471.600 27.600 477.600 ;
        RECT 28.800 471.000 30.600 477.600 ;
        RECT 41.400 471.000 43.200 477.600 ;
        RECT 44.400 471.600 46.200 477.600 ;
        RECT 49.500 471.000 51.300 483.600 ;
        RECT 61.800 471.600 63.600 483.600 ;
        RECT 64.800 482.700 72.600 483.600 ;
        RECT 64.800 471.600 66.600 482.700 ;
        RECT 67.800 471.000 69.600 481.800 ;
        RECT 70.800 471.600 72.600 482.700 ;
        RECT 86.850 477.600 88.050 490.950 ;
        RECT 92.100 489.150 93.900 490.950 ;
        RECT 98.550 490.050 99.450 493.950 ;
        RECT 107.400 493.050 108.300 503.400 ;
        RECT 122.400 493.050 123.600 503.400 ;
        RECT 139.500 500.400 141.300 507.000 ;
        RECT 144.000 500.400 145.800 506.400 ;
        RECT 148.500 500.400 150.300 507.000 ;
        RECT 158.700 500.400 160.500 507.000 ;
        RECT 137.100 493.200 138.900 495.000 ;
        RECT 144.000 493.200 145.050 500.400 ;
        RECT 163.800 499.200 165.600 506.400 ;
        RECT 176.700 500.400 178.500 507.000 ;
        RECT 181.800 499.200 183.600 506.400 ;
        RECT 161.400 498.300 165.600 499.200 ;
        RECT 179.400 498.300 183.600 499.200 ;
        RECT 197.400 499.200 199.200 506.400 ;
        RECT 202.500 500.400 204.300 507.000 ;
        RECT 214.800 500.400 216.600 506.400 ;
        RECT 222.600 501.000 224.400 506.400 ;
        RECT 214.800 499.500 219.300 500.400 ;
        RECT 197.400 498.300 201.600 499.200 ;
        RECT 149.100 493.200 150.900 495.000 ;
        RECT 158.100 493.200 159.900 495.000 ;
        RECT 161.400 493.200 162.600 498.300 ;
        RECT 164.100 493.200 165.900 495.000 ;
        RECT 176.100 493.200 177.900 495.000 ;
        RECT 179.400 493.200 180.600 498.300 ;
        RECT 192.000 495.450 196.050 496.050 ;
        RECT 182.100 493.200 183.900 495.000 ;
        RECT 191.550 493.950 196.050 495.450 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 121.950 490.950 124.050 493.050 ;
        RECT 124.950 490.950 127.050 493.050 ;
        RECT 136.950 491.100 139.050 493.200 ;
        RECT 139.950 491.100 142.050 493.200 ;
        RECT 142.950 491.100 145.050 493.200 ;
        RECT 145.950 491.100 148.050 493.200 ;
        RECT 148.950 491.100 151.050 493.200 ;
        RECT 157.950 491.100 160.050 493.200 ;
        RECT 160.950 491.100 163.050 493.200 ;
        RECT 163.950 491.100 166.050 493.200 ;
        RECT 175.950 491.100 178.050 493.200 ;
        RECT 178.950 491.100 181.050 493.200 ;
        RECT 181.950 491.100 184.050 493.200 ;
        RECT 94.950 488.550 99.450 490.050 ;
        RECT 104.100 489.150 105.900 490.950 ;
        RECT 94.950 487.950 99.000 488.550 ;
        RECT 107.400 483.600 108.300 490.950 ;
        RECT 110.100 489.150 111.900 490.950 ;
        RECT 83.400 471.000 85.200 477.600 ;
        RECT 86.400 471.600 88.200 477.600 ;
        RECT 91.500 471.000 93.300 483.600 ;
        RECT 104.700 482.400 108.300 483.600 ;
        RECT 104.700 471.600 106.500 482.400 ;
        RECT 109.800 471.000 111.600 483.600 ;
        RECT 122.400 477.600 123.600 490.950 ;
        RECT 125.100 489.150 126.900 490.950 ;
        RECT 140.100 489.300 141.900 491.100 ;
        RECT 144.000 485.400 144.900 491.100 ;
        RECT 146.100 489.300 147.900 491.100 ;
        RECT 148.950 489.450 151.050 490.050 ;
        RECT 157.950 489.450 160.050 490.050 ;
        RECT 148.950 488.550 160.050 489.450 ;
        RECT 148.950 487.950 151.050 488.550 ;
        RECT 157.950 487.950 160.050 488.550 ;
        RECT 139.800 484.500 144.900 485.400 ;
        RECT 121.800 471.600 123.600 477.600 ;
        RECT 124.800 471.000 126.600 477.600 ;
        RECT 136.800 472.500 138.600 483.600 ;
        RECT 139.800 473.400 141.600 484.500 ;
        RECT 142.800 482.400 150.600 483.300 ;
        RECT 142.800 472.500 144.600 482.400 ;
        RECT 136.800 471.600 144.600 472.500 ;
        RECT 145.800 471.000 147.600 481.500 ;
        RECT 148.800 471.600 150.600 482.400 ;
        RECT 161.400 477.600 162.600 491.100 ;
        RECT 163.950 489.450 166.050 490.050 ;
        RECT 169.950 489.450 172.050 490.050 ;
        RECT 163.950 488.550 172.050 489.450 ;
        RECT 163.950 487.950 166.050 488.550 ;
        RECT 169.950 487.950 172.050 488.550 ;
        RECT 179.400 477.600 180.600 491.100 ;
        RECT 191.550 489.900 192.450 493.950 ;
        RECT 197.100 493.200 198.900 495.000 ;
        RECT 200.400 493.200 201.600 498.300 ;
        RECT 217.200 497.100 219.300 499.500 ;
        RECT 222.750 498.900 223.650 501.000 ;
        RECT 229.800 500.400 231.600 506.400 ;
        RECT 230.100 499.500 231.600 500.400 ;
        RECT 239.400 501.300 241.200 506.400 ;
        RECT 242.400 502.200 244.200 507.000 ;
        RECT 245.400 501.300 247.200 506.400 ;
        RECT 239.400 499.950 247.200 501.300 ;
        RECT 248.400 500.400 250.200 506.400 ;
        RECT 220.650 496.800 223.650 498.900 ;
        RECT 227.250 498.000 231.600 499.500 ;
        RECT 248.400 498.300 249.600 500.400 ;
        RECT 205.950 495.450 210.000 496.050 ;
        RECT 203.100 493.200 204.900 495.000 ;
        RECT 205.950 493.950 210.450 495.450 ;
        RECT 196.950 491.100 199.050 493.200 ;
        RECT 199.950 491.100 202.050 493.200 ;
        RECT 202.950 491.100 205.050 493.200 ;
        RECT 190.950 487.800 193.050 489.900 ;
        RECT 200.400 477.600 201.600 491.100 ;
        RECT 209.550 490.050 210.450 493.950 ;
        RECT 214.950 491.100 217.050 493.200 ;
        RECT 219.750 492.900 221.850 495.000 ;
        RECT 219.900 491.100 221.700 492.900 ;
        RECT 205.950 488.550 210.450 490.050 ;
        RECT 215.100 489.300 216.900 491.100 ;
        RECT 222.750 490.200 223.650 496.800 ;
        RECT 224.550 495.900 226.350 497.700 ;
        RECT 227.250 497.400 229.350 498.000 ;
        RECT 245.850 497.250 249.600 498.300 ;
        RECT 260.400 497.400 262.200 507.000 ;
        RECT 267.000 498.000 268.800 506.400 ;
        RECT 283.800 503.400 285.600 507.000 ;
        RECT 286.800 503.400 288.600 506.400 ;
        RECT 289.800 503.400 291.600 507.000 ;
        RECT 271.950 501.450 274.050 501.900 ;
        RECT 280.950 501.450 283.050 502.050 ;
        RECT 271.950 500.550 283.050 501.450 ;
        RECT 271.950 499.800 274.050 500.550 ;
        RECT 280.950 499.950 283.050 500.550 ;
        RECT 274.950 498.450 277.050 499.050 ;
        RECT 283.950 498.450 286.050 498.900 ;
        RECT 224.700 495.000 226.800 495.900 ;
        RECT 224.700 493.800 231.750 495.000 ;
        RECT 229.950 493.200 231.750 493.800 ;
        RECT 224.700 490.800 226.800 492.900 ;
        RECT 229.950 491.100 232.050 493.200 ;
        RECT 242.100 493.050 243.900 494.850 ;
        RECT 245.850 493.050 247.050 497.250 ;
        RECT 267.000 496.800 270.300 498.000 ;
        RECT 274.950 497.550 286.050 498.450 ;
        RECT 274.950 496.950 277.050 497.550 ;
        RECT 283.950 496.800 286.050 497.550 ;
        RECT 255.000 495.450 259.050 496.050 ;
        RECT 248.100 493.050 249.900 494.850 ;
        RECT 254.550 493.950 259.050 495.450 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 241.950 490.950 244.050 493.050 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 247.950 490.950 250.050 493.050 ;
        RECT 220.650 488.700 223.650 490.200 ;
        RECT 225.000 489.000 226.800 490.800 ;
        RECT 239.100 489.150 240.900 490.950 ;
        RECT 205.950 487.950 210.000 488.550 ;
        RECT 220.650 488.100 222.750 488.700 ;
        RECT 217.800 483.600 219.900 484.500 ;
        RECT 214.800 482.400 219.900 483.600 ;
        RECT 220.800 483.600 222.000 488.100 ;
        RECT 223.650 485.700 225.450 487.800 ;
        RECT 223.650 484.800 228.900 485.700 ;
        RECT 226.800 483.900 228.900 484.800 ;
        RECT 220.800 482.700 224.100 483.600 ;
        RECT 226.800 482.700 231.600 483.900 ;
        RECT 158.400 471.000 160.200 477.600 ;
        RECT 161.400 471.600 163.200 477.600 ;
        RECT 164.400 471.000 166.200 477.600 ;
        RECT 176.400 471.000 178.200 477.600 ;
        RECT 179.400 471.600 181.200 477.600 ;
        RECT 182.400 471.000 184.200 477.600 ;
        RECT 196.800 471.000 198.600 477.600 ;
        RECT 199.800 471.600 201.600 477.600 ;
        RECT 202.800 471.000 204.600 477.600 ;
        RECT 214.800 471.600 216.600 482.400 ;
        RECT 222.300 471.600 224.100 482.700 ;
        RECT 229.800 471.600 231.600 482.700 ;
        RECT 239.700 471.000 241.500 483.600 ;
        RECT 244.950 477.600 246.150 490.950 ;
        RECT 254.550 489.450 255.450 493.950 ;
        RECT 260.100 493.200 261.900 495.000 ;
        RECT 266.100 493.200 267.900 495.000 ;
        RECT 269.400 493.200 270.300 496.800 ;
        RECT 259.950 491.100 262.050 493.200 ;
        RECT 262.950 491.100 265.050 493.200 ;
        RECT 265.950 491.100 268.050 493.200 ;
        RECT 268.950 491.100 271.050 493.200 ;
        RECT 287.400 493.050 288.300 503.400 ;
        RECT 299.400 497.400 301.200 507.000 ;
        RECT 306.000 498.000 307.800 506.400 ;
        RECT 322.800 500.400 324.600 506.400 ;
        RECT 323.400 498.300 324.600 500.400 ;
        RECT 325.800 501.300 327.600 506.400 ;
        RECT 328.800 502.200 330.600 507.000 ;
        RECT 331.800 501.300 333.600 506.400 ;
        RECT 325.800 499.950 333.600 501.300 ;
        RECT 344.400 499.200 346.200 506.400 ;
        RECT 349.500 500.400 351.300 507.000 ;
        RECT 363.300 502.200 365.100 506.400 ;
        RECT 362.400 500.400 365.100 502.200 ;
        RECT 366.300 500.400 368.100 507.000 ;
        RECT 306.000 496.800 309.300 498.000 ;
        RECT 323.400 497.250 327.150 498.300 ;
        RECT 299.100 493.200 300.900 495.000 ;
        RECT 305.100 493.200 306.900 495.000 ;
        RECT 308.400 493.200 309.300 496.800 ;
        RECT 254.550 488.550 261.450 489.450 ;
        RECT 263.100 489.300 264.900 491.100 ;
        RECT 260.550 486.450 261.450 488.550 ;
        RECT 265.950 486.450 268.050 487.050 ;
        RECT 260.550 485.550 268.050 486.450 ;
        RECT 265.950 484.950 268.050 485.550 ;
        RECT 269.400 478.800 270.300 491.100 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 286.950 490.950 289.050 493.050 ;
        RECT 289.950 490.950 292.050 493.050 ;
        RECT 298.950 491.100 301.050 493.200 ;
        RECT 301.950 491.100 304.050 493.200 ;
        RECT 304.950 491.100 307.050 493.200 ;
        RECT 307.950 491.100 310.050 493.200 ;
        RECT 323.100 493.050 324.900 494.850 ;
        RECT 325.950 493.050 327.150 497.250 ;
        RECT 337.950 496.950 340.050 499.050 ;
        RECT 344.400 498.300 348.600 499.200 ;
        RECT 329.100 493.050 330.900 494.850 ;
        RECT 284.100 489.150 285.900 490.950 ;
        RECT 287.400 483.600 288.300 490.950 ;
        RECT 290.100 489.150 291.900 490.950 ;
        RECT 302.100 489.300 303.900 491.100 ;
        RECT 292.950 486.450 295.050 487.050 ;
        RECT 304.950 486.450 307.050 487.050 ;
        RECT 292.950 485.550 307.050 486.450 ;
        RECT 292.950 484.950 295.050 485.550 ;
        RECT 304.950 484.950 307.050 485.550 ;
        RECT 263.700 477.900 270.300 478.800 ;
        RECT 263.700 477.600 265.200 477.900 ;
        RECT 244.800 471.600 246.600 477.600 ;
        RECT 247.800 471.000 249.600 477.600 ;
        RECT 260.400 471.000 262.200 477.600 ;
        RECT 263.400 471.600 265.200 477.600 ;
        RECT 269.400 477.600 270.300 477.900 ;
        RECT 284.700 482.400 288.300 483.600 ;
        RECT 266.400 471.000 268.200 477.000 ;
        RECT 269.400 471.600 271.200 477.600 ;
        RECT 284.700 471.600 286.500 482.400 ;
        RECT 289.800 471.000 291.600 483.600 ;
        RECT 308.400 478.800 309.300 491.100 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 325.950 490.950 328.050 493.050 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 331.950 490.950 334.050 493.050 ;
        RECT 316.950 483.450 321.000 484.050 ;
        RECT 316.950 483.000 321.450 483.450 ;
        RECT 316.950 481.950 322.050 483.000 ;
        RECT 310.950 480.450 313.050 481.050 ;
        RECT 316.800 480.450 318.900 480.900 ;
        RECT 310.950 479.550 318.900 480.450 ;
        RECT 310.950 478.950 313.050 479.550 ;
        RECT 316.800 478.800 318.900 479.550 ;
        RECT 319.950 478.800 322.050 481.950 ;
        RECT 302.700 477.900 309.300 478.800 ;
        RECT 302.700 477.600 304.200 477.900 ;
        RECT 299.400 471.000 301.200 477.600 ;
        RECT 302.400 471.600 304.200 477.600 ;
        RECT 308.400 477.600 309.300 477.900 ;
        RECT 326.850 477.600 328.050 490.950 ;
        RECT 332.100 489.150 333.900 490.950 ;
        RECT 338.550 490.050 339.450 496.950 ;
        RECT 344.100 493.200 345.900 495.000 ;
        RECT 347.400 493.200 348.600 498.300 ;
        RECT 352.950 495.450 357.000 496.050 ;
        RECT 350.100 493.200 351.900 495.000 ;
        RECT 352.950 493.950 357.450 495.450 ;
        RECT 343.950 491.100 346.050 493.200 ;
        RECT 346.950 491.100 349.050 493.200 ;
        RECT 349.950 491.100 352.050 493.200 ;
        RECT 334.950 488.550 339.450 490.050 ;
        RECT 334.950 487.950 339.000 488.550 ;
        RECT 305.400 471.000 307.200 477.000 ;
        RECT 308.400 471.600 310.200 477.600 ;
        RECT 323.400 471.000 325.200 477.600 ;
        RECT 326.400 471.600 328.200 477.600 ;
        RECT 331.500 471.000 333.300 483.600 ;
        RECT 347.400 477.600 348.600 491.100 ;
        RECT 356.550 490.050 357.450 493.950 ;
        RECT 362.400 493.200 363.300 500.400 ;
        RECT 365.100 498.600 366.900 499.500 ;
        RECT 370.800 498.600 372.600 506.400 ;
        RECT 380.700 500.400 382.500 507.000 ;
        RECT 385.800 499.200 387.600 506.400 ;
        RECT 365.100 497.700 372.600 498.600 ;
        RECT 383.400 498.300 387.600 499.200 ;
        RECT 401.400 499.200 403.200 506.400 ;
        RECT 406.500 500.400 408.300 507.000 ;
        RECT 416.400 501.300 418.200 506.400 ;
        RECT 419.400 502.200 421.200 507.000 ;
        RECT 422.400 501.300 424.200 506.400 ;
        RECT 416.400 499.950 424.200 501.300 ;
        RECT 425.400 500.400 427.200 506.400 ;
        RECT 438.000 500.400 439.800 507.000 ;
        RECT 442.500 501.600 444.300 506.400 ;
        RECT 445.500 503.400 447.300 507.000 ;
        RECT 442.500 500.400 447.600 501.600 ;
        RECT 401.400 498.300 405.600 499.200 ;
        RECT 425.400 498.300 426.600 500.400 ;
        RECT 361.950 491.100 364.050 493.200 ;
        RECT 364.950 491.100 367.050 493.200 ;
        RECT 356.550 488.550 361.050 490.050 ;
        RECT 357.000 487.950 361.050 488.550 ;
        RECT 362.400 483.600 363.300 491.100 ;
        RECT 365.100 489.300 366.900 491.100 ;
        RECT 343.800 471.000 345.600 477.600 ;
        RECT 346.800 471.600 348.600 477.600 ;
        RECT 349.800 471.000 351.600 477.600 ;
        RECT 361.800 471.600 363.600 483.600 ;
        RECT 368.700 477.600 369.600 497.700 ;
        RECT 371.100 493.200 372.900 495.000 ;
        RECT 380.100 493.200 381.900 495.000 ;
        RECT 383.400 493.200 384.600 498.300 ;
        RECT 386.100 493.200 387.900 495.000 ;
        RECT 401.100 493.200 402.900 495.000 ;
        RECT 404.400 493.200 405.600 498.300 ;
        RECT 422.850 497.250 426.600 498.300 ;
        RECT 407.100 493.200 408.900 495.000 ;
        RECT 370.950 491.100 373.050 493.200 ;
        RECT 379.950 491.100 382.050 493.200 ;
        RECT 382.950 491.100 385.050 493.200 ;
        RECT 385.950 491.100 388.050 493.200 ;
        RECT 400.950 491.100 403.050 493.200 ;
        RECT 403.950 491.100 406.050 493.200 ;
        RECT 406.950 491.100 409.050 493.200 ;
        RECT 419.100 493.050 420.900 494.850 ;
        RECT 422.850 493.050 424.050 497.250 ;
        RECT 425.100 493.050 426.900 494.850 ;
        RECT 437.100 493.200 438.900 495.000 ;
        RECT 443.100 493.200 444.900 495.000 ;
        RECT 446.700 493.200 447.600 500.400 ;
        RECT 452.550 500.400 454.350 506.400 ;
        RECT 455.850 503.400 457.650 507.000 ;
        RECT 460.650 503.400 462.450 506.400 ;
        RECT 464.850 503.400 466.650 507.000 ;
        RECT 468.450 503.400 470.250 506.400 ;
        RECT 471.750 503.400 473.550 507.000 ;
        RECT 476.250 504.300 478.050 506.400 ;
        RECT 476.250 503.400 480.000 504.300 ;
        RECT 481.050 503.400 482.850 507.000 ;
        RECT 460.650 502.500 461.700 503.400 ;
        RECT 457.950 501.300 461.700 502.500 ;
        RECT 469.200 502.500 470.250 503.400 ;
        RECT 478.950 502.500 480.000 503.400 ;
        RECT 469.200 501.450 474.150 502.500 ;
        RECT 457.950 500.400 460.050 501.300 ;
        RECT 472.350 500.700 474.150 501.450 ;
        RECT 383.400 477.600 384.600 491.100 ;
        RECT 404.400 477.600 405.600 491.100 ;
        RECT 415.950 490.950 418.050 493.050 ;
        RECT 418.950 490.950 421.050 493.050 ;
        RECT 421.950 490.950 424.050 493.050 ;
        RECT 424.950 490.950 427.050 493.050 ;
        RECT 436.950 491.100 439.050 493.200 ;
        RECT 439.950 491.100 442.050 493.200 ;
        RECT 442.950 491.100 445.050 493.200 ;
        RECT 445.950 491.100 448.050 493.200 ;
        RECT 452.550 493.050 453.750 500.400 ;
        RECT 475.650 499.800 477.450 501.600 ;
        RECT 478.950 500.400 481.050 502.500 ;
        RECT 484.050 500.400 485.850 506.400 ;
        RECT 494.700 500.400 496.500 507.000 ;
        RECT 465.150 498.000 466.950 498.600 ;
        RECT 476.100 498.000 477.150 499.800 ;
        RECT 465.150 496.800 477.150 498.000 ;
        RECT 452.550 491.250 458.850 493.050 ;
        RECT 416.100 489.150 417.900 490.950 ;
        RECT 364.800 471.000 366.600 477.600 ;
        RECT 367.800 471.600 369.600 477.600 ;
        RECT 370.800 471.000 372.600 477.600 ;
        RECT 380.400 471.000 382.200 477.600 ;
        RECT 383.400 471.600 385.200 477.600 ;
        RECT 386.400 471.000 388.200 477.600 ;
        RECT 400.800 471.000 402.600 477.600 ;
        RECT 403.800 471.600 405.600 477.600 ;
        RECT 406.800 471.000 408.600 477.600 ;
        RECT 416.700 471.000 418.500 483.600 ;
        RECT 421.950 477.600 423.150 490.950 ;
        RECT 440.100 489.300 441.900 491.100 ;
        RECT 446.700 483.600 447.600 491.100 ;
        RECT 452.550 490.950 457.050 491.250 ;
        RECT 452.550 483.600 453.750 490.950 ;
        RECT 454.950 485.400 456.750 487.200 ;
        RECT 455.850 484.200 460.050 485.400 ;
        RECT 465.150 484.200 466.050 496.800 ;
        RECT 476.100 495.600 483.000 496.800 ;
        RECT 476.100 495.000 477.900 495.600 ;
        RECT 482.100 494.850 483.000 495.600 ;
        RECT 479.100 493.800 480.900 494.400 ;
        RECT 472.950 492.600 480.900 493.800 ;
        RECT 482.100 493.050 483.900 494.850 ;
        RECT 472.950 490.950 475.050 492.600 ;
        RECT 481.950 490.950 484.050 493.050 ;
        RECT 474.750 485.700 476.550 486.000 ;
        RECT 484.950 485.700 485.850 500.400 ;
        RECT 499.800 499.200 501.600 506.400 ;
        RECT 514.800 500.400 516.600 506.400 ;
        RECT 497.400 498.300 501.600 499.200 ;
        RECT 515.400 498.300 516.600 500.400 ;
        RECT 517.800 501.300 519.600 506.400 ;
        RECT 520.800 502.200 522.600 507.000 ;
        RECT 523.800 501.300 525.600 506.400 ;
        RECT 517.800 499.950 525.600 501.300 ;
        RECT 533.400 501.300 535.200 506.400 ;
        RECT 536.400 502.200 538.200 507.000 ;
        RECT 539.400 501.300 541.200 506.400 ;
        RECT 533.400 499.950 541.200 501.300 ;
        RECT 542.400 500.400 544.200 506.400 ;
        RECT 556.800 503.400 558.600 506.400 ;
        RECT 559.800 503.400 561.600 507.000 ;
        RECT 569.400 503.400 571.200 507.000 ;
        RECT 572.400 503.400 574.200 506.400 ;
        RECT 575.400 503.400 577.200 507.000 ;
        RECT 587.400 506.400 588.600 507.000 ;
        RECT 587.400 503.400 589.200 506.400 ;
        RECT 590.400 503.400 592.200 506.400 ;
        RECT 593.400 503.400 595.200 507.000 ;
        RECT 542.400 498.300 543.600 500.400 ;
        RECT 494.100 493.200 495.900 495.000 ;
        RECT 497.400 493.200 498.600 498.300 ;
        RECT 515.400 497.250 519.150 498.300 ;
        RECT 500.100 493.200 501.900 495.000 ;
        RECT 493.950 491.100 496.050 493.200 ;
        RECT 496.950 491.100 499.050 493.200 ;
        RECT 499.950 491.100 502.050 493.200 ;
        RECT 515.100 493.050 516.900 494.850 ;
        RECT 517.950 493.050 519.150 497.250 ;
        RECT 539.850 497.250 543.600 498.300 ;
        RECT 521.100 493.050 522.900 494.850 ;
        RECT 536.100 493.050 537.900 494.850 ;
        RECT 539.850 493.050 541.050 497.250 ;
        RECT 552.000 495.450 556.050 496.050 ;
        RECT 542.100 493.050 543.900 494.850 ;
        RECT 551.550 493.950 556.050 495.450 ;
        RECT 474.750 485.100 485.850 485.700 ;
        RECT 437.400 482.700 445.200 483.600 ;
        RECT 421.800 471.600 423.600 477.600 ;
        RECT 424.800 471.000 426.600 477.600 ;
        RECT 437.400 471.600 439.200 482.700 ;
        RECT 440.400 471.000 442.200 481.800 ;
        RECT 443.400 471.600 445.200 482.700 ;
        RECT 446.400 471.600 448.200 483.600 ;
        RECT 452.550 471.600 454.350 483.600 ;
        RECT 457.950 483.300 460.050 484.200 ;
        RECT 460.950 483.300 466.050 484.200 ;
        RECT 468.150 484.500 485.850 485.100 ;
        RECT 468.150 484.200 476.550 484.500 ;
        RECT 460.950 482.400 461.850 483.300 ;
        RECT 459.150 480.600 461.850 482.400 ;
        RECT 462.750 482.100 464.550 482.400 ;
        RECT 468.150 482.100 469.050 484.200 ;
        RECT 484.950 483.600 485.850 484.500 ;
        RECT 462.750 481.200 469.050 482.100 ;
        RECT 469.950 482.700 471.750 483.300 ;
        RECT 469.950 481.500 477.450 482.700 ;
        RECT 462.750 480.600 464.550 481.200 ;
        RECT 476.250 480.600 477.450 481.500 ;
        RECT 457.950 477.600 461.850 479.700 ;
        RECT 466.950 479.550 468.750 480.300 ;
        RECT 471.750 479.550 473.550 480.300 ;
        RECT 466.950 478.500 473.550 479.550 ;
        RECT 476.250 478.500 481.050 480.600 ;
        RECT 455.550 471.000 457.350 474.600 ;
        RECT 460.050 471.600 461.850 477.600 ;
        RECT 464.250 471.000 466.050 477.600 ;
        RECT 467.850 471.600 469.650 478.500 ;
        RECT 476.250 477.600 477.450 478.500 ;
        RECT 470.850 471.000 472.650 477.600 ;
        RECT 475.650 471.600 477.450 477.600 ;
        RECT 481.050 471.000 482.850 477.600 ;
        RECT 484.050 471.600 485.850 483.600 ;
        RECT 497.400 477.600 498.600 491.100 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 520.950 490.950 523.050 493.050 ;
        RECT 523.950 490.950 526.050 493.050 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 538.950 490.950 541.050 493.050 ;
        RECT 541.950 490.950 544.050 493.050 ;
        RECT 518.850 477.600 520.050 490.950 ;
        RECT 524.100 489.150 525.900 490.950 ;
        RECT 533.100 489.150 534.900 490.950 ;
        RECT 494.400 471.000 496.200 477.600 ;
        RECT 497.400 471.600 499.200 477.600 ;
        RECT 500.400 471.000 502.200 477.600 ;
        RECT 515.400 471.000 517.200 477.600 ;
        RECT 518.400 471.600 520.200 477.600 ;
        RECT 523.500 471.000 525.300 483.600 ;
        RECT 533.700 471.000 535.500 483.600 ;
        RECT 538.950 477.600 540.150 490.950 ;
        RECT 551.550 490.050 552.450 493.950 ;
        RECT 557.400 493.050 558.600 503.400 ;
        RECT 572.700 493.050 573.600 503.400 ;
        RECT 574.950 501.450 577.050 502.050 ;
        RECT 583.950 501.450 586.050 502.050 ;
        RECT 574.950 500.550 586.050 501.450 ;
        RECT 574.950 499.950 577.050 500.550 ;
        RECT 583.950 499.950 586.050 500.550 ;
        RECT 591.300 499.200 592.200 503.400 ;
        RECT 596.400 500.400 598.200 506.400 ;
        RECT 608.400 501.300 610.200 506.400 ;
        RECT 611.400 502.200 613.200 507.000 ;
        RECT 614.400 501.300 616.200 506.400 ;
        RECT 591.300 498.300 594.600 499.200 ;
        RECT 592.800 497.400 594.600 498.300 ;
        RECT 587.100 493.050 588.900 494.850 ;
        RECT 556.950 490.950 559.050 493.050 ;
        RECT 559.950 490.950 562.050 493.050 ;
        RECT 568.950 490.950 571.050 493.050 ;
        RECT 571.950 490.950 574.050 493.050 ;
        RECT 574.950 490.950 577.050 493.050 ;
        RECT 586.950 490.950 589.050 493.050 ;
        RECT 589.950 490.950 592.050 493.050 ;
        RECT 551.550 488.550 556.050 490.050 ;
        RECT 552.000 487.950 556.050 488.550 ;
        RECT 557.400 477.600 558.600 490.950 ;
        RECT 560.100 489.150 561.900 490.950 ;
        RECT 569.100 489.150 570.900 490.950 ;
        RECT 572.700 483.600 573.600 490.950 ;
        RECT 575.100 489.150 576.900 490.950 ;
        RECT 590.100 489.150 591.900 490.950 ;
        RECT 593.700 486.900 594.600 497.400 ;
        RECT 597.000 493.050 598.050 500.400 ;
        RECT 608.400 499.950 616.200 501.300 ;
        RECT 617.400 500.400 619.200 506.400 ;
        RECT 617.400 498.300 618.600 500.400 ;
        RECT 614.850 497.250 618.600 498.300 ;
        RECT 629.400 498.600 631.200 506.400 ;
        RECT 633.900 500.400 635.700 507.000 ;
        RECT 636.900 502.200 638.700 506.400 ;
        RECT 636.900 500.400 639.600 502.200 ;
        RECT 635.100 498.600 636.900 499.500 ;
        RECT 629.400 497.700 636.900 498.600 ;
        RECT 611.100 493.050 612.900 494.850 ;
        RECT 614.850 493.050 616.050 497.250 ;
        RECT 617.100 493.050 618.900 494.850 ;
        RECT 629.100 493.200 630.900 495.000 ;
        RECT 592.800 486.300 594.600 486.900 ;
        RECT 587.400 485.100 594.600 486.300 ;
        RECT 595.950 490.950 598.050 493.050 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 610.950 490.950 613.050 493.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 616.950 490.950 619.050 493.050 ;
        RECT 628.950 491.100 631.050 493.200 ;
        RECT 587.400 483.600 588.600 485.100 ;
        RECT 595.950 483.600 597.300 490.950 ;
        RECT 608.100 489.150 609.900 490.950 ;
        RECT 538.800 471.600 540.600 477.600 ;
        RECT 541.800 471.000 543.600 477.600 ;
        RECT 556.800 471.600 558.600 477.600 ;
        RECT 559.800 471.000 561.600 477.600 ;
        RECT 569.400 471.000 571.200 483.600 ;
        RECT 572.700 482.400 576.300 483.600 ;
        RECT 574.500 471.600 576.300 482.400 ;
        RECT 583.950 480.450 586.050 480.900 ;
        RECT 578.550 480.000 586.050 480.450 ;
        RECT 577.950 479.550 586.050 480.000 ;
        RECT 577.950 475.950 580.050 479.550 ;
        RECT 583.950 478.800 586.050 479.550 ;
        RECT 587.400 471.600 589.200 483.600 ;
        RECT 591.900 471.000 593.700 483.600 ;
        RECT 594.900 482.100 597.300 483.600 ;
        RECT 594.900 471.600 596.700 482.100 ;
        RECT 608.700 471.000 610.500 483.600 ;
        RECT 613.950 477.600 615.150 490.950 ;
        RECT 632.400 477.600 633.300 497.700 ;
        RECT 638.700 493.200 639.600 500.400 ;
        RECT 653.400 499.200 655.200 506.400 ;
        RECT 658.500 500.400 660.300 507.000 ;
        RECT 668.400 500.400 670.200 506.400 ;
        RECT 675.600 501.000 677.400 506.400 ;
        RECT 668.400 499.500 669.900 500.400 ;
        RECT 653.400 498.300 657.600 499.200 ;
        RECT 653.100 493.200 654.900 495.000 ;
        RECT 656.400 493.200 657.600 498.300 ;
        RECT 668.400 498.000 672.750 499.500 ;
        RECT 670.650 497.400 672.750 498.000 ;
        RECT 676.350 498.900 677.250 501.000 ;
        RECT 683.400 500.400 685.200 506.400 ;
        RECT 697.800 503.400 699.600 507.000 ;
        RECT 700.800 503.400 702.600 506.400 ;
        RECT 703.800 503.400 705.600 507.000 ;
        RECT 716.700 503.400 718.500 507.000 ;
        RECT 680.700 499.500 685.200 500.400 ;
        RECT 673.650 495.900 675.450 497.700 ;
        RECT 676.350 496.800 679.350 498.900 ;
        RECT 680.700 497.100 682.800 499.500 ;
        RECT 673.200 495.000 675.300 495.900 ;
        RECT 659.100 493.200 660.900 495.000 ;
        RECT 668.250 493.800 675.300 495.000 ;
        RECT 668.250 493.200 670.050 493.800 ;
        RECT 634.950 491.100 637.050 493.200 ;
        RECT 637.950 491.100 640.050 493.200 ;
        RECT 652.950 491.100 655.050 493.200 ;
        RECT 655.950 491.100 658.050 493.200 ;
        RECT 658.950 491.100 661.050 493.200 ;
        RECT 667.950 491.100 670.050 493.200 ;
        RECT 635.100 489.300 636.900 491.100 ;
        RECT 638.700 483.600 639.600 491.100 ;
        RECT 613.800 471.600 615.600 477.600 ;
        RECT 616.800 471.000 618.600 477.600 ;
        RECT 629.400 471.000 631.200 477.600 ;
        RECT 632.400 471.600 634.200 477.600 ;
        RECT 635.400 471.000 637.200 477.600 ;
        RECT 638.400 471.600 640.200 483.600 ;
        RECT 656.400 477.600 657.600 491.100 ;
        RECT 673.200 490.800 675.300 492.900 ;
        RECT 673.200 489.000 675.000 490.800 ;
        RECT 676.350 490.200 677.250 496.800 ;
        RECT 694.950 495.450 697.050 496.050 ;
        RECT 678.150 492.900 680.250 495.000 ;
        RECT 689.550 494.550 697.050 495.450 ;
        RECT 678.300 491.100 680.100 492.900 ;
        RECT 682.950 491.100 685.050 493.200 ;
        RECT 676.350 488.700 679.350 490.200 ;
        RECT 683.100 489.450 684.900 491.100 ;
        RECT 689.550 489.450 690.450 494.550 ;
        RECT 694.950 493.950 697.050 494.550 ;
        RECT 701.400 493.050 702.300 503.400 ;
        RECT 719.700 501.600 721.500 506.400 ;
        RECT 716.400 500.400 721.500 501.600 ;
        RECT 724.200 500.400 726.000 507.000 ;
        RECT 734.400 503.400 736.200 507.000 ;
        RECT 737.400 503.400 739.200 506.400 ;
        RECT 740.400 503.400 742.200 507.000 ;
        RECT 716.400 493.200 717.300 500.400 ;
        RECT 721.950 498.450 724.050 499.350 ;
        RECT 730.950 498.450 733.050 499.050 ;
        RECT 721.950 497.550 733.050 498.450 ;
        RECT 721.950 497.250 724.050 497.550 ;
        RECT 730.950 496.950 733.050 497.550 ;
        RECT 719.100 493.200 720.900 495.000 ;
        RECT 725.100 493.200 726.900 495.000 ;
        RECT 697.950 490.950 700.050 493.050 ;
        RECT 700.950 490.950 703.050 493.050 ;
        RECT 703.950 490.950 706.050 493.050 ;
        RECT 715.950 491.100 718.050 493.200 ;
        RECT 718.950 491.100 721.050 493.200 ;
        RECT 721.950 491.100 724.050 493.200 ;
        RECT 724.950 491.100 727.050 493.200 ;
        RECT 737.700 493.050 738.600 503.400 ;
        RECT 752.400 500.400 754.200 506.400 ;
        RECT 759.900 500.400 761.700 506.400 ;
        RECT 767.400 500.400 769.200 506.400 ;
        RECT 779.400 503.400 781.200 507.000 ;
        RECT 782.400 503.400 784.200 506.400 ;
        RECT 785.400 503.400 787.200 507.000 ;
        RECT 747.000 498.450 751.050 499.050 ;
        RECT 746.550 496.950 751.050 498.450 ;
        RECT 753.000 498.600 754.200 500.400 ;
        RECT 760.200 498.900 761.400 500.400 ;
        RECT 764.400 499.500 769.200 500.400 ;
        RECT 753.000 497.700 759.300 498.600 ;
        RECT 683.100 489.300 690.450 489.450 ;
        RECT 677.250 488.100 679.350 488.700 ;
        RECT 683.550 488.550 690.450 489.300 ;
        RECT 698.100 489.150 699.900 490.950 ;
        RECT 658.950 486.450 661.050 486.900 ;
        RECT 667.950 486.450 670.050 487.050 ;
        RECT 658.950 485.550 670.050 486.450 ;
        RECT 674.550 485.700 676.350 487.800 ;
        RECT 658.950 484.800 661.050 485.550 ;
        RECT 667.950 484.950 670.050 485.550 ;
        RECT 671.100 484.800 676.350 485.700 ;
        RECT 671.100 483.900 673.200 484.800 ;
        RECT 668.400 482.700 673.200 483.900 ;
        RECT 678.000 483.600 679.200 488.100 ;
        RECT 675.900 482.700 679.200 483.600 ;
        RECT 680.100 483.600 682.200 484.500 ;
        RECT 701.400 483.600 702.300 490.950 ;
        RECT 704.100 489.150 705.900 490.950 ;
        RECT 716.400 483.600 717.300 491.100 ;
        RECT 722.100 489.300 723.900 491.100 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 739.950 490.950 742.050 493.050 ;
        RECT 734.100 489.150 735.900 490.950 ;
        RECT 737.700 483.600 738.600 490.950 ;
        RECT 740.100 489.150 741.900 490.950 ;
        RECT 746.550 489.450 747.450 496.950 ;
        RECT 757.200 495.600 759.300 497.700 ;
        RECT 752.250 493.200 754.050 495.000 ;
        RECT 757.500 493.800 759.300 495.600 ;
        RECT 760.200 496.800 763.050 498.900 ;
        RECT 764.400 498.300 766.500 499.500 ;
        RECT 751.950 492.300 754.050 493.200 ;
        RECT 751.950 491.100 759.300 492.300 ;
        RECT 757.500 490.500 759.300 491.100 ;
        RECT 760.200 491.100 761.250 496.800 ;
        RECT 762.150 493.800 764.250 495.900 ;
        RECT 762.600 492.000 764.400 493.800 ;
        RECT 766.950 491.100 769.050 493.200 ;
        RECT 782.700 493.050 783.600 503.400 ;
        RECT 797.700 500.400 799.500 507.000 ;
        RECT 802.800 499.200 804.600 506.400 ;
        RECT 816.000 500.400 817.800 507.000 ;
        RECT 820.500 501.600 822.300 506.400 ;
        RECT 823.500 503.400 825.300 507.000 ;
        RECT 838.800 503.400 840.600 506.400 ;
        RECT 841.800 503.400 843.600 507.000 ;
        RECT 820.500 500.400 825.600 501.600 ;
        RECT 800.400 498.300 804.600 499.200 ;
        RECT 797.100 493.200 798.900 495.000 ;
        RECT 800.400 493.200 801.600 498.300 ;
        RECT 810.000 495.450 814.050 496.050 ;
        RECT 803.100 493.200 804.900 495.000 ;
        RECT 809.550 493.950 814.050 495.450 ;
        RECT 760.200 490.200 762.600 491.100 ;
        RECT 743.550 488.550 747.450 489.450 ;
        RECT 743.550 487.050 744.450 488.550 ;
        RECT 756.300 487.500 760.050 489.300 ;
        RECT 760.950 488.100 763.050 490.200 ;
        RECT 767.100 489.450 768.900 491.100 ;
        RECT 778.950 490.950 781.050 493.050 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 796.950 491.100 799.050 493.200 ;
        RECT 799.950 491.100 802.050 493.200 ;
        RECT 802.950 491.100 805.050 493.200 ;
        RECT 772.950 489.450 775.050 490.050 ;
        RECT 767.100 489.300 775.050 489.450 ;
        RECT 767.550 488.550 775.050 489.300 ;
        RECT 779.100 489.150 780.900 490.950 ;
        RECT 757.950 487.200 760.050 487.500 ;
        RECT 739.950 485.550 744.450 487.050 ;
        RECT 761.100 486.000 762.000 488.100 ;
        RECT 772.950 487.950 775.050 488.550 ;
        RECT 739.950 484.950 744.000 485.550 ;
        RECT 754.800 483.600 756.900 485.700 ;
        RECT 760.500 485.100 762.000 486.000 ;
        RECT 760.500 483.600 761.700 485.100 ;
        RECT 652.800 471.000 654.600 477.600 ;
        RECT 655.800 471.600 657.600 477.600 ;
        RECT 658.800 471.000 660.600 477.600 ;
        RECT 668.400 471.600 670.200 482.700 ;
        RECT 675.900 471.600 677.700 482.700 ;
        RECT 680.100 482.400 685.200 483.600 ;
        RECT 683.400 471.600 685.200 482.400 ;
        RECT 698.700 482.400 702.300 483.600 ;
        RECT 698.700 471.600 700.500 482.400 ;
        RECT 703.800 471.000 705.600 483.600 ;
        RECT 715.800 471.600 717.600 483.600 ;
        RECT 718.800 482.700 726.600 483.600 ;
        RECT 718.800 471.600 720.600 482.700 ;
        RECT 721.800 471.000 723.600 481.800 ;
        RECT 724.800 471.600 726.600 482.700 ;
        RECT 734.400 471.000 736.200 483.600 ;
        RECT 737.700 482.400 741.300 483.600 ;
        RECT 739.500 471.600 741.300 482.400 ;
        RECT 752.400 482.700 756.900 483.600 ;
        RECT 752.400 471.600 754.200 482.700 ;
        RECT 759.900 478.050 761.700 483.600 ;
        RECT 764.400 483.600 766.500 484.500 ;
        RECT 782.700 483.600 783.600 490.950 ;
        RECT 785.100 489.150 786.900 490.950 ;
        RECT 764.400 482.400 769.200 483.600 ;
        RECT 759.900 475.950 763.050 478.050 ;
        RECT 759.900 471.600 761.700 475.950 ;
        RECT 767.400 471.600 769.200 482.400 ;
        RECT 779.400 471.000 781.200 483.600 ;
        RECT 782.700 482.400 786.300 483.600 ;
        RECT 784.500 471.600 786.300 482.400 ;
        RECT 800.400 477.600 801.600 491.100 ;
        RECT 809.550 490.050 810.450 493.950 ;
        RECT 815.100 493.200 816.900 495.000 ;
        RECT 821.100 493.200 822.900 495.000 ;
        RECT 824.700 493.200 825.600 500.400 ;
        RECT 826.950 495.450 831.000 496.050 ;
        RECT 826.950 493.950 831.450 495.450 ;
        RECT 814.950 491.100 817.050 493.200 ;
        RECT 817.950 491.100 820.050 493.200 ;
        RECT 820.950 491.100 823.050 493.200 ;
        RECT 823.950 491.100 826.050 493.200 ;
        RECT 805.950 488.550 810.450 490.050 ;
        RECT 818.100 489.300 819.900 491.100 ;
        RECT 805.950 487.950 810.000 488.550 ;
        RECT 824.700 483.600 825.600 491.100 ;
        RECT 830.550 490.050 831.450 493.950 ;
        RECT 839.400 493.050 840.600 503.400 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 826.950 488.550 831.450 490.050 ;
        RECT 826.950 487.950 831.000 488.550 ;
        RECT 815.400 482.700 823.200 483.600 ;
        RECT 797.400 471.000 799.200 477.600 ;
        RECT 800.400 471.600 802.200 477.600 ;
        RECT 803.400 471.000 805.200 477.600 ;
        RECT 815.400 471.600 817.200 482.700 ;
        RECT 818.400 471.000 820.200 481.800 ;
        RECT 821.400 471.600 823.200 482.700 ;
        RECT 824.400 471.600 826.200 483.600 ;
        RECT 839.400 477.600 840.600 490.950 ;
        RECT 842.100 489.150 843.900 490.950 ;
        RECT 838.800 471.600 840.600 477.600 ;
        RECT 841.800 471.000 843.600 477.600 ;
        RECT 11.400 461.400 13.200 468.000 ;
        RECT 14.400 461.400 16.200 467.400 ;
        RECT 14.850 448.050 16.050 461.400 ;
        RECT 19.500 455.400 21.300 468.000 ;
        RECT 31.800 461.400 33.600 467.400 ;
        RECT 34.800 462.000 36.600 468.000 ;
        RECT 32.700 461.100 33.600 461.400 ;
        RECT 37.800 461.400 39.600 467.400 ;
        RECT 40.800 461.400 42.600 468.000 ;
        RECT 52.800 461.400 54.600 467.400 ;
        RECT 55.800 462.000 57.600 468.000 ;
        RECT 37.800 461.100 39.300 461.400 ;
        RECT 32.700 460.200 39.300 461.100 ;
        RECT 53.700 461.100 54.600 461.400 ;
        RECT 58.800 461.400 60.600 467.400 ;
        RECT 61.800 461.400 63.600 468.000 ;
        RECT 73.800 461.400 75.600 467.400 ;
        RECT 76.800 462.000 78.600 468.000 ;
        RECT 58.800 461.100 60.300 461.400 ;
        RECT 53.700 460.200 60.300 461.100 ;
        RECT 74.700 461.100 75.600 461.400 ;
        RECT 79.800 461.400 81.600 467.400 ;
        RECT 82.800 461.400 84.600 468.000 ;
        RECT 79.800 461.100 81.300 461.400 ;
        RECT 74.700 460.200 81.300 461.100 ;
        RECT 20.100 448.050 21.900 449.850 ;
        RECT 10.950 445.950 13.050 448.050 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 16.950 445.950 19.050 448.050 ;
        RECT 19.950 445.950 22.050 448.050 ;
        RECT 32.700 447.900 33.600 460.200 ;
        RECT 38.100 447.900 39.900 449.700 ;
        RECT 53.700 447.900 54.600 460.200 ;
        RECT 59.100 447.900 60.900 449.700 ;
        RECT 74.700 447.900 75.600 460.200 ;
        RECT 92.700 455.400 94.500 468.000 ;
        RECT 97.800 461.400 99.600 467.400 ;
        RECT 100.800 461.400 102.600 468.000 ;
        RECT 116.400 461.400 118.200 468.000 ;
        RECT 119.400 461.400 121.200 467.400 ;
        RECT 79.950 453.450 82.050 454.050 ;
        RECT 85.950 453.450 88.050 454.050 ;
        RECT 79.950 452.550 88.050 453.450 ;
        RECT 79.950 451.950 82.050 452.550 ;
        RECT 85.950 451.950 88.050 452.550 ;
        RECT 80.100 447.900 81.900 449.700 ;
        RECT 92.100 448.050 93.900 449.850 ;
        RECT 97.950 448.050 99.150 461.400 ;
        RECT 119.850 448.050 121.050 461.400 ;
        RECT 124.500 455.400 126.300 468.000 ;
        RECT 136.800 461.400 138.600 468.000 ;
        RECT 139.800 461.400 141.600 467.400 ;
        RECT 142.800 461.400 144.600 468.000 ;
        RECT 136.950 450.450 139.050 451.050 ;
        RECT 125.100 448.050 126.900 449.850 ;
        RECT 131.550 449.550 139.050 450.450 ;
        RECT 11.100 444.150 12.900 445.950 ;
        RECT 13.950 441.750 15.150 445.950 ;
        RECT 17.100 444.150 18.900 445.950 ;
        RECT 31.950 445.800 34.050 447.900 ;
        RECT 34.950 445.800 37.050 447.900 ;
        RECT 37.950 445.800 40.050 447.900 ;
        RECT 40.950 445.800 43.050 447.900 ;
        RECT 52.950 445.800 55.050 447.900 ;
        RECT 55.950 445.800 58.050 447.900 ;
        RECT 58.950 445.800 61.050 447.900 ;
        RECT 61.950 445.800 64.050 447.900 ;
        RECT 73.950 445.800 76.050 447.900 ;
        RECT 76.950 445.800 79.050 447.900 ;
        RECT 79.950 445.800 82.050 447.900 ;
        RECT 82.950 445.800 85.050 447.900 ;
        RECT 91.950 445.950 94.050 448.050 ;
        RECT 94.950 445.950 97.050 448.050 ;
        RECT 97.950 445.950 100.050 448.050 ;
        RECT 100.950 445.950 103.050 448.050 ;
        RECT 115.950 445.950 118.050 448.050 ;
        RECT 118.950 445.950 121.050 448.050 ;
        RECT 121.950 445.950 124.050 448.050 ;
        RECT 124.950 445.950 127.050 448.050 ;
        RECT 11.400 440.700 15.150 441.750 ;
        RECT 32.700 442.200 33.600 445.800 ;
        RECT 35.100 444.000 36.900 445.800 ;
        RECT 41.100 444.000 42.900 445.800 ;
        RECT 53.700 442.200 54.600 445.800 ;
        RECT 56.100 444.000 57.900 445.800 ;
        RECT 62.100 444.000 63.900 445.800 ;
        RECT 74.700 442.200 75.600 445.800 ;
        RECT 77.100 444.000 78.900 445.800 ;
        RECT 83.100 444.000 84.900 445.800 ;
        RECT 95.100 444.150 96.900 445.950 ;
        RECT 32.700 441.000 36.000 442.200 ;
        RECT 11.400 438.600 12.600 440.700 ;
        RECT 10.800 432.600 12.600 438.600 ;
        RECT 13.800 437.700 21.600 439.050 ;
        RECT 13.800 432.600 15.600 437.700 ;
        RECT 16.800 432.000 18.600 436.800 ;
        RECT 19.800 432.600 21.600 437.700 ;
        RECT 34.200 432.600 36.000 441.000 ;
        RECT 40.800 432.000 42.600 441.600 ;
        RECT 53.700 441.000 57.000 442.200 ;
        RECT 55.200 432.600 57.000 441.000 ;
        RECT 61.800 432.000 63.600 441.600 ;
        RECT 74.700 441.000 78.000 442.200 ;
        RECT 98.850 441.750 100.050 445.950 ;
        RECT 101.100 444.150 102.900 445.950 ;
        RECT 116.100 444.150 117.900 445.950 ;
        RECT 118.950 441.750 120.150 445.950 ;
        RECT 122.100 444.150 123.900 445.950 ;
        RECT 131.550 445.050 132.450 449.550 ;
        RECT 136.950 448.950 139.050 449.550 ;
        RECT 140.400 447.900 141.600 461.400 ;
        RECT 152.400 456.300 154.200 467.400 ;
        RECT 159.900 456.300 161.700 467.400 ;
        RECT 167.400 456.600 169.200 467.400 ;
        RECT 181.800 461.400 183.600 468.000 ;
        RECT 184.800 461.400 186.600 467.400 ;
        RECT 187.800 461.400 189.600 468.000 ;
        RECT 197.400 461.400 199.200 468.000 ;
        RECT 200.400 461.400 202.200 467.400 ;
        RECT 203.400 461.400 205.200 468.000 ;
        RECT 152.400 455.100 157.200 456.300 ;
        RECT 159.900 455.400 163.200 456.300 ;
        RECT 155.100 454.200 157.200 455.100 ;
        RECT 155.100 453.300 160.350 454.200 ;
        RECT 158.550 451.200 160.350 453.300 ;
        RECT 162.000 450.900 163.200 455.400 ;
        RECT 164.100 455.400 169.200 456.600 ;
        RECT 164.100 454.500 166.200 455.400 ;
        RECT 161.250 450.300 163.350 450.900 ;
        RECT 168.000 450.450 172.050 451.050 ;
        RECT 157.200 448.200 159.000 450.000 ;
        RECT 160.350 448.800 163.350 450.300 ;
        RECT 167.550 449.700 172.050 450.450 ;
        RECT 167.100 448.950 172.050 449.700 ;
        RECT 136.950 445.800 139.050 447.900 ;
        RECT 139.950 445.800 142.050 447.900 ;
        RECT 142.950 445.800 145.050 447.900 ;
        RECT 151.950 445.800 154.050 447.900 ;
        RECT 157.200 446.100 159.300 448.200 ;
        RECT 127.950 443.550 132.450 445.050 ;
        RECT 137.100 444.000 138.900 445.800 ;
        RECT 127.950 442.950 132.000 443.550 ;
        RECT 76.200 432.600 78.000 441.000 ;
        RECT 82.800 432.000 84.600 441.600 ;
        RECT 98.850 440.700 102.600 441.750 ;
        RECT 92.400 437.700 100.200 439.050 ;
        RECT 92.400 432.600 94.200 437.700 ;
        RECT 95.400 432.000 97.200 436.800 ;
        RECT 98.400 432.600 100.200 437.700 ;
        RECT 101.400 438.600 102.600 440.700 ;
        RECT 116.400 440.700 120.150 441.750 ;
        RECT 140.400 440.700 141.600 445.800 ;
        RECT 143.100 444.000 144.900 445.800 ;
        RECT 152.250 445.200 154.050 445.800 ;
        RECT 152.250 444.000 159.300 445.200 ;
        RECT 157.200 443.100 159.300 444.000 ;
        RECT 154.650 441.000 156.750 441.600 ;
        RECT 157.650 441.300 159.450 443.100 ;
        RECT 160.350 442.200 161.250 448.800 ;
        RECT 167.100 447.900 168.900 448.950 ;
        RECT 185.400 447.900 186.600 461.400 ;
        RECT 162.300 446.100 164.100 447.900 ;
        RECT 162.150 444.000 164.250 446.100 ;
        RECT 166.950 445.800 169.050 447.900 ;
        RECT 181.950 445.800 184.050 447.900 ;
        RECT 184.950 445.800 187.050 447.900 ;
        RECT 187.950 445.800 190.050 447.900 ;
        RECT 196.950 445.800 199.050 447.900 ;
        RECT 182.100 444.000 183.900 445.800 ;
        RECT 116.400 438.600 117.600 440.700 ;
        RECT 137.400 439.800 141.600 440.700 ;
        RECT 101.400 432.600 103.200 438.600 ;
        RECT 115.800 432.600 117.600 438.600 ;
        RECT 118.800 437.700 126.600 439.050 ;
        RECT 118.800 432.600 120.600 437.700 ;
        RECT 121.800 432.000 123.600 436.800 ;
        RECT 124.800 432.600 126.600 437.700 ;
        RECT 137.400 432.600 139.200 439.800 ;
        RECT 152.400 439.500 156.750 441.000 ;
        RECT 160.350 440.100 163.350 442.200 ;
        RECT 152.400 438.600 153.900 439.500 ;
        RECT 142.500 432.000 144.300 438.600 ;
        RECT 152.400 432.600 154.200 438.600 ;
        RECT 160.350 438.000 161.250 440.100 ;
        RECT 164.700 439.500 166.800 441.900 ;
        RECT 185.400 440.700 186.600 445.800 ;
        RECT 188.100 444.000 189.900 445.800 ;
        RECT 197.100 444.000 198.900 445.800 ;
        RECT 200.400 441.300 201.300 461.400 ;
        RECT 206.400 455.400 208.200 467.400 ;
        RECT 220.800 461.400 222.600 468.000 ;
        RECT 223.800 461.400 225.600 467.400 ;
        RECT 226.800 461.400 228.600 468.000 ;
        RECT 203.100 447.900 204.900 449.700 ;
        RECT 206.700 447.900 207.600 455.400 ;
        RECT 224.400 447.900 225.600 461.400 ;
        RECT 238.800 455.400 240.600 467.400 ;
        RECT 241.800 461.400 243.600 468.000 ;
        RECT 244.800 461.400 246.600 467.400 ;
        RECT 247.800 461.400 249.600 468.000 ;
        RECT 226.950 450.450 229.050 451.050 ;
        RECT 235.950 450.450 238.050 451.050 ;
        RECT 226.950 449.550 238.050 450.450 ;
        RECT 226.950 448.950 229.050 449.550 ;
        RECT 235.950 448.950 238.050 449.550 ;
        RECT 239.400 447.900 240.300 455.400 ;
        RECT 242.100 447.900 243.900 449.700 ;
        RECT 202.950 445.800 205.050 447.900 ;
        RECT 205.950 445.800 208.050 447.900 ;
        RECT 220.950 445.800 223.050 447.900 ;
        RECT 223.950 445.800 226.050 447.900 ;
        RECT 226.950 445.800 229.050 447.900 ;
        RECT 238.950 445.800 241.050 447.900 ;
        RECT 241.950 445.800 244.050 447.900 ;
        RECT 182.400 439.800 186.600 440.700 ;
        RECT 197.400 440.400 204.900 441.300 ;
        RECT 164.700 438.600 169.200 439.500 ;
        RECT 159.600 432.600 161.400 438.000 ;
        RECT 167.400 432.600 169.200 438.600 ;
        RECT 182.400 432.600 184.200 439.800 ;
        RECT 187.500 432.000 189.300 438.600 ;
        RECT 197.400 432.600 199.200 440.400 ;
        RECT 203.100 439.500 204.900 440.400 ;
        RECT 206.700 438.600 207.600 445.800 ;
        RECT 221.100 444.000 222.900 445.800 ;
        RECT 224.400 440.700 225.600 445.800 ;
        RECT 227.100 444.000 228.900 445.800 ;
        RECT 201.900 432.000 203.700 438.600 ;
        RECT 204.900 436.800 207.600 438.600 ;
        RECT 221.400 439.800 225.600 440.700 ;
        RECT 204.900 432.600 206.700 436.800 ;
        RECT 221.400 432.600 223.200 439.800 ;
        RECT 239.400 438.600 240.300 445.800 ;
        RECT 245.700 441.300 246.600 461.400 ;
        RECT 257.400 456.300 259.200 467.400 ;
        RECT 257.400 455.400 261.900 456.300 ;
        RECT 264.900 455.400 266.700 467.400 ;
        RECT 272.400 456.600 274.200 467.400 ;
        RECT 286.800 461.400 288.600 468.000 ;
        RECT 289.800 461.400 291.600 467.400 ;
        RECT 292.800 461.400 294.600 468.000 ;
        RECT 259.800 453.300 261.900 455.400 ;
        RECT 265.500 453.900 266.700 455.400 ;
        RECT 269.400 455.400 274.200 456.600 ;
        RECT 269.400 454.500 271.500 455.400 ;
        RECT 265.500 453.000 267.000 453.900 ;
        RECT 262.950 451.500 265.050 451.800 ;
        RECT 250.950 450.450 253.050 451.050 ;
        RECT 256.950 450.450 259.050 451.050 ;
        RECT 250.950 449.550 259.050 450.450 ;
        RECT 261.300 449.700 265.050 451.500 ;
        RECT 266.100 450.900 267.000 453.000 ;
        RECT 280.950 453.450 283.050 454.050 ;
        RECT 286.950 453.450 289.050 454.050 ;
        RECT 280.950 452.550 289.050 453.450 ;
        RECT 280.950 451.950 283.050 452.550 ;
        RECT 286.950 451.950 289.050 452.550 ;
        RECT 250.950 448.950 253.050 449.550 ;
        RECT 256.950 448.950 259.050 449.550 ;
        RECT 265.950 448.800 268.050 450.900 ;
        RECT 274.950 450.450 277.050 451.050 ;
        RECT 286.950 450.450 289.050 450.900 ;
        RECT 262.500 447.900 264.300 448.500 ;
        RECT 247.950 445.800 250.050 447.900 ;
        RECT 256.950 446.700 264.300 447.900 ;
        RECT 265.200 447.900 267.600 448.800 ;
        RECT 272.100 447.900 273.900 449.700 ;
        RECT 274.950 449.550 289.050 450.450 ;
        RECT 274.950 448.950 277.050 449.550 ;
        RECT 286.950 448.800 289.050 449.550 ;
        RECT 290.400 447.900 291.600 461.400 ;
        RECT 304.800 455.400 306.600 467.400 ;
        RECT 307.800 461.400 309.600 468.000 ;
        RECT 310.800 461.400 312.600 467.400 ;
        RECT 304.800 448.050 306.000 455.400 ;
        RECT 311.400 454.500 312.600 461.400 ;
        RECT 320.700 455.400 322.500 468.000 ;
        RECT 325.800 461.400 327.600 467.400 ;
        RECT 328.800 461.400 330.600 468.000 ;
        RECT 341.400 461.400 343.200 468.000 ;
        RECT 344.400 461.400 346.200 467.400 ;
        RECT 347.400 461.400 349.200 468.000 ;
        RECT 306.900 453.600 312.600 454.500 ;
        RECT 306.900 452.700 308.850 453.600 ;
        RECT 256.950 445.800 259.050 446.700 ;
        RECT 248.100 444.000 249.900 445.800 ;
        RECT 257.250 444.000 259.050 445.800 ;
        RECT 262.500 443.400 264.300 445.200 ;
        RECT 262.200 441.300 264.300 443.400 ;
        RECT 242.100 440.400 249.600 441.300 ;
        RECT 242.100 439.500 243.900 440.400 ;
        RECT 226.500 432.000 228.300 438.600 ;
        RECT 239.400 436.800 242.100 438.600 ;
        RECT 240.300 432.600 242.100 436.800 ;
        RECT 243.300 432.000 245.100 438.600 ;
        RECT 247.800 432.600 249.600 440.400 ;
        RECT 258.000 440.400 264.300 441.300 ;
        RECT 265.200 442.200 266.250 447.900 ;
        RECT 267.600 445.200 269.400 447.000 ;
        RECT 271.950 445.800 274.050 447.900 ;
        RECT 286.950 445.800 289.050 447.900 ;
        RECT 289.950 445.800 292.050 447.900 ;
        RECT 292.950 445.800 295.050 447.900 ;
        RECT 304.800 445.950 307.050 448.050 ;
        RECT 267.150 443.100 269.250 445.200 ;
        RECT 287.100 444.000 288.900 445.800 ;
        RECT 258.000 438.600 259.200 440.400 ;
        RECT 265.200 440.100 268.050 442.200 ;
        RECT 290.400 440.700 291.600 445.800 ;
        RECT 293.100 444.000 294.900 445.800 ;
        RECT 265.200 438.600 266.400 440.100 ;
        RECT 269.400 439.500 271.500 440.700 ;
        RECT 287.400 439.800 291.600 440.700 ;
        RECT 269.400 438.600 274.200 439.500 ;
        RECT 257.400 432.600 259.200 438.600 ;
        RECT 264.900 432.600 266.700 438.600 ;
        RECT 272.400 432.600 274.200 438.600 ;
        RECT 287.400 432.600 289.200 439.800 ;
        RECT 304.800 438.600 306.000 445.950 ;
        RECT 307.950 441.300 308.850 452.700 ;
        RECT 311.100 448.050 312.900 449.850 ;
        RECT 320.100 448.050 321.900 449.850 ;
        RECT 325.950 448.050 327.150 461.400 ;
        RECT 328.950 453.450 331.050 454.050 ;
        RECT 334.950 453.450 337.050 454.050 ;
        RECT 328.950 452.550 337.050 453.450 ;
        RECT 328.950 451.950 331.050 452.550 ;
        RECT 334.950 451.950 337.050 452.550 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 322.950 445.950 325.050 448.050 ;
        RECT 325.950 445.950 328.050 448.050 ;
        RECT 328.950 445.950 331.050 448.050 ;
        RECT 344.400 447.900 345.600 461.400 ;
        RECT 354.150 455.400 355.950 467.400 ;
        RECT 357.150 461.400 358.950 468.000 ;
        RECT 362.550 461.400 364.350 467.400 ;
        RECT 367.350 461.400 369.150 468.000 ;
        RECT 362.550 460.500 363.750 461.400 ;
        RECT 370.350 460.500 372.150 467.400 ;
        RECT 373.950 461.400 375.750 468.000 ;
        RECT 378.150 461.400 379.950 467.400 ;
        RECT 382.650 464.400 384.450 468.000 ;
        RECT 358.950 458.400 363.750 460.500 ;
        RECT 366.450 459.450 373.050 460.500 ;
        RECT 366.450 458.700 368.250 459.450 ;
        RECT 371.250 458.700 373.050 459.450 ;
        RECT 378.150 459.300 382.050 461.400 ;
        RECT 362.550 457.500 363.750 458.400 ;
        RECT 375.450 457.800 377.250 458.400 ;
        RECT 362.550 456.300 370.050 457.500 ;
        RECT 368.250 455.700 370.050 456.300 ;
        RECT 370.950 456.900 377.250 457.800 ;
        RECT 354.150 454.500 355.050 455.400 ;
        RECT 370.950 454.800 371.850 456.900 ;
        RECT 375.450 456.600 377.250 456.900 ;
        RECT 378.150 456.600 380.850 458.400 ;
        RECT 378.150 455.700 379.050 456.600 ;
        RECT 363.450 454.500 371.850 454.800 ;
        RECT 354.150 453.900 371.850 454.500 ;
        RECT 373.950 454.800 379.050 455.700 ;
        RECT 379.950 454.800 382.050 455.700 ;
        RECT 385.650 455.400 387.450 467.400 ;
        RECT 354.150 453.300 365.250 453.900 ;
        RECT 323.100 444.150 324.900 445.950 ;
        RECT 306.900 440.400 308.850 441.300 ;
        RECT 326.850 441.750 328.050 445.950 ;
        RECT 329.100 444.150 330.900 445.950 ;
        RECT 340.950 445.800 343.050 447.900 ;
        RECT 343.950 445.800 346.050 447.900 ;
        RECT 346.950 445.800 349.050 447.900 ;
        RECT 341.100 444.000 342.900 445.800 ;
        RECT 326.850 440.700 330.600 441.750 ;
        RECT 306.900 439.500 312.600 440.400 ;
        RECT 292.500 432.000 294.300 438.600 ;
        RECT 304.800 432.600 306.600 438.600 ;
        RECT 311.400 435.600 312.600 439.500 ;
        RECT 307.800 432.000 309.600 435.600 ;
        RECT 310.800 432.600 312.600 435.600 ;
        RECT 320.400 437.700 328.200 439.050 ;
        RECT 320.400 432.600 322.200 437.700 ;
        RECT 323.400 432.000 325.200 436.800 ;
        RECT 326.400 432.600 328.200 437.700 ;
        RECT 329.400 438.600 330.600 440.700 ;
        RECT 344.400 440.700 345.600 445.800 ;
        RECT 347.100 444.000 348.900 445.800 ;
        RECT 344.400 439.800 348.600 440.700 ;
        RECT 329.400 432.600 331.200 438.600 ;
        RECT 341.700 432.000 343.500 438.600 ;
        RECT 346.800 432.600 348.600 439.800 ;
        RECT 354.150 438.600 355.050 453.300 ;
        RECT 363.450 453.000 365.250 453.300 ;
        RECT 355.950 445.950 358.050 448.050 ;
        RECT 364.950 446.400 367.050 448.050 ;
        RECT 356.100 444.150 357.900 445.950 ;
        RECT 359.100 445.200 367.050 446.400 ;
        RECT 359.100 444.600 360.900 445.200 ;
        RECT 357.000 443.400 357.900 444.150 ;
        RECT 362.100 443.400 363.900 444.000 ;
        RECT 357.000 442.200 363.900 443.400 ;
        RECT 373.950 442.200 374.850 454.800 ;
        RECT 379.950 453.600 384.150 454.800 ;
        RECT 383.250 451.800 385.050 453.600 ;
        RECT 386.250 448.050 387.450 455.400 ;
        RECT 395.400 461.400 397.200 467.400 ;
        RECT 398.400 461.400 400.200 468.000 ;
        RECT 395.400 454.500 396.600 461.400 ;
        RECT 401.400 455.400 403.200 467.400 ;
        RECT 413.400 461.400 415.200 468.000 ;
        RECT 416.400 461.400 418.200 467.400 ;
        RECT 419.400 461.400 421.200 468.000 ;
        RECT 431.400 461.400 433.200 468.000 ;
        RECT 434.400 461.400 436.200 467.400 ;
        RECT 437.400 461.400 439.200 468.000 ;
        RECT 452.400 461.400 454.200 468.000 ;
        RECT 455.400 461.400 457.200 467.400 ;
        RECT 395.400 453.600 401.100 454.500 ;
        RECT 399.150 452.700 401.100 453.600 ;
        RECT 395.100 448.050 396.900 449.850 ;
        RECT 382.950 447.750 387.450 448.050 ;
        RECT 381.150 445.950 387.450 447.750 ;
        RECT 394.950 445.950 397.050 448.050 ;
        RECT 362.850 441.000 374.850 442.200 ;
        RECT 362.850 439.200 363.900 441.000 ;
        RECT 373.050 440.400 374.850 441.000 ;
        RECT 354.150 432.600 355.950 438.600 ;
        RECT 358.950 436.500 361.050 438.600 ;
        RECT 362.550 437.400 364.350 439.200 ;
        RECT 386.250 438.600 387.450 445.950 ;
        RECT 399.150 441.300 400.050 452.700 ;
        RECT 402.000 448.050 403.200 455.400 ;
        RECT 400.950 445.950 403.200 448.050 ;
        RECT 416.400 447.900 417.600 461.400 ;
        RECT 434.400 447.900 435.600 461.400 ;
        RECT 442.950 453.450 445.050 454.050 ;
        RECT 451.950 453.450 454.050 454.050 ;
        RECT 442.950 452.550 454.050 453.450 ;
        RECT 442.950 451.950 445.050 452.550 ;
        RECT 451.950 451.950 454.050 452.550 ;
        RECT 455.850 448.050 457.050 461.400 ;
        RECT 460.500 455.400 462.300 468.000 ;
        RECT 465.150 455.400 466.950 467.400 ;
        RECT 468.150 461.400 469.950 468.000 ;
        RECT 473.550 461.400 475.350 467.400 ;
        RECT 478.350 461.400 480.150 468.000 ;
        RECT 473.550 460.500 474.750 461.400 ;
        RECT 481.350 460.500 483.150 467.400 ;
        RECT 484.950 461.400 486.750 468.000 ;
        RECT 489.150 461.400 490.950 467.400 ;
        RECT 493.650 464.400 495.450 468.000 ;
        RECT 469.950 458.400 474.750 460.500 ;
        RECT 477.450 459.450 484.050 460.500 ;
        RECT 477.450 458.700 479.250 459.450 ;
        RECT 482.250 458.700 484.050 459.450 ;
        RECT 489.150 459.300 493.050 461.400 ;
        RECT 473.550 457.500 474.750 458.400 ;
        RECT 486.450 457.800 488.250 458.400 ;
        RECT 473.550 456.300 481.050 457.500 ;
        RECT 479.250 455.700 481.050 456.300 ;
        RECT 481.950 456.900 488.250 457.800 ;
        RECT 465.150 454.500 466.050 455.400 ;
        RECT 481.950 454.800 482.850 456.900 ;
        RECT 486.450 456.600 488.250 456.900 ;
        RECT 489.150 456.600 491.850 458.400 ;
        RECT 489.150 455.700 490.050 456.600 ;
        RECT 474.450 454.500 482.850 454.800 ;
        RECT 465.150 453.900 482.850 454.500 ;
        RECT 484.950 454.800 490.050 455.700 ;
        RECT 490.950 454.800 493.050 455.700 ;
        RECT 496.650 455.400 498.450 467.400 ;
        RECT 509.400 461.400 511.200 468.000 ;
        RECT 512.400 461.400 514.200 467.400 ;
        RECT 465.150 453.300 476.250 453.900 ;
        RECT 461.100 448.050 462.900 449.850 ;
        RECT 399.150 440.400 401.100 441.300 ;
        RECT 365.850 437.550 367.650 438.300 ;
        RECT 379.950 437.700 382.050 438.600 ;
        RECT 365.850 436.500 370.800 437.550 ;
        RECT 360.000 435.600 361.050 436.500 ;
        RECT 369.750 435.600 370.800 436.500 ;
        RECT 378.300 436.500 382.050 437.700 ;
        RECT 378.300 435.600 379.350 436.500 ;
        RECT 357.150 432.000 358.950 435.600 ;
        RECT 360.000 434.700 363.750 435.600 ;
        RECT 361.950 432.600 363.750 434.700 ;
        RECT 366.450 432.000 368.250 435.600 ;
        RECT 369.750 432.600 371.550 435.600 ;
        RECT 373.350 432.000 375.150 435.600 ;
        RECT 377.550 432.600 379.350 435.600 ;
        RECT 382.350 432.000 384.150 435.600 ;
        RECT 385.650 432.600 387.450 438.600 ;
        RECT 395.400 439.500 401.100 440.400 ;
        RECT 395.400 435.600 396.600 439.500 ;
        RECT 402.000 438.600 403.200 445.950 ;
        RECT 412.950 445.800 415.050 447.900 ;
        RECT 415.950 445.800 418.050 447.900 ;
        RECT 418.950 445.800 421.050 447.900 ;
        RECT 430.950 445.800 433.050 447.900 ;
        RECT 433.950 445.800 436.050 447.900 ;
        RECT 436.950 445.800 439.050 447.900 ;
        RECT 451.950 445.950 454.050 448.050 ;
        RECT 454.950 445.950 457.050 448.050 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 413.100 444.000 414.900 445.800 ;
        RECT 416.400 440.700 417.600 445.800 ;
        RECT 419.100 444.000 420.900 445.800 ;
        RECT 431.100 444.000 432.900 445.800 ;
        RECT 434.400 440.700 435.600 445.800 ;
        RECT 437.100 444.000 438.900 445.800 ;
        RECT 452.100 444.150 453.900 445.950 ;
        RECT 454.950 441.750 456.150 445.950 ;
        RECT 458.100 444.150 459.900 445.950 ;
        RECT 452.400 440.700 456.150 441.750 ;
        RECT 416.400 439.800 420.600 440.700 ;
        RECT 434.400 439.800 438.600 440.700 ;
        RECT 395.400 432.600 397.200 435.600 ;
        RECT 398.400 432.000 400.200 435.600 ;
        RECT 401.400 432.600 403.200 438.600 ;
        RECT 413.700 432.000 415.500 438.600 ;
        RECT 418.800 432.600 420.600 439.800 ;
        RECT 431.700 432.000 433.500 438.600 ;
        RECT 436.800 432.600 438.600 439.800 ;
        RECT 452.400 438.600 453.600 440.700 ;
        RECT 451.800 432.600 453.600 438.600 ;
        RECT 454.800 437.700 462.600 439.050 ;
        RECT 454.800 432.600 456.600 437.700 ;
        RECT 457.800 432.000 459.600 436.800 ;
        RECT 460.800 432.600 462.600 437.700 ;
        RECT 465.150 438.600 466.050 453.300 ;
        RECT 474.450 453.000 476.250 453.300 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 475.950 446.400 478.050 448.050 ;
        RECT 467.100 444.150 468.900 445.950 ;
        RECT 470.100 445.200 478.050 446.400 ;
        RECT 470.100 444.600 471.900 445.200 ;
        RECT 468.000 443.400 468.900 444.150 ;
        RECT 473.100 443.400 474.900 444.000 ;
        RECT 468.000 442.200 474.900 443.400 ;
        RECT 484.950 442.200 485.850 454.800 ;
        RECT 490.950 453.600 495.150 454.800 ;
        RECT 494.250 451.800 496.050 453.600 ;
        RECT 497.250 448.050 498.450 455.400 ;
        RECT 499.950 450.450 502.050 451.050 ;
        RECT 505.950 450.450 508.050 450.900 ;
        RECT 499.950 449.550 508.050 450.450 ;
        RECT 499.950 448.950 502.050 449.550 ;
        RECT 505.950 448.800 508.050 449.550 ;
        RECT 512.850 448.050 514.050 461.400 ;
        RECT 517.500 455.400 519.300 468.000 ;
        RECT 529.800 455.400 531.600 467.400 ;
        RECT 532.800 455.400 534.600 468.000 ;
        RECT 545.400 461.400 547.200 468.000 ;
        RECT 548.400 461.400 550.200 467.400 ;
        RECT 518.100 448.050 519.900 449.850 ;
        RECT 493.950 447.750 498.450 448.050 ;
        RECT 492.150 445.950 498.450 447.750 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 511.950 445.950 514.050 448.050 ;
        RECT 514.950 445.950 517.050 448.050 ;
        RECT 517.950 445.950 520.050 448.050 ;
        RECT 530.400 447.900 531.600 455.400 ;
        RECT 548.850 448.050 550.050 461.400 ;
        RECT 553.500 455.400 555.300 468.000 ;
        RECT 563.400 455.400 565.200 467.400 ;
        RECT 567.900 455.400 569.700 468.000 ;
        RECT 570.900 456.900 572.700 467.400 ;
        RECT 586.800 461.400 588.600 467.400 ;
        RECT 589.800 461.400 591.600 468.000 ;
        RECT 570.900 455.400 573.300 456.900 ;
        RECT 563.400 453.900 564.600 455.400 ;
        RECT 563.400 452.700 570.600 453.900 ;
        RECT 568.800 452.100 570.600 452.700 ;
        RECT 554.100 448.050 555.900 449.850 ;
        RECT 566.100 448.050 567.900 449.850 ;
        RECT 473.850 441.000 485.850 442.200 ;
        RECT 473.850 439.200 474.900 441.000 ;
        RECT 484.050 440.400 485.850 441.000 ;
        RECT 465.150 432.600 466.950 438.600 ;
        RECT 469.950 436.500 472.050 438.600 ;
        RECT 473.550 437.400 475.350 439.200 ;
        RECT 497.250 438.600 498.450 445.950 ;
        RECT 509.100 444.150 510.900 445.950 ;
        RECT 511.950 441.750 513.150 445.950 ;
        RECT 515.100 444.150 516.900 445.950 ;
        RECT 529.950 445.800 532.050 447.900 ;
        RECT 532.950 445.800 535.050 447.900 ;
        RECT 544.950 445.950 547.050 448.050 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 553.950 445.950 556.050 448.050 ;
        RECT 562.950 445.950 565.050 448.050 ;
        RECT 565.950 445.950 568.050 448.050 ;
        RECT 509.400 440.700 513.150 441.750 ;
        RECT 509.400 438.600 510.600 440.700 ;
        RECT 476.850 437.550 478.650 438.300 ;
        RECT 490.950 437.700 493.050 438.600 ;
        RECT 476.850 436.500 481.800 437.550 ;
        RECT 471.000 435.600 472.050 436.500 ;
        RECT 480.750 435.600 481.800 436.500 ;
        RECT 489.300 436.500 493.050 437.700 ;
        RECT 489.300 435.600 490.350 436.500 ;
        RECT 468.150 432.000 469.950 435.600 ;
        RECT 471.000 434.700 474.750 435.600 ;
        RECT 472.950 432.600 474.750 434.700 ;
        RECT 477.450 432.000 479.250 435.600 ;
        RECT 480.750 432.600 482.550 435.600 ;
        RECT 484.350 432.000 486.150 435.600 ;
        RECT 488.550 432.600 490.350 435.600 ;
        RECT 493.350 432.000 495.150 435.600 ;
        RECT 496.650 432.600 498.450 438.600 ;
        RECT 508.800 432.600 510.600 438.600 ;
        RECT 511.800 437.700 519.600 439.050 ;
        RECT 530.400 438.600 531.600 445.800 ;
        RECT 533.100 444.000 534.900 445.800 ;
        RECT 545.100 444.150 546.900 445.950 ;
        RECT 547.950 441.750 549.150 445.950 ;
        RECT 551.100 444.150 552.900 445.950 ;
        RECT 563.100 444.150 564.900 445.950 ;
        RECT 545.400 440.700 549.150 441.750 ;
        RECT 569.700 441.600 570.600 452.100 ;
        RECT 571.950 448.050 573.300 455.400 ;
        RECT 587.400 448.050 588.600 461.400 ;
        RECT 601.800 455.400 603.600 467.400 ;
        RECT 604.800 456.300 606.600 467.400 ;
        RECT 607.800 457.200 609.600 468.000 ;
        RECT 610.800 456.300 612.600 467.400 ;
        RECT 604.800 455.400 612.600 456.300 ;
        RECT 622.800 455.400 624.600 467.400 ;
        RECT 625.800 456.300 627.600 467.400 ;
        RECT 628.800 457.200 630.600 468.000 ;
        RECT 631.800 456.300 633.600 467.400 ;
        RECT 643.800 461.400 645.600 467.400 ;
        RECT 646.800 461.400 648.600 468.000 ;
        RECT 625.800 455.400 633.600 456.300 ;
        RECT 590.100 448.050 591.900 449.850 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 586.950 445.950 589.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 602.400 447.900 603.300 455.400 ;
        RECT 610.950 450.450 613.050 451.050 ;
        RECT 616.950 450.450 619.050 451.050 ;
        RECT 608.100 447.900 609.900 449.700 ;
        RECT 610.950 449.550 619.050 450.450 ;
        RECT 610.950 448.950 613.050 449.550 ;
        RECT 616.950 448.950 619.050 449.550 ;
        RECT 623.400 447.900 624.300 455.400 ;
        RECT 625.950 453.450 628.050 454.050 ;
        RECT 637.950 453.450 640.050 454.050 ;
        RECT 625.950 452.550 640.050 453.450 ;
        RECT 625.950 451.950 628.050 452.550 ;
        RECT 637.950 451.950 640.050 452.550 ;
        RECT 629.100 447.900 630.900 449.700 ;
        RECT 644.400 448.050 645.600 461.400 ;
        RECT 656.700 455.400 658.500 468.000 ;
        RECT 661.800 461.400 663.600 467.400 ;
        RECT 664.800 461.400 666.600 468.000 ;
        RECT 680.400 461.400 682.200 468.000 ;
        RECT 683.400 461.400 685.200 467.400 ;
        RECT 647.100 448.050 648.900 449.850 ;
        RECT 656.100 448.050 657.900 449.850 ;
        RECT 661.950 448.050 663.150 461.400 ;
        RECT 683.850 448.050 685.050 461.400 ;
        RECT 688.500 455.400 690.300 468.000 ;
        RECT 700.800 461.400 702.600 467.400 ;
        RECT 703.800 462.000 705.600 468.000 ;
        RECT 701.700 461.100 702.600 461.400 ;
        RECT 706.800 461.400 708.600 467.400 ;
        RECT 709.800 461.400 711.600 468.000 ;
        RECT 721.800 461.400 723.600 468.000 ;
        RECT 724.800 461.400 726.600 467.400 ;
        RECT 727.800 461.400 729.600 468.000 ;
        RECT 739.800 461.400 741.600 468.000 ;
        RECT 742.800 461.400 744.600 467.400 ;
        RECT 745.800 461.400 747.600 468.000 ;
        RECT 755.400 461.400 757.200 468.000 ;
        RECT 758.400 461.400 760.200 467.400 ;
        RECT 773.400 461.400 775.200 468.000 ;
        RECT 776.400 461.400 778.200 467.400 ;
        RECT 706.800 461.100 708.300 461.400 ;
        RECT 701.700 460.200 708.300 461.100 ;
        RECT 689.100 448.050 690.900 449.850 ;
        RECT 568.800 440.700 570.600 441.600 ;
        RECT 545.400 438.600 546.600 440.700 ;
        RECT 567.300 439.800 570.600 440.700 ;
        RECT 511.800 432.600 513.600 437.700 ;
        RECT 514.800 432.000 516.600 436.800 ;
        RECT 517.800 432.600 519.600 437.700 ;
        RECT 529.800 432.600 531.600 438.600 ;
        RECT 532.800 432.000 534.600 438.600 ;
        RECT 544.800 432.600 546.600 438.600 ;
        RECT 547.800 437.700 555.600 439.050 ;
        RECT 547.800 432.600 549.600 437.700 ;
        RECT 550.800 432.000 552.600 436.800 ;
        RECT 553.800 432.600 555.600 437.700 ;
        RECT 567.300 435.600 568.200 439.800 ;
        RECT 573.000 438.600 574.050 445.950 ;
        RECT 563.400 432.600 565.200 435.600 ;
        RECT 566.400 432.600 568.200 435.600 ;
        RECT 563.400 432.000 564.600 432.600 ;
        RECT 569.400 432.000 571.200 435.600 ;
        RECT 572.400 432.600 574.200 438.600 ;
        RECT 587.400 435.600 588.600 445.950 ;
        RECT 601.950 445.800 604.050 447.900 ;
        RECT 604.950 445.800 607.050 447.900 ;
        RECT 607.950 445.800 610.050 447.900 ;
        RECT 610.950 445.800 613.050 447.900 ;
        RECT 622.950 445.800 625.050 447.900 ;
        RECT 625.950 445.800 628.050 447.900 ;
        RECT 628.950 445.800 631.050 447.900 ;
        RECT 631.950 445.800 634.050 447.900 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 646.950 445.950 649.050 448.050 ;
        RECT 655.950 445.950 658.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 679.950 445.950 682.050 448.050 ;
        RECT 682.950 445.950 685.050 448.050 ;
        RECT 685.950 445.950 688.050 448.050 ;
        RECT 688.950 445.950 691.050 448.050 ;
        RECT 701.700 447.900 702.600 460.200 ;
        RECT 709.950 453.450 712.050 454.050 ;
        RECT 721.950 453.450 724.050 454.050 ;
        RECT 709.950 452.550 724.050 453.450 ;
        RECT 709.950 451.950 712.050 452.550 ;
        RECT 721.950 451.950 724.050 452.550 ;
        RECT 709.950 450.450 712.050 450.900 ;
        RECT 718.950 450.450 721.050 451.050 ;
        RECT 707.100 447.900 708.900 449.700 ;
        RECT 709.950 449.550 721.050 450.450 ;
        RECT 709.950 448.800 712.050 449.550 ;
        RECT 718.950 448.950 721.050 449.550 ;
        RECT 725.400 447.900 726.600 461.400 ;
        RECT 727.950 453.450 730.050 454.050 ;
        RECT 739.950 453.450 742.050 454.050 ;
        RECT 727.950 452.550 742.050 453.450 ;
        RECT 727.950 451.950 730.050 452.550 ;
        RECT 739.950 451.950 742.050 452.550 ;
        RECT 739.950 450.450 742.050 450.900 ;
        RECT 734.550 449.550 742.050 450.450 ;
        RECT 602.400 438.600 603.300 445.800 ;
        RECT 605.100 444.000 606.900 445.800 ;
        RECT 611.100 444.000 612.900 445.800 ;
        RECT 623.400 438.600 624.300 445.800 ;
        RECT 626.100 444.000 627.900 445.800 ;
        RECT 632.100 444.000 633.900 445.800 ;
        RECT 602.400 437.400 607.500 438.600 ;
        RECT 586.800 432.600 588.600 435.600 ;
        RECT 589.800 432.000 591.600 435.600 ;
        RECT 602.700 432.000 604.500 435.600 ;
        RECT 605.700 432.600 607.500 437.400 ;
        RECT 610.200 432.000 612.000 438.600 ;
        RECT 623.400 437.400 628.500 438.600 ;
        RECT 623.700 432.000 625.500 435.600 ;
        RECT 626.700 432.600 628.500 437.400 ;
        RECT 631.200 432.000 633.000 438.600 ;
        RECT 644.400 435.600 645.600 445.950 ;
        RECT 659.100 444.150 660.900 445.950 ;
        RECT 662.850 441.750 664.050 445.950 ;
        RECT 665.100 444.150 666.900 445.950 ;
        RECT 680.100 444.150 681.900 445.950 ;
        RECT 682.950 441.750 684.150 445.950 ;
        RECT 686.100 444.150 687.900 445.950 ;
        RECT 700.950 445.800 703.050 447.900 ;
        RECT 703.950 445.800 706.050 447.900 ;
        RECT 706.950 445.800 709.050 447.900 ;
        RECT 709.950 445.800 712.050 447.900 ;
        RECT 721.950 445.800 724.050 447.900 ;
        RECT 724.950 445.800 727.050 447.900 ;
        RECT 727.950 445.800 730.050 447.900 ;
        RECT 662.850 440.700 666.600 441.750 ;
        RECT 656.400 437.700 664.200 439.050 ;
        RECT 643.800 432.600 645.600 435.600 ;
        RECT 646.800 432.000 648.600 435.600 ;
        RECT 656.400 432.600 658.200 437.700 ;
        RECT 659.400 432.000 661.200 436.800 ;
        RECT 662.400 432.600 664.200 437.700 ;
        RECT 665.400 438.600 666.600 440.700 ;
        RECT 680.400 440.700 684.150 441.750 ;
        RECT 701.700 442.200 702.600 445.800 ;
        RECT 704.100 444.000 705.900 445.800 ;
        RECT 710.100 444.000 711.900 445.800 ;
        RECT 722.100 444.000 723.900 445.800 ;
        RECT 701.700 441.000 705.000 442.200 ;
        RECT 680.400 438.600 681.600 440.700 ;
        RECT 665.400 432.600 667.200 438.600 ;
        RECT 679.800 432.600 681.600 438.600 ;
        RECT 682.800 437.700 690.600 439.050 ;
        RECT 682.800 432.600 684.600 437.700 ;
        RECT 685.800 432.000 687.600 436.800 ;
        RECT 688.800 432.600 690.600 437.700 ;
        RECT 703.200 432.600 705.000 441.000 ;
        RECT 709.800 432.000 711.600 441.600 ;
        RECT 725.400 440.700 726.600 445.800 ;
        RECT 728.100 444.000 729.900 445.800 ;
        RECT 734.550 445.050 735.450 449.550 ;
        RECT 739.950 448.800 742.050 449.550 ;
        RECT 743.400 447.900 744.600 461.400 ;
        RECT 755.100 448.050 756.900 449.850 ;
        RECT 758.400 448.050 759.600 461.400 ;
        RECT 760.950 453.450 763.050 454.050 ;
        RECT 772.950 453.450 775.050 454.050 ;
        RECT 760.950 452.550 775.050 453.450 ;
        RECT 760.950 451.950 763.050 452.550 ;
        RECT 772.950 451.950 775.050 452.550 ;
        RECT 776.850 448.050 778.050 461.400 ;
        RECT 781.500 455.400 783.300 468.000 ;
        RECT 791.400 456.300 793.200 467.400 ;
        RECT 794.400 457.200 796.200 468.000 ;
        RECT 797.400 456.300 799.200 467.400 ;
        RECT 791.400 455.400 799.200 456.300 ;
        RECT 800.400 455.400 802.200 467.400 ;
        RECT 812.400 461.400 814.200 467.400 ;
        RECT 815.400 461.400 817.200 468.000 ;
        RECT 782.100 448.050 783.900 449.850 ;
        RECT 739.950 445.800 742.050 447.900 ;
        RECT 742.950 445.800 745.050 447.900 ;
        RECT 745.950 445.800 748.050 447.900 ;
        RECT 754.950 445.950 757.050 448.050 ;
        RECT 757.950 445.950 760.050 448.050 ;
        RECT 772.950 445.950 775.050 448.050 ;
        RECT 775.950 445.950 778.050 448.050 ;
        RECT 778.950 445.950 781.050 448.050 ;
        RECT 781.950 445.950 784.050 448.050 ;
        RECT 794.100 447.900 795.900 449.700 ;
        RECT 800.700 447.900 801.600 455.400 ;
        RECT 812.400 454.500 813.600 461.400 ;
        RECT 818.400 455.400 820.200 467.400 ;
        RECT 832.800 456.600 834.600 467.400 ;
        RECT 832.800 455.400 837.600 456.600 ;
        RECT 812.400 453.600 818.100 454.500 ;
        RECT 816.150 452.700 818.100 453.600 ;
        RECT 812.100 448.050 813.900 449.850 ;
        RECT 734.550 443.550 739.050 445.050 ;
        RECT 740.100 444.000 741.900 445.800 ;
        RECT 735.000 442.950 739.050 443.550 ;
        RECT 743.400 440.700 744.600 445.800 ;
        RECT 746.100 444.000 747.900 445.800 ;
        RECT 722.400 439.800 726.600 440.700 ;
        RECT 740.400 439.800 744.600 440.700 ;
        RECT 722.400 432.600 724.200 439.800 ;
        RECT 727.500 432.000 729.300 438.600 ;
        RECT 740.400 432.600 742.200 439.800 ;
        RECT 745.500 432.000 747.300 438.600 ;
        RECT 758.400 435.600 759.600 445.950 ;
        RECT 773.100 444.150 774.900 445.950 ;
        RECT 775.950 441.750 777.150 445.950 ;
        RECT 779.100 444.150 780.900 445.950 ;
        RECT 790.950 445.800 793.050 447.900 ;
        RECT 793.950 445.800 796.050 447.900 ;
        RECT 796.950 445.800 799.050 447.900 ;
        RECT 799.950 445.800 802.050 447.900 ;
        RECT 811.950 445.950 814.050 448.050 ;
        RECT 791.100 444.000 792.900 445.800 ;
        RECT 797.100 444.000 798.900 445.800 ;
        RECT 773.400 440.700 777.150 441.750 ;
        RECT 773.400 438.600 774.600 440.700 ;
        RECT 755.400 432.000 757.200 435.600 ;
        RECT 758.400 432.600 760.200 435.600 ;
        RECT 772.800 432.600 774.600 438.600 ;
        RECT 775.800 437.700 783.600 439.050 ;
        RECT 800.700 438.600 801.600 445.800 ;
        RECT 816.150 441.300 817.050 452.700 ;
        RECT 819.000 448.050 820.200 455.400 ;
        RECT 835.500 454.500 837.600 455.400 ;
        RECT 840.300 455.400 842.100 467.400 ;
        RECT 847.800 456.300 849.600 467.400 ;
        RECT 845.100 455.400 849.600 456.300 ;
        RECT 840.300 453.900 841.500 455.400 ;
        RECT 840.000 453.000 841.500 453.900 ;
        RECT 845.100 453.300 847.200 455.400 ;
        RECT 829.950 450.450 834.000 451.050 ;
        RECT 840.000 450.900 840.900 453.000 ;
        RECT 841.950 451.500 844.050 451.800 ;
        RECT 829.950 449.700 834.450 450.450 ;
        RECT 829.950 448.950 834.900 449.700 ;
        RECT 817.950 445.950 820.200 448.050 ;
        RECT 833.100 447.900 834.900 448.950 ;
        RECT 838.950 448.800 841.050 450.900 ;
        RECT 841.950 449.700 845.700 451.500 ;
        RECT 847.950 450.450 850.050 451.050 ;
        RECT 853.950 450.450 856.050 451.050 ;
        RECT 847.950 449.550 856.050 450.450 ;
        RECT 847.950 448.950 850.050 449.550 ;
        RECT 853.950 448.950 856.050 449.550 ;
        RECT 839.400 447.900 841.800 448.800 ;
        RECT 816.150 440.400 818.100 441.300 ;
        RECT 775.800 432.600 777.600 437.700 ;
        RECT 778.800 432.000 780.600 436.800 ;
        RECT 781.800 432.600 783.600 437.700 ;
        RECT 792.000 432.000 793.800 438.600 ;
        RECT 796.500 437.400 801.600 438.600 ;
        RECT 812.400 439.500 818.100 440.400 ;
        RECT 796.500 432.600 798.300 437.400 ;
        RECT 812.400 435.600 813.600 439.500 ;
        RECT 819.000 438.600 820.200 445.950 ;
        RECT 832.950 445.800 835.050 447.900 ;
        RECT 837.600 445.200 839.400 447.000 ;
        RECT 837.750 443.100 839.850 445.200 ;
        RECT 840.750 442.200 841.800 447.900 ;
        RECT 842.700 447.900 844.500 448.500 ;
        RECT 842.700 446.700 850.050 447.900 ;
        RECT 847.950 445.800 850.050 446.700 ;
        RECT 835.500 439.500 837.600 440.700 ;
        RECT 838.950 440.100 841.800 442.200 ;
        RECT 842.700 443.400 844.500 445.200 ;
        RECT 847.950 444.000 849.750 445.800 ;
        RECT 842.700 441.300 844.800 443.400 ;
        RECT 842.700 440.400 849.000 441.300 ;
        RECT 799.500 432.000 801.300 435.600 ;
        RECT 812.400 432.600 814.200 435.600 ;
        RECT 815.400 432.000 817.200 435.600 ;
        RECT 818.400 432.600 820.200 438.600 ;
        RECT 832.800 438.600 837.600 439.500 ;
        RECT 840.600 438.600 841.800 440.100 ;
        RECT 847.800 438.600 849.000 440.400 ;
        RECT 832.800 432.600 834.600 438.600 ;
        RECT 840.300 432.600 842.100 438.600 ;
        RECT 847.800 432.600 849.600 438.600 ;
        RECT 11.700 425.400 13.500 429.000 ;
        RECT 14.700 423.600 16.500 428.400 ;
        RECT 11.400 422.400 16.500 423.600 ;
        RECT 19.200 422.400 21.000 429.000 ;
        RECT 31.800 425.400 33.600 428.400 ;
        RECT 34.800 425.400 36.600 429.000 ;
        RECT 11.400 415.200 12.300 422.400 ;
        RECT 13.950 420.450 16.050 420.900 ;
        RECT 28.950 420.450 31.050 421.050 ;
        RECT 13.950 419.550 31.050 420.450 ;
        RECT 13.950 418.800 16.050 419.550 ;
        RECT 28.950 418.950 31.050 419.550 ;
        RECT 14.100 415.200 15.900 417.000 ;
        RECT 20.100 415.200 21.900 417.000 ;
        RECT 10.950 413.100 13.050 415.200 ;
        RECT 13.950 413.100 16.050 415.200 ;
        RECT 16.950 413.100 19.050 415.200 ;
        RECT 19.950 413.100 22.050 415.200 ;
        RECT 32.400 415.050 33.600 425.400 ;
        RECT 49.200 420.000 51.000 428.400 ;
        RECT 47.700 418.800 51.000 420.000 ;
        RECT 55.800 419.400 57.600 429.000 ;
        RECT 67.800 422.400 69.600 428.400 ;
        RECT 68.400 420.300 69.600 422.400 ;
        RECT 70.800 423.300 72.600 428.400 ;
        RECT 73.800 424.200 75.600 429.000 ;
        RECT 76.800 423.300 78.600 428.400 ;
        RECT 89.700 425.400 91.500 429.000 ;
        RECT 92.700 423.600 94.500 428.400 ;
        RECT 70.800 421.950 78.600 423.300 ;
        RECT 89.400 422.400 94.500 423.600 ;
        RECT 97.200 422.400 99.000 429.000 ;
        RECT 68.400 419.250 72.150 420.300 ;
        RECT 42.000 417.450 46.050 418.050 ;
        RECT 41.550 415.950 46.050 417.450 ;
        RECT 11.400 405.600 12.300 413.100 ;
        RECT 17.100 411.300 18.900 413.100 ;
        RECT 31.950 412.950 34.050 415.050 ;
        RECT 34.950 412.950 37.050 415.050 ;
        RECT 16.950 408.450 19.050 409.050 ;
        RECT 28.950 408.450 31.050 409.050 ;
        RECT 16.950 407.550 31.050 408.450 ;
        RECT 16.950 406.950 19.050 407.550 ;
        RECT 28.950 406.950 31.050 407.550 ;
        RECT 10.800 393.600 12.600 405.600 ;
        RECT 13.800 404.700 21.600 405.600 ;
        RECT 13.800 393.600 15.600 404.700 ;
        RECT 16.800 393.000 18.600 403.800 ;
        RECT 19.800 393.600 21.600 404.700 ;
        RECT 32.400 399.600 33.600 412.950 ;
        RECT 35.100 411.150 36.900 412.950 ;
        RECT 41.550 412.050 42.450 415.950 ;
        RECT 47.700 415.200 48.600 418.800 ;
        RECT 50.100 415.200 51.900 417.000 ;
        RECT 56.100 415.200 57.900 417.000 ;
        RECT 46.950 413.100 49.050 415.200 ;
        RECT 49.950 413.100 52.050 415.200 ;
        RECT 52.950 413.100 55.050 415.200 ;
        RECT 55.950 413.100 58.050 415.200 ;
        RECT 68.100 415.050 69.900 416.850 ;
        RECT 70.950 415.050 72.150 419.250 ;
        RECT 79.950 417.450 84.000 418.050 ;
        RECT 74.100 415.050 75.900 416.850 ;
        RECT 79.950 415.950 84.450 417.450 ;
        RECT 41.550 410.550 46.050 412.050 ;
        RECT 42.000 409.950 46.050 410.550 ;
        RECT 47.700 400.800 48.600 413.100 ;
        RECT 53.100 411.300 54.900 413.100 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 70.950 412.950 73.050 415.050 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 76.950 412.950 79.050 415.050 ;
        RECT 47.700 399.900 54.300 400.800 ;
        RECT 47.700 399.600 48.600 399.900 ;
        RECT 31.800 393.600 33.600 399.600 ;
        RECT 34.800 393.000 36.600 399.600 ;
        RECT 46.800 393.600 48.600 399.600 ;
        RECT 52.800 399.600 54.300 399.900 ;
        RECT 71.850 399.600 73.050 412.950 ;
        RECT 77.100 411.150 78.900 412.950 ;
        RECT 83.550 412.050 84.450 415.950 ;
        RECT 89.400 415.200 90.300 422.400 ;
        RECT 112.200 420.000 114.000 428.400 ;
        RECT 110.700 418.800 114.000 420.000 ;
        RECT 118.800 419.400 120.600 429.000 ;
        RECT 128.400 425.400 130.200 429.000 ;
        RECT 131.400 425.400 133.200 428.400 ;
        RECT 92.100 415.200 93.900 417.000 ;
        RECT 98.100 415.200 99.900 417.000 ;
        RECT 110.700 415.200 111.600 418.800 ;
        RECT 113.100 415.200 114.900 417.000 ;
        RECT 119.100 415.200 120.900 417.000 ;
        RECT 88.950 413.100 91.050 415.200 ;
        RECT 91.950 413.100 94.050 415.200 ;
        RECT 94.950 413.100 97.050 415.200 ;
        RECT 97.950 413.100 100.050 415.200 ;
        RECT 109.950 413.100 112.050 415.200 ;
        RECT 112.950 413.100 115.050 415.200 ;
        RECT 115.950 413.100 118.050 415.200 ;
        RECT 118.950 413.100 121.050 415.200 ;
        RECT 131.400 415.050 132.600 425.400 ;
        RECT 143.400 423.300 145.200 428.400 ;
        RECT 146.400 424.200 148.200 429.000 ;
        RECT 149.400 423.300 151.200 428.400 ;
        RECT 143.400 421.950 151.200 423.300 ;
        RECT 152.400 422.400 154.200 428.400 ;
        RECT 164.400 425.400 166.200 429.000 ;
        RECT 167.400 425.400 169.200 428.400 ;
        RECT 170.400 425.400 172.200 429.000 ;
        RECT 152.400 420.300 153.600 422.400 ;
        RECT 149.850 419.250 153.600 420.300 ;
        RECT 146.100 415.050 147.900 416.850 ;
        RECT 149.850 415.050 151.050 419.250 ;
        RECT 152.100 415.050 153.900 416.850 ;
        RECT 167.700 415.050 168.600 425.400 ;
        RECT 185.400 421.200 187.200 428.400 ;
        RECT 190.500 422.400 192.300 429.000 ;
        RECT 200.700 422.400 202.500 429.000 ;
        RECT 205.200 422.400 207.000 428.400 ;
        RECT 209.700 422.400 211.500 429.000 ;
        RECT 224.700 422.400 226.500 429.000 ;
        RECT 185.400 420.300 189.600 421.200 ;
        RECT 185.100 415.200 186.900 417.000 ;
        RECT 188.400 415.200 189.600 420.300 ;
        RECT 191.100 415.200 192.900 417.000 ;
        RECT 200.100 415.200 201.900 417.000 ;
        RECT 205.950 415.200 207.000 422.400 ;
        RECT 229.800 421.200 231.600 428.400 ;
        RECT 227.400 420.300 231.600 421.200 ;
        RECT 245.400 421.200 247.200 428.400 ;
        RECT 250.500 422.400 252.300 429.000 ;
        RECT 262.800 422.400 264.600 428.400 ;
        RECT 245.400 420.300 249.600 421.200 ;
        RECT 212.100 415.200 213.900 417.000 ;
        RECT 224.100 415.200 225.900 417.000 ;
        RECT 227.400 415.200 228.600 420.300 ;
        RECT 230.100 415.200 231.900 417.000 ;
        RECT 245.100 415.200 246.900 417.000 ;
        RECT 248.400 415.200 249.600 420.300 ;
        RECT 263.400 420.300 264.600 422.400 ;
        RECT 265.800 423.300 267.600 428.400 ;
        RECT 268.800 424.200 270.600 429.000 ;
        RECT 271.800 423.300 273.600 428.400 ;
        RECT 281.400 425.400 283.200 429.000 ;
        RECT 284.400 425.400 286.200 428.400 ;
        RECT 265.800 421.950 273.600 423.300 ;
        RECT 263.400 419.250 267.150 420.300 ;
        RECT 253.950 417.450 258.000 418.050 ;
        RECT 251.100 415.200 252.900 417.000 ;
        RECT 253.950 415.950 258.450 417.450 ;
        RECT 79.950 410.550 84.450 412.050 ;
        RECT 79.950 409.950 84.000 410.550 ;
        RECT 89.400 405.600 90.300 413.100 ;
        RECT 95.100 411.300 96.900 413.100 ;
        RECT 49.800 393.000 51.600 399.000 ;
        RECT 52.800 393.600 54.600 399.600 ;
        RECT 55.800 393.000 57.600 399.600 ;
        RECT 68.400 393.000 70.200 399.600 ;
        RECT 71.400 393.600 73.200 399.600 ;
        RECT 76.500 393.000 78.300 405.600 ;
        RECT 88.800 393.600 90.600 405.600 ;
        RECT 91.800 404.700 99.600 405.600 ;
        RECT 91.800 393.600 93.600 404.700 ;
        RECT 94.800 393.000 96.600 403.800 ;
        RECT 97.800 393.600 99.600 404.700 ;
        RECT 110.700 400.800 111.600 413.100 ;
        RECT 116.100 411.300 117.900 413.100 ;
        RECT 127.950 412.950 130.050 415.050 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 142.950 412.950 145.050 415.050 ;
        RECT 145.950 412.950 148.050 415.050 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 163.950 412.950 166.050 415.050 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 184.950 413.100 187.050 415.200 ;
        RECT 187.950 413.100 190.050 415.200 ;
        RECT 190.950 413.100 193.050 415.200 ;
        RECT 199.950 413.100 202.050 415.200 ;
        RECT 202.950 413.100 205.050 415.200 ;
        RECT 205.950 413.100 208.050 415.200 ;
        RECT 208.950 413.100 211.050 415.200 ;
        RECT 211.950 413.100 214.050 415.200 ;
        RECT 223.950 413.100 226.050 415.200 ;
        RECT 226.950 413.100 229.050 415.200 ;
        RECT 229.950 413.100 232.050 415.200 ;
        RECT 244.950 413.100 247.050 415.200 ;
        RECT 247.950 413.100 250.050 415.200 ;
        RECT 250.950 413.100 253.050 415.200 ;
        RECT 118.950 411.450 121.050 412.050 ;
        RECT 124.950 411.450 127.050 412.050 ;
        RECT 118.950 410.550 127.050 411.450 ;
        RECT 128.100 411.150 129.900 412.950 ;
        RECT 118.950 409.950 121.050 410.550 ;
        RECT 124.950 409.950 127.050 410.550 ;
        RECT 110.700 399.900 117.300 400.800 ;
        RECT 110.700 399.600 111.600 399.900 ;
        RECT 109.800 393.600 111.600 399.600 ;
        RECT 115.800 399.600 117.300 399.900 ;
        RECT 131.400 399.600 132.600 412.950 ;
        RECT 143.100 411.150 144.900 412.950 ;
        RECT 112.800 393.000 114.600 399.000 ;
        RECT 115.800 393.600 117.600 399.600 ;
        RECT 118.800 393.000 120.600 399.600 ;
        RECT 128.400 393.000 130.200 399.600 ;
        RECT 131.400 393.600 133.200 399.600 ;
        RECT 143.700 393.000 145.500 405.600 ;
        RECT 148.950 399.600 150.150 412.950 ;
        RECT 164.100 411.150 165.900 412.950 ;
        RECT 167.700 405.600 168.600 412.950 ;
        RECT 170.100 411.150 171.900 412.950 ;
        RECT 148.800 393.600 150.600 399.600 ;
        RECT 151.800 393.000 153.600 399.600 ;
        RECT 164.400 393.000 166.200 405.600 ;
        RECT 167.700 404.400 171.300 405.600 ;
        RECT 169.500 393.600 171.300 404.400 ;
        RECT 188.400 399.600 189.600 413.100 ;
        RECT 203.100 411.300 204.900 413.100 ;
        RECT 206.100 407.400 207.000 413.100 ;
        RECT 209.100 411.300 210.900 413.100 ;
        RECT 206.100 406.500 211.200 407.400 ;
        RECT 200.400 404.400 208.200 405.300 ;
        RECT 184.800 393.000 186.600 399.600 ;
        RECT 187.800 393.600 189.600 399.600 ;
        RECT 190.800 393.000 192.600 399.600 ;
        RECT 200.400 393.600 202.200 404.400 ;
        RECT 203.400 393.000 205.200 403.500 ;
        RECT 206.400 394.500 208.200 404.400 ;
        RECT 209.400 395.400 211.200 406.500 ;
        RECT 212.400 394.500 214.200 405.600 ;
        RECT 227.400 399.600 228.600 413.100 ;
        RECT 248.400 399.600 249.600 413.100 ;
        RECT 257.550 412.050 258.450 415.950 ;
        RECT 263.100 415.050 264.900 416.850 ;
        RECT 265.950 415.050 267.150 419.250 ;
        RECT 269.100 415.050 270.900 416.850 ;
        RECT 284.400 415.050 285.600 425.400 ;
        RECT 296.400 419.400 298.200 429.000 ;
        RECT 303.000 420.000 304.800 428.400 ;
        RECT 317.400 425.400 319.200 429.000 ;
        RECT 320.400 425.400 322.200 428.400 ;
        RECT 303.000 418.800 306.300 420.000 ;
        RECT 291.000 417.450 295.050 418.050 ;
        RECT 290.550 415.950 295.050 417.450 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 257.550 410.550 262.050 412.050 ;
        RECT 258.000 409.950 262.050 410.550 ;
        RECT 266.850 399.600 268.050 412.950 ;
        RECT 272.100 411.150 273.900 412.950 ;
        RECT 281.100 411.150 282.900 412.950 ;
        RECT 206.400 393.600 214.200 394.500 ;
        RECT 224.400 393.000 226.200 399.600 ;
        RECT 227.400 393.600 229.200 399.600 ;
        RECT 230.400 393.000 232.200 399.600 ;
        RECT 244.800 393.000 246.600 399.600 ;
        RECT 247.800 393.600 249.600 399.600 ;
        RECT 250.800 393.000 252.600 399.600 ;
        RECT 263.400 393.000 265.200 399.600 ;
        RECT 266.400 393.600 268.200 399.600 ;
        RECT 271.500 393.000 273.300 405.600 ;
        RECT 284.400 399.600 285.600 412.950 ;
        RECT 290.550 412.050 291.450 415.950 ;
        RECT 296.100 415.200 297.900 417.000 ;
        RECT 302.100 415.200 303.900 417.000 ;
        RECT 305.400 415.200 306.300 418.800 ;
        RECT 295.950 413.100 298.050 415.200 ;
        RECT 298.950 413.100 301.050 415.200 ;
        RECT 301.950 413.100 304.050 415.200 ;
        RECT 304.950 413.100 307.050 415.200 ;
        RECT 320.400 415.050 321.600 425.400 ;
        RECT 334.800 422.400 336.600 428.400 ;
        RECT 335.400 420.300 336.600 422.400 ;
        RECT 337.800 423.300 339.600 428.400 ;
        RECT 340.800 424.200 342.600 429.000 ;
        RECT 343.800 423.300 345.600 428.400 ;
        RECT 337.800 421.950 345.600 423.300 ;
        RECT 348.150 422.400 349.950 428.400 ;
        RECT 351.150 425.400 352.950 429.000 ;
        RECT 355.950 426.300 357.750 428.400 ;
        RECT 354.000 425.400 357.750 426.300 ;
        RECT 360.450 425.400 362.250 429.000 ;
        RECT 363.750 425.400 365.550 428.400 ;
        RECT 367.350 425.400 369.150 429.000 ;
        RECT 371.550 425.400 373.350 428.400 ;
        RECT 376.350 425.400 378.150 429.000 ;
        RECT 354.000 424.500 355.050 425.400 ;
        RECT 363.750 424.500 364.800 425.400 ;
        RECT 352.950 422.400 355.050 424.500 ;
        RECT 335.400 419.250 339.150 420.300 ;
        RECT 335.100 415.050 336.900 416.850 ;
        RECT 337.950 415.050 339.150 419.250 ;
        RECT 341.100 415.050 342.900 416.850 ;
        RECT 290.550 410.550 295.050 412.050 ;
        RECT 299.100 411.300 300.900 413.100 ;
        RECT 291.000 409.950 295.050 410.550 ;
        RECT 305.400 400.800 306.300 413.100 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 334.950 412.950 337.050 415.050 ;
        RECT 337.950 412.950 340.050 415.050 ;
        RECT 340.950 412.950 343.050 415.050 ;
        RECT 343.950 412.950 346.050 415.050 ;
        RECT 317.100 411.150 318.900 412.950 ;
        RECT 299.700 399.900 306.300 400.800 ;
        RECT 299.700 399.600 301.200 399.900 ;
        RECT 281.400 393.000 283.200 399.600 ;
        RECT 284.400 393.600 286.200 399.600 ;
        RECT 296.400 393.000 298.200 399.600 ;
        RECT 299.400 393.600 301.200 399.600 ;
        RECT 305.400 399.600 306.300 399.900 ;
        RECT 320.400 399.600 321.600 412.950 ;
        RECT 338.850 399.600 340.050 412.950 ;
        RECT 344.100 411.150 345.900 412.950 ;
        RECT 348.150 407.700 349.050 422.400 ;
        RECT 356.550 421.800 358.350 423.600 ;
        RECT 359.850 423.450 364.800 424.500 ;
        RECT 372.300 424.500 373.350 425.400 ;
        RECT 359.850 422.700 361.650 423.450 ;
        RECT 372.300 423.300 376.050 424.500 ;
        RECT 373.950 422.400 376.050 423.300 ;
        RECT 379.650 422.400 381.450 428.400 ;
        RECT 389.400 425.400 391.200 429.000 ;
        RECT 392.400 425.400 394.200 428.400 ;
        RECT 356.850 420.000 357.900 421.800 ;
        RECT 367.050 420.000 368.850 420.600 ;
        RECT 356.850 418.800 368.850 420.000 ;
        RECT 351.000 417.600 357.900 418.800 ;
        RECT 351.000 416.850 351.900 417.600 ;
        RECT 356.100 417.000 357.900 417.600 ;
        RECT 350.100 415.050 351.900 416.850 ;
        RECT 353.100 415.800 354.900 416.400 ;
        RECT 349.950 412.950 352.050 415.050 ;
        RECT 353.100 414.600 361.050 415.800 ;
        RECT 358.950 412.950 361.050 414.600 ;
        RECT 357.450 407.700 359.250 408.000 ;
        RECT 348.150 407.100 359.250 407.700 ;
        RECT 348.150 406.500 365.850 407.100 ;
        RECT 348.150 405.600 349.050 406.500 ;
        RECT 357.450 406.200 365.850 406.500 ;
        RECT 302.400 393.000 304.200 399.000 ;
        RECT 305.400 393.600 307.200 399.600 ;
        RECT 317.400 393.000 319.200 399.600 ;
        RECT 320.400 393.600 322.200 399.600 ;
        RECT 335.400 393.000 337.200 399.600 ;
        RECT 338.400 393.600 340.200 399.600 ;
        RECT 343.500 393.000 345.300 405.600 ;
        RECT 348.150 393.600 349.950 405.600 ;
        RECT 362.250 404.700 364.050 405.300 ;
        RECT 356.550 403.500 364.050 404.700 ;
        RECT 364.950 404.100 365.850 406.200 ;
        RECT 367.950 406.200 368.850 418.800 ;
        RECT 380.250 415.050 381.450 422.400 ;
        RECT 392.400 415.050 393.600 425.400 ;
        RECT 404.400 423.300 406.200 428.400 ;
        RECT 407.400 424.200 409.200 429.000 ;
        RECT 410.400 423.300 412.200 428.400 ;
        RECT 404.400 421.950 412.200 423.300 ;
        RECT 413.400 422.400 415.200 428.400 ;
        RECT 420.150 422.400 421.950 428.400 ;
        RECT 423.150 425.400 424.950 429.000 ;
        RECT 427.950 426.300 429.750 428.400 ;
        RECT 426.000 425.400 429.750 426.300 ;
        RECT 432.450 425.400 434.250 429.000 ;
        RECT 435.750 425.400 437.550 428.400 ;
        RECT 439.350 425.400 441.150 429.000 ;
        RECT 443.550 425.400 445.350 428.400 ;
        RECT 448.350 425.400 450.150 429.000 ;
        RECT 426.000 424.500 427.050 425.400 ;
        RECT 435.750 424.500 436.800 425.400 ;
        RECT 424.950 422.400 427.050 424.500 ;
        RECT 413.400 420.300 414.600 422.400 ;
        RECT 410.850 419.250 414.600 420.300 ;
        RECT 407.100 415.050 408.900 416.850 ;
        RECT 410.850 415.050 412.050 419.250 ;
        RECT 413.100 415.050 414.900 416.850 ;
        RECT 375.150 413.250 381.450 415.050 ;
        RECT 376.950 412.950 381.450 413.250 ;
        RECT 388.950 412.950 391.050 415.050 ;
        RECT 391.950 412.950 394.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 412.950 412.950 415.050 415.050 ;
        RECT 377.250 407.400 379.050 409.200 ;
        RECT 373.950 406.200 378.150 407.400 ;
        RECT 367.950 405.300 373.050 406.200 ;
        RECT 373.950 405.300 376.050 406.200 ;
        RECT 380.250 405.600 381.450 412.950 ;
        RECT 389.100 411.150 390.900 412.950 ;
        RECT 372.150 404.400 373.050 405.300 ;
        RECT 369.450 404.100 371.250 404.400 ;
        RECT 356.550 402.600 357.750 403.500 ;
        RECT 364.950 403.200 371.250 404.100 ;
        RECT 369.450 402.600 371.250 403.200 ;
        RECT 372.150 402.600 374.850 404.400 ;
        RECT 352.950 400.500 357.750 402.600 ;
        RECT 360.450 401.550 362.250 402.300 ;
        RECT 365.250 401.550 367.050 402.300 ;
        RECT 360.450 400.500 367.050 401.550 ;
        RECT 356.550 399.600 357.750 400.500 ;
        RECT 351.150 393.000 352.950 399.600 ;
        RECT 356.550 393.600 358.350 399.600 ;
        RECT 361.350 393.000 363.150 399.600 ;
        RECT 364.350 393.600 366.150 400.500 ;
        RECT 372.150 399.600 376.050 401.700 ;
        RECT 367.950 393.000 369.750 399.600 ;
        RECT 372.150 393.600 373.950 399.600 ;
        RECT 376.650 393.000 378.450 396.600 ;
        RECT 379.650 393.600 381.450 405.600 ;
        RECT 392.400 399.600 393.600 412.950 ;
        RECT 404.100 411.150 405.900 412.950 ;
        RECT 389.400 393.000 391.200 399.600 ;
        RECT 392.400 393.600 394.200 399.600 ;
        RECT 404.700 393.000 406.500 405.600 ;
        RECT 409.950 399.600 411.150 412.950 ;
        RECT 420.150 407.700 421.050 422.400 ;
        RECT 428.550 421.800 430.350 423.600 ;
        RECT 431.850 423.450 436.800 424.500 ;
        RECT 444.300 424.500 445.350 425.400 ;
        RECT 431.850 422.700 433.650 423.450 ;
        RECT 444.300 423.300 448.050 424.500 ;
        RECT 445.950 422.400 448.050 423.300 ;
        RECT 451.650 422.400 453.450 428.400 ;
        RECT 428.850 420.000 429.900 421.800 ;
        RECT 439.050 420.000 440.850 420.600 ;
        RECT 428.850 418.800 440.850 420.000 ;
        RECT 423.000 417.600 429.900 418.800 ;
        RECT 423.000 416.850 423.900 417.600 ;
        RECT 428.100 417.000 429.900 417.600 ;
        RECT 422.100 415.050 423.900 416.850 ;
        RECT 425.100 415.800 426.900 416.400 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 425.100 414.600 433.050 415.800 ;
        RECT 430.950 412.950 433.050 414.600 ;
        RECT 429.450 407.700 431.250 408.000 ;
        RECT 420.150 407.100 431.250 407.700 ;
        RECT 420.150 406.500 437.850 407.100 ;
        RECT 420.150 405.600 421.050 406.500 ;
        RECT 429.450 406.200 437.850 406.500 ;
        RECT 409.800 393.600 411.600 399.600 ;
        RECT 412.800 393.000 414.600 399.600 ;
        RECT 420.150 393.600 421.950 405.600 ;
        RECT 434.250 404.700 436.050 405.300 ;
        RECT 428.550 403.500 436.050 404.700 ;
        RECT 436.950 404.100 437.850 406.200 ;
        RECT 439.950 406.200 440.850 418.800 ;
        RECT 452.250 415.050 453.450 422.400 ;
        RECT 464.400 421.200 466.200 428.400 ;
        RECT 469.500 422.400 471.300 429.000 ;
        RECT 481.800 422.400 483.600 429.000 ;
        RECT 484.800 421.500 486.600 428.400 ;
        RECT 487.800 422.400 489.600 429.000 ;
        RECT 490.800 421.500 492.600 428.400 ;
        RECT 493.800 422.400 495.600 429.000 ;
        RECT 496.800 421.500 498.600 428.400 ;
        RECT 499.800 422.400 501.600 429.000 ;
        RECT 502.800 421.500 504.600 428.400 ;
        RECT 505.800 422.400 507.600 429.000 ;
        RECT 515.400 422.400 517.200 429.000 ;
        RECT 464.400 420.300 468.600 421.200 ;
        RECT 464.100 415.200 465.900 417.000 ;
        RECT 467.400 415.200 468.600 420.300 ;
        RECT 483.900 420.300 486.600 421.500 ;
        RECT 488.700 420.300 492.600 421.500 ;
        RECT 494.700 420.300 498.600 421.500 ;
        RECT 500.700 420.300 504.600 421.500 ;
        RECT 518.400 421.500 520.200 428.400 ;
        RECT 521.400 422.400 523.200 429.000 ;
        RECT 524.400 421.500 526.200 428.400 ;
        RECT 527.400 422.400 529.200 429.000 ;
        RECT 530.400 421.500 532.200 428.400 ;
        RECT 533.400 422.400 535.200 429.000 ;
        RECT 536.400 421.500 538.200 428.400 ;
        RECT 539.400 422.400 541.200 429.000 ;
        RECT 555.300 424.200 557.100 428.400 ;
        RECT 554.400 422.400 557.100 424.200 ;
        RECT 558.300 422.400 560.100 429.000 ;
        RECT 518.400 420.300 522.300 421.500 ;
        RECT 524.400 420.300 528.300 421.500 ;
        RECT 530.400 420.300 534.300 421.500 ;
        RECT 536.400 420.300 539.100 421.500 ;
        RECT 470.100 415.200 471.900 417.000 ;
        RECT 483.900 415.200 484.800 420.300 ;
        RECT 488.700 419.400 489.900 420.300 ;
        RECT 494.700 419.400 495.900 420.300 ;
        RECT 500.700 419.400 501.900 420.300 ;
        RECT 485.700 418.200 489.900 419.400 ;
        RECT 485.700 417.600 487.500 418.200 ;
        RECT 447.150 413.250 453.450 415.050 ;
        RECT 448.950 412.950 453.450 413.250 ;
        RECT 463.950 413.100 466.050 415.200 ;
        RECT 466.950 413.100 469.050 415.200 ;
        RECT 469.950 413.100 472.050 415.200 ;
        RECT 481.950 413.100 484.800 415.200 ;
        RECT 449.250 407.400 451.050 409.200 ;
        RECT 445.950 406.200 450.150 407.400 ;
        RECT 439.950 405.300 445.050 406.200 ;
        RECT 445.950 405.300 448.050 406.200 ;
        RECT 452.250 405.600 453.450 412.950 ;
        RECT 444.150 404.400 445.050 405.300 ;
        RECT 441.450 404.100 443.250 404.400 ;
        RECT 428.550 402.600 429.750 403.500 ;
        RECT 436.950 403.200 443.250 404.100 ;
        RECT 441.450 402.600 443.250 403.200 ;
        RECT 444.150 402.600 446.850 404.400 ;
        RECT 424.950 400.500 429.750 402.600 ;
        RECT 432.450 401.550 434.250 402.300 ;
        RECT 437.250 401.550 439.050 402.300 ;
        RECT 432.450 400.500 439.050 401.550 ;
        RECT 428.550 399.600 429.750 400.500 ;
        RECT 423.150 393.000 424.950 399.600 ;
        RECT 428.550 393.600 430.350 399.600 ;
        RECT 433.350 393.000 435.150 399.600 ;
        RECT 436.350 393.600 438.150 400.500 ;
        RECT 444.150 399.600 448.050 401.700 ;
        RECT 439.950 393.000 441.750 399.600 ;
        RECT 444.150 393.600 445.950 399.600 ;
        RECT 448.650 393.000 450.450 396.600 ;
        RECT 451.650 393.600 453.450 405.600 ;
        RECT 467.400 399.600 468.600 413.100 ;
        RECT 483.900 407.700 484.800 413.100 ;
        RECT 488.700 407.700 489.900 418.200 ;
        RECT 491.700 418.200 495.900 419.400 ;
        RECT 491.700 417.600 493.500 418.200 ;
        RECT 494.700 407.700 495.900 418.200 ;
        RECT 497.700 418.200 501.900 419.400 ;
        RECT 497.700 417.600 499.500 418.200 ;
        RECT 500.700 407.700 501.900 418.200 ;
        RECT 521.100 419.400 522.300 420.300 ;
        RECT 527.100 419.400 528.300 420.300 ;
        RECT 533.100 419.400 534.300 420.300 ;
        RECT 521.100 418.200 525.300 419.400 ;
        RECT 503.100 415.200 504.900 417.000 ;
        RECT 518.100 415.200 519.900 417.000 ;
        RECT 502.950 413.100 505.050 415.200 ;
        RECT 517.950 413.100 520.050 415.200 ;
        RECT 521.100 407.700 522.300 418.200 ;
        RECT 523.500 417.600 525.300 418.200 ;
        RECT 527.100 418.200 531.300 419.400 ;
        RECT 527.100 407.700 528.300 418.200 ;
        RECT 529.500 417.600 531.300 418.200 ;
        RECT 533.100 418.200 537.300 419.400 ;
        RECT 533.100 407.700 534.300 418.200 ;
        RECT 535.500 417.600 537.300 418.200 ;
        RECT 538.200 415.200 539.100 420.300 ;
        RECT 554.400 415.200 555.300 422.400 ;
        RECT 557.100 420.600 558.900 421.500 ;
        RECT 562.800 420.600 564.600 428.400 ;
        RECT 572.400 425.400 574.200 428.400 ;
        RECT 575.400 425.400 577.200 429.000 ;
        RECT 572.400 421.500 573.600 425.400 ;
        RECT 578.400 422.400 580.200 428.400 ;
        RECT 590.400 425.400 592.200 429.000 ;
        RECT 593.400 425.400 595.200 428.400 ;
        RECT 605.400 425.400 607.200 429.000 ;
        RECT 608.400 425.400 610.200 428.400 ;
        RECT 611.400 425.400 613.200 429.000 ;
        RECT 572.400 420.600 578.100 421.500 ;
        RECT 557.100 419.700 564.600 420.600 ;
        RECT 576.150 419.700 578.100 420.600 ;
        RECT 538.200 413.100 541.050 415.200 ;
        RECT 553.950 413.100 556.050 415.200 ;
        RECT 556.950 413.100 559.050 415.200 ;
        RECT 538.200 407.700 539.100 413.100 ;
        RECT 483.900 406.500 486.600 407.700 ;
        RECT 488.700 406.500 492.600 407.700 ;
        RECT 494.700 406.500 498.600 407.700 ;
        RECT 500.700 406.500 504.600 407.700 ;
        RECT 463.800 393.000 465.600 399.600 ;
        RECT 466.800 393.600 468.600 399.600 ;
        RECT 469.800 393.000 471.600 399.600 ;
        RECT 481.800 393.000 483.600 405.600 ;
        RECT 484.800 393.600 486.600 406.500 ;
        RECT 487.800 393.000 489.600 405.600 ;
        RECT 490.800 393.600 492.600 406.500 ;
        RECT 493.800 393.000 495.600 405.600 ;
        RECT 496.800 393.600 498.600 406.500 ;
        RECT 499.800 393.000 501.600 405.600 ;
        RECT 502.800 393.600 504.600 406.500 ;
        RECT 518.400 406.500 522.300 407.700 ;
        RECT 524.400 406.500 528.300 407.700 ;
        RECT 530.400 406.500 534.300 407.700 ;
        RECT 536.400 406.500 539.100 407.700 ;
        RECT 505.800 393.000 507.600 405.600 ;
        RECT 515.400 393.000 517.200 405.600 ;
        RECT 518.400 393.600 520.200 406.500 ;
        RECT 521.400 393.000 523.200 405.600 ;
        RECT 524.400 393.600 526.200 406.500 ;
        RECT 527.400 393.000 529.200 405.600 ;
        RECT 530.400 393.600 532.200 406.500 ;
        RECT 533.400 393.000 535.200 405.600 ;
        RECT 536.400 393.600 538.200 406.500 ;
        RECT 554.400 405.600 555.300 413.100 ;
        RECT 557.100 411.300 558.900 413.100 ;
        RECT 539.400 393.000 541.200 405.600 ;
        RECT 553.800 393.600 555.600 405.600 ;
        RECT 560.700 399.600 561.600 419.700 ;
        RECT 563.100 415.200 564.900 417.000 ;
        RECT 562.950 413.100 565.050 415.200 ;
        RECT 571.950 412.950 574.050 415.050 ;
        RECT 572.100 411.150 573.900 412.950 ;
        RECT 576.150 408.300 577.050 419.700 ;
        RECT 579.000 415.050 580.200 422.400 ;
        RECT 593.400 415.050 594.600 425.400 ;
        RECT 600.000 417.450 604.050 418.050 ;
        RECT 599.550 415.950 604.050 417.450 ;
        RECT 577.950 412.950 580.200 415.050 ;
        RECT 589.950 412.950 592.050 415.050 ;
        RECT 592.950 412.950 595.050 415.050 ;
        RECT 576.150 407.400 578.100 408.300 ;
        RECT 572.400 406.500 578.100 407.400 ;
        RECT 572.400 399.600 573.600 406.500 ;
        RECT 579.000 405.600 580.200 412.950 ;
        RECT 590.100 411.150 591.900 412.950 ;
        RECT 556.800 393.000 558.600 399.600 ;
        RECT 559.800 393.600 561.600 399.600 ;
        RECT 562.800 393.000 564.600 399.600 ;
        RECT 572.400 393.600 574.200 399.600 ;
        RECT 575.400 393.000 577.200 399.600 ;
        RECT 578.400 393.600 580.200 405.600 ;
        RECT 593.400 399.600 594.600 412.950 ;
        RECT 599.550 412.050 600.450 415.950 ;
        RECT 608.700 415.050 609.600 425.400 ;
        RECT 623.400 423.300 625.200 428.400 ;
        RECT 626.400 424.200 628.200 429.000 ;
        RECT 629.400 423.300 631.200 428.400 ;
        RECT 623.400 421.950 631.200 423.300 ;
        RECT 632.400 422.400 634.200 428.400 ;
        RECT 638.550 422.400 640.350 428.400 ;
        RECT 641.850 425.400 643.650 429.000 ;
        RECT 646.650 425.400 648.450 428.400 ;
        RECT 650.850 425.400 652.650 429.000 ;
        RECT 654.450 425.400 656.250 428.400 ;
        RECT 657.750 425.400 659.550 429.000 ;
        RECT 662.250 426.300 664.050 428.400 ;
        RECT 662.250 425.400 666.000 426.300 ;
        RECT 667.050 425.400 668.850 429.000 ;
        RECT 646.650 424.500 647.700 425.400 ;
        RECT 643.950 423.300 647.700 424.500 ;
        RECT 655.200 424.500 656.250 425.400 ;
        RECT 664.950 424.500 666.000 425.400 ;
        RECT 655.200 423.450 660.150 424.500 ;
        RECT 643.950 422.400 646.050 423.300 ;
        RECT 658.350 422.700 660.150 423.450 ;
        RECT 632.400 420.300 633.600 422.400 ;
        RECT 629.850 419.250 633.600 420.300 ;
        RECT 626.100 415.050 627.900 416.850 ;
        RECT 629.850 415.050 631.050 419.250 ;
        RECT 632.100 415.050 633.900 416.850 ;
        RECT 638.550 415.050 639.750 422.400 ;
        RECT 661.650 421.800 663.450 423.600 ;
        RECT 664.950 422.400 667.050 424.500 ;
        RECT 670.050 422.400 671.850 428.400 ;
        RECT 680.700 422.400 682.500 429.000 ;
        RECT 651.150 420.000 652.950 420.600 ;
        RECT 662.100 420.000 663.150 421.800 ;
        RECT 651.150 418.800 663.150 420.000 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 638.550 413.250 644.850 415.050 ;
        RECT 638.550 412.950 643.050 413.250 ;
        RECT 599.550 410.550 604.050 412.050 ;
        RECT 605.100 411.150 606.900 412.950 ;
        RECT 600.000 409.950 604.050 410.550 ;
        RECT 608.700 405.600 609.600 412.950 ;
        RECT 611.100 411.150 612.900 412.950 ;
        RECT 623.100 411.150 624.900 412.950 ;
        RECT 590.400 393.000 592.200 399.600 ;
        RECT 593.400 393.600 595.200 399.600 ;
        RECT 605.400 393.000 607.200 405.600 ;
        RECT 608.700 404.400 612.300 405.600 ;
        RECT 610.500 393.600 612.300 404.400 ;
        RECT 623.700 393.000 625.500 405.600 ;
        RECT 628.950 399.600 630.150 412.950 ;
        RECT 638.550 405.600 639.750 412.950 ;
        RECT 640.950 407.400 642.750 409.200 ;
        RECT 641.850 406.200 646.050 407.400 ;
        RECT 651.150 406.200 652.050 418.800 ;
        RECT 662.100 417.600 669.000 418.800 ;
        RECT 662.100 417.000 663.900 417.600 ;
        RECT 668.100 416.850 669.000 417.600 ;
        RECT 665.100 415.800 666.900 416.400 ;
        RECT 658.950 414.600 666.900 415.800 ;
        RECT 668.100 415.050 669.900 416.850 ;
        RECT 658.950 412.950 661.050 414.600 ;
        RECT 667.950 412.950 670.050 415.050 ;
        RECT 660.750 407.700 662.550 408.000 ;
        RECT 670.950 407.700 671.850 422.400 ;
        RECT 685.800 421.200 687.600 428.400 ;
        RECT 698.400 423.300 700.200 428.400 ;
        RECT 701.400 424.200 703.200 429.000 ;
        RECT 704.400 423.300 706.200 428.400 ;
        RECT 698.400 421.950 706.200 423.300 ;
        RECT 707.400 422.400 709.200 428.400 ;
        RECT 721.800 422.400 723.600 428.400 ;
        RECT 683.400 420.300 687.600 421.200 ;
        RECT 707.400 420.300 708.600 422.400 ;
        RECT 680.100 415.200 681.900 417.000 ;
        RECT 683.400 415.200 684.600 420.300 ;
        RECT 704.850 419.250 708.600 420.300 ;
        RECT 722.400 420.300 723.600 422.400 ;
        RECT 724.800 423.300 726.600 428.400 ;
        RECT 727.800 424.200 729.600 429.000 ;
        RECT 730.800 423.300 732.600 428.400 ;
        RECT 724.800 421.950 732.600 423.300 ;
        RECT 743.400 421.200 745.200 428.400 ;
        RECT 748.500 422.400 750.300 429.000 ;
        RECT 743.400 420.300 747.600 421.200 ;
        RECT 722.400 419.250 726.150 420.300 ;
        RECT 686.100 415.200 687.900 417.000 ;
        RECT 679.950 413.100 682.050 415.200 ;
        RECT 682.950 413.100 685.050 415.200 ;
        RECT 685.950 413.100 688.050 415.200 ;
        RECT 701.100 415.050 702.900 416.850 ;
        RECT 704.850 415.050 706.050 419.250 ;
        RECT 717.000 417.450 721.050 418.050 ;
        RECT 707.100 415.050 708.900 416.850 ;
        RECT 716.550 415.950 721.050 417.450 ;
        RECT 660.750 407.100 671.850 407.700 ;
        RECT 628.800 393.600 630.600 399.600 ;
        RECT 631.800 393.000 633.600 399.600 ;
        RECT 638.550 393.600 640.350 405.600 ;
        RECT 643.950 405.300 646.050 406.200 ;
        RECT 646.950 405.300 652.050 406.200 ;
        RECT 654.150 406.500 671.850 407.100 ;
        RECT 654.150 406.200 662.550 406.500 ;
        RECT 646.950 404.400 647.850 405.300 ;
        RECT 645.150 402.600 647.850 404.400 ;
        RECT 648.750 404.100 650.550 404.400 ;
        RECT 654.150 404.100 655.050 406.200 ;
        RECT 670.950 405.600 671.850 406.500 ;
        RECT 648.750 403.200 655.050 404.100 ;
        RECT 655.950 404.700 657.750 405.300 ;
        RECT 655.950 403.500 663.450 404.700 ;
        RECT 648.750 402.600 650.550 403.200 ;
        RECT 662.250 402.600 663.450 403.500 ;
        RECT 643.950 399.600 647.850 401.700 ;
        RECT 652.950 401.550 654.750 402.300 ;
        RECT 657.750 401.550 659.550 402.300 ;
        RECT 652.950 400.500 659.550 401.550 ;
        RECT 662.250 400.500 667.050 402.600 ;
        RECT 641.550 393.000 643.350 396.600 ;
        RECT 646.050 393.600 647.850 399.600 ;
        RECT 650.250 393.000 652.050 399.600 ;
        RECT 653.850 393.600 655.650 400.500 ;
        RECT 662.250 399.600 663.450 400.500 ;
        RECT 656.850 393.000 658.650 399.600 ;
        RECT 661.650 393.600 663.450 399.600 ;
        RECT 667.050 393.000 668.850 399.600 ;
        RECT 670.050 393.600 671.850 405.600 ;
        RECT 683.400 399.600 684.600 413.100 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 706.950 412.950 709.050 415.050 ;
        RECT 698.100 411.150 699.900 412.950 ;
        RECT 680.400 393.000 682.200 399.600 ;
        RECT 683.400 393.600 685.200 399.600 ;
        RECT 686.400 393.000 688.200 399.600 ;
        RECT 698.700 393.000 700.500 405.600 ;
        RECT 703.950 399.600 705.150 412.950 ;
        RECT 716.550 412.050 717.450 415.950 ;
        RECT 722.100 415.050 723.900 416.850 ;
        RECT 724.950 415.050 726.150 419.250 ;
        RECT 728.100 415.050 729.900 416.850 ;
        RECT 743.100 415.200 744.900 417.000 ;
        RECT 746.400 415.200 747.600 420.300 ;
        RECT 758.400 419.400 760.200 429.000 ;
        RECT 765.000 420.000 766.800 428.400 ;
        RECT 765.000 418.800 768.300 420.000 ;
        RECT 779.400 419.400 781.200 429.000 ;
        RECT 786.000 420.000 787.800 428.400 ;
        RECT 786.000 418.800 789.300 420.000 ;
        RECT 800.400 419.400 802.200 429.000 ;
        RECT 807.000 420.000 808.800 428.400 ;
        RECT 821.400 425.400 823.200 429.000 ;
        RECT 824.400 425.400 826.200 428.400 ;
        RECT 836.400 425.400 838.200 428.400 ;
        RECT 839.400 425.400 841.200 429.000 ;
        RECT 807.000 418.800 810.300 420.000 ;
        RECT 749.100 415.200 750.900 417.000 ;
        RECT 758.100 415.200 759.900 417.000 ;
        RECT 764.100 415.200 765.900 417.000 ;
        RECT 767.400 415.200 768.300 418.800 ;
        RECT 774.000 417.450 778.050 418.050 ;
        RECT 773.550 415.950 778.050 417.450 ;
        RECT 721.950 412.950 724.050 415.050 ;
        RECT 724.950 412.950 727.050 415.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 742.950 413.100 745.050 415.200 ;
        RECT 745.950 413.100 748.050 415.200 ;
        RECT 748.950 413.100 751.050 415.200 ;
        RECT 757.950 413.100 760.050 415.200 ;
        RECT 760.950 413.100 763.050 415.200 ;
        RECT 763.950 413.100 766.050 415.200 ;
        RECT 766.950 413.100 769.050 415.200 ;
        RECT 716.550 410.550 721.050 412.050 ;
        RECT 717.000 409.950 721.050 410.550 ;
        RECT 725.850 399.600 727.050 412.950 ;
        RECT 731.100 411.150 732.900 412.950 ;
        RECT 703.800 393.600 705.600 399.600 ;
        RECT 706.800 393.000 708.600 399.600 ;
        RECT 722.400 393.000 724.200 399.600 ;
        RECT 725.400 393.600 727.200 399.600 ;
        RECT 730.500 393.000 732.300 405.600 ;
        RECT 746.400 399.600 747.600 413.100 ;
        RECT 761.100 411.300 762.900 413.100 ;
        RECT 767.400 400.800 768.300 413.100 ;
        RECT 773.550 411.450 774.450 415.950 ;
        RECT 779.100 415.200 780.900 417.000 ;
        RECT 785.100 415.200 786.900 417.000 ;
        RECT 788.400 415.200 789.300 418.800 ;
        RECT 800.100 415.200 801.900 417.000 ;
        RECT 806.100 415.200 807.900 417.000 ;
        RECT 809.400 415.200 810.300 418.800 ;
        RECT 811.950 417.450 816.000 418.050 ;
        RECT 811.950 415.950 816.450 417.450 ;
        RECT 778.950 413.100 781.050 415.200 ;
        RECT 781.950 413.100 784.050 415.200 ;
        RECT 784.950 413.100 787.050 415.200 ;
        RECT 787.950 413.100 790.050 415.200 ;
        RECT 799.950 413.100 802.050 415.200 ;
        RECT 802.950 413.100 805.050 415.200 ;
        RECT 805.950 413.100 808.050 415.200 ;
        RECT 808.950 413.100 811.050 415.200 ;
        RECT 770.550 411.000 780.450 411.450 ;
        RECT 782.100 411.300 783.900 413.100 ;
        RECT 769.950 410.550 780.450 411.000 ;
        RECT 769.950 406.950 772.050 410.550 ;
        RECT 779.550 408.450 780.450 410.550 ;
        RECT 784.950 408.450 787.050 409.050 ;
        RECT 779.550 407.550 787.050 408.450 ;
        RECT 784.950 406.950 787.050 407.550 ;
        RECT 788.400 400.800 789.300 413.100 ;
        RECT 803.100 411.300 804.900 413.100 ;
        RECT 809.400 400.800 810.300 413.100 ;
        RECT 815.550 412.050 816.450 415.950 ;
        RECT 824.400 415.050 825.600 425.400 ;
        RECT 836.400 421.500 837.600 425.400 ;
        RECT 842.400 422.400 844.200 428.400 ;
        RECT 836.400 420.600 842.100 421.500 ;
        RECT 840.150 419.700 842.100 420.600 ;
        RECT 826.950 417.450 831.000 418.050 ;
        RECT 826.950 415.950 831.450 417.450 ;
        RECT 820.950 412.950 823.050 415.050 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 815.550 410.550 820.050 412.050 ;
        RECT 821.100 411.150 822.900 412.950 ;
        RECT 816.000 409.950 820.050 410.550 ;
        RECT 761.700 399.900 768.300 400.800 ;
        RECT 761.700 399.600 763.200 399.900 ;
        RECT 742.800 393.000 744.600 399.600 ;
        RECT 745.800 393.600 747.600 399.600 ;
        RECT 748.800 393.000 750.600 399.600 ;
        RECT 758.400 393.000 760.200 399.600 ;
        RECT 761.400 393.600 763.200 399.600 ;
        RECT 767.400 399.600 768.300 399.900 ;
        RECT 782.700 399.900 789.300 400.800 ;
        RECT 782.700 399.600 784.200 399.900 ;
        RECT 764.400 393.000 766.200 399.000 ;
        RECT 767.400 393.600 769.200 399.600 ;
        RECT 779.400 393.000 781.200 399.600 ;
        RECT 782.400 393.600 784.200 399.600 ;
        RECT 788.400 399.600 789.300 399.900 ;
        RECT 803.700 399.900 810.300 400.800 ;
        RECT 803.700 399.600 805.200 399.900 ;
        RECT 785.400 393.000 787.200 399.000 ;
        RECT 788.400 393.600 790.200 399.600 ;
        RECT 800.400 393.000 802.200 399.600 ;
        RECT 803.400 393.600 805.200 399.600 ;
        RECT 809.400 399.600 810.300 399.900 ;
        RECT 824.400 399.600 825.600 412.950 ;
        RECT 830.550 412.050 831.450 415.950 ;
        RECT 835.950 412.950 838.050 415.050 ;
        RECT 826.950 410.550 831.450 412.050 ;
        RECT 836.100 411.150 837.900 412.950 ;
        RECT 826.950 409.950 831.000 410.550 ;
        RECT 840.150 408.300 841.050 419.700 ;
        RECT 843.000 415.050 844.200 422.400 ;
        RECT 841.950 412.950 844.200 415.050 ;
        RECT 840.150 407.400 842.100 408.300 ;
        RECT 836.400 406.500 842.100 407.400 ;
        RECT 836.400 399.600 837.600 406.500 ;
        RECT 843.000 405.600 844.200 412.950 ;
        RECT 806.400 393.000 808.200 399.000 ;
        RECT 809.400 393.600 811.200 399.600 ;
        RECT 821.400 393.000 823.200 399.600 ;
        RECT 824.400 393.600 826.200 399.600 ;
        RECT 836.400 393.600 838.200 399.600 ;
        RECT 839.400 393.000 841.200 399.600 ;
        RECT 842.400 393.600 844.200 405.600 ;
        RECT 10.800 383.400 12.600 389.400 ;
        RECT 13.800 384.000 15.600 390.000 ;
        RECT 11.700 383.100 12.600 383.400 ;
        RECT 16.800 383.400 18.600 389.400 ;
        RECT 19.800 383.400 21.600 390.000 ;
        RECT 16.800 383.100 18.300 383.400 ;
        RECT 11.700 382.200 18.300 383.100 ;
        RECT 11.700 369.900 12.600 382.200 ;
        RECT 29.400 378.300 31.200 389.400 ;
        RECT 32.400 379.200 34.200 390.000 ;
        RECT 35.400 378.300 37.200 389.400 ;
        RECT 29.400 377.400 37.200 378.300 ;
        RECT 38.400 377.400 40.200 389.400 ;
        RECT 45.150 377.400 46.950 389.400 ;
        RECT 48.150 383.400 49.950 390.000 ;
        RECT 53.550 383.400 55.350 389.400 ;
        RECT 58.350 383.400 60.150 390.000 ;
        RECT 53.550 382.500 54.750 383.400 ;
        RECT 61.350 382.500 63.150 389.400 ;
        RECT 64.950 383.400 66.750 390.000 ;
        RECT 69.150 383.400 70.950 389.400 ;
        RECT 73.650 386.400 75.450 390.000 ;
        RECT 49.950 380.400 54.750 382.500 ;
        RECT 57.450 381.450 64.050 382.500 ;
        RECT 57.450 380.700 59.250 381.450 ;
        RECT 62.250 380.700 64.050 381.450 ;
        RECT 69.150 381.300 73.050 383.400 ;
        RECT 53.550 379.500 54.750 380.400 ;
        RECT 66.450 379.800 68.250 380.400 ;
        RECT 53.550 378.300 61.050 379.500 ;
        RECT 59.250 377.700 61.050 378.300 ;
        RECT 61.950 378.900 68.250 379.800 ;
        RECT 13.950 375.450 16.050 376.050 ;
        RECT 34.950 375.450 37.050 376.050 ;
        RECT 13.950 374.550 37.050 375.450 ;
        RECT 13.950 373.950 16.050 374.550 ;
        RECT 34.950 373.950 37.050 374.550 ;
        RECT 17.100 369.900 18.900 371.700 ;
        RECT 32.100 369.900 33.900 371.700 ;
        RECT 38.700 369.900 39.600 377.400 ;
        RECT 45.150 376.500 46.050 377.400 ;
        RECT 61.950 376.800 62.850 378.900 ;
        RECT 66.450 378.600 68.250 378.900 ;
        RECT 69.150 378.600 71.850 380.400 ;
        RECT 69.150 377.700 70.050 378.600 ;
        RECT 54.450 376.500 62.850 376.800 ;
        RECT 45.150 375.900 62.850 376.500 ;
        RECT 64.950 376.800 70.050 377.700 ;
        RECT 70.950 376.800 73.050 377.700 ;
        RECT 76.650 377.400 78.450 389.400 ;
        RECT 88.800 377.400 90.600 389.400 ;
        RECT 91.800 378.300 93.600 389.400 ;
        RECT 94.800 379.200 96.600 390.000 ;
        RECT 97.800 378.300 99.600 389.400 ;
        RECT 109.800 383.400 111.600 389.400 ;
        RECT 112.800 384.000 114.600 390.000 ;
        RECT 91.800 377.400 99.600 378.300 ;
        RECT 110.700 383.100 111.600 383.400 ;
        RECT 115.800 383.400 117.600 389.400 ;
        RECT 118.800 383.400 120.600 390.000 ;
        RECT 115.800 383.100 117.300 383.400 ;
        RECT 110.700 382.200 117.300 383.100 ;
        RECT 45.150 375.300 56.250 375.900 ;
        RECT 10.950 367.800 13.050 369.900 ;
        RECT 13.950 367.800 16.050 369.900 ;
        RECT 16.950 367.800 19.050 369.900 ;
        RECT 19.950 367.800 22.050 369.900 ;
        RECT 28.950 367.800 31.050 369.900 ;
        RECT 31.950 367.800 34.050 369.900 ;
        RECT 34.950 367.800 37.050 369.900 ;
        RECT 37.950 367.800 40.050 369.900 ;
        RECT 11.700 364.200 12.600 367.800 ;
        RECT 14.100 366.000 15.900 367.800 ;
        RECT 20.100 366.000 21.900 367.800 ;
        RECT 29.100 366.000 30.900 367.800 ;
        RECT 35.100 366.000 36.900 367.800 ;
        RECT 11.700 363.000 15.000 364.200 ;
        RECT 13.200 354.600 15.000 363.000 ;
        RECT 19.800 354.000 21.600 363.600 ;
        RECT 38.700 360.600 39.600 367.800 ;
        RECT 30.000 354.000 31.800 360.600 ;
        RECT 34.500 359.400 39.600 360.600 ;
        RECT 45.150 360.600 46.050 375.300 ;
        RECT 54.450 375.000 56.250 375.300 ;
        RECT 46.950 367.950 49.050 370.050 ;
        RECT 55.950 368.400 58.050 370.050 ;
        RECT 47.100 366.150 48.900 367.950 ;
        RECT 50.100 367.200 58.050 368.400 ;
        RECT 50.100 366.600 51.900 367.200 ;
        RECT 48.000 365.400 48.900 366.150 ;
        RECT 53.100 365.400 54.900 366.000 ;
        RECT 48.000 364.200 54.900 365.400 ;
        RECT 64.950 364.200 65.850 376.800 ;
        RECT 70.950 375.600 75.150 376.800 ;
        RECT 74.250 373.800 76.050 375.600 ;
        RECT 77.250 370.050 78.450 377.400 ;
        RECT 73.950 369.750 78.450 370.050 ;
        RECT 89.400 369.900 90.300 377.400 ;
        RECT 95.100 369.900 96.900 371.700 ;
        RECT 110.700 369.900 111.600 382.200 ;
        RECT 131.700 378.600 133.500 389.400 ;
        RECT 131.700 377.400 135.300 378.600 ;
        RECT 136.800 377.400 138.600 390.000 ;
        RECT 148.800 378.600 150.600 389.400 ;
        RECT 148.800 377.400 153.900 378.600 ;
        RECT 156.300 378.300 158.100 389.400 ;
        RECT 163.800 378.300 165.600 389.400 ;
        RECT 175.800 383.400 177.600 390.000 ;
        RECT 178.800 383.400 180.600 389.400 ;
        RECT 181.800 383.400 183.600 390.000 ;
        RECT 191.400 383.400 193.200 390.000 ;
        RECT 194.400 383.400 196.200 389.400 ;
        RECT 116.100 369.900 117.900 371.700 ;
        RECT 131.100 370.050 132.900 371.850 ;
        RECT 134.400 370.050 135.300 377.400 ;
        RECT 151.800 376.500 153.900 377.400 ;
        RECT 154.800 377.400 158.100 378.300 ;
        RECT 142.950 372.450 145.050 373.050 ;
        RECT 154.800 372.900 156.000 377.400 ;
        RECT 160.800 377.100 165.600 378.300 ;
        RECT 160.800 376.200 162.900 377.100 ;
        RECT 157.650 375.300 162.900 376.200 ;
        RECT 157.650 373.200 159.450 375.300 ;
        RECT 137.100 370.050 138.900 371.850 ;
        RECT 142.950 371.700 150.450 372.450 ;
        RECT 154.650 372.300 156.750 372.900 ;
        RECT 142.950 371.550 150.900 371.700 ;
        RECT 142.950 370.950 145.050 371.550 ;
        RECT 72.150 367.950 78.450 369.750 ;
        RECT 53.850 363.000 65.850 364.200 ;
        RECT 53.850 361.200 54.900 363.000 ;
        RECT 64.050 362.400 65.850 363.000 ;
        RECT 34.500 354.600 36.300 359.400 ;
        RECT 37.500 354.000 39.300 357.600 ;
        RECT 45.150 354.600 46.950 360.600 ;
        RECT 49.950 358.500 52.050 360.600 ;
        RECT 53.550 359.400 55.350 361.200 ;
        RECT 77.250 360.600 78.450 367.950 ;
        RECT 88.950 367.800 91.050 369.900 ;
        RECT 91.950 367.800 94.050 369.900 ;
        RECT 94.950 367.800 97.050 369.900 ;
        RECT 97.950 367.800 100.050 369.900 ;
        RECT 109.950 367.800 112.050 369.900 ;
        RECT 112.950 367.800 115.050 369.900 ;
        RECT 115.950 367.800 118.050 369.900 ;
        RECT 118.950 367.800 121.050 369.900 ;
        RECT 130.950 367.950 133.050 370.050 ;
        RECT 133.950 367.950 136.050 370.050 ;
        RECT 136.950 367.950 139.050 370.050 ;
        RECT 149.100 369.900 150.900 371.550 ;
        RECT 154.650 370.800 157.650 372.300 ;
        RECT 56.850 359.550 58.650 360.300 ;
        RECT 70.950 359.700 73.050 360.600 ;
        RECT 56.850 358.500 61.800 359.550 ;
        RECT 51.000 357.600 52.050 358.500 ;
        RECT 60.750 357.600 61.800 358.500 ;
        RECT 69.300 358.500 73.050 359.700 ;
        RECT 69.300 357.600 70.350 358.500 ;
        RECT 48.150 354.000 49.950 357.600 ;
        RECT 51.000 356.700 54.750 357.600 ;
        RECT 52.950 354.600 54.750 356.700 ;
        RECT 57.450 354.000 59.250 357.600 ;
        RECT 60.750 354.600 62.550 357.600 ;
        RECT 64.350 354.000 66.150 357.600 ;
        RECT 68.550 354.600 70.350 357.600 ;
        RECT 73.350 354.000 75.150 357.600 ;
        RECT 76.650 354.600 78.450 360.600 ;
        RECT 89.400 360.600 90.300 367.800 ;
        RECT 92.100 366.000 93.900 367.800 ;
        RECT 98.100 366.000 99.900 367.800 ;
        RECT 110.700 364.200 111.600 367.800 ;
        RECT 113.100 366.000 114.900 367.800 ;
        RECT 119.100 366.000 120.900 367.800 ;
        RECT 110.700 363.000 114.000 364.200 ;
        RECT 89.400 359.400 94.500 360.600 ;
        RECT 89.700 354.000 91.500 357.600 ;
        RECT 92.700 354.600 94.500 359.400 ;
        RECT 97.200 354.000 99.000 360.600 ;
        RECT 112.200 354.600 114.000 363.000 ;
        RECT 118.800 354.000 120.600 363.600 ;
        RECT 134.400 357.600 135.300 367.950 ;
        RECT 148.950 367.800 151.050 369.900 ;
        RECT 153.900 368.100 155.700 369.900 ;
        RECT 153.750 366.000 155.850 368.100 ;
        RECT 156.750 364.200 157.650 370.800 ;
        RECT 159.000 370.200 160.800 372.000 ;
        RECT 158.700 368.100 160.800 370.200 ;
        RECT 179.400 369.900 180.600 383.400 ;
        RECT 191.100 370.050 192.900 371.850 ;
        RECT 194.400 370.050 195.600 383.400 ;
        RECT 201.150 377.400 202.950 389.400 ;
        RECT 204.150 383.400 205.950 390.000 ;
        RECT 209.550 383.400 211.350 389.400 ;
        RECT 214.350 383.400 216.150 390.000 ;
        RECT 209.550 382.500 210.750 383.400 ;
        RECT 217.350 382.500 219.150 389.400 ;
        RECT 220.950 383.400 222.750 390.000 ;
        RECT 225.150 383.400 226.950 389.400 ;
        RECT 229.650 386.400 231.450 390.000 ;
        RECT 205.950 380.400 210.750 382.500 ;
        RECT 213.450 381.450 220.050 382.500 ;
        RECT 213.450 380.700 215.250 381.450 ;
        RECT 218.250 380.700 220.050 381.450 ;
        RECT 225.150 381.300 229.050 383.400 ;
        RECT 209.550 379.500 210.750 380.400 ;
        RECT 222.450 379.800 224.250 380.400 ;
        RECT 209.550 378.300 217.050 379.500 ;
        RECT 215.250 377.700 217.050 378.300 ;
        RECT 217.950 378.900 224.250 379.800 ;
        RECT 201.150 376.500 202.050 377.400 ;
        RECT 217.950 376.800 218.850 378.900 ;
        RECT 222.450 378.600 224.250 378.900 ;
        RECT 225.150 378.600 227.850 380.400 ;
        RECT 225.150 377.700 226.050 378.600 ;
        RECT 210.450 376.500 218.850 376.800 ;
        RECT 201.150 375.900 218.850 376.500 ;
        RECT 220.950 376.800 226.050 377.700 ;
        RECT 226.950 376.800 229.050 377.700 ;
        RECT 232.650 377.400 234.450 389.400 ;
        RECT 242.400 383.400 244.200 390.000 ;
        RECT 245.400 383.400 247.200 389.400 ;
        RECT 248.400 383.400 250.200 390.000 ;
        RECT 201.150 375.300 212.250 375.900 ;
        RECT 163.950 367.800 166.050 369.900 ;
        RECT 175.950 367.800 178.050 369.900 ;
        RECT 178.950 367.800 181.050 369.900 ;
        RECT 181.950 367.800 184.050 369.900 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 163.950 367.200 165.750 367.800 ;
        RECT 158.700 366.000 165.750 367.200 ;
        RECT 176.100 366.000 177.900 367.800 ;
        RECT 158.700 365.100 160.800 366.000 ;
        RECT 151.200 361.500 153.300 363.900 ;
        RECT 154.650 362.100 157.650 364.200 ;
        RECT 158.550 363.300 160.350 365.100 ;
        RECT 148.800 360.600 153.300 361.500 ;
        RECT 130.800 354.000 132.600 357.600 ;
        RECT 133.800 354.600 135.600 357.600 ;
        RECT 136.800 354.000 138.600 357.600 ;
        RECT 148.800 354.600 150.600 360.600 ;
        RECT 156.750 360.000 157.650 362.100 ;
        RECT 161.250 363.000 163.350 363.600 ;
        RECT 161.250 361.500 165.600 363.000 ;
        RECT 179.400 362.700 180.600 367.800 ;
        RECT 182.100 366.000 183.900 367.800 ;
        RECT 164.100 360.600 165.600 361.500 ;
        RECT 156.600 354.600 158.400 360.000 ;
        RECT 163.800 354.600 165.600 360.600 ;
        RECT 176.400 361.800 180.600 362.700 ;
        RECT 176.400 354.600 178.200 361.800 ;
        RECT 181.500 354.000 183.300 360.600 ;
        RECT 194.400 357.600 195.600 367.950 ;
        RECT 201.150 360.600 202.050 375.300 ;
        RECT 210.450 375.000 212.250 375.300 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 211.950 368.400 214.050 370.050 ;
        RECT 203.100 366.150 204.900 367.950 ;
        RECT 206.100 367.200 214.050 368.400 ;
        RECT 206.100 366.600 207.900 367.200 ;
        RECT 204.000 365.400 204.900 366.150 ;
        RECT 209.100 365.400 210.900 366.000 ;
        RECT 204.000 364.200 210.900 365.400 ;
        RECT 220.950 364.200 221.850 376.800 ;
        RECT 226.950 375.600 231.150 376.800 ;
        RECT 230.250 373.800 232.050 375.600 ;
        RECT 233.250 370.050 234.450 377.400 ;
        RECT 229.950 369.750 234.450 370.050 ;
        RECT 228.150 367.950 234.450 369.750 ;
        RECT 209.850 363.000 221.850 364.200 ;
        RECT 209.850 361.200 210.900 363.000 ;
        RECT 220.050 362.400 221.850 363.000 ;
        RECT 191.400 354.000 193.200 357.600 ;
        RECT 194.400 354.600 196.200 357.600 ;
        RECT 201.150 354.600 202.950 360.600 ;
        RECT 205.950 358.500 208.050 360.600 ;
        RECT 209.550 359.400 211.350 361.200 ;
        RECT 233.250 360.600 234.450 367.950 ;
        RECT 241.950 367.800 244.050 369.900 ;
        RECT 242.100 366.000 243.900 367.800 ;
        RECT 245.400 363.300 246.300 383.400 ;
        RECT 251.400 377.400 253.200 389.400 ;
        RECT 263.400 383.400 265.200 390.000 ;
        RECT 266.400 383.400 268.200 389.400 ;
        RECT 248.100 369.900 249.900 371.700 ;
        RECT 251.700 369.900 252.600 377.400 ;
        RECT 263.100 370.050 264.900 371.850 ;
        RECT 266.400 370.050 267.600 383.400 ;
        RECT 278.400 377.400 280.200 390.000 ;
        RECT 282.900 377.400 286.200 389.400 ;
        RECT 288.900 377.400 290.700 390.000 ;
        RECT 305.700 378.600 307.500 389.400 ;
        RECT 305.700 377.400 309.300 378.600 ;
        RECT 310.800 377.400 312.600 390.000 ;
        RECT 320.700 377.400 322.500 390.000 ;
        RECT 325.800 383.400 327.600 389.400 ;
        RECT 328.800 383.400 330.600 390.000 ;
        RECT 344.400 383.400 346.200 390.000 ;
        RECT 347.400 383.400 349.200 389.400 ;
        RECT 247.950 367.800 250.050 369.900 ;
        RECT 250.950 367.800 253.050 369.900 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 278.100 369.900 279.900 371.700 ;
        RECT 284.100 369.900 285.300 377.400 ;
        RECT 290.100 369.900 291.900 371.700 ;
        RECT 305.100 370.050 306.900 371.850 ;
        RECT 308.400 370.050 309.300 377.400 ;
        RECT 311.100 370.050 312.900 371.850 ;
        RECT 320.100 370.050 321.900 371.850 ;
        RECT 325.950 370.050 327.150 383.400 ;
        RECT 347.850 370.050 349.050 383.400 ;
        RECT 352.500 377.400 354.300 390.000 ;
        RECT 362.700 377.400 364.500 390.000 ;
        RECT 367.800 383.400 369.600 389.400 ;
        RECT 370.800 383.400 372.600 390.000 ;
        RECT 383.400 383.400 385.200 390.000 ;
        RECT 386.400 383.400 388.200 389.400 ;
        RECT 353.100 370.050 354.900 371.850 ;
        RECT 362.100 370.050 363.900 371.850 ;
        RECT 367.950 370.050 369.150 383.400 ;
        RECT 383.100 370.050 384.900 371.850 ;
        RECT 386.400 370.050 387.600 383.400 ;
        RECT 400.800 377.400 402.600 389.400 ;
        RECT 403.800 383.400 405.600 390.000 ;
        RECT 406.800 383.400 408.600 389.400 ;
        RECT 400.800 370.050 402.000 377.400 ;
        RECT 407.400 376.500 408.600 383.400 ;
        RECT 418.800 377.400 420.600 389.400 ;
        RECT 421.800 383.400 423.600 390.000 ;
        RECT 424.800 383.400 426.600 389.400 ;
        RECT 427.800 383.400 429.600 390.000 ;
        RECT 402.900 375.600 408.600 376.500 ;
        RECT 402.900 374.700 404.850 375.600 ;
        RECT 212.850 359.550 214.650 360.300 ;
        RECT 226.950 359.700 229.050 360.600 ;
        RECT 212.850 358.500 217.800 359.550 ;
        RECT 207.000 357.600 208.050 358.500 ;
        RECT 216.750 357.600 217.800 358.500 ;
        RECT 225.300 358.500 229.050 359.700 ;
        RECT 225.300 357.600 226.350 358.500 ;
        RECT 204.150 354.000 205.950 357.600 ;
        RECT 207.000 356.700 210.750 357.600 ;
        RECT 208.950 354.600 210.750 356.700 ;
        RECT 213.450 354.000 215.250 357.600 ;
        RECT 216.750 354.600 218.550 357.600 ;
        RECT 220.350 354.000 222.150 357.600 ;
        RECT 224.550 354.600 226.350 357.600 ;
        RECT 229.350 354.000 231.150 357.600 ;
        RECT 232.650 354.600 234.450 360.600 ;
        RECT 242.400 362.400 249.900 363.300 ;
        RECT 242.400 354.600 244.200 362.400 ;
        RECT 248.100 361.500 249.900 362.400 ;
        RECT 251.700 360.600 252.600 367.800 ;
        RECT 246.900 354.000 248.700 360.600 ;
        RECT 249.900 358.800 252.600 360.600 ;
        RECT 249.900 354.600 251.700 358.800 ;
        RECT 266.400 357.600 267.600 367.950 ;
        RECT 277.950 367.800 280.050 369.900 ;
        RECT 280.950 367.800 283.050 369.900 ;
        RECT 283.950 367.800 286.050 369.900 ;
        RECT 286.950 367.800 289.050 369.900 ;
        RECT 289.950 367.800 292.050 369.900 ;
        RECT 304.950 367.950 307.050 370.050 ;
        RECT 307.950 367.950 310.050 370.050 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 322.950 367.950 325.050 370.050 ;
        RECT 325.950 367.950 328.050 370.050 ;
        RECT 328.950 367.950 331.050 370.050 ;
        RECT 343.950 367.950 346.050 370.050 ;
        RECT 346.950 367.950 349.050 370.050 ;
        RECT 349.950 367.950 352.050 370.050 ;
        RECT 352.950 367.950 355.050 370.050 ;
        RECT 361.950 367.950 364.050 370.050 ;
        RECT 364.950 367.950 367.050 370.050 ;
        RECT 367.950 367.950 370.050 370.050 ;
        RECT 370.950 367.950 373.050 370.050 ;
        RECT 382.950 367.950 385.050 370.050 ;
        RECT 385.950 367.950 388.050 370.050 ;
        RECT 400.800 367.950 403.050 370.050 ;
        RECT 281.100 366.000 282.900 367.800 ;
        RECT 283.950 365.400 285.000 367.800 ;
        RECT 287.100 366.000 288.900 367.800 ;
        RECT 284.100 363.300 285.300 365.400 ;
        RECT 284.100 362.100 288.600 363.300 ;
        RECT 278.400 360.000 286.200 360.900 ;
        RECT 287.700 360.600 288.600 362.100 ;
        RECT 263.400 354.000 265.200 357.600 ;
        RECT 266.400 354.600 268.200 357.600 ;
        RECT 278.400 354.600 280.200 360.000 ;
        RECT 281.400 354.000 283.200 359.100 ;
        RECT 284.400 355.500 286.200 360.000 ;
        RECT 287.400 356.400 289.200 360.600 ;
        RECT 290.400 355.500 292.200 360.600 ;
        RECT 308.400 357.600 309.300 367.950 ;
        RECT 323.100 366.150 324.900 367.950 ;
        RECT 326.850 363.750 328.050 367.950 ;
        RECT 329.100 366.150 330.900 367.950 ;
        RECT 344.100 366.150 345.900 367.950 ;
        RECT 346.950 363.750 348.150 367.950 ;
        RECT 350.100 366.150 351.900 367.950 ;
        RECT 365.100 366.150 366.900 367.950 ;
        RECT 326.850 362.700 330.600 363.750 ;
        RECT 320.400 359.700 328.200 361.050 ;
        RECT 284.400 354.600 292.200 355.500 ;
        RECT 304.800 354.000 306.600 357.600 ;
        RECT 307.800 354.600 309.600 357.600 ;
        RECT 310.800 354.000 312.600 357.600 ;
        RECT 320.400 354.600 322.200 359.700 ;
        RECT 323.400 354.000 325.200 358.800 ;
        RECT 326.400 354.600 328.200 359.700 ;
        RECT 329.400 360.600 330.600 362.700 ;
        RECT 344.400 362.700 348.150 363.750 ;
        RECT 368.850 363.750 370.050 367.950 ;
        RECT 371.100 366.150 372.900 367.950 ;
        RECT 368.850 362.700 372.600 363.750 ;
        RECT 344.400 360.600 345.600 362.700 ;
        RECT 329.400 354.600 331.200 360.600 ;
        RECT 343.800 354.600 345.600 360.600 ;
        RECT 346.800 359.700 354.600 361.050 ;
        RECT 346.800 354.600 348.600 359.700 ;
        RECT 349.800 354.000 351.600 358.800 ;
        RECT 352.800 354.600 354.600 359.700 ;
        RECT 362.400 359.700 370.200 361.050 ;
        RECT 362.400 354.600 364.200 359.700 ;
        RECT 365.400 354.000 367.200 358.800 ;
        RECT 368.400 354.600 370.200 359.700 ;
        RECT 371.400 360.600 372.600 362.700 ;
        RECT 371.400 354.600 373.200 360.600 ;
        RECT 386.400 357.600 387.600 367.950 ;
        RECT 400.800 360.600 402.000 367.950 ;
        RECT 403.950 363.300 404.850 374.700 ;
        RECT 407.100 370.050 408.900 371.850 ;
        RECT 406.950 367.950 409.050 370.050 ;
        RECT 419.400 369.900 420.300 377.400 ;
        RECT 422.100 369.900 423.900 371.700 ;
        RECT 418.950 367.800 421.050 369.900 ;
        RECT 421.950 367.800 424.050 369.900 ;
        RECT 402.900 362.400 404.850 363.300 ;
        RECT 402.900 361.500 408.600 362.400 ;
        RECT 383.400 354.000 385.200 357.600 ;
        RECT 386.400 354.600 388.200 357.600 ;
        RECT 400.800 354.600 402.600 360.600 ;
        RECT 407.400 357.600 408.600 361.500 ;
        RECT 419.400 360.600 420.300 367.800 ;
        RECT 425.700 363.300 426.600 383.400 ;
        RECT 441.300 378.900 443.100 389.400 ;
        RECT 440.700 377.400 443.100 378.900 ;
        RECT 444.300 377.400 446.100 390.000 ;
        RECT 448.800 377.400 450.600 389.400 ;
        RECT 458.400 383.400 460.200 390.000 ;
        RECT 461.400 383.400 463.200 389.400 ;
        RECT 464.400 383.400 466.200 390.000 ;
        RECT 479.400 383.400 481.200 390.000 ;
        RECT 482.400 383.400 484.200 389.400 ;
        RECT 427.950 372.450 430.050 373.050 ;
        RECT 436.950 372.450 439.050 373.050 ;
        RECT 427.950 371.550 439.050 372.450 ;
        RECT 427.950 370.950 430.050 371.550 ;
        RECT 436.950 370.950 439.050 371.550 ;
        RECT 440.700 370.050 442.050 377.400 ;
        RECT 449.400 375.900 450.600 377.400 ;
        RECT 427.950 367.800 430.050 369.900 ;
        RECT 439.950 367.950 442.050 370.050 ;
        RECT 443.400 374.700 450.600 375.900 ;
        RECT 443.400 374.100 445.200 374.700 ;
        RECT 428.100 366.000 429.900 367.800 ;
        RECT 422.100 362.400 429.600 363.300 ;
        RECT 422.100 361.500 423.900 362.400 ;
        RECT 419.400 358.800 422.100 360.600 ;
        RECT 403.800 354.000 405.600 357.600 ;
        RECT 406.800 354.600 408.600 357.600 ;
        RECT 420.300 354.600 422.100 358.800 ;
        RECT 423.300 354.000 425.100 360.600 ;
        RECT 427.800 354.600 429.600 362.400 ;
        RECT 439.950 360.600 441.000 367.950 ;
        RECT 443.400 363.600 444.300 374.100 ;
        RECT 451.950 372.450 454.050 373.050 ;
        RECT 457.950 372.450 460.050 373.050 ;
        RECT 446.100 370.050 447.900 371.850 ;
        RECT 451.950 371.550 460.050 372.450 ;
        RECT 451.950 370.950 454.050 371.550 ;
        RECT 457.950 370.950 460.050 371.550 ;
        RECT 445.950 367.950 448.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 461.400 369.900 462.600 383.400 ;
        RECT 474.000 372.450 478.050 373.050 ;
        RECT 473.550 370.950 478.050 372.450 ;
        RECT 449.100 366.150 450.900 367.950 ;
        RECT 457.950 367.800 460.050 369.900 ;
        RECT 460.950 367.800 463.050 369.900 ;
        RECT 463.950 367.800 466.050 369.900 ;
        RECT 458.100 366.000 459.900 367.800 ;
        RECT 443.400 362.700 445.200 363.600 ;
        RECT 461.400 362.700 462.600 367.800 ;
        RECT 464.100 366.000 465.900 367.800 ;
        RECT 473.550 367.050 474.450 370.950 ;
        RECT 482.850 370.050 484.050 383.400 ;
        RECT 487.500 377.400 489.300 390.000 ;
        RECT 497.400 383.400 499.200 390.000 ;
        RECT 500.400 383.400 502.200 389.400 ;
        RECT 503.400 383.400 505.200 390.000 ;
        RECT 488.100 370.050 489.900 371.850 ;
        RECT 478.950 367.950 481.050 370.050 ;
        RECT 481.950 367.950 484.050 370.050 ;
        RECT 484.950 367.950 487.050 370.050 ;
        RECT 487.950 367.950 490.050 370.050 ;
        RECT 500.400 369.900 501.600 383.400 ;
        RECT 509.550 377.400 511.350 389.400 ;
        RECT 512.550 386.400 514.350 390.000 ;
        RECT 517.050 383.400 518.850 389.400 ;
        RECT 521.250 383.400 523.050 390.000 ;
        RECT 514.950 381.300 518.850 383.400 ;
        RECT 524.850 382.500 526.650 389.400 ;
        RECT 527.850 383.400 529.650 390.000 ;
        RECT 532.650 383.400 534.450 389.400 ;
        RECT 538.050 383.400 539.850 390.000 ;
        RECT 533.250 382.500 534.450 383.400 ;
        RECT 523.950 381.450 530.550 382.500 ;
        RECT 523.950 380.700 525.750 381.450 ;
        RECT 528.750 380.700 530.550 381.450 ;
        RECT 533.250 380.400 538.050 382.500 ;
        RECT 516.150 378.600 518.850 380.400 ;
        RECT 519.750 379.800 521.550 380.400 ;
        RECT 519.750 378.900 526.050 379.800 ;
        RECT 533.250 379.500 534.450 380.400 ;
        RECT 519.750 378.600 521.550 378.900 ;
        RECT 517.950 377.700 518.850 378.600 ;
        RECT 509.550 370.050 510.750 377.400 ;
        RECT 514.950 376.800 517.050 377.700 ;
        RECT 517.950 376.800 523.050 377.700 ;
        RECT 512.850 375.600 517.050 376.800 ;
        RECT 511.950 373.800 513.750 375.600 ;
        RECT 473.550 365.550 478.050 367.050 ;
        RECT 479.100 366.150 480.900 367.950 ;
        RECT 474.000 364.950 478.050 365.550 ;
        RECT 481.950 363.750 483.150 367.950 ;
        RECT 485.100 366.150 486.900 367.950 ;
        RECT 496.950 367.800 499.050 369.900 ;
        RECT 499.950 367.800 502.050 369.900 ;
        RECT 502.950 367.800 505.050 369.900 ;
        RECT 509.550 369.750 514.050 370.050 ;
        RECT 509.550 367.950 515.850 369.750 ;
        RECT 497.100 366.000 498.900 367.800 ;
        RECT 479.400 362.700 483.150 363.750 ;
        RECT 500.400 362.700 501.600 367.800 ;
        RECT 503.100 366.000 504.900 367.800 ;
        RECT 443.400 361.800 446.700 362.700 ;
        RECT 461.400 361.800 465.600 362.700 ;
        RECT 439.800 354.600 441.600 360.600 ;
        RECT 445.800 357.600 446.700 361.800 ;
        RECT 442.800 354.000 444.600 357.600 ;
        RECT 445.800 354.600 447.600 357.600 ;
        RECT 448.800 354.600 450.600 357.600 ;
        RECT 449.400 354.000 450.600 354.600 ;
        RECT 458.700 354.000 460.500 360.600 ;
        RECT 463.800 354.600 465.600 361.800 ;
        RECT 479.400 360.600 480.600 362.700 ;
        RECT 500.400 361.800 504.600 362.700 ;
        RECT 478.800 354.600 480.600 360.600 ;
        RECT 481.800 359.700 489.600 361.050 ;
        RECT 481.800 354.600 483.600 359.700 ;
        RECT 484.800 354.000 486.600 358.800 ;
        RECT 487.800 354.600 489.600 359.700 ;
        RECT 497.700 354.000 499.500 360.600 ;
        RECT 502.800 354.600 504.600 361.800 ;
        RECT 509.550 360.600 510.750 367.950 ;
        RECT 522.150 364.200 523.050 376.800 ;
        RECT 525.150 376.800 526.050 378.900 ;
        RECT 526.950 378.300 534.450 379.500 ;
        RECT 526.950 377.700 528.750 378.300 ;
        RECT 541.050 377.400 542.850 389.400 ;
        RECT 525.150 376.500 533.550 376.800 ;
        RECT 541.950 376.500 542.850 377.400 ;
        RECT 525.150 375.900 542.850 376.500 ;
        RECT 531.750 375.300 542.850 375.900 ;
        RECT 531.750 375.000 533.550 375.300 ;
        RECT 529.950 368.400 532.050 370.050 ;
        RECT 529.950 367.200 537.900 368.400 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 536.100 366.600 537.900 367.200 ;
        RECT 539.100 366.150 540.900 367.950 ;
        RECT 533.100 365.400 534.900 366.000 ;
        RECT 539.100 365.400 540.000 366.150 ;
        RECT 533.100 364.200 540.000 365.400 ;
        RECT 522.150 363.000 534.150 364.200 ;
        RECT 522.150 362.400 523.950 363.000 ;
        RECT 533.100 361.200 534.150 363.000 ;
        RECT 509.550 354.600 511.350 360.600 ;
        RECT 514.950 359.700 517.050 360.600 ;
        RECT 514.950 358.500 518.700 359.700 ;
        RECT 529.350 359.550 531.150 360.300 ;
        RECT 517.650 357.600 518.700 358.500 ;
        RECT 526.200 358.500 531.150 359.550 ;
        RECT 532.650 359.400 534.450 361.200 ;
        RECT 541.950 360.600 542.850 375.300 ;
        RECT 535.950 358.500 538.050 360.600 ;
        RECT 526.200 357.600 527.250 358.500 ;
        RECT 535.950 357.600 537.000 358.500 ;
        RECT 512.850 354.000 514.650 357.600 ;
        RECT 517.650 354.600 519.450 357.600 ;
        RECT 521.850 354.000 523.650 357.600 ;
        RECT 525.450 354.600 527.250 357.600 ;
        RECT 528.750 354.000 530.550 357.600 ;
        RECT 533.250 356.700 537.000 357.600 ;
        RECT 533.250 354.600 535.050 356.700 ;
        RECT 538.050 354.000 539.850 357.600 ;
        RECT 541.050 354.600 542.850 360.600 ;
        RECT 546.150 377.400 547.950 389.400 ;
        RECT 549.150 383.400 550.950 390.000 ;
        RECT 554.550 383.400 556.350 389.400 ;
        RECT 559.350 383.400 561.150 390.000 ;
        RECT 554.550 382.500 555.750 383.400 ;
        RECT 562.350 382.500 564.150 389.400 ;
        RECT 565.950 383.400 567.750 390.000 ;
        RECT 570.150 383.400 571.950 389.400 ;
        RECT 574.650 386.400 576.450 390.000 ;
        RECT 550.950 380.400 555.750 382.500 ;
        RECT 558.450 381.450 565.050 382.500 ;
        RECT 558.450 380.700 560.250 381.450 ;
        RECT 563.250 380.700 565.050 381.450 ;
        RECT 570.150 381.300 574.050 383.400 ;
        RECT 554.550 379.500 555.750 380.400 ;
        RECT 567.450 379.800 569.250 380.400 ;
        RECT 554.550 378.300 562.050 379.500 ;
        RECT 560.250 377.700 562.050 378.300 ;
        RECT 562.950 378.900 569.250 379.800 ;
        RECT 546.150 376.500 547.050 377.400 ;
        RECT 562.950 376.800 563.850 378.900 ;
        RECT 567.450 378.600 569.250 378.900 ;
        RECT 570.150 378.600 572.850 380.400 ;
        RECT 570.150 377.700 571.050 378.600 ;
        RECT 555.450 376.500 563.850 376.800 ;
        RECT 546.150 375.900 563.850 376.500 ;
        RECT 565.950 376.800 571.050 377.700 ;
        RECT 571.950 376.800 574.050 377.700 ;
        RECT 577.650 377.400 579.450 389.400 ;
        RECT 587.400 383.400 589.200 390.000 ;
        RECT 590.400 383.400 592.200 389.400 ;
        RECT 546.150 375.300 557.250 375.900 ;
        RECT 546.150 360.600 547.050 375.300 ;
        RECT 555.450 375.000 557.250 375.300 ;
        RECT 547.950 367.950 550.050 370.050 ;
        RECT 556.950 368.400 559.050 370.050 ;
        RECT 548.100 366.150 549.900 367.950 ;
        RECT 551.100 367.200 559.050 368.400 ;
        RECT 551.100 366.600 552.900 367.200 ;
        RECT 549.000 365.400 549.900 366.150 ;
        RECT 554.100 365.400 555.900 366.000 ;
        RECT 549.000 364.200 555.900 365.400 ;
        RECT 565.950 364.200 566.850 376.800 ;
        RECT 571.950 375.600 576.150 376.800 ;
        RECT 575.250 373.800 577.050 375.600 ;
        RECT 578.250 370.050 579.450 377.400 ;
        RECT 587.100 370.050 588.900 371.850 ;
        RECT 590.400 370.050 591.600 383.400 ;
        RECT 602.400 377.400 604.200 390.000 ;
        RECT 606.900 377.400 610.200 389.400 ;
        RECT 612.900 377.400 614.700 390.000 ;
        RECT 626.400 383.400 628.200 390.000 ;
        RECT 629.400 383.400 631.200 389.400 ;
        RECT 632.400 383.400 634.200 390.000 ;
        RECT 574.950 369.750 579.450 370.050 ;
        RECT 573.150 367.950 579.450 369.750 ;
        RECT 586.950 367.950 589.050 370.050 ;
        RECT 589.950 367.950 592.050 370.050 ;
        RECT 602.100 369.900 603.900 371.700 ;
        RECT 608.100 369.900 609.300 377.400 ;
        RECT 614.100 369.900 615.900 371.700 ;
        RECT 554.850 363.000 566.850 364.200 ;
        RECT 554.850 361.200 555.900 363.000 ;
        RECT 565.050 362.400 566.850 363.000 ;
        RECT 546.150 354.600 547.950 360.600 ;
        RECT 550.950 358.500 553.050 360.600 ;
        RECT 554.550 359.400 556.350 361.200 ;
        RECT 578.250 360.600 579.450 367.950 ;
        RECT 557.850 359.550 559.650 360.300 ;
        RECT 571.950 359.700 574.050 360.600 ;
        RECT 557.850 358.500 562.800 359.550 ;
        RECT 552.000 357.600 553.050 358.500 ;
        RECT 561.750 357.600 562.800 358.500 ;
        RECT 570.300 358.500 574.050 359.700 ;
        RECT 570.300 357.600 571.350 358.500 ;
        RECT 549.150 354.000 550.950 357.600 ;
        RECT 552.000 356.700 555.750 357.600 ;
        RECT 553.950 354.600 555.750 356.700 ;
        RECT 558.450 354.000 560.250 357.600 ;
        RECT 561.750 354.600 563.550 357.600 ;
        RECT 565.350 354.000 567.150 357.600 ;
        RECT 569.550 354.600 571.350 357.600 ;
        RECT 574.350 354.000 576.150 357.600 ;
        RECT 577.650 354.600 579.450 360.600 ;
        RECT 590.400 357.600 591.600 367.950 ;
        RECT 601.950 367.800 604.050 369.900 ;
        RECT 604.950 367.800 607.050 369.900 ;
        RECT 607.950 367.800 610.050 369.900 ;
        RECT 610.950 367.800 613.050 369.900 ;
        RECT 613.950 367.800 616.050 369.900 ;
        RECT 625.950 367.800 628.050 369.900 ;
        RECT 605.100 366.000 606.900 367.800 ;
        RECT 607.950 365.400 609.000 367.800 ;
        RECT 611.100 366.000 612.900 367.800 ;
        RECT 626.100 366.000 627.900 367.800 ;
        RECT 608.100 363.300 609.300 365.400 ;
        RECT 629.400 363.300 630.300 383.400 ;
        RECT 635.400 377.400 637.200 389.400 ;
        RECT 649.800 388.500 657.600 389.400 ;
        RECT 649.800 377.400 651.600 388.500 ;
        RECT 632.100 369.900 633.900 371.700 ;
        RECT 635.700 369.900 636.600 377.400 ;
        RECT 652.800 376.500 654.600 387.600 ;
        RECT 655.800 378.600 657.600 388.500 ;
        RECT 658.800 379.500 660.600 390.000 ;
        RECT 661.800 378.600 663.600 389.400 ;
        RECT 655.800 377.700 663.600 378.600 ;
        RECT 666.150 377.400 667.950 389.400 ;
        RECT 669.150 383.400 670.950 390.000 ;
        RECT 674.550 383.400 676.350 389.400 ;
        RECT 679.350 383.400 681.150 390.000 ;
        RECT 674.550 382.500 675.750 383.400 ;
        RECT 682.350 382.500 684.150 389.400 ;
        RECT 685.950 383.400 687.750 390.000 ;
        RECT 690.150 383.400 691.950 389.400 ;
        RECT 694.650 386.400 696.450 390.000 ;
        RECT 670.950 380.400 675.750 382.500 ;
        RECT 678.450 381.450 685.050 382.500 ;
        RECT 678.450 380.700 680.250 381.450 ;
        RECT 683.250 380.700 685.050 381.450 ;
        RECT 690.150 381.300 694.050 383.400 ;
        RECT 674.550 379.500 675.750 380.400 ;
        RECT 687.450 379.800 689.250 380.400 ;
        RECT 674.550 378.300 682.050 379.500 ;
        RECT 680.250 377.700 682.050 378.300 ;
        RECT 682.950 378.900 689.250 379.800 ;
        RECT 666.150 376.500 667.050 377.400 ;
        RECT 682.950 376.800 683.850 378.900 ;
        RECT 687.450 378.600 689.250 378.900 ;
        RECT 690.150 378.600 692.850 380.400 ;
        RECT 690.150 377.700 691.050 378.600 ;
        RECT 675.450 376.500 683.850 376.800 ;
        RECT 652.800 375.600 657.900 376.500 ;
        RECT 653.100 369.900 654.900 371.700 ;
        RECT 657.000 369.900 657.900 375.600 ;
        RECT 666.150 375.900 683.850 376.500 ;
        RECT 685.950 376.800 691.050 377.700 ;
        RECT 691.950 376.800 694.050 377.700 ;
        RECT 697.650 377.400 699.450 389.400 ;
        RECT 666.150 375.300 677.250 375.900 ;
        RECT 659.100 369.900 660.900 371.700 ;
        RECT 631.950 367.800 634.050 369.900 ;
        RECT 634.950 367.800 637.050 369.900 ;
        RECT 649.950 367.800 652.050 369.900 ;
        RECT 652.950 367.800 655.050 369.900 ;
        RECT 655.950 367.800 658.050 369.900 ;
        RECT 658.950 367.800 661.050 369.900 ;
        RECT 661.950 367.800 664.050 369.900 ;
        RECT 608.100 362.100 612.600 363.300 ;
        RECT 602.400 360.000 610.200 360.900 ;
        RECT 611.700 360.600 612.600 362.100 ;
        RECT 626.400 362.400 633.900 363.300 ;
        RECT 587.400 354.000 589.200 357.600 ;
        RECT 590.400 354.600 592.200 357.600 ;
        RECT 602.400 354.600 604.200 360.000 ;
        RECT 605.400 354.000 607.200 359.100 ;
        RECT 608.400 355.500 610.200 360.000 ;
        RECT 611.400 356.400 613.200 360.600 ;
        RECT 614.400 355.500 616.200 360.600 ;
        RECT 608.400 354.600 616.200 355.500 ;
        RECT 626.400 354.600 628.200 362.400 ;
        RECT 632.100 361.500 633.900 362.400 ;
        RECT 635.700 360.600 636.600 367.800 ;
        RECT 650.100 366.000 651.900 367.800 ;
        RECT 657.000 360.600 658.050 367.800 ;
        RECT 662.100 366.000 663.900 367.800 ;
        RECT 666.150 360.600 667.050 375.300 ;
        RECT 675.450 375.000 677.250 375.300 ;
        RECT 667.950 367.950 670.050 370.050 ;
        RECT 676.950 368.400 679.050 370.050 ;
        RECT 668.100 366.150 669.900 367.950 ;
        RECT 671.100 367.200 679.050 368.400 ;
        RECT 671.100 366.600 672.900 367.200 ;
        RECT 669.000 365.400 669.900 366.150 ;
        RECT 674.100 365.400 675.900 366.000 ;
        RECT 669.000 364.200 675.900 365.400 ;
        RECT 685.950 364.200 686.850 376.800 ;
        RECT 691.950 375.600 696.150 376.800 ;
        RECT 695.250 373.800 697.050 375.600 ;
        RECT 698.250 370.050 699.450 377.400 ;
        RECT 694.950 369.750 699.450 370.050 ;
        RECT 693.150 367.950 699.450 369.750 ;
        RECT 674.850 363.000 686.850 364.200 ;
        RECT 674.850 361.200 675.900 363.000 ;
        RECT 685.050 362.400 686.850 363.000 ;
        RECT 630.900 354.000 632.700 360.600 ;
        RECT 633.900 358.800 636.600 360.600 ;
        RECT 633.900 354.600 635.700 358.800 ;
        RECT 652.500 354.000 654.300 360.600 ;
        RECT 657.000 354.600 658.800 360.600 ;
        RECT 661.500 354.000 663.300 360.600 ;
        RECT 666.150 354.600 667.950 360.600 ;
        RECT 670.950 358.500 673.050 360.600 ;
        RECT 674.550 359.400 676.350 361.200 ;
        RECT 698.250 360.600 699.450 367.950 ;
        RECT 677.850 359.550 679.650 360.300 ;
        RECT 691.950 359.700 694.050 360.600 ;
        RECT 677.850 358.500 682.800 359.550 ;
        RECT 672.000 357.600 673.050 358.500 ;
        RECT 681.750 357.600 682.800 358.500 ;
        RECT 690.300 358.500 694.050 359.700 ;
        RECT 690.300 357.600 691.350 358.500 ;
        RECT 669.150 354.000 670.950 357.600 ;
        RECT 672.000 356.700 675.750 357.600 ;
        RECT 673.950 354.600 675.750 356.700 ;
        RECT 678.450 354.000 680.250 357.600 ;
        RECT 681.750 354.600 683.550 357.600 ;
        RECT 685.350 354.000 687.150 357.600 ;
        RECT 689.550 354.600 691.350 357.600 ;
        RECT 694.350 354.000 696.150 357.600 ;
        RECT 697.650 354.600 699.450 360.600 ;
        RECT 702.150 377.400 703.950 389.400 ;
        RECT 705.150 383.400 706.950 390.000 ;
        RECT 710.550 383.400 712.350 389.400 ;
        RECT 715.350 383.400 717.150 390.000 ;
        RECT 710.550 382.500 711.750 383.400 ;
        RECT 718.350 382.500 720.150 389.400 ;
        RECT 721.950 383.400 723.750 390.000 ;
        RECT 726.150 383.400 727.950 389.400 ;
        RECT 730.650 386.400 732.450 390.000 ;
        RECT 706.950 380.400 711.750 382.500 ;
        RECT 714.450 381.450 721.050 382.500 ;
        RECT 714.450 380.700 716.250 381.450 ;
        RECT 719.250 380.700 721.050 381.450 ;
        RECT 726.150 381.300 730.050 383.400 ;
        RECT 710.550 379.500 711.750 380.400 ;
        RECT 723.450 379.800 725.250 380.400 ;
        RECT 710.550 378.300 718.050 379.500 ;
        RECT 716.250 377.700 718.050 378.300 ;
        RECT 718.950 378.900 725.250 379.800 ;
        RECT 702.150 376.500 703.050 377.400 ;
        RECT 718.950 376.800 719.850 378.900 ;
        RECT 723.450 378.600 725.250 378.900 ;
        RECT 726.150 378.600 728.850 380.400 ;
        RECT 726.150 377.700 727.050 378.600 ;
        RECT 711.450 376.500 719.850 376.800 ;
        RECT 702.150 375.900 719.850 376.500 ;
        RECT 721.950 376.800 727.050 377.700 ;
        RECT 727.950 376.800 730.050 377.700 ;
        RECT 733.650 377.400 735.450 389.400 ;
        RECT 745.800 383.400 747.600 389.400 ;
        RECT 748.800 383.400 750.600 390.000 ;
        RECT 702.150 375.300 713.250 375.900 ;
        RECT 702.150 360.600 703.050 375.300 ;
        RECT 711.450 375.000 713.250 375.300 ;
        RECT 703.950 367.950 706.050 370.050 ;
        RECT 712.950 368.400 715.050 370.050 ;
        RECT 704.100 366.150 705.900 367.950 ;
        RECT 707.100 367.200 715.050 368.400 ;
        RECT 707.100 366.600 708.900 367.200 ;
        RECT 705.000 365.400 705.900 366.150 ;
        RECT 710.100 365.400 711.900 366.000 ;
        RECT 705.000 364.200 711.900 365.400 ;
        RECT 721.950 364.200 722.850 376.800 ;
        RECT 727.950 375.600 732.150 376.800 ;
        RECT 731.250 373.800 733.050 375.600 ;
        RECT 734.250 370.050 735.450 377.400 ;
        RECT 746.400 370.050 747.600 383.400 ;
        RECT 758.700 377.400 760.500 390.000 ;
        RECT 763.800 383.400 765.600 389.400 ;
        RECT 766.800 383.400 768.600 390.000 ;
        RECT 749.100 370.050 750.900 371.850 ;
        RECT 758.100 370.050 759.900 371.850 ;
        RECT 763.950 370.050 765.150 383.400 ;
        RECT 774.150 377.400 775.950 389.400 ;
        RECT 777.150 383.400 778.950 390.000 ;
        RECT 782.550 383.400 784.350 389.400 ;
        RECT 787.350 383.400 789.150 390.000 ;
        RECT 782.550 382.500 783.750 383.400 ;
        RECT 790.350 382.500 792.150 389.400 ;
        RECT 793.950 383.400 795.750 390.000 ;
        RECT 798.150 383.400 799.950 389.400 ;
        RECT 802.650 386.400 804.450 390.000 ;
        RECT 778.950 380.400 783.750 382.500 ;
        RECT 786.450 381.450 793.050 382.500 ;
        RECT 786.450 380.700 788.250 381.450 ;
        RECT 791.250 380.700 793.050 381.450 ;
        RECT 798.150 381.300 802.050 383.400 ;
        RECT 782.550 379.500 783.750 380.400 ;
        RECT 795.450 379.800 797.250 380.400 ;
        RECT 782.550 378.300 790.050 379.500 ;
        RECT 788.250 377.700 790.050 378.300 ;
        RECT 790.950 378.900 797.250 379.800 ;
        RECT 774.150 376.500 775.050 377.400 ;
        RECT 790.950 376.800 791.850 378.900 ;
        RECT 795.450 378.600 797.250 378.900 ;
        RECT 798.150 378.600 800.850 380.400 ;
        RECT 798.150 377.700 799.050 378.600 ;
        RECT 783.450 376.500 791.850 376.800 ;
        RECT 774.150 375.900 791.850 376.500 ;
        RECT 793.950 376.800 799.050 377.700 ;
        RECT 799.950 376.800 802.050 377.700 ;
        RECT 805.650 377.400 807.450 389.400 ;
        RECT 817.800 383.400 819.600 390.000 ;
        RECT 820.800 383.400 822.600 389.400 ;
        RECT 823.800 383.400 825.600 390.000 ;
        RECT 833.400 383.400 835.200 390.000 ;
        RECT 836.400 383.400 838.200 389.400 ;
        RECT 839.400 383.400 841.200 390.000 ;
        RECT 774.150 375.300 785.250 375.900 ;
        RECT 730.950 369.750 735.450 370.050 ;
        RECT 729.150 367.950 735.450 369.750 ;
        RECT 745.950 367.950 748.050 370.050 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 763.950 367.950 766.050 370.050 ;
        RECT 766.950 367.950 769.050 370.050 ;
        RECT 710.850 363.000 722.850 364.200 ;
        RECT 710.850 361.200 711.900 363.000 ;
        RECT 721.050 362.400 722.850 363.000 ;
        RECT 702.150 354.600 703.950 360.600 ;
        RECT 706.950 358.500 709.050 360.600 ;
        RECT 710.550 359.400 712.350 361.200 ;
        RECT 734.250 360.600 735.450 367.950 ;
        RECT 713.850 359.550 715.650 360.300 ;
        RECT 727.950 359.700 730.050 360.600 ;
        RECT 713.850 358.500 718.800 359.550 ;
        RECT 708.000 357.600 709.050 358.500 ;
        RECT 717.750 357.600 718.800 358.500 ;
        RECT 726.300 358.500 730.050 359.700 ;
        RECT 726.300 357.600 727.350 358.500 ;
        RECT 705.150 354.000 706.950 357.600 ;
        RECT 708.000 356.700 711.750 357.600 ;
        RECT 709.950 354.600 711.750 356.700 ;
        RECT 714.450 354.000 716.250 357.600 ;
        RECT 717.750 354.600 719.550 357.600 ;
        RECT 721.350 354.000 723.150 357.600 ;
        RECT 725.550 354.600 727.350 357.600 ;
        RECT 730.350 354.000 732.150 357.600 ;
        RECT 733.650 354.600 735.450 360.600 ;
        RECT 746.400 357.600 747.600 367.950 ;
        RECT 761.100 366.150 762.900 367.950 ;
        RECT 764.850 363.750 766.050 367.950 ;
        RECT 767.100 366.150 768.900 367.950 ;
        RECT 764.850 362.700 768.600 363.750 ;
        RECT 758.400 359.700 766.200 361.050 ;
        RECT 745.800 354.600 747.600 357.600 ;
        RECT 748.800 354.000 750.600 357.600 ;
        RECT 758.400 354.600 760.200 359.700 ;
        RECT 761.400 354.000 763.200 358.800 ;
        RECT 764.400 354.600 766.200 359.700 ;
        RECT 767.400 360.600 768.600 362.700 ;
        RECT 774.150 360.600 775.050 375.300 ;
        RECT 783.450 375.000 785.250 375.300 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 784.950 368.400 787.050 370.050 ;
        RECT 776.100 366.150 777.900 367.950 ;
        RECT 779.100 367.200 787.050 368.400 ;
        RECT 779.100 366.600 780.900 367.200 ;
        RECT 777.000 365.400 777.900 366.150 ;
        RECT 782.100 365.400 783.900 366.000 ;
        RECT 777.000 364.200 783.900 365.400 ;
        RECT 793.950 364.200 794.850 376.800 ;
        RECT 799.950 375.600 804.150 376.800 ;
        RECT 803.250 373.800 805.050 375.600 ;
        RECT 806.250 370.050 807.450 377.400 ;
        RECT 802.950 369.750 807.450 370.050 ;
        RECT 821.400 369.900 822.600 383.400 ;
        RECT 836.400 369.900 837.600 383.400 ;
        RECT 801.150 367.950 807.450 369.750 ;
        RECT 782.850 363.000 794.850 364.200 ;
        RECT 782.850 361.200 783.900 363.000 ;
        RECT 793.050 362.400 794.850 363.000 ;
        RECT 767.400 354.600 769.200 360.600 ;
        RECT 774.150 354.600 775.950 360.600 ;
        RECT 778.950 358.500 781.050 360.600 ;
        RECT 782.550 359.400 784.350 361.200 ;
        RECT 806.250 360.600 807.450 367.950 ;
        RECT 817.950 367.800 820.050 369.900 ;
        RECT 820.950 367.800 823.050 369.900 ;
        RECT 823.950 367.800 826.050 369.900 ;
        RECT 832.950 367.800 835.050 369.900 ;
        RECT 835.950 367.800 838.050 369.900 ;
        RECT 838.950 367.800 841.050 369.900 ;
        RECT 818.100 366.000 819.900 367.800 ;
        RECT 821.400 362.700 822.600 367.800 ;
        RECT 824.100 366.000 825.900 367.800 ;
        RECT 833.100 366.000 834.900 367.800 ;
        RECT 785.850 359.550 787.650 360.300 ;
        RECT 799.950 359.700 802.050 360.600 ;
        RECT 785.850 358.500 790.800 359.550 ;
        RECT 780.000 357.600 781.050 358.500 ;
        RECT 789.750 357.600 790.800 358.500 ;
        RECT 798.300 358.500 802.050 359.700 ;
        RECT 798.300 357.600 799.350 358.500 ;
        RECT 777.150 354.000 778.950 357.600 ;
        RECT 780.000 356.700 783.750 357.600 ;
        RECT 781.950 354.600 783.750 356.700 ;
        RECT 786.450 354.000 788.250 357.600 ;
        RECT 789.750 354.600 791.550 357.600 ;
        RECT 793.350 354.000 795.150 357.600 ;
        RECT 797.550 354.600 799.350 357.600 ;
        RECT 802.350 354.000 804.150 357.600 ;
        RECT 805.650 354.600 807.450 360.600 ;
        RECT 818.400 361.800 822.600 362.700 ;
        RECT 836.400 362.700 837.600 367.800 ;
        RECT 839.100 366.000 840.900 367.800 ;
        RECT 836.400 361.800 840.600 362.700 ;
        RECT 818.400 354.600 820.200 361.800 ;
        RECT 823.500 354.000 825.300 360.600 ;
        RECT 833.700 354.000 835.500 360.600 ;
        RECT 838.800 354.600 840.600 361.800 ;
        RECT 10.800 347.400 12.600 350.400 ;
        RECT 13.800 347.400 15.600 351.000 ;
        RECT 11.400 337.050 12.600 347.400 ;
        RECT 28.200 342.000 30.000 350.400 ;
        RECT 26.700 340.800 30.000 342.000 ;
        RECT 34.800 341.400 36.600 351.000 ;
        RECT 45.000 344.400 46.800 351.000 ;
        RECT 49.500 345.600 51.300 350.400 ;
        RECT 52.500 347.400 54.300 351.000 ;
        RECT 49.500 344.400 54.600 345.600 ;
        RECT 67.800 344.400 69.600 350.400 ;
        RECT 26.700 337.200 27.600 340.800 ;
        RECT 29.100 337.200 30.900 339.000 ;
        RECT 35.100 337.200 36.900 339.000 ;
        RECT 44.100 337.200 45.900 339.000 ;
        RECT 50.100 337.200 51.900 339.000 ;
        RECT 53.700 337.200 54.600 344.400 ;
        RECT 68.400 342.300 69.600 344.400 ;
        RECT 70.800 345.300 72.600 350.400 ;
        RECT 73.800 346.200 75.600 351.000 ;
        RECT 76.800 345.300 78.600 350.400 ;
        RECT 88.800 347.400 90.600 350.400 ;
        RECT 91.800 347.400 93.600 351.000 ;
        RECT 103.800 349.500 111.600 350.400 ;
        RECT 70.800 343.950 78.600 345.300 ;
        RECT 68.400 341.250 72.150 342.300 ;
        RECT 10.950 334.950 13.050 337.050 ;
        RECT 13.950 334.950 16.050 337.050 ;
        RECT 25.950 335.100 28.050 337.200 ;
        RECT 28.950 335.100 31.050 337.200 ;
        RECT 31.950 335.100 34.050 337.200 ;
        RECT 34.950 335.100 37.050 337.200 ;
        RECT 43.950 335.100 46.050 337.200 ;
        RECT 46.950 335.100 49.050 337.200 ;
        RECT 49.950 335.100 52.050 337.200 ;
        RECT 52.950 335.100 55.050 337.200 ;
        RECT 68.100 337.050 69.900 338.850 ;
        RECT 70.950 337.050 72.150 341.250 ;
        RECT 74.100 337.050 75.900 338.850 ;
        RECT 89.400 337.050 90.600 347.400 ;
        RECT 103.800 344.400 105.600 349.500 ;
        RECT 106.800 344.400 108.600 348.600 ;
        RECT 109.800 345.000 111.600 349.500 ;
        RECT 112.800 345.900 114.600 351.000 ;
        RECT 115.800 345.000 117.600 350.400 ;
        RECT 107.400 342.900 108.300 344.400 ;
        RECT 109.800 344.100 117.600 345.000 ;
        RECT 125.700 344.400 127.500 351.000 ;
        RECT 130.800 343.200 132.600 350.400 ;
        RECT 145.800 347.400 147.600 350.400 ;
        RECT 148.800 347.400 150.600 351.000 ;
        RECT 107.400 341.700 111.900 342.900 ;
        RECT 110.700 339.600 111.900 341.700 ;
        RECT 128.400 342.300 132.600 343.200 ;
        RECT 107.100 337.200 108.900 339.000 ;
        RECT 111.000 337.200 112.050 339.600 ;
        RECT 113.100 337.200 114.900 339.000 ;
        RECT 125.100 337.200 126.900 339.000 ;
        RECT 128.400 337.200 129.600 342.300 ;
        RECT 131.100 337.200 132.900 339.000 ;
        RECT 11.400 321.600 12.600 334.950 ;
        RECT 14.100 333.150 15.900 334.950 ;
        RECT 26.700 322.800 27.600 335.100 ;
        RECT 32.100 333.300 33.900 335.100 ;
        RECT 47.100 333.300 48.900 335.100 ;
        RECT 34.950 330.450 37.050 331.050 ;
        RECT 49.950 330.450 52.050 331.050 ;
        RECT 34.950 329.550 52.050 330.450 ;
        RECT 34.950 328.950 37.050 329.550 ;
        RECT 49.950 328.950 52.050 329.550 ;
        RECT 53.700 327.600 54.600 335.100 ;
        RECT 67.950 334.950 70.050 337.050 ;
        RECT 70.950 334.950 73.050 337.050 ;
        RECT 73.950 334.950 76.050 337.050 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 88.950 334.950 91.050 337.050 ;
        RECT 91.950 334.950 94.050 337.050 ;
        RECT 103.950 335.100 106.050 337.200 ;
        RECT 106.950 335.100 109.050 337.200 ;
        RECT 109.950 335.100 112.050 337.200 ;
        RECT 112.950 335.100 115.050 337.200 ;
        RECT 115.950 335.100 118.050 337.200 ;
        RECT 124.950 335.100 127.050 337.200 ;
        RECT 127.950 335.100 130.050 337.200 ;
        RECT 130.950 335.100 133.050 337.200 ;
        RECT 146.400 337.050 147.600 347.400 ;
        RECT 153.150 344.400 154.950 350.400 ;
        RECT 156.150 347.400 157.950 351.000 ;
        RECT 160.950 348.300 162.750 350.400 ;
        RECT 159.000 347.400 162.750 348.300 ;
        RECT 165.450 347.400 167.250 351.000 ;
        RECT 168.750 347.400 170.550 350.400 ;
        RECT 172.350 347.400 174.150 351.000 ;
        RECT 176.550 347.400 178.350 350.400 ;
        RECT 181.350 347.400 183.150 351.000 ;
        RECT 159.000 346.500 160.050 347.400 ;
        RECT 168.750 346.500 169.800 347.400 ;
        RECT 157.950 344.400 160.050 346.500 ;
        RECT 44.400 326.700 52.200 327.600 ;
        RECT 26.700 321.900 33.300 322.800 ;
        RECT 26.700 321.600 27.600 321.900 ;
        RECT 10.800 315.600 12.600 321.600 ;
        RECT 13.800 315.000 15.600 321.600 ;
        RECT 25.800 315.600 27.600 321.600 ;
        RECT 31.800 321.600 33.300 321.900 ;
        RECT 28.800 315.000 30.600 321.000 ;
        RECT 31.800 315.600 33.600 321.600 ;
        RECT 34.800 315.000 36.600 321.600 ;
        RECT 44.400 315.600 46.200 326.700 ;
        RECT 47.400 315.000 49.200 325.800 ;
        RECT 50.400 315.600 52.200 326.700 ;
        RECT 53.400 315.600 55.200 327.600 ;
        RECT 71.850 321.600 73.050 334.950 ;
        RECT 77.100 333.150 78.900 334.950 ;
        RECT 68.400 315.000 70.200 321.600 ;
        RECT 71.400 315.600 73.200 321.600 ;
        RECT 76.500 315.000 78.300 327.600 ;
        RECT 89.400 321.600 90.600 334.950 ;
        RECT 92.100 333.150 93.900 334.950 ;
        RECT 104.100 333.300 105.900 335.100 ;
        RECT 110.700 327.600 111.900 335.100 ;
        RECT 116.100 333.300 117.900 335.100 ;
        RECT 88.800 315.600 90.600 321.600 ;
        RECT 91.800 315.000 93.600 321.600 ;
        RECT 105.300 315.000 107.100 327.600 ;
        RECT 109.800 315.600 113.100 327.600 ;
        RECT 115.800 315.000 117.600 327.600 ;
        RECT 128.400 321.600 129.600 335.100 ;
        RECT 145.950 334.950 148.050 337.050 ;
        RECT 148.950 334.950 151.050 337.050 ;
        RECT 146.400 321.600 147.600 334.950 ;
        RECT 149.100 333.150 150.900 334.950 ;
        RECT 153.150 329.700 154.050 344.400 ;
        RECT 161.550 343.800 163.350 345.600 ;
        RECT 164.850 345.450 169.800 346.500 ;
        RECT 177.300 346.500 178.350 347.400 ;
        RECT 164.850 344.700 166.650 345.450 ;
        RECT 177.300 345.300 181.050 346.500 ;
        RECT 178.950 344.400 181.050 345.300 ;
        RECT 184.650 344.400 186.450 350.400 ;
        RECT 161.850 342.000 162.900 343.800 ;
        RECT 172.050 342.000 173.850 342.600 ;
        RECT 161.850 340.800 173.850 342.000 ;
        RECT 156.000 339.600 162.900 340.800 ;
        RECT 156.000 338.850 156.900 339.600 ;
        RECT 161.100 339.000 162.900 339.600 ;
        RECT 155.100 337.050 156.900 338.850 ;
        RECT 158.100 337.800 159.900 338.400 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 158.100 336.600 166.050 337.800 ;
        RECT 163.950 334.950 166.050 336.600 ;
        RECT 162.450 329.700 164.250 330.000 ;
        RECT 153.150 329.100 164.250 329.700 ;
        RECT 153.150 328.500 170.850 329.100 ;
        RECT 153.150 327.600 154.050 328.500 ;
        RECT 162.450 328.200 170.850 328.500 ;
        RECT 125.400 315.000 127.200 321.600 ;
        RECT 128.400 315.600 130.200 321.600 ;
        RECT 131.400 315.000 133.200 321.600 ;
        RECT 145.800 315.600 147.600 321.600 ;
        RECT 148.800 315.000 150.600 321.600 ;
        RECT 153.150 315.600 154.950 327.600 ;
        RECT 167.250 326.700 169.050 327.300 ;
        RECT 161.550 325.500 169.050 326.700 ;
        RECT 169.950 326.100 170.850 328.200 ;
        RECT 172.950 328.200 173.850 340.800 ;
        RECT 185.250 337.050 186.450 344.400 ;
        RECT 194.400 345.300 196.200 350.400 ;
        RECT 197.400 346.200 199.200 351.000 ;
        RECT 200.400 345.300 202.200 350.400 ;
        RECT 194.400 343.950 202.200 345.300 ;
        RECT 203.400 344.400 205.200 350.400 ;
        RECT 203.400 342.300 204.600 344.400 ;
        RECT 218.400 343.200 220.200 350.400 ;
        RECT 223.500 344.400 225.300 351.000 ;
        RECT 233.400 345.300 235.200 350.400 ;
        RECT 236.400 346.200 238.200 351.000 ;
        RECT 239.400 345.300 241.200 350.400 ;
        RECT 233.400 343.950 241.200 345.300 ;
        RECT 242.400 344.400 244.200 350.400 ;
        RECT 254.700 344.400 256.500 351.000 ;
        RECT 218.400 342.300 222.600 343.200 ;
        RECT 242.400 342.300 243.600 344.400 ;
        RECT 259.800 343.200 261.600 350.400 ;
        RECT 272.400 347.400 274.200 351.000 ;
        RECT 275.400 347.400 277.200 350.400 ;
        RECT 287.400 347.400 289.200 351.000 ;
        RECT 290.400 347.400 292.200 350.400 ;
        RECT 200.850 341.250 204.600 342.300 ;
        RECT 197.100 337.050 198.900 338.850 ;
        RECT 200.850 337.050 202.050 341.250 ;
        RECT 203.100 337.050 204.900 338.850 ;
        RECT 218.100 337.200 219.900 339.000 ;
        RECT 221.400 337.200 222.600 342.300 ;
        RECT 239.850 341.250 243.600 342.300 ;
        RECT 257.400 342.300 261.600 343.200 ;
        RECT 224.100 337.200 225.900 339.000 ;
        RECT 180.150 335.250 186.450 337.050 ;
        RECT 181.950 334.950 186.450 335.250 ;
        RECT 193.950 334.950 196.050 337.050 ;
        RECT 196.950 334.950 199.050 337.050 ;
        RECT 199.950 334.950 202.050 337.050 ;
        RECT 202.950 334.950 205.050 337.050 ;
        RECT 217.950 335.100 220.050 337.200 ;
        RECT 220.950 335.100 223.050 337.200 ;
        RECT 223.950 335.100 226.050 337.200 ;
        RECT 236.100 337.050 237.900 338.850 ;
        RECT 239.850 337.050 241.050 341.250 ;
        RECT 242.100 337.050 243.900 338.850 ;
        RECT 254.100 337.200 255.900 339.000 ;
        RECT 257.400 337.200 258.600 342.300 ;
        RECT 260.100 337.200 261.900 339.000 ;
        RECT 182.250 329.400 184.050 331.200 ;
        RECT 178.950 328.200 183.150 329.400 ;
        RECT 172.950 327.300 178.050 328.200 ;
        RECT 178.950 327.300 181.050 328.200 ;
        RECT 185.250 327.600 186.450 334.950 ;
        RECT 194.100 333.150 195.900 334.950 ;
        RECT 177.150 326.400 178.050 327.300 ;
        RECT 174.450 326.100 176.250 326.400 ;
        RECT 161.550 324.600 162.750 325.500 ;
        RECT 169.950 325.200 176.250 326.100 ;
        RECT 174.450 324.600 176.250 325.200 ;
        RECT 177.150 324.600 179.850 326.400 ;
        RECT 157.950 322.500 162.750 324.600 ;
        RECT 165.450 323.550 167.250 324.300 ;
        RECT 170.250 323.550 172.050 324.300 ;
        RECT 165.450 322.500 172.050 323.550 ;
        RECT 161.550 321.600 162.750 322.500 ;
        RECT 156.150 315.000 157.950 321.600 ;
        RECT 161.550 315.600 163.350 321.600 ;
        RECT 166.350 315.000 168.150 321.600 ;
        RECT 169.350 315.600 171.150 322.500 ;
        RECT 177.150 321.600 181.050 323.700 ;
        RECT 172.950 315.000 174.750 321.600 ;
        RECT 177.150 315.600 178.950 321.600 ;
        RECT 181.650 315.000 183.450 318.600 ;
        RECT 184.650 315.600 186.450 327.600 ;
        RECT 194.700 315.000 196.500 327.600 ;
        RECT 199.950 321.600 201.150 334.950 ;
        RECT 221.400 321.600 222.600 335.100 ;
        RECT 232.950 334.950 235.050 337.050 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 238.950 334.950 241.050 337.050 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 253.950 335.100 256.050 337.200 ;
        RECT 256.950 335.100 259.050 337.200 ;
        RECT 259.950 335.100 262.050 337.200 ;
        RECT 275.400 337.050 276.600 347.400 ;
        RECT 277.950 339.450 282.000 340.050 ;
        RECT 277.950 337.950 282.450 339.450 ;
        RECT 233.100 333.150 234.900 334.950 ;
        RECT 199.800 315.600 201.600 321.600 ;
        RECT 202.800 315.000 204.600 321.600 ;
        RECT 217.800 315.000 219.600 321.600 ;
        RECT 220.800 315.600 222.600 321.600 ;
        RECT 223.800 315.000 225.600 321.600 ;
        RECT 233.700 315.000 235.500 327.600 ;
        RECT 238.950 321.600 240.150 334.950 ;
        RECT 257.400 321.600 258.600 335.100 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 272.100 333.150 273.900 334.950 ;
        RECT 275.400 321.600 276.600 334.950 ;
        RECT 281.550 334.050 282.450 337.950 ;
        RECT 290.400 337.050 291.600 347.400 ;
        RECT 305.400 343.200 307.200 350.400 ;
        RECT 310.500 344.400 312.300 351.000 ;
        RECT 320.700 344.400 322.500 351.000 ;
        RECT 325.800 343.200 327.600 350.400 ;
        RECT 338.400 347.400 340.200 351.000 ;
        RECT 341.400 347.400 343.200 350.400 ;
        RECT 355.800 347.400 357.600 351.000 ;
        RECT 358.800 347.400 360.600 350.400 ;
        RECT 361.800 347.400 363.600 351.000 ;
        RECT 305.400 342.300 309.600 343.200 ;
        RECT 301.950 339.450 304.050 340.050 ;
        RECT 296.550 338.550 304.050 339.450 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 289.950 334.950 292.050 337.050 ;
        RECT 277.950 332.550 282.450 334.050 ;
        RECT 287.100 333.150 288.900 334.950 ;
        RECT 277.950 331.950 282.000 332.550 ;
        RECT 290.400 321.600 291.600 334.950 ;
        RECT 296.550 334.050 297.450 338.550 ;
        RECT 301.950 337.950 304.050 338.550 ;
        RECT 305.100 337.200 306.900 339.000 ;
        RECT 308.400 337.200 309.600 342.300 ;
        RECT 323.400 342.300 327.600 343.200 ;
        RECT 311.100 337.200 312.900 339.000 ;
        RECT 320.100 337.200 321.900 339.000 ;
        RECT 323.400 337.200 324.600 342.300 ;
        RECT 326.100 337.200 327.900 339.000 ;
        RECT 304.950 335.100 307.050 337.200 ;
        RECT 307.950 335.100 310.050 337.200 ;
        RECT 310.950 335.100 313.050 337.200 ;
        RECT 319.950 335.100 322.050 337.200 ;
        RECT 322.950 335.100 325.050 337.200 ;
        RECT 325.950 335.100 328.050 337.200 ;
        RECT 341.400 337.050 342.600 347.400 ;
        RECT 359.400 337.050 360.300 347.400 ;
        RECT 371.400 345.300 373.200 350.400 ;
        RECT 374.400 346.200 376.200 351.000 ;
        RECT 377.400 345.300 379.200 350.400 ;
        RECT 371.400 343.950 379.200 345.300 ;
        RECT 380.400 344.400 382.200 350.400 ;
        RECT 392.400 347.400 394.200 350.400 ;
        RECT 395.400 347.400 397.200 351.000 ;
        RECT 380.400 342.300 381.600 344.400 ;
        RECT 392.400 343.500 393.600 347.400 ;
        RECT 398.400 344.400 400.200 350.400 ;
        RECT 412.800 344.400 414.600 350.400 ;
        RECT 392.400 342.600 398.100 343.500 ;
        RECT 377.850 341.250 381.600 342.300 ;
        RECT 396.150 341.700 398.100 342.600 ;
        RECT 374.100 337.050 375.900 338.850 ;
        RECT 377.850 337.050 379.050 341.250 ;
        RECT 380.100 337.050 381.900 338.850 ;
        RECT 292.950 332.550 297.450 334.050 ;
        RECT 292.950 331.950 297.000 332.550 ;
        RECT 308.400 321.600 309.600 335.100 ;
        RECT 323.400 321.600 324.600 335.100 ;
        RECT 337.950 334.950 340.050 337.050 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 355.950 334.950 358.050 337.050 ;
        RECT 358.950 334.950 361.050 337.050 ;
        RECT 361.950 334.950 364.050 337.050 ;
        RECT 370.950 334.950 373.050 337.050 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 379.950 334.950 382.050 337.050 ;
        RECT 391.950 334.950 394.050 337.050 ;
        RECT 338.100 333.150 339.900 334.950 ;
        RECT 341.400 321.600 342.600 334.950 ;
        RECT 356.100 333.150 357.900 334.950 ;
        RECT 359.400 327.600 360.300 334.950 ;
        RECT 362.100 333.150 363.900 334.950 ;
        RECT 371.100 333.150 372.900 334.950 ;
        RECT 356.700 326.400 360.300 327.600 ;
        RECT 238.800 315.600 240.600 321.600 ;
        RECT 241.800 315.000 243.600 321.600 ;
        RECT 254.400 315.000 256.200 321.600 ;
        RECT 257.400 315.600 259.200 321.600 ;
        RECT 260.400 315.000 262.200 321.600 ;
        RECT 272.400 315.000 274.200 321.600 ;
        RECT 275.400 315.600 277.200 321.600 ;
        RECT 287.400 315.000 289.200 321.600 ;
        RECT 290.400 315.600 292.200 321.600 ;
        RECT 304.800 315.000 306.600 321.600 ;
        RECT 307.800 315.600 309.600 321.600 ;
        RECT 310.800 315.000 312.600 321.600 ;
        RECT 320.400 315.000 322.200 321.600 ;
        RECT 323.400 315.600 325.200 321.600 ;
        RECT 326.400 315.000 328.200 321.600 ;
        RECT 338.400 315.000 340.200 321.600 ;
        RECT 341.400 315.600 343.200 321.600 ;
        RECT 356.700 315.600 358.500 326.400 ;
        RECT 361.800 315.000 363.600 327.600 ;
        RECT 371.700 315.000 373.500 327.600 ;
        RECT 376.950 321.600 378.150 334.950 ;
        RECT 392.100 333.150 393.900 334.950 ;
        RECT 396.150 330.300 397.050 341.700 ;
        RECT 399.000 337.050 400.200 344.400 ;
        RECT 413.400 342.300 414.600 344.400 ;
        RECT 415.800 345.300 417.600 350.400 ;
        RECT 418.800 346.200 420.600 351.000 ;
        RECT 421.800 345.300 423.600 350.400 ;
        RECT 433.800 347.400 435.600 350.400 ;
        RECT 436.800 347.400 438.600 351.000 ;
        RECT 415.800 343.950 423.600 345.300 ;
        RECT 413.400 341.250 417.150 342.300 ;
        RECT 413.100 337.050 414.900 338.850 ;
        RECT 415.950 337.050 417.150 341.250 ;
        RECT 419.100 337.050 420.900 338.850 ;
        RECT 434.400 337.050 435.600 347.400 ;
        RECT 440.550 344.400 442.350 350.400 ;
        RECT 443.850 347.400 445.650 351.000 ;
        RECT 448.650 347.400 450.450 350.400 ;
        RECT 452.850 347.400 454.650 351.000 ;
        RECT 456.450 347.400 458.250 350.400 ;
        RECT 459.750 347.400 461.550 351.000 ;
        RECT 464.250 348.300 466.050 350.400 ;
        RECT 464.250 347.400 468.000 348.300 ;
        RECT 469.050 347.400 470.850 351.000 ;
        RECT 448.650 346.500 449.700 347.400 ;
        RECT 445.950 345.300 449.700 346.500 ;
        RECT 457.200 346.500 458.250 347.400 ;
        RECT 466.950 346.500 468.000 347.400 ;
        RECT 457.200 345.450 462.150 346.500 ;
        RECT 445.950 344.400 448.050 345.300 ;
        RECT 460.350 344.700 462.150 345.450 ;
        RECT 440.550 337.050 441.750 344.400 ;
        RECT 463.650 343.800 465.450 345.600 ;
        RECT 466.950 344.400 469.050 346.500 ;
        RECT 472.050 344.400 473.850 350.400 ;
        RECT 453.150 342.000 454.950 342.600 ;
        RECT 464.100 342.000 465.150 343.800 ;
        RECT 453.150 340.800 465.150 342.000 ;
        RECT 397.950 334.950 400.200 337.050 ;
        RECT 412.950 334.950 415.050 337.050 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 418.950 334.950 421.050 337.050 ;
        RECT 421.950 334.950 424.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 436.950 334.950 439.050 337.050 ;
        RECT 440.550 335.250 446.850 337.050 ;
        RECT 440.550 334.950 445.050 335.250 ;
        RECT 396.150 329.400 398.100 330.300 ;
        RECT 392.400 328.500 398.100 329.400 ;
        RECT 392.400 321.600 393.600 328.500 ;
        RECT 399.000 327.600 400.200 334.950 ;
        RECT 376.800 315.600 378.600 321.600 ;
        RECT 379.800 315.000 381.600 321.600 ;
        RECT 392.400 315.600 394.200 321.600 ;
        RECT 395.400 315.000 397.200 321.600 ;
        RECT 398.400 315.600 400.200 327.600 ;
        RECT 416.850 321.600 418.050 334.950 ;
        RECT 422.100 333.150 423.900 334.950 ;
        RECT 413.400 315.000 415.200 321.600 ;
        RECT 416.400 315.600 418.200 321.600 ;
        RECT 421.500 315.000 423.300 327.600 ;
        RECT 434.400 321.600 435.600 334.950 ;
        RECT 437.100 333.150 438.900 334.950 ;
        RECT 440.550 327.600 441.750 334.950 ;
        RECT 442.950 329.400 444.750 331.200 ;
        RECT 443.850 328.200 448.050 329.400 ;
        RECT 453.150 328.200 454.050 340.800 ;
        RECT 464.100 339.600 471.000 340.800 ;
        RECT 464.100 339.000 465.900 339.600 ;
        RECT 470.100 338.850 471.000 339.600 ;
        RECT 467.100 337.800 468.900 338.400 ;
        RECT 460.950 336.600 468.900 337.800 ;
        RECT 470.100 337.050 471.900 338.850 ;
        RECT 460.950 334.950 463.050 336.600 ;
        RECT 469.950 334.950 472.050 337.050 ;
        RECT 462.750 329.700 464.550 330.000 ;
        RECT 472.950 329.700 473.850 344.400 ;
        RECT 462.750 329.100 473.850 329.700 ;
        RECT 433.800 315.600 435.600 321.600 ;
        RECT 436.800 315.000 438.600 321.600 ;
        RECT 440.550 315.600 442.350 327.600 ;
        RECT 445.950 327.300 448.050 328.200 ;
        RECT 448.950 327.300 454.050 328.200 ;
        RECT 456.150 328.500 473.850 329.100 ;
        RECT 456.150 328.200 464.550 328.500 ;
        RECT 448.950 326.400 449.850 327.300 ;
        RECT 447.150 324.600 449.850 326.400 ;
        RECT 450.750 326.100 452.550 326.400 ;
        RECT 456.150 326.100 457.050 328.200 ;
        RECT 472.950 327.600 473.850 328.500 ;
        RECT 450.750 325.200 457.050 326.100 ;
        RECT 457.950 326.700 459.750 327.300 ;
        RECT 457.950 325.500 465.450 326.700 ;
        RECT 450.750 324.600 452.550 325.200 ;
        RECT 464.250 324.600 465.450 325.500 ;
        RECT 445.950 321.600 449.850 323.700 ;
        RECT 454.950 323.550 456.750 324.300 ;
        RECT 459.750 323.550 461.550 324.300 ;
        RECT 454.950 322.500 461.550 323.550 ;
        RECT 464.250 322.500 469.050 324.600 ;
        RECT 443.550 315.000 445.350 318.600 ;
        RECT 448.050 315.600 449.850 321.600 ;
        RECT 452.250 315.000 454.050 321.600 ;
        RECT 455.850 315.600 457.650 322.500 ;
        RECT 464.250 321.600 465.450 322.500 ;
        RECT 458.850 315.000 460.650 321.600 ;
        RECT 463.650 315.600 465.450 321.600 ;
        RECT 469.050 315.000 470.850 321.600 ;
        RECT 472.050 315.600 473.850 327.600 ;
        RECT 484.800 344.400 486.600 350.400 ;
        RECT 487.800 347.400 489.600 351.000 ;
        RECT 490.800 347.400 492.600 350.400 ;
        RECT 484.800 337.050 486.000 344.400 ;
        RECT 491.400 343.500 492.600 347.400 ;
        RECT 500.400 345.300 502.200 350.400 ;
        RECT 503.400 346.200 505.200 351.000 ;
        RECT 506.400 345.300 508.200 350.400 ;
        RECT 500.400 343.950 508.200 345.300 ;
        RECT 509.400 344.400 511.200 350.400 ;
        RECT 486.900 342.600 492.600 343.500 ;
        RECT 486.900 341.700 488.850 342.600 ;
        RECT 509.400 342.300 510.600 344.400 ;
        RECT 524.400 343.200 526.200 350.400 ;
        RECT 529.500 344.400 531.300 351.000 ;
        RECT 533.550 344.400 535.350 350.400 ;
        RECT 536.850 347.400 538.650 351.000 ;
        RECT 541.650 347.400 543.450 350.400 ;
        RECT 545.850 347.400 547.650 351.000 ;
        RECT 549.450 347.400 551.250 350.400 ;
        RECT 552.750 347.400 554.550 351.000 ;
        RECT 557.250 348.300 559.050 350.400 ;
        RECT 557.250 347.400 561.000 348.300 ;
        RECT 562.050 347.400 563.850 351.000 ;
        RECT 541.650 346.500 542.700 347.400 ;
        RECT 538.950 345.300 542.700 346.500 ;
        RECT 550.200 346.500 551.250 347.400 ;
        RECT 559.950 346.500 561.000 347.400 ;
        RECT 550.200 345.450 555.150 346.500 ;
        RECT 538.950 344.400 541.050 345.300 ;
        RECT 553.350 344.700 555.150 345.450 ;
        RECT 524.400 342.300 528.600 343.200 ;
        RECT 484.800 334.950 487.050 337.050 ;
        RECT 484.800 327.600 486.000 334.950 ;
        RECT 487.950 330.300 488.850 341.700 ;
        RECT 506.850 341.250 510.600 342.300 ;
        RECT 503.100 337.050 504.900 338.850 ;
        RECT 506.850 337.050 508.050 341.250 ;
        RECT 511.950 339.450 514.050 340.050 ;
        RECT 517.950 339.450 520.050 340.050 ;
        RECT 509.100 337.050 510.900 338.850 ;
        RECT 511.950 338.550 520.050 339.450 ;
        RECT 511.950 337.950 514.050 338.550 ;
        RECT 517.950 337.950 520.050 338.550 ;
        RECT 524.100 337.200 525.900 339.000 ;
        RECT 527.400 337.200 528.600 342.300 ;
        RECT 530.100 337.200 531.900 339.000 ;
        RECT 490.950 334.950 493.050 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 505.950 334.950 508.050 337.050 ;
        RECT 508.950 334.950 511.050 337.050 ;
        RECT 523.950 335.100 526.050 337.200 ;
        RECT 526.950 335.100 529.050 337.200 ;
        RECT 529.950 335.100 532.050 337.200 ;
        RECT 533.550 337.050 534.750 344.400 ;
        RECT 556.650 343.800 558.450 345.600 ;
        RECT 559.950 344.400 562.050 346.500 ;
        RECT 565.050 344.400 566.850 350.400 ;
        RECT 546.150 342.000 547.950 342.600 ;
        RECT 557.100 342.000 558.150 343.800 ;
        RECT 546.150 340.800 558.150 342.000 ;
        RECT 533.550 335.250 539.850 337.050 ;
        RECT 491.100 333.150 492.900 334.950 ;
        RECT 500.100 333.150 501.900 334.950 ;
        RECT 486.900 329.400 488.850 330.300 ;
        RECT 486.900 328.500 492.600 329.400 ;
        RECT 484.800 315.600 486.600 327.600 ;
        RECT 491.400 321.600 492.600 328.500 ;
        RECT 487.800 315.000 489.600 321.600 ;
        RECT 490.800 315.600 492.600 321.600 ;
        RECT 500.700 315.000 502.500 327.600 ;
        RECT 505.950 321.600 507.150 334.950 ;
        RECT 527.400 321.600 528.600 335.100 ;
        RECT 533.550 334.950 538.050 335.250 ;
        RECT 533.550 327.600 534.750 334.950 ;
        RECT 535.950 329.400 537.750 331.200 ;
        RECT 536.850 328.200 541.050 329.400 ;
        RECT 546.150 328.200 547.050 340.800 ;
        RECT 557.100 339.600 564.000 340.800 ;
        RECT 557.100 339.000 558.900 339.600 ;
        RECT 563.100 338.850 564.000 339.600 ;
        RECT 560.100 337.800 561.900 338.400 ;
        RECT 553.950 336.600 561.900 337.800 ;
        RECT 563.100 337.050 564.900 338.850 ;
        RECT 553.950 334.950 556.050 336.600 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 555.750 329.700 557.550 330.000 ;
        RECT 565.950 329.700 566.850 344.400 ;
        RECT 575.400 345.300 577.200 350.400 ;
        RECT 578.400 346.200 580.200 351.000 ;
        RECT 581.400 345.300 583.200 350.400 ;
        RECT 575.400 343.950 583.200 345.300 ;
        RECT 584.400 344.400 586.200 350.400 ;
        RECT 598.800 347.400 600.600 350.400 ;
        RECT 601.800 347.400 603.600 351.000 ;
        RECT 584.400 342.300 585.600 344.400 ;
        RECT 581.850 341.250 585.600 342.300 ;
        RECT 578.100 337.050 579.900 338.850 ;
        RECT 581.850 337.050 583.050 341.250 ;
        RECT 584.100 337.050 585.900 338.850 ;
        RECT 599.400 337.050 600.600 347.400 ;
        RECT 606.150 344.400 607.950 350.400 ;
        RECT 609.150 347.400 610.950 351.000 ;
        RECT 613.950 348.300 615.750 350.400 ;
        RECT 612.000 347.400 615.750 348.300 ;
        RECT 618.450 347.400 620.250 351.000 ;
        RECT 621.750 347.400 623.550 350.400 ;
        RECT 625.350 347.400 627.150 351.000 ;
        RECT 629.550 347.400 631.350 350.400 ;
        RECT 634.350 347.400 636.150 351.000 ;
        RECT 612.000 346.500 613.050 347.400 ;
        RECT 621.750 346.500 622.800 347.400 ;
        RECT 610.950 344.400 613.050 346.500 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 601.950 334.950 604.050 337.050 ;
        RECT 575.100 333.150 576.900 334.950 ;
        RECT 555.750 329.100 566.850 329.700 ;
        RECT 505.800 315.600 507.600 321.600 ;
        RECT 508.800 315.000 510.600 321.600 ;
        RECT 523.800 315.000 525.600 321.600 ;
        RECT 526.800 315.600 528.600 321.600 ;
        RECT 529.800 315.000 531.600 321.600 ;
        RECT 533.550 315.600 535.350 327.600 ;
        RECT 538.950 327.300 541.050 328.200 ;
        RECT 541.950 327.300 547.050 328.200 ;
        RECT 549.150 328.500 566.850 329.100 ;
        RECT 549.150 328.200 557.550 328.500 ;
        RECT 541.950 326.400 542.850 327.300 ;
        RECT 540.150 324.600 542.850 326.400 ;
        RECT 543.750 326.100 545.550 326.400 ;
        RECT 549.150 326.100 550.050 328.200 ;
        RECT 565.950 327.600 566.850 328.500 ;
        RECT 543.750 325.200 550.050 326.100 ;
        RECT 550.950 326.700 552.750 327.300 ;
        RECT 550.950 325.500 558.450 326.700 ;
        RECT 543.750 324.600 545.550 325.200 ;
        RECT 557.250 324.600 558.450 325.500 ;
        RECT 538.950 321.600 542.850 323.700 ;
        RECT 547.950 323.550 549.750 324.300 ;
        RECT 552.750 323.550 554.550 324.300 ;
        RECT 547.950 322.500 554.550 323.550 ;
        RECT 557.250 322.500 562.050 324.600 ;
        RECT 536.550 315.000 538.350 318.600 ;
        RECT 541.050 315.600 542.850 321.600 ;
        RECT 545.250 315.000 547.050 321.600 ;
        RECT 548.850 315.600 550.650 322.500 ;
        RECT 557.250 321.600 558.450 322.500 ;
        RECT 551.850 315.000 553.650 321.600 ;
        RECT 556.650 315.600 558.450 321.600 ;
        RECT 562.050 315.000 563.850 321.600 ;
        RECT 565.050 315.600 566.850 327.600 ;
        RECT 575.700 315.000 577.500 327.600 ;
        RECT 580.950 321.600 582.150 334.950 ;
        RECT 583.950 324.450 586.050 325.050 ;
        RECT 589.950 324.450 592.050 324.900 ;
        RECT 583.950 323.550 592.050 324.450 ;
        RECT 583.950 322.950 586.050 323.550 ;
        RECT 589.950 322.800 592.050 323.550 ;
        RECT 599.400 321.600 600.600 334.950 ;
        RECT 602.100 333.150 603.900 334.950 ;
        RECT 606.150 329.700 607.050 344.400 ;
        RECT 614.550 343.800 616.350 345.600 ;
        RECT 617.850 345.450 622.800 346.500 ;
        RECT 630.300 346.500 631.350 347.400 ;
        RECT 617.850 344.700 619.650 345.450 ;
        RECT 630.300 345.300 634.050 346.500 ;
        RECT 631.950 344.400 634.050 345.300 ;
        RECT 637.650 344.400 639.450 350.400 ;
        RECT 614.850 342.000 615.900 343.800 ;
        RECT 625.050 342.000 626.850 342.600 ;
        RECT 614.850 340.800 626.850 342.000 ;
        RECT 609.000 339.600 615.900 340.800 ;
        RECT 609.000 338.850 609.900 339.600 ;
        RECT 614.100 339.000 615.900 339.600 ;
        RECT 608.100 337.050 609.900 338.850 ;
        RECT 611.100 337.800 612.900 338.400 ;
        RECT 607.950 334.950 610.050 337.050 ;
        RECT 611.100 336.600 619.050 337.800 ;
        RECT 616.950 334.950 619.050 336.600 ;
        RECT 615.450 329.700 617.250 330.000 ;
        RECT 606.150 329.100 617.250 329.700 ;
        RECT 606.150 328.500 623.850 329.100 ;
        RECT 606.150 327.600 607.050 328.500 ;
        RECT 615.450 328.200 623.850 328.500 ;
        RECT 580.800 315.600 582.600 321.600 ;
        RECT 583.800 315.000 585.600 321.600 ;
        RECT 598.800 315.600 600.600 321.600 ;
        RECT 601.800 315.000 603.600 321.600 ;
        RECT 606.150 315.600 607.950 327.600 ;
        RECT 620.250 326.700 622.050 327.300 ;
        RECT 614.550 325.500 622.050 326.700 ;
        RECT 622.950 326.100 623.850 328.200 ;
        RECT 625.950 328.200 626.850 340.800 ;
        RECT 638.250 337.050 639.450 344.400 ;
        RECT 650.400 343.200 652.200 350.400 ;
        RECT 655.500 344.400 657.300 351.000 ;
        RECT 665.400 350.400 666.600 351.000 ;
        RECT 665.400 347.400 667.200 350.400 ;
        RECT 668.400 347.400 670.200 350.400 ;
        RECT 671.400 347.400 673.200 351.000 ;
        RECT 669.300 343.200 670.200 347.400 ;
        RECT 674.400 344.400 676.200 350.400 ;
        RECT 643.950 340.950 646.050 343.050 ;
        RECT 650.400 342.300 654.600 343.200 ;
        RECT 669.300 342.300 672.600 343.200 ;
        RECT 633.150 335.250 639.450 337.050 ;
        RECT 634.950 334.950 639.450 335.250 ;
        RECT 635.250 329.400 637.050 331.200 ;
        RECT 631.950 328.200 636.150 329.400 ;
        RECT 625.950 327.300 631.050 328.200 ;
        RECT 631.950 327.300 634.050 328.200 ;
        RECT 638.250 327.600 639.450 334.950 ;
        RECT 644.550 334.050 645.450 340.950 ;
        RECT 650.100 337.200 651.900 339.000 ;
        RECT 653.400 337.200 654.600 342.300 ;
        RECT 670.800 341.400 672.600 342.300 ;
        RECT 656.100 337.200 657.900 339.000 ;
        RECT 649.950 335.100 652.050 337.200 ;
        RECT 652.950 335.100 655.050 337.200 ;
        RECT 655.950 335.100 658.050 337.200 ;
        RECT 665.100 337.050 666.900 338.850 ;
        RECT 644.550 332.550 649.050 334.050 ;
        RECT 645.000 331.950 649.050 332.550 ;
        RECT 630.150 326.400 631.050 327.300 ;
        RECT 627.450 326.100 629.250 326.400 ;
        RECT 614.550 324.600 615.750 325.500 ;
        RECT 622.950 325.200 629.250 326.100 ;
        RECT 627.450 324.600 629.250 325.200 ;
        RECT 630.150 324.600 632.850 326.400 ;
        RECT 610.950 322.500 615.750 324.600 ;
        RECT 618.450 323.550 620.250 324.300 ;
        RECT 623.250 323.550 625.050 324.300 ;
        RECT 618.450 322.500 625.050 323.550 ;
        RECT 614.550 321.600 615.750 322.500 ;
        RECT 609.150 315.000 610.950 321.600 ;
        RECT 614.550 315.600 616.350 321.600 ;
        RECT 619.350 315.000 621.150 321.600 ;
        RECT 622.350 315.600 624.150 322.500 ;
        RECT 630.150 321.600 634.050 323.700 ;
        RECT 625.950 315.000 627.750 321.600 ;
        RECT 630.150 315.600 631.950 321.600 ;
        RECT 634.650 315.000 636.450 318.600 ;
        RECT 637.650 315.600 639.450 327.600 ;
        RECT 653.400 321.600 654.600 335.100 ;
        RECT 664.950 334.950 667.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 668.100 333.150 669.900 334.950 ;
        RECT 671.700 330.900 672.600 341.400 ;
        RECT 675.000 337.050 676.050 344.400 ;
        RECT 686.400 342.600 688.200 350.400 ;
        RECT 690.900 344.400 692.700 351.000 ;
        RECT 693.900 346.200 695.700 350.400 ;
        RECT 693.900 344.400 696.600 346.200 ;
        RECT 709.800 344.400 711.600 350.400 ;
        RECT 692.100 342.600 693.900 343.500 ;
        RECT 686.400 341.700 693.900 342.600 ;
        RECT 686.100 337.200 687.900 339.000 ;
        RECT 670.800 330.300 672.600 330.900 ;
        RECT 665.400 329.100 672.600 330.300 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 685.950 335.100 688.050 337.200 ;
        RECT 665.400 327.600 666.600 329.100 ;
        RECT 673.950 327.600 675.300 334.950 ;
        RECT 649.800 315.000 651.600 321.600 ;
        RECT 652.800 315.600 654.600 321.600 ;
        RECT 655.800 315.000 657.600 321.600 ;
        RECT 665.400 315.600 667.200 327.600 ;
        RECT 669.900 315.000 671.700 327.600 ;
        RECT 672.900 326.100 675.300 327.600 ;
        RECT 672.900 315.600 674.700 326.100 ;
        RECT 689.400 321.600 690.300 341.700 ;
        RECT 695.700 337.200 696.600 344.400 ;
        RECT 710.400 342.300 711.600 344.400 ;
        RECT 712.800 345.300 714.600 350.400 ;
        RECT 715.800 346.200 717.600 351.000 ;
        RECT 718.800 345.300 720.600 350.400 ;
        RECT 730.800 347.400 732.600 350.400 ;
        RECT 733.800 347.400 735.600 351.000 ;
        RECT 743.400 347.400 745.200 351.000 ;
        RECT 746.400 347.400 748.200 350.400 ;
        RECT 749.400 347.400 751.200 351.000 ;
        RECT 761.400 347.400 763.200 351.000 ;
        RECT 764.400 347.400 766.200 350.400 ;
        RECT 767.400 347.400 769.200 351.000 ;
        RECT 779.400 347.400 781.200 351.000 ;
        RECT 782.400 347.400 784.200 350.400 ;
        RECT 785.400 347.400 787.200 351.000 ;
        RECT 797.400 347.400 799.200 351.000 ;
        RECT 800.400 347.400 802.200 350.400 ;
        RECT 803.400 347.400 805.200 351.000 ;
        RECT 817.800 347.400 819.600 350.400 ;
        RECT 820.800 347.400 822.600 351.000 ;
        RECT 712.800 343.950 720.600 345.300 ;
        RECT 710.400 341.250 714.150 342.300 ;
        RECT 691.950 335.100 694.050 337.200 ;
        RECT 694.950 335.100 697.050 337.200 ;
        RECT 710.100 337.050 711.900 338.850 ;
        RECT 712.950 337.050 714.150 341.250 ;
        RECT 716.100 337.050 717.900 338.850 ;
        RECT 731.400 337.050 732.600 347.400 ;
        RECT 746.700 337.050 747.600 347.400 ;
        RECT 748.950 342.450 751.050 343.050 ;
        RECT 757.950 342.450 760.050 343.050 ;
        RECT 748.950 341.550 760.050 342.450 ;
        RECT 748.950 340.950 751.050 341.550 ;
        RECT 757.950 340.950 760.050 341.550 ;
        RECT 764.700 337.050 765.600 347.400 ;
        RECT 782.700 337.050 783.600 347.400 ;
        RECT 800.700 337.050 801.600 347.400 ;
        RECT 818.400 337.050 819.600 347.400 ;
        RECT 833.400 343.200 835.200 350.400 ;
        RECT 838.500 344.400 840.300 351.000 ;
        RECT 848.700 344.400 850.500 351.000 ;
        RECT 853.800 343.200 855.600 350.400 ;
        RECT 833.400 342.300 837.600 343.200 ;
        RECT 833.100 337.200 834.900 339.000 ;
        RECT 836.400 337.200 837.600 342.300 ;
        RECT 851.400 342.300 855.600 343.200 ;
        RECT 839.100 337.200 840.900 339.000 ;
        RECT 848.100 337.200 849.900 339.000 ;
        RECT 851.400 337.200 852.600 342.300 ;
        RECT 854.100 337.200 855.900 339.000 ;
        RECT 692.100 333.300 693.900 335.100 ;
        RECT 695.700 327.600 696.600 335.100 ;
        RECT 709.950 334.950 712.050 337.050 ;
        RECT 712.950 334.950 715.050 337.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 730.950 334.950 733.050 337.050 ;
        RECT 733.950 334.950 736.050 337.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 778.950 334.950 781.050 337.050 ;
        RECT 781.950 334.950 784.050 337.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 799.950 334.950 802.050 337.050 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 817.950 334.950 820.050 337.050 ;
        RECT 820.950 334.950 823.050 337.050 ;
        RECT 832.950 335.100 835.050 337.200 ;
        RECT 835.950 335.100 838.050 337.200 ;
        RECT 838.950 335.100 841.050 337.200 ;
        RECT 847.950 335.100 850.050 337.200 ;
        RECT 850.950 335.100 853.050 337.200 ;
        RECT 853.950 335.100 856.050 337.200 ;
        RECT 686.400 315.000 688.200 321.600 ;
        RECT 689.400 315.600 691.200 321.600 ;
        RECT 692.400 315.000 694.200 321.600 ;
        RECT 695.400 315.600 697.200 327.600 ;
        RECT 713.850 321.600 715.050 334.950 ;
        RECT 719.100 333.150 720.900 334.950 ;
        RECT 710.400 315.000 712.200 321.600 ;
        RECT 713.400 315.600 715.200 321.600 ;
        RECT 718.500 315.000 720.300 327.600 ;
        RECT 731.400 321.600 732.600 334.950 ;
        RECT 734.100 333.150 735.900 334.950 ;
        RECT 743.100 333.150 744.900 334.950 ;
        RECT 746.700 327.600 747.600 334.950 ;
        RECT 749.100 333.150 750.900 334.950 ;
        RECT 761.100 333.150 762.900 334.950 ;
        RECT 764.700 327.600 765.600 334.950 ;
        RECT 767.100 333.150 768.900 334.950 ;
        RECT 779.100 333.150 780.900 334.950 ;
        RECT 782.700 327.600 783.600 334.950 ;
        RECT 785.100 333.150 786.900 334.950 ;
        RECT 797.100 333.150 798.900 334.950 ;
        RECT 800.700 327.600 801.600 334.950 ;
        RECT 803.100 333.150 804.900 334.950 ;
        RECT 730.800 315.600 732.600 321.600 ;
        RECT 733.800 315.000 735.600 321.600 ;
        RECT 743.400 315.000 745.200 327.600 ;
        RECT 746.700 326.400 750.300 327.600 ;
        RECT 748.500 315.600 750.300 326.400 ;
        RECT 761.400 315.000 763.200 327.600 ;
        RECT 764.700 326.400 768.300 327.600 ;
        RECT 766.500 315.600 768.300 326.400 ;
        RECT 779.400 315.000 781.200 327.600 ;
        RECT 782.700 326.400 786.300 327.600 ;
        RECT 784.500 315.600 786.300 326.400 ;
        RECT 797.400 315.000 799.200 327.600 ;
        RECT 800.700 326.400 804.300 327.600 ;
        RECT 802.500 315.600 804.300 326.400 ;
        RECT 818.400 321.600 819.600 334.950 ;
        RECT 821.100 333.150 822.900 334.950 ;
        RECT 823.950 333.450 826.050 334.050 ;
        RECT 832.950 333.450 835.050 334.050 ;
        RECT 823.950 332.550 835.050 333.450 ;
        RECT 823.950 331.950 826.050 332.550 ;
        RECT 832.950 331.950 835.050 332.550 ;
        RECT 836.400 321.600 837.600 335.100 ;
        RECT 851.400 321.600 852.600 335.100 ;
        RECT 817.800 315.600 819.600 321.600 ;
        RECT 820.800 315.000 822.600 321.600 ;
        RECT 832.800 315.000 834.600 321.600 ;
        RECT 835.800 315.600 837.600 321.600 ;
        RECT 838.800 315.000 840.600 321.600 ;
        RECT 848.400 315.000 850.200 321.600 ;
        RECT 851.400 315.600 853.200 321.600 ;
        RECT 854.400 315.000 856.200 321.600 ;
        RECT 10.800 305.400 12.600 312.000 ;
        RECT 13.800 305.400 15.600 311.400 ;
        RECT 16.800 305.400 18.600 312.000 ;
        RECT 14.400 291.900 15.600 305.400 ;
        RECT 26.400 299.400 28.200 312.000 ;
        RECT 30.900 299.400 34.200 311.400 ;
        RECT 36.900 299.400 38.700 312.000 ;
        RECT 45.150 299.400 46.950 311.400 ;
        RECT 48.150 305.400 49.950 312.000 ;
        RECT 53.550 305.400 55.350 311.400 ;
        RECT 58.350 305.400 60.150 312.000 ;
        RECT 53.550 304.500 54.750 305.400 ;
        RECT 61.350 304.500 63.150 311.400 ;
        RECT 64.950 305.400 66.750 312.000 ;
        RECT 69.150 305.400 70.950 311.400 ;
        RECT 73.650 308.400 75.450 312.000 ;
        RECT 49.950 302.400 54.750 304.500 ;
        RECT 57.450 303.450 64.050 304.500 ;
        RECT 57.450 302.700 59.250 303.450 ;
        RECT 62.250 302.700 64.050 303.450 ;
        RECT 69.150 303.300 73.050 305.400 ;
        RECT 53.550 301.500 54.750 302.400 ;
        RECT 66.450 301.800 68.250 302.400 ;
        RECT 53.550 300.300 61.050 301.500 ;
        RECT 59.250 299.700 61.050 300.300 ;
        RECT 61.950 300.900 68.250 301.800 ;
        RECT 26.100 291.900 27.900 293.700 ;
        RECT 32.100 291.900 33.300 299.400 ;
        RECT 45.150 298.500 46.050 299.400 ;
        RECT 61.950 298.800 62.850 300.900 ;
        RECT 66.450 300.600 68.250 300.900 ;
        RECT 69.150 300.600 71.850 302.400 ;
        RECT 69.150 299.700 70.050 300.600 ;
        RECT 54.450 298.500 62.850 298.800 ;
        RECT 45.150 297.900 62.850 298.500 ;
        RECT 64.950 298.800 70.050 299.700 ;
        RECT 70.950 298.800 73.050 299.700 ;
        RECT 76.650 299.400 78.450 311.400 ;
        RECT 45.150 297.300 56.250 297.900 ;
        RECT 38.100 291.900 39.900 293.700 ;
        RECT 10.950 289.800 13.050 291.900 ;
        RECT 13.950 289.800 16.050 291.900 ;
        RECT 16.950 289.800 19.050 291.900 ;
        RECT 25.950 289.800 28.050 291.900 ;
        RECT 28.950 289.800 31.050 291.900 ;
        RECT 31.950 289.800 34.050 291.900 ;
        RECT 34.950 289.800 37.050 291.900 ;
        RECT 37.950 289.800 40.050 291.900 ;
        RECT 11.100 288.000 12.900 289.800 ;
        RECT 14.400 284.700 15.600 289.800 ;
        RECT 17.100 288.000 18.900 289.800 ;
        RECT 29.100 288.000 30.900 289.800 ;
        RECT 31.950 287.400 33.000 289.800 ;
        RECT 35.100 288.000 36.900 289.800 ;
        RECT 11.400 283.800 15.600 284.700 ;
        RECT 32.100 285.300 33.300 287.400 ;
        RECT 32.100 284.100 36.600 285.300 ;
        RECT 11.400 276.600 13.200 283.800 ;
        RECT 16.500 276.000 18.300 282.600 ;
        RECT 26.400 282.000 34.200 282.900 ;
        RECT 35.700 282.600 36.600 284.100 ;
        RECT 45.150 282.600 46.050 297.300 ;
        RECT 54.450 297.000 56.250 297.300 ;
        RECT 46.950 289.950 49.050 292.050 ;
        RECT 55.950 290.400 58.050 292.050 ;
        RECT 47.100 288.150 48.900 289.950 ;
        RECT 50.100 289.200 58.050 290.400 ;
        RECT 50.100 288.600 51.900 289.200 ;
        RECT 48.000 287.400 48.900 288.150 ;
        RECT 53.100 287.400 54.900 288.000 ;
        RECT 48.000 286.200 54.900 287.400 ;
        RECT 64.950 286.200 65.850 298.800 ;
        RECT 70.950 297.600 75.150 298.800 ;
        RECT 74.250 295.800 76.050 297.600 ;
        RECT 77.250 292.050 78.450 299.400 ;
        RECT 73.950 291.750 78.450 292.050 ;
        RECT 72.150 289.950 78.450 291.750 ;
        RECT 53.850 285.000 65.850 286.200 ;
        RECT 53.850 283.200 54.900 285.000 ;
        RECT 64.050 284.400 65.850 285.000 ;
        RECT 26.400 276.600 28.200 282.000 ;
        RECT 29.400 276.000 31.200 281.100 ;
        RECT 32.400 277.500 34.200 282.000 ;
        RECT 35.400 278.400 37.200 282.600 ;
        RECT 38.400 277.500 40.200 282.600 ;
        RECT 32.400 276.600 40.200 277.500 ;
        RECT 45.150 276.600 46.950 282.600 ;
        RECT 49.950 280.500 52.050 282.600 ;
        RECT 53.550 281.400 55.350 283.200 ;
        RECT 77.250 282.600 78.450 289.950 ;
        RECT 56.850 281.550 58.650 282.300 ;
        RECT 70.950 281.700 73.050 282.600 ;
        RECT 56.850 280.500 61.800 281.550 ;
        RECT 51.000 279.600 52.050 280.500 ;
        RECT 60.750 279.600 61.800 280.500 ;
        RECT 69.300 280.500 73.050 281.700 ;
        RECT 69.300 279.600 70.350 280.500 ;
        RECT 48.150 276.000 49.950 279.600 ;
        RECT 51.000 278.700 54.750 279.600 ;
        RECT 52.950 276.600 54.750 278.700 ;
        RECT 57.450 276.000 59.250 279.600 ;
        RECT 60.750 276.600 62.550 279.600 ;
        RECT 64.350 276.000 66.150 279.600 ;
        RECT 68.550 276.600 70.350 279.600 ;
        RECT 73.350 276.000 75.150 279.600 ;
        RECT 76.650 276.600 78.450 282.600 ;
        RECT 81.150 299.400 82.950 311.400 ;
        RECT 84.150 305.400 85.950 312.000 ;
        RECT 89.550 305.400 91.350 311.400 ;
        RECT 94.350 305.400 96.150 312.000 ;
        RECT 89.550 304.500 90.750 305.400 ;
        RECT 97.350 304.500 99.150 311.400 ;
        RECT 100.950 305.400 102.750 312.000 ;
        RECT 105.150 305.400 106.950 311.400 ;
        RECT 109.650 308.400 111.450 312.000 ;
        RECT 85.950 302.400 90.750 304.500 ;
        RECT 93.450 303.450 100.050 304.500 ;
        RECT 93.450 302.700 95.250 303.450 ;
        RECT 98.250 302.700 100.050 303.450 ;
        RECT 105.150 303.300 109.050 305.400 ;
        RECT 89.550 301.500 90.750 302.400 ;
        RECT 102.450 301.800 104.250 302.400 ;
        RECT 89.550 300.300 97.050 301.500 ;
        RECT 95.250 299.700 97.050 300.300 ;
        RECT 97.950 300.900 104.250 301.800 ;
        RECT 81.150 298.500 82.050 299.400 ;
        RECT 97.950 298.800 98.850 300.900 ;
        RECT 102.450 300.600 104.250 300.900 ;
        RECT 105.150 300.600 107.850 302.400 ;
        RECT 105.150 299.700 106.050 300.600 ;
        RECT 90.450 298.500 98.850 298.800 ;
        RECT 81.150 297.900 98.850 298.500 ;
        RECT 100.950 298.800 106.050 299.700 ;
        RECT 106.950 298.800 109.050 299.700 ;
        RECT 112.650 299.400 114.450 311.400 ;
        RECT 124.800 305.400 126.600 312.000 ;
        RECT 127.800 305.400 129.600 311.400 ;
        RECT 130.800 305.400 132.600 312.000 ;
        RECT 143.400 305.400 145.200 312.000 ;
        RECT 146.400 305.400 148.200 311.400 ;
        RECT 81.150 297.300 92.250 297.900 ;
        RECT 81.150 282.600 82.050 297.300 ;
        RECT 90.450 297.000 92.250 297.300 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 91.950 290.400 94.050 292.050 ;
        RECT 83.100 288.150 84.900 289.950 ;
        RECT 86.100 289.200 94.050 290.400 ;
        RECT 86.100 288.600 87.900 289.200 ;
        RECT 84.000 287.400 84.900 288.150 ;
        RECT 89.100 287.400 90.900 288.000 ;
        RECT 84.000 286.200 90.900 287.400 ;
        RECT 100.950 286.200 101.850 298.800 ;
        RECT 106.950 297.600 111.150 298.800 ;
        RECT 110.250 295.800 112.050 297.600 ;
        RECT 113.250 292.050 114.450 299.400 ;
        RECT 109.950 291.750 114.450 292.050 ;
        RECT 128.400 291.900 129.600 305.400 ;
        RECT 146.850 292.050 148.050 305.400 ;
        RECT 151.500 299.400 153.300 312.000 ;
        RECT 161.400 305.400 163.200 312.000 ;
        RECT 164.400 305.400 166.200 311.400 ;
        RECT 179.400 305.400 181.200 312.000 ;
        RECT 182.400 305.400 184.200 311.400 ;
        RECT 152.100 292.050 153.900 293.850 ;
        RECT 161.100 292.050 162.900 293.850 ;
        RECT 164.400 292.050 165.600 305.400 ;
        RECT 169.950 297.450 172.050 298.050 ;
        RECT 178.950 297.450 181.050 298.050 ;
        RECT 169.950 296.550 181.050 297.450 ;
        RECT 169.950 295.950 172.050 296.550 ;
        RECT 178.950 295.950 181.050 296.550 ;
        RECT 166.950 294.450 169.050 295.050 ;
        RECT 166.950 293.550 174.450 294.450 ;
        RECT 166.950 292.950 169.050 293.550 ;
        RECT 108.150 289.950 114.450 291.750 ;
        RECT 89.850 285.000 101.850 286.200 ;
        RECT 89.850 283.200 90.900 285.000 ;
        RECT 100.050 284.400 101.850 285.000 ;
        RECT 81.150 276.600 82.950 282.600 ;
        RECT 85.950 280.500 88.050 282.600 ;
        RECT 89.550 281.400 91.350 283.200 ;
        RECT 113.250 282.600 114.450 289.950 ;
        RECT 124.950 289.800 127.050 291.900 ;
        RECT 127.950 289.800 130.050 291.900 ;
        RECT 130.950 289.800 133.050 291.900 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 160.950 289.950 163.050 292.050 ;
        RECT 163.950 289.950 166.050 292.050 ;
        RECT 125.100 288.000 126.900 289.800 ;
        RECT 128.400 284.700 129.600 289.800 ;
        RECT 131.100 288.000 132.900 289.800 ;
        RECT 143.100 288.150 144.900 289.950 ;
        RECT 145.950 285.750 147.150 289.950 ;
        RECT 149.100 288.150 150.900 289.950 ;
        RECT 92.850 281.550 94.650 282.300 ;
        RECT 106.950 281.700 109.050 282.600 ;
        RECT 92.850 280.500 97.800 281.550 ;
        RECT 87.000 279.600 88.050 280.500 ;
        RECT 96.750 279.600 97.800 280.500 ;
        RECT 105.300 280.500 109.050 281.700 ;
        RECT 105.300 279.600 106.350 280.500 ;
        RECT 84.150 276.000 85.950 279.600 ;
        RECT 87.000 278.700 90.750 279.600 ;
        RECT 88.950 276.600 90.750 278.700 ;
        RECT 93.450 276.000 95.250 279.600 ;
        RECT 96.750 276.600 98.550 279.600 ;
        RECT 100.350 276.000 102.150 279.600 ;
        RECT 104.550 276.600 106.350 279.600 ;
        RECT 109.350 276.000 111.150 279.600 ;
        RECT 112.650 276.600 114.450 282.600 ;
        RECT 125.400 283.800 129.600 284.700 ;
        RECT 143.400 284.700 147.150 285.750 ;
        RECT 125.400 276.600 127.200 283.800 ;
        RECT 143.400 282.600 144.600 284.700 ;
        RECT 130.500 276.000 132.300 282.600 ;
        RECT 142.800 276.600 144.600 282.600 ;
        RECT 145.800 281.700 153.600 283.050 ;
        RECT 145.800 276.600 147.600 281.700 ;
        RECT 148.800 276.000 150.600 280.800 ;
        RECT 151.800 276.600 153.600 281.700 ;
        RECT 164.400 279.600 165.600 289.950 ;
        RECT 173.550 289.050 174.450 293.550 ;
        RECT 182.850 292.050 184.050 305.400 ;
        RECT 187.500 299.400 189.300 312.000 ;
        RECT 199.800 305.400 201.600 312.000 ;
        RECT 202.800 305.400 204.600 311.400 ;
        RECT 205.800 305.400 207.600 312.000 ;
        RECT 217.800 305.400 219.600 312.000 ;
        RECT 220.800 305.400 222.600 311.400 ;
        RECT 223.800 305.400 225.600 312.000 ;
        RECT 188.100 292.050 189.900 293.850 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 184.950 289.950 187.050 292.050 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 203.400 291.900 204.600 305.400 ;
        RECT 205.950 294.450 208.050 295.050 ;
        RECT 211.950 294.450 214.050 295.050 ;
        RECT 205.950 293.550 214.050 294.450 ;
        RECT 205.950 292.950 208.050 293.550 ;
        RECT 211.950 292.950 214.050 293.550 ;
        RECT 221.400 291.900 222.600 305.400 ;
        RECT 233.400 300.300 235.200 311.400 ;
        RECT 233.400 299.400 237.900 300.300 ;
        RECT 240.900 299.400 242.700 311.400 ;
        RECT 248.400 300.600 250.200 311.400 ;
        RECT 235.800 297.300 237.900 299.400 ;
        RECT 241.500 297.900 242.700 299.400 ;
        RECT 245.400 299.400 250.200 300.600 ;
        RECT 262.800 299.400 264.600 311.400 ;
        RECT 265.800 300.300 267.600 311.400 ;
        RECT 268.800 301.200 270.600 312.000 ;
        RECT 271.800 300.300 273.600 311.400 ;
        RECT 283.800 305.400 285.600 311.400 ;
        RECT 286.800 306.000 288.600 312.000 ;
        RECT 265.800 299.400 273.600 300.300 ;
        RECT 284.700 305.100 285.600 305.400 ;
        RECT 289.800 305.400 291.600 311.400 ;
        RECT 292.800 305.400 294.600 312.000 ;
        RECT 302.400 305.400 304.200 312.000 ;
        RECT 305.400 305.400 307.200 311.400 ;
        RECT 308.400 305.400 310.200 312.000 ;
        RECT 289.800 305.100 291.300 305.400 ;
        RECT 284.700 304.200 291.300 305.100 ;
        RECT 245.400 298.500 247.500 299.400 ;
        RECT 241.500 297.000 243.000 297.900 ;
        RECT 238.950 295.500 241.050 295.800 ;
        RECT 237.300 293.700 241.050 295.500 ;
        RECT 242.100 294.900 243.000 297.000 ;
        RECT 241.950 292.800 244.050 294.900 ;
        RECT 238.500 291.900 240.300 292.500 ;
        RECT 173.550 287.550 178.050 289.050 ;
        RECT 179.100 288.150 180.900 289.950 ;
        RECT 174.000 286.950 178.050 287.550 ;
        RECT 181.950 285.750 183.150 289.950 ;
        RECT 185.100 288.150 186.900 289.950 ;
        RECT 199.950 289.800 202.050 291.900 ;
        RECT 202.950 289.800 205.050 291.900 ;
        RECT 205.950 289.800 208.050 291.900 ;
        RECT 217.950 289.800 220.050 291.900 ;
        RECT 220.950 289.800 223.050 291.900 ;
        RECT 223.950 289.800 226.050 291.900 ;
        RECT 232.950 290.700 240.300 291.900 ;
        RECT 241.200 291.900 243.600 292.800 ;
        RECT 248.100 291.900 249.900 293.700 ;
        RECT 263.400 291.900 264.300 299.400 ;
        RECT 269.100 291.900 270.900 293.700 ;
        RECT 284.700 291.900 285.600 304.200 ;
        RECT 290.100 291.900 291.900 293.700 ;
        RECT 305.400 291.900 306.600 305.400 ;
        RECT 322.800 299.400 324.600 311.400 ;
        RECT 325.800 305.400 327.600 312.000 ;
        RECT 328.800 305.400 330.600 311.400 ;
        RECT 338.400 305.400 340.200 312.000 ;
        RECT 341.400 305.400 343.200 311.400 ;
        RECT 344.400 305.400 346.200 312.000 ;
        RECT 322.800 292.050 324.000 299.400 ;
        RECT 329.400 298.500 330.600 305.400 ;
        RECT 324.900 297.600 330.600 298.500 ;
        RECT 324.900 296.700 326.850 297.600 ;
        RECT 232.950 289.800 235.050 290.700 ;
        RECT 200.100 288.000 201.900 289.800 ;
        RECT 179.400 284.700 183.150 285.750 ;
        RECT 203.400 284.700 204.600 289.800 ;
        RECT 206.100 288.000 207.900 289.800 ;
        RECT 218.100 288.000 219.900 289.800 ;
        RECT 221.400 284.700 222.600 289.800 ;
        RECT 224.100 288.000 225.900 289.800 ;
        RECT 233.250 288.000 235.050 289.800 ;
        RECT 238.500 287.400 240.300 289.200 ;
        RECT 238.200 285.300 240.300 287.400 ;
        RECT 179.400 282.600 180.600 284.700 ;
        RECT 200.400 283.800 204.600 284.700 ;
        RECT 218.400 283.800 222.600 284.700 ;
        RECT 234.000 284.400 240.300 285.300 ;
        RECT 241.200 286.200 242.250 291.900 ;
        RECT 243.600 289.200 245.400 291.000 ;
        RECT 247.950 289.800 250.050 291.900 ;
        RECT 262.950 289.800 265.050 291.900 ;
        RECT 265.950 289.800 268.050 291.900 ;
        RECT 268.950 289.800 271.050 291.900 ;
        RECT 271.950 289.800 274.050 291.900 ;
        RECT 283.950 289.800 286.050 291.900 ;
        RECT 286.950 289.800 289.050 291.900 ;
        RECT 289.950 289.800 292.050 291.900 ;
        RECT 292.950 289.800 295.050 291.900 ;
        RECT 301.950 289.800 304.050 291.900 ;
        RECT 304.950 289.800 307.050 291.900 ;
        RECT 307.950 289.800 310.050 291.900 ;
        RECT 322.800 289.950 325.050 292.050 ;
        RECT 243.150 287.100 245.250 289.200 ;
        RECT 161.400 276.000 163.200 279.600 ;
        RECT 164.400 276.600 166.200 279.600 ;
        RECT 178.800 276.600 180.600 282.600 ;
        RECT 181.800 281.700 189.600 283.050 ;
        RECT 181.800 276.600 183.600 281.700 ;
        RECT 184.800 276.000 186.600 280.800 ;
        RECT 187.800 276.600 189.600 281.700 ;
        RECT 200.400 276.600 202.200 283.800 ;
        RECT 205.500 276.000 207.300 282.600 ;
        RECT 218.400 276.600 220.200 283.800 ;
        RECT 234.000 282.600 235.200 284.400 ;
        RECT 241.200 284.100 244.050 286.200 ;
        RECT 241.200 282.600 242.400 284.100 ;
        RECT 245.400 283.500 247.500 284.700 ;
        RECT 245.400 282.600 250.200 283.500 ;
        RECT 223.500 276.000 225.300 282.600 ;
        RECT 233.400 276.600 235.200 282.600 ;
        RECT 240.900 276.600 242.700 282.600 ;
        RECT 248.400 276.600 250.200 282.600 ;
        RECT 263.400 282.600 264.300 289.800 ;
        RECT 266.100 288.000 267.900 289.800 ;
        RECT 272.100 288.000 273.900 289.800 ;
        RECT 284.700 286.200 285.600 289.800 ;
        RECT 287.100 288.000 288.900 289.800 ;
        RECT 293.100 288.000 294.900 289.800 ;
        RECT 302.100 288.000 303.900 289.800 ;
        RECT 265.950 285.450 268.050 286.050 ;
        RECT 277.950 285.450 280.050 286.050 ;
        RECT 265.950 284.550 280.050 285.450 ;
        RECT 284.700 285.000 288.000 286.200 ;
        RECT 265.950 283.950 268.050 284.550 ;
        RECT 277.950 283.950 280.050 284.550 ;
        RECT 263.400 281.400 268.500 282.600 ;
        RECT 263.700 276.000 265.500 279.600 ;
        RECT 266.700 276.600 268.500 281.400 ;
        RECT 271.200 276.000 273.000 282.600 ;
        RECT 286.200 276.600 288.000 285.000 ;
        RECT 292.800 276.000 294.600 285.600 ;
        RECT 305.400 284.700 306.600 289.800 ;
        RECT 308.100 288.000 309.900 289.800 ;
        RECT 305.400 283.800 309.600 284.700 ;
        RECT 302.700 276.000 304.500 282.600 ;
        RECT 307.800 276.600 309.600 283.800 ;
        RECT 322.800 282.600 324.000 289.950 ;
        RECT 325.950 285.300 326.850 296.700 ;
        RECT 329.100 292.050 330.900 293.850 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 341.400 291.900 342.600 305.400 ;
        RECT 359.700 300.600 361.500 311.400 ;
        RECT 359.700 299.400 363.300 300.600 ;
        RECT 364.800 299.400 366.600 312.000 ;
        RECT 376.800 305.400 378.600 312.000 ;
        RECT 379.800 305.400 381.600 311.400 ;
        RECT 382.800 305.400 384.600 312.000 ;
        RECT 394.800 305.400 396.600 312.000 ;
        RECT 397.800 305.400 399.600 311.400 ;
        RECT 400.800 305.400 402.600 312.000 ;
        RECT 413.400 305.400 415.200 312.000 ;
        RECT 416.400 305.400 418.200 311.400 ;
        RECT 354.000 294.450 358.050 295.050 ;
        RECT 353.550 292.950 358.050 294.450 ;
        RECT 337.950 289.800 340.050 291.900 ;
        RECT 340.950 289.800 343.050 291.900 ;
        RECT 343.950 289.800 346.050 291.900 ;
        RECT 338.100 288.000 339.900 289.800 ;
        RECT 324.900 284.400 326.850 285.300 ;
        RECT 341.400 284.700 342.600 289.800 ;
        RECT 344.100 288.000 345.900 289.800 ;
        RECT 353.550 289.050 354.450 292.950 ;
        RECT 359.100 292.050 360.900 293.850 ;
        RECT 362.400 292.050 363.300 299.400 ;
        RECT 365.100 292.050 366.900 293.850 ;
        RECT 358.950 289.950 361.050 292.050 ;
        RECT 361.950 289.950 364.050 292.050 ;
        RECT 364.950 289.950 367.050 292.050 ;
        RECT 380.400 291.900 381.600 305.400 ;
        RECT 385.950 294.450 390.000 295.050 ;
        RECT 385.950 292.950 390.450 294.450 ;
        RECT 353.550 287.550 358.050 289.050 ;
        RECT 354.000 286.950 358.050 287.550 ;
        RECT 324.900 283.500 330.600 284.400 ;
        RECT 341.400 283.800 345.600 284.700 ;
        RECT 322.800 276.600 324.600 282.600 ;
        RECT 329.400 279.600 330.600 283.500 ;
        RECT 325.800 276.000 327.600 279.600 ;
        RECT 328.800 276.600 330.600 279.600 ;
        RECT 338.700 276.000 340.500 282.600 ;
        RECT 343.800 276.600 345.600 283.800 ;
        RECT 362.400 279.600 363.300 289.950 ;
        RECT 376.950 289.800 379.050 291.900 ;
        RECT 379.950 289.800 382.050 291.900 ;
        RECT 382.950 289.800 385.050 291.900 ;
        RECT 377.100 288.000 378.900 289.800 ;
        RECT 380.400 284.700 381.600 289.800 ;
        RECT 383.100 288.000 384.900 289.800 ;
        RECT 389.550 289.050 390.450 292.950 ;
        RECT 398.400 291.900 399.600 305.400 ;
        RECT 416.850 292.050 418.050 305.400 ;
        RECT 421.500 299.400 423.300 312.000 ;
        RECT 433.800 305.400 435.600 311.400 ;
        RECT 436.800 305.400 438.600 312.000 ;
        RECT 422.100 292.050 423.900 293.850 ;
        RECT 434.400 292.050 435.600 305.400 ;
        RECT 440.550 299.400 442.350 311.400 ;
        RECT 443.550 308.400 445.350 312.000 ;
        RECT 448.050 305.400 449.850 311.400 ;
        RECT 452.250 305.400 454.050 312.000 ;
        RECT 445.950 303.300 449.850 305.400 ;
        RECT 455.850 304.500 457.650 311.400 ;
        RECT 458.850 305.400 460.650 312.000 ;
        RECT 463.650 305.400 465.450 311.400 ;
        RECT 469.050 305.400 470.850 312.000 ;
        RECT 464.250 304.500 465.450 305.400 ;
        RECT 454.950 303.450 461.550 304.500 ;
        RECT 454.950 302.700 456.750 303.450 ;
        RECT 459.750 302.700 461.550 303.450 ;
        RECT 464.250 302.400 469.050 304.500 ;
        RECT 447.150 300.600 449.850 302.400 ;
        RECT 450.750 301.800 452.550 302.400 ;
        RECT 450.750 300.900 457.050 301.800 ;
        RECT 464.250 301.500 465.450 302.400 ;
        RECT 450.750 300.600 452.550 300.900 ;
        RECT 448.950 299.700 449.850 300.600 ;
        RECT 437.100 292.050 438.900 293.850 ;
        RECT 440.550 292.050 441.750 299.400 ;
        RECT 445.950 298.800 448.050 299.700 ;
        RECT 448.950 298.800 454.050 299.700 ;
        RECT 443.850 297.600 448.050 298.800 ;
        RECT 442.950 295.800 444.750 297.600 ;
        RECT 394.950 289.800 397.050 291.900 ;
        RECT 397.950 289.800 400.050 291.900 ;
        RECT 400.950 289.800 403.050 291.900 ;
        RECT 412.950 289.950 415.050 292.050 ;
        RECT 415.950 289.950 418.050 292.050 ;
        RECT 418.950 289.950 421.050 292.050 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 433.950 289.950 436.050 292.050 ;
        RECT 436.950 289.950 439.050 292.050 ;
        RECT 440.550 291.750 445.050 292.050 ;
        RECT 440.550 289.950 446.850 291.750 ;
        RECT 389.550 287.550 394.050 289.050 ;
        RECT 395.100 288.000 396.900 289.800 ;
        RECT 390.000 286.950 394.050 287.550 ;
        RECT 398.400 284.700 399.600 289.800 ;
        RECT 401.100 288.000 402.900 289.800 ;
        RECT 413.100 288.150 414.900 289.950 ;
        RECT 415.950 285.750 417.150 289.950 ;
        RECT 419.100 288.150 420.900 289.950 ;
        RECT 377.400 283.800 381.600 284.700 ;
        RECT 395.400 283.800 399.600 284.700 ;
        RECT 413.400 284.700 417.150 285.750 ;
        RECT 358.800 276.000 360.600 279.600 ;
        RECT 361.800 276.600 363.600 279.600 ;
        RECT 364.800 276.000 366.600 279.600 ;
        RECT 377.400 276.600 379.200 283.800 ;
        RECT 382.500 276.000 384.300 282.600 ;
        RECT 395.400 276.600 397.200 283.800 ;
        RECT 413.400 282.600 414.600 284.700 ;
        RECT 400.500 276.000 402.300 282.600 ;
        RECT 412.800 276.600 414.600 282.600 ;
        RECT 415.800 281.700 423.600 283.050 ;
        RECT 415.800 276.600 417.600 281.700 ;
        RECT 418.800 276.000 420.600 280.800 ;
        RECT 421.800 276.600 423.600 281.700 ;
        RECT 434.400 279.600 435.600 289.950 ;
        RECT 440.550 282.600 441.750 289.950 ;
        RECT 453.150 286.200 454.050 298.800 ;
        RECT 456.150 298.800 457.050 300.900 ;
        RECT 457.950 300.300 465.450 301.500 ;
        RECT 457.950 299.700 459.750 300.300 ;
        RECT 472.050 299.400 473.850 311.400 ;
        RECT 482.400 299.400 484.200 312.000 ;
        RECT 456.150 298.500 464.550 298.800 ;
        RECT 472.950 298.500 473.850 299.400 ;
        RECT 456.150 297.900 473.850 298.500 ;
        RECT 462.750 297.300 473.850 297.900 ;
        RECT 485.400 298.500 487.200 311.400 ;
        RECT 488.400 299.400 490.200 312.000 ;
        RECT 491.400 299.400 493.200 311.400 ;
        RECT 494.400 299.400 496.200 312.000 ;
        RECT 506.400 299.400 508.200 312.000 ;
        RECT 491.400 298.500 492.600 299.400 ;
        RECT 485.400 297.600 492.600 298.500 ;
        RECT 462.750 297.000 464.550 297.300 ;
        RECT 460.950 290.400 463.050 292.050 ;
        RECT 460.950 289.200 468.900 290.400 ;
        RECT 469.950 289.950 472.050 292.050 ;
        RECT 467.100 288.600 468.900 289.200 ;
        RECT 470.100 288.150 471.900 289.950 ;
        RECT 464.100 287.400 465.900 288.000 ;
        RECT 470.100 287.400 471.000 288.150 ;
        RECT 464.100 286.200 471.000 287.400 ;
        RECT 453.150 285.000 465.150 286.200 ;
        RECT 453.150 284.400 454.950 285.000 ;
        RECT 464.100 283.200 465.150 285.000 ;
        RECT 433.800 276.600 435.600 279.600 ;
        RECT 436.800 276.000 438.600 279.600 ;
        RECT 440.550 276.600 442.350 282.600 ;
        RECT 445.950 281.700 448.050 282.600 ;
        RECT 445.950 280.500 449.700 281.700 ;
        RECT 460.350 281.550 462.150 282.300 ;
        RECT 448.650 279.600 449.700 280.500 ;
        RECT 457.200 280.500 462.150 281.550 ;
        RECT 463.650 281.400 465.450 283.200 ;
        RECT 472.950 282.600 473.850 297.300 ;
        RECT 485.100 291.900 486.900 293.700 ;
        RECT 491.400 291.900 492.600 297.600 ;
        RECT 509.400 298.500 511.200 311.400 ;
        RECT 512.400 299.400 514.200 312.000 ;
        RECT 515.400 298.500 517.200 311.400 ;
        RECT 518.400 299.400 520.200 312.000 ;
        RECT 521.400 298.500 523.200 311.400 ;
        RECT 524.400 299.400 526.200 312.000 ;
        RECT 527.400 298.500 529.200 311.400 ;
        RECT 530.400 299.400 532.200 312.000 ;
        RECT 544.800 305.400 546.600 312.000 ;
        RECT 547.800 305.400 549.600 311.400 ;
        RECT 550.800 305.400 552.600 312.000 ;
        RECT 509.400 297.300 513.300 298.500 ;
        RECT 515.400 297.300 519.300 298.500 ;
        RECT 521.400 297.300 525.300 298.500 ;
        RECT 527.400 297.300 530.100 298.500 ;
        RECT 484.950 289.800 487.050 291.900 ;
        RECT 490.950 289.800 493.050 291.900 ;
        RECT 508.950 289.800 511.050 291.900 ;
        RECT 491.400 284.700 492.600 289.800 ;
        RECT 509.100 288.000 510.900 289.800 ;
        RECT 512.100 286.800 513.300 297.300 ;
        RECT 514.500 286.800 516.300 287.400 ;
        RECT 512.100 285.600 516.300 286.800 ;
        RECT 518.100 286.800 519.300 297.300 ;
        RECT 520.500 286.800 522.300 287.400 ;
        RECT 518.100 285.600 522.300 286.800 ;
        RECT 524.100 286.800 525.300 297.300 ;
        RECT 529.200 291.900 530.100 297.300 ;
        RECT 548.400 291.900 549.600 305.400 ;
        RECT 554.550 299.400 556.350 311.400 ;
        RECT 557.550 308.400 559.350 312.000 ;
        RECT 562.050 305.400 563.850 311.400 ;
        RECT 566.250 305.400 568.050 312.000 ;
        RECT 559.950 303.300 563.850 305.400 ;
        RECT 569.850 304.500 571.650 311.400 ;
        RECT 572.850 305.400 574.650 312.000 ;
        RECT 577.650 305.400 579.450 311.400 ;
        RECT 583.050 305.400 584.850 312.000 ;
        RECT 578.250 304.500 579.450 305.400 ;
        RECT 568.950 303.450 575.550 304.500 ;
        RECT 568.950 302.700 570.750 303.450 ;
        RECT 573.750 302.700 575.550 303.450 ;
        RECT 578.250 302.400 583.050 304.500 ;
        RECT 561.150 300.600 563.850 302.400 ;
        RECT 564.750 301.800 566.550 302.400 ;
        RECT 564.750 300.900 571.050 301.800 ;
        RECT 578.250 301.500 579.450 302.400 ;
        RECT 564.750 300.600 566.550 300.900 ;
        RECT 562.950 299.700 563.850 300.600 ;
        RECT 554.550 292.050 555.750 299.400 ;
        RECT 559.950 298.800 562.050 299.700 ;
        RECT 562.950 298.800 568.050 299.700 ;
        RECT 557.850 297.600 562.050 298.800 ;
        RECT 556.950 295.800 558.750 297.600 ;
        RECT 529.200 289.800 532.050 291.900 ;
        RECT 544.950 289.800 547.050 291.900 ;
        RECT 547.950 289.800 550.050 291.900 ;
        RECT 550.950 289.800 553.050 291.900 ;
        RECT 554.550 291.750 559.050 292.050 ;
        RECT 554.550 289.950 560.850 291.750 ;
        RECT 526.500 286.800 528.300 287.400 ;
        RECT 524.100 285.600 528.300 286.800 ;
        RECT 512.100 284.700 513.300 285.600 ;
        RECT 518.100 284.700 519.300 285.600 ;
        RECT 524.100 284.700 525.300 285.600 ;
        RECT 529.200 284.700 530.100 289.800 ;
        RECT 545.100 288.000 546.900 289.800 ;
        RECT 548.400 284.700 549.600 289.800 ;
        RECT 551.100 288.000 552.900 289.800 ;
        RECT 485.400 283.500 492.600 284.700 ;
        RECT 485.400 282.600 486.600 283.500 ;
        RECT 491.400 282.600 492.600 283.500 ;
        RECT 509.400 283.500 513.300 284.700 ;
        RECT 515.400 283.500 519.300 284.700 ;
        RECT 521.400 283.500 525.300 284.700 ;
        RECT 527.400 283.500 530.100 284.700 ;
        RECT 545.400 283.800 549.600 284.700 ;
        RECT 466.950 280.500 469.050 282.600 ;
        RECT 457.200 279.600 458.250 280.500 ;
        RECT 466.950 279.600 468.000 280.500 ;
        RECT 443.850 276.000 445.650 279.600 ;
        RECT 448.650 276.600 450.450 279.600 ;
        RECT 452.850 276.000 454.650 279.600 ;
        RECT 456.450 276.600 458.250 279.600 ;
        RECT 459.750 276.000 461.550 279.600 ;
        RECT 464.250 278.700 468.000 279.600 ;
        RECT 464.250 276.600 466.050 278.700 ;
        RECT 469.050 276.000 470.850 279.600 ;
        RECT 472.050 276.600 473.850 282.600 ;
        RECT 482.400 276.000 484.200 282.600 ;
        RECT 485.400 276.600 487.200 282.600 ;
        RECT 488.400 276.000 490.200 282.600 ;
        RECT 491.400 276.600 493.200 282.600 ;
        RECT 494.400 276.000 496.200 282.600 ;
        RECT 506.400 276.000 508.200 282.600 ;
        RECT 509.400 276.600 511.200 283.500 ;
        RECT 512.400 276.000 514.200 282.600 ;
        RECT 515.400 276.600 517.200 283.500 ;
        RECT 518.400 276.000 520.200 282.600 ;
        RECT 521.400 276.600 523.200 283.500 ;
        RECT 524.400 276.000 526.200 282.600 ;
        RECT 527.400 276.600 529.200 283.500 ;
        RECT 530.400 276.000 532.200 282.600 ;
        RECT 545.400 276.600 547.200 283.800 ;
        RECT 554.550 282.600 555.750 289.950 ;
        RECT 567.150 286.200 568.050 298.800 ;
        RECT 570.150 298.800 571.050 300.900 ;
        RECT 571.950 300.300 579.450 301.500 ;
        RECT 571.950 299.700 573.750 300.300 ;
        RECT 586.050 299.400 587.850 311.400 ;
        RECT 599.400 305.400 601.200 312.000 ;
        RECT 602.400 305.400 604.200 311.400 ;
        RECT 570.150 298.500 578.550 298.800 ;
        RECT 586.950 298.500 587.850 299.400 ;
        RECT 570.150 297.900 587.850 298.500 ;
        RECT 576.750 297.300 587.850 297.900 ;
        RECT 576.750 297.000 578.550 297.300 ;
        RECT 574.950 290.400 577.050 292.050 ;
        RECT 574.950 289.200 582.900 290.400 ;
        RECT 583.950 289.950 586.050 292.050 ;
        RECT 581.100 288.600 582.900 289.200 ;
        RECT 584.100 288.150 585.900 289.950 ;
        RECT 578.100 287.400 579.900 288.000 ;
        RECT 584.100 287.400 585.000 288.150 ;
        RECT 578.100 286.200 585.000 287.400 ;
        RECT 567.150 285.000 579.150 286.200 ;
        RECT 567.150 284.400 568.950 285.000 ;
        RECT 578.100 283.200 579.150 285.000 ;
        RECT 550.500 276.000 552.300 282.600 ;
        RECT 554.550 276.600 556.350 282.600 ;
        RECT 559.950 281.700 562.050 282.600 ;
        RECT 559.950 280.500 563.700 281.700 ;
        RECT 574.350 281.550 576.150 282.300 ;
        RECT 562.650 279.600 563.700 280.500 ;
        RECT 571.200 280.500 576.150 281.550 ;
        RECT 577.650 281.400 579.450 283.200 ;
        RECT 586.950 282.600 587.850 297.300 ;
        RECT 602.850 292.050 604.050 305.400 ;
        RECT 607.500 299.400 609.300 312.000 ;
        RECT 619.800 299.400 621.600 311.400 ;
        RECT 622.800 305.400 624.600 312.000 ;
        RECT 625.800 305.400 627.600 311.400 ;
        RECT 608.100 292.050 609.900 293.850 ;
        RECT 619.800 292.050 621.000 299.400 ;
        RECT 626.400 298.500 627.600 305.400 ;
        RECT 621.900 297.600 627.600 298.500 ;
        RECT 630.150 299.400 631.950 311.400 ;
        RECT 633.150 305.400 634.950 312.000 ;
        RECT 638.550 305.400 640.350 311.400 ;
        RECT 643.350 305.400 645.150 312.000 ;
        RECT 638.550 304.500 639.750 305.400 ;
        RECT 646.350 304.500 648.150 311.400 ;
        RECT 649.950 305.400 651.750 312.000 ;
        RECT 654.150 305.400 655.950 311.400 ;
        RECT 658.650 308.400 660.450 312.000 ;
        RECT 634.950 302.400 639.750 304.500 ;
        RECT 642.450 303.450 649.050 304.500 ;
        RECT 642.450 302.700 644.250 303.450 ;
        RECT 647.250 302.700 649.050 303.450 ;
        RECT 654.150 303.300 658.050 305.400 ;
        RECT 638.550 301.500 639.750 302.400 ;
        RECT 651.450 301.800 653.250 302.400 ;
        RECT 638.550 300.300 646.050 301.500 ;
        RECT 644.250 299.700 646.050 300.300 ;
        RECT 646.950 300.900 653.250 301.800 ;
        RECT 630.150 298.500 631.050 299.400 ;
        RECT 646.950 298.800 647.850 300.900 ;
        RECT 651.450 300.600 653.250 300.900 ;
        RECT 654.150 300.600 656.850 302.400 ;
        RECT 654.150 299.700 655.050 300.600 ;
        RECT 639.450 298.500 647.850 298.800 ;
        RECT 630.150 297.900 647.850 298.500 ;
        RECT 649.950 298.800 655.050 299.700 ;
        RECT 655.950 298.800 658.050 299.700 ;
        RECT 661.650 299.400 663.450 311.400 ;
        RECT 673.800 300.600 675.600 311.400 ;
        RECT 681.300 310.050 683.100 311.400 ;
        RECT 679.950 307.950 683.100 310.050 ;
        RECT 673.800 299.400 678.600 300.600 ;
        RECT 621.900 296.700 623.850 297.600 ;
        RECT 598.950 289.950 601.050 292.050 ;
        RECT 601.950 289.950 604.050 292.050 ;
        RECT 604.950 289.950 607.050 292.050 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 619.800 289.950 622.050 292.050 ;
        RECT 599.100 288.150 600.900 289.950 ;
        RECT 601.950 285.750 603.150 289.950 ;
        RECT 605.100 288.150 606.900 289.950 ;
        RECT 599.400 284.700 603.150 285.750 ;
        RECT 599.400 282.600 600.600 284.700 ;
        RECT 580.950 280.500 583.050 282.600 ;
        RECT 571.200 279.600 572.250 280.500 ;
        RECT 580.950 279.600 582.000 280.500 ;
        RECT 557.850 276.000 559.650 279.600 ;
        RECT 562.650 276.600 564.450 279.600 ;
        RECT 566.850 276.000 568.650 279.600 ;
        RECT 570.450 276.600 572.250 279.600 ;
        RECT 573.750 276.000 575.550 279.600 ;
        RECT 578.250 278.700 582.000 279.600 ;
        RECT 578.250 276.600 580.050 278.700 ;
        RECT 583.050 276.000 584.850 279.600 ;
        RECT 586.050 276.600 587.850 282.600 ;
        RECT 598.800 276.600 600.600 282.600 ;
        RECT 601.800 281.700 609.600 283.050 ;
        RECT 601.800 276.600 603.600 281.700 ;
        RECT 604.800 276.000 606.600 280.800 ;
        RECT 607.800 276.600 609.600 281.700 ;
        RECT 619.800 282.600 621.000 289.950 ;
        RECT 622.950 285.300 623.850 296.700 ;
        RECT 630.150 297.300 641.250 297.900 ;
        RECT 626.100 292.050 627.900 293.850 ;
        RECT 625.950 289.950 628.050 292.050 ;
        RECT 621.900 284.400 623.850 285.300 ;
        RECT 621.900 283.500 627.600 284.400 ;
        RECT 619.800 276.600 621.600 282.600 ;
        RECT 626.400 279.600 627.600 283.500 ;
        RECT 622.800 276.000 624.600 279.600 ;
        RECT 625.800 276.600 627.600 279.600 ;
        RECT 630.150 282.600 631.050 297.300 ;
        RECT 639.450 297.000 641.250 297.300 ;
        RECT 631.950 289.950 634.050 292.050 ;
        RECT 640.950 290.400 643.050 292.050 ;
        RECT 632.100 288.150 633.900 289.950 ;
        RECT 635.100 289.200 643.050 290.400 ;
        RECT 635.100 288.600 636.900 289.200 ;
        RECT 633.000 287.400 633.900 288.150 ;
        RECT 638.100 287.400 639.900 288.000 ;
        RECT 633.000 286.200 639.900 287.400 ;
        RECT 649.950 286.200 650.850 298.800 ;
        RECT 655.950 297.600 660.150 298.800 ;
        RECT 659.250 295.800 661.050 297.600 ;
        RECT 662.250 292.050 663.450 299.400 ;
        RECT 676.500 298.500 678.600 299.400 ;
        RECT 681.300 299.400 683.100 307.950 ;
        RECT 688.800 300.300 690.600 311.400 ;
        RECT 698.400 305.400 700.200 312.000 ;
        RECT 701.400 305.400 703.200 311.400 ;
        RECT 686.100 299.400 690.600 300.300 ;
        RECT 681.300 297.900 682.500 299.400 ;
        RECT 681.000 297.000 682.500 297.900 ;
        RECT 686.100 297.300 688.200 299.400 ;
        RECT 670.950 294.450 675.000 295.050 ;
        RECT 681.000 294.900 681.900 297.000 ;
        RECT 682.950 295.500 685.050 295.800 ;
        RECT 670.950 293.700 675.450 294.450 ;
        RECT 670.950 292.950 675.900 293.700 ;
        RECT 658.950 291.750 663.450 292.050 ;
        RECT 674.100 291.900 675.900 292.950 ;
        RECT 679.950 292.800 682.050 294.900 ;
        RECT 682.950 293.700 686.700 295.500 ;
        RECT 680.400 291.900 682.800 292.800 ;
        RECT 657.150 289.950 663.450 291.750 ;
        RECT 638.850 285.000 650.850 286.200 ;
        RECT 638.850 283.200 639.900 285.000 ;
        RECT 649.050 284.400 650.850 285.000 ;
        RECT 630.150 276.600 631.950 282.600 ;
        RECT 634.950 280.500 637.050 282.600 ;
        RECT 638.550 281.400 640.350 283.200 ;
        RECT 662.250 282.600 663.450 289.950 ;
        RECT 673.950 289.800 676.050 291.900 ;
        RECT 678.600 289.200 680.400 291.000 ;
        RECT 678.750 287.100 680.850 289.200 ;
        RECT 681.750 286.200 682.800 291.900 ;
        RECT 683.700 291.900 685.500 292.500 ;
        RECT 698.100 292.050 699.900 293.850 ;
        RECT 701.400 292.050 702.600 305.400 ;
        RECT 713.700 299.400 715.500 312.000 ;
        RECT 718.800 305.400 720.600 311.400 ;
        RECT 721.800 305.400 723.600 312.000 ;
        RECT 703.950 294.450 708.000 295.050 ;
        RECT 703.950 292.950 708.450 294.450 ;
        RECT 683.700 290.700 691.050 291.900 ;
        RECT 688.950 289.800 691.050 290.700 ;
        RECT 697.950 289.950 700.050 292.050 ;
        RECT 700.950 289.950 703.050 292.050 ;
        RECT 676.500 283.500 678.600 284.700 ;
        RECT 679.950 284.100 682.800 286.200 ;
        RECT 683.700 287.400 685.500 289.200 ;
        RECT 688.950 288.000 690.750 289.800 ;
        RECT 683.700 285.300 685.800 287.400 ;
        RECT 683.700 284.400 690.000 285.300 ;
        RECT 641.850 281.550 643.650 282.300 ;
        RECT 655.950 281.700 658.050 282.600 ;
        RECT 641.850 280.500 646.800 281.550 ;
        RECT 636.000 279.600 637.050 280.500 ;
        RECT 645.750 279.600 646.800 280.500 ;
        RECT 654.300 280.500 658.050 281.700 ;
        RECT 654.300 279.600 655.350 280.500 ;
        RECT 633.150 276.000 634.950 279.600 ;
        RECT 636.000 278.700 639.750 279.600 ;
        RECT 637.950 276.600 639.750 278.700 ;
        RECT 642.450 276.000 644.250 279.600 ;
        RECT 645.750 276.600 647.550 279.600 ;
        RECT 649.350 276.000 651.150 279.600 ;
        RECT 653.550 276.600 655.350 279.600 ;
        RECT 658.350 276.000 660.150 279.600 ;
        RECT 661.650 276.600 663.450 282.600 ;
        RECT 673.800 282.600 678.600 283.500 ;
        RECT 681.600 282.600 682.800 284.100 ;
        RECT 688.800 282.600 690.000 284.400 ;
        RECT 673.800 276.600 675.600 282.600 ;
        RECT 681.300 276.600 683.100 282.600 ;
        RECT 688.800 276.600 690.600 282.600 ;
        RECT 701.400 279.600 702.600 289.950 ;
        RECT 707.550 289.050 708.450 292.950 ;
        RECT 713.100 292.050 714.900 293.850 ;
        RECT 718.950 292.050 720.150 305.400 ;
        RECT 737.700 300.600 739.500 311.400 ;
        RECT 737.700 299.400 741.300 300.600 ;
        RECT 742.800 299.400 744.600 312.000 ;
        RECT 752.400 300.300 754.200 311.400 ;
        RECT 755.400 301.200 757.200 312.000 ;
        RECT 758.400 300.300 760.200 311.400 ;
        RECT 752.400 299.400 760.200 300.300 ;
        RECT 761.400 299.400 763.200 311.400 ;
        RECT 776.700 300.600 778.500 311.400 ;
        RECT 776.700 299.400 780.300 300.600 ;
        RECT 781.800 299.400 783.600 312.000 ;
        RECT 791.400 305.400 793.200 312.000 ;
        RECT 794.400 305.400 796.200 311.400 ;
        RECT 797.400 305.400 799.200 312.000 ;
        RECT 737.100 292.050 738.900 293.850 ;
        RECT 740.400 292.050 741.300 299.400 ;
        RECT 743.100 292.050 744.900 293.850 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 715.950 289.950 718.050 292.050 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 755.100 291.900 756.900 293.700 ;
        RECT 761.700 291.900 762.600 299.400 ;
        RECT 776.100 292.050 777.900 293.850 ;
        RECT 779.400 292.050 780.300 299.400 ;
        RECT 782.100 292.050 783.900 293.850 ;
        RECT 707.550 287.550 712.050 289.050 ;
        RECT 716.100 288.150 717.900 289.950 ;
        RECT 708.000 286.950 712.050 287.550 ;
        RECT 719.850 285.750 721.050 289.950 ;
        RECT 722.100 288.150 723.900 289.950 ;
        RECT 719.850 284.700 723.600 285.750 ;
        RECT 713.400 281.700 721.200 283.050 ;
        RECT 698.400 276.000 700.200 279.600 ;
        RECT 701.400 276.600 703.200 279.600 ;
        RECT 713.400 276.600 715.200 281.700 ;
        RECT 716.400 276.000 718.200 280.800 ;
        RECT 719.400 276.600 721.200 281.700 ;
        RECT 722.400 282.600 723.600 284.700 ;
        RECT 722.400 276.600 724.200 282.600 ;
        RECT 740.400 279.600 741.300 289.950 ;
        RECT 751.950 289.800 754.050 291.900 ;
        RECT 754.950 289.800 757.050 291.900 ;
        RECT 757.950 289.800 760.050 291.900 ;
        RECT 760.950 289.800 763.050 291.900 ;
        RECT 775.950 289.950 778.050 292.050 ;
        RECT 778.950 289.950 781.050 292.050 ;
        RECT 781.950 289.950 784.050 292.050 ;
        RECT 794.400 291.900 795.600 305.400 ;
        RECT 809.700 299.400 811.500 312.000 ;
        RECT 814.800 305.400 816.600 311.400 ;
        RECT 817.800 305.400 819.600 312.000 ;
        RECT 833.400 305.400 835.200 312.000 ;
        RECT 836.400 305.400 838.200 311.400 ;
        RECT 799.950 294.450 804.000 295.050 ;
        RECT 799.950 292.950 804.450 294.450 ;
        RECT 752.100 288.000 753.900 289.800 ;
        RECT 758.100 288.000 759.900 289.800 ;
        RECT 761.700 282.600 762.600 289.800 ;
        RECT 736.800 276.000 738.600 279.600 ;
        RECT 739.800 276.600 741.600 279.600 ;
        RECT 742.800 276.000 744.600 279.600 ;
        RECT 753.000 276.000 754.800 282.600 ;
        RECT 757.500 281.400 762.600 282.600 ;
        RECT 757.500 276.600 759.300 281.400 ;
        RECT 779.400 279.600 780.300 289.950 ;
        RECT 790.950 289.800 793.050 291.900 ;
        RECT 793.950 289.800 796.050 291.900 ;
        RECT 796.950 289.800 799.050 291.900 ;
        RECT 791.100 288.000 792.900 289.800 ;
        RECT 794.400 284.700 795.600 289.800 ;
        RECT 797.100 288.000 798.900 289.800 ;
        RECT 803.550 289.050 804.450 292.950 ;
        RECT 809.100 292.050 810.900 293.850 ;
        RECT 814.950 292.050 816.150 305.400 ;
        RECT 836.850 292.050 838.050 305.400 ;
        RECT 841.500 299.400 843.300 312.000 ;
        RECT 842.100 292.050 843.900 293.850 ;
        RECT 808.950 289.950 811.050 292.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 814.950 289.950 817.050 292.050 ;
        RECT 817.950 289.950 820.050 292.050 ;
        RECT 832.950 289.950 835.050 292.050 ;
        RECT 835.950 289.950 838.050 292.050 ;
        RECT 838.950 289.950 841.050 292.050 ;
        RECT 841.950 289.950 844.050 292.050 ;
        RECT 803.550 287.550 808.050 289.050 ;
        RECT 812.100 288.150 813.900 289.950 ;
        RECT 804.000 286.950 808.050 287.550 ;
        RECT 815.850 285.750 817.050 289.950 ;
        RECT 818.100 288.150 819.900 289.950 ;
        RECT 833.100 288.150 834.900 289.950 ;
        RECT 835.950 285.750 837.150 289.950 ;
        RECT 839.100 288.150 840.900 289.950 ;
        RECT 815.850 284.700 819.600 285.750 ;
        RECT 794.400 283.800 798.600 284.700 ;
        RECT 760.500 276.000 762.300 279.600 ;
        RECT 775.800 276.000 777.600 279.600 ;
        RECT 778.800 276.600 780.600 279.600 ;
        RECT 781.800 276.000 783.600 279.600 ;
        RECT 791.700 276.000 793.500 282.600 ;
        RECT 796.800 276.600 798.600 283.800 ;
        RECT 809.400 281.700 817.200 283.050 ;
        RECT 809.400 276.600 811.200 281.700 ;
        RECT 812.400 276.000 814.200 280.800 ;
        RECT 815.400 276.600 817.200 281.700 ;
        RECT 818.400 282.600 819.600 284.700 ;
        RECT 833.400 284.700 837.150 285.750 ;
        RECT 833.400 282.600 834.600 284.700 ;
        RECT 818.400 276.600 820.200 282.600 ;
        RECT 832.800 276.600 834.600 282.600 ;
        RECT 835.800 281.700 843.600 283.050 ;
        RECT 835.800 276.600 837.600 281.700 ;
        RECT 838.800 276.000 840.600 280.800 ;
        RECT 841.800 276.600 843.600 281.700 ;
        RECT 2.550 266.400 4.350 272.400 ;
        RECT 5.850 269.400 7.650 273.000 ;
        RECT 10.650 269.400 12.450 272.400 ;
        RECT 14.850 269.400 16.650 273.000 ;
        RECT 18.450 269.400 20.250 272.400 ;
        RECT 21.750 269.400 23.550 273.000 ;
        RECT 26.250 270.300 28.050 272.400 ;
        RECT 26.250 269.400 30.000 270.300 ;
        RECT 31.050 269.400 32.850 273.000 ;
        RECT 10.650 268.500 11.700 269.400 ;
        RECT 7.950 267.300 11.700 268.500 ;
        RECT 19.200 268.500 20.250 269.400 ;
        RECT 28.950 268.500 30.000 269.400 ;
        RECT 19.200 267.450 24.150 268.500 ;
        RECT 7.950 266.400 10.050 267.300 ;
        RECT 22.350 266.700 24.150 267.450 ;
        RECT 2.550 259.050 3.750 266.400 ;
        RECT 25.650 265.800 27.450 267.600 ;
        RECT 28.950 266.400 31.050 268.500 ;
        RECT 34.050 266.400 35.850 272.400 ;
        RECT 15.150 264.000 16.950 264.600 ;
        RECT 26.100 264.000 27.150 265.800 ;
        RECT 15.150 262.800 27.150 264.000 ;
        RECT 2.550 257.250 8.850 259.050 ;
        RECT 2.550 256.950 7.050 257.250 ;
        RECT 2.550 249.600 3.750 256.950 ;
        RECT 4.950 251.400 6.750 253.200 ;
        RECT 5.850 250.200 10.050 251.400 ;
        RECT 15.150 250.200 16.050 262.800 ;
        RECT 26.100 261.600 33.000 262.800 ;
        RECT 26.100 261.000 27.900 261.600 ;
        RECT 32.100 260.850 33.000 261.600 ;
        RECT 29.100 259.800 30.900 260.400 ;
        RECT 22.950 258.600 30.900 259.800 ;
        RECT 32.100 259.050 33.900 260.850 ;
        RECT 22.950 256.950 25.050 258.600 ;
        RECT 31.950 256.950 34.050 259.050 ;
        RECT 24.750 251.700 26.550 252.000 ;
        RECT 34.950 251.700 35.850 266.400 ;
        RECT 24.750 251.100 35.850 251.700 ;
        RECT 2.550 237.600 4.350 249.600 ;
        RECT 7.950 249.300 10.050 250.200 ;
        RECT 10.950 249.300 16.050 250.200 ;
        RECT 18.150 250.500 35.850 251.100 ;
        RECT 18.150 250.200 26.550 250.500 ;
        RECT 10.950 248.400 11.850 249.300 ;
        RECT 9.150 246.600 11.850 248.400 ;
        RECT 12.750 248.100 14.550 248.400 ;
        RECT 18.150 248.100 19.050 250.200 ;
        RECT 34.950 249.600 35.850 250.500 ;
        RECT 12.750 247.200 19.050 248.100 ;
        RECT 19.950 248.700 21.750 249.300 ;
        RECT 19.950 247.500 27.450 248.700 ;
        RECT 12.750 246.600 14.550 247.200 ;
        RECT 26.250 246.600 27.450 247.500 ;
        RECT 7.950 243.600 11.850 245.700 ;
        RECT 16.950 245.550 18.750 246.300 ;
        RECT 21.750 245.550 23.550 246.300 ;
        RECT 16.950 244.500 23.550 245.550 ;
        RECT 26.250 244.500 31.050 246.600 ;
        RECT 5.550 237.000 7.350 240.600 ;
        RECT 10.050 237.600 11.850 243.600 ;
        RECT 14.250 237.000 16.050 243.600 ;
        RECT 17.850 237.600 19.650 244.500 ;
        RECT 26.250 243.600 27.450 244.500 ;
        RECT 20.850 237.000 22.650 243.600 ;
        RECT 25.650 237.600 27.450 243.600 ;
        RECT 31.050 237.000 32.850 243.600 ;
        RECT 34.050 237.600 35.850 249.600 ;
        RECT 39.150 266.400 40.950 272.400 ;
        RECT 42.150 269.400 43.950 273.000 ;
        RECT 46.950 270.300 48.750 272.400 ;
        RECT 45.000 269.400 48.750 270.300 ;
        RECT 51.450 269.400 53.250 273.000 ;
        RECT 54.750 269.400 56.550 272.400 ;
        RECT 58.350 269.400 60.150 273.000 ;
        RECT 62.550 269.400 64.350 272.400 ;
        RECT 67.350 269.400 69.150 273.000 ;
        RECT 45.000 268.500 46.050 269.400 ;
        RECT 54.750 268.500 55.800 269.400 ;
        RECT 43.950 266.400 46.050 268.500 ;
        RECT 39.150 251.700 40.050 266.400 ;
        RECT 47.550 265.800 49.350 267.600 ;
        RECT 50.850 267.450 55.800 268.500 ;
        RECT 63.300 268.500 64.350 269.400 ;
        RECT 50.850 266.700 52.650 267.450 ;
        RECT 63.300 267.300 67.050 268.500 ;
        RECT 64.950 266.400 67.050 267.300 ;
        RECT 70.650 266.400 72.450 272.400 ;
        RECT 80.700 266.400 82.500 273.000 ;
        RECT 47.850 264.000 48.900 265.800 ;
        RECT 58.050 264.000 59.850 264.600 ;
        RECT 47.850 262.800 59.850 264.000 ;
        RECT 42.000 261.600 48.900 262.800 ;
        RECT 42.000 260.850 42.900 261.600 ;
        RECT 47.100 261.000 48.900 261.600 ;
        RECT 41.100 259.050 42.900 260.850 ;
        RECT 44.100 259.800 45.900 260.400 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 44.100 258.600 52.050 259.800 ;
        RECT 49.950 256.950 52.050 258.600 ;
        RECT 48.450 251.700 50.250 252.000 ;
        RECT 39.150 251.100 50.250 251.700 ;
        RECT 39.150 250.500 56.850 251.100 ;
        RECT 39.150 249.600 40.050 250.500 ;
        RECT 48.450 250.200 56.850 250.500 ;
        RECT 39.150 237.600 40.950 249.600 ;
        RECT 53.250 248.700 55.050 249.300 ;
        RECT 47.550 247.500 55.050 248.700 ;
        RECT 55.950 248.100 56.850 250.200 ;
        RECT 58.950 250.200 59.850 262.800 ;
        RECT 71.250 259.050 72.450 266.400 ;
        RECT 85.800 265.200 87.600 272.400 ;
        RECT 100.800 266.400 102.600 272.400 ;
        RECT 83.400 264.300 87.600 265.200 ;
        RECT 101.400 264.300 102.600 266.400 ;
        RECT 103.800 267.300 105.600 272.400 ;
        RECT 106.800 268.200 108.600 273.000 ;
        RECT 109.800 267.300 111.600 272.400 ;
        RECT 103.800 265.950 111.600 267.300 ;
        RECT 121.800 266.400 123.600 273.000 ;
        RECT 124.800 265.500 126.600 272.400 ;
        RECT 127.800 266.400 129.600 273.000 ;
        RECT 130.800 265.500 132.600 272.400 ;
        RECT 133.800 266.400 135.600 273.000 ;
        RECT 136.800 265.500 138.600 272.400 ;
        RECT 139.800 266.400 141.600 273.000 ;
        RECT 142.800 265.500 144.600 272.400 ;
        RECT 145.800 266.400 147.600 273.000 ;
        RECT 123.900 264.300 126.600 265.500 ;
        RECT 128.700 264.300 132.600 265.500 ;
        RECT 134.700 264.300 138.600 265.500 ;
        RECT 140.700 264.300 144.600 265.500 ;
        RECT 158.400 265.200 160.200 272.400 ;
        RECT 163.500 266.400 165.300 273.000 ;
        RECT 173.400 269.400 175.200 273.000 ;
        RECT 176.400 269.400 178.200 272.400 ;
        RECT 179.400 269.400 181.200 273.000 ;
        RECT 191.400 269.400 193.200 273.000 ;
        RECT 194.400 269.400 196.200 272.400 ;
        RECT 197.400 269.400 199.200 273.000 ;
        RECT 158.400 264.300 162.600 265.200 ;
        RECT 80.100 259.200 81.900 261.000 ;
        RECT 83.400 259.200 84.600 264.300 ;
        RECT 101.400 263.250 105.150 264.300 ;
        RECT 88.950 261.450 91.050 262.050 ;
        RECT 86.100 259.200 87.900 261.000 ;
        RECT 88.950 260.550 96.450 261.450 ;
        RECT 88.950 259.950 91.050 260.550 ;
        RECT 66.150 257.250 72.450 259.050 ;
        RECT 67.950 256.950 72.450 257.250 ;
        RECT 79.950 257.100 82.050 259.200 ;
        RECT 82.950 257.100 85.050 259.200 ;
        RECT 85.950 257.100 88.050 259.200 ;
        RECT 68.250 251.400 70.050 253.200 ;
        RECT 64.950 250.200 69.150 251.400 ;
        RECT 58.950 249.300 64.050 250.200 ;
        RECT 64.950 249.300 67.050 250.200 ;
        RECT 71.250 249.600 72.450 256.950 ;
        RECT 63.150 248.400 64.050 249.300 ;
        RECT 60.450 248.100 62.250 248.400 ;
        RECT 47.550 246.600 48.750 247.500 ;
        RECT 55.950 247.200 62.250 248.100 ;
        RECT 60.450 246.600 62.250 247.200 ;
        RECT 63.150 246.600 65.850 248.400 ;
        RECT 43.950 244.500 48.750 246.600 ;
        RECT 51.450 245.550 53.250 246.300 ;
        RECT 56.250 245.550 58.050 246.300 ;
        RECT 51.450 244.500 58.050 245.550 ;
        RECT 47.550 243.600 48.750 244.500 ;
        RECT 42.150 237.000 43.950 243.600 ;
        RECT 47.550 237.600 49.350 243.600 ;
        RECT 52.350 237.000 54.150 243.600 ;
        RECT 55.350 237.600 57.150 244.500 ;
        RECT 63.150 243.600 67.050 245.700 ;
        RECT 58.950 237.000 60.750 243.600 ;
        RECT 63.150 237.600 64.950 243.600 ;
        RECT 67.650 237.000 69.450 240.600 ;
        RECT 70.650 237.600 72.450 249.600 ;
        RECT 83.400 243.600 84.600 257.100 ;
        RECT 95.550 256.050 96.450 260.550 ;
        RECT 101.100 259.050 102.900 260.850 ;
        RECT 103.950 259.050 105.150 263.250 ;
        RECT 107.100 259.050 108.900 260.850 ;
        RECT 123.900 259.200 124.800 264.300 ;
        RECT 128.700 263.400 129.900 264.300 ;
        RECT 134.700 263.400 135.900 264.300 ;
        RECT 140.700 263.400 141.900 264.300 ;
        RECT 125.700 262.200 129.900 263.400 ;
        RECT 125.700 261.600 127.500 262.200 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 121.950 257.100 124.800 259.200 ;
        RECT 95.550 254.550 100.050 256.050 ;
        RECT 96.000 253.950 100.050 254.550 ;
        RECT 104.850 243.600 106.050 256.950 ;
        RECT 110.100 255.150 111.900 256.950 ;
        RECT 123.900 251.700 124.800 257.100 ;
        RECT 128.700 251.700 129.900 262.200 ;
        RECT 131.700 262.200 135.900 263.400 ;
        RECT 131.700 261.600 133.500 262.200 ;
        RECT 134.700 251.700 135.900 262.200 ;
        RECT 137.700 262.200 141.900 263.400 ;
        RECT 137.700 261.600 139.500 262.200 ;
        RECT 140.700 251.700 141.900 262.200 ;
        RECT 143.100 259.200 144.900 261.000 ;
        RECT 158.100 259.200 159.900 261.000 ;
        RECT 161.400 259.200 162.600 264.300 ;
        RECT 164.100 259.200 165.900 261.000 ;
        RECT 142.950 257.100 145.050 259.200 ;
        RECT 157.950 257.100 160.050 259.200 ;
        RECT 160.950 257.100 163.050 259.200 ;
        RECT 163.950 257.100 166.050 259.200 ;
        RECT 176.700 259.050 177.600 269.400 ;
        RECT 194.700 259.050 195.600 269.400 ;
        RECT 203.550 266.400 205.350 272.400 ;
        RECT 206.850 269.400 208.650 273.000 ;
        RECT 211.650 269.400 213.450 272.400 ;
        RECT 215.850 269.400 217.650 273.000 ;
        RECT 219.450 269.400 221.250 272.400 ;
        RECT 222.750 269.400 224.550 273.000 ;
        RECT 227.250 270.300 229.050 272.400 ;
        RECT 227.250 269.400 231.000 270.300 ;
        RECT 232.050 269.400 233.850 273.000 ;
        RECT 211.650 268.500 212.700 269.400 ;
        RECT 208.950 267.300 212.700 268.500 ;
        RECT 220.200 268.500 221.250 269.400 ;
        RECT 229.950 268.500 231.000 269.400 ;
        RECT 220.200 267.450 225.150 268.500 ;
        RECT 208.950 266.400 211.050 267.300 ;
        RECT 223.350 266.700 225.150 267.450 ;
        RECT 203.550 259.050 204.750 266.400 ;
        RECT 226.650 265.800 228.450 267.600 ;
        RECT 229.950 266.400 232.050 268.500 ;
        RECT 235.050 266.400 236.850 272.400 ;
        RECT 245.400 269.400 247.200 273.000 ;
        RECT 248.400 269.400 250.200 272.400 ;
        RECT 216.150 264.000 217.950 264.600 ;
        RECT 227.100 264.000 228.150 265.800 ;
        RECT 216.150 262.800 228.150 264.000 ;
        RECT 123.900 250.500 126.600 251.700 ;
        RECT 128.700 250.500 132.600 251.700 ;
        RECT 134.700 250.500 138.600 251.700 ;
        RECT 140.700 250.500 144.600 251.700 ;
        RECT 80.400 237.000 82.200 243.600 ;
        RECT 83.400 237.600 85.200 243.600 ;
        RECT 86.400 237.000 88.200 243.600 ;
        RECT 101.400 237.000 103.200 243.600 ;
        RECT 104.400 237.600 106.200 243.600 ;
        RECT 109.500 237.000 111.300 249.600 ;
        RECT 121.800 237.000 123.600 249.600 ;
        RECT 124.800 237.600 126.600 250.500 ;
        RECT 127.800 237.000 129.600 249.600 ;
        RECT 130.800 237.600 132.600 250.500 ;
        RECT 133.800 237.000 135.600 249.600 ;
        RECT 136.800 237.600 138.600 250.500 ;
        RECT 139.800 237.000 141.600 249.600 ;
        RECT 142.800 237.600 144.600 250.500 ;
        RECT 145.800 237.000 147.600 249.600 ;
        RECT 161.400 243.600 162.600 257.100 ;
        RECT 172.950 256.950 175.050 259.050 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 178.950 256.950 181.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 196.950 256.950 199.050 259.050 ;
        RECT 203.550 257.250 209.850 259.050 ;
        RECT 203.550 256.950 208.050 257.250 ;
        RECT 173.100 255.150 174.900 256.950 ;
        RECT 176.700 249.600 177.600 256.950 ;
        RECT 179.100 255.150 180.900 256.950 ;
        RECT 191.100 255.150 192.900 256.950 ;
        RECT 194.700 249.600 195.600 256.950 ;
        RECT 197.100 255.150 198.900 256.950 ;
        RECT 203.550 249.600 204.750 256.950 ;
        RECT 205.950 251.400 207.750 253.200 ;
        RECT 206.850 250.200 211.050 251.400 ;
        RECT 216.150 250.200 217.050 262.800 ;
        RECT 227.100 261.600 234.000 262.800 ;
        RECT 227.100 261.000 228.900 261.600 ;
        RECT 233.100 260.850 234.000 261.600 ;
        RECT 230.100 259.800 231.900 260.400 ;
        RECT 223.950 258.600 231.900 259.800 ;
        RECT 233.100 259.050 234.900 260.850 ;
        RECT 223.950 256.950 226.050 258.600 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 225.750 251.700 227.550 252.000 ;
        RECT 235.950 251.700 236.850 266.400 ;
        RECT 248.400 259.050 249.600 269.400 ;
        RECT 260.400 264.600 262.200 272.400 ;
        RECT 264.900 266.400 266.700 273.000 ;
        RECT 267.900 268.200 269.700 272.400 ;
        RECT 267.900 266.400 270.600 268.200 ;
        RECT 283.800 266.400 285.600 272.400 ;
        RECT 266.100 264.600 267.900 265.500 ;
        RECT 260.400 263.700 267.900 264.600 ;
        RECT 260.100 259.200 261.900 261.000 ;
        RECT 244.950 256.950 247.050 259.050 ;
        RECT 247.950 256.950 250.050 259.050 ;
        RECT 259.950 257.100 262.050 259.200 ;
        RECT 245.100 255.150 246.900 256.950 ;
        RECT 225.750 251.100 236.850 251.700 ;
        RECT 157.800 237.000 159.600 243.600 ;
        RECT 160.800 237.600 162.600 243.600 ;
        RECT 163.800 237.000 165.600 243.600 ;
        RECT 173.400 237.000 175.200 249.600 ;
        RECT 176.700 248.400 180.300 249.600 ;
        RECT 178.500 237.600 180.300 248.400 ;
        RECT 191.400 237.000 193.200 249.600 ;
        RECT 194.700 248.400 198.300 249.600 ;
        RECT 196.500 237.600 198.300 248.400 ;
        RECT 203.550 237.600 205.350 249.600 ;
        RECT 208.950 249.300 211.050 250.200 ;
        RECT 211.950 249.300 217.050 250.200 ;
        RECT 219.150 250.500 236.850 251.100 ;
        RECT 219.150 250.200 227.550 250.500 ;
        RECT 211.950 248.400 212.850 249.300 ;
        RECT 210.150 246.600 212.850 248.400 ;
        RECT 213.750 248.100 215.550 248.400 ;
        RECT 219.150 248.100 220.050 250.200 ;
        RECT 235.950 249.600 236.850 250.500 ;
        RECT 213.750 247.200 220.050 248.100 ;
        RECT 220.950 248.700 222.750 249.300 ;
        RECT 220.950 247.500 228.450 248.700 ;
        RECT 213.750 246.600 215.550 247.200 ;
        RECT 227.250 246.600 228.450 247.500 ;
        RECT 208.950 243.600 212.850 245.700 ;
        RECT 217.950 245.550 219.750 246.300 ;
        RECT 222.750 245.550 224.550 246.300 ;
        RECT 217.950 244.500 224.550 245.550 ;
        RECT 227.250 244.500 232.050 246.600 ;
        RECT 206.550 237.000 208.350 240.600 ;
        RECT 211.050 237.600 212.850 243.600 ;
        RECT 215.250 237.000 217.050 243.600 ;
        RECT 218.850 237.600 220.650 244.500 ;
        RECT 227.250 243.600 228.450 244.500 ;
        RECT 221.850 237.000 223.650 243.600 ;
        RECT 226.650 237.600 228.450 243.600 ;
        RECT 232.050 237.000 233.850 243.600 ;
        RECT 235.050 237.600 236.850 249.600 ;
        RECT 248.400 243.600 249.600 256.950 ;
        RECT 263.400 243.600 264.300 263.700 ;
        RECT 269.700 259.200 270.600 266.400 ;
        RECT 284.400 264.300 285.600 266.400 ;
        RECT 286.800 267.300 288.600 272.400 ;
        RECT 289.800 268.200 291.600 273.000 ;
        RECT 292.800 267.300 294.600 272.400 ;
        RECT 286.800 265.950 294.600 267.300 ;
        RECT 302.400 267.300 304.200 272.400 ;
        RECT 305.400 268.200 307.200 273.000 ;
        RECT 308.400 267.300 310.200 272.400 ;
        RECT 302.400 265.950 310.200 267.300 ;
        RECT 311.400 266.400 313.200 272.400 ;
        RECT 323.700 266.400 325.500 273.000 ;
        RECT 311.400 264.300 312.600 266.400 ;
        RECT 328.800 265.200 330.600 272.400 ;
        RECT 341.400 269.400 343.200 273.000 ;
        RECT 344.400 269.400 346.200 272.400 ;
        RECT 347.400 269.400 349.200 273.000 ;
        RECT 359.400 269.400 361.200 273.000 ;
        RECT 362.400 269.400 364.200 272.400 ;
        RECT 284.400 263.250 288.150 264.300 ;
        RECT 280.950 261.450 283.050 262.050 ;
        RECT 275.550 260.550 283.050 261.450 ;
        RECT 265.950 257.100 268.050 259.200 ;
        RECT 268.950 257.100 271.050 259.200 ;
        RECT 266.100 255.300 267.900 257.100 ;
        RECT 269.700 249.600 270.600 257.100 ;
        RECT 275.550 256.050 276.450 260.550 ;
        RECT 280.950 259.950 283.050 260.550 ;
        RECT 284.100 259.050 285.900 260.850 ;
        RECT 286.950 259.050 288.150 263.250 ;
        RECT 308.850 263.250 312.600 264.300 ;
        RECT 326.400 264.300 330.600 265.200 ;
        RECT 340.950 264.450 343.050 265.050 ;
        RECT 290.100 259.050 291.900 260.850 ;
        RECT 305.100 259.050 306.900 260.850 ;
        RECT 308.850 259.050 310.050 263.250 ;
        RECT 311.100 259.050 312.900 260.850 ;
        RECT 323.100 259.200 324.900 261.000 ;
        RECT 326.400 259.200 327.600 264.300 ;
        RECT 335.550 263.550 343.050 264.450 ;
        RECT 329.100 259.200 330.900 261.000 ;
        RECT 283.950 256.950 286.050 259.050 ;
        RECT 286.950 256.950 289.050 259.050 ;
        RECT 289.950 256.950 292.050 259.050 ;
        RECT 292.950 256.950 295.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 304.950 256.950 307.050 259.050 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 310.950 256.950 313.050 259.050 ;
        RECT 322.950 257.100 325.050 259.200 ;
        RECT 325.950 257.100 328.050 259.200 ;
        RECT 328.950 257.100 331.050 259.200 ;
        RECT 271.950 254.550 276.450 256.050 ;
        RECT 271.950 253.950 276.000 254.550 ;
        RECT 245.400 237.000 247.200 243.600 ;
        RECT 248.400 237.600 250.200 243.600 ;
        RECT 260.400 237.000 262.200 243.600 ;
        RECT 263.400 237.600 265.200 243.600 ;
        RECT 266.400 237.000 268.200 243.600 ;
        RECT 269.400 237.600 271.200 249.600 ;
        RECT 287.850 243.600 289.050 256.950 ;
        RECT 293.100 255.150 294.900 256.950 ;
        RECT 302.100 255.150 303.900 256.950 ;
        RECT 284.400 237.000 286.200 243.600 ;
        RECT 287.400 237.600 289.200 243.600 ;
        RECT 292.500 237.000 294.300 249.600 ;
        RECT 302.700 237.000 304.500 249.600 ;
        RECT 307.950 243.600 309.150 256.950 ;
        RECT 310.950 252.450 313.050 253.050 ;
        RECT 322.950 252.450 325.050 252.900 ;
        RECT 310.950 251.550 325.050 252.450 ;
        RECT 310.950 250.950 313.050 251.550 ;
        RECT 322.950 250.800 325.050 251.550 ;
        RECT 326.400 243.600 327.600 257.100 ;
        RECT 328.950 255.450 331.050 256.050 ;
        RECT 335.550 255.450 336.450 263.550 ;
        RECT 340.950 262.950 343.050 263.550 ;
        RECT 344.700 259.050 345.600 269.400 ;
        RECT 362.400 259.050 363.600 269.400 ;
        RECT 377.400 265.200 379.200 272.400 ;
        RECT 382.500 266.400 384.300 273.000 ;
        RECT 392.700 266.400 394.500 273.000 ;
        RECT 397.800 265.200 399.600 272.400 ;
        RECT 410.700 266.400 412.500 273.000 ;
        RECT 415.800 265.200 417.600 272.400 ;
        RECT 377.400 264.300 381.600 265.200 ;
        RECT 377.100 259.200 378.900 261.000 ;
        RECT 380.400 259.200 381.600 264.300 ;
        RECT 395.400 264.300 399.600 265.200 ;
        RECT 413.400 264.300 417.600 265.200 ;
        RECT 428.400 269.400 430.200 272.400 ;
        RECT 431.400 269.400 433.200 273.000 ;
        RECT 428.400 265.500 429.600 269.400 ;
        RECT 434.400 266.400 436.200 272.400 ;
        RECT 423.000 264.450 427.050 265.050 ;
        RECT 428.400 264.600 434.100 265.500 ;
        RECT 383.100 259.200 384.900 261.000 ;
        RECT 392.100 259.200 393.900 261.000 ;
        RECT 395.400 259.200 396.600 264.300 ;
        RECT 398.100 259.200 399.900 261.000 ;
        RECT 410.100 259.200 411.900 261.000 ;
        RECT 413.400 259.200 414.600 264.300 ;
        RECT 422.550 262.950 427.050 264.450 ;
        RECT 432.150 263.700 434.100 264.600 ;
        RECT 416.100 259.200 417.900 261.000 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 376.950 257.100 379.050 259.200 ;
        RECT 379.950 257.100 382.050 259.200 ;
        RECT 382.950 257.100 385.050 259.200 ;
        RECT 391.950 257.100 394.050 259.200 ;
        RECT 394.950 257.100 397.050 259.200 ;
        RECT 397.950 257.100 400.050 259.200 ;
        RECT 409.950 257.100 412.050 259.200 ;
        RECT 412.950 257.100 415.050 259.200 ;
        RECT 415.950 257.100 418.050 259.200 ;
        RECT 328.950 254.550 336.450 255.450 ;
        RECT 341.100 255.150 342.900 256.950 ;
        RECT 328.950 253.950 331.050 254.550 ;
        RECT 344.700 249.600 345.600 256.950 ;
        RECT 347.100 255.150 348.900 256.950 ;
        RECT 359.100 255.150 360.900 256.950 ;
        RECT 307.800 237.600 309.600 243.600 ;
        RECT 310.800 237.000 312.600 243.600 ;
        RECT 323.400 237.000 325.200 243.600 ;
        RECT 326.400 237.600 328.200 243.600 ;
        RECT 329.400 237.000 331.200 243.600 ;
        RECT 341.400 237.000 343.200 249.600 ;
        RECT 344.700 248.400 348.300 249.600 ;
        RECT 346.500 237.600 348.300 248.400 ;
        RECT 362.400 243.600 363.600 256.950 ;
        RECT 380.400 243.600 381.600 257.100 ;
        RECT 395.400 243.600 396.600 257.100 ;
        RECT 413.400 243.600 414.600 257.100 ;
        RECT 415.950 255.450 418.050 256.050 ;
        RECT 422.550 255.450 423.450 262.950 ;
        RECT 427.950 256.950 430.050 259.050 ;
        RECT 415.950 254.550 423.450 255.450 ;
        RECT 428.100 255.150 429.900 256.950 ;
        RECT 415.950 253.950 418.050 254.550 ;
        RECT 432.150 252.300 433.050 263.700 ;
        RECT 435.000 259.050 436.200 266.400 ;
        RECT 446.400 267.300 448.200 272.400 ;
        RECT 449.400 268.200 451.200 273.000 ;
        RECT 452.400 267.300 454.200 272.400 ;
        RECT 446.400 265.950 454.200 267.300 ;
        RECT 455.400 266.400 457.200 272.400 ;
        RECT 455.400 264.300 456.600 266.400 ;
        RECT 470.400 265.200 472.200 272.400 ;
        RECT 475.500 266.400 477.300 273.000 ;
        RECT 480.150 266.400 481.950 272.400 ;
        RECT 483.150 269.400 484.950 273.000 ;
        RECT 487.950 270.300 489.750 272.400 ;
        RECT 486.000 269.400 489.750 270.300 ;
        RECT 492.450 269.400 494.250 273.000 ;
        RECT 495.750 269.400 497.550 272.400 ;
        RECT 499.350 269.400 501.150 273.000 ;
        RECT 503.550 269.400 505.350 272.400 ;
        RECT 508.350 269.400 510.150 273.000 ;
        RECT 486.000 268.500 487.050 269.400 ;
        RECT 495.750 268.500 496.800 269.400 ;
        RECT 484.950 266.400 487.050 268.500 ;
        RECT 470.400 264.300 474.600 265.200 ;
        RECT 452.850 263.250 456.600 264.300 ;
        RECT 449.100 259.050 450.900 260.850 ;
        RECT 452.850 259.050 454.050 263.250 ;
        RECT 455.100 259.050 456.900 260.850 ;
        RECT 470.100 259.200 471.900 261.000 ;
        RECT 473.400 259.200 474.600 264.300 ;
        RECT 476.100 259.200 477.900 261.000 ;
        RECT 433.950 256.950 436.200 259.050 ;
        RECT 445.950 256.950 448.050 259.050 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 451.950 256.950 454.050 259.050 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 469.950 257.100 472.050 259.200 ;
        RECT 472.950 257.100 475.050 259.200 ;
        RECT 475.950 257.100 478.050 259.200 ;
        RECT 432.150 251.400 434.100 252.300 ;
        RECT 428.400 250.500 434.100 251.400 ;
        RECT 428.400 243.600 429.600 250.500 ;
        RECT 435.000 249.600 436.200 256.950 ;
        RECT 446.100 255.150 447.900 256.950 ;
        RECT 359.400 237.000 361.200 243.600 ;
        RECT 362.400 237.600 364.200 243.600 ;
        RECT 376.800 237.000 378.600 243.600 ;
        RECT 379.800 237.600 381.600 243.600 ;
        RECT 382.800 237.000 384.600 243.600 ;
        RECT 392.400 237.000 394.200 243.600 ;
        RECT 395.400 237.600 397.200 243.600 ;
        RECT 398.400 237.000 400.200 243.600 ;
        RECT 410.400 237.000 412.200 243.600 ;
        RECT 413.400 237.600 415.200 243.600 ;
        RECT 416.400 237.000 418.200 243.600 ;
        RECT 428.400 237.600 430.200 243.600 ;
        RECT 431.400 237.000 433.200 243.600 ;
        RECT 434.400 237.600 436.200 249.600 ;
        RECT 446.700 237.000 448.500 249.600 ;
        RECT 451.950 243.600 453.150 256.950 ;
        RECT 473.400 243.600 474.600 257.100 ;
        RECT 480.150 251.700 481.050 266.400 ;
        RECT 488.550 265.800 490.350 267.600 ;
        RECT 491.850 267.450 496.800 268.500 ;
        RECT 504.300 268.500 505.350 269.400 ;
        RECT 491.850 266.700 493.650 267.450 ;
        RECT 504.300 267.300 508.050 268.500 ;
        RECT 505.950 266.400 508.050 267.300 ;
        RECT 511.650 266.400 513.450 272.400 ;
        RECT 521.700 266.400 523.500 273.000 ;
        RECT 526.200 266.400 528.000 272.400 ;
        RECT 530.700 266.400 532.500 273.000 ;
        RECT 540.150 266.400 541.950 272.400 ;
        RECT 543.150 269.400 544.950 273.000 ;
        RECT 547.950 270.300 549.750 272.400 ;
        RECT 546.000 269.400 549.750 270.300 ;
        RECT 552.450 269.400 554.250 273.000 ;
        RECT 555.750 269.400 557.550 272.400 ;
        RECT 559.350 269.400 561.150 273.000 ;
        RECT 563.550 269.400 565.350 272.400 ;
        RECT 568.350 269.400 570.150 273.000 ;
        RECT 546.000 268.500 547.050 269.400 ;
        RECT 555.750 268.500 556.800 269.400 ;
        RECT 544.950 266.400 547.050 268.500 ;
        RECT 488.850 264.000 489.900 265.800 ;
        RECT 499.050 264.000 500.850 264.600 ;
        RECT 488.850 262.800 500.850 264.000 ;
        RECT 483.000 261.600 489.900 262.800 ;
        RECT 483.000 260.850 483.900 261.600 ;
        RECT 488.100 261.000 489.900 261.600 ;
        RECT 482.100 259.050 483.900 260.850 ;
        RECT 485.100 259.800 486.900 260.400 ;
        RECT 481.950 256.950 484.050 259.050 ;
        RECT 485.100 258.600 493.050 259.800 ;
        RECT 490.950 256.950 493.050 258.600 ;
        RECT 489.450 251.700 491.250 252.000 ;
        RECT 480.150 251.100 491.250 251.700 ;
        RECT 480.150 250.500 497.850 251.100 ;
        RECT 480.150 249.600 481.050 250.500 ;
        RECT 489.450 250.200 497.850 250.500 ;
        RECT 451.800 237.600 453.600 243.600 ;
        RECT 454.800 237.000 456.600 243.600 ;
        RECT 469.800 237.000 471.600 243.600 ;
        RECT 472.800 237.600 474.600 243.600 ;
        RECT 475.800 237.000 477.600 243.600 ;
        RECT 480.150 237.600 481.950 249.600 ;
        RECT 494.250 248.700 496.050 249.300 ;
        RECT 488.550 247.500 496.050 248.700 ;
        RECT 496.950 248.100 497.850 250.200 ;
        RECT 499.950 250.200 500.850 262.800 ;
        RECT 512.250 259.050 513.450 266.400 ;
        RECT 521.100 259.200 522.900 261.000 ;
        RECT 526.950 259.200 528.000 266.400 ;
        RECT 533.100 259.200 534.900 261.000 ;
        RECT 507.150 257.250 513.450 259.050 ;
        RECT 508.950 256.950 513.450 257.250 ;
        RECT 520.950 257.100 523.050 259.200 ;
        RECT 523.950 257.100 526.050 259.200 ;
        RECT 526.950 257.100 529.050 259.200 ;
        RECT 529.950 257.100 532.050 259.200 ;
        RECT 532.950 257.100 535.050 259.200 ;
        RECT 509.250 251.400 511.050 253.200 ;
        RECT 505.950 250.200 510.150 251.400 ;
        RECT 499.950 249.300 505.050 250.200 ;
        RECT 505.950 249.300 508.050 250.200 ;
        RECT 512.250 249.600 513.450 256.950 ;
        RECT 514.950 255.450 517.050 256.050 ;
        RECT 520.950 255.450 523.050 256.050 ;
        RECT 514.950 254.550 523.050 255.450 ;
        RECT 524.100 255.300 525.900 257.100 ;
        RECT 514.950 253.950 517.050 254.550 ;
        RECT 520.950 253.950 523.050 254.550 ;
        RECT 527.100 251.400 528.000 257.100 ;
        RECT 530.100 255.300 531.900 257.100 ;
        RECT 540.150 251.700 541.050 266.400 ;
        RECT 548.550 265.800 550.350 267.600 ;
        RECT 551.850 267.450 556.800 268.500 ;
        RECT 564.300 268.500 565.350 269.400 ;
        RECT 551.850 266.700 553.650 267.450 ;
        RECT 564.300 267.300 568.050 268.500 ;
        RECT 565.950 266.400 568.050 267.300 ;
        RECT 571.650 266.400 573.450 272.400 ;
        RECT 548.850 264.000 549.900 265.800 ;
        RECT 559.050 264.000 560.850 264.600 ;
        RECT 548.850 262.800 560.850 264.000 ;
        RECT 543.000 261.600 549.900 262.800 ;
        RECT 543.000 260.850 543.900 261.600 ;
        RECT 548.100 261.000 549.900 261.600 ;
        RECT 542.100 259.050 543.900 260.850 ;
        RECT 545.100 259.800 546.900 260.400 ;
        RECT 541.950 256.950 544.050 259.050 ;
        RECT 545.100 258.600 553.050 259.800 ;
        RECT 550.950 256.950 553.050 258.600 ;
        RECT 549.450 251.700 551.250 252.000 ;
        RECT 527.100 250.500 532.200 251.400 ;
        RECT 504.150 248.400 505.050 249.300 ;
        RECT 501.450 248.100 503.250 248.400 ;
        RECT 488.550 246.600 489.750 247.500 ;
        RECT 496.950 247.200 503.250 248.100 ;
        RECT 501.450 246.600 503.250 247.200 ;
        RECT 504.150 246.600 506.850 248.400 ;
        RECT 484.950 244.500 489.750 246.600 ;
        RECT 492.450 245.550 494.250 246.300 ;
        RECT 497.250 245.550 499.050 246.300 ;
        RECT 492.450 244.500 499.050 245.550 ;
        RECT 488.550 243.600 489.750 244.500 ;
        RECT 483.150 237.000 484.950 243.600 ;
        RECT 488.550 237.600 490.350 243.600 ;
        RECT 493.350 237.000 495.150 243.600 ;
        RECT 496.350 237.600 498.150 244.500 ;
        RECT 504.150 243.600 508.050 245.700 ;
        RECT 499.950 237.000 501.750 243.600 ;
        RECT 504.150 237.600 505.950 243.600 ;
        RECT 508.650 237.000 510.450 240.600 ;
        RECT 511.650 237.600 513.450 249.600 ;
        RECT 521.400 248.400 529.200 249.300 ;
        RECT 521.400 237.600 523.200 248.400 ;
        RECT 524.400 237.000 526.200 247.500 ;
        RECT 527.400 238.500 529.200 248.400 ;
        RECT 530.400 239.400 532.200 250.500 ;
        RECT 540.150 251.100 551.250 251.700 ;
        RECT 540.150 250.500 557.850 251.100 ;
        RECT 540.150 249.600 541.050 250.500 ;
        RECT 549.450 250.200 557.850 250.500 ;
        RECT 533.400 238.500 535.200 249.600 ;
        RECT 527.400 237.600 535.200 238.500 ;
        RECT 540.150 237.600 541.950 249.600 ;
        RECT 554.250 248.700 556.050 249.300 ;
        RECT 548.550 247.500 556.050 248.700 ;
        RECT 556.950 248.100 557.850 250.200 ;
        RECT 559.950 250.200 560.850 262.800 ;
        RECT 572.250 259.050 573.450 266.400 ;
        RECT 584.400 265.200 586.200 272.400 ;
        RECT 589.500 266.400 591.300 273.000 ;
        RECT 599.400 267.300 601.200 272.400 ;
        RECT 602.400 268.200 604.200 273.000 ;
        RECT 605.400 267.300 607.200 272.400 ;
        RECT 599.400 265.950 607.200 267.300 ;
        RECT 608.400 266.400 610.200 272.400 ;
        RECT 622.800 269.400 624.600 272.400 ;
        RECT 625.800 269.400 627.600 273.000 ;
        RECT 584.400 264.300 588.600 265.200 ;
        RECT 608.400 264.300 609.600 266.400 ;
        RECT 584.100 259.200 585.900 261.000 ;
        RECT 587.400 259.200 588.600 264.300 ;
        RECT 605.850 263.250 609.600 264.300 ;
        RECT 590.100 259.200 591.900 261.000 ;
        RECT 567.150 257.250 573.450 259.050 ;
        RECT 568.950 256.950 573.450 257.250 ;
        RECT 583.950 257.100 586.050 259.200 ;
        RECT 586.950 257.100 589.050 259.200 ;
        RECT 589.950 257.100 592.050 259.200 ;
        RECT 602.100 259.050 603.900 260.850 ;
        RECT 605.850 259.050 607.050 263.250 ;
        RECT 608.100 259.050 609.900 260.850 ;
        RECT 623.400 259.050 624.600 269.400 ;
        RECT 630.150 266.400 631.950 272.400 ;
        RECT 633.150 269.400 634.950 273.000 ;
        RECT 637.950 270.300 639.750 272.400 ;
        RECT 636.000 269.400 639.750 270.300 ;
        RECT 642.450 269.400 644.250 273.000 ;
        RECT 645.750 269.400 647.550 272.400 ;
        RECT 649.350 269.400 651.150 273.000 ;
        RECT 653.550 269.400 655.350 272.400 ;
        RECT 658.350 269.400 660.150 273.000 ;
        RECT 636.000 268.500 637.050 269.400 ;
        RECT 645.750 268.500 646.800 269.400 ;
        RECT 634.950 266.400 637.050 268.500 ;
        RECT 569.250 251.400 571.050 253.200 ;
        RECT 565.950 250.200 570.150 251.400 ;
        RECT 559.950 249.300 565.050 250.200 ;
        RECT 565.950 249.300 568.050 250.200 ;
        RECT 572.250 249.600 573.450 256.950 ;
        RECT 564.150 248.400 565.050 249.300 ;
        RECT 561.450 248.100 563.250 248.400 ;
        RECT 548.550 246.600 549.750 247.500 ;
        RECT 556.950 247.200 563.250 248.100 ;
        RECT 561.450 246.600 563.250 247.200 ;
        RECT 564.150 246.600 566.850 248.400 ;
        RECT 544.950 244.500 549.750 246.600 ;
        RECT 552.450 245.550 554.250 246.300 ;
        RECT 557.250 245.550 559.050 246.300 ;
        RECT 552.450 244.500 559.050 245.550 ;
        RECT 548.550 243.600 549.750 244.500 ;
        RECT 543.150 237.000 544.950 243.600 ;
        RECT 548.550 237.600 550.350 243.600 ;
        RECT 553.350 237.000 555.150 243.600 ;
        RECT 556.350 237.600 558.150 244.500 ;
        RECT 564.150 243.600 568.050 245.700 ;
        RECT 559.950 237.000 561.750 243.600 ;
        RECT 564.150 237.600 565.950 243.600 ;
        RECT 568.650 237.000 570.450 240.600 ;
        RECT 571.650 237.600 573.450 249.600 ;
        RECT 587.400 243.600 588.600 257.100 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 622.950 256.950 625.050 259.050 ;
        RECT 625.950 256.950 628.050 259.050 ;
        RECT 599.100 255.150 600.900 256.950 ;
        RECT 583.800 237.000 585.600 243.600 ;
        RECT 586.800 237.600 588.600 243.600 ;
        RECT 589.800 237.000 591.600 243.600 ;
        RECT 599.700 237.000 601.500 249.600 ;
        RECT 604.950 243.600 606.150 256.950 ;
        RECT 623.400 243.600 624.600 256.950 ;
        RECT 626.100 255.150 627.900 256.950 ;
        RECT 630.150 251.700 631.050 266.400 ;
        RECT 638.550 265.800 640.350 267.600 ;
        RECT 641.850 267.450 646.800 268.500 ;
        RECT 654.300 268.500 655.350 269.400 ;
        RECT 641.850 266.700 643.650 267.450 ;
        RECT 654.300 267.300 658.050 268.500 ;
        RECT 655.950 266.400 658.050 267.300 ;
        RECT 661.650 266.400 663.450 272.400 ;
        RECT 673.800 269.400 675.600 273.000 ;
        RECT 676.800 269.400 678.600 272.400 ;
        RECT 679.800 269.400 681.600 273.000 ;
        RECT 638.850 264.000 639.900 265.800 ;
        RECT 649.050 264.000 650.850 264.600 ;
        RECT 638.850 262.800 650.850 264.000 ;
        RECT 633.000 261.600 639.900 262.800 ;
        RECT 633.000 260.850 633.900 261.600 ;
        RECT 638.100 261.000 639.900 261.600 ;
        RECT 632.100 259.050 633.900 260.850 ;
        RECT 635.100 259.800 636.900 260.400 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 635.100 258.600 643.050 259.800 ;
        RECT 640.950 256.950 643.050 258.600 ;
        RECT 639.450 251.700 641.250 252.000 ;
        RECT 630.150 251.100 641.250 251.700 ;
        RECT 630.150 250.500 647.850 251.100 ;
        RECT 630.150 249.600 631.050 250.500 ;
        RECT 639.450 250.200 647.850 250.500 ;
        RECT 604.800 237.600 606.600 243.600 ;
        RECT 607.800 237.000 609.600 243.600 ;
        RECT 622.800 237.600 624.600 243.600 ;
        RECT 625.800 237.000 627.600 243.600 ;
        RECT 630.150 237.600 631.950 249.600 ;
        RECT 644.250 248.700 646.050 249.300 ;
        RECT 638.550 247.500 646.050 248.700 ;
        RECT 646.950 248.100 647.850 250.200 ;
        RECT 649.950 250.200 650.850 262.800 ;
        RECT 662.250 259.050 663.450 266.400 ;
        RECT 677.400 259.050 678.300 269.400 ;
        RECT 691.800 266.400 693.600 272.400 ;
        RECT 692.400 264.300 693.600 266.400 ;
        RECT 694.800 267.300 696.600 272.400 ;
        RECT 697.800 268.200 699.600 273.000 ;
        RECT 700.800 267.300 702.600 272.400 ;
        RECT 712.800 269.400 714.600 272.400 ;
        RECT 715.800 269.400 717.600 273.000 ;
        RECT 727.800 269.400 729.600 273.000 ;
        RECT 730.800 269.400 732.600 272.400 ;
        RECT 733.800 269.400 735.600 273.000 ;
        RECT 694.800 265.950 702.600 267.300 ;
        RECT 692.400 263.250 696.150 264.300 ;
        RECT 692.100 259.050 693.900 260.850 ;
        RECT 694.950 259.050 696.150 263.250 ;
        RECT 708.000 261.450 712.050 262.050 ;
        RECT 707.550 261.000 712.050 261.450 ;
        RECT 698.100 259.050 699.900 260.850 ;
        RECT 706.950 259.950 712.050 261.000 ;
        RECT 657.150 257.250 663.450 259.050 ;
        RECT 658.950 256.950 663.450 257.250 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 691.950 256.950 694.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 700.950 256.950 703.050 259.050 ;
        RECT 659.250 251.400 661.050 253.200 ;
        RECT 655.950 250.200 660.150 251.400 ;
        RECT 649.950 249.300 655.050 250.200 ;
        RECT 655.950 249.300 658.050 250.200 ;
        RECT 662.250 249.600 663.450 256.950 ;
        RECT 674.100 255.150 675.900 256.950 ;
        RECT 667.950 252.450 670.050 253.050 ;
        RECT 673.950 252.450 676.050 253.050 ;
        RECT 667.950 251.550 676.050 252.450 ;
        RECT 667.950 250.950 670.050 251.550 ;
        RECT 673.950 250.950 676.050 251.550 ;
        RECT 677.400 249.600 678.300 256.950 ;
        RECT 680.100 255.150 681.900 256.950 ;
        RECT 654.150 248.400 655.050 249.300 ;
        RECT 651.450 248.100 653.250 248.400 ;
        RECT 638.550 246.600 639.750 247.500 ;
        RECT 646.950 247.200 653.250 248.100 ;
        RECT 651.450 246.600 653.250 247.200 ;
        RECT 654.150 246.600 656.850 248.400 ;
        RECT 634.950 244.500 639.750 246.600 ;
        RECT 642.450 245.550 644.250 246.300 ;
        RECT 647.250 245.550 649.050 246.300 ;
        RECT 642.450 244.500 649.050 245.550 ;
        RECT 638.550 243.600 639.750 244.500 ;
        RECT 633.150 237.000 634.950 243.600 ;
        RECT 638.550 237.600 640.350 243.600 ;
        RECT 643.350 237.000 645.150 243.600 ;
        RECT 646.350 237.600 648.150 244.500 ;
        RECT 654.150 243.600 658.050 245.700 ;
        RECT 649.950 237.000 651.750 243.600 ;
        RECT 654.150 237.600 655.950 243.600 ;
        RECT 658.650 237.000 660.450 240.600 ;
        RECT 661.650 237.600 663.450 249.600 ;
        RECT 674.700 248.400 678.300 249.600 ;
        RECT 674.700 237.600 676.500 248.400 ;
        RECT 679.800 237.000 681.600 249.600 ;
        RECT 695.850 243.600 697.050 256.950 ;
        RECT 701.100 255.150 702.900 256.950 ;
        RECT 706.950 256.800 709.050 259.950 ;
        RECT 713.400 259.050 714.600 269.400 ;
        RECT 718.950 261.450 723.000 262.050 ;
        RECT 718.950 259.950 723.450 261.450 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 692.400 237.000 694.200 243.600 ;
        RECT 695.400 237.600 697.200 243.600 ;
        RECT 700.500 237.000 702.300 249.600 ;
        RECT 713.400 243.600 714.600 256.950 ;
        RECT 716.100 255.150 717.900 256.950 ;
        RECT 722.550 256.050 723.450 259.950 ;
        RECT 731.400 259.050 732.300 269.400 ;
        RECT 744.000 266.400 745.800 273.000 ;
        RECT 748.500 267.600 750.300 272.400 ;
        RECT 751.500 269.400 753.300 273.000 ;
        RECT 764.400 269.400 766.200 273.000 ;
        RECT 767.400 269.400 769.200 272.400 ;
        RECT 770.400 269.400 772.200 273.000 ;
        RECT 748.500 266.400 753.600 267.600 ;
        RECT 743.100 259.200 744.900 261.000 ;
        RECT 749.100 259.200 750.900 261.000 ;
        RECT 752.700 259.200 753.600 266.400 ;
        RECT 754.950 261.450 759.000 262.050 ;
        RECT 754.950 259.950 759.450 261.450 ;
        RECT 727.950 256.950 730.050 259.050 ;
        RECT 730.950 256.950 733.050 259.050 ;
        RECT 733.950 256.950 736.050 259.050 ;
        RECT 742.950 257.100 745.050 259.200 ;
        RECT 745.950 257.100 748.050 259.200 ;
        RECT 748.950 257.100 751.050 259.200 ;
        RECT 751.950 257.100 754.050 259.200 ;
        RECT 718.950 254.550 723.450 256.050 ;
        RECT 728.100 255.150 729.900 256.950 ;
        RECT 718.950 253.950 723.000 254.550 ;
        RECT 731.400 249.600 732.300 256.950 ;
        RECT 734.100 255.150 735.900 256.950 ;
        RECT 746.100 255.300 747.900 257.100 ;
        RECT 752.700 249.600 753.600 257.100 ;
        RECT 758.550 256.050 759.450 259.950 ;
        RECT 767.700 259.050 768.600 269.400 ;
        RECT 784.800 266.400 786.600 272.400 ;
        RECT 785.400 264.300 786.600 266.400 ;
        RECT 787.800 267.300 789.600 272.400 ;
        RECT 790.800 268.200 792.600 273.000 ;
        RECT 793.800 267.300 795.600 272.400 ;
        RECT 803.400 269.400 805.200 273.000 ;
        RECT 806.400 269.400 808.200 272.400 ;
        RECT 787.800 265.950 795.600 267.300 ;
        RECT 785.400 263.250 789.150 264.300 ;
        RECT 785.100 259.050 786.900 260.850 ;
        RECT 787.950 259.050 789.150 263.250 ;
        RECT 791.100 259.050 792.900 260.850 ;
        RECT 806.400 259.050 807.600 269.400 ;
        RECT 813.150 266.400 814.950 272.400 ;
        RECT 816.150 269.400 817.950 273.000 ;
        RECT 820.950 270.300 822.750 272.400 ;
        RECT 819.000 269.400 822.750 270.300 ;
        RECT 825.450 269.400 827.250 273.000 ;
        RECT 828.750 269.400 830.550 272.400 ;
        RECT 832.350 269.400 834.150 273.000 ;
        RECT 836.550 269.400 838.350 272.400 ;
        RECT 841.350 269.400 843.150 273.000 ;
        RECT 819.000 268.500 820.050 269.400 ;
        RECT 828.750 268.500 829.800 269.400 ;
        RECT 817.950 266.400 820.050 268.500 ;
        RECT 763.950 256.950 766.050 259.050 ;
        RECT 766.950 256.950 769.050 259.050 ;
        RECT 769.950 256.950 772.050 259.050 ;
        RECT 784.950 256.950 787.050 259.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 754.950 254.550 759.450 256.050 ;
        RECT 764.100 255.150 765.900 256.950 ;
        RECT 754.950 253.950 759.000 254.550 ;
        RECT 767.700 249.600 768.600 256.950 ;
        RECT 770.100 255.150 771.900 256.950 ;
        RECT 728.700 248.400 732.300 249.600 ;
        RECT 712.800 237.600 714.600 243.600 ;
        RECT 715.800 237.000 717.600 243.600 ;
        RECT 728.700 237.600 730.500 248.400 ;
        RECT 733.800 237.000 735.600 249.600 ;
        RECT 743.400 248.700 751.200 249.600 ;
        RECT 743.400 237.600 745.200 248.700 ;
        RECT 746.400 237.000 748.200 247.800 ;
        RECT 749.400 237.600 751.200 248.700 ;
        RECT 752.400 237.600 754.200 249.600 ;
        RECT 764.400 237.000 766.200 249.600 ;
        RECT 767.700 248.400 771.300 249.600 ;
        RECT 769.500 237.600 771.300 248.400 ;
        RECT 788.850 243.600 790.050 256.950 ;
        RECT 794.100 255.150 795.900 256.950 ;
        RECT 803.100 255.150 804.900 256.950 ;
        RECT 785.400 237.000 787.200 243.600 ;
        RECT 788.400 237.600 790.200 243.600 ;
        RECT 793.500 237.000 795.300 249.600 ;
        RECT 806.400 243.600 807.600 256.950 ;
        RECT 813.150 251.700 814.050 266.400 ;
        RECT 821.550 265.800 823.350 267.600 ;
        RECT 824.850 267.450 829.800 268.500 ;
        RECT 837.300 268.500 838.350 269.400 ;
        RECT 824.850 266.700 826.650 267.450 ;
        RECT 837.300 267.300 841.050 268.500 ;
        RECT 838.950 266.400 841.050 267.300 ;
        RECT 844.650 266.400 846.450 272.400 ;
        RECT 821.850 264.000 822.900 265.800 ;
        RECT 832.050 264.000 833.850 264.600 ;
        RECT 821.850 262.800 833.850 264.000 ;
        RECT 816.000 261.600 822.900 262.800 ;
        RECT 816.000 260.850 816.900 261.600 ;
        RECT 821.100 261.000 822.900 261.600 ;
        RECT 815.100 259.050 816.900 260.850 ;
        RECT 818.100 259.800 819.900 260.400 ;
        RECT 814.950 256.950 817.050 259.050 ;
        RECT 818.100 258.600 826.050 259.800 ;
        RECT 823.950 256.950 826.050 258.600 ;
        RECT 822.450 251.700 824.250 252.000 ;
        RECT 813.150 251.100 824.250 251.700 ;
        RECT 813.150 250.500 830.850 251.100 ;
        RECT 813.150 249.600 814.050 250.500 ;
        RECT 822.450 250.200 830.850 250.500 ;
        RECT 803.400 237.000 805.200 243.600 ;
        RECT 806.400 237.600 808.200 243.600 ;
        RECT 813.150 237.600 814.950 249.600 ;
        RECT 827.250 248.700 829.050 249.300 ;
        RECT 821.550 247.500 829.050 248.700 ;
        RECT 829.950 248.100 830.850 250.200 ;
        RECT 832.950 250.200 833.850 262.800 ;
        RECT 845.250 259.050 846.450 266.400 ;
        RECT 840.150 257.250 846.450 259.050 ;
        RECT 841.950 256.950 846.450 257.250 ;
        RECT 842.250 251.400 844.050 253.200 ;
        RECT 838.950 250.200 843.150 251.400 ;
        RECT 832.950 249.300 838.050 250.200 ;
        RECT 838.950 249.300 841.050 250.200 ;
        RECT 845.250 249.600 846.450 256.950 ;
        RECT 837.150 248.400 838.050 249.300 ;
        RECT 834.450 248.100 836.250 248.400 ;
        RECT 821.550 246.600 822.750 247.500 ;
        RECT 829.950 247.200 836.250 248.100 ;
        RECT 834.450 246.600 836.250 247.200 ;
        RECT 837.150 246.600 839.850 248.400 ;
        RECT 817.950 244.500 822.750 246.600 ;
        RECT 825.450 245.550 827.250 246.300 ;
        RECT 830.250 245.550 832.050 246.300 ;
        RECT 825.450 244.500 832.050 245.550 ;
        RECT 821.550 243.600 822.750 244.500 ;
        RECT 816.150 237.000 817.950 243.600 ;
        RECT 821.550 237.600 823.350 243.600 ;
        RECT 826.350 237.000 828.150 243.600 ;
        RECT 829.350 237.600 831.150 244.500 ;
        RECT 837.150 243.600 841.050 245.700 ;
        RECT 832.950 237.000 834.750 243.600 ;
        RECT 837.150 237.600 838.950 243.600 ;
        RECT 841.650 237.000 843.450 240.600 ;
        RECT 844.650 237.600 846.450 249.600 ;
        RECT 2.550 221.400 4.350 233.400 ;
        RECT 5.550 230.400 7.350 234.000 ;
        RECT 10.050 227.400 11.850 233.400 ;
        RECT 14.250 227.400 16.050 234.000 ;
        RECT 7.950 225.300 11.850 227.400 ;
        RECT 17.850 226.500 19.650 233.400 ;
        RECT 20.850 227.400 22.650 234.000 ;
        RECT 25.650 227.400 27.450 233.400 ;
        RECT 31.050 227.400 32.850 234.000 ;
        RECT 26.250 226.500 27.450 227.400 ;
        RECT 16.950 225.450 23.550 226.500 ;
        RECT 16.950 224.700 18.750 225.450 ;
        RECT 21.750 224.700 23.550 225.450 ;
        RECT 26.250 224.400 31.050 226.500 ;
        RECT 9.150 222.600 11.850 224.400 ;
        RECT 12.750 223.800 14.550 224.400 ;
        RECT 12.750 222.900 19.050 223.800 ;
        RECT 26.250 223.500 27.450 224.400 ;
        RECT 12.750 222.600 14.550 222.900 ;
        RECT 10.950 221.700 11.850 222.600 ;
        RECT 2.550 214.050 3.750 221.400 ;
        RECT 7.950 220.800 10.050 221.700 ;
        RECT 10.950 220.800 16.050 221.700 ;
        RECT 5.850 219.600 10.050 220.800 ;
        RECT 4.950 217.800 6.750 219.600 ;
        RECT 2.550 213.750 7.050 214.050 ;
        RECT 2.550 211.950 8.850 213.750 ;
        RECT 2.550 204.600 3.750 211.950 ;
        RECT 15.150 208.200 16.050 220.800 ;
        RECT 18.150 220.800 19.050 222.900 ;
        RECT 19.950 222.300 27.450 223.500 ;
        RECT 19.950 221.700 21.750 222.300 ;
        RECT 34.050 221.400 35.850 233.400 ;
        RECT 46.800 221.400 48.600 233.400 ;
        RECT 49.800 227.400 51.600 234.000 ;
        RECT 52.800 227.400 54.600 233.400 ;
        RECT 55.800 227.400 57.600 234.000 ;
        RECT 18.150 220.500 26.550 220.800 ;
        RECT 34.950 220.500 35.850 221.400 ;
        RECT 18.150 219.900 35.850 220.500 ;
        RECT 24.750 219.300 35.850 219.900 ;
        RECT 24.750 219.000 26.550 219.300 ;
        RECT 22.950 212.400 25.050 214.050 ;
        RECT 22.950 211.200 30.900 212.400 ;
        RECT 31.950 211.950 34.050 214.050 ;
        RECT 29.100 210.600 30.900 211.200 ;
        RECT 32.100 210.150 33.900 211.950 ;
        RECT 26.100 209.400 27.900 210.000 ;
        RECT 32.100 209.400 33.000 210.150 ;
        RECT 26.100 208.200 33.000 209.400 ;
        RECT 15.150 207.000 27.150 208.200 ;
        RECT 15.150 206.400 16.950 207.000 ;
        RECT 26.100 205.200 27.150 207.000 ;
        RECT 2.550 198.600 4.350 204.600 ;
        RECT 7.950 203.700 10.050 204.600 ;
        RECT 7.950 202.500 11.700 203.700 ;
        RECT 22.350 203.550 24.150 204.300 ;
        RECT 10.650 201.600 11.700 202.500 ;
        RECT 19.200 202.500 24.150 203.550 ;
        RECT 25.650 203.400 27.450 205.200 ;
        RECT 34.950 204.600 35.850 219.300 ;
        RECT 47.400 213.900 48.300 221.400 ;
        RECT 50.100 213.900 51.900 215.700 ;
        RECT 46.950 211.800 49.050 213.900 ;
        RECT 49.950 211.800 52.050 213.900 ;
        RECT 28.950 202.500 31.050 204.600 ;
        RECT 19.200 201.600 20.250 202.500 ;
        RECT 28.950 201.600 30.000 202.500 ;
        RECT 5.850 198.000 7.650 201.600 ;
        RECT 10.650 198.600 12.450 201.600 ;
        RECT 14.850 198.000 16.650 201.600 ;
        RECT 18.450 198.600 20.250 201.600 ;
        RECT 21.750 198.000 23.550 201.600 ;
        RECT 26.250 200.700 30.000 201.600 ;
        RECT 26.250 198.600 28.050 200.700 ;
        RECT 31.050 198.000 32.850 201.600 ;
        RECT 34.050 198.600 35.850 204.600 ;
        RECT 47.400 204.600 48.300 211.800 ;
        RECT 53.700 207.300 54.600 227.400 ;
        RECT 65.400 221.400 67.200 234.000 ;
        RECT 70.500 222.600 72.300 233.400 ;
        RECT 83.400 227.400 85.200 234.000 ;
        RECT 86.400 227.400 88.200 233.400 ;
        RECT 100.800 227.400 102.600 233.400 ;
        RECT 103.800 227.400 105.600 234.000 ;
        RECT 68.700 221.400 72.300 222.600 ;
        RECT 65.100 214.050 66.900 215.850 ;
        RECT 68.700 214.050 69.600 221.400 ;
        RECT 71.100 214.050 72.900 215.850 ;
        RECT 83.100 214.050 84.900 215.850 ;
        RECT 86.400 214.050 87.600 227.400 ;
        RECT 101.400 214.050 102.600 227.400 ;
        RECT 113.700 221.400 115.500 234.000 ;
        RECT 118.800 227.400 120.600 233.400 ;
        RECT 121.800 227.400 123.600 234.000 ;
        RECT 103.950 219.450 106.050 220.050 ;
        RECT 112.950 219.450 115.050 220.050 ;
        RECT 103.950 218.550 115.050 219.450 ;
        RECT 103.950 217.950 106.050 218.550 ;
        RECT 112.950 217.950 115.050 218.550 ;
        RECT 104.100 214.050 105.900 215.850 ;
        RECT 113.100 214.050 114.900 215.850 ;
        RECT 118.950 214.050 120.150 227.400 ;
        RECT 129.150 221.400 130.950 233.400 ;
        RECT 132.150 227.400 133.950 234.000 ;
        RECT 137.550 227.400 139.350 233.400 ;
        RECT 142.350 227.400 144.150 234.000 ;
        RECT 137.550 226.500 138.750 227.400 ;
        RECT 145.350 226.500 147.150 233.400 ;
        RECT 148.950 227.400 150.750 234.000 ;
        RECT 153.150 227.400 154.950 233.400 ;
        RECT 157.650 230.400 159.450 234.000 ;
        RECT 133.950 224.400 138.750 226.500 ;
        RECT 141.450 225.450 148.050 226.500 ;
        RECT 141.450 224.700 143.250 225.450 ;
        RECT 146.250 224.700 148.050 225.450 ;
        RECT 153.150 225.300 157.050 227.400 ;
        RECT 137.550 223.500 138.750 224.400 ;
        RECT 150.450 223.800 152.250 224.400 ;
        RECT 137.550 222.300 145.050 223.500 ;
        RECT 143.250 221.700 145.050 222.300 ;
        RECT 145.950 222.900 152.250 223.800 ;
        RECT 129.150 220.500 130.050 221.400 ;
        RECT 145.950 220.800 146.850 222.900 ;
        RECT 150.450 222.600 152.250 222.900 ;
        RECT 153.150 222.600 155.850 224.400 ;
        RECT 153.150 221.700 154.050 222.600 ;
        RECT 138.450 220.500 146.850 220.800 ;
        RECT 129.150 219.900 146.850 220.500 ;
        RECT 148.950 220.800 154.050 221.700 ;
        RECT 154.950 220.800 157.050 221.700 ;
        RECT 160.650 221.400 162.450 233.400 ;
        RECT 173.700 222.600 175.500 233.400 ;
        RECT 173.700 221.400 177.300 222.600 ;
        RECT 178.800 221.400 180.600 234.000 ;
        RECT 188.700 221.400 190.500 234.000 ;
        RECT 193.800 227.400 195.600 233.400 ;
        RECT 196.800 227.400 198.600 234.000 ;
        RECT 211.800 227.400 213.600 234.000 ;
        RECT 214.800 227.400 216.600 233.400 ;
        RECT 217.800 227.400 219.600 234.000 ;
        RECT 129.150 219.300 140.250 219.900 ;
        RECT 55.950 211.800 58.050 213.900 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 82.950 211.950 85.050 214.050 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 103.950 211.950 106.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 121.950 211.950 124.050 214.050 ;
        RECT 56.100 210.000 57.900 211.800 ;
        RECT 50.100 206.400 57.600 207.300 ;
        RECT 50.100 205.500 51.900 206.400 ;
        RECT 47.400 202.800 50.100 204.600 ;
        RECT 48.300 198.600 50.100 202.800 ;
        RECT 51.300 198.000 53.100 204.600 ;
        RECT 55.800 198.600 57.600 206.400 ;
        RECT 68.700 201.600 69.600 211.950 ;
        RECT 86.400 201.600 87.600 211.950 ;
        RECT 101.400 201.600 102.600 211.950 ;
        RECT 116.100 210.150 117.900 211.950 ;
        RECT 119.850 207.750 121.050 211.950 ;
        RECT 122.100 210.150 123.900 211.950 ;
        RECT 119.850 206.700 123.600 207.750 ;
        RECT 113.400 203.700 121.200 205.050 ;
        RECT 65.400 198.000 67.200 201.600 ;
        RECT 68.400 198.600 70.200 201.600 ;
        RECT 71.400 198.000 73.200 201.600 ;
        RECT 83.400 198.000 85.200 201.600 ;
        RECT 86.400 198.600 88.200 201.600 ;
        RECT 100.800 198.600 102.600 201.600 ;
        RECT 103.800 198.000 105.600 201.600 ;
        RECT 113.400 198.600 115.200 203.700 ;
        RECT 116.400 198.000 118.200 202.800 ;
        RECT 119.400 198.600 121.200 203.700 ;
        RECT 122.400 204.600 123.600 206.700 ;
        RECT 129.150 204.600 130.050 219.300 ;
        RECT 138.450 219.000 140.250 219.300 ;
        RECT 130.950 211.950 133.050 214.050 ;
        RECT 139.950 212.400 142.050 214.050 ;
        RECT 131.100 210.150 132.900 211.950 ;
        RECT 134.100 211.200 142.050 212.400 ;
        RECT 134.100 210.600 135.900 211.200 ;
        RECT 132.000 209.400 132.900 210.150 ;
        RECT 137.100 209.400 138.900 210.000 ;
        RECT 132.000 208.200 138.900 209.400 ;
        RECT 148.950 208.200 149.850 220.800 ;
        RECT 154.950 219.600 159.150 220.800 ;
        RECT 158.250 217.800 160.050 219.600 ;
        RECT 161.250 214.050 162.450 221.400 ;
        RECT 173.100 214.050 174.900 215.850 ;
        RECT 176.400 214.050 177.300 221.400 ;
        RECT 179.100 214.050 180.900 215.850 ;
        RECT 188.100 214.050 189.900 215.850 ;
        RECT 193.950 214.050 195.150 227.400 ;
        RECT 157.950 213.750 162.450 214.050 ;
        RECT 156.150 211.950 162.450 213.750 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 187.950 211.950 190.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 196.950 211.950 199.050 214.050 ;
        RECT 215.400 213.900 216.600 227.400 ;
        RECT 221.550 221.400 223.350 233.400 ;
        RECT 224.550 230.400 226.350 234.000 ;
        RECT 229.050 227.400 230.850 233.400 ;
        RECT 233.250 227.400 235.050 234.000 ;
        RECT 226.950 225.300 230.850 227.400 ;
        RECT 236.850 226.500 238.650 233.400 ;
        RECT 239.850 227.400 241.650 234.000 ;
        RECT 244.650 227.400 246.450 233.400 ;
        RECT 250.050 227.400 251.850 234.000 ;
        RECT 245.250 226.500 246.450 227.400 ;
        RECT 235.950 225.450 242.550 226.500 ;
        RECT 235.950 224.700 237.750 225.450 ;
        RECT 240.750 224.700 242.550 225.450 ;
        RECT 245.250 224.400 250.050 226.500 ;
        RECT 228.150 222.600 230.850 224.400 ;
        RECT 231.750 223.800 233.550 224.400 ;
        RECT 231.750 222.900 238.050 223.800 ;
        RECT 245.250 223.500 246.450 224.400 ;
        RECT 231.750 222.600 233.550 222.900 ;
        RECT 229.950 221.700 230.850 222.600 ;
        RECT 221.550 214.050 222.750 221.400 ;
        RECT 226.950 220.800 229.050 221.700 ;
        RECT 229.950 220.800 235.050 221.700 ;
        RECT 224.850 219.600 229.050 220.800 ;
        RECT 223.950 217.800 225.750 219.600 ;
        RECT 137.850 207.000 149.850 208.200 ;
        RECT 137.850 205.200 138.900 207.000 ;
        RECT 148.050 206.400 149.850 207.000 ;
        RECT 122.400 198.600 124.200 204.600 ;
        RECT 129.150 198.600 130.950 204.600 ;
        RECT 133.950 202.500 136.050 204.600 ;
        RECT 137.550 203.400 139.350 205.200 ;
        RECT 161.250 204.600 162.450 211.950 ;
        RECT 140.850 203.550 142.650 204.300 ;
        RECT 154.950 203.700 157.050 204.600 ;
        RECT 140.850 202.500 145.800 203.550 ;
        RECT 135.000 201.600 136.050 202.500 ;
        RECT 144.750 201.600 145.800 202.500 ;
        RECT 153.300 202.500 157.050 203.700 ;
        RECT 153.300 201.600 154.350 202.500 ;
        RECT 132.150 198.000 133.950 201.600 ;
        RECT 135.000 200.700 138.750 201.600 ;
        RECT 136.950 198.600 138.750 200.700 ;
        RECT 141.450 198.000 143.250 201.600 ;
        RECT 144.750 198.600 146.550 201.600 ;
        RECT 148.350 198.000 150.150 201.600 ;
        RECT 152.550 198.600 154.350 201.600 ;
        RECT 157.350 198.000 159.150 201.600 ;
        RECT 160.650 198.600 162.450 204.600 ;
        RECT 176.400 201.600 177.300 211.950 ;
        RECT 191.100 210.150 192.900 211.950 ;
        RECT 194.850 207.750 196.050 211.950 ;
        RECT 197.100 210.150 198.900 211.950 ;
        RECT 211.950 211.800 214.050 213.900 ;
        RECT 214.950 211.800 217.050 213.900 ;
        RECT 217.950 211.800 220.050 213.900 ;
        RECT 221.550 213.750 226.050 214.050 ;
        RECT 221.550 211.950 227.850 213.750 ;
        RECT 212.100 210.000 213.900 211.800 ;
        RECT 194.850 206.700 198.600 207.750 ;
        RECT 215.400 206.700 216.600 211.800 ;
        RECT 218.100 210.000 219.900 211.800 ;
        RECT 188.400 203.700 196.200 205.050 ;
        RECT 172.800 198.000 174.600 201.600 ;
        RECT 175.800 198.600 177.600 201.600 ;
        RECT 178.800 198.000 180.600 201.600 ;
        RECT 188.400 198.600 190.200 203.700 ;
        RECT 191.400 198.000 193.200 202.800 ;
        RECT 194.400 198.600 196.200 203.700 ;
        RECT 197.400 204.600 198.600 206.700 ;
        RECT 212.400 205.800 216.600 206.700 ;
        RECT 197.400 198.600 199.200 204.600 ;
        RECT 212.400 198.600 214.200 205.800 ;
        RECT 221.550 204.600 222.750 211.950 ;
        RECT 234.150 208.200 235.050 220.800 ;
        RECT 237.150 220.800 238.050 222.900 ;
        RECT 238.950 222.300 246.450 223.500 ;
        RECT 238.950 221.700 240.750 222.300 ;
        RECT 253.050 221.400 254.850 233.400 ;
        RECT 265.800 222.600 267.600 233.400 ;
        RECT 265.800 221.400 270.900 222.600 ;
        RECT 273.300 222.300 275.100 233.400 ;
        RECT 280.800 222.300 282.600 233.400 ;
        RECT 292.800 227.400 294.600 234.000 ;
        RECT 295.800 227.400 297.600 233.400 ;
        RECT 298.800 227.400 300.600 234.000 ;
        RECT 311.400 227.400 313.200 234.000 ;
        RECT 314.400 227.400 316.200 233.400 ;
        RECT 237.150 220.500 245.550 220.800 ;
        RECT 253.950 220.500 254.850 221.400 ;
        RECT 268.800 220.500 270.900 221.400 ;
        RECT 271.800 221.400 275.100 222.300 ;
        RECT 237.150 219.900 254.850 220.500 ;
        RECT 243.750 219.300 254.850 219.900 ;
        RECT 243.750 219.000 245.550 219.300 ;
        RECT 241.950 212.400 244.050 214.050 ;
        RECT 241.950 211.200 249.900 212.400 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 248.100 210.600 249.900 211.200 ;
        RECT 251.100 210.150 252.900 211.950 ;
        RECT 245.100 209.400 246.900 210.000 ;
        RECT 251.100 209.400 252.000 210.150 ;
        RECT 245.100 208.200 252.000 209.400 ;
        RECT 234.150 207.000 246.150 208.200 ;
        RECT 234.150 206.400 235.950 207.000 ;
        RECT 245.100 205.200 246.150 207.000 ;
        RECT 217.500 198.000 219.300 204.600 ;
        RECT 221.550 198.600 223.350 204.600 ;
        RECT 226.950 203.700 229.050 204.600 ;
        RECT 226.950 202.500 230.700 203.700 ;
        RECT 241.350 203.550 243.150 204.300 ;
        RECT 229.650 201.600 230.700 202.500 ;
        RECT 238.200 202.500 243.150 203.550 ;
        RECT 244.650 203.400 246.450 205.200 ;
        RECT 253.950 204.600 254.850 219.300 ;
        RECT 262.950 216.450 267.000 217.050 ;
        RECT 271.800 216.900 273.000 221.400 ;
        RECT 277.800 221.100 282.600 222.300 ;
        RECT 277.800 220.200 279.900 221.100 ;
        RECT 274.650 219.300 279.900 220.200 ;
        RECT 274.650 217.200 276.450 219.300 ;
        RECT 262.950 215.700 267.450 216.450 ;
        RECT 271.650 216.300 273.750 216.900 ;
        RECT 262.950 214.950 267.900 215.700 ;
        RECT 266.100 213.900 267.900 214.950 ;
        RECT 271.650 214.800 274.650 216.300 ;
        RECT 265.950 211.800 268.050 213.900 ;
        RECT 270.900 212.100 272.700 213.900 ;
        RECT 270.750 210.000 272.850 212.100 ;
        RECT 273.750 208.200 274.650 214.800 ;
        RECT 276.000 214.200 277.800 216.000 ;
        RECT 275.700 212.100 277.800 214.200 ;
        RECT 296.400 213.900 297.600 227.400 ;
        RECT 314.850 214.050 316.050 227.400 ;
        RECT 319.500 221.400 321.300 234.000 ;
        RECT 324.150 221.400 325.950 233.400 ;
        RECT 327.150 227.400 328.950 234.000 ;
        RECT 332.550 227.400 334.350 233.400 ;
        RECT 337.350 227.400 339.150 234.000 ;
        RECT 332.550 226.500 333.750 227.400 ;
        RECT 340.350 226.500 342.150 233.400 ;
        RECT 343.950 227.400 345.750 234.000 ;
        RECT 348.150 227.400 349.950 233.400 ;
        RECT 352.650 230.400 354.450 234.000 ;
        RECT 328.950 224.400 333.750 226.500 ;
        RECT 336.450 225.450 343.050 226.500 ;
        RECT 336.450 224.700 338.250 225.450 ;
        RECT 341.250 224.700 343.050 225.450 ;
        RECT 348.150 225.300 352.050 227.400 ;
        RECT 332.550 223.500 333.750 224.400 ;
        RECT 345.450 223.800 347.250 224.400 ;
        RECT 332.550 222.300 340.050 223.500 ;
        RECT 338.250 221.700 340.050 222.300 ;
        RECT 340.950 222.900 347.250 223.800 ;
        RECT 324.150 220.500 325.050 221.400 ;
        RECT 340.950 220.800 341.850 222.900 ;
        RECT 345.450 222.600 347.250 222.900 ;
        RECT 348.150 222.600 350.850 224.400 ;
        RECT 348.150 221.700 349.050 222.600 ;
        RECT 333.450 220.500 341.850 220.800 ;
        RECT 324.150 219.900 341.850 220.500 ;
        RECT 343.950 220.800 349.050 221.700 ;
        RECT 349.950 220.800 352.050 221.700 ;
        RECT 355.650 221.400 357.450 233.400 ;
        RECT 324.150 219.300 335.250 219.900 ;
        RECT 320.100 214.050 321.900 215.850 ;
        RECT 280.950 211.800 283.050 213.900 ;
        RECT 292.950 211.800 295.050 213.900 ;
        RECT 295.950 211.800 298.050 213.900 ;
        RECT 298.950 211.800 301.050 213.900 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 280.950 211.200 282.750 211.800 ;
        RECT 275.700 210.000 282.750 211.200 ;
        RECT 293.100 210.000 294.900 211.800 ;
        RECT 275.700 209.100 277.800 210.000 ;
        RECT 268.200 205.500 270.300 207.900 ;
        RECT 271.650 206.100 274.650 208.200 ;
        RECT 275.550 207.300 277.350 209.100 ;
        RECT 247.950 202.500 250.050 204.600 ;
        RECT 238.200 201.600 239.250 202.500 ;
        RECT 247.950 201.600 249.000 202.500 ;
        RECT 224.850 198.000 226.650 201.600 ;
        RECT 229.650 198.600 231.450 201.600 ;
        RECT 233.850 198.000 235.650 201.600 ;
        RECT 237.450 198.600 239.250 201.600 ;
        RECT 240.750 198.000 242.550 201.600 ;
        RECT 245.250 200.700 249.000 201.600 ;
        RECT 245.250 198.600 247.050 200.700 ;
        RECT 250.050 198.000 251.850 201.600 ;
        RECT 253.050 198.600 254.850 204.600 ;
        RECT 265.800 204.600 270.300 205.500 ;
        RECT 265.800 198.600 267.600 204.600 ;
        RECT 273.750 204.000 274.650 206.100 ;
        RECT 278.250 207.000 280.350 207.600 ;
        RECT 278.250 205.500 282.600 207.000 ;
        RECT 296.400 206.700 297.600 211.800 ;
        RECT 299.100 210.000 300.900 211.800 ;
        RECT 311.100 210.150 312.900 211.950 ;
        RECT 313.950 207.750 315.150 211.950 ;
        RECT 317.100 210.150 318.900 211.950 ;
        RECT 281.100 204.600 282.600 205.500 ;
        RECT 273.600 198.600 275.400 204.000 ;
        RECT 280.800 198.600 282.600 204.600 ;
        RECT 293.400 205.800 297.600 206.700 ;
        RECT 311.400 206.700 315.150 207.750 ;
        RECT 293.400 198.600 295.200 205.800 ;
        RECT 311.400 204.600 312.600 206.700 ;
        RECT 298.500 198.000 300.300 204.600 ;
        RECT 310.800 198.600 312.600 204.600 ;
        RECT 313.800 203.700 321.600 205.050 ;
        RECT 313.800 198.600 315.600 203.700 ;
        RECT 316.800 198.000 318.600 202.800 ;
        RECT 319.800 198.600 321.600 203.700 ;
        RECT 324.150 204.600 325.050 219.300 ;
        RECT 333.450 219.000 335.250 219.300 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 334.950 212.400 337.050 214.050 ;
        RECT 326.100 210.150 327.900 211.950 ;
        RECT 329.100 211.200 337.050 212.400 ;
        RECT 329.100 210.600 330.900 211.200 ;
        RECT 327.000 209.400 327.900 210.150 ;
        RECT 332.100 209.400 333.900 210.000 ;
        RECT 327.000 208.200 333.900 209.400 ;
        RECT 343.950 208.200 344.850 220.800 ;
        RECT 349.950 219.600 354.150 220.800 ;
        RECT 353.250 217.800 355.050 219.600 ;
        RECT 356.250 214.050 357.450 221.400 ;
        RECT 352.950 213.750 357.450 214.050 ;
        RECT 351.150 211.950 357.450 213.750 ;
        RECT 332.850 207.000 344.850 208.200 ;
        RECT 332.850 205.200 333.900 207.000 ;
        RECT 343.050 206.400 344.850 207.000 ;
        RECT 324.150 198.600 325.950 204.600 ;
        RECT 328.950 202.500 331.050 204.600 ;
        RECT 332.550 203.400 334.350 205.200 ;
        RECT 356.250 204.600 357.450 211.950 ;
        RECT 335.850 203.550 337.650 204.300 ;
        RECT 349.950 203.700 352.050 204.600 ;
        RECT 335.850 202.500 340.800 203.550 ;
        RECT 330.000 201.600 331.050 202.500 ;
        RECT 339.750 201.600 340.800 202.500 ;
        RECT 348.300 202.500 352.050 203.700 ;
        RECT 348.300 201.600 349.350 202.500 ;
        RECT 327.150 198.000 328.950 201.600 ;
        RECT 330.000 200.700 333.750 201.600 ;
        RECT 331.950 198.600 333.750 200.700 ;
        RECT 336.450 198.000 338.250 201.600 ;
        RECT 339.750 198.600 341.550 201.600 ;
        RECT 343.350 198.000 345.150 201.600 ;
        RECT 347.550 198.600 349.350 201.600 ;
        RECT 352.350 198.000 354.150 201.600 ;
        RECT 355.650 198.600 357.450 204.600 ;
        RECT 360.150 221.400 361.950 233.400 ;
        RECT 363.150 227.400 364.950 234.000 ;
        RECT 368.550 227.400 370.350 233.400 ;
        RECT 373.350 227.400 375.150 234.000 ;
        RECT 368.550 226.500 369.750 227.400 ;
        RECT 376.350 226.500 378.150 233.400 ;
        RECT 379.950 227.400 381.750 234.000 ;
        RECT 384.150 227.400 385.950 233.400 ;
        RECT 388.650 230.400 390.450 234.000 ;
        RECT 364.950 224.400 369.750 226.500 ;
        RECT 372.450 225.450 379.050 226.500 ;
        RECT 372.450 224.700 374.250 225.450 ;
        RECT 377.250 224.700 379.050 225.450 ;
        RECT 384.150 225.300 388.050 227.400 ;
        RECT 368.550 223.500 369.750 224.400 ;
        RECT 381.450 223.800 383.250 224.400 ;
        RECT 368.550 222.300 376.050 223.500 ;
        RECT 374.250 221.700 376.050 222.300 ;
        RECT 376.950 222.900 383.250 223.800 ;
        RECT 360.150 220.500 361.050 221.400 ;
        RECT 376.950 220.800 377.850 222.900 ;
        RECT 381.450 222.600 383.250 222.900 ;
        RECT 384.150 222.600 386.850 224.400 ;
        RECT 384.150 221.700 385.050 222.600 ;
        RECT 369.450 220.500 377.850 220.800 ;
        RECT 360.150 219.900 377.850 220.500 ;
        RECT 379.950 220.800 385.050 221.700 ;
        RECT 385.950 220.800 388.050 221.700 ;
        RECT 391.650 221.400 393.450 233.400 ;
        RECT 404.700 222.600 406.500 233.400 ;
        RECT 404.700 221.400 408.300 222.600 ;
        RECT 409.800 221.400 411.600 234.000 ;
        RECT 419.400 222.300 421.200 233.400 ;
        RECT 422.400 223.200 424.200 234.000 ;
        RECT 425.400 222.300 427.200 233.400 ;
        RECT 419.400 221.400 427.200 222.300 ;
        RECT 428.400 221.400 430.200 233.400 ;
        RECT 434.550 221.400 436.350 233.400 ;
        RECT 437.550 230.400 439.350 234.000 ;
        RECT 442.050 227.400 443.850 233.400 ;
        RECT 446.250 227.400 448.050 234.000 ;
        RECT 439.950 225.300 443.850 227.400 ;
        RECT 449.850 226.500 451.650 233.400 ;
        RECT 452.850 227.400 454.650 234.000 ;
        RECT 457.650 227.400 459.450 233.400 ;
        RECT 463.050 227.400 464.850 234.000 ;
        RECT 458.250 226.500 459.450 227.400 ;
        RECT 448.950 225.450 455.550 226.500 ;
        RECT 448.950 224.700 450.750 225.450 ;
        RECT 453.750 224.700 455.550 225.450 ;
        RECT 458.250 224.400 463.050 226.500 ;
        RECT 441.150 222.600 443.850 224.400 ;
        RECT 444.750 223.800 446.550 224.400 ;
        RECT 444.750 222.900 451.050 223.800 ;
        RECT 458.250 223.500 459.450 224.400 ;
        RECT 444.750 222.600 446.550 222.900 ;
        RECT 442.950 221.700 443.850 222.600 ;
        RECT 360.150 219.300 371.250 219.900 ;
        RECT 360.150 204.600 361.050 219.300 ;
        RECT 369.450 219.000 371.250 219.300 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 370.950 212.400 373.050 214.050 ;
        RECT 362.100 210.150 363.900 211.950 ;
        RECT 365.100 211.200 373.050 212.400 ;
        RECT 365.100 210.600 366.900 211.200 ;
        RECT 363.000 209.400 363.900 210.150 ;
        RECT 368.100 209.400 369.900 210.000 ;
        RECT 363.000 208.200 369.900 209.400 ;
        RECT 379.950 208.200 380.850 220.800 ;
        RECT 385.950 219.600 390.150 220.800 ;
        RECT 389.250 217.800 391.050 219.600 ;
        RECT 392.250 214.050 393.450 221.400 ;
        RECT 404.100 214.050 405.900 215.850 ;
        RECT 407.400 214.050 408.300 221.400 ;
        RECT 410.100 214.050 411.900 215.850 ;
        RECT 388.950 213.750 393.450 214.050 ;
        RECT 387.150 211.950 393.450 213.750 ;
        RECT 403.950 211.950 406.050 214.050 ;
        RECT 406.950 211.950 409.050 214.050 ;
        RECT 409.950 211.950 412.050 214.050 ;
        RECT 422.100 213.900 423.900 215.700 ;
        RECT 428.700 213.900 429.600 221.400 ;
        RECT 434.550 214.050 435.750 221.400 ;
        RECT 439.950 220.800 442.050 221.700 ;
        RECT 442.950 220.800 448.050 221.700 ;
        RECT 437.850 219.600 442.050 220.800 ;
        RECT 436.950 217.800 438.750 219.600 ;
        RECT 368.850 207.000 380.850 208.200 ;
        RECT 368.850 205.200 369.900 207.000 ;
        RECT 379.050 206.400 380.850 207.000 ;
        RECT 360.150 198.600 361.950 204.600 ;
        RECT 364.950 202.500 367.050 204.600 ;
        RECT 368.550 203.400 370.350 205.200 ;
        RECT 392.250 204.600 393.450 211.950 ;
        RECT 371.850 203.550 373.650 204.300 ;
        RECT 385.950 203.700 388.050 204.600 ;
        RECT 371.850 202.500 376.800 203.550 ;
        RECT 366.000 201.600 367.050 202.500 ;
        RECT 375.750 201.600 376.800 202.500 ;
        RECT 384.300 202.500 388.050 203.700 ;
        RECT 384.300 201.600 385.350 202.500 ;
        RECT 363.150 198.000 364.950 201.600 ;
        RECT 366.000 200.700 369.750 201.600 ;
        RECT 367.950 198.600 369.750 200.700 ;
        RECT 372.450 198.000 374.250 201.600 ;
        RECT 375.750 198.600 377.550 201.600 ;
        RECT 379.350 198.000 381.150 201.600 ;
        RECT 383.550 198.600 385.350 201.600 ;
        RECT 388.350 198.000 390.150 201.600 ;
        RECT 391.650 198.600 393.450 204.600 ;
        RECT 407.400 201.600 408.300 211.950 ;
        RECT 418.950 211.800 421.050 213.900 ;
        RECT 421.950 211.800 424.050 213.900 ;
        RECT 424.950 211.800 427.050 213.900 ;
        RECT 427.950 211.800 430.050 213.900 ;
        RECT 434.550 213.750 439.050 214.050 ;
        RECT 434.550 211.950 440.850 213.750 ;
        RECT 419.100 210.000 420.900 211.800 ;
        RECT 425.100 210.000 426.900 211.800 ;
        RECT 428.700 204.600 429.600 211.800 ;
        RECT 403.800 198.000 405.600 201.600 ;
        RECT 406.800 198.600 408.600 201.600 ;
        RECT 409.800 198.000 411.600 201.600 ;
        RECT 420.000 198.000 421.800 204.600 ;
        RECT 424.500 203.400 429.600 204.600 ;
        RECT 434.550 204.600 435.750 211.950 ;
        RECT 447.150 208.200 448.050 220.800 ;
        RECT 450.150 220.800 451.050 222.900 ;
        RECT 451.950 222.300 459.450 223.500 ;
        RECT 451.950 221.700 453.750 222.300 ;
        RECT 466.050 221.400 467.850 233.400 ;
        RECT 476.400 221.400 478.200 234.000 ;
        RECT 450.150 220.500 458.550 220.800 ;
        RECT 466.950 220.500 467.850 221.400 ;
        RECT 450.150 219.900 467.850 220.500 ;
        RECT 456.750 219.300 467.850 219.900 ;
        RECT 479.400 220.500 481.200 233.400 ;
        RECT 482.400 221.400 484.200 234.000 ;
        RECT 485.400 220.500 487.200 233.400 ;
        RECT 488.400 221.400 490.200 234.000 ;
        RECT 491.400 220.500 493.200 233.400 ;
        RECT 494.400 221.400 496.200 234.000 ;
        RECT 497.400 220.500 499.200 233.400 ;
        RECT 500.400 221.400 502.200 234.000 ;
        RECT 512.400 222.300 514.200 233.400 ;
        RECT 515.400 223.200 517.200 234.000 ;
        RECT 518.400 222.300 520.200 233.400 ;
        RECT 512.400 221.400 520.200 222.300 ;
        RECT 521.400 221.400 523.200 233.400 ;
        RECT 536.700 222.600 538.500 233.400 ;
        RECT 536.700 221.400 540.300 222.600 ;
        RECT 541.800 221.400 543.600 234.000 ;
        RECT 551.400 222.300 553.200 233.400 ;
        RECT 554.400 223.200 556.200 234.000 ;
        RECT 557.400 222.300 559.200 233.400 ;
        RECT 551.400 221.400 559.200 222.300 ;
        RECT 560.400 221.400 562.200 233.400 ;
        RECT 567.150 221.400 568.950 233.400 ;
        RECT 570.150 227.400 571.950 234.000 ;
        RECT 575.550 227.400 577.350 233.400 ;
        RECT 580.350 227.400 582.150 234.000 ;
        RECT 575.550 226.500 576.750 227.400 ;
        RECT 583.350 226.500 585.150 233.400 ;
        RECT 586.950 227.400 588.750 234.000 ;
        RECT 591.150 227.400 592.950 233.400 ;
        RECT 595.650 230.400 597.450 234.000 ;
        RECT 571.950 224.400 576.750 226.500 ;
        RECT 579.450 225.450 586.050 226.500 ;
        RECT 579.450 224.700 581.250 225.450 ;
        RECT 584.250 224.700 586.050 225.450 ;
        RECT 591.150 225.300 595.050 227.400 ;
        RECT 575.550 223.500 576.750 224.400 ;
        RECT 588.450 223.800 590.250 224.400 ;
        RECT 575.550 222.300 583.050 223.500 ;
        RECT 581.250 221.700 583.050 222.300 ;
        RECT 583.950 222.900 590.250 223.800 ;
        RECT 479.400 219.300 483.300 220.500 ;
        RECT 485.400 219.300 489.300 220.500 ;
        RECT 491.400 219.300 495.300 220.500 ;
        RECT 497.400 219.300 500.100 220.500 ;
        RECT 456.750 219.000 458.550 219.300 ;
        RECT 454.950 212.400 457.050 214.050 ;
        RECT 454.950 211.200 462.900 212.400 ;
        RECT 463.950 211.950 466.050 214.050 ;
        RECT 461.100 210.600 462.900 211.200 ;
        RECT 464.100 210.150 465.900 211.950 ;
        RECT 458.100 209.400 459.900 210.000 ;
        RECT 464.100 209.400 465.000 210.150 ;
        RECT 458.100 208.200 465.000 209.400 ;
        RECT 447.150 207.000 459.150 208.200 ;
        RECT 447.150 206.400 448.950 207.000 ;
        RECT 458.100 205.200 459.150 207.000 ;
        RECT 424.500 198.600 426.300 203.400 ;
        RECT 427.500 198.000 429.300 201.600 ;
        RECT 434.550 198.600 436.350 204.600 ;
        RECT 439.950 203.700 442.050 204.600 ;
        RECT 439.950 202.500 443.700 203.700 ;
        RECT 454.350 203.550 456.150 204.300 ;
        RECT 442.650 201.600 443.700 202.500 ;
        RECT 451.200 202.500 456.150 203.550 ;
        RECT 457.650 203.400 459.450 205.200 ;
        RECT 466.950 204.600 467.850 219.300 ;
        RECT 478.950 211.800 481.050 213.900 ;
        RECT 479.100 210.000 480.900 211.800 ;
        RECT 482.100 208.800 483.300 219.300 ;
        RECT 484.500 208.800 486.300 209.400 ;
        RECT 482.100 207.600 486.300 208.800 ;
        RECT 488.100 208.800 489.300 219.300 ;
        RECT 490.500 208.800 492.300 209.400 ;
        RECT 488.100 207.600 492.300 208.800 ;
        RECT 494.100 208.800 495.300 219.300 ;
        RECT 499.200 213.900 500.100 219.300 ;
        RECT 515.100 213.900 516.900 215.700 ;
        RECT 521.700 213.900 522.600 221.400 ;
        RECT 536.100 214.050 537.900 215.850 ;
        RECT 539.400 214.050 540.300 221.400 ;
        RECT 542.100 214.050 543.900 215.850 ;
        RECT 499.200 211.800 502.050 213.900 ;
        RECT 511.950 211.800 514.050 213.900 ;
        RECT 514.950 211.800 517.050 213.900 ;
        RECT 517.950 211.800 520.050 213.900 ;
        RECT 520.950 211.800 523.050 213.900 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 538.950 211.950 541.050 214.050 ;
        RECT 541.950 211.950 544.050 214.050 ;
        RECT 554.100 213.900 555.900 215.700 ;
        RECT 560.700 213.900 561.600 221.400 ;
        RECT 567.150 220.500 568.050 221.400 ;
        RECT 583.950 220.800 584.850 222.900 ;
        RECT 588.450 222.600 590.250 222.900 ;
        RECT 591.150 222.600 593.850 224.400 ;
        RECT 591.150 221.700 592.050 222.600 ;
        RECT 576.450 220.500 584.850 220.800 ;
        RECT 567.150 219.900 584.850 220.500 ;
        RECT 586.950 220.800 592.050 221.700 ;
        RECT 592.950 220.800 595.050 221.700 ;
        RECT 598.650 221.400 600.450 233.400 ;
        RECT 608.400 221.400 610.200 234.000 ;
        RECT 613.500 222.600 615.300 233.400 ;
        RECT 611.700 221.400 615.300 222.600 ;
        RECT 621.150 221.400 622.950 233.400 ;
        RECT 624.150 227.400 625.950 234.000 ;
        RECT 629.550 227.400 631.350 233.400 ;
        RECT 634.350 227.400 636.150 234.000 ;
        RECT 629.550 226.500 630.750 227.400 ;
        RECT 637.350 226.500 639.150 233.400 ;
        RECT 640.950 227.400 642.750 234.000 ;
        RECT 645.150 227.400 646.950 233.400 ;
        RECT 649.650 230.400 651.450 234.000 ;
        RECT 625.950 224.400 630.750 226.500 ;
        RECT 633.450 225.450 640.050 226.500 ;
        RECT 633.450 224.700 635.250 225.450 ;
        RECT 638.250 224.700 640.050 225.450 ;
        RECT 645.150 225.300 649.050 227.400 ;
        RECT 629.550 223.500 630.750 224.400 ;
        RECT 642.450 223.800 644.250 224.400 ;
        RECT 629.550 222.300 637.050 223.500 ;
        RECT 635.250 221.700 637.050 222.300 ;
        RECT 637.950 222.900 644.250 223.800 ;
        RECT 567.150 219.300 578.250 219.900 ;
        RECT 496.500 208.800 498.300 209.400 ;
        RECT 494.100 207.600 498.300 208.800 ;
        RECT 482.100 206.700 483.300 207.600 ;
        RECT 488.100 206.700 489.300 207.600 ;
        RECT 494.100 206.700 495.300 207.600 ;
        RECT 499.200 206.700 500.100 211.800 ;
        RECT 512.100 210.000 513.900 211.800 ;
        RECT 518.100 210.000 519.900 211.800 ;
        RECT 479.400 205.500 483.300 206.700 ;
        RECT 485.400 205.500 489.300 206.700 ;
        RECT 491.400 205.500 495.300 206.700 ;
        RECT 497.400 205.500 500.100 206.700 ;
        RECT 460.950 202.500 463.050 204.600 ;
        RECT 451.200 201.600 452.250 202.500 ;
        RECT 460.950 201.600 462.000 202.500 ;
        RECT 437.850 198.000 439.650 201.600 ;
        RECT 442.650 198.600 444.450 201.600 ;
        RECT 446.850 198.000 448.650 201.600 ;
        RECT 450.450 198.600 452.250 201.600 ;
        RECT 453.750 198.000 455.550 201.600 ;
        RECT 458.250 200.700 462.000 201.600 ;
        RECT 458.250 198.600 460.050 200.700 ;
        RECT 463.050 198.000 464.850 201.600 ;
        RECT 466.050 198.600 467.850 204.600 ;
        RECT 476.400 198.000 478.200 204.600 ;
        RECT 479.400 198.600 481.200 205.500 ;
        RECT 482.400 198.000 484.200 204.600 ;
        RECT 485.400 198.600 487.200 205.500 ;
        RECT 488.400 198.000 490.200 204.600 ;
        RECT 491.400 198.600 493.200 205.500 ;
        RECT 494.400 198.000 496.200 204.600 ;
        RECT 497.400 198.600 499.200 205.500 ;
        RECT 521.700 204.600 522.600 211.800 ;
        RECT 500.400 198.000 502.200 204.600 ;
        RECT 513.000 198.000 514.800 204.600 ;
        RECT 517.500 203.400 522.600 204.600 ;
        RECT 517.500 198.600 519.300 203.400 ;
        RECT 539.400 201.600 540.300 211.950 ;
        RECT 550.950 211.800 553.050 213.900 ;
        RECT 553.950 211.800 556.050 213.900 ;
        RECT 556.950 211.800 559.050 213.900 ;
        RECT 559.950 211.800 562.050 213.900 ;
        RECT 551.100 210.000 552.900 211.800 ;
        RECT 557.100 210.000 558.900 211.800 ;
        RECT 560.700 204.600 561.600 211.800 ;
        RECT 520.500 198.000 522.300 201.600 ;
        RECT 535.800 198.000 537.600 201.600 ;
        RECT 538.800 198.600 540.600 201.600 ;
        RECT 541.800 198.000 543.600 201.600 ;
        RECT 552.000 198.000 553.800 204.600 ;
        RECT 556.500 203.400 561.600 204.600 ;
        RECT 567.150 204.600 568.050 219.300 ;
        RECT 576.450 219.000 578.250 219.300 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 577.950 212.400 580.050 214.050 ;
        RECT 569.100 210.150 570.900 211.950 ;
        RECT 572.100 211.200 580.050 212.400 ;
        RECT 572.100 210.600 573.900 211.200 ;
        RECT 570.000 209.400 570.900 210.150 ;
        RECT 575.100 209.400 576.900 210.000 ;
        RECT 570.000 208.200 576.900 209.400 ;
        RECT 586.950 208.200 587.850 220.800 ;
        RECT 592.950 219.600 597.150 220.800 ;
        RECT 596.250 217.800 598.050 219.600 ;
        RECT 599.250 214.050 600.450 221.400 ;
        RECT 608.100 214.050 609.900 215.850 ;
        RECT 611.700 214.050 612.600 221.400 ;
        RECT 621.150 220.500 622.050 221.400 ;
        RECT 637.950 220.800 638.850 222.900 ;
        RECT 642.450 222.600 644.250 222.900 ;
        RECT 645.150 222.600 647.850 224.400 ;
        RECT 645.150 221.700 646.050 222.600 ;
        RECT 630.450 220.500 638.850 220.800 ;
        RECT 621.150 219.900 638.850 220.500 ;
        RECT 640.950 220.800 646.050 221.700 ;
        RECT 646.950 220.800 649.050 221.700 ;
        RECT 652.650 221.400 654.450 233.400 ;
        RECT 662.400 227.400 664.200 234.000 ;
        RECT 665.400 227.400 667.200 233.400 ;
        RECT 668.400 227.400 670.200 234.000 ;
        RECT 683.400 227.400 685.200 234.000 ;
        RECT 686.400 227.400 688.200 233.400 ;
        RECT 621.150 219.300 632.250 219.900 ;
        RECT 614.100 214.050 615.900 215.850 ;
        RECT 595.950 213.750 600.450 214.050 ;
        RECT 594.150 211.950 600.450 213.750 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 613.950 211.950 616.050 214.050 ;
        RECT 575.850 207.000 587.850 208.200 ;
        RECT 575.850 205.200 576.900 207.000 ;
        RECT 586.050 206.400 587.850 207.000 ;
        RECT 556.500 198.600 558.300 203.400 ;
        RECT 559.500 198.000 561.300 201.600 ;
        RECT 567.150 198.600 568.950 204.600 ;
        RECT 571.950 202.500 574.050 204.600 ;
        RECT 575.550 203.400 577.350 205.200 ;
        RECT 599.250 204.600 600.450 211.950 ;
        RECT 578.850 203.550 580.650 204.300 ;
        RECT 592.950 203.700 595.050 204.600 ;
        RECT 578.850 202.500 583.800 203.550 ;
        RECT 573.000 201.600 574.050 202.500 ;
        RECT 582.750 201.600 583.800 202.500 ;
        RECT 591.300 202.500 595.050 203.700 ;
        RECT 591.300 201.600 592.350 202.500 ;
        RECT 570.150 198.000 571.950 201.600 ;
        RECT 573.000 200.700 576.750 201.600 ;
        RECT 574.950 198.600 576.750 200.700 ;
        RECT 579.450 198.000 581.250 201.600 ;
        RECT 582.750 198.600 584.550 201.600 ;
        RECT 586.350 198.000 588.150 201.600 ;
        RECT 590.550 198.600 592.350 201.600 ;
        RECT 595.350 198.000 597.150 201.600 ;
        RECT 598.650 198.600 600.450 204.600 ;
        RECT 611.700 201.600 612.600 211.950 ;
        RECT 621.150 204.600 622.050 219.300 ;
        RECT 630.450 219.000 632.250 219.300 ;
        RECT 622.950 211.950 625.050 214.050 ;
        RECT 631.950 212.400 634.050 214.050 ;
        RECT 623.100 210.150 624.900 211.950 ;
        RECT 626.100 211.200 634.050 212.400 ;
        RECT 626.100 210.600 627.900 211.200 ;
        RECT 624.000 209.400 624.900 210.150 ;
        RECT 629.100 209.400 630.900 210.000 ;
        RECT 624.000 208.200 630.900 209.400 ;
        RECT 640.950 208.200 641.850 220.800 ;
        RECT 646.950 219.600 651.150 220.800 ;
        RECT 650.250 217.800 652.050 219.600 ;
        RECT 653.250 214.050 654.450 221.400 ;
        RECT 649.950 213.750 654.450 214.050 ;
        RECT 665.400 213.900 666.600 227.400 ;
        RECT 678.000 216.450 682.050 217.050 ;
        RECT 677.550 214.950 682.050 216.450 ;
        RECT 648.150 211.950 654.450 213.750 ;
        RECT 629.850 207.000 641.850 208.200 ;
        RECT 629.850 205.200 630.900 207.000 ;
        RECT 640.050 206.400 641.850 207.000 ;
        RECT 608.400 198.000 610.200 201.600 ;
        RECT 611.400 198.600 613.200 201.600 ;
        RECT 614.400 198.000 616.200 201.600 ;
        RECT 621.150 198.600 622.950 204.600 ;
        RECT 625.950 202.500 628.050 204.600 ;
        RECT 629.550 203.400 631.350 205.200 ;
        RECT 653.250 204.600 654.450 211.950 ;
        RECT 661.950 211.800 664.050 213.900 ;
        RECT 664.950 211.800 667.050 213.900 ;
        RECT 667.950 211.800 670.050 213.900 ;
        RECT 662.100 210.000 663.900 211.800 ;
        RECT 665.400 206.700 666.600 211.800 ;
        RECT 668.100 210.000 669.900 211.800 ;
        RECT 677.550 211.050 678.450 214.950 ;
        RECT 686.850 214.050 688.050 227.400 ;
        RECT 691.500 221.400 693.300 234.000 ;
        RECT 703.800 227.400 705.600 234.000 ;
        RECT 706.800 227.400 708.600 233.400 ;
        RECT 709.800 227.400 711.600 234.000 ;
        RECT 692.100 214.050 693.900 215.850 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 691.950 211.950 694.050 214.050 ;
        RECT 707.400 213.900 708.600 227.400 ;
        RECT 719.400 222.300 721.200 233.400 ;
        RECT 719.400 221.400 723.900 222.300 ;
        RECT 726.900 221.400 728.700 233.400 ;
        RECT 734.400 222.600 736.200 233.400 ;
        RECT 721.800 219.300 723.900 221.400 ;
        RECT 727.500 219.900 728.700 221.400 ;
        RECT 731.400 221.400 736.200 222.600 ;
        RECT 746.400 227.400 748.200 233.400 ;
        RECT 749.400 227.400 751.200 234.000 ;
        RECT 731.400 220.500 733.500 221.400 ;
        RECT 746.400 220.500 747.600 227.400 ;
        RECT 752.400 221.400 754.200 233.400 ;
        RECT 766.800 227.400 768.600 233.400 ;
        RECT 769.800 227.400 771.600 234.000 ;
        RECT 727.500 219.000 729.000 219.900 ;
        RECT 746.400 219.600 752.100 220.500 ;
        RECT 724.950 217.500 727.050 217.800 ;
        RECT 723.300 215.700 727.050 217.500 ;
        RECT 728.100 216.900 729.000 219.000 ;
        RECT 750.150 218.700 752.100 219.600 ;
        RECT 727.950 214.800 730.050 216.900 ;
        RECT 735.000 216.450 739.050 217.050 ;
        RECT 734.550 215.700 739.050 216.450 ;
        RECT 734.100 214.950 739.050 215.700 ;
        RECT 724.500 213.900 726.300 214.500 ;
        RECT 677.550 209.550 682.050 211.050 ;
        RECT 683.100 210.150 684.900 211.950 ;
        RECT 678.000 208.950 682.050 209.550 ;
        RECT 685.950 207.750 687.150 211.950 ;
        RECT 689.100 210.150 690.900 211.950 ;
        RECT 703.950 211.800 706.050 213.900 ;
        RECT 706.950 211.800 709.050 213.900 ;
        RECT 709.950 211.800 712.050 213.900 ;
        RECT 718.950 212.700 726.300 213.900 ;
        RECT 727.200 213.900 729.600 214.800 ;
        RECT 734.100 213.900 735.900 214.950 ;
        RECT 746.100 214.050 747.900 215.850 ;
        RECT 718.950 211.800 721.050 212.700 ;
        RECT 704.100 210.000 705.900 211.800 ;
        RECT 683.400 206.700 687.150 207.750 ;
        RECT 707.400 206.700 708.600 211.800 ;
        RECT 710.100 210.000 711.900 211.800 ;
        RECT 719.250 210.000 721.050 211.800 ;
        RECT 724.500 209.400 726.300 211.200 ;
        RECT 724.200 207.300 726.300 209.400 ;
        RECT 665.400 205.800 669.600 206.700 ;
        RECT 632.850 203.550 634.650 204.300 ;
        RECT 646.950 203.700 649.050 204.600 ;
        RECT 632.850 202.500 637.800 203.550 ;
        RECT 627.000 201.600 628.050 202.500 ;
        RECT 636.750 201.600 637.800 202.500 ;
        RECT 645.300 202.500 649.050 203.700 ;
        RECT 645.300 201.600 646.350 202.500 ;
        RECT 624.150 198.000 625.950 201.600 ;
        RECT 627.000 200.700 630.750 201.600 ;
        RECT 628.950 198.600 630.750 200.700 ;
        RECT 633.450 198.000 635.250 201.600 ;
        RECT 636.750 198.600 638.550 201.600 ;
        RECT 640.350 198.000 642.150 201.600 ;
        RECT 644.550 198.600 646.350 201.600 ;
        RECT 649.350 198.000 651.150 201.600 ;
        RECT 652.650 198.600 654.450 204.600 ;
        RECT 662.700 198.000 664.500 204.600 ;
        RECT 667.800 198.600 669.600 205.800 ;
        RECT 683.400 204.600 684.600 206.700 ;
        RECT 704.400 205.800 708.600 206.700 ;
        RECT 720.000 206.400 726.300 207.300 ;
        RECT 727.200 208.200 728.250 213.900 ;
        RECT 729.600 211.200 731.400 213.000 ;
        RECT 733.950 211.800 736.050 213.900 ;
        RECT 745.950 211.950 748.050 214.050 ;
        RECT 729.150 209.100 731.250 211.200 ;
        RECT 682.800 198.600 684.600 204.600 ;
        RECT 685.800 203.700 693.600 205.050 ;
        RECT 685.800 198.600 687.600 203.700 ;
        RECT 688.800 198.000 690.600 202.800 ;
        RECT 691.800 198.600 693.600 203.700 ;
        RECT 704.400 198.600 706.200 205.800 ;
        RECT 720.000 204.600 721.200 206.400 ;
        RECT 727.200 206.100 730.050 208.200 ;
        RECT 750.150 207.300 751.050 218.700 ;
        RECT 753.000 214.050 754.200 221.400 ;
        RECT 767.400 214.050 768.600 227.400 ;
        RECT 779.400 221.400 781.200 234.000 ;
        RECT 784.500 222.600 786.300 233.400 ;
        RECT 799.800 227.400 801.600 233.400 ;
        RECT 802.800 227.400 804.600 234.000 ;
        RECT 814.800 227.400 816.600 234.000 ;
        RECT 817.800 227.400 819.600 233.400 ;
        RECT 820.800 227.400 822.600 234.000 ;
        RECT 833.400 227.400 835.200 234.000 ;
        RECT 836.400 227.400 838.200 233.400 ;
        RECT 782.700 221.400 786.300 222.600 ;
        RECT 770.100 214.050 771.900 215.850 ;
        RECT 779.100 214.050 780.900 215.850 ;
        RECT 782.700 214.050 783.600 221.400 ;
        RECT 785.100 214.050 786.900 215.850 ;
        RECT 800.400 214.050 801.600 227.400 ;
        RECT 803.100 214.050 804.900 215.850 ;
        RECT 751.950 211.950 754.200 214.050 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 769.950 211.950 772.050 214.050 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 818.400 213.900 819.600 227.400 ;
        RECT 836.850 214.050 838.050 227.400 ;
        RECT 841.500 221.400 843.300 234.000 ;
        RECT 842.100 214.050 843.900 215.850 ;
        RECT 727.200 204.600 728.400 206.100 ;
        RECT 731.400 205.500 733.500 206.700 ;
        RECT 750.150 206.400 752.100 207.300 ;
        RECT 746.400 205.500 752.100 206.400 ;
        RECT 731.400 204.600 736.200 205.500 ;
        RECT 709.500 198.000 711.300 204.600 ;
        RECT 719.400 198.600 721.200 204.600 ;
        RECT 726.900 198.600 728.700 204.600 ;
        RECT 734.400 198.600 736.200 204.600 ;
        RECT 746.400 201.600 747.600 205.500 ;
        RECT 753.000 204.600 754.200 211.950 ;
        RECT 746.400 198.600 748.200 201.600 ;
        RECT 749.400 198.000 751.200 201.600 ;
        RECT 752.400 198.600 754.200 204.600 ;
        RECT 767.400 201.600 768.600 211.950 ;
        RECT 782.700 201.600 783.600 211.950 ;
        RECT 800.400 201.600 801.600 211.950 ;
        RECT 814.950 211.800 817.050 213.900 ;
        RECT 817.950 211.800 820.050 213.900 ;
        RECT 820.950 211.800 823.050 213.900 ;
        RECT 832.950 211.950 835.050 214.050 ;
        RECT 835.950 211.950 838.050 214.050 ;
        RECT 838.950 211.950 841.050 214.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 815.100 210.000 816.900 211.800 ;
        RECT 818.400 206.700 819.600 211.800 ;
        RECT 821.100 210.000 822.900 211.800 ;
        RECT 833.100 210.150 834.900 211.950 ;
        RECT 835.950 207.750 837.150 211.950 ;
        RECT 839.100 210.150 840.900 211.950 ;
        RECT 815.400 205.800 819.600 206.700 ;
        RECT 833.400 206.700 837.150 207.750 ;
        RECT 766.800 198.600 768.600 201.600 ;
        RECT 769.800 198.000 771.600 201.600 ;
        RECT 779.400 198.000 781.200 201.600 ;
        RECT 782.400 198.600 784.200 201.600 ;
        RECT 785.400 198.000 787.200 201.600 ;
        RECT 799.800 198.600 801.600 201.600 ;
        RECT 802.800 198.000 804.600 201.600 ;
        RECT 815.400 198.600 817.200 205.800 ;
        RECT 833.400 204.600 834.600 206.700 ;
        RECT 820.500 198.000 822.300 204.600 ;
        RECT 832.800 198.600 834.600 204.600 ;
        RECT 835.800 203.700 843.600 205.050 ;
        RECT 835.800 198.600 837.600 203.700 ;
        RECT 838.800 198.000 840.600 202.800 ;
        RECT 841.800 198.600 843.600 203.700 ;
        RECT 8.400 191.400 10.200 195.000 ;
        RECT 11.400 191.400 13.200 194.400 ;
        RECT 11.400 181.050 12.600 191.400 ;
        RECT 17.550 188.400 19.350 194.400 ;
        RECT 20.850 191.400 22.650 195.000 ;
        RECT 25.650 191.400 27.450 194.400 ;
        RECT 29.850 191.400 31.650 195.000 ;
        RECT 33.450 191.400 35.250 194.400 ;
        RECT 36.750 191.400 38.550 195.000 ;
        RECT 41.250 192.300 43.050 194.400 ;
        RECT 41.250 191.400 45.000 192.300 ;
        RECT 46.050 191.400 47.850 195.000 ;
        RECT 25.650 190.500 26.700 191.400 ;
        RECT 22.950 189.300 26.700 190.500 ;
        RECT 34.200 190.500 35.250 191.400 ;
        RECT 43.950 190.500 45.000 191.400 ;
        RECT 34.200 189.450 39.150 190.500 ;
        RECT 22.950 188.400 25.050 189.300 ;
        RECT 37.350 188.700 39.150 189.450 ;
        RECT 17.550 181.050 18.750 188.400 ;
        RECT 40.650 187.800 42.450 189.600 ;
        RECT 43.950 188.400 46.050 190.500 ;
        RECT 49.050 188.400 50.850 194.400 ;
        RECT 59.700 188.400 61.500 195.000 ;
        RECT 30.150 186.000 31.950 186.600 ;
        RECT 41.100 186.000 42.150 187.800 ;
        RECT 30.150 184.800 42.150 186.000 ;
        RECT 7.950 178.950 10.050 181.050 ;
        RECT 10.950 178.950 13.050 181.050 ;
        RECT 17.550 179.250 23.850 181.050 ;
        RECT 17.550 178.950 22.050 179.250 ;
        RECT 8.100 177.150 9.900 178.950 ;
        RECT 11.400 165.600 12.600 178.950 ;
        RECT 17.550 171.600 18.750 178.950 ;
        RECT 19.950 173.400 21.750 175.200 ;
        RECT 20.850 172.200 25.050 173.400 ;
        RECT 30.150 172.200 31.050 184.800 ;
        RECT 41.100 183.600 48.000 184.800 ;
        RECT 41.100 183.000 42.900 183.600 ;
        RECT 47.100 182.850 48.000 183.600 ;
        RECT 44.100 181.800 45.900 182.400 ;
        RECT 37.950 180.600 45.900 181.800 ;
        RECT 47.100 181.050 48.900 182.850 ;
        RECT 37.950 178.950 40.050 180.600 ;
        RECT 46.950 178.950 49.050 181.050 ;
        RECT 39.750 173.700 41.550 174.000 ;
        RECT 49.950 173.700 50.850 188.400 ;
        RECT 64.800 187.200 66.600 194.400 ;
        RECT 77.400 191.400 79.200 195.000 ;
        RECT 80.400 191.400 82.200 194.400 ;
        RECT 62.400 186.300 66.600 187.200 ;
        RECT 59.100 181.200 60.900 183.000 ;
        RECT 62.400 181.200 63.600 186.300 ;
        RECT 65.100 181.200 66.900 183.000 ;
        RECT 58.950 179.100 61.050 181.200 ;
        RECT 61.950 179.100 64.050 181.200 ;
        RECT 64.950 179.100 67.050 181.200 ;
        RECT 80.400 181.050 81.600 191.400 ;
        RECT 92.400 189.300 94.200 194.400 ;
        RECT 95.400 190.200 97.200 195.000 ;
        RECT 98.400 189.300 100.200 194.400 ;
        RECT 92.400 187.950 100.200 189.300 ;
        RECT 101.400 188.400 103.200 194.400 ;
        RECT 113.400 189.300 115.200 194.400 ;
        RECT 116.400 190.200 118.200 195.000 ;
        RECT 119.400 189.300 121.200 194.400 ;
        RECT 101.400 186.300 102.600 188.400 ;
        RECT 113.400 187.950 121.200 189.300 ;
        RECT 122.400 188.400 124.200 194.400 ;
        RECT 134.400 191.400 136.200 195.000 ;
        RECT 137.400 191.400 139.200 194.400 ;
        RECT 140.400 191.400 142.200 195.000 ;
        RECT 122.400 186.300 123.600 188.400 ;
        RECT 98.850 185.250 102.600 186.300 ;
        RECT 119.850 185.250 123.600 186.300 ;
        RECT 95.100 181.050 96.900 182.850 ;
        RECT 98.850 181.050 100.050 185.250 ;
        RECT 108.000 183.450 112.050 184.050 ;
        RECT 101.100 181.050 102.900 182.850 ;
        RECT 107.550 181.950 112.050 183.450 ;
        RECT 39.750 173.100 50.850 173.700 ;
        RECT 8.400 159.000 10.200 165.600 ;
        RECT 11.400 159.600 13.200 165.600 ;
        RECT 17.550 159.600 19.350 171.600 ;
        RECT 22.950 171.300 25.050 172.200 ;
        RECT 25.950 171.300 31.050 172.200 ;
        RECT 33.150 172.500 50.850 173.100 ;
        RECT 33.150 172.200 41.550 172.500 ;
        RECT 25.950 170.400 26.850 171.300 ;
        RECT 24.150 168.600 26.850 170.400 ;
        RECT 27.750 170.100 29.550 170.400 ;
        RECT 33.150 170.100 34.050 172.200 ;
        RECT 49.950 171.600 50.850 172.500 ;
        RECT 27.750 169.200 34.050 170.100 ;
        RECT 34.950 170.700 36.750 171.300 ;
        RECT 34.950 169.500 42.450 170.700 ;
        RECT 27.750 168.600 29.550 169.200 ;
        RECT 41.250 168.600 42.450 169.500 ;
        RECT 22.950 165.600 26.850 167.700 ;
        RECT 31.950 167.550 33.750 168.300 ;
        RECT 36.750 167.550 38.550 168.300 ;
        RECT 31.950 166.500 38.550 167.550 ;
        RECT 41.250 166.500 46.050 168.600 ;
        RECT 20.550 159.000 22.350 162.600 ;
        RECT 25.050 159.600 26.850 165.600 ;
        RECT 29.250 159.000 31.050 165.600 ;
        RECT 32.850 159.600 34.650 166.500 ;
        RECT 41.250 165.600 42.450 166.500 ;
        RECT 35.850 159.000 37.650 165.600 ;
        RECT 40.650 159.600 42.450 165.600 ;
        RECT 46.050 159.000 47.850 165.600 ;
        RECT 49.050 159.600 50.850 171.600 ;
        RECT 62.400 165.600 63.600 179.100 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 77.100 177.150 78.900 178.950 ;
        RECT 80.400 165.600 81.600 178.950 ;
        RECT 92.100 177.150 93.900 178.950 ;
        RECT 59.400 159.000 61.200 165.600 ;
        RECT 62.400 159.600 64.200 165.600 ;
        RECT 65.400 159.000 67.200 165.600 ;
        RECT 77.400 159.000 79.200 165.600 ;
        RECT 80.400 159.600 82.200 165.600 ;
        RECT 92.700 159.000 94.500 171.600 ;
        RECT 97.950 165.600 99.150 178.950 ;
        RECT 107.550 178.050 108.450 181.950 ;
        RECT 116.100 181.050 117.900 182.850 ;
        RECT 119.850 181.050 121.050 185.250 ;
        RECT 122.100 181.050 123.900 182.850 ;
        RECT 137.700 181.050 138.600 191.400 ;
        RECT 154.800 188.400 156.600 195.000 ;
        RECT 157.800 187.500 159.600 194.400 ;
        RECT 160.800 188.400 162.600 195.000 ;
        RECT 163.800 187.500 165.600 194.400 ;
        RECT 166.800 188.400 168.600 195.000 ;
        RECT 169.800 187.500 171.600 194.400 ;
        RECT 172.800 188.400 174.600 195.000 ;
        RECT 175.800 187.500 177.600 194.400 ;
        RECT 178.800 188.400 180.600 195.000 ;
        RECT 190.800 188.400 192.600 194.400 ;
        RECT 193.800 191.400 195.600 195.000 ;
        RECT 196.800 191.400 198.600 194.400 ;
        RECT 156.900 186.300 159.600 187.500 ;
        RECT 161.700 186.300 165.600 187.500 ;
        RECT 167.700 186.300 171.600 187.500 ;
        RECT 173.700 186.300 177.600 187.500 ;
        RECT 156.900 181.200 157.800 186.300 ;
        RECT 161.700 185.400 162.900 186.300 ;
        RECT 167.700 185.400 168.900 186.300 ;
        RECT 173.700 185.400 174.900 186.300 ;
        RECT 158.700 184.200 162.900 185.400 ;
        RECT 158.700 183.600 160.500 184.200 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 121.950 178.950 124.050 181.050 ;
        RECT 133.950 178.950 136.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 154.950 179.100 157.800 181.200 ;
        RECT 103.950 176.550 108.450 178.050 ;
        RECT 113.100 177.150 114.900 178.950 ;
        RECT 103.950 175.950 108.000 176.550 ;
        RECT 97.800 159.600 99.600 165.600 ;
        RECT 100.800 159.000 102.600 165.600 ;
        RECT 113.700 159.000 115.500 171.600 ;
        RECT 118.950 165.600 120.150 178.950 ;
        RECT 134.100 177.150 135.900 178.950 ;
        RECT 137.700 171.600 138.600 178.950 ;
        RECT 140.100 177.150 141.900 178.950 ;
        RECT 156.900 173.700 157.800 179.100 ;
        RECT 161.700 173.700 162.900 184.200 ;
        RECT 164.700 184.200 168.900 185.400 ;
        RECT 164.700 183.600 166.500 184.200 ;
        RECT 167.700 173.700 168.900 184.200 ;
        RECT 170.700 184.200 174.900 185.400 ;
        RECT 170.700 183.600 172.500 184.200 ;
        RECT 173.700 173.700 174.900 184.200 ;
        RECT 176.100 181.200 177.900 183.000 ;
        RECT 175.950 179.100 178.050 181.200 ;
        RECT 190.800 181.050 192.000 188.400 ;
        RECT 197.400 187.500 198.600 191.400 ;
        RECT 206.700 188.400 208.500 195.000 ;
        RECT 192.900 186.600 198.600 187.500 ;
        RECT 211.800 187.200 213.600 194.400 ;
        RECT 226.800 188.400 228.600 194.400 ;
        RECT 192.900 185.700 194.850 186.600 ;
        RECT 190.800 178.950 193.050 181.050 ;
        RECT 178.950 177.450 181.050 178.050 ;
        RECT 184.950 177.450 187.050 178.050 ;
        RECT 178.950 176.550 187.050 177.450 ;
        RECT 178.950 175.950 181.050 176.550 ;
        RECT 184.950 175.950 187.050 176.550 ;
        RECT 156.900 172.500 159.600 173.700 ;
        RECT 161.700 172.500 165.600 173.700 ;
        RECT 167.700 172.500 171.600 173.700 ;
        RECT 173.700 172.500 177.600 173.700 ;
        RECT 118.800 159.600 120.600 165.600 ;
        RECT 121.800 159.000 123.600 165.600 ;
        RECT 134.400 159.000 136.200 171.600 ;
        RECT 137.700 170.400 141.300 171.600 ;
        RECT 139.500 159.600 141.300 170.400 ;
        RECT 154.800 159.000 156.600 171.600 ;
        RECT 157.800 159.600 159.600 172.500 ;
        RECT 160.800 159.000 162.600 171.600 ;
        RECT 163.800 159.600 165.600 172.500 ;
        RECT 166.800 159.000 168.600 171.600 ;
        RECT 169.800 159.600 171.600 172.500 ;
        RECT 172.800 159.000 174.600 171.600 ;
        RECT 175.800 159.600 177.600 172.500 ;
        RECT 190.800 171.600 192.000 178.950 ;
        RECT 193.950 174.300 194.850 185.700 ;
        RECT 209.400 186.300 213.600 187.200 ;
        RECT 227.400 186.300 228.600 188.400 ;
        RECT 229.800 189.300 231.600 194.400 ;
        RECT 232.800 190.200 234.600 195.000 ;
        RECT 235.800 189.300 237.600 194.400 ;
        RECT 229.800 187.950 237.600 189.300 ;
        RECT 240.150 188.400 241.950 194.400 ;
        RECT 243.150 191.400 244.950 195.000 ;
        RECT 247.950 192.300 249.750 194.400 ;
        RECT 246.000 191.400 249.750 192.300 ;
        RECT 252.450 191.400 254.250 195.000 ;
        RECT 255.750 191.400 257.550 194.400 ;
        RECT 259.350 191.400 261.150 195.000 ;
        RECT 263.550 191.400 265.350 194.400 ;
        RECT 268.350 191.400 270.150 195.000 ;
        RECT 246.000 190.500 247.050 191.400 ;
        RECT 255.750 190.500 256.800 191.400 ;
        RECT 244.950 188.400 247.050 190.500 ;
        RECT 206.100 181.200 207.900 183.000 ;
        RECT 209.400 181.200 210.600 186.300 ;
        RECT 227.400 185.250 231.150 186.300 ;
        RECT 212.100 181.200 213.900 183.000 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 205.950 179.100 208.050 181.200 ;
        RECT 208.950 179.100 211.050 181.200 ;
        RECT 211.950 179.100 214.050 181.200 ;
        RECT 227.100 181.050 228.900 182.850 ;
        RECT 229.950 181.050 231.150 185.250 ;
        RECT 233.100 181.050 234.900 182.850 ;
        RECT 197.100 177.150 198.900 178.950 ;
        RECT 192.900 173.400 194.850 174.300 ;
        RECT 192.900 172.500 198.600 173.400 ;
        RECT 178.800 159.000 180.600 171.600 ;
        RECT 190.800 159.600 192.600 171.600 ;
        RECT 197.400 165.600 198.600 172.500 ;
        RECT 209.400 165.600 210.600 179.100 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 229.950 178.950 232.050 181.050 ;
        RECT 232.950 178.950 235.050 181.050 ;
        RECT 235.950 178.950 238.050 181.050 ;
        RECT 230.850 165.600 232.050 178.950 ;
        RECT 236.100 177.150 237.900 178.950 ;
        RECT 240.150 173.700 241.050 188.400 ;
        RECT 248.550 187.800 250.350 189.600 ;
        RECT 251.850 189.450 256.800 190.500 ;
        RECT 264.300 190.500 265.350 191.400 ;
        RECT 251.850 188.700 253.650 189.450 ;
        RECT 264.300 189.300 268.050 190.500 ;
        RECT 265.950 188.400 268.050 189.300 ;
        RECT 271.650 188.400 273.450 194.400 ;
        RECT 281.700 188.400 283.500 195.000 ;
        RECT 248.850 186.000 249.900 187.800 ;
        RECT 259.050 186.000 260.850 186.600 ;
        RECT 248.850 184.800 260.850 186.000 ;
        RECT 243.000 183.600 249.900 184.800 ;
        RECT 243.000 182.850 243.900 183.600 ;
        RECT 248.100 183.000 249.900 183.600 ;
        RECT 242.100 181.050 243.900 182.850 ;
        RECT 245.100 181.800 246.900 182.400 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 245.100 180.600 253.050 181.800 ;
        RECT 250.950 178.950 253.050 180.600 ;
        RECT 249.450 173.700 251.250 174.000 ;
        RECT 240.150 173.100 251.250 173.700 ;
        RECT 240.150 172.500 257.850 173.100 ;
        RECT 240.150 171.600 241.050 172.500 ;
        RECT 249.450 172.200 257.850 172.500 ;
        RECT 193.800 159.000 195.600 165.600 ;
        RECT 196.800 159.600 198.600 165.600 ;
        RECT 206.400 159.000 208.200 165.600 ;
        RECT 209.400 159.600 211.200 165.600 ;
        RECT 212.400 159.000 214.200 165.600 ;
        RECT 227.400 159.000 229.200 165.600 ;
        RECT 230.400 159.600 232.200 165.600 ;
        RECT 235.500 159.000 237.300 171.600 ;
        RECT 240.150 159.600 241.950 171.600 ;
        RECT 254.250 170.700 256.050 171.300 ;
        RECT 248.550 169.500 256.050 170.700 ;
        RECT 256.950 170.100 257.850 172.200 ;
        RECT 259.950 172.200 260.850 184.800 ;
        RECT 272.250 181.050 273.450 188.400 ;
        RECT 286.800 187.200 288.600 194.400 ;
        RECT 301.800 188.400 303.600 194.400 ;
        RECT 284.400 186.300 288.600 187.200 ;
        RECT 302.400 186.300 303.600 188.400 ;
        RECT 304.800 189.300 306.600 194.400 ;
        RECT 307.800 190.200 309.600 195.000 ;
        RECT 310.800 189.300 312.600 194.400 ;
        RECT 304.800 187.950 312.600 189.300 ;
        RECT 322.800 188.400 324.600 194.400 ;
        RECT 323.400 186.300 324.600 188.400 ;
        RECT 325.800 189.300 327.600 194.400 ;
        RECT 328.800 190.200 330.600 195.000 ;
        RECT 331.800 189.300 333.600 194.400 ;
        RECT 325.800 187.950 333.600 189.300 ;
        RECT 336.150 188.400 337.950 194.400 ;
        RECT 339.150 191.400 340.950 195.000 ;
        RECT 343.950 192.300 345.750 194.400 ;
        RECT 342.000 191.400 345.750 192.300 ;
        RECT 348.450 191.400 350.250 195.000 ;
        RECT 351.750 191.400 353.550 194.400 ;
        RECT 355.350 191.400 357.150 195.000 ;
        RECT 359.550 191.400 361.350 194.400 ;
        RECT 364.350 191.400 366.150 195.000 ;
        RECT 342.000 190.500 343.050 191.400 ;
        RECT 351.750 190.500 352.800 191.400 ;
        RECT 340.950 188.400 343.050 190.500 ;
        RECT 281.100 181.200 282.900 183.000 ;
        RECT 284.400 181.200 285.600 186.300 ;
        RECT 302.400 185.250 306.150 186.300 ;
        RECT 323.400 185.250 327.150 186.300 ;
        RECT 289.950 183.450 294.000 184.050 ;
        RECT 287.100 181.200 288.900 183.000 ;
        RECT 289.950 181.950 294.450 183.450 ;
        RECT 267.150 179.250 273.450 181.050 ;
        RECT 268.950 178.950 273.450 179.250 ;
        RECT 280.950 179.100 283.050 181.200 ;
        RECT 283.950 179.100 286.050 181.200 ;
        RECT 286.950 179.100 289.050 181.200 ;
        RECT 269.250 173.400 271.050 175.200 ;
        RECT 265.950 172.200 270.150 173.400 ;
        RECT 259.950 171.300 265.050 172.200 ;
        RECT 265.950 171.300 268.050 172.200 ;
        RECT 272.250 171.600 273.450 178.950 ;
        RECT 264.150 170.400 265.050 171.300 ;
        RECT 261.450 170.100 263.250 170.400 ;
        RECT 248.550 168.600 249.750 169.500 ;
        RECT 256.950 169.200 263.250 170.100 ;
        RECT 261.450 168.600 263.250 169.200 ;
        RECT 264.150 168.600 266.850 170.400 ;
        RECT 244.950 166.500 249.750 168.600 ;
        RECT 252.450 167.550 254.250 168.300 ;
        RECT 257.250 167.550 259.050 168.300 ;
        RECT 252.450 166.500 259.050 167.550 ;
        RECT 248.550 165.600 249.750 166.500 ;
        RECT 243.150 159.000 244.950 165.600 ;
        RECT 248.550 159.600 250.350 165.600 ;
        RECT 253.350 159.000 255.150 165.600 ;
        RECT 256.350 159.600 258.150 166.500 ;
        RECT 264.150 165.600 268.050 167.700 ;
        RECT 259.950 159.000 261.750 165.600 ;
        RECT 264.150 159.600 265.950 165.600 ;
        RECT 268.650 159.000 270.450 162.600 ;
        RECT 271.650 159.600 273.450 171.600 ;
        RECT 284.400 165.600 285.600 179.100 ;
        RECT 293.550 178.050 294.450 181.950 ;
        RECT 302.100 181.050 303.900 182.850 ;
        RECT 304.950 181.050 306.150 185.250 ;
        RECT 308.100 181.050 309.900 182.850 ;
        RECT 323.100 181.050 324.900 182.850 ;
        RECT 325.950 181.050 327.150 185.250 ;
        RECT 329.100 181.050 330.900 182.850 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 304.950 178.950 307.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 325.950 178.950 328.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 289.950 176.550 294.450 178.050 ;
        RECT 289.950 175.950 294.000 176.550 ;
        RECT 305.850 165.600 307.050 178.950 ;
        RECT 311.100 177.150 312.900 178.950 ;
        RECT 310.950 174.450 313.050 175.050 ;
        RECT 319.950 174.450 322.050 175.050 ;
        RECT 310.950 173.550 322.050 174.450 ;
        RECT 310.950 172.950 313.050 173.550 ;
        RECT 319.950 172.950 322.050 173.550 ;
        RECT 281.400 159.000 283.200 165.600 ;
        RECT 284.400 159.600 286.200 165.600 ;
        RECT 287.400 159.000 289.200 165.600 ;
        RECT 302.400 159.000 304.200 165.600 ;
        RECT 305.400 159.600 307.200 165.600 ;
        RECT 310.500 159.000 312.300 171.600 ;
        RECT 313.950 171.450 316.050 172.050 ;
        RECT 319.950 171.450 322.050 171.900 ;
        RECT 313.950 170.550 322.050 171.450 ;
        RECT 313.950 169.950 316.050 170.550 ;
        RECT 319.950 169.800 322.050 170.550 ;
        RECT 326.850 165.600 328.050 178.950 ;
        RECT 332.100 177.150 333.900 178.950 ;
        RECT 336.150 173.700 337.050 188.400 ;
        RECT 344.550 187.800 346.350 189.600 ;
        RECT 347.850 189.450 352.800 190.500 ;
        RECT 360.300 190.500 361.350 191.400 ;
        RECT 347.850 188.700 349.650 189.450 ;
        RECT 360.300 189.300 364.050 190.500 ;
        RECT 361.950 188.400 364.050 189.300 ;
        RECT 367.650 188.400 369.450 194.400 ;
        RECT 344.850 186.000 345.900 187.800 ;
        RECT 355.050 186.000 356.850 186.600 ;
        RECT 344.850 184.800 356.850 186.000 ;
        RECT 339.000 183.600 345.900 184.800 ;
        RECT 339.000 182.850 339.900 183.600 ;
        RECT 344.100 183.000 345.900 183.600 ;
        RECT 338.100 181.050 339.900 182.850 ;
        RECT 341.100 181.800 342.900 182.400 ;
        RECT 337.950 178.950 340.050 181.050 ;
        RECT 341.100 180.600 349.050 181.800 ;
        RECT 346.950 178.950 349.050 180.600 ;
        RECT 345.450 173.700 347.250 174.000 ;
        RECT 336.150 173.100 347.250 173.700 ;
        RECT 336.150 172.500 353.850 173.100 ;
        RECT 336.150 171.600 337.050 172.500 ;
        RECT 345.450 172.200 353.850 172.500 ;
        RECT 323.400 159.000 325.200 165.600 ;
        RECT 326.400 159.600 328.200 165.600 ;
        RECT 331.500 159.000 333.300 171.600 ;
        RECT 336.150 159.600 337.950 171.600 ;
        RECT 350.250 170.700 352.050 171.300 ;
        RECT 344.550 169.500 352.050 170.700 ;
        RECT 352.950 170.100 353.850 172.200 ;
        RECT 355.950 172.200 356.850 184.800 ;
        RECT 368.250 181.050 369.450 188.400 ;
        RECT 377.400 189.300 379.200 194.400 ;
        RECT 380.400 190.200 382.200 195.000 ;
        RECT 383.400 189.300 385.200 194.400 ;
        RECT 377.400 187.950 385.200 189.300 ;
        RECT 386.400 188.400 388.200 194.400 ;
        RECT 400.800 188.400 402.600 194.400 ;
        RECT 386.400 186.300 387.600 188.400 ;
        RECT 383.850 185.250 387.600 186.300 ;
        RECT 401.400 186.300 402.600 188.400 ;
        RECT 403.800 189.300 405.600 194.400 ;
        RECT 406.800 190.200 408.600 195.000 ;
        RECT 409.800 189.300 411.600 194.400 ;
        RECT 419.400 191.400 421.200 195.000 ;
        RECT 422.400 191.400 424.200 194.400 ;
        RECT 425.400 191.400 427.200 195.000 ;
        RECT 403.800 187.950 411.600 189.300 ;
        RECT 401.400 185.250 405.150 186.300 ;
        RECT 380.100 181.050 381.900 182.850 ;
        RECT 383.850 181.050 385.050 185.250 ;
        RECT 386.100 181.050 387.900 182.850 ;
        RECT 401.100 181.050 402.900 182.850 ;
        RECT 403.950 181.050 405.150 185.250 ;
        RECT 407.100 181.050 408.900 182.850 ;
        RECT 422.700 181.050 423.600 191.400 ;
        RECT 437.700 188.400 439.500 195.000 ;
        RECT 442.200 188.400 444.000 194.400 ;
        RECT 446.700 188.400 448.500 195.000 ;
        RECT 461.400 188.400 463.200 195.000 ;
        RECT 437.100 181.200 438.900 183.000 ;
        RECT 442.950 181.200 444.000 188.400 ;
        RECT 464.400 187.500 466.200 194.400 ;
        RECT 467.400 188.400 469.200 195.000 ;
        RECT 470.400 187.500 472.200 194.400 ;
        RECT 473.400 188.400 475.200 195.000 ;
        RECT 476.400 187.500 478.200 194.400 ;
        RECT 479.400 188.400 481.200 195.000 ;
        RECT 482.400 187.500 484.200 194.400 ;
        RECT 485.400 188.400 487.200 195.000 ;
        RECT 498.000 188.400 499.800 195.000 ;
        RECT 502.500 189.600 504.300 194.400 ;
        RECT 505.500 191.400 507.300 195.000 ;
        RECT 502.500 188.400 507.600 189.600 ;
        RECT 464.400 186.300 468.300 187.500 ;
        RECT 470.400 186.300 474.300 187.500 ;
        RECT 476.400 186.300 480.300 187.500 ;
        RECT 482.400 186.300 485.100 187.500 ;
        RECT 467.100 185.400 468.300 186.300 ;
        RECT 473.100 185.400 474.300 186.300 ;
        RECT 479.100 185.400 480.300 186.300 ;
        RECT 467.100 184.200 471.300 185.400 ;
        RECT 449.100 181.200 450.900 183.000 ;
        RECT 464.100 181.200 465.900 183.000 ;
        RECT 363.150 179.250 369.450 181.050 ;
        RECT 364.950 178.950 369.450 179.250 ;
        RECT 376.950 178.950 379.050 181.050 ;
        RECT 379.950 178.950 382.050 181.050 ;
        RECT 382.950 178.950 385.050 181.050 ;
        RECT 385.950 178.950 388.050 181.050 ;
        RECT 400.950 178.950 403.050 181.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 418.950 178.950 421.050 181.050 ;
        RECT 421.950 178.950 424.050 181.050 ;
        RECT 424.950 178.950 427.050 181.050 ;
        RECT 436.950 179.100 439.050 181.200 ;
        RECT 439.950 179.100 442.050 181.200 ;
        RECT 442.950 179.100 445.050 181.200 ;
        RECT 445.950 179.100 448.050 181.200 ;
        RECT 448.950 179.100 451.050 181.200 ;
        RECT 463.950 179.100 466.050 181.200 ;
        RECT 365.250 173.400 367.050 175.200 ;
        RECT 361.950 172.200 366.150 173.400 ;
        RECT 355.950 171.300 361.050 172.200 ;
        RECT 361.950 171.300 364.050 172.200 ;
        RECT 368.250 171.600 369.450 178.950 ;
        RECT 377.100 177.150 378.900 178.950 ;
        RECT 360.150 170.400 361.050 171.300 ;
        RECT 357.450 170.100 359.250 170.400 ;
        RECT 344.550 168.600 345.750 169.500 ;
        RECT 352.950 169.200 359.250 170.100 ;
        RECT 357.450 168.600 359.250 169.200 ;
        RECT 360.150 168.600 362.850 170.400 ;
        RECT 340.950 166.500 345.750 168.600 ;
        RECT 348.450 167.550 350.250 168.300 ;
        RECT 353.250 167.550 355.050 168.300 ;
        RECT 348.450 166.500 355.050 167.550 ;
        RECT 344.550 165.600 345.750 166.500 ;
        RECT 339.150 159.000 340.950 165.600 ;
        RECT 344.550 159.600 346.350 165.600 ;
        RECT 349.350 159.000 351.150 165.600 ;
        RECT 352.350 159.600 354.150 166.500 ;
        RECT 360.150 165.600 364.050 167.700 ;
        RECT 355.950 159.000 357.750 165.600 ;
        RECT 360.150 159.600 361.950 165.600 ;
        RECT 364.650 159.000 366.450 162.600 ;
        RECT 367.650 159.600 369.450 171.600 ;
        RECT 377.700 159.000 379.500 171.600 ;
        RECT 382.950 165.600 384.150 178.950 ;
        RECT 404.850 165.600 406.050 178.950 ;
        RECT 410.100 177.150 411.900 178.950 ;
        RECT 419.100 177.150 420.900 178.950 ;
        RECT 422.700 171.600 423.600 178.950 ;
        RECT 425.100 177.150 426.900 178.950 ;
        RECT 440.100 177.300 441.900 179.100 ;
        RECT 443.100 173.400 444.000 179.100 ;
        RECT 446.100 177.300 447.900 179.100 ;
        RECT 467.100 173.700 468.300 184.200 ;
        RECT 469.500 183.600 471.300 184.200 ;
        RECT 473.100 184.200 477.300 185.400 ;
        RECT 473.100 173.700 474.300 184.200 ;
        RECT 475.500 183.600 477.300 184.200 ;
        RECT 479.100 184.200 483.300 185.400 ;
        RECT 479.100 173.700 480.300 184.200 ;
        RECT 481.500 183.600 483.300 184.200 ;
        RECT 484.200 181.200 485.100 186.300 ;
        RECT 497.100 181.200 498.900 183.000 ;
        RECT 503.100 181.200 504.900 183.000 ;
        RECT 506.700 181.200 507.600 188.400 ;
        RECT 513.150 188.400 514.950 194.400 ;
        RECT 516.150 191.400 517.950 195.000 ;
        RECT 520.950 192.300 522.750 194.400 ;
        RECT 519.000 191.400 522.750 192.300 ;
        RECT 525.450 191.400 527.250 195.000 ;
        RECT 528.750 191.400 530.550 194.400 ;
        RECT 532.350 191.400 534.150 195.000 ;
        RECT 536.550 191.400 538.350 194.400 ;
        RECT 541.350 191.400 543.150 195.000 ;
        RECT 519.000 190.500 520.050 191.400 ;
        RECT 528.750 190.500 529.800 191.400 ;
        RECT 517.950 188.400 520.050 190.500 ;
        RECT 484.200 179.100 487.050 181.200 ;
        RECT 496.950 179.100 499.050 181.200 ;
        RECT 499.950 179.100 502.050 181.200 ;
        RECT 502.950 179.100 505.050 181.200 ;
        RECT 505.950 179.100 508.050 181.200 ;
        RECT 484.200 173.700 485.100 179.100 ;
        RECT 500.100 177.300 501.900 179.100 ;
        RECT 443.100 172.500 448.200 173.400 ;
        RECT 382.800 159.600 384.600 165.600 ;
        RECT 385.800 159.000 387.600 165.600 ;
        RECT 401.400 159.000 403.200 165.600 ;
        RECT 404.400 159.600 406.200 165.600 ;
        RECT 409.500 159.000 411.300 171.600 ;
        RECT 419.400 159.000 421.200 171.600 ;
        RECT 422.700 170.400 426.300 171.600 ;
        RECT 424.500 159.600 426.300 170.400 ;
        RECT 437.400 170.400 445.200 171.300 ;
        RECT 437.400 159.600 439.200 170.400 ;
        RECT 440.400 159.000 442.200 169.500 ;
        RECT 443.400 160.500 445.200 170.400 ;
        RECT 446.400 161.400 448.200 172.500 ;
        RECT 464.400 172.500 468.300 173.700 ;
        RECT 470.400 172.500 474.300 173.700 ;
        RECT 476.400 172.500 480.300 173.700 ;
        RECT 482.400 172.500 485.100 173.700 ;
        RECT 449.400 160.500 451.200 171.600 ;
        RECT 443.400 159.600 451.200 160.500 ;
        RECT 461.400 159.000 463.200 171.600 ;
        RECT 464.400 159.600 466.200 172.500 ;
        RECT 467.400 159.000 469.200 171.600 ;
        RECT 470.400 159.600 472.200 172.500 ;
        RECT 473.400 159.000 475.200 171.600 ;
        RECT 476.400 159.600 478.200 172.500 ;
        RECT 479.400 159.000 481.200 171.600 ;
        RECT 482.400 159.600 484.200 172.500 ;
        RECT 506.700 171.600 507.600 179.100 ;
        RECT 513.150 173.700 514.050 188.400 ;
        RECT 521.550 187.800 523.350 189.600 ;
        RECT 524.850 189.450 529.800 190.500 ;
        RECT 537.300 190.500 538.350 191.400 ;
        RECT 524.850 188.700 526.650 189.450 ;
        RECT 537.300 189.300 541.050 190.500 ;
        RECT 538.950 188.400 541.050 189.300 ;
        RECT 544.650 188.400 546.450 194.400 ;
        RECT 554.400 191.400 556.200 195.000 ;
        RECT 557.400 191.400 559.200 194.400 ;
        RECT 560.400 191.400 562.200 195.000 ;
        RECT 521.850 186.000 522.900 187.800 ;
        RECT 532.050 186.000 533.850 186.600 ;
        RECT 521.850 184.800 533.850 186.000 ;
        RECT 516.000 183.600 522.900 184.800 ;
        RECT 516.000 182.850 516.900 183.600 ;
        RECT 521.100 183.000 522.900 183.600 ;
        RECT 515.100 181.050 516.900 182.850 ;
        RECT 518.100 181.800 519.900 182.400 ;
        RECT 514.950 178.950 517.050 181.050 ;
        RECT 518.100 180.600 526.050 181.800 ;
        RECT 523.950 178.950 526.050 180.600 ;
        RECT 522.450 173.700 524.250 174.000 ;
        RECT 513.150 173.100 524.250 173.700 ;
        RECT 513.150 172.500 530.850 173.100 ;
        RECT 513.150 171.600 514.050 172.500 ;
        RECT 522.450 172.200 530.850 172.500 ;
        RECT 485.400 159.000 487.200 171.600 ;
        RECT 497.400 170.700 505.200 171.600 ;
        RECT 497.400 159.600 499.200 170.700 ;
        RECT 500.400 159.000 502.200 169.800 ;
        RECT 503.400 159.600 505.200 170.700 ;
        RECT 506.400 159.600 508.200 171.600 ;
        RECT 513.150 159.600 514.950 171.600 ;
        RECT 527.250 170.700 529.050 171.300 ;
        RECT 521.550 169.500 529.050 170.700 ;
        RECT 529.950 170.100 530.850 172.200 ;
        RECT 532.950 172.200 533.850 184.800 ;
        RECT 545.250 181.050 546.450 188.400 ;
        RECT 557.700 181.050 558.600 191.400 ;
        RECT 572.400 188.400 574.200 195.000 ;
        RECT 575.400 187.500 577.200 194.400 ;
        RECT 578.400 188.400 580.200 195.000 ;
        RECT 581.400 187.500 583.200 194.400 ;
        RECT 584.400 188.400 586.200 195.000 ;
        RECT 587.400 187.500 589.200 194.400 ;
        RECT 590.400 188.400 592.200 195.000 ;
        RECT 593.400 187.500 595.200 194.400 ;
        RECT 596.400 188.400 598.200 195.000 ;
        RECT 575.400 186.300 579.300 187.500 ;
        RECT 581.400 186.300 585.300 187.500 ;
        RECT 587.400 186.300 591.300 187.500 ;
        RECT 593.400 186.300 596.100 187.500 ;
        RECT 611.400 187.200 613.200 194.400 ;
        RECT 616.500 188.400 618.300 195.000 ;
        RECT 627.000 188.400 628.800 195.000 ;
        RECT 631.500 189.600 633.300 194.400 ;
        RECT 634.500 191.400 636.300 195.000 ;
        RECT 649.800 191.400 651.600 195.000 ;
        RECT 652.800 191.400 654.600 194.400 ;
        RECT 655.800 191.400 657.600 195.000 ;
        RECT 631.500 188.400 636.600 189.600 ;
        RECT 611.400 186.300 615.600 187.200 ;
        RECT 578.100 185.400 579.300 186.300 ;
        RECT 584.100 185.400 585.300 186.300 ;
        RECT 590.100 185.400 591.300 186.300 ;
        RECT 578.100 184.200 582.300 185.400 ;
        RECT 575.100 181.200 576.900 183.000 ;
        RECT 540.150 179.250 546.450 181.050 ;
        RECT 541.950 178.950 546.450 179.250 ;
        RECT 553.950 178.950 556.050 181.050 ;
        RECT 556.950 178.950 559.050 181.050 ;
        RECT 559.950 178.950 562.050 181.050 ;
        RECT 574.950 179.100 577.050 181.200 ;
        RECT 542.250 173.400 544.050 175.200 ;
        RECT 538.950 172.200 543.150 173.400 ;
        RECT 532.950 171.300 538.050 172.200 ;
        RECT 538.950 171.300 541.050 172.200 ;
        RECT 545.250 171.600 546.450 178.950 ;
        RECT 554.100 177.150 555.900 178.950 ;
        RECT 557.700 171.600 558.600 178.950 ;
        RECT 560.100 177.150 561.900 178.950 ;
        RECT 578.100 173.700 579.300 184.200 ;
        RECT 580.500 183.600 582.300 184.200 ;
        RECT 584.100 184.200 588.300 185.400 ;
        RECT 584.100 173.700 585.300 184.200 ;
        RECT 586.500 183.600 588.300 184.200 ;
        RECT 590.100 184.200 594.300 185.400 ;
        RECT 590.100 173.700 591.300 184.200 ;
        RECT 592.500 183.600 594.300 184.200 ;
        RECT 595.200 181.200 596.100 186.300 ;
        RECT 611.100 181.200 612.900 183.000 ;
        RECT 614.400 181.200 615.600 186.300 ;
        RECT 617.100 181.200 618.900 183.000 ;
        RECT 626.100 181.200 627.900 183.000 ;
        RECT 632.100 181.200 633.900 183.000 ;
        RECT 635.700 181.200 636.600 188.400 ;
        RECT 595.200 179.100 598.050 181.200 ;
        RECT 610.950 179.100 613.050 181.200 ;
        RECT 613.950 179.100 616.050 181.200 ;
        RECT 616.950 179.100 619.050 181.200 ;
        RECT 625.950 179.100 628.050 181.200 ;
        RECT 628.950 179.100 631.050 181.200 ;
        RECT 631.950 179.100 634.050 181.200 ;
        RECT 634.950 179.100 637.050 181.200 ;
        RECT 653.400 181.050 654.300 191.400 ;
        RECT 659.550 188.400 661.350 194.400 ;
        RECT 662.850 191.400 664.650 195.000 ;
        RECT 667.650 191.400 669.450 194.400 ;
        RECT 671.850 191.400 673.650 195.000 ;
        RECT 675.450 191.400 677.250 194.400 ;
        RECT 678.750 191.400 680.550 195.000 ;
        RECT 683.250 192.300 685.050 194.400 ;
        RECT 683.250 191.400 687.000 192.300 ;
        RECT 688.050 191.400 689.850 195.000 ;
        RECT 667.650 190.500 668.700 191.400 ;
        RECT 664.950 189.300 668.700 190.500 ;
        RECT 676.200 190.500 677.250 191.400 ;
        RECT 685.950 190.500 687.000 191.400 ;
        RECT 676.200 189.450 681.150 190.500 ;
        RECT 664.950 188.400 667.050 189.300 ;
        RECT 679.350 188.700 681.150 189.450 ;
        RECT 659.550 181.050 660.750 188.400 ;
        RECT 682.650 187.800 684.450 189.600 ;
        RECT 685.950 188.400 688.050 190.500 ;
        RECT 691.050 188.400 692.850 194.400 ;
        RECT 672.150 186.000 673.950 186.600 ;
        RECT 683.100 186.000 684.150 187.800 ;
        RECT 672.150 184.800 684.150 186.000 ;
        RECT 595.200 173.700 596.100 179.100 ;
        RECT 575.400 172.500 579.300 173.700 ;
        RECT 581.400 172.500 585.300 173.700 ;
        RECT 587.400 172.500 591.300 173.700 ;
        RECT 593.400 172.500 596.100 173.700 ;
        RECT 537.150 170.400 538.050 171.300 ;
        RECT 534.450 170.100 536.250 170.400 ;
        RECT 521.550 168.600 522.750 169.500 ;
        RECT 529.950 169.200 536.250 170.100 ;
        RECT 534.450 168.600 536.250 169.200 ;
        RECT 537.150 168.600 539.850 170.400 ;
        RECT 517.950 166.500 522.750 168.600 ;
        RECT 525.450 167.550 527.250 168.300 ;
        RECT 530.250 167.550 532.050 168.300 ;
        RECT 525.450 166.500 532.050 167.550 ;
        RECT 521.550 165.600 522.750 166.500 ;
        RECT 516.150 159.000 517.950 165.600 ;
        RECT 521.550 159.600 523.350 165.600 ;
        RECT 526.350 159.000 528.150 165.600 ;
        RECT 529.350 159.600 531.150 166.500 ;
        RECT 537.150 165.600 541.050 167.700 ;
        RECT 532.950 159.000 534.750 165.600 ;
        RECT 537.150 159.600 538.950 165.600 ;
        RECT 541.650 159.000 543.450 162.600 ;
        RECT 544.650 159.600 546.450 171.600 ;
        RECT 554.400 159.000 556.200 171.600 ;
        RECT 557.700 170.400 561.300 171.600 ;
        RECT 559.500 159.600 561.300 170.400 ;
        RECT 572.400 159.000 574.200 171.600 ;
        RECT 575.400 159.600 577.200 172.500 ;
        RECT 578.400 159.000 580.200 171.600 ;
        RECT 581.400 159.600 583.200 172.500 ;
        RECT 584.400 159.000 586.200 171.600 ;
        RECT 587.400 159.600 589.200 172.500 ;
        RECT 590.400 159.000 592.200 171.600 ;
        RECT 593.400 159.600 595.200 172.500 ;
        RECT 596.400 159.000 598.200 171.600 ;
        RECT 614.400 165.600 615.600 179.100 ;
        RECT 629.100 177.300 630.900 179.100 ;
        RECT 635.700 171.600 636.600 179.100 ;
        RECT 649.950 178.950 652.050 181.050 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 655.950 178.950 658.050 181.050 ;
        RECT 659.550 179.250 665.850 181.050 ;
        RECT 659.550 178.950 664.050 179.250 ;
        RECT 650.100 177.150 651.900 178.950 ;
        RECT 653.400 171.600 654.300 178.950 ;
        RECT 656.100 177.150 657.900 178.950 ;
        RECT 659.550 171.600 660.750 178.950 ;
        RECT 661.950 173.400 663.750 175.200 ;
        RECT 662.850 172.200 667.050 173.400 ;
        RECT 672.150 172.200 673.050 184.800 ;
        RECT 683.100 183.600 690.000 184.800 ;
        RECT 683.100 183.000 684.900 183.600 ;
        RECT 689.100 182.850 690.000 183.600 ;
        RECT 686.100 181.800 687.900 182.400 ;
        RECT 679.950 180.600 687.900 181.800 ;
        RECT 689.100 181.050 690.900 182.850 ;
        RECT 679.950 178.950 682.050 180.600 ;
        RECT 688.950 178.950 691.050 181.050 ;
        RECT 681.750 173.700 683.550 174.000 ;
        RECT 691.950 173.700 692.850 188.400 ;
        RECT 704.400 187.200 706.200 194.400 ;
        RECT 709.500 188.400 711.300 195.000 ;
        RECT 721.800 188.400 723.600 194.400 ;
        RECT 704.400 186.300 708.600 187.200 ;
        RECT 699.000 183.450 703.050 184.050 ;
        RECT 698.550 181.950 703.050 183.450 ;
        RECT 698.550 177.450 699.450 181.950 ;
        RECT 704.100 181.200 705.900 183.000 ;
        RECT 707.400 181.200 708.600 186.300 ;
        RECT 722.400 186.300 723.600 188.400 ;
        RECT 724.800 189.300 726.600 194.400 ;
        RECT 727.800 190.200 729.600 195.000 ;
        RECT 730.800 189.300 732.600 194.400 ;
        RECT 724.800 187.950 732.600 189.300 ;
        RECT 742.800 188.400 744.600 194.400 ;
        RECT 743.400 186.300 744.600 188.400 ;
        RECT 745.800 189.300 747.600 194.400 ;
        RECT 748.800 190.200 750.600 195.000 ;
        RECT 751.800 189.300 753.600 194.400 ;
        RECT 745.800 187.950 753.600 189.300 ;
        RECT 761.400 186.600 763.200 194.400 ;
        RECT 765.900 188.400 767.700 195.000 ;
        RECT 768.900 190.200 770.700 194.400 ;
        RECT 768.900 188.400 771.600 190.200 ;
        RECT 784.800 188.400 786.600 194.400 ;
        RECT 767.100 186.600 768.900 187.500 ;
        RECT 722.400 185.250 726.150 186.300 ;
        RECT 743.400 185.250 747.150 186.300 ;
        RECT 761.400 185.700 768.900 186.600 ;
        RECT 710.100 181.200 711.900 183.000 ;
        RECT 703.950 179.100 706.050 181.200 ;
        RECT 706.950 179.100 709.050 181.200 ;
        RECT 709.950 179.100 712.050 181.200 ;
        RECT 722.100 181.050 723.900 182.850 ;
        RECT 724.950 181.050 726.150 185.250 ;
        RECT 728.100 181.050 729.900 182.850 ;
        RECT 743.100 181.050 744.900 182.850 ;
        RECT 745.950 181.050 747.150 185.250 ;
        RECT 749.100 181.050 750.900 182.850 ;
        RECT 761.100 181.200 762.900 183.000 ;
        RECT 703.950 177.450 706.050 178.050 ;
        RECT 698.550 176.550 706.050 177.450 ;
        RECT 703.950 175.950 706.050 176.550 ;
        RECT 681.750 173.100 692.850 173.700 ;
        RECT 626.400 170.700 634.200 171.600 ;
        RECT 610.800 159.000 612.600 165.600 ;
        RECT 613.800 159.600 615.600 165.600 ;
        RECT 616.800 159.000 618.600 165.600 ;
        RECT 626.400 159.600 628.200 170.700 ;
        RECT 629.400 159.000 631.200 169.800 ;
        RECT 632.400 159.600 634.200 170.700 ;
        RECT 635.400 159.600 637.200 171.600 ;
        RECT 650.700 170.400 654.300 171.600 ;
        RECT 650.700 159.600 652.500 170.400 ;
        RECT 655.800 159.000 657.600 171.600 ;
        RECT 659.550 159.600 661.350 171.600 ;
        RECT 664.950 171.300 667.050 172.200 ;
        RECT 667.950 171.300 673.050 172.200 ;
        RECT 675.150 172.500 692.850 173.100 ;
        RECT 675.150 172.200 683.550 172.500 ;
        RECT 667.950 170.400 668.850 171.300 ;
        RECT 666.150 168.600 668.850 170.400 ;
        RECT 669.750 170.100 671.550 170.400 ;
        RECT 675.150 170.100 676.050 172.200 ;
        RECT 691.950 171.600 692.850 172.500 ;
        RECT 669.750 169.200 676.050 170.100 ;
        RECT 676.950 170.700 678.750 171.300 ;
        RECT 676.950 169.500 684.450 170.700 ;
        RECT 669.750 168.600 671.550 169.200 ;
        RECT 683.250 168.600 684.450 169.500 ;
        RECT 664.950 165.600 668.850 167.700 ;
        RECT 673.950 167.550 675.750 168.300 ;
        RECT 678.750 167.550 680.550 168.300 ;
        RECT 673.950 166.500 680.550 167.550 ;
        RECT 683.250 166.500 688.050 168.600 ;
        RECT 662.550 159.000 664.350 162.600 ;
        RECT 667.050 159.600 668.850 165.600 ;
        RECT 671.250 159.000 673.050 165.600 ;
        RECT 674.850 159.600 676.650 166.500 ;
        RECT 683.250 165.600 684.450 166.500 ;
        RECT 677.850 159.000 679.650 165.600 ;
        RECT 682.650 159.600 684.450 165.600 ;
        RECT 688.050 159.000 689.850 165.600 ;
        RECT 691.050 159.600 692.850 171.600 ;
        RECT 707.400 165.600 708.600 179.100 ;
        RECT 715.950 178.050 718.050 181.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 727.950 178.950 730.050 181.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 742.950 178.950 745.050 181.050 ;
        RECT 745.950 178.950 748.050 181.050 ;
        RECT 748.950 178.950 751.050 181.050 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 760.950 179.100 763.050 181.200 ;
        RECT 715.950 177.000 721.050 178.050 ;
        RECT 716.550 176.550 721.050 177.000 ;
        RECT 717.000 175.950 721.050 176.550 ;
        RECT 725.850 165.600 727.050 178.950 ;
        RECT 731.100 177.150 732.900 178.950 ;
        RECT 703.800 159.000 705.600 165.600 ;
        RECT 706.800 159.600 708.600 165.600 ;
        RECT 709.800 159.000 711.600 165.600 ;
        RECT 722.400 159.000 724.200 165.600 ;
        RECT 725.400 159.600 727.200 165.600 ;
        RECT 730.500 159.000 732.300 171.600 ;
        RECT 736.950 171.450 739.050 175.050 ;
        RECT 742.950 171.450 745.050 171.900 ;
        RECT 736.950 171.000 745.050 171.450 ;
        RECT 737.550 170.550 745.050 171.000 ;
        RECT 742.950 169.800 745.050 170.550 ;
        RECT 746.850 165.600 748.050 178.950 ;
        RECT 752.100 177.150 753.900 178.950 ;
        RECT 743.400 159.000 745.200 165.600 ;
        RECT 746.400 159.600 748.200 165.600 ;
        RECT 751.500 159.000 753.300 171.600 ;
        RECT 764.400 165.600 765.300 185.700 ;
        RECT 770.700 181.200 771.600 188.400 ;
        RECT 785.400 186.300 786.600 188.400 ;
        RECT 787.800 189.300 789.600 194.400 ;
        RECT 790.800 190.200 792.600 195.000 ;
        RECT 793.800 189.300 795.600 194.400 ;
        RECT 787.800 187.950 795.600 189.300 ;
        RECT 798.150 188.400 799.950 194.400 ;
        RECT 801.150 191.400 802.950 195.000 ;
        RECT 805.950 192.300 807.750 194.400 ;
        RECT 804.000 191.400 807.750 192.300 ;
        RECT 810.450 191.400 812.250 195.000 ;
        RECT 813.750 191.400 815.550 194.400 ;
        RECT 817.350 191.400 819.150 195.000 ;
        RECT 821.550 191.400 823.350 194.400 ;
        RECT 826.350 191.400 828.150 195.000 ;
        RECT 804.000 190.500 805.050 191.400 ;
        RECT 813.750 190.500 814.800 191.400 ;
        RECT 802.950 188.400 805.050 190.500 ;
        RECT 785.400 185.250 789.150 186.300 ;
        RECT 780.000 183.450 784.050 184.050 ;
        RECT 779.550 181.950 784.050 183.450 ;
        RECT 766.950 179.100 769.050 181.200 ;
        RECT 769.950 179.100 772.050 181.200 ;
        RECT 767.100 177.300 768.900 179.100 ;
        RECT 770.700 171.600 771.600 179.100 ;
        RECT 779.550 178.050 780.450 181.950 ;
        RECT 785.100 181.050 786.900 182.850 ;
        RECT 787.950 181.050 789.150 185.250 ;
        RECT 791.100 181.050 792.900 182.850 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 793.950 178.950 796.050 181.050 ;
        RECT 779.550 176.550 784.050 178.050 ;
        RECT 780.000 175.950 784.050 176.550 ;
        RECT 772.950 174.450 775.050 175.050 ;
        RECT 784.950 174.450 787.050 175.050 ;
        RECT 772.950 173.550 787.050 174.450 ;
        RECT 772.950 172.950 775.050 173.550 ;
        RECT 784.950 172.950 787.050 173.550 ;
        RECT 761.400 159.000 763.200 165.600 ;
        RECT 764.400 159.600 766.200 165.600 ;
        RECT 767.400 159.000 769.200 165.600 ;
        RECT 770.400 159.600 772.200 171.600 ;
        RECT 788.850 165.600 790.050 178.950 ;
        RECT 794.100 177.150 795.900 178.950 ;
        RECT 798.150 173.700 799.050 188.400 ;
        RECT 806.550 187.800 808.350 189.600 ;
        RECT 809.850 189.450 814.800 190.500 ;
        RECT 822.300 190.500 823.350 191.400 ;
        RECT 809.850 188.700 811.650 189.450 ;
        RECT 822.300 189.300 826.050 190.500 ;
        RECT 823.950 188.400 826.050 189.300 ;
        RECT 829.650 188.400 831.450 194.400 ;
        RECT 839.400 191.400 841.200 195.000 ;
        RECT 842.400 191.400 844.200 194.400 ;
        RECT 806.850 186.000 807.900 187.800 ;
        RECT 817.050 186.000 818.850 186.600 ;
        RECT 806.850 184.800 818.850 186.000 ;
        RECT 801.000 183.600 807.900 184.800 ;
        RECT 801.000 182.850 801.900 183.600 ;
        RECT 806.100 183.000 807.900 183.600 ;
        RECT 800.100 181.050 801.900 182.850 ;
        RECT 803.100 181.800 804.900 182.400 ;
        RECT 799.950 178.950 802.050 181.050 ;
        RECT 803.100 180.600 811.050 181.800 ;
        RECT 808.950 178.950 811.050 180.600 ;
        RECT 807.450 173.700 809.250 174.000 ;
        RECT 798.150 173.100 809.250 173.700 ;
        RECT 798.150 172.500 815.850 173.100 ;
        RECT 798.150 171.600 799.050 172.500 ;
        RECT 807.450 172.200 815.850 172.500 ;
        RECT 785.400 159.000 787.200 165.600 ;
        RECT 788.400 159.600 790.200 165.600 ;
        RECT 793.500 159.000 795.300 171.600 ;
        RECT 798.150 159.600 799.950 171.600 ;
        RECT 812.250 170.700 814.050 171.300 ;
        RECT 806.550 169.500 814.050 170.700 ;
        RECT 814.950 170.100 815.850 172.200 ;
        RECT 817.950 172.200 818.850 184.800 ;
        RECT 830.250 181.050 831.450 188.400 ;
        RECT 842.400 181.050 843.600 191.400 ;
        RECT 825.150 179.250 831.450 181.050 ;
        RECT 826.950 178.950 831.450 179.250 ;
        RECT 838.950 178.950 841.050 181.050 ;
        RECT 841.950 178.950 844.050 181.050 ;
        RECT 827.250 173.400 829.050 175.200 ;
        RECT 823.950 172.200 828.150 173.400 ;
        RECT 817.950 171.300 823.050 172.200 ;
        RECT 823.950 171.300 826.050 172.200 ;
        RECT 830.250 171.600 831.450 178.950 ;
        RECT 839.100 177.150 840.900 178.950 ;
        RECT 822.150 170.400 823.050 171.300 ;
        RECT 819.450 170.100 821.250 170.400 ;
        RECT 806.550 168.600 807.750 169.500 ;
        RECT 814.950 169.200 821.250 170.100 ;
        RECT 819.450 168.600 821.250 169.200 ;
        RECT 822.150 168.600 824.850 170.400 ;
        RECT 802.950 166.500 807.750 168.600 ;
        RECT 810.450 167.550 812.250 168.300 ;
        RECT 815.250 167.550 817.050 168.300 ;
        RECT 810.450 166.500 817.050 167.550 ;
        RECT 806.550 165.600 807.750 166.500 ;
        RECT 801.150 159.000 802.950 165.600 ;
        RECT 806.550 159.600 808.350 165.600 ;
        RECT 811.350 159.000 813.150 165.600 ;
        RECT 814.350 159.600 816.150 166.500 ;
        RECT 822.150 165.600 826.050 167.700 ;
        RECT 817.950 159.000 819.750 165.600 ;
        RECT 822.150 159.600 823.950 165.600 ;
        RECT 826.650 159.000 828.450 162.600 ;
        RECT 829.650 159.600 831.450 171.600 ;
        RECT 842.400 165.600 843.600 178.950 ;
        RECT 839.400 159.000 841.200 165.600 ;
        RECT 842.400 159.600 844.200 165.600 ;
        RECT 11.700 144.600 13.500 155.400 ;
        RECT 11.700 143.400 15.300 144.600 ;
        RECT 16.800 143.400 18.600 156.000 ;
        RECT 29.700 144.600 31.500 155.400 ;
        RECT 29.700 143.400 33.300 144.600 ;
        RECT 34.800 143.400 36.600 156.000 ;
        RECT 47.700 144.600 49.500 155.400 ;
        RECT 47.700 143.400 51.300 144.600 ;
        RECT 52.800 143.400 54.600 156.000 ;
        RECT 62.400 149.400 64.200 156.000 ;
        RECT 65.400 149.400 67.200 155.400 ;
        RECT 11.100 136.050 12.900 137.850 ;
        RECT 14.400 136.050 15.300 143.400 ;
        RECT 17.100 136.050 18.900 137.850 ;
        RECT 29.100 136.050 30.900 137.850 ;
        RECT 32.400 136.050 33.300 143.400 ;
        RECT 35.100 136.050 36.900 137.850 ;
        RECT 47.100 136.050 48.900 137.850 ;
        RECT 50.400 136.050 51.300 143.400 ;
        RECT 53.100 136.050 54.900 137.850 ;
        RECT 62.100 136.050 63.900 137.850 ;
        RECT 65.400 136.050 66.600 149.400 ;
        RECT 77.700 143.400 79.500 156.000 ;
        RECT 82.800 149.400 84.600 155.400 ;
        RECT 85.800 149.400 87.600 156.000 ;
        RECT 77.100 136.050 78.900 137.850 ;
        RECT 82.950 136.050 84.150 149.400 ;
        RECT 98.400 144.300 100.200 155.400 ;
        RECT 98.400 143.400 102.900 144.300 ;
        RECT 105.900 143.400 107.700 155.400 ;
        RECT 113.400 144.600 115.200 155.400 ;
        RECT 100.800 141.300 102.900 143.400 ;
        RECT 106.500 141.900 107.700 143.400 ;
        RECT 110.400 143.400 115.200 144.600 ;
        RECT 125.400 149.400 127.200 155.400 ;
        RECT 128.400 149.400 130.200 156.000 ;
        RECT 110.400 142.500 112.500 143.400 ;
        RECT 125.400 142.500 126.600 149.400 ;
        RECT 131.400 143.400 133.200 155.400 ;
        RECT 143.700 143.400 145.500 156.000 ;
        RECT 148.800 149.400 150.600 155.400 ;
        RECT 151.800 149.400 153.600 156.000 ;
        RECT 106.500 141.000 108.000 141.900 ;
        RECT 103.950 139.500 106.050 139.800 ;
        RECT 88.950 138.450 93.000 139.050 ;
        RECT 88.950 136.950 93.450 138.450 ;
        RECT 102.300 137.700 106.050 139.500 ;
        RECT 107.100 138.900 108.000 141.000 ;
        RECT 115.950 141.450 120.000 142.050 ;
        RECT 125.400 141.600 131.100 142.500 ;
        RECT 115.950 139.950 120.450 141.450 ;
        RECT 114.000 138.900 117.000 139.050 ;
        RECT 10.950 133.950 13.050 136.050 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 28.950 133.950 31.050 136.050 ;
        RECT 31.950 133.950 34.050 136.050 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 46.950 133.950 49.050 136.050 ;
        RECT 49.950 133.950 52.050 136.050 ;
        RECT 52.950 133.950 55.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 14.400 123.600 15.300 133.950 ;
        RECT 32.400 123.600 33.300 133.950 ;
        RECT 50.400 123.600 51.300 133.950 ;
        RECT 65.400 123.600 66.600 133.950 ;
        RECT 80.100 132.150 81.900 133.950 ;
        RECT 83.850 129.750 85.050 133.950 ;
        RECT 86.100 132.150 87.900 133.950 ;
        RECT 92.550 133.050 93.450 136.950 ;
        RECT 106.950 136.800 109.050 138.900 ;
        RECT 114.000 138.450 118.050 138.900 ;
        RECT 113.550 137.700 118.050 138.450 ;
        RECT 113.100 136.950 118.050 137.700 ;
        RECT 103.500 135.900 105.300 136.500 ;
        RECT 97.950 134.700 105.300 135.900 ;
        RECT 106.200 135.900 108.600 136.800 ;
        RECT 113.100 135.900 114.900 136.950 ;
        RECT 115.950 136.800 118.050 136.950 ;
        RECT 97.950 133.800 100.050 134.700 ;
        RECT 88.950 131.550 93.450 133.050 ;
        RECT 98.250 132.000 100.050 133.800 ;
        RECT 88.950 130.950 93.000 131.550 ;
        RECT 103.500 131.400 105.300 133.200 ;
        RECT 83.850 128.700 87.600 129.750 ;
        RECT 103.200 129.300 105.300 131.400 ;
        RECT 77.400 125.700 85.200 127.050 ;
        RECT 10.800 120.000 12.600 123.600 ;
        RECT 13.800 120.600 15.600 123.600 ;
        RECT 16.800 120.000 18.600 123.600 ;
        RECT 28.800 120.000 30.600 123.600 ;
        RECT 31.800 120.600 33.600 123.600 ;
        RECT 34.800 120.000 36.600 123.600 ;
        RECT 46.800 120.000 48.600 123.600 ;
        RECT 49.800 120.600 51.600 123.600 ;
        RECT 52.800 120.000 54.600 123.600 ;
        RECT 62.400 120.000 64.200 123.600 ;
        RECT 65.400 120.600 67.200 123.600 ;
        RECT 77.400 120.600 79.200 125.700 ;
        RECT 80.400 120.000 82.200 124.800 ;
        RECT 83.400 120.600 85.200 125.700 ;
        RECT 86.400 126.600 87.600 128.700 ;
        RECT 99.000 128.400 105.300 129.300 ;
        RECT 106.200 130.200 107.250 135.900 ;
        RECT 108.600 133.200 110.400 135.000 ;
        RECT 112.950 133.800 115.050 135.900 ;
        RECT 108.150 131.100 110.250 133.200 ;
        RECT 119.550 133.050 120.450 139.950 ;
        RECT 129.150 140.700 131.100 141.600 ;
        RECT 125.100 136.050 126.900 137.850 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 119.550 131.550 124.050 133.050 ;
        RECT 120.000 130.950 124.050 131.550 ;
        RECT 99.000 126.600 100.200 128.400 ;
        RECT 106.200 128.100 109.050 130.200 ;
        RECT 129.150 129.300 130.050 140.700 ;
        RECT 132.000 136.050 133.200 143.400 ;
        RECT 139.950 138.450 142.050 142.050 ;
        RECT 130.950 133.950 133.200 136.050 ;
        RECT 106.200 126.600 107.400 128.100 ;
        RECT 110.400 127.500 112.500 128.700 ;
        RECT 129.150 128.400 131.100 129.300 ;
        RECT 125.400 127.500 131.100 128.400 ;
        RECT 110.400 126.600 115.200 127.500 ;
        RECT 86.400 120.600 88.200 126.600 ;
        RECT 98.400 120.600 100.200 126.600 ;
        RECT 105.900 120.600 107.700 126.600 ;
        RECT 113.400 120.600 115.200 126.600 ;
        RECT 125.400 123.600 126.600 127.500 ;
        RECT 132.000 126.600 133.200 133.950 ;
        RECT 137.550 138.000 142.050 138.450 ;
        RECT 137.550 137.550 141.450 138.000 ;
        RECT 137.550 130.050 138.450 137.550 ;
        RECT 143.100 136.050 144.900 137.850 ;
        RECT 148.950 136.050 150.150 149.400 ;
        RECT 159.150 143.400 160.950 155.400 ;
        RECT 162.150 149.400 163.950 156.000 ;
        RECT 167.550 149.400 169.350 155.400 ;
        RECT 172.350 149.400 174.150 156.000 ;
        RECT 167.550 148.500 168.750 149.400 ;
        RECT 175.350 148.500 177.150 155.400 ;
        RECT 178.950 149.400 180.750 156.000 ;
        RECT 183.150 149.400 184.950 155.400 ;
        RECT 187.650 152.400 189.450 156.000 ;
        RECT 163.950 146.400 168.750 148.500 ;
        RECT 171.450 147.450 178.050 148.500 ;
        RECT 171.450 146.700 173.250 147.450 ;
        RECT 176.250 146.700 178.050 147.450 ;
        RECT 183.150 147.300 187.050 149.400 ;
        RECT 167.550 145.500 168.750 146.400 ;
        RECT 180.450 145.800 182.250 146.400 ;
        RECT 167.550 144.300 175.050 145.500 ;
        RECT 173.250 143.700 175.050 144.300 ;
        RECT 175.950 144.900 182.250 145.800 ;
        RECT 159.150 142.500 160.050 143.400 ;
        RECT 175.950 142.800 176.850 144.900 ;
        RECT 180.450 144.600 182.250 144.900 ;
        RECT 183.150 144.600 185.850 146.400 ;
        RECT 183.150 143.700 184.050 144.600 ;
        RECT 168.450 142.500 176.850 142.800 ;
        RECT 159.150 141.900 176.850 142.500 ;
        RECT 178.950 142.800 184.050 143.700 ;
        RECT 184.950 142.800 187.050 143.700 ;
        RECT 190.650 143.400 192.450 155.400 ;
        RECT 200.400 149.400 202.200 156.000 ;
        RECT 203.400 149.400 205.200 155.400 ;
        RECT 206.400 149.400 208.200 156.000 ;
        RECT 159.150 141.300 170.250 141.900 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 146.100 132.150 147.900 133.950 ;
        RECT 136.950 127.950 139.050 130.050 ;
        RECT 149.850 129.750 151.050 133.950 ;
        RECT 152.100 132.150 153.900 133.950 ;
        RECT 149.850 128.700 153.600 129.750 ;
        RECT 125.400 120.600 127.200 123.600 ;
        RECT 128.400 120.000 130.200 123.600 ;
        RECT 131.400 120.600 133.200 126.600 ;
        RECT 143.400 125.700 151.200 127.050 ;
        RECT 143.400 120.600 145.200 125.700 ;
        RECT 146.400 120.000 148.200 124.800 ;
        RECT 149.400 120.600 151.200 125.700 ;
        RECT 152.400 126.600 153.600 128.700 ;
        RECT 159.150 126.600 160.050 141.300 ;
        RECT 168.450 141.000 170.250 141.300 ;
        RECT 160.950 133.950 163.050 136.050 ;
        RECT 169.950 134.400 172.050 136.050 ;
        RECT 161.100 132.150 162.900 133.950 ;
        RECT 164.100 133.200 172.050 134.400 ;
        RECT 164.100 132.600 165.900 133.200 ;
        RECT 162.000 131.400 162.900 132.150 ;
        RECT 167.100 131.400 168.900 132.000 ;
        RECT 162.000 130.200 168.900 131.400 ;
        RECT 178.950 130.200 179.850 142.800 ;
        RECT 184.950 141.600 189.150 142.800 ;
        RECT 188.250 139.800 190.050 141.600 ;
        RECT 191.250 136.050 192.450 143.400 ;
        RECT 187.950 135.750 192.450 136.050 ;
        RECT 203.400 135.900 204.600 149.400 ;
        RECT 218.700 143.400 220.500 156.000 ;
        RECT 223.800 149.400 225.600 155.400 ;
        RECT 226.800 149.400 228.600 156.000 ;
        RECT 242.400 149.400 244.200 156.000 ;
        RECT 245.400 149.400 247.200 155.400 ;
        RECT 208.950 138.450 213.000 139.050 ;
        RECT 208.950 136.950 213.450 138.450 ;
        RECT 186.150 133.950 192.450 135.750 ;
        RECT 167.850 129.000 179.850 130.200 ;
        RECT 167.850 127.200 168.900 129.000 ;
        RECT 178.050 128.400 179.850 129.000 ;
        RECT 152.400 120.600 154.200 126.600 ;
        RECT 159.150 120.600 160.950 126.600 ;
        RECT 163.950 124.500 166.050 126.600 ;
        RECT 167.550 125.400 169.350 127.200 ;
        RECT 191.250 126.600 192.450 133.950 ;
        RECT 199.950 133.800 202.050 135.900 ;
        RECT 202.950 133.800 205.050 135.900 ;
        RECT 205.950 133.800 208.050 135.900 ;
        RECT 200.100 132.000 201.900 133.800 ;
        RECT 203.400 128.700 204.600 133.800 ;
        RECT 206.100 132.000 207.900 133.800 ;
        RECT 212.550 133.050 213.450 136.950 ;
        RECT 218.100 136.050 219.900 137.850 ;
        RECT 223.950 136.050 225.150 149.400 ;
        RECT 245.850 136.050 247.050 149.400 ;
        RECT 250.500 143.400 252.300 156.000 ;
        RECT 263.400 149.400 265.200 156.000 ;
        RECT 266.400 149.400 268.200 155.400 ;
        RECT 251.100 136.050 252.900 137.850 ;
        RECT 266.850 136.050 268.050 149.400 ;
        RECT 271.500 143.400 273.300 156.000 ;
        RECT 276.150 143.400 277.950 155.400 ;
        RECT 279.150 149.400 280.950 156.000 ;
        RECT 284.550 149.400 286.350 155.400 ;
        RECT 289.350 149.400 291.150 156.000 ;
        RECT 284.550 148.500 285.750 149.400 ;
        RECT 292.350 148.500 294.150 155.400 ;
        RECT 295.950 149.400 297.750 156.000 ;
        RECT 300.150 149.400 301.950 155.400 ;
        RECT 304.650 152.400 306.450 156.000 ;
        RECT 280.950 146.400 285.750 148.500 ;
        RECT 288.450 147.450 295.050 148.500 ;
        RECT 288.450 146.700 290.250 147.450 ;
        RECT 293.250 146.700 295.050 147.450 ;
        RECT 300.150 147.300 304.050 149.400 ;
        RECT 284.550 145.500 285.750 146.400 ;
        RECT 297.450 145.800 299.250 146.400 ;
        RECT 284.550 144.300 292.050 145.500 ;
        RECT 290.250 143.700 292.050 144.300 ;
        RECT 292.950 144.900 299.250 145.800 ;
        RECT 276.150 142.500 277.050 143.400 ;
        RECT 292.950 142.800 293.850 144.900 ;
        RECT 297.450 144.600 299.250 144.900 ;
        RECT 300.150 144.600 302.850 146.400 ;
        RECT 300.150 143.700 301.050 144.600 ;
        RECT 285.450 142.500 293.850 142.800 ;
        RECT 276.150 141.900 293.850 142.500 ;
        RECT 295.950 142.800 301.050 143.700 ;
        RECT 301.950 142.800 304.050 143.700 ;
        RECT 307.650 143.400 309.450 155.400 ;
        RECT 317.400 149.400 319.200 156.000 ;
        RECT 320.400 149.400 322.200 155.400 ;
        RECT 323.400 149.400 325.200 156.000 ;
        RECT 276.150 141.300 287.250 141.900 ;
        RECT 272.100 136.050 273.900 137.850 ;
        RECT 217.950 133.950 220.050 136.050 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 250.950 133.950 253.050 136.050 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 208.950 131.550 213.450 133.050 ;
        RECT 221.100 132.150 222.900 133.950 ;
        RECT 208.950 130.950 213.000 131.550 ;
        RECT 224.850 129.750 226.050 133.950 ;
        RECT 227.100 132.150 228.900 133.950 ;
        RECT 242.100 132.150 243.900 133.950 ;
        RECT 244.950 129.750 246.150 133.950 ;
        RECT 248.100 132.150 249.900 133.950 ;
        RECT 263.100 132.150 264.900 133.950 ;
        RECT 265.950 129.750 267.150 133.950 ;
        RECT 269.100 132.150 270.900 133.950 ;
        RECT 224.850 128.700 228.600 129.750 ;
        RECT 203.400 127.800 207.600 128.700 ;
        RECT 170.850 125.550 172.650 126.300 ;
        RECT 184.950 125.700 187.050 126.600 ;
        RECT 170.850 124.500 175.800 125.550 ;
        RECT 165.000 123.600 166.050 124.500 ;
        RECT 174.750 123.600 175.800 124.500 ;
        RECT 183.300 124.500 187.050 125.700 ;
        RECT 183.300 123.600 184.350 124.500 ;
        RECT 162.150 120.000 163.950 123.600 ;
        RECT 165.000 122.700 168.750 123.600 ;
        RECT 166.950 120.600 168.750 122.700 ;
        RECT 171.450 120.000 173.250 123.600 ;
        RECT 174.750 120.600 176.550 123.600 ;
        RECT 178.350 120.000 180.150 123.600 ;
        RECT 182.550 120.600 184.350 123.600 ;
        RECT 187.350 120.000 189.150 123.600 ;
        RECT 190.650 120.600 192.450 126.600 ;
        RECT 200.700 120.000 202.500 126.600 ;
        RECT 205.800 120.600 207.600 127.800 ;
        RECT 218.400 125.700 226.200 127.050 ;
        RECT 218.400 120.600 220.200 125.700 ;
        RECT 221.400 120.000 223.200 124.800 ;
        RECT 224.400 120.600 226.200 125.700 ;
        RECT 227.400 126.600 228.600 128.700 ;
        RECT 242.400 128.700 246.150 129.750 ;
        RECT 263.400 128.700 267.150 129.750 ;
        RECT 242.400 126.600 243.600 128.700 ;
        RECT 227.400 120.600 229.200 126.600 ;
        RECT 241.800 120.600 243.600 126.600 ;
        RECT 244.800 125.700 252.600 127.050 ;
        RECT 263.400 126.600 264.600 128.700 ;
        RECT 244.800 120.600 246.600 125.700 ;
        RECT 247.800 120.000 249.600 124.800 ;
        RECT 250.800 120.600 252.600 125.700 ;
        RECT 262.800 120.600 264.600 126.600 ;
        RECT 265.800 125.700 273.600 127.050 ;
        RECT 265.800 120.600 267.600 125.700 ;
        RECT 268.800 120.000 270.600 124.800 ;
        RECT 271.800 120.600 273.600 125.700 ;
        RECT 276.150 126.600 277.050 141.300 ;
        RECT 285.450 141.000 287.250 141.300 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 286.950 134.400 289.050 136.050 ;
        RECT 278.100 132.150 279.900 133.950 ;
        RECT 281.100 133.200 289.050 134.400 ;
        RECT 281.100 132.600 282.900 133.200 ;
        RECT 279.000 131.400 279.900 132.150 ;
        RECT 284.100 131.400 285.900 132.000 ;
        RECT 279.000 130.200 285.900 131.400 ;
        RECT 295.950 130.200 296.850 142.800 ;
        RECT 301.950 141.600 306.150 142.800 ;
        RECT 305.250 139.800 307.050 141.600 ;
        RECT 308.250 136.050 309.450 143.400 ;
        RECT 310.950 138.450 313.050 139.050 ;
        RECT 316.950 138.450 319.050 139.050 ;
        RECT 310.950 137.550 319.050 138.450 ;
        RECT 310.950 136.950 313.050 137.550 ;
        RECT 316.950 136.950 319.050 137.550 ;
        RECT 304.950 135.750 309.450 136.050 ;
        RECT 320.400 135.900 321.600 149.400 ;
        RECT 335.400 144.600 337.200 155.400 ;
        RECT 338.400 145.500 340.200 156.000 ;
        RECT 341.400 154.500 349.200 155.400 ;
        RECT 341.400 144.600 343.200 154.500 ;
        RECT 335.400 143.700 343.200 144.600 ;
        RECT 344.400 142.500 346.200 153.600 ;
        RECT 347.400 143.400 349.200 154.500 ;
        RECT 361.800 143.400 363.600 155.400 ;
        RECT 364.800 149.400 366.600 156.000 ;
        RECT 367.800 149.400 369.600 155.400 ;
        RECT 341.100 141.600 346.200 142.500 ;
        RECT 322.950 138.450 325.050 139.050 ;
        RECT 328.950 138.450 331.050 139.050 ;
        RECT 322.950 137.550 331.050 138.450 ;
        RECT 322.950 136.950 325.050 137.550 ;
        RECT 328.950 136.950 331.050 137.550 ;
        RECT 338.100 135.900 339.900 137.700 ;
        RECT 341.100 135.900 342.000 141.600 ;
        RECT 349.950 138.450 354.000 139.050 ;
        RECT 344.100 135.900 345.900 137.700 ;
        RECT 349.950 136.950 354.450 138.450 ;
        RECT 303.150 133.950 309.450 135.750 ;
        RECT 284.850 129.000 296.850 130.200 ;
        RECT 284.850 127.200 285.900 129.000 ;
        RECT 295.050 128.400 296.850 129.000 ;
        RECT 276.150 120.600 277.950 126.600 ;
        RECT 280.950 124.500 283.050 126.600 ;
        RECT 284.550 125.400 286.350 127.200 ;
        RECT 308.250 126.600 309.450 133.950 ;
        RECT 316.950 133.800 319.050 135.900 ;
        RECT 319.950 133.800 322.050 135.900 ;
        RECT 322.950 133.800 325.050 135.900 ;
        RECT 334.950 133.800 337.050 135.900 ;
        RECT 337.950 133.800 340.050 135.900 ;
        RECT 340.950 133.800 343.050 135.900 ;
        RECT 343.950 133.800 346.050 135.900 ;
        RECT 346.950 133.800 349.050 135.900 ;
        RECT 317.100 132.000 318.900 133.800 ;
        RECT 320.400 128.700 321.600 133.800 ;
        RECT 323.100 132.000 324.900 133.800 ;
        RECT 335.100 132.000 336.900 133.800 ;
        RECT 320.400 127.800 324.600 128.700 ;
        RECT 287.850 125.550 289.650 126.300 ;
        RECT 301.950 125.700 304.050 126.600 ;
        RECT 287.850 124.500 292.800 125.550 ;
        RECT 282.000 123.600 283.050 124.500 ;
        RECT 291.750 123.600 292.800 124.500 ;
        RECT 300.300 124.500 304.050 125.700 ;
        RECT 300.300 123.600 301.350 124.500 ;
        RECT 279.150 120.000 280.950 123.600 ;
        RECT 282.000 122.700 285.750 123.600 ;
        RECT 283.950 120.600 285.750 122.700 ;
        RECT 288.450 120.000 290.250 123.600 ;
        RECT 291.750 120.600 293.550 123.600 ;
        RECT 295.350 120.000 297.150 123.600 ;
        RECT 299.550 120.600 301.350 123.600 ;
        RECT 304.350 120.000 306.150 123.600 ;
        RECT 307.650 120.600 309.450 126.600 ;
        RECT 317.700 120.000 319.500 126.600 ;
        RECT 322.800 120.600 324.600 127.800 ;
        RECT 340.950 126.600 342.000 133.800 ;
        RECT 347.100 132.000 348.900 133.800 ;
        RECT 353.550 129.900 354.450 136.950 ;
        RECT 361.800 136.050 363.000 143.400 ;
        RECT 368.400 142.500 369.600 149.400 ;
        RECT 363.900 141.600 369.600 142.500 ;
        RECT 379.800 143.400 381.600 155.400 ;
        RECT 382.800 149.400 384.600 156.000 ;
        RECT 385.800 149.400 387.600 155.400 ;
        RECT 363.900 140.700 365.850 141.600 ;
        RECT 361.800 133.950 364.050 136.050 ;
        RECT 352.950 127.800 355.050 129.900 ;
        RECT 361.800 126.600 363.000 133.950 ;
        RECT 364.950 129.300 365.850 140.700 ;
        RECT 370.950 138.450 375.000 139.050 ;
        RECT 368.100 136.050 369.900 137.850 ;
        RECT 370.950 136.950 375.450 138.450 ;
        RECT 367.950 133.950 370.050 136.050 ;
        RECT 374.550 133.050 375.450 136.950 ;
        RECT 370.950 131.550 375.450 133.050 ;
        RECT 379.800 136.050 381.000 143.400 ;
        RECT 386.400 142.500 387.600 149.400 ;
        RECT 381.900 141.600 387.600 142.500 ;
        RECT 390.150 143.400 391.950 155.400 ;
        RECT 393.150 149.400 394.950 156.000 ;
        RECT 398.550 149.400 400.350 155.400 ;
        RECT 403.350 149.400 405.150 156.000 ;
        RECT 398.550 148.500 399.750 149.400 ;
        RECT 406.350 148.500 408.150 155.400 ;
        RECT 409.950 149.400 411.750 156.000 ;
        RECT 414.150 149.400 415.950 155.400 ;
        RECT 418.650 152.400 420.450 156.000 ;
        RECT 394.950 146.400 399.750 148.500 ;
        RECT 402.450 147.450 409.050 148.500 ;
        RECT 402.450 146.700 404.250 147.450 ;
        RECT 407.250 146.700 409.050 147.450 ;
        RECT 414.150 147.300 418.050 149.400 ;
        RECT 398.550 145.500 399.750 146.400 ;
        RECT 411.450 145.800 413.250 146.400 ;
        RECT 398.550 144.300 406.050 145.500 ;
        RECT 404.250 143.700 406.050 144.300 ;
        RECT 406.950 144.900 413.250 145.800 ;
        RECT 390.150 142.500 391.050 143.400 ;
        RECT 406.950 142.800 407.850 144.900 ;
        RECT 411.450 144.600 413.250 144.900 ;
        RECT 414.150 144.600 416.850 146.400 ;
        RECT 414.150 143.700 415.050 144.600 ;
        RECT 399.450 142.500 407.850 142.800 ;
        RECT 390.150 141.900 407.850 142.500 ;
        RECT 409.950 142.800 415.050 143.700 ;
        RECT 415.950 142.800 418.050 143.700 ;
        RECT 421.650 143.400 423.450 155.400 ;
        RECT 433.800 149.400 435.600 156.000 ;
        RECT 436.800 149.400 438.600 155.400 ;
        RECT 439.800 149.400 441.600 156.000 ;
        RECT 381.900 140.700 383.850 141.600 ;
        RECT 379.800 133.950 382.050 136.050 ;
        RECT 370.950 130.950 375.000 131.550 ;
        RECT 363.900 128.400 365.850 129.300 ;
        RECT 363.900 127.500 369.600 128.400 ;
        RECT 335.700 120.000 337.500 126.600 ;
        RECT 340.200 120.600 342.000 126.600 ;
        RECT 344.700 120.000 346.500 126.600 ;
        RECT 361.800 120.600 363.600 126.600 ;
        RECT 368.400 123.600 369.600 127.500 ;
        RECT 364.800 120.000 366.600 123.600 ;
        RECT 367.800 120.600 369.600 123.600 ;
        RECT 379.800 126.600 381.000 133.950 ;
        RECT 382.950 129.300 383.850 140.700 ;
        RECT 390.150 141.300 401.250 141.900 ;
        RECT 386.100 136.050 387.900 137.850 ;
        RECT 385.950 133.950 388.050 136.050 ;
        RECT 381.900 128.400 383.850 129.300 ;
        RECT 381.900 127.500 387.600 128.400 ;
        RECT 379.800 120.600 381.600 126.600 ;
        RECT 386.400 123.600 387.600 127.500 ;
        RECT 382.800 120.000 384.600 123.600 ;
        RECT 385.800 120.600 387.600 123.600 ;
        RECT 390.150 126.600 391.050 141.300 ;
        RECT 399.450 141.000 401.250 141.300 ;
        RECT 391.950 133.950 394.050 136.050 ;
        RECT 400.950 134.400 403.050 136.050 ;
        RECT 392.100 132.150 393.900 133.950 ;
        RECT 395.100 133.200 403.050 134.400 ;
        RECT 395.100 132.600 396.900 133.200 ;
        RECT 393.000 131.400 393.900 132.150 ;
        RECT 398.100 131.400 399.900 132.000 ;
        RECT 393.000 130.200 399.900 131.400 ;
        RECT 409.950 130.200 410.850 142.800 ;
        RECT 415.950 141.600 420.150 142.800 ;
        RECT 419.250 139.800 421.050 141.600 ;
        RECT 422.250 136.050 423.450 143.400 ;
        RECT 418.950 135.750 423.450 136.050 ;
        RECT 437.400 135.900 438.600 149.400 ;
        RECT 444.150 143.400 445.950 155.400 ;
        RECT 447.150 149.400 448.950 156.000 ;
        RECT 452.550 149.400 454.350 155.400 ;
        RECT 457.350 149.400 459.150 156.000 ;
        RECT 452.550 148.500 453.750 149.400 ;
        RECT 460.350 148.500 462.150 155.400 ;
        RECT 463.950 149.400 465.750 156.000 ;
        RECT 468.150 149.400 469.950 155.400 ;
        RECT 472.650 152.400 474.450 156.000 ;
        RECT 448.950 146.400 453.750 148.500 ;
        RECT 456.450 147.450 463.050 148.500 ;
        RECT 456.450 146.700 458.250 147.450 ;
        RECT 461.250 146.700 463.050 147.450 ;
        RECT 468.150 147.300 472.050 149.400 ;
        RECT 452.550 145.500 453.750 146.400 ;
        RECT 465.450 145.800 467.250 146.400 ;
        RECT 452.550 144.300 460.050 145.500 ;
        RECT 458.250 143.700 460.050 144.300 ;
        RECT 460.950 144.900 467.250 145.800 ;
        RECT 444.150 142.500 445.050 143.400 ;
        RECT 460.950 142.800 461.850 144.900 ;
        RECT 465.450 144.600 467.250 144.900 ;
        RECT 468.150 144.600 470.850 146.400 ;
        RECT 468.150 143.700 469.050 144.600 ;
        RECT 453.450 142.500 461.850 142.800 ;
        RECT 444.150 141.900 461.850 142.500 ;
        RECT 463.950 142.800 469.050 143.700 ;
        RECT 469.950 142.800 472.050 143.700 ;
        RECT 475.650 143.400 477.450 155.400 ;
        RECT 488.700 144.600 490.500 155.400 ;
        RECT 488.700 143.400 492.300 144.600 ;
        RECT 493.800 143.400 495.600 156.000 ;
        RECT 503.700 143.400 505.500 156.000 ;
        RECT 508.800 149.400 510.600 155.400 ;
        RECT 511.800 149.400 513.600 156.000 ;
        RECT 444.150 141.300 455.250 141.900 ;
        RECT 417.150 133.950 423.450 135.750 ;
        RECT 398.850 129.000 410.850 130.200 ;
        RECT 398.850 127.200 399.900 129.000 ;
        RECT 409.050 128.400 410.850 129.000 ;
        RECT 390.150 120.600 391.950 126.600 ;
        RECT 394.950 124.500 397.050 126.600 ;
        RECT 398.550 125.400 400.350 127.200 ;
        RECT 422.250 126.600 423.450 133.950 ;
        RECT 433.950 133.800 436.050 135.900 ;
        RECT 436.950 133.800 439.050 135.900 ;
        RECT 439.950 133.800 442.050 135.900 ;
        RECT 434.100 132.000 435.900 133.800 ;
        RECT 437.400 128.700 438.600 133.800 ;
        RECT 440.100 132.000 441.900 133.800 ;
        RECT 401.850 125.550 403.650 126.300 ;
        RECT 415.950 125.700 418.050 126.600 ;
        RECT 401.850 124.500 406.800 125.550 ;
        RECT 396.000 123.600 397.050 124.500 ;
        RECT 405.750 123.600 406.800 124.500 ;
        RECT 414.300 124.500 418.050 125.700 ;
        RECT 414.300 123.600 415.350 124.500 ;
        RECT 393.150 120.000 394.950 123.600 ;
        RECT 396.000 122.700 399.750 123.600 ;
        RECT 397.950 120.600 399.750 122.700 ;
        RECT 402.450 120.000 404.250 123.600 ;
        RECT 405.750 120.600 407.550 123.600 ;
        RECT 409.350 120.000 411.150 123.600 ;
        RECT 413.550 120.600 415.350 123.600 ;
        RECT 418.350 120.000 420.150 123.600 ;
        RECT 421.650 120.600 423.450 126.600 ;
        RECT 434.400 127.800 438.600 128.700 ;
        RECT 434.400 120.600 436.200 127.800 ;
        RECT 444.150 126.600 445.050 141.300 ;
        RECT 453.450 141.000 455.250 141.300 ;
        RECT 445.950 133.950 448.050 136.050 ;
        RECT 454.950 134.400 457.050 136.050 ;
        RECT 446.100 132.150 447.900 133.950 ;
        RECT 449.100 133.200 457.050 134.400 ;
        RECT 449.100 132.600 450.900 133.200 ;
        RECT 447.000 131.400 447.900 132.150 ;
        RECT 452.100 131.400 453.900 132.000 ;
        RECT 447.000 130.200 453.900 131.400 ;
        RECT 463.950 130.200 464.850 142.800 ;
        RECT 469.950 141.600 474.150 142.800 ;
        RECT 473.250 139.800 475.050 141.600 ;
        RECT 476.250 136.050 477.450 143.400 ;
        RECT 488.100 136.050 489.900 137.850 ;
        RECT 491.400 136.050 492.300 143.400 ;
        RECT 494.100 136.050 495.900 137.850 ;
        RECT 503.100 136.050 504.900 137.850 ;
        RECT 508.950 136.050 510.150 149.400 ;
        RECT 519.150 143.400 520.950 155.400 ;
        RECT 522.150 149.400 523.950 156.000 ;
        RECT 527.550 149.400 529.350 155.400 ;
        RECT 532.350 149.400 534.150 156.000 ;
        RECT 527.550 148.500 528.750 149.400 ;
        RECT 535.350 148.500 537.150 155.400 ;
        RECT 538.950 149.400 540.750 156.000 ;
        RECT 543.150 149.400 544.950 155.400 ;
        RECT 547.650 152.400 549.450 156.000 ;
        RECT 523.950 146.400 528.750 148.500 ;
        RECT 531.450 147.450 538.050 148.500 ;
        RECT 531.450 146.700 533.250 147.450 ;
        RECT 536.250 146.700 538.050 147.450 ;
        RECT 543.150 147.300 547.050 149.400 ;
        RECT 527.550 145.500 528.750 146.400 ;
        RECT 540.450 145.800 542.250 146.400 ;
        RECT 527.550 144.300 535.050 145.500 ;
        RECT 533.250 143.700 535.050 144.300 ;
        RECT 535.950 144.900 542.250 145.800 ;
        RECT 519.150 142.500 520.050 143.400 ;
        RECT 535.950 142.800 536.850 144.900 ;
        RECT 540.450 144.600 542.250 144.900 ;
        RECT 543.150 144.600 545.850 146.400 ;
        RECT 543.150 143.700 544.050 144.600 ;
        RECT 528.450 142.500 536.850 142.800 ;
        RECT 519.150 141.900 536.850 142.500 ;
        RECT 538.950 142.800 544.050 143.700 ;
        RECT 544.950 142.800 547.050 143.700 ;
        RECT 550.650 143.400 552.450 155.400 ;
        RECT 560.700 143.400 562.500 156.000 ;
        RECT 565.800 149.400 567.600 155.400 ;
        RECT 568.800 149.400 570.600 156.000 ;
        RECT 519.150 141.300 530.250 141.900 ;
        RECT 472.950 135.750 477.450 136.050 ;
        RECT 471.150 133.950 477.450 135.750 ;
        RECT 487.950 133.950 490.050 136.050 ;
        RECT 490.950 133.950 493.050 136.050 ;
        RECT 493.950 133.950 496.050 136.050 ;
        RECT 502.950 133.950 505.050 136.050 ;
        RECT 505.950 133.950 508.050 136.050 ;
        RECT 508.950 133.950 511.050 136.050 ;
        RECT 511.950 133.950 514.050 136.050 ;
        RECT 452.850 129.000 464.850 130.200 ;
        RECT 452.850 127.200 453.900 129.000 ;
        RECT 463.050 128.400 464.850 129.000 ;
        RECT 439.500 120.000 441.300 126.600 ;
        RECT 444.150 120.600 445.950 126.600 ;
        RECT 448.950 124.500 451.050 126.600 ;
        RECT 452.550 125.400 454.350 127.200 ;
        RECT 476.250 126.600 477.450 133.950 ;
        RECT 455.850 125.550 457.650 126.300 ;
        RECT 469.950 125.700 472.050 126.600 ;
        RECT 455.850 124.500 460.800 125.550 ;
        RECT 450.000 123.600 451.050 124.500 ;
        RECT 459.750 123.600 460.800 124.500 ;
        RECT 468.300 124.500 472.050 125.700 ;
        RECT 468.300 123.600 469.350 124.500 ;
        RECT 447.150 120.000 448.950 123.600 ;
        RECT 450.000 122.700 453.750 123.600 ;
        RECT 451.950 120.600 453.750 122.700 ;
        RECT 456.450 120.000 458.250 123.600 ;
        RECT 459.750 120.600 461.550 123.600 ;
        RECT 463.350 120.000 465.150 123.600 ;
        RECT 467.550 120.600 469.350 123.600 ;
        RECT 472.350 120.000 474.150 123.600 ;
        RECT 475.650 120.600 477.450 126.600 ;
        RECT 491.400 123.600 492.300 133.950 ;
        RECT 506.100 132.150 507.900 133.950 ;
        RECT 509.850 129.750 511.050 133.950 ;
        RECT 512.100 132.150 513.900 133.950 ;
        RECT 509.850 128.700 513.600 129.750 ;
        RECT 503.400 125.700 511.200 127.050 ;
        RECT 487.800 120.000 489.600 123.600 ;
        RECT 490.800 120.600 492.600 123.600 ;
        RECT 493.800 120.000 495.600 123.600 ;
        RECT 503.400 120.600 505.200 125.700 ;
        RECT 506.400 120.000 508.200 124.800 ;
        RECT 509.400 120.600 511.200 125.700 ;
        RECT 512.400 126.600 513.600 128.700 ;
        RECT 519.150 126.600 520.050 141.300 ;
        RECT 528.450 141.000 530.250 141.300 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 529.950 134.400 532.050 136.050 ;
        RECT 521.100 132.150 522.900 133.950 ;
        RECT 524.100 133.200 532.050 134.400 ;
        RECT 524.100 132.600 525.900 133.200 ;
        RECT 522.000 131.400 522.900 132.150 ;
        RECT 527.100 131.400 528.900 132.000 ;
        RECT 522.000 130.200 528.900 131.400 ;
        RECT 538.950 130.200 539.850 142.800 ;
        RECT 544.950 141.600 549.150 142.800 ;
        RECT 548.250 139.800 550.050 141.600 ;
        RECT 551.250 136.050 552.450 143.400 ;
        RECT 560.100 136.050 561.900 137.850 ;
        RECT 565.950 136.050 567.150 149.400 ;
        RECT 581.400 143.400 583.200 156.000 ;
        RECT 586.500 144.600 588.300 155.400 ;
        RECT 584.700 143.400 588.300 144.600 ;
        RECT 599.700 143.400 601.500 156.000 ;
        RECT 604.800 149.400 606.600 155.400 ;
        RECT 607.800 149.400 609.600 156.000 ;
        RECT 581.100 136.050 582.900 137.850 ;
        RECT 584.700 136.050 585.600 143.400 ;
        RECT 586.950 141.450 589.050 142.050 ;
        RECT 595.950 141.450 598.050 142.050 ;
        RECT 586.950 140.550 598.050 141.450 ;
        RECT 586.950 139.950 589.050 140.550 ;
        RECT 595.950 139.950 598.050 140.550 ;
        RECT 587.100 136.050 588.900 137.850 ;
        RECT 599.100 136.050 600.900 137.850 ;
        RECT 604.950 136.050 606.150 149.400 ;
        RECT 620.400 143.400 622.200 156.000 ;
        RECT 625.500 144.600 627.300 155.400 ;
        RECT 641.400 149.400 643.200 156.000 ;
        RECT 644.400 149.400 646.200 155.400 ;
        RECT 623.700 143.400 627.300 144.600 ;
        RECT 620.100 136.050 621.900 137.850 ;
        RECT 623.700 136.050 624.600 143.400 ;
        RECT 628.950 138.450 631.050 139.050 ;
        RECT 634.950 138.450 637.050 139.050 ;
        RECT 626.100 136.050 627.900 137.850 ;
        RECT 628.950 137.550 637.050 138.450 ;
        RECT 628.950 136.950 631.050 137.550 ;
        RECT 634.950 136.950 637.050 137.550 ;
        RECT 644.850 136.050 646.050 149.400 ;
        RECT 649.500 143.400 651.300 156.000 ;
        RECT 659.700 143.400 661.500 156.000 ;
        RECT 664.800 149.400 666.600 155.400 ;
        RECT 667.800 149.400 669.600 156.000 ;
        RECT 680.400 149.400 682.200 156.000 ;
        RECT 683.400 149.400 685.200 155.400 ;
        RECT 695.400 149.400 697.200 156.000 ;
        RECT 698.400 149.400 700.200 155.400 ;
        RECT 650.100 136.050 651.900 137.850 ;
        RECT 659.100 136.050 660.900 137.850 ;
        RECT 664.950 136.050 666.150 149.400 ;
        RECT 670.950 144.450 673.050 144.900 ;
        RECT 679.950 144.450 682.050 145.050 ;
        RECT 670.950 143.550 682.050 144.450 ;
        RECT 670.950 142.800 673.050 143.550 ;
        RECT 679.950 142.950 682.050 143.550 ;
        RECT 680.100 136.050 681.900 137.850 ;
        RECT 683.400 136.050 684.600 149.400 ;
        RECT 695.100 136.050 696.900 137.850 ;
        RECT 698.400 136.050 699.600 149.400 ;
        RECT 704.550 143.400 706.350 155.400 ;
        RECT 707.550 152.400 709.350 156.000 ;
        RECT 712.050 149.400 713.850 155.400 ;
        RECT 716.250 149.400 718.050 156.000 ;
        RECT 709.950 147.300 713.850 149.400 ;
        RECT 719.850 148.500 721.650 155.400 ;
        RECT 722.850 149.400 724.650 156.000 ;
        RECT 727.650 149.400 729.450 155.400 ;
        RECT 733.050 149.400 734.850 156.000 ;
        RECT 728.250 148.500 729.450 149.400 ;
        RECT 718.950 147.450 725.550 148.500 ;
        RECT 718.950 146.700 720.750 147.450 ;
        RECT 723.750 146.700 725.550 147.450 ;
        RECT 728.250 146.400 733.050 148.500 ;
        RECT 711.150 144.600 713.850 146.400 ;
        RECT 714.750 145.800 716.550 146.400 ;
        RECT 714.750 144.900 721.050 145.800 ;
        RECT 728.250 145.500 729.450 146.400 ;
        RECT 714.750 144.600 716.550 144.900 ;
        RECT 712.950 143.700 713.850 144.600 ;
        RECT 704.550 136.050 705.750 143.400 ;
        RECT 709.950 142.800 712.050 143.700 ;
        RECT 712.950 142.800 718.050 143.700 ;
        RECT 707.850 141.600 712.050 142.800 ;
        RECT 706.950 139.800 708.750 141.600 ;
        RECT 547.950 135.750 552.450 136.050 ;
        RECT 546.150 133.950 552.450 135.750 ;
        RECT 559.950 133.950 562.050 136.050 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 565.950 133.950 568.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 583.950 133.950 586.050 136.050 ;
        RECT 586.950 133.950 589.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 604.950 133.950 607.050 136.050 ;
        RECT 607.950 133.950 610.050 136.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 625.950 133.950 628.050 136.050 ;
        RECT 640.950 133.950 643.050 136.050 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 658.950 133.950 661.050 136.050 ;
        RECT 661.950 133.950 664.050 136.050 ;
        RECT 664.950 133.950 667.050 136.050 ;
        RECT 667.950 133.950 670.050 136.050 ;
        RECT 679.950 133.950 682.050 136.050 ;
        RECT 682.950 133.950 685.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 697.950 133.950 700.050 136.050 ;
        RECT 704.550 135.750 709.050 136.050 ;
        RECT 704.550 133.950 710.850 135.750 ;
        RECT 527.850 129.000 539.850 130.200 ;
        RECT 527.850 127.200 528.900 129.000 ;
        RECT 538.050 128.400 539.850 129.000 ;
        RECT 512.400 120.600 514.200 126.600 ;
        RECT 519.150 120.600 520.950 126.600 ;
        RECT 523.950 124.500 526.050 126.600 ;
        RECT 527.550 125.400 529.350 127.200 ;
        RECT 551.250 126.600 552.450 133.950 ;
        RECT 563.100 132.150 564.900 133.950 ;
        RECT 566.850 129.750 568.050 133.950 ;
        RECT 569.100 132.150 570.900 133.950 ;
        RECT 566.850 128.700 570.600 129.750 ;
        RECT 530.850 125.550 532.650 126.300 ;
        RECT 544.950 125.700 547.050 126.600 ;
        RECT 530.850 124.500 535.800 125.550 ;
        RECT 525.000 123.600 526.050 124.500 ;
        RECT 534.750 123.600 535.800 124.500 ;
        RECT 543.300 124.500 547.050 125.700 ;
        RECT 543.300 123.600 544.350 124.500 ;
        RECT 522.150 120.000 523.950 123.600 ;
        RECT 525.000 122.700 528.750 123.600 ;
        RECT 526.950 120.600 528.750 122.700 ;
        RECT 531.450 120.000 533.250 123.600 ;
        RECT 534.750 120.600 536.550 123.600 ;
        RECT 538.350 120.000 540.150 123.600 ;
        RECT 542.550 120.600 544.350 123.600 ;
        RECT 547.350 120.000 549.150 123.600 ;
        RECT 550.650 120.600 552.450 126.600 ;
        RECT 560.400 125.700 568.200 127.050 ;
        RECT 560.400 120.600 562.200 125.700 ;
        RECT 563.400 120.000 565.200 124.800 ;
        RECT 566.400 120.600 568.200 125.700 ;
        RECT 569.400 126.600 570.600 128.700 ;
        RECT 569.400 120.600 571.200 126.600 ;
        RECT 584.700 123.600 585.600 133.950 ;
        RECT 602.100 132.150 603.900 133.950 ;
        RECT 605.850 129.750 607.050 133.950 ;
        RECT 608.100 132.150 609.900 133.950 ;
        RECT 605.850 128.700 609.600 129.750 ;
        RECT 599.400 125.700 607.200 127.050 ;
        RECT 581.400 120.000 583.200 123.600 ;
        RECT 584.400 120.600 586.200 123.600 ;
        RECT 587.400 120.000 589.200 123.600 ;
        RECT 599.400 120.600 601.200 125.700 ;
        RECT 602.400 120.000 604.200 124.800 ;
        RECT 605.400 120.600 607.200 125.700 ;
        RECT 608.400 126.600 609.600 128.700 ;
        RECT 608.400 120.600 610.200 126.600 ;
        RECT 623.700 123.600 624.600 133.950 ;
        RECT 641.100 132.150 642.900 133.950 ;
        RECT 643.950 129.750 645.150 133.950 ;
        RECT 647.100 132.150 648.900 133.950 ;
        RECT 662.100 132.150 663.900 133.950 ;
        RECT 641.400 128.700 645.150 129.750 ;
        RECT 665.850 129.750 667.050 133.950 ;
        RECT 668.100 132.150 669.900 133.950 ;
        RECT 665.850 128.700 669.600 129.750 ;
        RECT 641.400 126.600 642.600 128.700 ;
        RECT 620.400 120.000 622.200 123.600 ;
        RECT 623.400 120.600 625.200 123.600 ;
        RECT 626.400 120.000 628.200 123.600 ;
        RECT 640.800 120.600 642.600 126.600 ;
        RECT 643.800 125.700 651.600 127.050 ;
        RECT 643.800 120.600 645.600 125.700 ;
        RECT 646.800 120.000 648.600 124.800 ;
        RECT 649.800 120.600 651.600 125.700 ;
        RECT 659.400 125.700 667.200 127.050 ;
        RECT 659.400 120.600 661.200 125.700 ;
        RECT 662.400 120.000 664.200 124.800 ;
        RECT 665.400 120.600 667.200 125.700 ;
        RECT 668.400 126.600 669.600 128.700 ;
        RECT 668.400 120.600 670.200 126.600 ;
        RECT 683.400 123.600 684.600 133.950 ;
        RECT 698.400 123.600 699.600 133.950 ;
        RECT 704.550 126.600 705.750 133.950 ;
        RECT 717.150 130.200 718.050 142.800 ;
        RECT 720.150 142.800 721.050 144.900 ;
        RECT 721.950 144.300 729.450 145.500 ;
        RECT 721.950 143.700 723.750 144.300 ;
        RECT 736.050 143.400 737.850 155.400 ;
        RECT 720.150 142.500 728.550 142.800 ;
        RECT 736.950 142.500 737.850 143.400 ;
        RECT 720.150 141.900 737.850 142.500 ;
        RECT 726.750 141.300 737.850 141.900 ;
        RECT 746.400 149.400 748.200 155.400 ;
        RECT 749.400 149.400 751.200 156.000 ;
        RECT 746.400 142.500 747.600 149.400 ;
        RECT 752.400 143.400 754.200 155.400 ;
        RECT 764.700 143.400 766.500 156.000 ;
        RECT 769.800 149.400 771.600 155.400 ;
        RECT 772.800 149.400 774.600 156.000 ;
        RECT 787.800 149.400 789.600 156.000 ;
        RECT 790.800 149.400 792.600 155.400 ;
        RECT 793.800 149.400 795.600 156.000 ;
        RECT 746.400 141.600 752.100 142.500 ;
        RECT 726.750 141.000 728.550 141.300 ;
        RECT 724.950 134.400 727.050 136.050 ;
        RECT 724.950 133.200 732.900 134.400 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 731.100 132.600 732.900 133.200 ;
        RECT 734.100 132.150 735.900 133.950 ;
        RECT 728.100 131.400 729.900 132.000 ;
        RECT 734.100 131.400 735.000 132.150 ;
        RECT 728.100 130.200 735.000 131.400 ;
        RECT 717.150 129.000 729.150 130.200 ;
        RECT 717.150 128.400 718.950 129.000 ;
        RECT 728.100 127.200 729.150 129.000 ;
        RECT 680.400 120.000 682.200 123.600 ;
        RECT 683.400 120.600 685.200 123.600 ;
        RECT 695.400 120.000 697.200 123.600 ;
        RECT 698.400 120.600 700.200 123.600 ;
        RECT 704.550 120.600 706.350 126.600 ;
        RECT 709.950 125.700 712.050 126.600 ;
        RECT 709.950 124.500 713.700 125.700 ;
        RECT 724.350 125.550 726.150 126.300 ;
        RECT 712.650 123.600 713.700 124.500 ;
        RECT 721.200 124.500 726.150 125.550 ;
        RECT 727.650 125.400 729.450 127.200 ;
        RECT 736.950 126.600 737.850 141.300 ;
        RECT 750.150 140.700 752.100 141.600 ;
        RECT 746.100 136.050 747.900 137.850 ;
        RECT 745.950 133.950 748.050 136.050 ;
        RECT 750.150 129.300 751.050 140.700 ;
        RECT 753.000 136.050 754.200 143.400 ;
        RECT 764.100 136.050 765.900 137.850 ;
        RECT 769.950 136.050 771.150 149.400 ;
        RECT 751.950 133.950 754.200 136.050 ;
        RECT 763.950 133.950 766.050 136.050 ;
        RECT 766.950 133.950 769.050 136.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 791.400 135.900 792.600 149.400 ;
        RECT 803.700 143.400 805.500 156.000 ;
        RECT 808.800 149.400 810.600 155.400 ;
        RECT 811.800 149.400 813.600 156.000 ;
        RECT 803.100 136.050 804.900 137.850 ;
        RECT 808.950 136.050 810.150 149.400 ;
        RECT 818.550 143.400 820.350 155.400 ;
        RECT 821.550 152.400 823.350 156.000 ;
        RECT 826.050 149.400 827.850 155.400 ;
        RECT 830.250 149.400 832.050 156.000 ;
        RECT 823.950 147.300 827.850 149.400 ;
        RECT 833.850 148.500 835.650 155.400 ;
        RECT 836.850 149.400 838.650 156.000 ;
        RECT 841.650 149.400 843.450 155.400 ;
        RECT 847.050 149.400 848.850 156.000 ;
        RECT 842.250 148.500 843.450 149.400 ;
        RECT 832.950 147.450 839.550 148.500 ;
        RECT 832.950 146.700 834.750 147.450 ;
        RECT 837.750 146.700 839.550 147.450 ;
        RECT 842.250 146.400 847.050 148.500 ;
        RECT 825.150 144.600 827.850 146.400 ;
        RECT 828.750 145.800 830.550 146.400 ;
        RECT 828.750 144.900 835.050 145.800 ;
        RECT 842.250 145.500 843.450 146.400 ;
        RECT 828.750 144.600 830.550 144.900 ;
        RECT 826.950 143.700 827.850 144.600 ;
        RECT 818.550 136.050 819.750 143.400 ;
        RECT 823.950 142.800 826.050 143.700 ;
        RECT 826.950 142.800 832.050 143.700 ;
        RECT 821.850 141.600 826.050 142.800 ;
        RECT 820.950 139.800 822.750 141.600 ;
        RECT 750.150 128.400 752.100 129.300 ;
        RECT 730.950 124.500 733.050 126.600 ;
        RECT 721.200 123.600 722.250 124.500 ;
        RECT 730.950 123.600 732.000 124.500 ;
        RECT 707.850 120.000 709.650 123.600 ;
        RECT 712.650 120.600 714.450 123.600 ;
        RECT 716.850 120.000 718.650 123.600 ;
        RECT 720.450 120.600 722.250 123.600 ;
        RECT 723.750 120.000 725.550 123.600 ;
        RECT 728.250 122.700 732.000 123.600 ;
        RECT 728.250 120.600 730.050 122.700 ;
        RECT 733.050 120.000 734.850 123.600 ;
        RECT 736.050 120.600 737.850 126.600 ;
        RECT 746.400 127.500 752.100 128.400 ;
        RECT 746.400 123.600 747.600 127.500 ;
        RECT 753.000 126.600 754.200 133.950 ;
        RECT 767.100 132.150 768.900 133.950 ;
        RECT 770.850 129.750 772.050 133.950 ;
        RECT 773.100 132.150 774.900 133.950 ;
        RECT 787.950 133.800 790.050 135.900 ;
        RECT 790.950 133.800 793.050 135.900 ;
        RECT 793.950 133.800 796.050 135.900 ;
        RECT 802.950 133.950 805.050 136.050 ;
        RECT 805.950 133.950 808.050 136.050 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 818.550 135.750 823.050 136.050 ;
        RECT 818.550 133.950 824.850 135.750 ;
        RECT 788.100 132.000 789.900 133.800 ;
        RECT 770.850 128.700 774.600 129.750 ;
        RECT 791.400 128.700 792.600 133.800 ;
        RECT 794.100 132.000 795.900 133.800 ;
        RECT 806.100 132.150 807.900 133.950 ;
        RECT 809.850 129.750 811.050 133.950 ;
        RECT 812.100 132.150 813.900 133.950 ;
        RECT 809.850 128.700 813.600 129.750 ;
        RECT 746.400 120.600 748.200 123.600 ;
        RECT 749.400 120.000 751.200 123.600 ;
        RECT 752.400 120.600 754.200 126.600 ;
        RECT 764.400 125.700 772.200 127.050 ;
        RECT 764.400 120.600 766.200 125.700 ;
        RECT 767.400 120.000 769.200 124.800 ;
        RECT 770.400 120.600 772.200 125.700 ;
        RECT 773.400 126.600 774.600 128.700 ;
        RECT 788.400 127.800 792.600 128.700 ;
        RECT 773.400 120.600 775.200 126.600 ;
        RECT 788.400 120.600 790.200 127.800 ;
        RECT 793.500 120.000 795.300 126.600 ;
        RECT 803.400 125.700 811.200 127.050 ;
        RECT 803.400 120.600 805.200 125.700 ;
        RECT 806.400 120.000 808.200 124.800 ;
        RECT 809.400 120.600 811.200 125.700 ;
        RECT 812.400 126.600 813.600 128.700 ;
        RECT 818.550 126.600 819.750 133.950 ;
        RECT 831.150 130.200 832.050 142.800 ;
        RECT 834.150 142.800 835.050 144.900 ;
        RECT 835.950 144.300 843.450 145.500 ;
        RECT 835.950 143.700 837.750 144.300 ;
        RECT 850.050 143.400 851.850 155.400 ;
        RECT 834.150 142.500 842.550 142.800 ;
        RECT 850.950 142.500 851.850 143.400 ;
        RECT 834.150 141.900 851.850 142.500 ;
        RECT 840.750 141.300 851.850 141.900 ;
        RECT 840.750 141.000 842.550 141.300 ;
        RECT 838.950 134.400 841.050 136.050 ;
        RECT 838.950 133.200 846.900 134.400 ;
        RECT 847.950 133.950 850.050 136.050 ;
        RECT 845.100 132.600 846.900 133.200 ;
        RECT 848.100 132.150 849.900 133.950 ;
        RECT 842.100 131.400 843.900 132.000 ;
        RECT 848.100 131.400 849.000 132.150 ;
        RECT 842.100 130.200 849.000 131.400 ;
        RECT 831.150 129.000 843.150 130.200 ;
        RECT 831.150 128.400 832.950 129.000 ;
        RECT 842.100 127.200 843.150 129.000 ;
        RECT 812.400 120.600 814.200 126.600 ;
        RECT 818.550 120.600 820.350 126.600 ;
        RECT 823.950 125.700 826.050 126.600 ;
        RECT 823.950 124.500 827.700 125.700 ;
        RECT 838.350 125.550 840.150 126.300 ;
        RECT 826.650 123.600 827.700 124.500 ;
        RECT 835.200 124.500 840.150 125.550 ;
        RECT 841.650 125.400 843.450 127.200 ;
        RECT 850.950 126.600 851.850 141.300 ;
        RECT 844.950 124.500 847.050 126.600 ;
        RECT 835.200 123.600 836.250 124.500 ;
        RECT 844.950 123.600 846.000 124.500 ;
        RECT 821.850 120.000 823.650 123.600 ;
        RECT 826.650 120.600 828.450 123.600 ;
        RECT 830.850 120.000 832.650 123.600 ;
        RECT 834.450 120.600 836.250 123.600 ;
        RECT 837.750 120.000 839.550 123.600 ;
        RECT 842.250 122.700 846.000 123.600 ;
        RECT 842.250 120.600 844.050 122.700 ;
        RECT 847.050 120.000 848.850 123.600 ;
        RECT 850.050 120.600 851.850 126.600 ;
        RECT 10.800 110.400 12.600 116.400 ;
        RECT 18.300 110.400 20.100 116.400 ;
        RECT 25.800 110.400 27.600 116.400 ;
        RECT 35.400 113.400 37.200 117.000 ;
        RECT 38.400 113.400 40.200 116.400 ;
        RECT 52.800 113.400 54.600 117.000 ;
        RECT 55.800 113.400 57.600 116.400 ;
        RECT 58.800 113.400 60.600 117.000 ;
        RECT 71.700 113.400 73.500 117.000 ;
        RECT 10.800 109.500 15.600 110.400 ;
        RECT 13.500 108.300 15.600 109.500 ;
        RECT 18.600 108.900 19.800 110.400 ;
        RECT 16.950 106.800 19.800 108.900 ;
        RECT 25.800 108.600 27.000 110.400 ;
        RECT 15.750 103.800 17.850 105.900 ;
        RECT 1.950 102.450 4.050 103.050 ;
        RECT 10.950 102.450 13.050 103.200 ;
        RECT 1.950 101.550 13.050 102.450 ;
        RECT 15.600 102.000 17.400 103.800 ;
        RECT 1.950 100.950 4.050 101.550 ;
        RECT 10.950 101.100 13.050 101.550 ;
        RECT 18.750 101.100 19.800 106.800 ;
        RECT 20.700 107.700 27.000 108.600 ;
        RECT 20.700 105.600 22.800 107.700 ;
        RECT 20.700 103.800 22.500 105.600 ;
        RECT 25.950 103.200 27.750 105.000 ;
        RECT 25.950 102.300 28.050 103.200 ;
        RECT 38.400 103.050 39.600 113.400 ;
        RECT 56.400 103.050 57.300 113.400 ;
        RECT 74.700 111.600 76.500 116.400 ;
        RECT 71.400 110.400 76.500 111.600 ;
        RECT 79.200 110.400 81.000 117.000 ;
        RECT 91.800 110.400 93.600 116.400 ;
        RECT 99.600 111.000 101.400 116.400 ;
        RECT 71.400 103.200 72.300 110.400 ;
        RECT 91.800 109.500 96.300 110.400 ;
        RECT 94.200 107.100 96.300 109.500 ;
        RECT 99.750 108.900 100.650 111.000 ;
        RECT 106.800 110.400 108.600 116.400 ;
        RECT 116.700 110.400 118.500 117.000 ;
        RECT 107.100 109.500 108.600 110.400 ;
        RECT 97.650 106.800 100.650 108.900 ;
        RECT 104.250 108.000 108.600 109.500 ;
        RECT 121.800 109.200 123.600 116.400 ;
        RECT 134.700 110.400 136.500 117.000 ;
        RECT 139.800 109.200 141.600 116.400 ;
        RECT 119.400 108.300 123.600 109.200 ;
        RECT 137.400 108.300 141.600 109.200 ;
        RECT 147.150 110.400 148.950 116.400 ;
        RECT 150.150 113.400 151.950 117.000 ;
        RECT 154.950 114.300 156.750 116.400 ;
        RECT 153.000 113.400 156.750 114.300 ;
        RECT 159.450 113.400 161.250 117.000 ;
        RECT 162.750 113.400 164.550 116.400 ;
        RECT 166.350 113.400 168.150 117.000 ;
        RECT 170.550 113.400 172.350 116.400 ;
        RECT 175.350 113.400 177.150 117.000 ;
        RECT 153.000 112.500 154.050 113.400 ;
        RECT 162.750 112.500 163.800 113.400 ;
        RECT 151.950 110.400 154.050 112.500 ;
        RECT 74.100 103.200 75.900 105.000 ;
        RECT 80.100 103.200 81.900 105.000 ;
        RECT 11.100 99.300 12.900 101.100 ;
        RECT 17.400 100.200 19.800 101.100 ;
        RECT 20.700 101.100 28.050 102.300 ;
        RECT 20.700 100.500 22.500 101.100 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 52.950 100.950 55.050 103.050 ;
        RECT 55.950 100.950 58.050 103.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 70.950 101.100 73.050 103.200 ;
        RECT 73.950 101.100 76.050 103.200 ;
        RECT 76.950 101.100 79.050 103.200 ;
        RECT 79.950 101.100 82.050 103.200 ;
        RECT 91.950 101.100 94.050 103.200 ;
        RECT 96.750 102.900 98.850 105.000 ;
        RECT 96.900 101.100 98.700 102.900 ;
        RECT 16.950 98.100 19.050 100.200 ;
        RECT 18.000 96.000 18.900 98.100 ;
        RECT 19.950 97.500 23.700 99.300 ;
        RECT 35.100 99.150 36.900 100.950 ;
        RECT 19.950 97.200 22.050 97.500 ;
        RECT 18.000 95.100 19.500 96.000 ;
        RECT 13.500 93.600 15.600 94.500 ;
        RECT 10.800 92.400 15.600 93.600 ;
        RECT 18.300 93.600 19.500 95.100 ;
        RECT 23.100 93.600 25.200 95.700 ;
        RECT 10.800 81.600 12.600 92.400 ;
        RECT 18.300 81.600 20.100 93.600 ;
        RECT 23.100 92.700 27.600 93.600 ;
        RECT 25.800 81.600 27.600 92.700 ;
        RECT 38.400 87.600 39.600 100.950 ;
        RECT 53.100 99.150 54.900 100.950 ;
        RECT 56.400 93.600 57.300 100.950 ;
        RECT 59.100 99.150 60.900 100.950 ;
        RECT 58.950 96.450 61.050 97.050 ;
        RECT 67.950 96.450 70.050 97.050 ;
        RECT 58.950 95.550 70.050 96.450 ;
        RECT 58.950 94.950 61.050 95.550 ;
        RECT 67.950 94.950 70.050 95.550 ;
        RECT 71.400 93.600 72.300 101.100 ;
        RECT 77.100 99.300 78.900 101.100 ;
        RECT 85.950 99.450 88.050 100.050 ;
        RECT 92.100 99.450 93.900 101.100 ;
        RECT 99.750 100.200 100.650 106.800 ;
        RECT 101.550 105.900 103.350 107.700 ;
        RECT 104.250 107.400 106.350 108.000 ;
        RECT 101.700 105.000 103.800 105.900 ;
        RECT 101.700 103.800 108.750 105.000 ;
        RECT 106.950 103.200 108.750 103.800 ;
        RECT 116.100 103.200 117.900 105.000 ;
        RECT 119.400 103.200 120.600 108.300 ;
        RECT 122.100 103.200 123.900 105.000 ;
        RECT 134.100 103.200 135.900 105.000 ;
        RECT 137.400 103.200 138.600 108.300 ;
        RECT 140.100 103.200 141.900 105.000 ;
        RECT 101.700 100.800 103.800 102.900 ;
        RECT 106.950 101.100 109.050 103.200 ;
        RECT 115.950 101.100 118.050 103.200 ;
        RECT 118.950 101.100 121.050 103.200 ;
        RECT 121.950 101.100 124.050 103.200 ;
        RECT 133.950 101.100 136.050 103.200 ;
        RECT 136.950 101.100 139.050 103.200 ;
        RECT 139.950 101.100 142.050 103.200 ;
        RECT 85.950 99.300 93.900 99.450 ;
        RECT 85.950 98.550 93.450 99.300 ;
        RECT 97.650 98.700 100.650 100.200 ;
        RECT 102.000 99.000 103.800 100.800 ;
        RECT 85.950 97.950 88.050 98.550 ;
        RECT 97.650 98.100 99.750 98.700 ;
        RECT 94.800 93.600 96.900 94.500 ;
        RECT 53.700 92.400 57.300 93.600 ;
        RECT 35.400 81.000 37.200 87.600 ;
        RECT 38.400 81.600 40.200 87.600 ;
        RECT 53.700 81.600 55.500 92.400 ;
        RECT 58.800 81.000 60.600 93.600 ;
        RECT 70.800 81.600 72.600 93.600 ;
        RECT 73.800 92.700 81.600 93.600 ;
        RECT 73.800 81.600 75.600 92.700 ;
        RECT 76.800 81.000 78.600 91.800 ;
        RECT 79.800 81.600 81.600 92.700 ;
        RECT 91.800 92.400 96.900 93.600 ;
        RECT 97.800 93.600 99.000 98.100 ;
        RECT 100.650 95.700 102.450 97.800 ;
        RECT 100.650 94.800 105.900 95.700 ;
        RECT 103.800 93.900 105.900 94.800 ;
        RECT 97.800 92.700 101.100 93.600 ;
        RECT 103.800 92.700 108.600 93.900 ;
        RECT 91.800 81.600 93.600 92.400 ;
        RECT 99.300 81.600 101.100 92.700 ;
        RECT 106.800 81.600 108.600 92.700 ;
        RECT 119.400 87.600 120.600 101.100 ;
        RECT 137.400 87.600 138.600 101.100 ;
        RECT 147.150 95.700 148.050 110.400 ;
        RECT 155.550 109.800 157.350 111.600 ;
        RECT 158.850 111.450 163.800 112.500 ;
        RECT 171.300 112.500 172.350 113.400 ;
        RECT 158.850 110.700 160.650 111.450 ;
        RECT 171.300 111.300 175.050 112.500 ;
        RECT 172.950 110.400 175.050 111.300 ;
        RECT 178.650 110.400 180.450 116.400 ;
        RECT 155.850 108.000 156.900 109.800 ;
        RECT 166.050 108.000 167.850 108.600 ;
        RECT 155.850 106.800 167.850 108.000 ;
        RECT 150.000 105.600 156.900 106.800 ;
        RECT 150.000 104.850 150.900 105.600 ;
        RECT 155.100 105.000 156.900 105.600 ;
        RECT 149.100 103.050 150.900 104.850 ;
        RECT 152.100 103.800 153.900 104.400 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 152.100 102.600 160.050 103.800 ;
        RECT 157.950 100.950 160.050 102.600 ;
        RECT 156.450 95.700 158.250 96.000 ;
        RECT 147.150 95.100 158.250 95.700 ;
        RECT 147.150 94.500 164.850 95.100 ;
        RECT 147.150 93.600 148.050 94.500 ;
        RECT 156.450 94.200 164.850 94.500 ;
        RECT 116.400 81.000 118.200 87.600 ;
        RECT 119.400 81.600 121.200 87.600 ;
        RECT 122.400 81.000 124.200 87.600 ;
        RECT 134.400 81.000 136.200 87.600 ;
        RECT 137.400 81.600 139.200 87.600 ;
        RECT 140.400 81.000 142.200 87.600 ;
        RECT 147.150 81.600 148.950 93.600 ;
        RECT 161.250 92.700 163.050 93.300 ;
        RECT 155.550 91.500 163.050 92.700 ;
        RECT 163.950 92.100 164.850 94.200 ;
        RECT 166.950 94.200 167.850 106.800 ;
        RECT 179.250 103.050 180.450 110.400 ;
        RECT 188.400 111.300 190.200 116.400 ;
        RECT 191.400 112.200 193.200 117.000 ;
        RECT 194.400 111.300 196.200 116.400 ;
        RECT 188.400 109.950 196.200 111.300 ;
        RECT 197.400 110.400 199.200 116.400 ;
        RECT 209.700 110.400 211.500 117.000 ;
        RECT 197.400 108.300 198.600 110.400 ;
        RECT 214.800 109.200 216.600 116.400 ;
        RECT 194.850 107.250 198.600 108.300 ;
        RECT 212.400 108.300 216.600 109.200 ;
        RECT 221.550 110.400 223.350 116.400 ;
        RECT 224.850 113.400 226.650 117.000 ;
        RECT 229.650 113.400 231.450 116.400 ;
        RECT 233.850 113.400 235.650 117.000 ;
        RECT 237.450 113.400 239.250 116.400 ;
        RECT 240.750 113.400 242.550 117.000 ;
        RECT 245.250 114.300 247.050 116.400 ;
        RECT 245.250 113.400 249.000 114.300 ;
        RECT 250.050 113.400 251.850 117.000 ;
        RECT 229.650 112.500 230.700 113.400 ;
        RECT 226.950 111.300 230.700 112.500 ;
        RECT 238.200 112.500 239.250 113.400 ;
        RECT 247.950 112.500 249.000 113.400 ;
        RECT 238.200 111.450 243.150 112.500 ;
        RECT 226.950 110.400 229.050 111.300 ;
        RECT 241.350 110.700 243.150 111.450 ;
        RECT 191.100 103.050 192.900 104.850 ;
        RECT 194.850 103.050 196.050 107.250 ;
        RECT 197.100 103.050 198.900 104.850 ;
        RECT 209.100 103.200 210.900 105.000 ;
        RECT 212.400 103.200 213.600 108.300 ;
        RECT 215.100 103.200 216.900 105.000 ;
        RECT 174.150 101.250 180.450 103.050 ;
        RECT 175.950 100.950 180.450 101.250 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 193.950 100.950 196.050 103.050 ;
        RECT 196.950 100.950 199.050 103.050 ;
        RECT 208.950 101.100 211.050 103.200 ;
        RECT 211.950 101.100 214.050 103.200 ;
        RECT 214.950 101.100 217.050 103.200 ;
        RECT 221.550 103.050 222.750 110.400 ;
        RECT 244.650 109.800 246.450 111.600 ;
        RECT 247.950 110.400 250.050 112.500 ;
        RECT 253.050 110.400 254.850 116.400 ;
        RECT 234.150 108.000 235.950 108.600 ;
        RECT 245.100 108.000 246.150 109.800 ;
        RECT 234.150 106.800 246.150 108.000 ;
        RECT 221.550 101.250 227.850 103.050 ;
        RECT 176.250 95.400 178.050 97.200 ;
        RECT 172.950 94.200 177.150 95.400 ;
        RECT 166.950 93.300 172.050 94.200 ;
        RECT 172.950 93.300 175.050 94.200 ;
        RECT 179.250 93.600 180.450 100.950 ;
        RECT 188.100 99.150 189.900 100.950 ;
        RECT 171.150 92.400 172.050 93.300 ;
        RECT 168.450 92.100 170.250 92.400 ;
        RECT 155.550 90.600 156.750 91.500 ;
        RECT 163.950 91.200 170.250 92.100 ;
        RECT 168.450 90.600 170.250 91.200 ;
        RECT 171.150 90.600 173.850 92.400 ;
        RECT 151.950 88.500 156.750 90.600 ;
        RECT 159.450 89.550 161.250 90.300 ;
        RECT 164.250 89.550 166.050 90.300 ;
        RECT 159.450 88.500 166.050 89.550 ;
        RECT 155.550 87.600 156.750 88.500 ;
        RECT 150.150 81.000 151.950 87.600 ;
        RECT 155.550 81.600 157.350 87.600 ;
        RECT 160.350 81.000 162.150 87.600 ;
        RECT 163.350 81.600 165.150 88.500 ;
        RECT 171.150 87.600 175.050 89.700 ;
        RECT 166.950 81.000 168.750 87.600 ;
        RECT 171.150 81.600 172.950 87.600 ;
        RECT 175.650 81.000 177.450 84.600 ;
        RECT 178.650 81.600 180.450 93.600 ;
        RECT 188.700 81.000 190.500 93.600 ;
        RECT 193.950 87.600 195.150 100.950 ;
        RECT 212.400 87.600 213.600 101.100 ;
        RECT 221.550 100.950 226.050 101.250 ;
        RECT 221.550 93.600 222.750 100.950 ;
        RECT 223.950 95.400 225.750 97.200 ;
        RECT 224.850 94.200 229.050 95.400 ;
        RECT 234.150 94.200 235.050 106.800 ;
        RECT 245.100 105.600 252.000 106.800 ;
        RECT 245.100 105.000 246.900 105.600 ;
        RECT 251.100 104.850 252.000 105.600 ;
        RECT 248.100 103.800 249.900 104.400 ;
        RECT 241.950 102.600 249.900 103.800 ;
        RECT 251.100 103.050 252.900 104.850 ;
        RECT 241.950 100.950 244.050 102.600 ;
        RECT 250.950 100.950 253.050 103.050 ;
        RECT 243.750 95.700 245.550 96.000 ;
        RECT 253.950 95.700 254.850 110.400 ;
        RECT 263.400 113.400 265.200 116.400 ;
        RECT 266.400 113.400 268.200 117.000 ;
        RECT 263.400 109.500 264.600 113.400 ;
        RECT 269.400 110.400 271.200 116.400 ;
        RECT 281.700 110.400 283.500 117.000 ;
        RECT 263.400 108.600 269.100 109.500 ;
        RECT 267.150 107.700 269.100 108.600 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 263.100 99.150 264.900 100.950 ;
        RECT 243.750 95.100 254.850 95.700 ;
        RECT 267.150 96.300 268.050 107.700 ;
        RECT 270.000 103.050 271.200 110.400 ;
        RECT 286.800 109.200 288.600 116.400 ;
        RECT 284.400 108.300 288.600 109.200 ;
        RECT 293.550 110.400 295.350 116.400 ;
        RECT 296.850 113.400 298.650 117.000 ;
        RECT 301.650 113.400 303.450 116.400 ;
        RECT 305.850 113.400 307.650 117.000 ;
        RECT 309.450 113.400 311.250 116.400 ;
        RECT 312.750 113.400 314.550 117.000 ;
        RECT 317.250 114.300 319.050 116.400 ;
        RECT 317.250 113.400 321.000 114.300 ;
        RECT 322.050 113.400 323.850 117.000 ;
        RECT 301.650 112.500 302.700 113.400 ;
        RECT 298.950 111.300 302.700 112.500 ;
        RECT 310.200 112.500 311.250 113.400 ;
        RECT 319.950 112.500 321.000 113.400 ;
        RECT 310.200 111.450 315.150 112.500 ;
        RECT 298.950 110.400 301.050 111.300 ;
        RECT 313.350 110.700 315.150 111.450 ;
        RECT 281.100 103.200 282.900 105.000 ;
        RECT 284.400 103.200 285.600 108.300 ;
        RECT 287.100 103.200 288.900 105.000 ;
        RECT 268.950 100.950 271.200 103.050 ;
        RECT 280.950 101.100 283.050 103.200 ;
        RECT 283.950 101.100 286.050 103.200 ;
        RECT 286.950 101.100 289.050 103.200 ;
        RECT 293.550 103.050 294.750 110.400 ;
        RECT 316.650 109.800 318.450 111.600 ;
        RECT 319.950 110.400 322.050 112.500 ;
        RECT 325.050 110.400 326.850 116.400 ;
        RECT 306.150 108.000 307.950 108.600 ;
        RECT 317.100 108.000 318.150 109.800 ;
        RECT 306.150 106.800 318.150 108.000 ;
        RECT 293.550 101.250 299.850 103.050 ;
        RECT 267.150 95.400 269.100 96.300 ;
        RECT 193.800 81.600 195.600 87.600 ;
        RECT 196.800 81.000 198.600 87.600 ;
        RECT 209.400 81.000 211.200 87.600 ;
        RECT 212.400 81.600 214.200 87.600 ;
        RECT 215.400 81.000 217.200 87.600 ;
        RECT 221.550 81.600 223.350 93.600 ;
        RECT 226.950 93.300 229.050 94.200 ;
        RECT 229.950 93.300 235.050 94.200 ;
        RECT 237.150 94.500 254.850 95.100 ;
        RECT 237.150 94.200 245.550 94.500 ;
        RECT 229.950 92.400 230.850 93.300 ;
        RECT 228.150 90.600 230.850 92.400 ;
        RECT 231.750 92.100 233.550 92.400 ;
        RECT 237.150 92.100 238.050 94.200 ;
        RECT 253.950 93.600 254.850 94.500 ;
        RECT 231.750 91.200 238.050 92.100 ;
        RECT 238.950 92.700 240.750 93.300 ;
        RECT 238.950 91.500 246.450 92.700 ;
        RECT 231.750 90.600 233.550 91.200 ;
        RECT 245.250 90.600 246.450 91.500 ;
        RECT 226.950 87.600 230.850 89.700 ;
        RECT 235.950 89.550 237.750 90.300 ;
        RECT 240.750 89.550 242.550 90.300 ;
        RECT 235.950 88.500 242.550 89.550 ;
        RECT 245.250 88.500 250.050 90.600 ;
        RECT 224.550 81.000 226.350 84.600 ;
        RECT 229.050 81.600 230.850 87.600 ;
        RECT 233.250 81.000 235.050 87.600 ;
        RECT 236.850 81.600 238.650 88.500 ;
        RECT 245.250 87.600 246.450 88.500 ;
        RECT 239.850 81.000 241.650 87.600 ;
        RECT 244.650 81.600 246.450 87.600 ;
        RECT 250.050 81.000 251.850 87.600 ;
        RECT 253.050 81.600 254.850 93.600 ;
        RECT 263.400 94.500 269.100 95.400 ;
        RECT 263.400 87.600 264.600 94.500 ;
        RECT 270.000 93.600 271.200 100.950 ;
        RECT 263.400 81.600 265.200 87.600 ;
        RECT 266.400 81.000 268.200 87.600 ;
        RECT 269.400 81.600 271.200 93.600 ;
        RECT 284.400 87.600 285.600 101.100 ;
        RECT 293.550 100.950 298.050 101.250 ;
        RECT 293.550 93.600 294.750 100.950 ;
        RECT 295.950 95.400 297.750 97.200 ;
        RECT 296.850 94.200 301.050 95.400 ;
        RECT 306.150 94.200 307.050 106.800 ;
        RECT 317.100 105.600 324.000 106.800 ;
        RECT 317.100 105.000 318.900 105.600 ;
        RECT 323.100 104.850 324.000 105.600 ;
        RECT 320.100 103.800 321.900 104.400 ;
        RECT 313.950 102.600 321.900 103.800 ;
        RECT 323.100 103.050 324.900 104.850 ;
        RECT 313.950 100.950 316.050 102.600 ;
        RECT 322.950 100.950 325.050 103.050 ;
        RECT 315.750 95.700 317.550 96.000 ;
        RECT 325.950 95.700 326.850 110.400 ;
        RECT 335.400 111.300 337.200 116.400 ;
        RECT 338.400 112.200 340.200 117.000 ;
        RECT 341.400 111.300 343.200 116.400 ;
        RECT 335.400 109.950 343.200 111.300 ;
        RECT 344.400 110.400 346.200 116.400 ;
        RECT 358.800 110.400 360.600 116.400 ;
        RECT 344.400 108.300 345.600 110.400 ;
        RECT 341.850 107.250 345.600 108.300 ;
        RECT 359.400 108.300 360.600 110.400 ;
        RECT 361.800 111.300 363.600 116.400 ;
        RECT 364.800 112.200 366.600 117.000 ;
        RECT 367.800 111.300 369.600 116.400 ;
        RECT 379.800 113.400 381.600 116.400 ;
        RECT 382.800 113.400 384.600 117.000 ;
        RECT 361.800 109.950 369.600 111.300 ;
        RECT 359.400 107.250 363.150 108.300 ;
        RECT 338.100 103.050 339.900 104.850 ;
        RECT 341.850 103.050 343.050 107.250 ;
        RECT 355.950 105.450 358.050 106.050 ;
        RECT 344.100 103.050 345.900 104.850 ;
        RECT 350.550 104.550 358.050 105.450 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 340.950 100.950 343.050 103.050 ;
        RECT 343.950 100.950 346.050 103.050 ;
        RECT 335.100 99.150 336.900 100.950 ;
        RECT 315.750 95.100 326.850 95.700 ;
        RECT 281.400 81.000 283.200 87.600 ;
        RECT 284.400 81.600 286.200 87.600 ;
        RECT 287.400 81.000 289.200 87.600 ;
        RECT 293.550 81.600 295.350 93.600 ;
        RECT 298.950 93.300 301.050 94.200 ;
        RECT 301.950 93.300 307.050 94.200 ;
        RECT 309.150 94.500 326.850 95.100 ;
        RECT 309.150 94.200 317.550 94.500 ;
        RECT 301.950 92.400 302.850 93.300 ;
        RECT 300.150 90.600 302.850 92.400 ;
        RECT 303.750 92.100 305.550 92.400 ;
        RECT 309.150 92.100 310.050 94.200 ;
        RECT 325.950 93.600 326.850 94.500 ;
        RECT 303.750 91.200 310.050 92.100 ;
        RECT 310.950 92.700 312.750 93.300 ;
        RECT 310.950 91.500 318.450 92.700 ;
        RECT 303.750 90.600 305.550 91.200 ;
        RECT 317.250 90.600 318.450 91.500 ;
        RECT 298.950 87.600 302.850 89.700 ;
        RECT 307.950 89.550 309.750 90.300 ;
        RECT 312.750 89.550 314.550 90.300 ;
        RECT 307.950 88.500 314.550 89.550 ;
        RECT 317.250 88.500 322.050 90.600 ;
        RECT 296.550 81.000 298.350 84.600 ;
        RECT 301.050 81.600 302.850 87.600 ;
        RECT 305.250 81.000 307.050 87.600 ;
        RECT 308.850 81.600 310.650 88.500 ;
        RECT 317.250 87.600 318.450 88.500 ;
        RECT 311.850 81.000 313.650 87.600 ;
        RECT 316.650 81.600 318.450 87.600 ;
        RECT 322.050 81.000 323.850 87.600 ;
        RECT 325.050 81.600 326.850 93.600 ;
        RECT 335.700 81.000 337.500 93.600 ;
        RECT 340.950 87.600 342.150 100.950 ;
        RECT 350.550 100.050 351.450 104.550 ;
        RECT 355.950 103.950 358.050 104.550 ;
        RECT 359.100 103.050 360.900 104.850 ;
        RECT 361.950 103.050 363.150 107.250 ;
        RECT 365.100 103.050 366.900 104.850 ;
        RECT 380.400 103.050 381.600 113.400 ;
        RECT 392.700 110.400 394.500 117.000 ;
        RECT 397.200 110.400 399.000 116.400 ;
        RECT 401.700 110.400 403.500 117.000 ;
        RECT 418.800 110.400 420.600 116.400 ;
        RECT 421.800 110.400 423.600 117.000 ;
        RECT 431.400 111.300 433.200 116.400 ;
        RECT 434.400 112.200 436.200 117.000 ;
        RECT 437.400 111.300 439.200 116.400 ;
        RECT 392.100 103.200 393.900 105.000 ;
        RECT 397.950 103.200 399.000 110.400 ;
        RECT 403.950 108.450 406.050 109.050 ;
        RECT 403.950 107.550 411.450 108.450 ;
        RECT 403.950 106.950 406.050 107.550 ;
        RECT 404.100 103.200 405.900 105.000 ;
        RECT 358.950 100.950 361.050 103.050 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 379.950 100.950 382.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 391.950 101.100 394.050 103.200 ;
        RECT 394.950 101.100 397.050 103.200 ;
        RECT 397.950 101.100 400.050 103.200 ;
        RECT 400.950 101.100 403.050 103.200 ;
        RECT 403.950 101.100 406.050 103.200 ;
        RECT 346.950 98.550 351.450 100.050 ;
        RECT 346.950 97.950 351.000 98.550 ;
        RECT 362.850 87.600 364.050 100.950 ;
        RECT 368.100 99.150 369.900 100.950 ;
        RECT 340.800 81.600 342.600 87.600 ;
        RECT 343.800 81.000 345.600 87.600 ;
        RECT 359.400 81.000 361.200 87.600 ;
        RECT 362.400 81.600 364.200 87.600 ;
        RECT 367.500 81.000 369.300 93.600 ;
        RECT 380.400 87.600 381.600 100.950 ;
        RECT 383.100 99.150 384.900 100.950 ;
        RECT 395.100 99.300 396.900 101.100 ;
        RECT 398.100 95.400 399.000 101.100 ;
        RECT 401.100 99.300 402.900 101.100 ;
        RECT 403.950 99.450 406.050 100.050 ;
        RECT 410.550 99.450 411.450 107.550 ;
        RECT 419.400 103.200 420.600 110.400 ;
        RECT 431.400 109.950 439.200 111.300 ;
        RECT 440.400 110.400 442.200 116.400 ;
        RECT 454.800 113.400 456.600 117.000 ;
        RECT 457.800 113.400 459.600 116.400 ;
        RECT 460.800 113.400 462.600 117.000 ;
        RECT 440.400 108.300 441.600 110.400 ;
        RECT 437.850 107.250 441.600 108.300 ;
        RECT 422.100 103.200 423.900 105.000 ;
        RECT 418.950 101.100 421.050 103.200 ;
        RECT 421.950 101.100 424.050 103.200 ;
        RECT 434.100 103.050 435.900 104.850 ;
        RECT 437.850 103.050 439.050 107.250 ;
        RECT 440.100 103.050 441.900 104.850 ;
        RECT 458.400 103.050 459.300 113.400 ;
        RECT 465.150 110.400 466.950 116.400 ;
        RECT 468.150 113.400 469.950 117.000 ;
        RECT 472.950 114.300 474.750 116.400 ;
        RECT 471.000 113.400 474.750 114.300 ;
        RECT 477.450 113.400 479.250 117.000 ;
        RECT 480.750 113.400 482.550 116.400 ;
        RECT 484.350 113.400 486.150 117.000 ;
        RECT 488.550 113.400 490.350 116.400 ;
        RECT 493.350 113.400 495.150 117.000 ;
        RECT 471.000 112.500 472.050 113.400 ;
        RECT 480.750 112.500 481.800 113.400 ;
        RECT 469.950 110.400 472.050 112.500 ;
        RECT 403.950 98.550 411.450 99.450 ;
        RECT 403.950 97.950 406.050 98.550 ;
        RECT 398.100 94.500 403.200 95.400 ;
        RECT 392.400 92.400 400.200 93.300 ;
        RECT 379.800 81.600 381.600 87.600 ;
        RECT 382.800 81.000 384.600 87.600 ;
        RECT 392.400 81.600 394.200 92.400 ;
        RECT 395.400 81.000 397.200 91.500 ;
        RECT 398.400 82.500 400.200 92.400 ;
        RECT 401.400 83.400 403.200 94.500 ;
        RECT 419.400 93.600 420.600 101.100 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 439.950 100.950 442.050 103.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 431.100 99.150 432.900 100.950 ;
        RECT 404.400 82.500 406.200 93.600 ;
        RECT 398.400 81.600 406.200 82.500 ;
        RECT 418.800 81.600 420.600 93.600 ;
        RECT 421.800 81.000 423.600 93.600 ;
        RECT 431.700 81.000 433.500 93.600 ;
        RECT 436.950 87.600 438.150 100.950 ;
        RECT 455.100 99.150 456.900 100.950 ;
        RECT 458.400 93.600 459.300 100.950 ;
        RECT 461.100 99.150 462.900 100.950 ;
        RECT 465.150 95.700 466.050 110.400 ;
        RECT 473.550 109.800 475.350 111.600 ;
        RECT 476.850 111.450 481.800 112.500 ;
        RECT 489.300 112.500 490.350 113.400 ;
        RECT 476.850 110.700 478.650 111.450 ;
        RECT 489.300 111.300 493.050 112.500 ;
        RECT 490.950 110.400 493.050 111.300 ;
        RECT 496.650 110.400 498.450 116.400 ;
        RECT 473.850 108.000 474.900 109.800 ;
        RECT 484.050 108.000 485.850 108.600 ;
        RECT 473.850 106.800 485.850 108.000 ;
        RECT 468.000 105.600 474.900 106.800 ;
        RECT 468.000 104.850 468.900 105.600 ;
        RECT 473.100 105.000 474.900 105.600 ;
        RECT 467.100 103.050 468.900 104.850 ;
        RECT 470.100 103.800 471.900 104.400 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 470.100 102.600 478.050 103.800 ;
        RECT 475.950 100.950 478.050 102.600 ;
        RECT 474.450 95.700 476.250 96.000 ;
        RECT 465.150 95.100 476.250 95.700 ;
        RECT 465.150 94.500 482.850 95.100 ;
        RECT 465.150 93.600 466.050 94.500 ;
        RECT 474.450 94.200 482.850 94.500 ;
        RECT 455.700 92.400 459.300 93.600 ;
        RECT 436.800 81.600 438.600 87.600 ;
        RECT 439.800 81.000 441.600 87.600 ;
        RECT 455.700 81.600 457.500 92.400 ;
        RECT 460.800 81.000 462.600 93.600 ;
        RECT 465.150 81.600 466.950 93.600 ;
        RECT 479.250 92.700 481.050 93.300 ;
        RECT 473.550 91.500 481.050 92.700 ;
        RECT 481.950 92.100 482.850 94.200 ;
        RECT 484.950 94.200 485.850 106.800 ;
        RECT 497.250 103.050 498.450 110.400 ;
        RECT 492.150 101.250 498.450 103.050 ;
        RECT 493.950 100.950 498.450 101.250 ;
        RECT 494.250 95.400 496.050 97.200 ;
        RECT 490.950 94.200 495.150 95.400 ;
        RECT 484.950 93.300 490.050 94.200 ;
        RECT 490.950 93.300 493.050 94.200 ;
        RECT 497.250 93.600 498.450 100.950 ;
        RECT 489.150 92.400 490.050 93.300 ;
        RECT 486.450 92.100 488.250 92.400 ;
        RECT 473.550 90.600 474.750 91.500 ;
        RECT 481.950 91.200 488.250 92.100 ;
        RECT 486.450 90.600 488.250 91.200 ;
        RECT 489.150 90.600 491.850 92.400 ;
        RECT 469.950 88.500 474.750 90.600 ;
        RECT 477.450 89.550 479.250 90.300 ;
        RECT 482.250 89.550 484.050 90.300 ;
        RECT 477.450 88.500 484.050 89.550 ;
        RECT 473.550 87.600 474.750 88.500 ;
        RECT 468.150 81.000 469.950 87.600 ;
        RECT 473.550 81.600 475.350 87.600 ;
        RECT 478.350 81.000 480.150 87.600 ;
        RECT 481.350 81.600 483.150 88.500 ;
        RECT 489.150 87.600 493.050 89.700 ;
        RECT 484.950 81.000 486.750 87.600 ;
        RECT 489.150 81.600 490.950 87.600 ;
        RECT 493.650 81.000 495.450 84.600 ;
        RECT 496.650 81.600 498.450 93.600 ;
        RECT 501.150 110.400 502.950 116.400 ;
        RECT 504.150 113.400 505.950 117.000 ;
        RECT 508.950 114.300 510.750 116.400 ;
        RECT 507.000 113.400 510.750 114.300 ;
        RECT 513.450 113.400 515.250 117.000 ;
        RECT 516.750 113.400 518.550 116.400 ;
        RECT 520.350 113.400 522.150 117.000 ;
        RECT 524.550 113.400 526.350 116.400 ;
        RECT 529.350 113.400 531.150 117.000 ;
        RECT 507.000 112.500 508.050 113.400 ;
        RECT 516.750 112.500 517.800 113.400 ;
        RECT 505.950 110.400 508.050 112.500 ;
        RECT 501.150 95.700 502.050 110.400 ;
        RECT 509.550 109.800 511.350 111.600 ;
        RECT 512.850 111.450 517.800 112.500 ;
        RECT 525.300 112.500 526.350 113.400 ;
        RECT 512.850 110.700 514.650 111.450 ;
        RECT 525.300 111.300 529.050 112.500 ;
        RECT 526.950 110.400 529.050 111.300 ;
        RECT 532.650 110.400 534.450 116.400 ;
        RECT 509.850 108.000 510.900 109.800 ;
        RECT 520.050 108.000 521.850 108.600 ;
        RECT 509.850 106.800 521.850 108.000 ;
        RECT 504.000 105.600 510.900 106.800 ;
        RECT 504.000 104.850 504.900 105.600 ;
        RECT 509.100 105.000 510.900 105.600 ;
        RECT 503.100 103.050 504.900 104.850 ;
        RECT 506.100 103.800 507.900 104.400 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 506.100 102.600 514.050 103.800 ;
        RECT 511.950 100.950 514.050 102.600 ;
        RECT 510.450 95.700 512.250 96.000 ;
        RECT 501.150 95.100 512.250 95.700 ;
        RECT 501.150 94.500 518.850 95.100 ;
        RECT 501.150 93.600 502.050 94.500 ;
        RECT 510.450 94.200 518.850 94.500 ;
        RECT 501.150 81.600 502.950 93.600 ;
        RECT 515.250 92.700 517.050 93.300 ;
        RECT 509.550 91.500 517.050 92.700 ;
        RECT 517.950 92.100 518.850 94.200 ;
        RECT 520.950 94.200 521.850 106.800 ;
        RECT 533.250 103.050 534.450 110.400 ;
        RECT 542.400 107.400 544.200 117.000 ;
        RECT 549.000 108.000 550.800 116.400 ;
        RECT 563.400 110.400 565.200 117.000 ;
        RECT 566.400 110.400 568.200 116.400 ;
        RECT 578.700 110.400 580.500 117.000 ;
        RECT 549.000 106.800 552.300 108.000 ;
        RECT 542.100 103.200 543.900 105.000 ;
        RECT 548.100 103.200 549.900 105.000 ;
        RECT 551.400 103.200 552.300 106.800 ;
        RECT 553.950 105.450 558.000 106.050 ;
        RECT 553.950 103.950 558.450 105.450 ;
        RECT 528.150 101.250 534.450 103.050 ;
        RECT 529.950 100.950 534.450 101.250 ;
        RECT 541.950 101.100 544.050 103.200 ;
        RECT 544.950 101.100 547.050 103.200 ;
        RECT 547.950 101.100 550.050 103.200 ;
        RECT 550.950 101.100 553.050 103.200 ;
        RECT 530.250 95.400 532.050 97.200 ;
        RECT 526.950 94.200 531.150 95.400 ;
        RECT 520.950 93.300 526.050 94.200 ;
        RECT 526.950 93.300 529.050 94.200 ;
        RECT 533.250 93.600 534.450 100.950 ;
        RECT 535.950 99.450 538.050 100.050 ;
        RECT 541.950 99.450 544.050 100.050 ;
        RECT 535.950 98.550 544.050 99.450 ;
        RECT 545.100 99.300 546.900 101.100 ;
        RECT 535.950 97.950 538.050 98.550 ;
        RECT 541.950 97.950 544.050 98.550 ;
        RECT 525.150 92.400 526.050 93.300 ;
        RECT 522.450 92.100 524.250 92.400 ;
        RECT 509.550 90.600 510.750 91.500 ;
        RECT 517.950 91.200 524.250 92.100 ;
        RECT 522.450 90.600 524.250 91.200 ;
        RECT 525.150 90.600 527.850 92.400 ;
        RECT 505.950 88.500 510.750 90.600 ;
        RECT 513.450 89.550 515.250 90.300 ;
        RECT 518.250 89.550 520.050 90.300 ;
        RECT 513.450 88.500 520.050 89.550 ;
        RECT 509.550 87.600 510.750 88.500 ;
        RECT 504.150 81.000 505.950 87.600 ;
        RECT 509.550 81.600 511.350 87.600 ;
        RECT 514.350 81.000 516.150 87.600 ;
        RECT 517.350 81.600 519.150 88.500 ;
        RECT 525.150 87.600 529.050 89.700 ;
        RECT 520.950 81.000 522.750 87.600 ;
        RECT 525.150 81.600 526.950 87.600 ;
        RECT 529.650 81.000 531.450 84.600 ;
        RECT 532.650 81.600 534.450 93.600 ;
        RECT 538.950 93.450 541.050 94.050 ;
        RECT 547.950 93.450 550.050 94.050 ;
        RECT 538.950 92.550 550.050 93.450 ;
        RECT 538.950 91.950 541.050 92.550 ;
        RECT 547.950 91.950 550.050 92.550 ;
        RECT 551.400 88.800 552.300 101.100 ;
        RECT 557.550 100.050 558.450 103.950 ;
        RECT 563.100 103.200 564.900 105.000 ;
        RECT 566.400 103.200 567.600 110.400 ;
        RECT 583.800 109.200 585.600 116.400 ;
        RECT 581.400 108.300 585.600 109.200 ;
        RECT 596.400 113.400 598.200 116.400 ;
        RECT 599.400 113.400 601.200 117.000 ;
        RECT 596.400 109.500 597.600 113.400 ;
        RECT 602.400 110.400 604.200 116.400 ;
        RECT 596.400 108.600 602.100 109.500 ;
        RECT 578.100 103.200 579.900 105.000 ;
        RECT 581.400 103.200 582.600 108.300 ;
        RECT 600.150 107.700 602.100 108.600 ;
        RECT 584.100 103.200 585.900 105.000 ;
        RECT 562.950 101.100 565.050 103.200 ;
        RECT 565.950 101.100 568.050 103.200 ;
        RECT 577.950 101.100 580.050 103.200 ;
        RECT 580.950 101.100 583.050 103.200 ;
        RECT 583.950 101.100 586.050 103.200 ;
        RECT 553.950 98.550 558.450 100.050 ;
        RECT 553.950 97.950 558.000 98.550 ;
        RECT 566.400 93.600 567.600 101.100 ;
        RECT 545.700 87.900 552.300 88.800 ;
        RECT 545.700 87.600 547.200 87.900 ;
        RECT 542.400 81.000 544.200 87.600 ;
        RECT 545.400 81.600 547.200 87.600 ;
        RECT 551.400 87.600 552.300 87.900 ;
        RECT 548.400 81.000 550.200 87.000 ;
        RECT 551.400 81.600 553.200 87.600 ;
        RECT 563.400 81.000 565.200 93.600 ;
        RECT 566.400 81.600 568.200 93.600 ;
        RECT 581.400 87.600 582.600 101.100 ;
        RECT 595.950 100.950 598.050 103.050 ;
        RECT 596.100 99.150 597.900 100.950 ;
        RECT 600.150 96.300 601.050 107.700 ;
        RECT 603.000 103.050 604.200 110.400 ;
        RECT 614.400 113.400 616.200 116.400 ;
        RECT 617.400 113.400 619.200 117.000 ;
        RECT 614.400 109.500 615.600 113.400 ;
        RECT 620.400 110.400 622.200 116.400 ;
        RECT 614.400 108.600 620.100 109.500 ;
        RECT 618.150 107.700 620.100 108.600 ;
        RECT 601.950 100.950 604.200 103.050 ;
        RECT 613.950 100.950 616.050 103.050 ;
        RECT 600.150 95.400 602.100 96.300 ;
        RECT 596.400 94.500 602.100 95.400 ;
        RECT 596.400 87.600 597.600 94.500 ;
        RECT 603.000 93.600 604.200 100.950 ;
        RECT 614.100 99.150 615.900 100.950 ;
        RECT 618.150 96.300 619.050 107.700 ;
        RECT 621.000 103.050 622.200 110.400 ;
        RECT 632.400 113.400 634.200 116.400 ;
        RECT 635.400 113.400 637.200 117.000 ;
        RECT 632.400 109.500 633.600 113.400 ;
        RECT 638.400 110.400 640.200 116.400 ;
        RECT 652.800 110.400 654.600 116.400 ;
        RECT 632.400 108.600 638.100 109.500 ;
        RECT 636.150 107.700 638.100 108.600 ;
        RECT 627.000 105.450 631.050 106.050 ;
        RECT 619.950 100.950 622.200 103.050 ;
        RECT 618.150 95.400 620.100 96.300 ;
        RECT 578.400 81.000 580.200 87.600 ;
        RECT 581.400 81.600 583.200 87.600 ;
        RECT 584.400 81.000 586.200 87.600 ;
        RECT 596.400 81.600 598.200 87.600 ;
        RECT 599.400 81.000 601.200 87.600 ;
        RECT 602.400 81.600 604.200 93.600 ;
        RECT 614.400 94.500 620.100 95.400 ;
        RECT 614.400 87.600 615.600 94.500 ;
        RECT 621.000 93.600 622.200 100.950 ;
        RECT 626.550 103.950 631.050 105.450 ;
        RECT 626.550 100.050 627.450 103.950 ;
        RECT 631.950 100.950 634.050 103.050 ;
        RECT 626.550 98.550 631.050 100.050 ;
        RECT 632.100 99.150 633.900 100.950 ;
        RECT 627.000 97.950 631.050 98.550 ;
        RECT 636.150 96.300 637.050 107.700 ;
        RECT 639.000 103.050 640.200 110.400 ;
        RECT 653.400 108.300 654.600 110.400 ;
        RECT 655.800 111.300 657.600 116.400 ;
        RECT 658.800 112.200 660.600 117.000 ;
        RECT 661.800 111.300 663.600 116.400 ;
        RECT 655.800 109.950 663.600 111.300 ;
        RECT 673.800 110.400 675.600 116.400 ;
        RECT 674.400 108.300 675.600 110.400 ;
        RECT 676.800 111.300 678.600 116.400 ;
        RECT 679.800 112.200 681.600 117.000 ;
        RECT 682.800 111.300 684.600 116.400 ;
        RECT 676.800 109.950 684.600 111.300 ;
        RECT 694.800 110.400 696.600 116.400 ;
        RECT 695.400 108.300 696.600 110.400 ;
        RECT 697.800 111.300 699.600 116.400 ;
        RECT 700.800 112.200 702.600 117.000 ;
        RECT 703.800 111.300 705.600 116.400 ;
        RECT 697.800 109.950 705.600 111.300 ;
        RECT 713.700 110.400 715.500 117.000 ;
        RECT 718.800 109.200 720.600 116.400 ;
        RECT 733.800 113.400 735.600 116.400 ;
        RECT 736.800 113.400 738.600 117.000 ;
        RECT 716.400 108.300 720.600 109.200 ;
        RECT 653.400 107.250 657.150 108.300 ;
        RECT 674.400 107.250 678.150 108.300 ;
        RECT 695.400 107.250 699.150 108.300 ;
        RECT 648.000 105.450 652.050 106.050 ;
        RECT 637.950 100.950 640.200 103.050 ;
        RECT 636.150 95.400 638.100 96.300 ;
        RECT 614.400 81.600 616.200 87.600 ;
        RECT 617.400 81.000 619.200 87.600 ;
        RECT 620.400 81.600 622.200 93.600 ;
        RECT 632.400 94.500 638.100 95.400 ;
        RECT 632.400 87.600 633.600 94.500 ;
        RECT 639.000 93.600 640.200 100.950 ;
        RECT 647.550 103.950 652.050 105.450 ;
        RECT 647.550 100.050 648.450 103.950 ;
        RECT 653.100 103.050 654.900 104.850 ;
        RECT 655.950 103.050 657.150 107.250 ;
        RECT 659.100 103.050 660.900 104.850 ;
        RECT 674.100 103.050 675.900 104.850 ;
        RECT 676.950 103.050 678.150 107.250 ;
        RECT 680.100 103.050 681.900 104.850 ;
        RECT 695.100 103.050 696.900 104.850 ;
        RECT 697.950 103.050 699.150 107.250 ;
        RECT 701.100 103.050 702.900 104.850 ;
        RECT 713.100 103.200 714.900 105.000 ;
        RECT 716.400 103.200 717.600 108.300 ;
        RECT 719.100 103.200 720.900 105.000 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 676.950 100.950 679.050 103.050 ;
        RECT 679.950 100.950 682.050 103.050 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 694.950 100.950 697.050 103.050 ;
        RECT 697.950 100.950 700.050 103.050 ;
        RECT 700.950 100.950 703.050 103.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 712.950 101.100 715.050 103.200 ;
        RECT 715.950 101.100 718.050 103.200 ;
        RECT 718.950 101.100 721.050 103.200 ;
        RECT 734.400 103.050 735.600 113.400 ;
        RECT 740.550 110.400 742.350 116.400 ;
        RECT 743.850 113.400 745.650 117.000 ;
        RECT 748.650 113.400 750.450 116.400 ;
        RECT 752.850 113.400 754.650 117.000 ;
        RECT 756.450 113.400 758.250 116.400 ;
        RECT 759.750 113.400 761.550 117.000 ;
        RECT 764.250 114.300 766.050 116.400 ;
        RECT 764.250 113.400 768.000 114.300 ;
        RECT 769.050 113.400 770.850 117.000 ;
        RECT 748.650 112.500 749.700 113.400 ;
        RECT 745.950 111.300 749.700 112.500 ;
        RECT 757.200 112.500 758.250 113.400 ;
        RECT 766.950 112.500 768.000 113.400 ;
        RECT 757.200 111.450 762.150 112.500 ;
        RECT 745.950 110.400 748.050 111.300 ;
        RECT 760.350 110.700 762.150 111.450 ;
        RECT 740.550 103.050 741.750 110.400 ;
        RECT 763.650 109.800 765.450 111.600 ;
        RECT 766.950 110.400 769.050 112.500 ;
        RECT 772.050 110.400 773.850 116.400 ;
        RECT 753.150 108.000 754.950 108.600 ;
        RECT 764.100 108.000 765.150 109.800 ;
        RECT 753.150 106.800 765.150 108.000 ;
        RECT 647.550 98.550 652.050 100.050 ;
        RECT 648.000 97.950 652.050 98.550 ;
        RECT 632.400 81.600 634.200 87.600 ;
        RECT 635.400 81.000 637.200 87.600 ;
        RECT 638.400 81.600 640.200 93.600 ;
        RECT 656.850 87.600 658.050 100.950 ;
        RECT 662.100 99.150 663.900 100.950 ;
        RECT 653.400 81.000 655.200 87.600 ;
        RECT 656.400 81.600 658.200 87.600 ;
        RECT 661.500 81.000 663.300 93.600 ;
        RECT 677.850 87.600 679.050 100.950 ;
        RECT 683.100 99.150 684.900 100.950 ;
        RECT 674.400 81.000 676.200 87.600 ;
        RECT 677.400 81.600 679.200 87.600 ;
        RECT 682.500 81.000 684.300 93.600 ;
        RECT 698.850 87.600 700.050 100.950 ;
        RECT 704.100 99.150 705.900 100.950 ;
        RECT 695.400 81.000 697.200 87.600 ;
        RECT 698.400 81.600 700.200 87.600 ;
        RECT 703.500 81.000 705.300 93.600 ;
        RECT 716.400 87.600 717.600 101.100 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 740.550 101.250 746.850 103.050 ;
        RECT 740.550 100.950 745.050 101.250 ;
        RECT 734.400 87.600 735.600 100.950 ;
        RECT 737.100 99.150 738.900 100.950 ;
        RECT 740.550 93.600 741.750 100.950 ;
        RECT 742.950 95.400 744.750 97.200 ;
        RECT 743.850 94.200 748.050 95.400 ;
        RECT 753.150 94.200 754.050 106.800 ;
        RECT 764.100 105.600 771.000 106.800 ;
        RECT 764.100 105.000 765.900 105.600 ;
        RECT 770.100 104.850 771.000 105.600 ;
        RECT 767.100 103.800 768.900 104.400 ;
        RECT 760.950 102.600 768.900 103.800 ;
        RECT 770.100 103.050 771.900 104.850 ;
        RECT 760.950 100.950 763.050 102.600 ;
        RECT 769.950 100.950 772.050 103.050 ;
        RECT 762.750 95.700 764.550 96.000 ;
        RECT 772.950 95.700 773.850 110.400 ;
        RECT 782.400 111.300 784.200 116.400 ;
        RECT 785.400 112.200 787.200 117.000 ;
        RECT 788.400 111.300 790.200 116.400 ;
        RECT 782.400 109.950 790.200 111.300 ;
        RECT 791.400 110.400 793.200 116.400 ;
        RECT 803.700 110.400 805.500 117.000 ;
        RECT 791.400 108.300 792.600 110.400 ;
        RECT 808.800 109.200 810.600 116.400 ;
        RECT 788.850 107.250 792.600 108.300 ;
        RECT 806.400 108.300 810.600 109.200 ;
        RECT 815.550 110.400 817.350 116.400 ;
        RECT 818.850 113.400 820.650 117.000 ;
        RECT 823.650 113.400 825.450 116.400 ;
        RECT 827.850 113.400 829.650 117.000 ;
        RECT 831.450 113.400 833.250 116.400 ;
        RECT 834.750 113.400 836.550 117.000 ;
        RECT 839.250 114.300 841.050 116.400 ;
        RECT 839.250 113.400 843.000 114.300 ;
        RECT 844.050 113.400 845.850 117.000 ;
        RECT 823.650 112.500 824.700 113.400 ;
        RECT 820.950 111.300 824.700 112.500 ;
        RECT 832.200 112.500 833.250 113.400 ;
        RECT 841.950 112.500 843.000 113.400 ;
        RECT 832.200 111.450 837.150 112.500 ;
        RECT 820.950 110.400 823.050 111.300 ;
        RECT 835.350 110.700 837.150 111.450 ;
        RECT 785.100 103.050 786.900 104.850 ;
        RECT 788.850 103.050 790.050 107.250 ;
        RECT 791.100 103.050 792.900 104.850 ;
        RECT 803.100 103.200 804.900 105.000 ;
        RECT 806.400 103.200 807.600 108.300 ;
        RECT 809.100 103.200 810.900 105.000 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 784.950 100.950 787.050 103.050 ;
        RECT 787.950 100.950 790.050 103.050 ;
        RECT 790.950 100.950 793.050 103.050 ;
        RECT 802.950 101.100 805.050 103.200 ;
        RECT 805.950 101.100 808.050 103.200 ;
        RECT 808.950 101.100 811.050 103.200 ;
        RECT 815.550 103.050 816.750 110.400 ;
        RECT 838.650 109.800 840.450 111.600 ;
        RECT 841.950 110.400 844.050 112.500 ;
        RECT 847.050 110.400 848.850 116.400 ;
        RECT 828.150 108.000 829.950 108.600 ;
        RECT 839.100 108.000 840.150 109.800 ;
        RECT 828.150 106.800 840.150 108.000 ;
        RECT 815.550 101.250 821.850 103.050 ;
        RECT 782.100 99.150 783.900 100.950 ;
        RECT 762.750 95.100 773.850 95.700 ;
        RECT 713.400 81.000 715.200 87.600 ;
        RECT 716.400 81.600 718.200 87.600 ;
        RECT 719.400 81.000 721.200 87.600 ;
        RECT 733.800 81.600 735.600 87.600 ;
        RECT 736.800 81.000 738.600 87.600 ;
        RECT 740.550 81.600 742.350 93.600 ;
        RECT 745.950 93.300 748.050 94.200 ;
        RECT 748.950 93.300 754.050 94.200 ;
        RECT 756.150 94.500 773.850 95.100 ;
        RECT 756.150 94.200 764.550 94.500 ;
        RECT 748.950 92.400 749.850 93.300 ;
        RECT 747.150 90.600 749.850 92.400 ;
        RECT 750.750 92.100 752.550 92.400 ;
        RECT 756.150 92.100 757.050 94.200 ;
        RECT 772.950 93.600 773.850 94.500 ;
        RECT 750.750 91.200 757.050 92.100 ;
        RECT 757.950 92.700 759.750 93.300 ;
        RECT 757.950 91.500 765.450 92.700 ;
        RECT 750.750 90.600 752.550 91.200 ;
        RECT 764.250 90.600 765.450 91.500 ;
        RECT 745.950 87.600 749.850 89.700 ;
        RECT 754.950 89.550 756.750 90.300 ;
        RECT 759.750 89.550 761.550 90.300 ;
        RECT 754.950 88.500 761.550 89.550 ;
        RECT 764.250 88.500 769.050 90.600 ;
        RECT 743.550 81.000 745.350 84.600 ;
        RECT 748.050 81.600 749.850 87.600 ;
        RECT 752.250 81.000 754.050 87.600 ;
        RECT 755.850 81.600 757.650 88.500 ;
        RECT 764.250 87.600 765.450 88.500 ;
        RECT 758.850 81.000 760.650 87.600 ;
        RECT 763.650 81.600 765.450 87.600 ;
        RECT 769.050 81.000 770.850 87.600 ;
        RECT 772.050 81.600 773.850 93.600 ;
        RECT 782.700 81.000 784.500 93.600 ;
        RECT 787.950 87.600 789.150 100.950 ;
        RECT 806.400 87.600 807.600 101.100 ;
        RECT 815.550 100.950 820.050 101.250 ;
        RECT 815.550 93.600 816.750 100.950 ;
        RECT 817.950 95.400 819.750 97.200 ;
        RECT 818.850 94.200 823.050 95.400 ;
        RECT 828.150 94.200 829.050 106.800 ;
        RECT 839.100 105.600 846.000 106.800 ;
        RECT 839.100 105.000 840.900 105.600 ;
        RECT 845.100 104.850 846.000 105.600 ;
        RECT 842.100 103.800 843.900 104.400 ;
        RECT 835.950 102.600 843.900 103.800 ;
        RECT 845.100 103.050 846.900 104.850 ;
        RECT 835.950 100.950 838.050 102.600 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 837.750 95.700 839.550 96.000 ;
        RECT 847.950 95.700 848.850 110.400 ;
        RECT 837.750 95.100 848.850 95.700 ;
        RECT 787.800 81.600 789.600 87.600 ;
        RECT 790.800 81.000 792.600 87.600 ;
        RECT 803.400 81.000 805.200 87.600 ;
        RECT 806.400 81.600 808.200 87.600 ;
        RECT 809.400 81.000 811.200 87.600 ;
        RECT 815.550 81.600 817.350 93.600 ;
        RECT 820.950 93.300 823.050 94.200 ;
        RECT 823.950 93.300 829.050 94.200 ;
        RECT 831.150 94.500 848.850 95.100 ;
        RECT 831.150 94.200 839.550 94.500 ;
        RECT 823.950 92.400 824.850 93.300 ;
        RECT 822.150 90.600 824.850 92.400 ;
        RECT 825.750 92.100 827.550 92.400 ;
        RECT 831.150 92.100 832.050 94.200 ;
        RECT 847.950 93.600 848.850 94.500 ;
        RECT 825.750 91.200 832.050 92.100 ;
        RECT 832.950 92.700 834.750 93.300 ;
        RECT 832.950 91.500 840.450 92.700 ;
        RECT 825.750 90.600 827.550 91.200 ;
        RECT 839.250 90.600 840.450 91.500 ;
        RECT 820.950 87.600 824.850 89.700 ;
        RECT 829.950 89.550 831.750 90.300 ;
        RECT 834.750 89.550 836.550 90.300 ;
        RECT 829.950 88.500 836.550 89.550 ;
        RECT 839.250 88.500 844.050 90.600 ;
        RECT 818.550 81.000 820.350 84.600 ;
        RECT 823.050 81.600 824.850 87.600 ;
        RECT 827.250 81.000 829.050 87.600 ;
        RECT 830.850 81.600 832.650 88.500 ;
        RECT 839.250 87.600 840.450 88.500 ;
        RECT 833.850 81.000 835.650 87.600 ;
        RECT 838.650 81.600 840.450 87.600 ;
        RECT 844.050 81.000 845.850 87.600 ;
        RECT 847.050 81.600 848.850 93.600 ;
        RECT 10.800 71.400 12.600 77.400 ;
        RECT 13.800 71.400 15.600 78.000 ;
        RECT 11.400 58.050 12.600 71.400 ;
        RECT 17.550 65.400 19.350 77.400 ;
        RECT 20.550 74.400 22.350 78.000 ;
        RECT 25.050 71.400 26.850 77.400 ;
        RECT 29.250 71.400 31.050 78.000 ;
        RECT 22.950 69.300 26.850 71.400 ;
        RECT 32.850 70.500 34.650 77.400 ;
        RECT 35.850 71.400 37.650 78.000 ;
        RECT 40.650 71.400 42.450 77.400 ;
        RECT 46.050 71.400 47.850 78.000 ;
        RECT 41.250 70.500 42.450 71.400 ;
        RECT 31.950 69.450 38.550 70.500 ;
        RECT 31.950 68.700 33.750 69.450 ;
        RECT 36.750 68.700 38.550 69.450 ;
        RECT 41.250 68.400 46.050 70.500 ;
        RECT 24.150 66.600 26.850 68.400 ;
        RECT 27.750 67.800 29.550 68.400 ;
        RECT 27.750 66.900 34.050 67.800 ;
        RECT 41.250 67.500 42.450 68.400 ;
        RECT 27.750 66.600 29.550 66.900 ;
        RECT 25.950 65.700 26.850 66.600 ;
        RECT 14.100 58.050 15.900 59.850 ;
        RECT 17.550 58.050 18.750 65.400 ;
        RECT 22.950 64.800 25.050 65.700 ;
        RECT 25.950 64.800 31.050 65.700 ;
        RECT 20.850 63.600 25.050 64.800 ;
        RECT 19.950 61.800 21.750 63.600 ;
        RECT 10.950 55.950 13.050 58.050 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 17.550 57.750 22.050 58.050 ;
        RECT 17.550 55.950 23.850 57.750 ;
        RECT 11.400 45.600 12.600 55.950 ;
        RECT 17.550 48.600 18.750 55.950 ;
        RECT 30.150 52.200 31.050 64.800 ;
        RECT 33.150 64.800 34.050 66.900 ;
        RECT 34.950 66.300 42.450 67.500 ;
        RECT 34.950 65.700 36.750 66.300 ;
        RECT 49.050 65.400 50.850 77.400 ;
        RECT 59.700 65.400 61.500 78.000 ;
        RECT 64.800 71.400 66.600 77.400 ;
        RECT 67.800 71.400 69.600 78.000 ;
        RECT 80.400 71.400 82.200 78.000 ;
        RECT 83.400 71.400 85.200 77.400 ;
        RECT 86.400 71.400 88.200 78.000 ;
        RECT 33.150 64.500 41.550 64.800 ;
        RECT 49.950 64.500 50.850 65.400 ;
        RECT 33.150 63.900 50.850 64.500 ;
        RECT 39.750 63.300 50.850 63.900 ;
        RECT 39.750 63.000 41.550 63.300 ;
        RECT 37.950 56.400 40.050 58.050 ;
        RECT 37.950 55.200 45.900 56.400 ;
        RECT 46.950 55.950 49.050 58.050 ;
        RECT 44.100 54.600 45.900 55.200 ;
        RECT 47.100 54.150 48.900 55.950 ;
        RECT 41.100 53.400 42.900 54.000 ;
        RECT 47.100 53.400 48.000 54.150 ;
        RECT 41.100 52.200 48.000 53.400 ;
        RECT 30.150 51.000 42.150 52.200 ;
        RECT 30.150 50.400 31.950 51.000 ;
        RECT 41.100 49.200 42.150 51.000 ;
        RECT 10.800 42.600 12.600 45.600 ;
        RECT 13.800 42.000 15.600 45.600 ;
        RECT 17.550 42.600 19.350 48.600 ;
        RECT 22.950 47.700 25.050 48.600 ;
        RECT 22.950 46.500 26.700 47.700 ;
        RECT 37.350 47.550 39.150 48.300 ;
        RECT 25.650 45.600 26.700 46.500 ;
        RECT 34.200 46.500 39.150 47.550 ;
        RECT 40.650 47.400 42.450 49.200 ;
        RECT 49.950 48.600 50.850 63.300 ;
        RECT 59.100 58.050 60.900 59.850 ;
        RECT 64.950 58.050 66.150 71.400 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 83.400 57.900 84.600 71.400 ;
        RECT 92.550 65.400 94.350 77.400 ;
        RECT 95.550 74.400 97.350 78.000 ;
        RECT 100.050 71.400 101.850 77.400 ;
        RECT 104.250 71.400 106.050 78.000 ;
        RECT 97.950 69.300 101.850 71.400 ;
        RECT 107.850 70.500 109.650 77.400 ;
        RECT 110.850 71.400 112.650 78.000 ;
        RECT 115.650 71.400 117.450 77.400 ;
        RECT 121.050 71.400 122.850 78.000 ;
        RECT 116.250 70.500 117.450 71.400 ;
        RECT 106.950 69.450 113.550 70.500 ;
        RECT 106.950 68.700 108.750 69.450 ;
        RECT 111.750 68.700 113.550 69.450 ;
        RECT 116.250 68.400 121.050 70.500 ;
        RECT 99.150 66.600 101.850 68.400 ;
        RECT 102.750 67.800 104.550 68.400 ;
        RECT 102.750 66.900 109.050 67.800 ;
        RECT 116.250 67.500 117.450 68.400 ;
        RECT 102.750 66.600 104.550 66.900 ;
        RECT 100.950 65.700 101.850 66.600 ;
        RECT 92.550 58.050 93.750 65.400 ;
        RECT 97.950 64.800 100.050 65.700 ;
        RECT 100.950 64.800 106.050 65.700 ;
        RECT 95.850 63.600 100.050 64.800 ;
        RECT 94.950 61.800 96.750 63.600 ;
        RECT 62.100 54.150 63.900 55.950 ;
        RECT 65.850 51.750 67.050 55.950 ;
        RECT 68.100 54.150 69.900 55.950 ;
        RECT 79.950 55.800 82.050 57.900 ;
        RECT 82.950 55.800 85.050 57.900 ;
        RECT 85.950 55.800 88.050 57.900 ;
        RECT 92.550 57.750 97.050 58.050 ;
        RECT 92.550 55.950 98.850 57.750 ;
        RECT 80.100 54.000 81.900 55.800 ;
        RECT 65.850 50.700 69.600 51.750 ;
        RECT 43.950 46.500 46.050 48.600 ;
        RECT 34.200 45.600 35.250 46.500 ;
        RECT 43.950 45.600 45.000 46.500 ;
        RECT 20.850 42.000 22.650 45.600 ;
        RECT 25.650 42.600 27.450 45.600 ;
        RECT 29.850 42.000 31.650 45.600 ;
        RECT 33.450 42.600 35.250 45.600 ;
        RECT 36.750 42.000 38.550 45.600 ;
        RECT 41.250 44.700 45.000 45.600 ;
        RECT 41.250 42.600 43.050 44.700 ;
        RECT 46.050 42.000 47.850 45.600 ;
        RECT 49.050 42.600 50.850 48.600 ;
        RECT 59.400 47.700 67.200 49.050 ;
        RECT 59.400 42.600 61.200 47.700 ;
        RECT 62.400 42.000 64.200 46.800 ;
        RECT 65.400 42.600 67.200 47.700 ;
        RECT 68.400 48.600 69.600 50.700 ;
        RECT 83.400 50.700 84.600 55.800 ;
        RECT 86.100 54.000 87.900 55.800 ;
        RECT 83.400 49.800 87.600 50.700 ;
        RECT 68.400 42.600 70.200 48.600 ;
        RECT 80.700 42.000 82.500 48.600 ;
        RECT 85.800 42.600 87.600 49.800 ;
        RECT 92.550 48.600 93.750 55.950 ;
        RECT 105.150 52.200 106.050 64.800 ;
        RECT 108.150 64.800 109.050 66.900 ;
        RECT 109.950 66.300 117.450 67.500 ;
        RECT 109.950 65.700 111.750 66.300 ;
        RECT 124.050 65.400 125.850 77.400 ;
        RECT 137.700 66.600 139.500 77.400 ;
        RECT 137.700 65.400 141.300 66.600 ;
        RECT 142.800 65.400 144.600 78.000 ;
        RECT 154.800 65.400 156.600 77.400 ;
        RECT 157.800 66.300 159.600 77.400 ;
        RECT 160.800 67.200 162.600 78.000 ;
        RECT 163.800 66.300 165.600 77.400 ;
        RECT 157.800 65.400 165.600 66.300 ;
        RECT 168.150 65.400 169.950 77.400 ;
        RECT 171.150 71.400 172.950 78.000 ;
        RECT 176.550 71.400 178.350 77.400 ;
        RECT 181.350 71.400 183.150 78.000 ;
        RECT 176.550 70.500 177.750 71.400 ;
        RECT 184.350 70.500 186.150 77.400 ;
        RECT 187.950 71.400 189.750 78.000 ;
        RECT 192.150 71.400 193.950 77.400 ;
        RECT 196.650 74.400 198.450 78.000 ;
        RECT 172.950 68.400 177.750 70.500 ;
        RECT 180.450 69.450 187.050 70.500 ;
        RECT 180.450 68.700 182.250 69.450 ;
        RECT 185.250 68.700 187.050 69.450 ;
        RECT 192.150 69.300 196.050 71.400 ;
        RECT 176.550 67.500 177.750 68.400 ;
        RECT 189.450 67.800 191.250 68.400 ;
        RECT 176.550 66.300 184.050 67.500 ;
        RECT 182.250 65.700 184.050 66.300 ;
        RECT 184.950 66.900 191.250 67.800 ;
        RECT 108.150 64.500 116.550 64.800 ;
        RECT 124.950 64.500 125.850 65.400 ;
        RECT 108.150 63.900 125.850 64.500 ;
        RECT 114.750 63.300 125.850 63.900 ;
        RECT 114.750 63.000 116.550 63.300 ;
        RECT 112.950 56.400 115.050 58.050 ;
        RECT 112.950 55.200 120.900 56.400 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 119.100 54.600 120.900 55.200 ;
        RECT 122.100 54.150 123.900 55.950 ;
        RECT 116.100 53.400 117.900 54.000 ;
        RECT 122.100 53.400 123.000 54.150 ;
        RECT 116.100 52.200 123.000 53.400 ;
        RECT 105.150 51.000 117.150 52.200 ;
        RECT 105.150 50.400 106.950 51.000 ;
        RECT 116.100 49.200 117.150 51.000 ;
        RECT 92.550 42.600 94.350 48.600 ;
        RECT 97.950 47.700 100.050 48.600 ;
        RECT 97.950 46.500 101.700 47.700 ;
        RECT 112.350 47.550 114.150 48.300 ;
        RECT 100.650 45.600 101.700 46.500 ;
        RECT 109.200 46.500 114.150 47.550 ;
        RECT 115.650 47.400 117.450 49.200 ;
        RECT 124.950 48.600 125.850 63.300 ;
        RECT 137.100 58.050 138.900 59.850 ;
        RECT 140.400 58.050 141.300 65.400 ;
        RECT 143.100 58.050 144.900 59.850 ;
        RECT 136.950 55.950 139.050 58.050 ;
        RECT 139.950 55.950 142.050 58.050 ;
        RECT 142.950 55.950 145.050 58.050 ;
        RECT 155.400 57.900 156.300 65.400 ;
        RECT 168.150 64.500 169.050 65.400 ;
        RECT 184.950 64.800 185.850 66.900 ;
        RECT 189.450 66.600 191.250 66.900 ;
        RECT 192.150 66.600 194.850 68.400 ;
        RECT 192.150 65.700 193.050 66.600 ;
        RECT 177.450 64.500 185.850 64.800 ;
        RECT 168.150 63.900 185.850 64.500 ;
        RECT 187.950 64.800 193.050 65.700 ;
        RECT 193.950 64.800 196.050 65.700 ;
        RECT 199.650 65.400 201.450 77.400 ;
        RECT 211.800 65.400 213.600 77.400 ;
        RECT 214.800 66.300 216.600 77.400 ;
        RECT 217.800 67.200 219.600 78.000 ;
        RECT 220.800 66.300 222.600 77.400 ;
        RECT 214.800 65.400 222.600 66.300 ;
        RECT 224.550 65.400 226.350 77.400 ;
        RECT 227.550 74.400 229.350 78.000 ;
        RECT 232.050 71.400 233.850 77.400 ;
        RECT 236.250 71.400 238.050 78.000 ;
        RECT 229.950 69.300 233.850 71.400 ;
        RECT 239.850 70.500 241.650 77.400 ;
        RECT 242.850 71.400 244.650 78.000 ;
        RECT 247.650 71.400 249.450 77.400 ;
        RECT 253.050 71.400 254.850 78.000 ;
        RECT 248.250 70.500 249.450 71.400 ;
        RECT 238.950 69.450 245.550 70.500 ;
        RECT 238.950 68.700 240.750 69.450 ;
        RECT 243.750 68.700 245.550 69.450 ;
        RECT 248.250 68.400 253.050 70.500 ;
        RECT 231.150 66.600 233.850 68.400 ;
        RECT 234.750 67.800 236.550 68.400 ;
        RECT 234.750 66.900 241.050 67.800 ;
        RECT 248.250 67.500 249.450 68.400 ;
        RECT 234.750 66.600 236.550 66.900 ;
        RECT 232.950 65.700 233.850 66.600 ;
        RECT 168.150 63.300 179.250 63.900 ;
        RECT 161.100 57.900 162.900 59.700 ;
        RECT 127.950 51.450 130.050 52.050 ;
        RECT 136.950 51.450 139.050 52.050 ;
        RECT 127.950 50.550 139.050 51.450 ;
        RECT 127.950 49.950 130.050 50.550 ;
        RECT 136.950 49.950 139.050 50.550 ;
        RECT 118.950 46.500 121.050 48.600 ;
        RECT 109.200 45.600 110.250 46.500 ;
        RECT 118.950 45.600 120.000 46.500 ;
        RECT 95.850 42.000 97.650 45.600 ;
        RECT 100.650 42.600 102.450 45.600 ;
        RECT 104.850 42.000 106.650 45.600 ;
        RECT 108.450 42.600 110.250 45.600 ;
        RECT 111.750 42.000 113.550 45.600 ;
        RECT 116.250 44.700 120.000 45.600 ;
        RECT 116.250 42.600 118.050 44.700 ;
        RECT 121.050 42.000 122.850 45.600 ;
        RECT 124.050 42.600 125.850 48.600 ;
        RECT 140.400 45.600 141.300 55.950 ;
        RECT 154.950 55.800 157.050 57.900 ;
        RECT 157.950 55.800 160.050 57.900 ;
        RECT 160.950 55.800 163.050 57.900 ;
        RECT 163.950 55.800 166.050 57.900 ;
        RECT 155.400 48.600 156.300 55.800 ;
        RECT 158.100 54.000 159.900 55.800 ;
        RECT 164.100 54.000 165.900 55.800 ;
        RECT 168.150 48.600 169.050 63.300 ;
        RECT 177.450 63.000 179.250 63.300 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 178.950 56.400 181.050 58.050 ;
        RECT 170.100 54.150 171.900 55.950 ;
        RECT 173.100 55.200 181.050 56.400 ;
        RECT 173.100 54.600 174.900 55.200 ;
        RECT 171.000 53.400 171.900 54.150 ;
        RECT 176.100 53.400 177.900 54.000 ;
        RECT 171.000 52.200 177.900 53.400 ;
        RECT 187.950 52.200 188.850 64.800 ;
        RECT 193.950 63.600 198.150 64.800 ;
        RECT 197.250 61.800 199.050 63.600 ;
        RECT 200.250 58.050 201.450 65.400 ;
        RECT 196.950 57.750 201.450 58.050 ;
        RECT 212.400 57.900 213.300 65.400 ;
        RECT 218.100 57.900 219.900 59.700 ;
        RECT 224.550 58.050 225.750 65.400 ;
        RECT 229.950 64.800 232.050 65.700 ;
        RECT 232.950 64.800 238.050 65.700 ;
        RECT 227.850 63.600 232.050 64.800 ;
        RECT 226.950 61.800 228.750 63.600 ;
        RECT 195.150 55.950 201.450 57.750 ;
        RECT 176.850 51.000 188.850 52.200 ;
        RECT 176.850 49.200 177.900 51.000 ;
        RECT 187.050 50.400 188.850 51.000 ;
        RECT 155.400 47.400 160.500 48.600 ;
        RECT 136.800 42.000 138.600 45.600 ;
        RECT 139.800 42.600 141.600 45.600 ;
        RECT 142.800 42.000 144.600 45.600 ;
        RECT 155.700 42.000 157.500 45.600 ;
        RECT 158.700 42.600 160.500 47.400 ;
        RECT 163.200 42.000 165.000 48.600 ;
        RECT 168.150 42.600 169.950 48.600 ;
        RECT 172.950 46.500 175.050 48.600 ;
        RECT 176.550 47.400 178.350 49.200 ;
        RECT 200.250 48.600 201.450 55.950 ;
        RECT 211.950 55.800 214.050 57.900 ;
        RECT 214.950 55.800 217.050 57.900 ;
        RECT 217.950 55.800 220.050 57.900 ;
        RECT 220.950 55.800 223.050 57.900 ;
        RECT 224.550 57.750 229.050 58.050 ;
        RECT 224.550 55.950 230.850 57.750 ;
        RECT 179.850 47.550 181.650 48.300 ;
        RECT 193.950 47.700 196.050 48.600 ;
        RECT 179.850 46.500 184.800 47.550 ;
        RECT 174.000 45.600 175.050 46.500 ;
        RECT 183.750 45.600 184.800 46.500 ;
        RECT 192.300 46.500 196.050 47.700 ;
        RECT 192.300 45.600 193.350 46.500 ;
        RECT 171.150 42.000 172.950 45.600 ;
        RECT 174.000 44.700 177.750 45.600 ;
        RECT 175.950 42.600 177.750 44.700 ;
        RECT 180.450 42.000 182.250 45.600 ;
        RECT 183.750 42.600 185.550 45.600 ;
        RECT 187.350 42.000 189.150 45.600 ;
        RECT 191.550 42.600 193.350 45.600 ;
        RECT 196.350 42.000 198.150 45.600 ;
        RECT 199.650 42.600 201.450 48.600 ;
        RECT 212.400 48.600 213.300 55.800 ;
        RECT 215.100 54.000 216.900 55.800 ;
        RECT 221.100 54.000 222.900 55.800 ;
        RECT 224.550 48.600 225.750 55.950 ;
        RECT 237.150 52.200 238.050 64.800 ;
        RECT 240.150 64.800 241.050 66.900 ;
        RECT 241.950 66.300 249.450 67.500 ;
        RECT 241.950 65.700 243.750 66.300 ;
        RECT 256.050 65.400 257.850 77.400 ;
        RECT 266.700 65.400 268.500 78.000 ;
        RECT 271.800 71.400 273.600 77.400 ;
        RECT 274.800 71.400 276.600 78.000 ;
        RECT 287.400 71.400 289.200 78.000 ;
        RECT 290.400 71.400 292.200 77.400 ;
        RECT 293.400 71.400 295.200 78.000 ;
        RECT 307.800 71.400 309.600 78.000 ;
        RECT 310.800 71.400 312.600 77.400 ;
        RECT 313.800 71.400 315.600 78.000 ;
        RECT 326.400 71.400 328.200 78.000 ;
        RECT 329.400 71.400 331.200 77.400 ;
        RECT 240.150 64.500 248.550 64.800 ;
        RECT 256.950 64.500 257.850 65.400 ;
        RECT 240.150 63.900 257.850 64.500 ;
        RECT 246.750 63.300 257.850 63.900 ;
        RECT 246.750 63.000 248.550 63.300 ;
        RECT 244.950 56.400 247.050 58.050 ;
        RECT 244.950 55.200 252.900 56.400 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 251.100 54.600 252.900 55.200 ;
        RECT 254.100 54.150 255.900 55.950 ;
        RECT 248.100 53.400 249.900 54.000 ;
        RECT 254.100 53.400 255.000 54.150 ;
        RECT 248.100 52.200 255.000 53.400 ;
        RECT 237.150 51.000 249.150 52.200 ;
        RECT 237.150 50.400 238.950 51.000 ;
        RECT 248.100 49.200 249.150 51.000 ;
        RECT 212.400 47.400 217.500 48.600 ;
        RECT 212.700 42.000 214.500 45.600 ;
        RECT 215.700 42.600 217.500 47.400 ;
        RECT 220.200 42.000 222.000 48.600 ;
        RECT 224.550 42.600 226.350 48.600 ;
        RECT 229.950 47.700 232.050 48.600 ;
        RECT 229.950 46.500 233.700 47.700 ;
        RECT 244.350 47.550 246.150 48.300 ;
        RECT 232.650 45.600 233.700 46.500 ;
        RECT 241.200 46.500 246.150 47.550 ;
        RECT 247.650 47.400 249.450 49.200 ;
        RECT 256.950 48.600 257.850 63.300 ;
        RECT 259.950 63.450 262.050 63.900 ;
        RECT 265.950 63.450 268.050 64.050 ;
        RECT 259.950 62.550 268.050 63.450 ;
        RECT 259.950 61.800 262.050 62.550 ;
        RECT 265.950 61.950 268.050 62.550 ;
        RECT 266.100 58.050 267.900 59.850 ;
        RECT 271.950 58.050 273.150 71.400 ;
        RECT 277.950 60.450 282.000 61.050 ;
        RECT 277.950 58.950 282.450 60.450 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 274.950 55.950 277.050 58.050 ;
        RECT 269.100 54.150 270.900 55.950 ;
        RECT 272.850 51.750 274.050 55.950 ;
        RECT 275.100 54.150 276.900 55.950 ;
        RECT 281.550 55.050 282.450 58.950 ;
        RECT 290.400 57.900 291.600 71.400 ;
        RECT 311.400 57.900 312.600 71.400 ;
        RECT 329.850 58.050 331.050 71.400 ;
        RECT 334.500 65.400 336.300 78.000 ;
        RECT 339.150 65.400 340.950 77.400 ;
        RECT 342.150 71.400 343.950 78.000 ;
        RECT 347.550 71.400 349.350 77.400 ;
        RECT 352.350 71.400 354.150 78.000 ;
        RECT 347.550 70.500 348.750 71.400 ;
        RECT 355.350 70.500 357.150 77.400 ;
        RECT 358.950 71.400 360.750 78.000 ;
        RECT 363.150 71.400 364.950 77.400 ;
        RECT 367.650 74.400 369.450 78.000 ;
        RECT 343.950 68.400 348.750 70.500 ;
        RECT 351.450 69.450 358.050 70.500 ;
        RECT 351.450 68.700 353.250 69.450 ;
        RECT 356.250 68.700 358.050 69.450 ;
        RECT 363.150 69.300 367.050 71.400 ;
        RECT 347.550 67.500 348.750 68.400 ;
        RECT 360.450 67.800 362.250 68.400 ;
        RECT 347.550 66.300 355.050 67.500 ;
        RECT 353.250 65.700 355.050 66.300 ;
        RECT 355.950 66.900 362.250 67.800 ;
        RECT 339.150 64.500 340.050 65.400 ;
        RECT 355.950 64.800 356.850 66.900 ;
        RECT 360.450 66.600 362.250 66.900 ;
        RECT 363.150 66.600 365.850 68.400 ;
        RECT 363.150 65.700 364.050 66.600 ;
        RECT 348.450 64.500 356.850 64.800 ;
        RECT 339.150 63.900 356.850 64.500 ;
        RECT 358.950 64.800 364.050 65.700 ;
        RECT 364.950 64.800 367.050 65.700 ;
        RECT 370.650 65.400 372.450 77.400 ;
        RECT 380.400 71.400 382.200 78.000 ;
        RECT 383.400 71.400 385.200 77.400 ;
        RECT 386.400 72.000 388.200 78.000 ;
        RECT 383.700 71.100 385.200 71.400 ;
        RECT 389.400 71.400 391.200 77.400 ;
        RECT 401.400 71.400 403.200 78.000 ;
        RECT 404.400 71.400 406.200 77.400 ;
        RECT 407.400 71.400 409.200 78.000 ;
        RECT 421.800 71.400 423.600 77.400 ;
        RECT 424.800 71.400 426.600 78.000 ;
        RECT 389.400 71.100 390.300 71.400 ;
        RECT 383.700 70.200 390.300 71.100 ;
        RECT 339.150 63.300 350.250 63.900 ;
        RECT 335.100 58.050 336.900 59.850 ;
        RECT 286.950 55.800 289.050 57.900 ;
        RECT 289.950 55.800 292.050 57.900 ;
        RECT 292.950 55.800 295.050 57.900 ;
        RECT 307.950 55.800 310.050 57.900 ;
        RECT 310.950 55.800 313.050 57.900 ;
        RECT 313.950 55.800 316.050 57.900 ;
        RECT 325.950 55.950 328.050 58.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 277.950 53.550 282.450 55.050 ;
        RECT 287.100 54.000 288.900 55.800 ;
        RECT 277.950 52.950 282.000 53.550 ;
        RECT 272.850 50.700 276.600 51.750 ;
        RECT 250.950 46.500 253.050 48.600 ;
        RECT 241.200 45.600 242.250 46.500 ;
        RECT 250.950 45.600 252.000 46.500 ;
        RECT 227.850 42.000 229.650 45.600 ;
        RECT 232.650 42.600 234.450 45.600 ;
        RECT 236.850 42.000 238.650 45.600 ;
        RECT 240.450 42.600 242.250 45.600 ;
        RECT 243.750 42.000 245.550 45.600 ;
        RECT 248.250 44.700 252.000 45.600 ;
        RECT 248.250 42.600 250.050 44.700 ;
        RECT 253.050 42.000 254.850 45.600 ;
        RECT 256.050 42.600 257.850 48.600 ;
        RECT 266.400 47.700 274.200 49.050 ;
        RECT 266.400 42.600 268.200 47.700 ;
        RECT 269.400 42.000 271.200 46.800 ;
        RECT 272.400 42.600 274.200 47.700 ;
        RECT 275.400 48.600 276.600 50.700 ;
        RECT 290.400 50.700 291.600 55.800 ;
        RECT 293.100 54.000 294.900 55.800 ;
        RECT 308.100 54.000 309.900 55.800 ;
        RECT 311.400 50.700 312.600 55.800 ;
        RECT 314.100 54.000 315.900 55.800 ;
        RECT 326.100 54.150 327.900 55.950 ;
        RECT 290.400 49.800 294.600 50.700 ;
        RECT 275.400 42.600 277.200 48.600 ;
        RECT 287.700 42.000 289.500 48.600 ;
        RECT 292.800 42.600 294.600 49.800 ;
        RECT 308.400 49.800 312.600 50.700 ;
        RECT 313.950 51.450 316.050 52.050 ;
        RECT 319.950 51.450 322.050 52.050 ;
        RECT 328.950 51.750 330.150 55.950 ;
        RECT 332.100 54.150 333.900 55.950 ;
        RECT 313.950 50.550 322.050 51.450 ;
        RECT 313.950 49.950 316.050 50.550 ;
        RECT 319.950 49.950 322.050 50.550 ;
        RECT 326.400 50.700 330.150 51.750 ;
        RECT 308.400 42.600 310.200 49.800 ;
        RECT 326.400 48.600 327.600 50.700 ;
        RECT 313.500 42.000 315.300 48.600 ;
        RECT 325.800 42.600 327.600 48.600 ;
        RECT 328.800 47.700 336.600 49.050 ;
        RECT 328.800 42.600 330.600 47.700 ;
        RECT 331.800 42.000 333.600 46.800 ;
        RECT 334.800 42.600 336.600 47.700 ;
        RECT 339.150 48.600 340.050 63.300 ;
        RECT 348.450 63.000 350.250 63.300 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 349.950 56.400 352.050 58.050 ;
        RECT 341.100 54.150 342.900 55.950 ;
        RECT 344.100 55.200 352.050 56.400 ;
        RECT 344.100 54.600 345.900 55.200 ;
        RECT 342.000 53.400 342.900 54.150 ;
        RECT 347.100 53.400 348.900 54.000 ;
        RECT 342.000 52.200 348.900 53.400 ;
        RECT 358.950 52.200 359.850 64.800 ;
        RECT 364.950 63.600 369.150 64.800 ;
        RECT 368.250 61.800 370.050 63.600 ;
        RECT 371.250 58.050 372.450 65.400 ;
        RECT 367.950 57.750 372.450 58.050 ;
        RECT 383.100 57.900 384.900 59.700 ;
        RECT 389.400 57.900 390.300 70.200 ;
        RECT 400.950 60.450 403.050 61.050 ;
        RECT 395.550 59.550 403.050 60.450 ;
        RECT 366.150 55.950 372.450 57.750 ;
        RECT 347.850 51.000 359.850 52.200 ;
        RECT 347.850 49.200 348.900 51.000 ;
        RECT 358.050 50.400 359.850 51.000 ;
        RECT 339.150 42.600 340.950 48.600 ;
        RECT 343.950 46.500 346.050 48.600 ;
        RECT 347.550 47.400 349.350 49.200 ;
        RECT 371.250 48.600 372.450 55.950 ;
        RECT 379.950 55.800 382.050 57.900 ;
        RECT 382.950 55.800 385.050 57.900 ;
        RECT 385.950 55.800 388.050 57.900 ;
        RECT 388.950 55.800 391.050 57.900 ;
        RECT 380.100 54.000 381.900 55.800 ;
        RECT 386.100 54.000 387.900 55.800 ;
        RECT 389.400 52.200 390.300 55.800 ;
        RECT 395.550 55.050 396.450 59.550 ;
        RECT 400.950 58.950 403.050 59.550 ;
        RECT 404.400 57.900 405.600 71.400 ;
        RECT 415.950 61.950 418.050 64.050 ;
        RECT 406.950 60.450 409.050 61.050 ;
        RECT 412.950 60.450 415.050 61.050 ;
        RECT 406.950 59.550 415.050 60.450 ;
        RECT 406.950 58.950 409.050 59.550 ;
        RECT 412.950 58.950 415.050 59.550 ;
        RECT 400.950 55.800 403.050 57.900 ;
        RECT 403.950 55.800 406.050 57.900 ;
        RECT 406.950 55.800 409.050 57.900 ;
        RECT 391.950 53.550 396.450 55.050 ;
        RECT 401.100 54.000 402.900 55.800 ;
        RECT 391.950 52.950 396.000 53.550 ;
        RECT 350.850 47.550 352.650 48.300 ;
        RECT 364.950 47.700 367.050 48.600 ;
        RECT 350.850 46.500 355.800 47.550 ;
        RECT 345.000 45.600 346.050 46.500 ;
        RECT 354.750 45.600 355.800 46.500 ;
        RECT 363.300 46.500 367.050 47.700 ;
        RECT 363.300 45.600 364.350 46.500 ;
        RECT 342.150 42.000 343.950 45.600 ;
        RECT 345.000 44.700 348.750 45.600 ;
        RECT 346.950 42.600 348.750 44.700 ;
        RECT 351.450 42.000 353.250 45.600 ;
        RECT 354.750 42.600 356.550 45.600 ;
        RECT 358.350 42.000 360.150 45.600 ;
        RECT 362.550 42.600 364.350 45.600 ;
        RECT 367.350 42.000 369.150 45.600 ;
        RECT 370.650 42.600 372.450 48.600 ;
        RECT 380.400 42.000 382.200 51.600 ;
        RECT 387.000 51.000 390.300 52.200 ;
        RECT 387.000 42.600 388.800 51.000 ;
        RECT 404.400 50.700 405.600 55.800 ;
        RECT 407.100 54.000 408.900 55.800 ;
        RECT 409.950 54.450 412.050 55.050 ;
        RECT 416.550 54.450 417.450 61.950 ;
        RECT 422.400 58.050 423.600 71.400 ;
        RECT 434.400 65.400 436.200 78.000 ;
        RECT 439.500 66.600 441.300 77.400 ;
        RECT 437.700 65.400 441.300 66.600 ;
        RECT 456.300 65.400 458.100 78.000 ;
        RECT 460.800 65.400 464.100 77.400 ;
        RECT 466.800 65.400 468.600 78.000 ;
        RECT 476.400 71.400 478.200 78.000 ;
        RECT 479.400 71.400 481.200 77.400 ;
        RECT 425.100 58.050 426.900 59.850 ;
        RECT 434.100 58.050 435.900 59.850 ;
        RECT 437.700 58.050 438.600 65.400 ;
        RECT 440.100 58.050 441.900 59.850 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 455.100 57.900 456.900 59.700 ;
        RECT 461.700 57.900 462.900 65.400 ;
        RECT 467.100 57.900 468.900 59.700 ;
        RECT 476.100 58.050 477.900 59.850 ;
        RECT 479.400 58.050 480.600 71.400 ;
        RECT 493.800 65.400 495.600 77.400 ;
        RECT 496.800 71.400 498.600 78.000 ;
        RECT 499.800 71.400 501.600 77.400 ;
        RECT 511.800 71.400 513.600 77.400 ;
        RECT 514.800 71.400 516.600 78.000 ;
        RECT 493.800 58.050 495.000 65.400 ;
        RECT 500.400 64.500 501.600 71.400 ;
        RECT 495.900 63.600 501.600 64.500 ;
        RECT 495.900 62.700 497.850 63.600 ;
        RECT 409.950 53.550 417.450 54.450 ;
        RECT 409.950 52.950 412.050 53.550 ;
        RECT 404.400 49.800 408.600 50.700 ;
        RECT 401.700 42.000 403.500 48.600 ;
        RECT 406.800 42.600 408.600 49.800 ;
        RECT 422.400 45.600 423.600 55.950 ;
        RECT 424.950 51.450 427.050 52.050 ;
        RECT 433.950 51.450 436.050 52.050 ;
        RECT 424.950 50.550 436.050 51.450 ;
        RECT 424.950 49.950 427.050 50.550 ;
        RECT 433.950 49.950 436.050 50.550 ;
        RECT 437.700 45.600 438.600 55.950 ;
        RECT 454.950 55.800 457.050 57.900 ;
        RECT 457.950 55.800 460.050 57.900 ;
        RECT 460.950 55.800 463.050 57.900 ;
        RECT 463.950 55.800 466.050 57.900 ;
        RECT 466.950 55.800 469.050 57.900 ;
        RECT 475.950 55.950 478.050 58.050 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 493.800 55.950 496.050 58.050 ;
        RECT 458.100 54.000 459.900 55.800 ;
        RECT 462.000 53.400 463.050 55.800 ;
        RECT 464.100 54.000 465.900 55.800 ;
        RECT 461.700 51.300 462.900 53.400 ;
        RECT 458.400 50.100 462.900 51.300 ;
        RECT 442.950 48.450 445.050 49.050 ;
        RECT 448.950 48.450 451.050 49.050 ;
        RECT 458.400 48.600 459.300 50.100 ;
        RECT 442.950 47.550 451.050 48.450 ;
        RECT 442.950 46.950 445.050 47.550 ;
        RECT 448.950 46.950 451.050 47.550 ;
        RECT 421.800 42.600 423.600 45.600 ;
        RECT 424.800 42.000 426.600 45.600 ;
        RECT 434.400 42.000 436.200 45.600 ;
        RECT 437.400 42.600 439.200 45.600 ;
        RECT 440.400 42.000 442.200 45.600 ;
        RECT 454.800 43.500 456.600 48.600 ;
        RECT 457.800 44.400 459.600 48.600 ;
        RECT 460.800 48.000 468.600 48.900 ;
        RECT 460.800 43.500 462.600 48.000 ;
        RECT 454.800 42.600 462.600 43.500 ;
        RECT 463.800 42.000 465.600 47.100 ;
        RECT 466.800 42.600 468.600 48.000 ;
        RECT 479.400 45.600 480.600 55.950 ;
        RECT 493.800 48.600 495.000 55.950 ;
        RECT 496.950 51.300 497.850 62.700 ;
        RECT 500.100 58.050 501.900 59.850 ;
        RECT 512.400 58.050 513.600 71.400 ;
        RECT 524.700 65.400 526.500 78.000 ;
        RECT 529.800 71.400 531.600 77.400 ;
        RECT 532.800 71.400 534.600 78.000 ;
        RECT 547.800 71.400 549.600 78.000 ;
        RECT 550.800 71.400 552.600 77.400 ;
        RECT 553.800 71.400 555.600 78.000 ;
        RECT 515.100 58.050 516.900 59.850 ;
        RECT 524.100 58.050 525.900 59.850 ;
        RECT 529.950 58.050 531.150 71.400 ;
        RECT 532.950 63.450 535.050 64.050 ;
        RECT 538.950 63.450 541.050 64.050 ;
        RECT 532.950 62.550 541.050 63.450 ;
        RECT 532.950 61.950 535.050 62.550 ;
        RECT 538.950 61.950 541.050 62.550 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 514.950 55.950 517.050 58.050 ;
        RECT 523.950 55.950 526.050 58.050 ;
        RECT 526.950 55.950 529.050 58.050 ;
        RECT 529.950 55.950 532.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 551.400 57.900 552.600 71.400 ;
        RECT 558.150 65.400 559.950 77.400 ;
        RECT 561.150 71.400 562.950 78.000 ;
        RECT 566.550 71.400 568.350 77.400 ;
        RECT 571.350 71.400 573.150 78.000 ;
        RECT 566.550 70.500 567.750 71.400 ;
        RECT 574.350 70.500 576.150 77.400 ;
        RECT 577.950 71.400 579.750 78.000 ;
        RECT 582.150 71.400 583.950 77.400 ;
        RECT 586.650 74.400 588.450 78.000 ;
        RECT 562.950 68.400 567.750 70.500 ;
        RECT 570.450 69.450 577.050 70.500 ;
        RECT 570.450 68.700 572.250 69.450 ;
        RECT 575.250 68.700 577.050 69.450 ;
        RECT 582.150 69.300 586.050 71.400 ;
        RECT 566.550 67.500 567.750 68.400 ;
        RECT 579.450 67.800 581.250 68.400 ;
        RECT 566.550 66.300 574.050 67.500 ;
        RECT 572.250 65.700 574.050 66.300 ;
        RECT 574.950 66.900 581.250 67.800 ;
        RECT 558.150 64.500 559.050 65.400 ;
        RECT 574.950 64.800 575.850 66.900 ;
        RECT 579.450 66.600 581.250 66.900 ;
        RECT 582.150 66.600 584.850 68.400 ;
        RECT 582.150 65.700 583.050 66.600 ;
        RECT 567.450 64.500 575.850 64.800 ;
        RECT 558.150 63.900 575.850 64.500 ;
        RECT 577.950 64.800 583.050 65.700 ;
        RECT 583.950 64.800 586.050 65.700 ;
        RECT 589.650 65.400 591.450 77.400 ;
        RECT 599.400 71.400 601.200 78.000 ;
        RECT 602.400 71.400 604.200 77.400 ;
        RECT 605.400 71.400 607.200 78.000 ;
        RECT 619.800 71.400 621.600 78.000 ;
        RECT 622.800 71.400 624.600 77.400 ;
        RECT 625.800 71.400 627.600 78.000 ;
        RECT 558.150 63.300 569.250 63.900 ;
        RECT 495.900 50.400 497.850 51.300 ;
        RECT 495.900 49.500 501.600 50.400 ;
        RECT 476.400 42.000 478.200 45.600 ;
        RECT 479.400 42.600 481.200 45.600 ;
        RECT 493.800 42.600 495.600 48.600 ;
        RECT 500.400 45.600 501.600 49.500 ;
        RECT 512.400 45.600 513.600 55.950 ;
        RECT 527.100 54.150 528.900 55.950 ;
        RECT 530.850 51.750 532.050 55.950 ;
        RECT 533.100 54.150 534.900 55.950 ;
        RECT 547.950 55.800 550.050 57.900 ;
        RECT 550.950 55.800 553.050 57.900 ;
        RECT 553.950 55.800 556.050 57.900 ;
        RECT 548.100 54.000 549.900 55.800 ;
        RECT 530.850 50.700 534.600 51.750 ;
        RECT 551.400 50.700 552.600 55.800 ;
        RECT 554.100 54.000 555.900 55.800 ;
        RECT 524.400 47.700 532.200 49.050 ;
        RECT 496.800 42.000 498.600 45.600 ;
        RECT 499.800 42.600 501.600 45.600 ;
        RECT 511.800 42.600 513.600 45.600 ;
        RECT 514.800 42.000 516.600 45.600 ;
        RECT 524.400 42.600 526.200 47.700 ;
        RECT 527.400 42.000 529.200 46.800 ;
        RECT 530.400 42.600 532.200 47.700 ;
        RECT 533.400 48.600 534.600 50.700 ;
        RECT 548.400 49.800 552.600 50.700 ;
        RECT 533.400 42.600 535.200 48.600 ;
        RECT 548.400 42.600 550.200 49.800 ;
        RECT 558.150 48.600 559.050 63.300 ;
        RECT 567.450 63.000 569.250 63.300 ;
        RECT 559.950 55.950 562.050 58.050 ;
        RECT 568.950 56.400 571.050 58.050 ;
        RECT 560.100 54.150 561.900 55.950 ;
        RECT 563.100 55.200 571.050 56.400 ;
        RECT 563.100 54.600 564.900 55.200 ;
        RECT 561.000 53.400 561.900 54.150 ;
        RECT 566.100 53.400 567.900 54.000 ;
        RECT 561.000 52.200 567.900 53.400 ;
        RECT 577.950 52.200 578.850 64.800 ;
        RECT 583.950 63.600 588.150 64.800 ;
        RECT 587.250 61.800 589.050 63.600 ;
        RECT 590.250 58.050 591.450 65.400 ;
        RECT 586.950 57.750 591.450 58.050 ;
        RECT 602.400 57.900 603.600 71.400 ;
        RECT 623.400 57.900 624.600 71.400 ;
        RECT 638.700 66.600 640.500 77.400 ;
        RECT 638.700 65.400 642.300 66.600 ;
        RECT 643.800 65.400 645.600 78.000 ;
        RECT 653.400 71.400 655.200 77.400 ;
        RECT 656.400 71.400 658.200 78.000 ;
        RECT 638.100 58.050 639.900 59.850 ;
        RECT 641.400 58.050 642.300 65.400 ;
        RECT 653.400 64.500 654.600 71.400 ;
        RECT 659.400 65.400 661.200 77.400 ;
        RECT 671.400 65.400 673.200 78.000 ;
        RECT 676.500 66.600 678.300 77.400 ;
        RECT 674.700 65.400 678.300 66.600 ;
        RECT 689.400 65.400 691.200 78.000 ;
        RECT 694.500 66.600 696.300 77.400 ;
        RECT 692.700 65.400 696.300 66.600 ;
        RECT 709.800 65.400 711.600 77.400 ;
        RECT 712.800 66.300 714.600 77.400 ;
        RECT 715.800 67.200 717.600 78.000 ;
        RECT 718.800 66.300 720.600 77.400 ;
        RECT 728.400 71.400 730.200 78.000 ;
        RECT 731.400 71.400 733.200 77.400 ;
        RECT 743.400 71.400 745.200 78.000 ;
        RECT 746.400 71.400 748.200 77.400 ;
        RECT 749.400 71.400 751.200 78.000 ;
        RECT 712.800 65.400 720.600 66.300 ;
        RECT 653.400 63.600 659.100 64.500 ;
        RECT 657.150 62.700 659.100 63.600 ;
        RECT 644.100 58.050 645.900 59.850 ;
        RECT 653.100 58.050 654.900 59.850 ;
        RECT 585.150 55.950 591.450 57.750 ;
        RECT 566.850 51.000 578.850 52.200 ;
        RECT 566.850 49.200 567.900 51.000 ;
        RECT 577.050 50.400 578.850 51.000 ;
        RECT 553.500 42.000 555.300 48.600 ;
        RECT 558.150 42.600 559.950 48.600 ;
        RECT 562.950 46.500 565.050 48.600 ;
        RECT 566.550 47.400 568.350 49.200 ;
        RECT 590.250 48.600 591.450 55.950 ;
        RECT 598.950 55.800 601.050 57.900 ;
        RECT 601.950 55.800 604.050 57.900 ;
        RECT 604.950 55.800 607.050 57.900 ;
        RECT 619.950 55.800 622.050 57.900 ;
        RECT 622.950 55.800 625.050 57.900 ;
        RECT 625.950 55.800 628.050 57.900 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 652.950 55.950 655.050 58.050 ;
        RECT 599.100 54.000 600.900 55.800 ;
        RECT 602.400 50.700 603.600 55.800 ;
        RECT 605.100 54.000 606.900 55.800 ;
        RECT 620.100 54.000 621.900 55.800 ;
        RECT 623.400 50.700 624.600 55.800 ;
        RECT 626.100 54.000 627.900 55.800 ;
        RECT 602.400 49.800 606.600 50.700 ;
        RECT 569.850 47.550 571.650 48.300 ;
        RECT 583.950 47.700 586.050 48.600 ;
        RECT 569.850 46.500 574.800 47.550 ;
        RECT 564.000 45.600 565.050 46.500 ;
        RECT 573.750 45.600 574.800 46.500 ;
        RECT 582.300 46.500 586.050 47.700 ;
        RECT 582.300 45.600 583.350 46.500 ;
        RECT 561.150 42.000 562.950 45.600 ;
        RECT 564.000 44.700 567.750 45.600 ;
        RECT 565.950 42.600 567.750 44.700 ;
        RECT 570.450 42.000 572.250 45.600 ;
        RECT 573.750 42.600 575.550 45.600 ;
        RECT 577.350 42.000 579.150 45.600 ;
        RECT 581.550 42.600 583.350 45.600 ;
        RECT 586.350 42.000 588.150 45.600 ;
        RECT 589.650 42.600 591.450 48.600 ;
        RECT 599.700 42.000 601.500 48.600 ;
        RECT 604.800 42.600 606.600 49.800 ;
        RECT 620.400 49.800 624.600 50.700 ;
        RECT 620.400 42.600 622.200 49.800 ;
        RECT 625.500 42.000 627.300 48.600 ;
        RECT 641.400 45.600 642.300 55.950 ;
        RECT 657.150 51.300 658.050 62.700 ;
        RECT 660.000 58.050 661.200 65.400 ;
        RECT 671.100 58.050 672.900 59.850 ;
        RECT 674.700 58.050 675.600 65.400 ;
        RECT 676.950 63.450 679.050 64.050 ;
        RECT 685.950 63.450 688.050 64.050 ;
        RECT 676.950 62.550 688.050 63.450 ;
        RECT 676.950 61.950 679.050 62.550 ;
        RECT 685.950 61.950 688.050 62.550 ;
        RECT 677.100 58.050 678.900 59.850 ;
        RECT 689.100 58.050 690.900 59.850 ;
        RECT 692.700 58.050 693.600 65.400 ;
        RECT 695.100 58.050 696.900 59.850 ;
        RECT 658.950 55.950 661.200 58.050 ;
        RECT 670.950 55.950 673.050 58.050 ;
        RECT 673.950 55.950 676.050 58.050 ;
        RECT 676.950 55.950 679.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 691.950 55.950 694.050 58.050 ;
        RECT 694.950 55.950 697.050 58.050 ;
        RECT 710.400 57.900 711.300 65.400 ;
        RECT 716.100 57.900 717.900 59.700 ;
        RECT 728.100 58.050 729.900 59.850 ;
        RECT 731.400 58.050 732.600 71.400 ;
        RECT 657.150 50.400 659.100 51.300 ;
        RECT 653.400 49.500 659.100 50.400 ;
        RECT 653.400 45.600 654.600 49.500 ;
        RECT 660.000 48.600 661.200 55.950 ;
        RECT 637.800 42.000 639.600 45.600 ;
        RECT 640.800 42.600 642.600 45.600 ;
        RECT 643.800 42.000 645.600 45.600 ;
        RECT 653.400 42.600 655.200 45.600 ;
        RECT 656.400 42.000 658.200 45.600 ;
        RECT 659.400 42.600 661.200 48.600 ;
        RECT 674.700 45.600 675.600 55.950 ;
        RECT 692.700 45.600 693.600 55.950 ;
        RECT 709.950 55.800 712.050 57.900 ;
        RECT 712.950 55.800 715.050 57.900 ;
        RECT 715.950 55.800 718.050 57.900 ;
        RECT 718.950 55.800 721.050 57.900 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 730.950 55.950 733.050 58.050 ;
        RECT 710.400 48.600 711.300 55.800 ;
        RECT 713.100 54.000 714.900 55.800 ;
        RECT 719.100 54.000 720.900 55.800 ;
        RECT 710.400 47.400 715.500 48.600 ;
        RECT 671.400 42.000 673.200 45.600 ;
        RECT 674.400 42.600 676.200 45.600 ;
        RECT 677.400 42.000 679.200 45.600 ;
        RECT 689.400 42.000 691.200 45.600 ;
        RECT 692.400 42.600 694.200 45.600 ;
        RECT 695.400 42.000 697.200 45.600 ;
        RECT 710.700 42.000 712.500 45.600 ;
        RECT 713.700 42.600 715.500 47.400 ;
        RECT 718.200 42.000 720.000 48.600 ;
        RECT 731.400 45.600 732.600 55.950 ;
        RECT 742.950 55.800 745.050 57.900 ;
        RECT 743.100 54.000 744.900 55.800 ;
        RECT 746.400 51.300 747.300 71.400 ;
        RECT 752.400 65.400 754.200 77.400 ;
        RECT 764.400 71.400 766.200 78.000 ;
        RECT 767.400 71.400 769.200 77.400 ;
        RECT 781.800 71.400 783.600 77.400 ;
        RECT 784.800 71.400 786.600 78.000 ;
        RECT 749.100 57.900 750.900 59.700 ;
        RECT 752.700 57.900 753.600 65.400 ;
        RECT 764.100 58.050 765.900 59.850 ;
        RECT 767.400 58.050 768.600 71.400 ;
        RECT 782.400 58.050 783.600 71.400 ;
        RECT 789.150 65.400 790.950 77.400 ;
        RECT 792.150 71.400 793.950 78.000 ;
        RECT 797.550 71.400 799.350 77.400 ;
        RECT 802.350 71.400 804.150 78.000 ;
        RECT 797.550 70.500 798.750 71.400 ;
        RECT 805.350 70.500 807.150 77.400 ;
        RECT 808.950 71.400 810.750 78.000 ;
        RECT 813.150 71.400 814.950 77.400 ;
        RECT 817.650 74.400 819.450 78.000 ;
        RECT 793.950 68.400 798.750 70.500 ;
        RECT 801.450 69.450 808.050 70.500 ;
        RECT 801.450 68.700 803.250 69.450 ;
        RECT 806.250 68.700 808.050 69.450 ;
        RECT 813.150 69.300 817.050 71.400 ;
        RECT 797.550 67.500 798.750 68.400 ;
        RECT 810.450 67.800 812.250 68.400 ;
        RECT 797.550 66.300 805.050 67.500 ;
        RECT 803.250 65.700 805.050 66.300 ;
        RECT 805.950 66.900 812.250 67.800 ;
        RECT 789.150 64.500 790.050 65.400 ;
        RECT 805.950 64.800 806.850 66.900 ;
        RECT 810.450 66.600 812.250 66.900 ;
        RECT 813.150 66.600 815.850 68.400 ;
        RECT 813.150 65.700 814.050 66.600 ;
        RECT 798.450 64.500 806.850 64.800 ;
        RECT 789.150 63.900 806.850 64.500 ;
        RECT 808.950 64.800 814.050 65.700 ;
        RECT 814.950 64.800 817.050 65.700 ;
        RECT 820.650 65.400 822.450 77.400 ;
        RECT 830.400 71.400 832.200 78.000 ;
        RECT 833.400 71.400 835.200 77.400 ;
        RECT 789.150 63.300 800.250 63.900 ;
        RECT 785.100 58.050 786.900 59.850 ;
        RECT 748.950 55.800 751.050 57.900 ;
        RECT 751.950 55.800 754.050 57.900 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 743.400 50.400 750.900 51.300 ;
        RECT 728.400 42.000 730.200 45.600 ;
        RECT 731.400 42.600 733.200 45.600 ;
        RECT 743.400 42.600 745.200 50.400 ;
        RECT 749.100 49.500 750.900 50.400 ;
        RECT 752.700 48.600 753.600 55.800 ;
        RECT 747.900 42.000 749.700 48.600 ;
        RECT 750.900 46.800 753.600 48.600 ;
        RECT 750.900 42.600 752.700 46.800 ;
        RECT 767.400 45.600 768.600 55.950 ;
        RECT 782.400 45.600 783.600 55.950 ;
        RECT 789.150 48.600 790.050 63.300 ;
        RECT 798.450 63.000 800.250 63.300 ;
        RECT 790.950 55.950 793.050 58.050 ;
        RECT 799.950 56.400 802.050 58.050 ;
        RECT 791.100 54.150 792.900 55.950 ;
        RECT 794.100 55.200 802.050 56.400 ;
        RECT 794.100 54.600 795.900 55.200 ;
        RECT 792.000 53.400 792.900 54.150 ;
        RECT 797.100 53.400 798.900 54.000 ;
        RECT 792.000 52.200 798.900 53.400 ;
        RECT 808.950 52.200 809.850 64.800 ;
        RECT 814.950 63.600 819.150 64.800 ;
        RECT 818.250 61.800 820.050 63.600 ;
        RECT 821.250 58.050 822.450 65.400 ;
        RECT 830.100 58.050 831.900 59.850 ;
        RECT 833.400 58.050 834.600 71.400 ;
        RECT 845.400 65.400 847.200 78.000 ;
        RECT 850.500 66.600 852.300 77.400 ;
        RECT 848.700 65.400 852.300 66.600 ;
        RECT 845.100 58.050 846.900 59.850 ;
        RECT 848.700 58.050 849.600 65.400 ;
        RECT 851.100 58.050 852.900 59.850 ;
        RECT 817.950 57.750 822.450 58.050 ;
        RECT 816.150 55.950 822.450 57.750 ;
        RECT 829.950 55.950 832.050 58.050 ;
        RECT 832.950 55.950 835.050 58.050 ;
        RECT 844.950 55.950 847.050 58.050 ;
        RECT 847.950 55.950 850.050 58.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 797.850 51.000 809.850 52.200 ;
        RECT 797.850 49.200 798.900 51.000 ;
        RECT 808.050 50.400 809.850 51.000 ;
        RECT 764.400 42.000 766.200 45.600 ;
        RECT 767.400 42.600 769.200 45.600 ;
        RECT 781.800 42.600 783.600 45.600 ;
        RECT 784.800 42.000 786.600 45.600 ;
        RECT 789.150 42.600 790.950 48.600 ;
        RECT 793.950 46.500 796.050 48.600 ;
        RECT 797.550 47.400 799.350 49.200 ;
        RECT 821.250 48.600 822.450 55.950 ;
        RECT 800.850 47.550 802.650 48.300 ;
        RECT 814.950 47.700 817.050 48.600 ;
        RECT 800.850 46.500 805.800 47.550 ;
        RECT 795.000 45.600 796.050 46.500 ;
        RECT 804.750 45.600 805.800 46.500 ;
        RECT 813.300 46.500 817.050 47.700 ;
        RECT 813.300 45.600 814.350 46.500 ;
        RECT 792.150 42.000 793.950 45.600 ;
        RECT 795.000 44.700 798.750 45.600 ;
        RECT 796.950 42.600 798.750 44.700 ;
        RECT 801.450 42.000 803.250 45.600 ;
        RECT 804.750 42.600 806.550 45.600 ;
        RECT 808.350 42.000 810.150 45.600 ;
        RECT 812.550 42.600 814.350 45.600 ;
        RECT 817.350 42.000 819.150 45.600 ;
        RECT 820.650 42.600 822.450 48.600 ;
        RECT 833.400 45.600 834.600 55.950 ;
        RECT 848.700 45.600 849.600 55.950 ;
        RECT 830.400 42.000 832.200 45.600 ;
        RECT 833.400 42.600 835.200 45.600 ;
        RECT 845.400 42.000 847.200 45.600 ;
        RECT 848.400 42.600 850.200 45.600 ;
        RECT 851.400 42.000 853.200 45.600 ;
        RECT 10.800 35.400 12.600 38.400 ;
        RECT 13.800 35.400 15.600 39.000 ;
        RECT 11.400 25.050 12.600 35.400 ;
        RECT 17.550 32.400 19.350 38.400 ;
        RECT 20.850 35.400 22.650 39.000 ;
        RECT 25.650 35.400 27.450 38.400 ;
        RECT 29.850 35.400 31.650 39.000 ;
        RECT 33.450 35.400 35.250 38.400 ;
        RECT 36.750 35.400 38.550 39.000 ;
        RECT 41.250 36.300 43.050 38.400 ;
        RECT 41.250 35.400 45.000 36.300 ;
        RECT 46.050 35.400 47.850 39.000 ;
        RECT 25.650 34.500 26.700 35.400 ;
        RECT 22.950 33.300 26.700 34.500 ;
        RECT 34.200 34.500 35.250 35.400 ;
        RECT 43.950 34.500 45.000 35.400 ;
        RECT 34.200 33.450 39.150 34.500 ;
        RECT 22.950 32.400 25.050 33.300 ;
        RECT 37.350 32.700 39.150 33.450 ;
        RECT 17.550 25.050 18.750 32.400 ;
        RECT 40.650 31.800 42.450 33.600 ;
        RECT 43.950 32.400 46.050 34.500 ;
        RECT 49.050 32.400 50.850 38.400 ;
        RECT 30.150 30.000 31.950 30.600 ;
        RECT 41.100 30.000 42.150 31.800 ;
        RECT 30.150 28.800 42.150 30.000 ;
        RECT 10.950 22.950 13.050 25.050 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 17.550 23.250 23.850 25.050 ;
        RECT 17.550 22.950 22.050 23.250 ;
        RECT 11.400 9.600 12.600 22.950 ;
        RECT 14.100 21.150 15.900 22.950 ;
        RECT 17.550 15.600 18.750 22.950 ;
        RECT 19.950 17.400 21.750 19.200 ;
        RECT 20.850 16.200 25.050 17.400 ;
        RECT 30.150 16.200 31.050 28.800 ;
        RECT 41.100 27.600 48.000 28.800 ;
        RECT 41.100 27.000 42.900 27.600 ;
        RECT 47.100 26.850 48.000 27.600 ;
        RECT 44.100 25.800 45.900 26.400 ;
        RECT 37.950 24.600 45.900 25.800 ;
        RECT 47.100 25.050 48.900 26.850 ;
        RECT 37.950 22.950 40.050 24.600 ;
        RECT 46.950 22.950 49.050 25.050 ;
        RECT 39.750 17.700 41.550 18.000 ;
        RECT 49.950 17.700 50.850 32.400 ;
        RECT 59.400 33.300 61.200 38.400 ;
        RECT 62.400 34.200 64.200 39.000 ;
        RECT 65.400 33.300 67.200 38.400 ;
        RECT 59.400 31.950 67.200 33.300 ;
        RECT 68.400 32.400 70.200 38.400 ;
        RECT 80.700 32.400 82.500 39.000 ;
        RECT 68.400 30.300 69.600 32.400 ;
        RECT 85.800 31.200 87.600 38.400 ;
        RECT 65.850 29.250 69.600 30.300 ;
        RECT 83.400 30.300 87.600 31.200 ;
        RECT 92.550 32.400 94.350 38.400 ;
        RECT 95.850 35.400 97.650 39.000 ;
        RECT 100.650 35.400 102.450 38.400 ;
        RECT 104.850 35.400 106.650 39.000 ;
        RECT 108.450 35.400 110.250 38.400 ;
        RECT 111.750 35.400 113.550 39.000 ;
        RECT 116.250 36.300 118.050 38.400 ;
        RECT 116.250 35.400 120.000 36.300 ;
        RECT 121.050 35.400 122.850 39.000 ;
        RECT 100.650 34.500 101.700 35.400 ;
        RECT 97.950 33.300 101.700 34.500 ;
        RECT 109.200 34.500 110.250 35.400 ;
        RECT 118.950 34.500 120.000 35.400 ;
        RECT 109.200 33.450 114.150 34.500 ;
        RECT 97.950 32.400 100.050 33.300 ;
        RECT 112.350 32.700 114.150 33.450 ;
        RECT 62.100 25.050 63.900 26.850 ;
        RECT 65.850 25.050 67.050 29.250 ;
        RECT 68.100 25.050 69.900 26.850 ;
        RECT 80.100 25.200 81.900 27.000 ;
        RECT 83.400 25.200 84.600 30.300 ;
        RECT 86.100 25.200 87.900 27.000 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 64.950 22.950 67.050 25.050 ;
        RECT 67.950 22.950 70.050 25.050 ;
        RECT 79.950 23.100 82.050 25.200 ;
        RECT 82.950 23.100 85.050 25.200 ;
        RECT 85.950 23.100 88.050 25.200 ;
        RECT 92.550 25.050 93.750 32.400 ;
        RECT 115.650 31.800 117.450 33.600 ;
        RECT 118.950 32.400 121.050 34.500 ;
        RECT 124.050 32.400 125.850 38.400 ;
        RECT 136.800 35.400 138.600 39.000 ;
        RECT 139.800 35.400 141.600 38.400 ;
        RECT 142.800 35.400 144.600 39.000 ;
        RECT 155.700 35.400 157.500 39.000 ;
        RECT 105.150 30.000 106.950 30.600 ;
        RECT 116.100 30.000 117.150 31.800 ;
        RECT 105.150 28.800 117.150 30.000 ;
        RECT 92.550 23.250 98.850 25.050 ;
        RECT 59.100 21.150 60.900 22.950 ;
        RECT 39.750 17.100 50.850 17.700 ;
        RECT 10.800 3.600 12.600 9.600 ;
        RECT 13.800 3.000 15.600 9.600 ;
        RECT 17.550 3.600 19.350 15.600 ;
        RECT 22.950 15.300 25.050 16.200 ;
        RECT 25.950 15.300 31.050 16.200 ;
        RECT 33.150 16.500 50.850 17.100 ;
        RECT 33.150 16.200 41.550 16.500 ;
        RECT 25.950 14.400 26.850 15.300 ;
        RECT 24.150 12.600 26.850 14.400 ;
        RECT 27.750 14.100 29.550 14.400 ;
        RECT 33.150 14.100 34.050 16.200 ;
        RECT 49.950 15.600 50.850 16.500 ;
        RECT 27.750 13.200 34.050 14.100 ;
        RECT 34.950 14.700 36.750 15.300 ;
        RECT 34.950 13.500 42.450 14.700 ;
        RECT 27.750 12.600 29.550 13.200 ;
        RECT 41.250 12.600 42.450 13.500 ;
        RECT 22.950 9.600 26.850 11.700 ;
        RECT 31.950 11.550 33.750 12.300 ;
        RECT 36.750 11.550 38.550 12.300 ;
        RECT 31.950 10.500 38.550 11.550 ;
        RECT 41.250 10.500 46.050 12.600 ;
        RECT 20.550 3.000 22.350 6.600 ;
        RECT 25.050 3.600 26.850 9.600 ;
        RECT 29.250 3.000 31.050 9.600 ;
        RECT 32.850 3.600 34.650 10.500 ;
        RECT 41.250 9.600 42.450 10.500 ;
        RECT 35.850 3.000 37.650 9.600 ;
        RECT 40.650 3.600 42.450 9.600 ;
        RECT 46.050 3.000 47.850 9.600 ;
        RECT 49.050 3.600 50.850 15.600 ;
        RECT 59.700 3.000 61.500 15.600 ;
        RECT 64.950 9.600 66.150 22.950 ;
        RECT 83.400 9.600 84.600 23.100 ;
        RECT 92.550 22.950 97.050 23.250 ;
        RECT 92.550 15.600 93.750 22.950 ;
        RECT 94.950 17.400 96.750 19.200 ;
        RECT 95.850 16.200 100.050 17.400 ;
        RECT 105.150 16.200 106.050 28.800 ;
        RECT 116.100 27.600 123.000 28.800 ;
        RECT 116.100 27.000 117.900 27.600 ;
        RECT 122.100 26.850 123.000 27.600 ;
        RECT 119.100 25.800 120.900 26.400 ;
        RECT 112.950 24.600 120.900 25.800 ;
        RECT 122.100 25.050 123.900 26.850 ;
        RECT 112.950 22.950 115.050 24.600 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 114.750 17.700 116.550 18.000 ;
        RECT 124.950 17.700 125.850 32.400 ;
        RECT 140.400 25.050 141.300 35.400 ;
        RECT 158.700 33.600 160.500 38.400 ;
        RECT 155.400 32.400 160.500 33.600 ;
        RECT 163.200 32.400 165.000 39.000 ;
        RECT 168.150 32.400 169.950 38.400 ;
        RECT 171.150 35.400 172.950 39.000 ;
        RECT 175.950 36.300 177.750 38.400 ;
        RECT 174.000 35.400 177.750 36.300 ;
        RECT 180.450 35.400 182.250 39.000 ;
        RECT 183.750 35.400 185.550 38.400 ;
        RECT 187.350 35.400 189.150 39.000 ;
        RECT 191.550 35.400 193.350 38.400 ;
        RECT 196.350 35.400 198.150 39.000 ;
        RECT 174.000 34.500 175.050 35.400 ;
        RECT 183.750 34.500 184.800 35.400 ;
        RECT 172.950 32.400 175.050 34.500 ;
        RECT 155.400 25.200 156.300 32.400 ;
        RECT 158.100 25.200 159.900 27.000 ;
        RECT 164.100 25.200 165.900 27.000 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 139.950 22.950 142.050 25.050 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 154.950 23.100 157.050 25.200 ;
        RECT 157.950 23.100 160.050 25.200 ;
        RECT 160.950 23.100 163.050 25.200 ;
        RECT 163.950 23.100 166.050 25.200 ;
        RECT 137.100 21.150 138.900 22.950 ;
        RECT 114.750 17.100 125.850 17.700 ;
        RECT 64.800 3.600 66.600 9.600 ;
        RECT 67.800 3.000 69.600 9.600 ;
        RECT 80.400 3.000 82.200 9.600 ;
        RECT 83.400 3.600 85.200 9.600 ;
        RECT 86.400 3.000 88.200 9.600 ;
        RECT 92.550 3.600 94.350 15.600 ;
        RECT 97.950 15.300 100.050 16.200 ;
        RECT 100.950 15.300 106.050 16.200 ;
        RECT 108.150 16.500 125.850 17.100 ;
        RECT 108.150 16.200 116.550 16.500 ;
        RECT 100.950 14.400 101.850 15.300 ;
        RECT 99.150 12.600 101.850 14.400 ;
        RECT 102.750 14.100 104.550 14.400 ;
        RECT 108.150 14.100 109.050 16.200 ;
        RECT 124.950 15.600 125.850 16.500 ;
        RECT 140.400 15.600 141.300 22.950 ;
        RECT 143.100 21.150 144.900 22.950 ;
        RECT 142.950 18.450 145.050 19.050 ;
        RECT 151.950 18.450 154.050 19.050 ;
        RECT 142.950 17.550 154.050 18.450 ;
        RECT 142.950 16.950 145.050 17.550 ;
        RECT 151.950 16.950 154.050 17.550 ;
        RECT 155.400 15.600 156.300 23.100 ;
        RECT 161.100 21.300 162.900 23.100 ;
        RECT 168.150 17.700 169.050 32.400 ;
        RECT 176.550 31.800 178.350 33.600 ;
        RECT 179.850 33.450 184.800 34.500 ;
        RECT 192.300 34.500 193.350 35.400 ;
        RECT 179.850 32.700 181.650 33.450 ;
        RECT 192.300 33.300 196.050 34.500 ;
        RECT 193.950 32.400 196.050 33.300 ;
        RECT 199.650 32.400 201.450 38.400 ;
        RECT 211.800 35.400 213.600 39.000 ;
        RECT 214.800 35.400 216.600 38.400 ;
        RECT 217.800 35.400 219.600 39.000 ;
        RECT 176.850 30.000 177.900 31.800 ;
        RECT 187.050 30.000 188.850 30.600 ;
        RECT 176.850 28.800 188.850 30.000 ;
        RECT 171.000 27.600 177.900 28.800 ;
        RECT 171.000 26.850 171.900 27.600 ;
        RECT 176.100 27.000 177.900 27.600 ;
        RECT 170.100 25.050 171.900 26.850 ;
        RECT 173.100 25.800 174.900 26.400 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 173.100 24.600 181.050 25.800 ;
        RECT 178.950 22.950 181.050 24.600 ;
        RECT 177.450 17.700 179.250 18.000 ;
        RECT 168.150 17.100 179.250 17.700 ;
        RECT 168.150 16.500 185.850 17.100 ;
        RECT 168.150 15.600 169.050 16.500 ;
        RECT 177.450 16.200 185.850 16.500 ;
        RECT 102.750 13.200 109.050 14.100 ;
        RECT 109.950 14.700 111.750 15.300 ;
        RECT 109.950 13.500 117.450 14.700 ;
        RECT 102.750 12.600 104.550 13.200 ;
        RECT 116.250 12.600 117.450 13.500 ;
        RECT 97.950 9.600 101.850 11.700 ;
        RECT 106.950 11.550 108.750 12.300 ;
        RECT 111.750 11.550 113.550 12.300 ;
        RECT 106.950 10.500 113.550 11.550 ;
        RECT 116.250 10.500 121.050 12.600 ;
        RECT 95.550 3.000 97.350 6.600 ;
        RECT 100.050 3.600 101.850 9.600 ;
        RECT 104.250 3.000 106.050 9.600 ;
        RECT 107.850 3.600 109.650 10.500 ;
        RECT 116.250 9.600 117.450 10.500 ;
        RECT 110.850 3.000 112.650 9.600 ;
        RECT 115.650 3.600 117.450 9.600 ;
        RECT 121.050 3.000 122.850 9.600 ;
        RECT 124.050 3.600 125.850 15.600 ;
        RECT 137.700 14.400 141.300 15.600 ;
        RECT 137.700 3.600 139.500 14.400 ;
        RECT 142.800 3.000 144.600 15.600 ;
        RECT 154.800 3.600 156.600 15.600 ;
        RECT 157.800 14.700 165.600 15.600 ;
        RECT 157.800 3.600 159.600 14.700 ;
        RECT 160.800 3.000 162.600 13.800 ;
        RECT 163.800 3.600 165.600 14.700 ;
        RECT 168.150 3.600 169.950 15.600 ;
        RECT 182.250 14.700 184.050 15.300 ;
        RECT 176.550 13.500 184.050 14.700 ;
        RECT 184.950 14.100 185.850 16.200 ;
        RECT 187.950 16.200 188.850 28.800 ;
        RECT 200.250 25.050 201.450 32.400 ;
        RECT 215.400 25.050 216.300 35.400 ;
        RECT 229.800 32.400 231.600 38.400 ;
        RECT 230.400 30.300 231.600 32.400 ;
        RECT 232.800 33.300 234.600 38.400 ;
        RECT 235.800 34.200 237.600 39.000 ;
        RECT 238.800 33.300 240.600 38.400 ;
        RECT 232.800 31.950 240.600 33.300 ;
        RECT 248.700 32.400 250.500 39.000 ;
        RECT 253.800 31.200 255.600 38.400 ;
        RECT 251.400 30.300 255.600 31.200 ;
        RECT 269.400 31.200 271.200 38.400 ;
        RECT 274.500 32.400 276.300 39.000 ;
        RECT 286.800 32.400 288.600 38.400 ;
        RECT 269.400 30.300 273.600 31.200 ;
        RECT 230.400 29.250 234.150 30.300 ;
        RECT 230.100 25.050 231.900 26.850 ;
        RECT 232.950 25.050 234.150 29.250 ;
        RECT 236.100 25.050 237.900 26.850 ;
        RECT 248.100 25.200 249.900 27.000 ;
        RECT 251.400 25.200 252.600 30.300 ;
        RECT 254.100 25.200 255.900 27.000 ;
        RECT 269.100 25.200 270.900 27.000 ;
        RECT 272.400 25.200 273.600 30.300 ;
        RECT 287.400 30.300 288.600 32.400 ;
        RECT 289.800 33.300 291.600 38.400 ;
        RECT 292.800 34.200 294.600 39.000 ;
        RECT 295.800 33.300 297.600 38.400 ;
        RECT 289.800 31.950 297.600 33.300 ;
        RECT 300.150 32.400 301.950 38.400 ;
        RECT 303.150 35.400 304.950 39.000 ;
        RECT 307.950 36.300 309.750 38.400 ;
        RECT 306.000 35.400 309.750 36.300 ;
        RECT 312.450 35.400 314.250 39.000 ;
        RECT 315.750 35.400 317.550 38.400 ;
        RECT 319.350 35.400 321.150 39.000 ;
        RECT 323.550 35.400 325.350 38.400 ;
        RECT 328.350 35.400 330.150 39.000 ;
        RECT 306.000 34.500 307.050 35.400 ;
        RECT 315.750 34.500 316.800 35.400 ;
        RECT 304.950 32.400 307.050 34.500 ;
        RECT 287.400 29.250 291.150 30.300 ;
        RECT 275.100 25.200 276.900 27.000 ;
        RECT 195.150 23.250 201.450 25.050 ;
        RECT 196.950 22.950 201.450 23.250 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 229.950 22.950 232.050 25.050 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 247.950 23.100 250.050 25.200 ;
        RECT 250.950 23.100 253.050 25.200 ;
        RECT 253.950 23.100 256.050 25.200 ;
        RECT 268.950 23.100 271.050 25.200 ;
        RECT 271.950 23.100 274.050 25.200 ;
        RECT 274.950 23.100 277.050 25.200 ;
        RECT 287.100 25.050 288.900 26.850 ;
        RECT 289.950 25.050 291.150 29.250 ;
        RECT 293.100 25.050 294.900 26.850 ;
        RECT 197.250 17.400 199.050 19.200 ;
        RECT 193.950 16.200 198.150 17.400 ;
        RECT 187.950 15.300 193.050 16.200 ;
        RECT 193.950 15.300 196.050 16.200 ;
        RECT 200.250 15.600 201.450 22.950 ;
        RECT 212.100 21.150 213.900 22.950 ;
        RECT 215.400 15.600 216.300 22.950 ;
        RECT 218.100 21.150 219.900 22.950 ;
        RECT 192.150 14.400 193.050 15.300 ;
        RECT 189.450 14.100 191.250 14.400 ;
        RECT 176.550 12.600 177.750 13.500 ;
        RECT 184.950 13.200 191.250 14.100 ;
        RECT 189.450 12.600 191.250 13.200 ;
        RECT 192.150 12.600 194.850 14.400 ;
        RECT 172.950 10.500 177.750 12.600 ;
        RECT 180.450 11.550 182.250 12.300 ;
        RECT 185.250 11.550 187.050 12.300 ;
        RECT 180.450 10.500 187.050 11.550 ;
        RECT 176.550 9.600 177.750 10.500 ;
        RECT 171.150 3.000 172.950 9.600 ;
        RECT 176.550 3.600 178.350 9.600 ;
        RECT 181.350 3.000 183.150 9.600 ;
        RECT 184.350 3.600 186.150 10.500 ;
        RECT 192.150 9.600 196.050 11.700 ;
        RECT 187.950 3.000 189.750 9.600 ;
        RECT 192.150 3.600 193.950 9.600 ;
        RECT 196.650 3.000 198.450 6.600 ;
        RECT 199.650 3.600 201.450 15.600 ;
        RECT 212.700 14.400 216.300 15.600 ;
        RECT 212.700 3.600 214.500 14.400 ;
        RECT 217.800 3.000 219.600 15.600 ;
        RECT 233.850 9.600 235.050 22.950 ;
        RECT 239.100 21.150 240.900 22.950 ;
        RECT 230.400 3.000 232.200 9.600 ;
        RECT 233.400 3.600 235.200 9.600 ;
        RECT 238.500 3.000 240.300 15.600 ;
        RECT 251.400 9.600 252.600 23.100 ;
        RECT 253.950 21.450 256.050 22.050 ;
        RECT 259.950 21.450 262.050 22.050 ;
        RECT 253.950 20.550 262.050 21.450 ;
        RECT 253.950 19.950 256.050 20.550 ;
        RECT 259.950 19.950 262.050 20.550 ;
        RECT 272.400 9.600 273.600 23.100 ;
        RECT 286.950 22.950 289.050 25.050 ;
        RECT 289.950 22.950 292.050 25.050 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 290.850 9.600 292.050 22.950 ;
        RECT 296.100 21.150 297.900 22.950 ;
        RECT 300.150 17.700 301.050 32.400 ;
        RECT 308.550 31.800 310.350 33.600 ;
        RECT 311.850 33.450 316.800 34.500 ;
        RECT 324.300 34.500 325.350 35.400 ;
        RECT 311.850 32.700 313.650 33.450 ;
        RECT 324.300 33.300 328.050 34.500 ;
        RECT 325.950 32.400 328.050 33.300 ;
        RECT 331.650 32.400 333.450 38.400 ;
        RECT 341.400 35.400 343.200 39.000 ;
        RECT 344.400 35.400 346.200 38.400 ;
        RECT 356.400 35.400 358.200 39.000 ;
        RECT 359.400 35.400 361.200 38.400 ;
        RECT 373.800 35.400 375.600 38.400 ;
        RECT 376.800 35.400 378.600 39.000 ;
        RECT 308.850 30.000 309.900 31.800 ;
        RECT 319.050 30.000 320.850 30.600 ;
        RECT 308.850 28.800 320.850 30.000 ;
        RECT 303.000 27.600 309.900 28.800 ;
        RECT 303.000 26.850 303.900 27.600 ;
        RECT 308.100 27.000 309.900 27.600 ;
        RECT 302.100 25.050 303.900 26.850 ;
        RECT 305.100 25.800 306.900 26.400 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 305.100 24.600 313.050 25.800 ;
        RECT 310.950 22.950 313.050 24.600 ;
        RECT 309.450 17.700 311.250 18.000 ;
        RECT 300.150 17.100 311.250 17.700 ;
        RECT 300.150 16.500 317.850 17.100 ;
        RECT 300.150 15.600 301.050 16.500 ;
        RECT 309.450 16.200 317.850 16.500 ;
        RECT 248.400 3.000 250.200 9.600 ;
        RECT 251.400 3.600 253.200 9.600 ;
        RECT 254.400 3.000 256.200 9.600 ;
        RECT 268.800 3.000 270.600 9.600 ;
        RECT 271.800 3.600 273.600 9.600 ;
        RECT 274.800 3.000 276.600 9.600 ;
        RECT 287.400 3.000 289.200 9.600 ;
        RECT 290.400 3.600 292.200 9.600 ;
        RECT 295.500 3.000 297.300 15.600 ;
        RECT 300.150 3.600 301.950 15.600 ;
        RECT 314.250 14.700 316.050 15.300 ;
        RECT 308.550 13.500 316.050 14.700 ;
        RECT 316.950 14.100 317.850 16.200 ;
        RECT 319.950 16.200 320.850 28.800 ;
        RECT 332.250 25.050 333.450 32.400 ;
        RECT 344.400 25.050 345.600 35.400 ;
        RECT 359.400 25.050 360.600 35.400 ;
        RECT 374.400 25.050 375.600 35.400 ;
        RECT 388.800 32.400 390.600 38.400 ;
        RECT 389.400 30.300 390.600 32.400 ;
        RECT 391.800 33.300 393.600 38.400 ;
        RECT 394.800 34.200 396.600 39.000 ;
        RECT 397.800 33.300 399.600 38.400 ;
        RECT 409.800 35.400 411.600 38.400 ;
        RECT 412.800 35.400 414.600 39.000 ;
        RECT 391.800 31.950 399.600 33.300 ;
        RECT 389.400 29.250 393.150 30.300 ;
        RECT 389.100 25.050 390.900 26.850 ;
        RECT 391.950 25.050 393.150 29.250 ;
        RECT 405.000 27.450 409.050 28.050 ;
        RECT 395.100 25.050 396.900 26.850 ;
        RECT 404.550 25.950 409.050 27.450 ;
        RECT 327.150 23.250 333.450 25.050 ;
        RECT 328.950 22.950 333.450 23.250 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 373.950 22.950 376.050 25.050 ;
        RECT 376.950 22.950 379.050 25.050 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 394.950 22.950 397.050 25.050 ;
        RECT 397.950 22.950 400.050 25.050 ;
        RECT 329.250 17.400 331.050 19.200 ;
        RECT 325.950 16.200 330.150 17.400 ;
        RECT 319.950 15.300 325.050 16.200 ;
        RECT 325.950 15.300 328.050 16.200 ;
        RECT 332.250 15.600 333.450 22.950 ;
        RECT 341.100 21.150 342.900 22.950 ;
        RECT 324.150 14.400 325.050 15.300 ;
        RECT 321.450 14.100 323.250 14.400 ;
        RECT 308.550 12.600 309.750 13.500 ;
        RECT 316.950 13.200 323.250 14.100 ;
        RECT 321.450 12.600 323.250 13.200 ;
        RECT 324.150 12.600 326.850 14.400 ;
        RECT 304.950 10.500 309.750 12.600 ;
        RECT 312.450 11.550 314.250 12.300 ;
        RECT 317.250 11.550 319.050 12.300 ;
        RECT 312.450 10.500 319.050 11.550 ;
        RECT 308.550 9.600 309.750 10.500 ;
        RECT 303.150 3.000 304.950 9.600 ;
        RECT 308.550 3.600 310.350 9.600 ;
        RECT 313.350 3.000 315.150 9.600 ;
        RECT 316.350 3.600 318.150 10.500 ;
        RECT 324.150 9.600 328.050 11.700 ;
        RECT 319.950 3.000 321.750 9.600 ;
        RECT 324.150 3.600 325.950 9.600 ;
        RECT 328.650 3.000 330.450 6.600 ;
        RECT 331.650 3.600 333.450 15.600 ;
        RECT 344.400 9.600 345.600 22.950 ;
        RECT 356.100 21.150 357.900 22.950 ;
        RECT 359.400 9.600 360.600 22.950 ;
        RECT 364.950 15.450 367.050 16.050 ;
        RECT 370.950 15.450 373.050 16.050 ;
        RECT 364.950 14.550 373.050 15.450 ;
        RECT 364.950 13.950 367.050 14.550 ;
        RECT 370.950 13.950 373.050 14.550 ;
        RECT 374.400 9.600 375.600 22.950 ;
        RECT 377.100 21.150 378.900 22.950 ;
        RECT 392.850 9.600 394.050 22.950 ;
        RECT 398.100 21.150 399.900 22.950 ;
        RECT 404.550 22.050 405.450 25.950 ;
        RECT 410.400 25.050 411.600 35.400 ;
        RECT 422.400 33.300 424.200 38.400 ;
        RECT 425.400 34.200 427.200 39.000 ;
        RECT 428.400 33.300 430.200 38.400 ;
        RECT 422.400 31.950 430.200 33.300 ;
        RECT 431.400 32.400 433.200 38.400 ;
        RECT 438.150 32.400 439.950 38.400 ;
        RECT 441.150 35.400 442.950 39.000 ;
        RECT 445.950 36.300 447.750 38.400 ;
        RECT 444.000 35.400 447.750 36.300 ;
        RECT 450.450 35.400 452.250 39.000 ;
        RECT 453.750 35.400 455.550 38.400 ;
        RECT 457.350 35.400 459.150 39.000 ;
        RECT 461.550 35.400 463.350 38.400 ;
        RECT 466.350 35.400 468.150 39.000 ;
        RECT 444.000 34.500 445.050 35.400 ;
        RECT 453.750 34.500 454.800 35.400 ;
        RECT 442.950 32.400 445.050 34.500 ;
        RECT 431.400 30.300 432.600 32.400 ;
        RECT 428.850 29.250 432.600 30.300 ;
        RECT 425.100 25.050 426.900 26.850 ;
        RECT 428.850 25.050 430.050 29.250 ;
        RECT 431.100 25.050 432.900 26.850 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 421.950 22.950 424.050 25.050 ;
        RECT 424.950 22.950 427.050 25.050 ;
        RECT 427.950 22.950 430.050 25.050 ;
        RECT 430.950 22.950 433.050 25.050 ;
        RECT 404.550 20.550 409.050 22.050 ;
        RECT 405.000 19.950 409.050 20.550 ;
        RECT 341.400 3.000 343.200 9.600 ;
        RECT 344.400 3.600 346.200 9.600 ;
        RECT 356.400 3.000 358.200 9.600 ;
        RECT 359.400 3.600 361.200 9.600 ;
        RECT 373.800 3.600 375.600 9.600 ;
        RECT 376.800 3.000 378.600 9.600 ;
        RECT 389.400 3.000 391.200 9.600 ;
        RECT 392.400 3.600 394.200 9.600 ;
        RECT 397.500 3.000 399.300 15.600 ;
        RECT 410.400 9.600 411.600 22.950 ;
        RECT 413.100 21.150 414.900 22.950 ;
        RECT 422.100 21.150 423.900 22.950 ;
        RECT 409.800 3.600 411.600 9.600 ;
        RECT 412.800 3.000 414.600 9.600 ;
        RECT 422.700 3.000 424.500 15.600 ;
        RECT 427.950 9.600 429.150 22.950 ;
        RECT 438.150 17.700 439.050 32.400 ;
        RECT 446.550 31.800 448.350 33.600 ;
        RECT 449.850 33.450 454.800 34.500 ;
        RECT 462.300 34.500 463.350 35.400 ;
        RECT 449.850 32.700 451.650 33.450 ;
        RECT 462.300 33.300 466.050 34.500 ;
        RECT 463.950 32.400 466.050 33.300 ;
        RECT 469.650 32.400 471.450 38.400 ;
        RECT 481.800 35.400 483.600 38.400 ;
        RECT 484.800 35.400 486.600 39.000 ;
        RECT 446.850 30.000 447.900 31.800 ;
        RECT 457.050 30.000 458.850 30.600 ;
        RECT 446.850 28.800 458.850 30.000 ;
        RECT 441.000 27.600 447.900 28.800 ;
        RECT 441.000 26.850 441.900 27.600 ;
        RECT 446.100 27.000 447.900 27.600 ;
        RECT 440.100 25.050 441.900 26.850 ;
        RECT 443.100 25.800 444.900 26.400 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 443.100 24.600 451.050 25.800 ;
        RECT 448.950 22.950 451.050 24.600 ;
        RECT 447.450 17.700 449.250 18.000 ;
        RECT 438.150 17.100 449.250 17.700 ;
        RECT 438.150 16.500 455.850 17.100 ;
        RECT 438.150 15.600 439.050 16.500 ;
        RECT 447.450 16.200 455.850 16.500 ;
        RECT 427.800 3.600 429.600 9.600 ;
        RECT 430.800 3.000 432.600 9.600 ;
        RECT 438.150 3.600 439.950 15.600 ;
        RECT 452.250 14.700 454.050 15.300 ;
        RECT 446.550 13.500 454.050 14.700 ;
        RECT 454.950 14.100 455.850 16.200 ;
        RECT 457.950 16.200 458.850 28.800 ;
        RECT 470.250 25.050 471.450 32.400 ;
        RECT 482.400 25.050 483.600 35.400 ;
        RECT 497.400 31.200 499.200 38.400 ;
        RECT 502.500 32.400 504.300 39.000 ;
        RECT 514.800 32.400 516.600 38.400 ;
        RECT 497.400 30.300 501.600 31.200 ;
        RECT 497.100 25.200 498.900 27.000 ;
        RECT 500.400 25.200 501.600 30.300 ;
        RECT 515.400 30.300 516.600 32.400 ;
        RECT 517.800 33.300 519.600 38.400 ;
        RECT 520.800 34.200 522.600 39.000 ;
        RECT 523.800 33.300 525.600 38.400 ;
        RECT 517.800 31.950 525.600 33.300 ;
        RECT 527.550 32.400 529.350 38.400 ;
        RECT 530.850 35.400 532.650 39.000 ;
        RECT 535.650 35.400 537.450 38.400 ;
        RECT 539.850 35.400 541.650 39.000 ;
        RECT 543.450 35.400 545.250 38.400 ;
        RECT 546.750 35.400 548.550 39.000 ;
        RECT 551.250 36.300 553.050 38.400 ;
        RECT 551.250 35.400 555.000 36.300 ;
        RECT 556.050 35.400 557.850 39.000 ;
        RECT 535.650 34.500 536.700 35.400 ;
        RECT 532.950 33.300 536.700 34.500 ;
        RECT 544.200 34.500 545.250 35.400 ;
        RECT 553.950 34.500 555.000 35.400 ;
        RECT 544.200 33.450 549.150 34.500 ;
        RECT 532.950 32.400 535.050 33.300 ;
        RECT 547.350 32.700 549.150 33.450 ;
        RECT 515.400 29.250 519.150 30.300 ;
        RECT 503.100 25.200 504.900 27.000 ;
        RECT 465.150 23.250 471.450 25.050 ;
        RECT 466.950 22.950 471.450 23.250 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 496.950 23.100 499.050 25.200 ;
        RECT 499.950 23.100 502.050 25.200 ;
        RECT 502.950 23.100 505.050 25.200 ;
        RECT 515.100 25.050 516.900 26.850 ;
        RECT 517.950 25.050 519.150 29.250 ;
        RECT 521.100 25.050 522.900 26.850 ;
        RECT 527.550 25.050 528.750 32.400 ;
        RECT 550.650 31.800 552.450 33.600 ;
        RECT 553.950 32.400 556.050 34.500 ;
        RECT 559.050 32.400 560.850 38.400 ;
        RECT 540.150 30.000 541.950 30.600 ;
        RECT 551.100 30.000 552.150 31.800 ;
        RECT 540.150 28.800 552.150 30.000 ;
        RECT 467.250 17.400 469.050 19.200 ;
        RECT 463.950 16.200 468.150 17.400 ;
        RECT 457.950 15.300 463.050 16.200 ;
        RECT 463.950 15.300 466.050 16.200 ;
        RECT 470.250 15.600 471.450 22.950 ;
        RECT 462.150 14.400 463.050 15.300 ;
        RECT 459.450 14.100 461.250 14.400 ;
        RECT 446.550 12.600 447.750 13.500 ;
        RECT 454.950 13.200 461.250 14.100 ;
        RECT 459.450 12.600 461.250 13.200 ;
        RECT 462.150 12.600 464.850 14.400 ;
        RECT 442.950 10.500 447.750 12.600 ;
        RECT 450.450 11.550 452.250 12.300 ;
        RECT 455.250 11.550 457.050 12.300 ;
        RECT 450.450 10.500 457.050 11.550 ;
        RECT 446.550 9.600 447.750 10.500 ;
        RECT 441.150 3.000 442.950 9.600 ;
        RECT 446.550 3.600 448.350 9.600 ;
        RECT 451.350 3.000 453.150 9.600 ;
        RECT 454.350 3.600 456.150 10.500 ;
        RECT 462.150 9.600 466.050 11.700 ;
        RECT 457.950 3.000 459.750 9.600 ;
        RECT 462.150 3.600 463.950 9.600 ;
        RECT 466.650 3.000 468.450 6.600 ;
        RECT 469.650 3.600 471.450 15.600 ;
        RECT 482.400 9.600 483.600 22.950 ;
        RECT 485.100 21.150 486.900 22.950 ;
        RECT 500.400 9.600 501.600 23.100 ;
        RECT 514.950 22.950 517.050 25.050 ;
        RECT 517.950 22.950 520.050 25.050 ;
        RECT 520.950 22.950 523.050 25.050 ;
        RECT 523.950 22.950 526.050 25.050 ;
        RECT 527.550 23.250 533.850 25.050 ;
        RECT 527.550 22.950 532.050 23.250 ;
        RECT 502.950 12.450 505.050 13.050 ;
        RECT 514.950 12.450 517.050 13.050 ;
        RECT 502.950 11.550 517.050 12.450 ;
        RECT 502.950 10.950 505.050 11.550 ;
        RECT 514.950 10.950 517.050 11.550 ;
        RECT 518.850 9.600 520.050 22.950 ;
        RECT 524.100 21.150 525.900 22.950 ;
        RECT 527.550 15.600 528.750 22.950 ;
        RECT 529.950 17.400 531.750 19.200 ;
        RECT 530.850 16.200 535.050 17.400 ;
        RECT 540.150 16.200 541.050 28.800 ;
        RECT 551.100 27.600 558.000 28.800 ;
        RECT 551.100 27.000 552.900 27.600 ;
        RECT 557.100 26.850 558.000 27.600 ;
        RECT 554.100 25.800 555.900 26.400 ;
        RECT 547.950 24.600 555.900 25.800 ;
        RECT 557.100 25.050 558.900 26.850 ;
        RECT 547.950 22.950 550.050 24.600 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 549.750 17.700 551.550 18.000 ;
        RECT 559.950 17.700 560.850 32.400 ;
        RECT 572.400 31.200 574.200 38.400 ;
        RECT 577.500 32.400 579.300 39.000 ;
        RECT 589.800 32.400 591.600 38.400 ;
        RECT 572.400 30.300 576.600 31.200 ;
        RECT 572.100 25.200 573.900 27.000 ;
        RECT 575.400 25.200 576.600 30.300 ;
        RECT 590.400 30.300 591.600 32.400 ;
        RECT 592.800 33.300 594.600 38.400 ;
        RECT 595.800 34.200 597.600 39.000 ;
        RECT 598.800 33.300 600.600 38.400 ;
        RECT 592.800 31.950 600.600 33.300 ;
        RECT 603.150 32.400 604.950 38.400 ;
        RECT 606.150 35.400 607.950 39.000 ;
        RECT 610.950 36.300 612.750 38.400 ;
        RECT 609.000 35.400 612.750 36.300 ;
        RECT 615.450 35.400 617.250 39.000 ;
        RECT 618.750 35.400 620.550 38.400 ;
        RECT 622.350 35.400 624.150 39.000 ;
        RECT 626.550 35.400 628.350 38.400 ;
        RECT 631.350 35.400 633.150 39.000 ;
        RECT 609.000 34.500 610.050 35.400 ;
        RECT 618.750 34.500 619.800 35.400 ;
        RECT 607.950 32.400 610.050 34.500 ;
        RECT 590.400 29.250 594.150 30.300 ;
        RECT 580.950 27.450 585.000 28.050 ;
        RECT 578.100 25.200 579.900 27.000 ;
        RECT 580.950 25.950 585.450 27.450 ;
        RECT 571.950 23.100 574.050 25.200 ;
        RECT 574.950 23.100 577.050 25.200 ;
        RECT 577.950 23.100 580.050 25.200 ;
        RECT 565.950 21.450 568.050 22.050 ;
        RECT 571.950 21.450 574.050 22.050 ;
        RECT 565.950 20.550 574.050 21.450 ;
        RECT 565.950 19.950 568.050 20.550 ;
        RECT 571.950 19.950 574.050 20.550 ;
        RECT 549.750 17.100 560.850 17.700 ;
        RECT 481.800 3.600 483.600 9.600 ;
        RECT 484.800 3.000 486.600 9.600 ;
        RECT 496.800 3.000 498.600 9.600 ;
        RECT 499.800 3.600 501.600 9.600 ;
        RECT 502.800 3.000 504.600 9.600 ;
        RECT 515.400 3.000 517.200 9.600 ;
        RECT 518.400 3.600 520.200 9.600 ;
        RECT 523.500 3.000 525.300 15.600 ;
        RECT 527.550 3.600 529.350 15.600 ;
        RECT 532.950 15.300 535.050 16.200 ;
        RECT 535.950 15.300 541.050 16.200 ;
        RECT 543.150 16.500 560.850 17.100 ;
        RECT 543.150 16.200 551.550 16.500 ;
        RECT 535.950 14.400 536.850 15.300 ;
        RECT 534.150 12.600 536.850 14.400 ;
        RECT 537.750 14.100 539.550 14.400 ;
        RECT 543.150 14.100 544.050 16.200 ;
        RECT 559.950 15.600 560.850 16.500 ;
        RECT 537.750 13.200 544.050 14.100 ;
        RECT 544.950 14.700 546.750 15.300 ;
        RECT 544.950 13.500 552.450 14.700 ;
        RECT 537.750 12.600 539.550 13.200 ;
        RECT 551.250 12.600 552.450 13.500 ;
        RECT 532.950 9.600 536.850 11.700 ;
        RECT 541.950 11.550 543.750 12.300 ;
        RECT 546.750 11.550 548.550 12.300 ;
        RECT 541.950 10.500 548.550 11.550 ;
        RECT 551.250 10.500 556.050 12.600 ;
        RECT 530.550 3.000 532.350 6.600 ;
        RECT 535.050 3.600 536.850 9.600 ;
        RECT 539.250 3.000 541.050 9.600 ;
        RECT 542.850 3.600 544.650 10.500 ;
        RECT 551.250 9.600 552.450 10.500 ;
        RECT 545.850 3.000 547.650 9.600 ;
        RECT 550.650 3.600 552.450 9.600 ;
        RECT 556.050 3.000 557.850 9.600 ;
        RECT 559.050 3.600 560.850 15.600 ;
        RECT 575.400 9.600 576.600 23.100 ;
        RECT 584.550 22.050 585.450 25.950 ;
        RECT 590.100 25.050 591.900 26.850 ;
        RECT 592.950 25.050 594.150 29.250 ;
        RECT 596.100 25.050 597.900 26.850 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 592.950 22.950 595.050 25.050 ;
        RECT 595.950 22.950 598.050 25.050 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 584.550 20.550 589.050 22.050 ;
        RECT 585.000 19.950 589.050 20.550 ;
        RECT 593.850 9.600 595.050 22.950 ;
        RECT 599.100 21.150 600.900 22.950 ;
        RECT 603.150 17.700 604.050 32.400 ;
        RECT 611.550 31.800 613.350 33.600 ;
        RECT 614.850 33.450 619.800 34.500 ;
        RECT 627.300 34.500 628.350 35.400 ;
        RECT 614.850 32.700 616.650 33.450 ;
        RECT 627.300 33.300 631.050 34.500 ;
        RECT 628.950 32.400 631.050 33.300 ;
        RECT 634.650 32.400 636.450 38.400 ;
        RECT 611.850 30.000 612.900 31.800 ;
        RECT 622.050 30.000 623.850 30.600 ;
        RECT 611.850 28.800 623.850 30.000 ;
        RECT 606.000 27.600 612.900 28.800 ;
        RECT 606.000 26.850 606.900 27.600 ;
        RECT 611.100 27.000 612.900 27.600 ;
        RECT 605.100 25.050 606.900 26.850 ;
        RECT 608.100 25.800 609.900 26.400 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 608.100 24.600 616.050 25.800 ;
        RECT 613.950 22.950 616.050 24.600 ;
        RECT 612.450 17.700 614.250 18.000 ;
        RECT 603.150 17.100 614.250 17.700 ;
        RECT 603.150 16.500 620.850 17.100 ;
        RECT 603.150 15.600 604.050 16.500 ;
        RECT 612.450 16.200 620.850 16.500 ;
        RECT 571.800 3.000 573.600 9.600 ;
        RECT 574.800 3.600 576.600 9.600 ;
        RECT 577.800 3.000 579.600 9.600 ;
        RECT 590.400 3.000 592.200 9.600 ;
        RECT 593.400 3.600 595.200 9.600 ;
        RECT 598.500 3.000 600.300 15.600 ;
        RECT 603.150 3.600 604.950 15.600 ;
        RECT 617.250 14.700 619.050 15.300 ;
        RECT 611.550 13.500 619.050 14.700 ;
        RECT 619.950 14.100 620.850 16.200 ;
        RECT 622.950 16.200 623.850 28.800 ;
        RECT 635.250 25.050 636.450 32.400 ;
        RECT 644.400 35.400 646.200 38.400 ;
        RECT 647.400 35.400 649.200 39.000 ;
        RECT 644.400 31.500 645.600 35.400 ;
        RECT 650.400 32.400 652.200 38.400 ;
        RECT 662.400 35.400 664.200 39.000 ;
        RECT 665.400 35.400 667.200 38.400 ;
        RECT 677.400 35.400 679.200 39.000 ;
        RECT 680.400 35.400 682.200 38.400 ;
        RECT 683.400 35.400 685.200 39.000 ;
        RECT 697.800 35.400 699.600 38.400 ;
        RECT 700.800 35.400 702.600 39.000 ;
        RECT 713.700 35.400 715.500 39.000 ;
        RECT 644.400 30.600 650.100 31.500 ;
        RECT 648.150 29.700 650.100 30.600 ;
        RECT 630.150 23.250 636.450 25.050 ;
        RECT 631.950 22.950 636.450 23.250 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 632.250 17.400 634.050 19.200 ;
        RECT 628.950 16.200 633.150 17.400 ;
        RECT 622.950 15.300 628.050 16.200 ;
        RECT 628.950 15.300 631.050 16.200 ;
        RECT 635.250 15.600 636.450 22.950 ;
        RECT 644.100 21.150 645.900 22.950 ;
        RECT 648.150 18.300 649.050 29.700 ;
        RECT 651.000 25.050 652.200 32.400 ;
        RECT 665.400 25.050 666.600 35.400 ;
        RECT 680.700 25.050 681.600 35.400 ;
        RECT 698.400 25.050 699.600 35.400 ;
        RECT 716.700 33.600 718.500 38.400 ;
        RECT 713.400 32.400 718.500 33.600 ;
        RECT 721.200 32.400 723.000 39.000 ;
        RECT 731.400 35.400 733.200 39.000 ;
        RECT 734.400 35.400 736.200 38.400 ;
        RECT 746.400 35.400 748.200 39.000 ;
        RECT 749.400 35.400 751.200 38.400 ;
        RECT 752.400 35.400 754.200 39.000 ;
        RECT 713.400 25.200 714.300 32.400 ;
        RECT 716.100 25.200 717.900 27.000 ;
        RECT 722.100 25.200 723.900 27.000 ;
        RECT 649.950 22.950 652.200 25.050 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 664.950 22.950 667.050 25.050 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 697.950 22.950 700.050 25.050 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 712.950 23.100 715.050 25.200 ;
        RECT 715.950 23.100 718.050 25.200 ;
        RECT 718.950 23.100 721.050 25.200 ;
        RECT 721.950 23.100 724.050 25.200 ;
        RECT 734.400 25.050 735.600 35.400 ;
        RECT 736.950 27.450 741.000 28.050 ;
        RECT 736.950 25.950 741.450 27.450 ;
        RECT 648.150 17.400 650.100 18.300 ;
        RECT 627.150 14.400 628.050 15.300 ;
        RECT 624.450 14.100 626.250 14.400 ;
        RECT 611.550 12.600 612.750 13.500 ;
        RECT 619.950 13.200 626.250 14.100 ;
        RECT 624.450 12.600 626.250 13.200 ;
        RECT 627.150 12.600 629.850 14.400 ;
        RECT 607.950 10.500 612.750 12.600 ;
        RECT 615.450 11.550 617.250 12.300 ;
        RECT 620.250 11.550 622.050 12.300 ;
        RECT 615.450 10.500 622.050 11.550 ;
        RECT 611.550 9.600 612.750 10.500 ;
        RECT 606.150 3.000 607.950 9.600 ;
        RECT 611.550 3.600 613.350 9.600 ;
        RECT 616.350 3.000 618.150 9.600 ;
        RECT 619.350 3.600 621.150 10.500 ;
        RECT 627.150 9.600 631.050 11.700 ;
        RECT 622.950 3.000 624.750 9.600 ;
        RECT 627.150 3.600 628.950 9.600 ;
        RECT 631.650 3.000 633.450 6.600 ;
        RECT 634.650 3.600 636.450 15.600 ;
        RECT 644.400 16.500 650.100 17.400 ;
        RECT 644.400 9.600 645.600 16.500 ;
        RECT 651.000 15.600 652.200 22.950 ;
        RECT 662.100 21.150 663.900 22.950 ;
        RECT 644.400 3.600 646.200 9.600 ;
        RECT 647.400 3.000 649.200 9.600 ;
        RECT 650.400 3.600 652.200 15.600 ;
        RECT 665.400 9.600 666.600 22.950 ;
        RECT 677.100 21.150 678.900 22.950 ;
        RECT 680.700 15.600 681.600 22.950 ;
        RECT 683.100 21.150 684.900 22.950 ;
        RECT 662.400 3.000 664.200 9.600 ;
        RECT 665.400 3.600 667.200 9.600 ;
        RECT 677.400 3.000 679.200 15.600 ;
        RECT 680.700 14.400 684.300 15.600 ;
        RECT 682.500 3.600 684.300 14.400 ;
        RECT 698.400 9.600 699.600 22.950 ;
        RECT 701.100 21.150 702.900 22.950 ;
        RECT 713.400 15.600 714.300 23.100 ;
        RECT 719.100 21.300 720.900 23.100 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 733.950 22.950 736.050 25.050 ;
        RECT 731.100 21.150 732.900 22.950 ;
        RECT 697.800 3.600 699.600 9.600 ;
        RECT 700.800 3.000 702.600 9.600 ;
        RECT 712.800 3.600 714.600 15.600 ;
        RECT 715.800 14.700 723.600 15.600 ;
        RECT 715.800 3.600 717.600 14.700 ;
        RECT 718.800 3.000 720.600 13.800 ;
        RECT 721.800 3.600 723.600 14.700 ;
        RECT 734.400 9.600 735.600 22.950 ;
        RECT 740.550 22.050 741.450 25.950 ;
        RECT 749.700 25.050 750.600 35.400 ;
        RECT 751.950 33.450 754.050 34.050 ;
        RECT 757.950 33.450 760.050 34.050 ;
        RECT 751.950 32.550 760.050 33.450 ;
        RECT 751.950 31.950 754.050 32.550 ;
        RECT 757.950 31.950 760.050 32.550 ;
        RECT 766.800 32.400 768.600 38.400 ;
        RECT 751.950 30.450 754.050 30.900 ;
        RECT 760.950 30.450 763.050 31.050 ;
        RECT 751.950 29.550 763.050 30.450 ;
        RECT 751.950 28.800 754.050 29.550 ;
        RECT 760.950 28.950 763.050 29.550 ;
        RECT 767.400 30.300 768.600 32.400 ;
        RECT 769.800 33.300 771.600 38.400 ;
        RECT 772.800 34.200 774.600 39.000 ;
        RECT 785.400 38.400 786.600 39.000 ;
        RECT 775.800 33.300 777.600 38.400 ;
        RECT 785.400 35.400 787.200 38.400 ;
        RECT 788.400 35.400 790.200 38.400 ;
        RECT 791.400 35.400 793.200 39.000 ;
        RECT 769.800 31.950 777.600 33.300 ;
        RECT 789.300 31.200 790.200 35.400 ;
        RECT 794.400 32.400 796.200 38.400 ;
        RECT 807.000 32.400 808.800 39.000 ;
        RECT 811.500 33.600 813.300 38.400 ;
        RECT 814.500 35.400 816.300 39.000 ;
        RECT 811.500 32.400 816.600 33.600 ;
        RECT 827.700 32.400 829.500 39.000 ;
        RECT 832.200 32.400 834.000 38.400 ;
        RECT 836.700 32.400 838.500 39.000 ;
        RECT 789.300 30.300 792.600 31.200 ;
        RECT 767.400 29.250 771.150 30.300 ;
        RECT 790.800 29.400 792.600 30.300 ;
        RECT 767.100 25.050 768.900 26.850 ;
        RECT 769.950 25.050 771.150 29.250 ;
        RECT 773.100 25.050 774.900 26.850 ;
        RECT 785.100 25.050 786.900 26.850 ;
        RECT 745.950 22.950 748.050 25.050 ;
        RECT 748.950 22.950 751.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 784.950 22.950 787.050 25.050 ;
        RECT 787.950 22.950 790.050 25.050 ;
        RECT 740.550 20.550 745.050 22.050 ;
        RECT 746.100 21.150 747.900 22.950 ;
        RECT 741.000 19.950 745.050 20.550 ;
        RECT 749.700 15.600 750.600 22.950 ;
        RECT 752.100 21.150 753.900 22.950 ;
        RECT 731.400 3.000 733.200 9.600 ;
        RECT 734.400 3.600 736.200 9.600 ;
        RECT 746.400 3.000 748.200 15.600 ;
        RECT 749.700 14.400 753.300 15.600 ;
        RECT 751.500 3.600 753.300 14.400 ;
        RECT 770.850 9.600 772.050 22.950 ;
        RECT 776.100 21.150 777.900 22.950 ;
        RECT 788.100 21.150 789.900 22.950 ;
        RECT 791.700 18.900 792.600 29.400 ;
        RECT 795.000 25.050 796.050 32.400 ;
        RECT 806.100 25.200 807.900 27.000 ;
        RECT 812.100 25.200 813.900 27.000 ;
        RECT 815.700 25.200 816.600 32.400 ;
        RECT 817.950 27.450 822.000 28.050 ;
        RECT 817.950 25.950 822.450 27.450 ;
        RECT 790.800 18.300 792.600 18.900 ;
        RECT 785.400 17.100 792.600 18.300 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 805.950 23.100 808.050 25.200 ;
        RECT 808.950 23.100 811.050 25.200 ;
        RECT 811.950 23.100 814.050 25.200 ;
        RECT 814.950 23.100 817.050 25.200 ;
        RECT 785.400 15.600 786.600 17.100 ;
        RECT 793.950 15.600 795.300 22.950 ;
        RECT 809.100 21.300 810.900 23.100 ;
        RECT 815.700 15.600 816.600 23.100 ;
        RECT 821.550 22.050 822.450 25.950 ;
        RECT 827.100 25.200 828.900 27.000 ;
        RECT 832.950 25.200 834.000 32.400 ;
        RECT 839.100 25.200 840.900 27.000 ;
        RECT 826.950 23.100 829.050 25.200 ;
        RECT 829.950 23.100 832.050 25.200 ;
        RECT 832.950 23.100 835.050 25.200 ;
        RECT 835.950 23.100 838.050 25.200 ;
        RECT 838.950 23.100 841.050 25.200 ;
        RECT 821.550 20.550 826.050 22.050 ;
        RECT 830.100 21.300 831.900 23.100 ;
        RECT 822.000 19.950 826.050 20.550 ;
        RECT 833.100 17.400 834.000 23.100 ;
        RECT 836.100 21.300 837.900 23.100 ;
        RECT 833.100 16.500 838.200 17.400 ;
        RECT 767.400 3.000 769.200 9.600 ;
        RECT 770.400 3.600 772.200 9.600 ;
        RECT 775.500 3.000 777.300 15.600 ;
        RECT 785.400 3.600 787.200 15.600 ;
        RECT 789.900 3.000 791.700 15.600 ;
        RECT 792.900 14.100 795.300 15.600 ;
        RECT 806.400 14.700 814.200 15.600 ;
        RECT 792.900 3.600 794.700 14.100 ;
        RECT 806.400 3.600 808.200 14.700 ;
        RECT 809.400 3.000 811.200 13.800 ;
        RECT 812.400 3.600 814.200 14.700 ;
        RECT 815.400 3.600 817.200 15.600 ;
        RECT 827.400 14.400 835.200 15.300 ;
        RECT 827.400 3.600 829.200 14.400 ;
        RECT 830.400 3.000 832.200 13.500 ;
        RECT 833.400 4.500 835.200 14.400 ;
        RECT 836.400 5.400 838.200 16.500 ;
        RECT 839.400 4.500 841.200 15.600 ;
        RECT 833.400 3.600 841.200 4.500 ;
      LAYER metal2 ;
        RECT 46.950 820.950 49.050 823.050 ;
        RECT 88.950 820.950 91.050 823.050 ;
        RECT 439.950 820.950 442.050 823.050 ;
        RECT 460.800 820.950 462.900 823.050 ;
        RECT 514.950 820.950 517.050 823.050 ;
        RECT 565.800 820.950 567.900 823.050 ;
        RECT 604.950 820.950 607.050 823.050 ;
        RECT 619.950 820.950 622.050 823.050 ;
        RECT 31.950 811.950 34.050 814.050 ;
        RECT 32.400 808.350 33.450 811.950 ;
        RECT 4.950 805.950 7.050 808.050 ;
        RECT 10.950 806.250 13.050 808.350 ;
        RECT 16.950 806.250 19.050 808.350 ;
        RECT 31.950 806.250 34.050 808.350 ;
        RECT 37.950 806.250 40.050 808.350 ;
        RECT 43.950 806.250 46.050 808.350 ;
        RECT 5.400 754.050 6.450 805.950 ;
        RECT 11.400 805.500 12.600 806.250 ;
        RECT 17.400 805.500 18.600 806.250 ;
        RECT 32.400 805.500 33.600 806.250 ;
        RECT 38.400 805.500 39.600 806.250 ;
        RECT 10.950 803.100 13.050 805.200 ;
        RECT 13.950 803.100 16.050 805.200 ;
        RECT 16.950 803.100 19.050 805.200 ;
        RECT 19.950 803.100 22.050 805.200 ;
        RECT 28.950 803.100 31.050 805.200 ;
        RECT 31.950 803.100 34.050 805.200 ;
        RECT 34.950 803.100 37.050 805.200 ;
        RECT 37.950 803.100 40.050 805.200 ;
        RECT 14.400 801.000 15.600 802.800 ;
        RECT 20.400 802.050 21.600 802.800 ;
        RECT 16.800 801.000 18.900 802.050 ;
        RECT 13.950 796.950 16.050 801.000 ;
        RECT 16.800 799.950 19.050 801.000 ;
        RECT 19.950 799.950 22.050 802.050 ;
        RECT 29.400 800.400 30.600 802.800 ;
        RECT 35.400 802.050 36.600 802.800 ;
        RECT 16.950 796.950 19.050 799.950 ;
        RECT 29.400 799.050 30.450 800.400 ;
        RECT 28.950 796.950 31.050 799.050 ;
        RECT 34.950 796.950 37.050 802.050 ;
        RECT 40.950 796.950 43.050 802.050 ;
        RECT 29.400 784.050 30.450 796.950 ;
        RECT 28.950 781.950 31.050 784.050 ;
        RECT 44.400 775.050 45.450 806.250 ;
        RECT 47.400 802.050 48.450 820.950 ;
        RECT 49.950 817.950 52.050 820.050 ;
        RECT 50.400 814.050 51.450 817.950 ;
        RECT 49.950 811.950 52.050 814.050 ;
        RECT 58.950 811.950 61.050 814.050 ;
        RECT 85.950 811.950 88.050 814.050 ;
        RECT 49.950 807.600 54.000 808.050 ;
        RECT 59.400 807.600 60.450 811.950 ;
        RECT 49.950 805.950 54.600 807.600 ;
        RECT 53.400 805.500 54.600 805.950 ;
        RECT 59.400 805.500 60.600 807.600 ;
        RECT 73.950 806.250 76.050 808.350 ;
        RECT 74.400 805.500 75.600 806.250 ;
        RECT 82.950 805.950 85.050 808.050 ;
        RECT 52.950 803.100 55.050 805.200 ;
        RECT 55.950 803.100 58.050 805.200 ;
        RECT 58.950 803.100 61.050 805.200 ;
        RECT 61.950 803.100 64.050 805.200 ;
        RECT 70.950 803.100 73.050 805.200 ;
        RECT 73.950 803.100 76.050 805.200 ;
        RECT 76.950 803.100 79.050 805.200 ;
        RECT 56.400 802.050 57.600 802.800 ;
        RECT 62.400 802.050 63.600 802.800 ;
        RECT 71.400 802.050 72.600 802.800 ;
        RECT 46.950 799.950 49.050 802.050 ;
        RECT 55.950 799.950 58.050 802.050 ;
        RECT 61.950 799.950 64.050 802.050 ;
        RECT 70.950 799.950 73.050 802.050 ;
        RECT 77.400 800.400 78.600 802.800 ;
        RECT 83.400 802.050 84.450 805.950 ;
        RECT 61.950 787.950 64.050 790.050 ;
        RECT 43.950 772.950 46.050 775.050 ;
        RECT 16.950 766.950 19.050 769.050 ;
        RECT 31.950 766.950 34.050 769.050 ;
        RECT 46.950 766.950 49.050 769.050 ;
        RECT 10.950 761.100 13.050 763.200 ;
        RECT 17.400 762.600 18.450 766.950 ;
        RECT 32.400 762.600 33.450 766.950 ;
        RECT 11.400 760.350 12.600 761.100 ;
        RECT 17.400 760.350 18.600 762.600 ;
        RECT 32.400 760.350 33.600 762.600 ;
        RECT 37.950 761.100 40.050 763.200 ;
        RECT 38.400 760.350 39.600 761.100 ;
        RECT 43.950 760.950 46.050 763.050 ;
        RECT 10.950 757.950 13.050 760.050 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 28.950 757.950 31.050 760.050 ;
        RECT 31.950 757.950 34.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 14.400 755.400 15.600 757.650 ;
        RECT 20.400 756.000 21.600 757.650 ;
        RECT 29.400 756.000 30.600 757.650 ;
        RECT 4.950 751.950 7.050 754.050 ;
        RECT 1.950 739.950 4.050 742.050 ;
        RECT 10.950 739.950 13.050 742.050 ;
        RECT 2.400 619.050 3.450 739.950 ;
        RECT 4.950 730.950 7.050 733.050 ;
        RECT 5.400 724.050 6.450 730.950 ;
        RECT 11.400 729.600 12.450 739.950 ;
        RECT 14.400 733.050 15.450 755.400 ;
        RECT 19.950 751.950 22.050 756.000 ;
        RECT 28.950 751.950 31.050 756.000 ;
        RECT 35.400 755.400 36.600 757.650 ;
        RECT 35.400 745.050 36.450 755.400 ;
        RECT 40.950 754.950 43.050 757.050 ;
        RECT 41.400 751.050 42.450 754.950 ;
        RECT 40.950 748.950 43.050 751.050 ;
        RECT 34.950 742.950 37.050 745.050 ;
        RECT 16.950 739.950 19.050 742.050 ;
        RECT 31.950 739.950 34.050 742.050 ;
        RECT 13.950 730.950 16.050 733.050 ;
        RECT 17.400 729.600 18.450 739.950 ;
        RECT 32.400 729.600 33.450 739.950 ;
        RECT 11.400 727.500 12.600 729.600 ;
        RECT 17.400 727.500 18.600 729.600 ;
        RECT 32.400 727.500 33.600 729.600 ;
        RECT 37.950 728.250 40.050 730.350 ;
        RECT 38.400 727.500 39.600 728.250 ;
        RECT 10.950 725.100 13.050 727.200 ;
        RECT 13.950 725.100 16.050 727.200 ;
        RECT 16.950 725.100 19.050 727.200 ;
        RECT 19.950 725.100 22.050 727.200 ;
        RECT 28.950 725.100 31.050 727.200 ;
        RECT 31.950 725.100 34.050 727.200 ;
        RECT 34.950 725.100 37.050 727.200 ;
        RECT 37.950 725.100 40.050 727.200 ;
        RECT 14.400 724.050 15.600 724.800 ;
        RECT 4.950 721.950 7.050 724.050 ;
        RECT 13.950 721.950 16.050 724.050 ;
        RECT 20.400 722.400 21.600 724.800 ;
        RECT 29.400 724.050 30.600 724.800 ;
        RECT 20.400 709.050 21.450 722.400 ;
        RECT 28.950 721.950 31.050 724.050 ;
        RECT 35.400 722.400 36.600 724.800 ;
        RECT 31.950 718.950 34.050 721.050 ;
        RECT 19.950 706.950 22.050 709.050 ;
        RECT 4.950 691.950 7.050 694.050 ;
        RECT 28.950 691.950 31.050 694.050 ;
        RECT 5.400 678.900 6.450 691.950 ;
        RECT 10.950 683.100 13.050 685.200 ;
        RECT 11.400 682.350 12.600 683.100 ;
        RECT 19.950 682.950 22.050 685.050 ;
        RECT 29.400 684.600 30.450 691.950 ;
        RECT 32.400 685.050 33.450 718.950 ;
        RECT 35.400 709.050 36.450 722.400 ;
        RECT 40.950 721.950 43.050 724.050 ;
        RECT 34.950 706.950 37.050 709.050 ;
        RECT 37.950 703.950 40.050 706.050 ;
        RECT 34.950 697.950 37.050 700.050 ;
        RECT 10.950 679.950 13.050 682.050 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 14.400 678.900 15.600 679.650 ;
        RECT 4.950 676.800 7.050 678.900 ;
        RECT 13.950 676.800 16.050 678.900 ;
        RECT 14.400 658.050 15.450 676.800 ;
        RECT 20.400 670.050 21.450 682.950 ;
        RECT 29.400 682.200 30.600 684.600 ;
        RECT 31.950 682.950 34.050 685.050 ;
        RECT 35.400 684.600 36.450 697.950 ;
        RECT 38.400 694.050 39.450 703.950 ;
        RECT 37.950 691.950 40.050 694.050 ;
        RECT 41.400 691.050 42.450 721.950 ;
        RECT 44.400 715.050 45.450 760.950 ;
        RECT 47.400 757.050 48.450 766.950 ;
        RECT 52.950 761.100 55.050 763.200 ;
        RECT 53.400 760.350 54.600 761.100 ;
        RECT 52.950 757.950 55.050 760.050 ;
        RECT 55.950 757.950 58.050 760.050 ;
        RECT 46.950 754.950 49.050 757.050 ;
        RECT 56.400 755.400 57.600 757.650 ;
        RECT 56.400 751.050 57.450 755.400 ;
        RECT 55.950 748.950 58.050 751.050 ;
        RECT 49.950 742.950 52.050 745.050 ;
        RECT 46.950 733.950 49.050 736.050 ;
        RECT 47.400 718.050 48.450 733.950 ;
        RECT 50.400 730.050 51.450 742.950 ;
        RECT 52.950 739.950 55.050 742.050 ;
        RECT 49.950 727.950 52.050 730.050 ;
        RECT 53.400 729.600 54.450 739.950 ;
        RECT 56.400 733.050 57.450 748.950 ;
        RECT 58.950 733.950 61.050 736.050 ;
        RECT 55.950 730.950 58.050 733.050 ;
        RECT 59.400 729.600 60.450 733.950 ;
        RECT 62.400 733.050 63.450 787.950 ;
        RECT 71.400 778.050 72.450 799.950 ;
        RECT 77.400 796.050 78.450 800.400 ;
        RECT 82.950 799.950 85.050 802.050 ;
        RECT 76.950 793.950 79.050 796.050 ;
        RECT 83.400 790.050 84.450 799.950 ;
        RECT 86.400 799.050 87.450 811.950 ;
        RECT 89.400 808.050 90.450 820.950 ;
        RECT 91.950 817.950 94.050 820.050 ;
        RECT 112.950 817.950 115.050 820.050 ;
        RECT 133.950 817.950 136.050 820.050 ;
        RECT 88.950 805.950 91.050 808.050 ;
        RECT 92.400 807.600 93.450 817.950 ;
        RECT 92.400 805.500 93.600 807.600 ;
        RECT 97.950 807.000 100.050 811.050 ;
        RECT 113.400 808.350 114.450 817.950 ;
        RECT 121.950 808.950 124.050 811.050 ;
        RECT 98.400 805.500 99.600 807.000 ;
        RECT 112.950 806.250 115.050 808.350 ;
        RECT 113.400 805.500 114.600 806.250 ;
        RECT 91.950 803.100 94.050 805.200 ;
        RECT 94.950 803.100 97.050 805.200 ;
        RECT 97.950 803.100 100.050 805.200 ;
        RECT 100.950 803.100 103.050 805.200 ;
        RECT 109.950 803.100 112.050 805.200 ;
        RECT 112.950 803.100 115.050 805.200 ;
        RECT 115.950 803.100 118.050 805.200 ;
        RECT 95.400 802.050 96.600 802.800 ;
        RECT 101.400 802.050 102.600 802.800 ;
        RECT 110.400 802.050 111.600 802.800 ;
        RECT 94.950 799.950 97.050 802.050 ;
        RECT 100.950 799.950 103.050 802.050 ;
        RECT 109.950 799.950 112.050 802.050 ;
        RECT 116.400 800.400 117.600 802.800 ;
        RECT 85.950 796.950 88.050 799.050 ;
        RECT 110.400 790.050 111.450 799.950 ;
        RECT 112.950 796.950 115.050 799.050 ;
        RECT 82.950 787.950 85.050 790.050 ;
        RECT 109.950 787.950 112.050 790.050 ;
        RECT 82.950 781.950 85.050 784.050 ;
        RECT 70.950 775.950 73.050 778.050 ;
        RECT 79.950 772.950 82.050 775.050 ;
        RECT 70.950 766.950 73.050 769.050 ;
        RECT 71.400 762.600 72.450 766.950 ;
        RECT 80.400 763.050 81.450 772.950 ;
        RECT 71.400 760.200 72.600 762.600 ;
        RECT 76.950 760.950 79.050 763.050 ;
        RECT 79.950 760.950 82.050 763.050 ;
        RECT 77.400 760.200 78.600 760.950 ;
        RECT 67.950 757.800 70.050 759.900 ;
        RECT 70.950 757.800 73.050 759.900 ;
        RECT 73.950 757.800 76.050 759.900 ;
        RECT 76.950 757.800 79.050 759.900 ;
        RECT 68.400 756.750 69.600 757.500 ;
        RECT 67.950 754.650 70.050 756.750 ;
        RECT 74.400 755.400 75.600 757.500 ;
        RECT 83.400 757.050 84.450 781.950 ;
        RECT 97.950 766.950 100.050 769.050 ;
        RECT 106.950 768.450 111.000 769.050 ;
        RECT 106.950 766.950 111.450 768.450 ;
        RECT 91.950 760.950 94.050 766.050 ;
        RECT 98.400 762.600 99.450 766.950 ;
        RECT 100.950 763.950 106.050 766.050 ;
        RECT 110.400 763.200 111.450 766.950 ;
        RECT 92.400 760.200 93.600 760.950 ;
        RECT 98.400 760.200 99.600 762.600 ;
        RECT 109.950 761.100 112.050 763.200 ;
        RECT 113.400 762.450 114.450 796.950 ;
        RECT 116.400 796.050 117.450 800.400 ;
        RECT 118.950 796.950 121.050 799.050 ;
        RECT 115.950 793.950 118.050 796.050 ;
        RECT 119.400 790.050 120.450 796.950 ;
        RECT 122.400 796.050 123.450 808.950 ;
        RECT 127.950 806.100 130.050 808.200 ;
        RECT 134.400 807.600 135.450 817.950 ;
        RECT 440.400 817.050 441.450 820.950 ;
        RECT 262.950 814.950 265.050 817.050 ;
        RECT 301.950 814.950 304.050 817.050 ;
        RECT 394.950 814.950 397.050 817.050 ;
        RECT 439.800 814.950 441.900 817.050 ;
        RECT 172.950 811.950 175.050 814.050 ;
        RECT 184.950 811.950 187.050 814.050 ;
        RECT 173.400 807.600 174.450 811.950 ;
        RECT 185.400 808.350 186.450 811.950 ;
        RECT 128.400 805.350 129.600 806.100 ;
        RECT 134.400 805.350 135.600 807.600 ;
        RECT 173.400 805.500 174.600 807.600 ;
        RECT 184.950 806.250 187.050 808.350 ;
        RECT 193.950 806.250 196.050 808.350 ;
        RECT 199.950 806.250 202.050 808.350 ;
        RECT 238.950 806.250 241.050 808.350 ;
        RECT 247.800 806.250 249.900 808.350 ;
        RECT 127.950 802.950 130.050 805.050 ;
        RECT 130.950 802.950 133.050 805.050 ;
        RECT 133.950 802.950 136.050 805.050 ;
        RECT 151.950 802.950 154.050 805.050 ;
        RECT 157.950 802.950 160.050 805.050 ;
        RECT 166.950 803.100 169.050 805.200 ;
        RECT 172.950 803.100 175.050 805.200 ;
        RECT 175.950 803.100 178.050 805.200 ;
        RECT 131.400 800.400 132.600 802.650 ;
        RECT 152.400 801.900 153.600 802.650 ;
        RECT 121.950 793.950 124.050 796.050 ;
        RECT 118.950 787.950 121.050 790.050 ;
        RECT 131.400 777.450 132.450 800.400 ;
        RECT 151.950 799.800 154.050 801.900 ;
        RECT 167.400 800.400 168.600 802.800 ;
        RECT 176.400 800.400 177.600 802.800 ;
        RECT 167.400 799.050 168.450 800.400 ;
        RECT 166.950 796.950 169.050 799.050 ;
        RECT 167.400 790.050 168.450 796.950 ;
        RECT 166.950 787.950 169.050 790.050 ;
        RECT 176.400 784.050 177.450 800.400 ;
        RECT 185.400 799.050 186.450 806.250 ;
        RECT 194.400 805.500 195.600 806.250 ;
        RECT 200.400 805.500 201.600 806.250 ;
        RECT 239.400 805.500 240.600 806.250 ;
        RECT 190.950 803.100 193.050 805.200 ;
        RECT 193.950 803.100 196.050 805.200 ;
        RECT 196.950 803.100 199.050 805.200 ;
        RECT 199.950 803.100 202.050 805.200 ;
        RECT 202.950 803.100 205.050 805.200 ;
        RECT 214.950 802.950 217.050 805.050 ;
        RECT 220.950 802.950 223.050 805.050 ;
        RECT 229.950 803.100 232.050 805.200 ;
        RECT 232.950 803.100 235.050 805.200 ;
        RECT 235.950 803.100 238.050 805.200 ;
        RECT 238.950 803.100 241.050 805.200 ;
        RECT 241.950 803.100 244.050 805.200 ;
        RECT 191.400 800.400 192.600 802.800 ;
        RECT 197.400 800.400 198.600 802.800 ;
        RECT 184.950 796.950 187.050 799.050 ;
        RECT 191.400 790.050 192.450 800.400 ;
        RECT 190.950 787.950 193.050 790.050 ;
        RECT 169.950 781.950 172.050 784.050 ;
        RECT 175.950 781.950 178.050 784.050 ;
        RECT 128.400 776.400 132.450 777.450 ;
        RECT 113.400 761.400 117.450 762.450 ;
        RECT 110.400 760.350 111.600 761.100 ;
        RECT 88.950 757.800 91.050 759.900 ;
        RECT 91.950 757.800 94.050 759.900 ;
        RECT 94.950 757.800 97.050 759.900 ;
        RECT 97.950 757.800 100.050 759.900 ;
        RECT 106.950 757.950 109.050 760.050 ;
        RECT 109.950 757.950 112.050 760.050 ;
        RECT 74.400 748.050 75.450 755.400 ;
        RECT 79.950 754.950 82.050 757.050 ;
        RECT 82.950 754.950 85.050 757.050 ;
        RECT 89.400 755.400 90.600 757.500 ;
        RECT 95.400 755.400 96.600 757.500 ;
        RECT 103.950 756.450 106.050 757.050 ;
        RECT 107.400 756.450 108.600 757.650 ;
        RECT 103.950 755.400 108.600 756.450 ;
        RECT 73.950 745.950 76.050 748.050 ;
        RECT 80.400 736.050 81.450 754.950 ;
        RECT 89.400 739.050 90.450 755.400 ;
        RECT 95.400 748.050 96.450 755.400 ;
        RECT 103.950 754.950 106.050 755.400 ;
        RECT 94.950 745.950 97.050 748.050 ;
        RECT 104.400 745.050 105.450 754.950 ;
        RECT 116.400 754.050 117.450 761.400 ;
        RECT 121.950 760.950 124.050 763.050 ;
        RECT 128.400 762.600 129.450 776.400 ;
        RECT 145.950 775.950 148.050 778.050 ;
        RECT 146.400 769.050 147.450 775.950 ;
        RECT 145.950 766.950 148.050 769.050 ;
        RECT 136.800 763.950 138.900 766.050 ;
        RECT 122.400 760.200 123.600 760.950 ;
        RECT 128.400 760.200 129.600 762.600 ;
        RECT 121.950 757.800 124.050 759.900 ;
        RECT 124.950 757.800 127.050 759.900 ;
        RECT 127.950 757.800 130.050 759.900 ;
        RECT 130.950 757.800 133.050 759.900 ;
        RECT 125.400 755.400 126.600 757.500 ;
        RECT 131.400 757.050 132.600 757.500 ;
        RECT 137.400 757.050 138.450 763.950 ;
        RECT 139.950 760.950 142.050 766.050 ;
        RECT 143.400 762.450 144.600 762.600 ;
        RECT 146.400 762.450 147.450 766.950 ;
        RECT 143.400 761.400 147.450 762.450 ;
        RECT 143.400 760.200 144.600 761.400 ;
        RECT 151.950 760.950 154.050 763.050 ;
        RECT 163.950 760.950 166.050 763.050 ;
        RECT 170.400 762.600 171.450 781.950 ;
        RECT 178.950 778.950 181.050 781.050 ;
        RECT 175.950 769.950 178.050 772.050 ;
        RECT 152.400 760.200 153.600 760.950 ;
        RECT 164.400 760.200 165.600 760.950 ;
        RECT 170.400 760.200 171.600 762.600 ;
        RECT 142.950 757.800 145.050 759.900 ;
        RECT 148.950 757.800 151.050 759.900 ;
        RECT 151.950 757.800 154.050 759.900 ;
        RECT 163.950 757.800 166.050 759.900 ;
        RECT 166.950 757.800 169.050 759.900 ;
        RECT 169.950 757.800 172.050 759.900 ;
        RECT 131.400 755.400 136.050 757.050 ;
        RECT 106.950 751.950 109.050 754.050 ;
        RECT 115.950 751.950 118.050 754.050 ;
        RECT 103.950 742.950 106.050 745.050 ;
        RECT 88.950 736.950 91.050 739.050 ;
        RECT 70.950 733.950 73.050 736.050 ;
        RECT 79.950 733.950 82.050 736.050 ;
        RECT 61.950 730.950 64.050 733.050 ;
        RECT 67.950 730.950 70.050 733.050 ;
        RECT 53.400 727.500 54.600 729.600 ;
        RECT 59.400 727.500 60.600 729.600 ;
        RECT 52.950 725.100 55.050 727.200 ;
        RECT 55.950 725.100 58.050 727.200 ;
        RECT 58.950 725.100 61.050 727.200 ;
        RECT 61.950 725.100 64.050 727.200 ;
        RECT 52.950 721.950 55.050 724.050 ;
        RECT 56.400 722.400 57.600 724.800 ;
        RECT 62.400 724.050 63.600 724.800 ;
        RECT 46.950 715.950 49.050 718.050 ;
        RECT 43.950 712.950 46.050 715.050 ;
        RECT 40.950 688.950 43.050 691.050 ;
        RECT 53.400 688.050 54.450 721.950 ;
        RECT 56.400 715.050 57.450 722.400 ;
        RECT 61.950 721.950 64.050 724.050 ;
        RECT 55.950 712.950 58.050 715.050 ;
        RECT 68.400 700.050 69.450 730.950 ;
        RECT 71.400 730.050 72.450 733.950 ;
        RECT 80.400 730.350 81.450 733.950 ;
        RECT 70.950 727.950 73.050 730.050 ;
        RECT 73.950 728.250 76.050 730.350 ;
        RECT 79.950 728.250 82.050 730.350 ;
        RECT 94.950 728.250 97.050 730.350 ;
        RECT 102.000 729.600 106.050 730.050 ;
        RECT 74.400 727.500 75.600 728.250 ;
        RECT 80.400 727.500 81.600 728.250 ;
        RECT 95.400 727.500 96.600 728.250 ;
        RECT 101.400 727.950 106.050 729.600 ;
        RECT 101.400 727.500 102.600 727.950 ;
        RECT 73.950 725.100 76.050 727.200 ;
        RECT 76.950 725.100 79.050 727.200 ;
        RECT 79.950 725.100 82.050 727.200 ;
        RECT 82.950 725.100 85.050 727.200 ;
        RECT 91.950 725.100 94.050 727.200 ;
        RECT 94.950 725.100 97.050 727.200 ;
        RECT 97.950 725.100 100.050 727.200 ;
        RECT 100.950 725.100 103.050 727.200 ;
        RECT 73.950 721.950 76.050 724.050 ;
        RECT 77.400 722.400 78.600 724.800 ;
        RECT 83.400 723.000 84.600 724.800 ;
        RECT 70.950 715.950 73.050 718.050 ;
        RECT 71.400 711.450 72.450 715.950 ;
        RECT 74.400 715.050 75.450 721.950 ;
        RECT 77.400 718.050 78.450 722.400 ;
        RECT 82.950 718.950 85.050 723.000 ;
        RECT 88.950 721.800 91.050 723.900 ;
        RECT 92.400 722.400 93.600 724.800 ;
        RECT 98.400 723.000 99.600 724.800 ;
        RECT 76.950 715.950 79.050 718.050 ;
        RECT 73.950 712.950 76.050 715.050 ;
        RECT 77.400 711.450 78.450 715.950 ;
        RECT 71.400 710.400 78.450 711.450 ;
        RECT 89.400 700.050 90.450 721.800 ;
        RECT 92.400 718.050 93.450 722.400 ;
        RECT 97.950 718.950 100.050 723.000 ;
        RECT 91.950 715.950 94.050 718.050 ;
        RECT 97.950 715.800 100.050 717.900 ;
        RECT 58.950 697.950 61.050 700.050 ;
        RECT 67.950 697.950 70.050 700.050 ;
        RECT 88.950 697.950 91.050 700.050 ;
        RECT 52.950 685.950 55.050 688.050 ;
        RECT 35.400 682.200 36.600 684.600 ;
        RECT 49.950 683.100 52.050 685.200 ;
        RECT 50.400 682.350 51.600 683.100 ;
        RECT 25.950 679.800 28.050 681.900 ;
        RECT 28.950 679.800 31.050 681.900 ;
        RECT 31.950 679.800 34.050 681.900 ;
        RECT 34.950 679.800 37.050 681.900 ;
        RECT 37.950 679.800 40.050 681.900 ;
        RECT 46.950 679.950 49.050 682.050 ;
        RECT 49.950 679.950 52.050 682.050 ;
        RECT 52.950 679.950 55.050 682.050 ;
        RECT 26.400 678.450 27.600 679.500 ;
        RECT 32.400 678.750 33.600 679.500 ;
        RECT 38.400 678.750 39.600 679.500 ;
        RECT 47.400 678.900 48.600 679.650 ;
        RECT 23.400 677.400 27.600 678.450 ;
        RECT 19.950 667.950 22.050 670.050 ;
        RECT 13.950 655.950 16.050 658.050 ;
        RECT 23.400 655.050 24.450 677.400 ;
        RECT 31.950 676.650 34.050 678.750 ;
        RECT 37.950 676.650 40.050 678.750 ;
        RECT 46.950 676.800 49.050 678.900 ;
        RECT 53.400 678.000 54.600 679.650 ;
        RECT 47.400 667.050 48.450 676.800 ;
        RECT 52.950 673.950 55.050 678.000 ;
        RECT 55.950 676.950 58.050 679.050 ;
        RECT 46.950 664.950 49.050 667.050 ;
        RECT 34.950 655.950 37.050 658.050 ;
        RECT 43.950 655.950 46.050 658.050 ;
        RECT 13.950 650.100 16.050 654.900 ;
        RECT 22.950 652.950 25.050 655.050 ;
        RECT 14.400 649.350 15.600 650.100 ;
        RECT 19.950 649.950 22.050 652.050 ;
        RECT 28.950 650.100 31.050 652.200 ;
        RECT 35.400 651.600 36.450 655.950 ;
        RECT 44.400 651.600 45.450 655.950 ;
        RECT 56.400 655.050 57.450 676.950 ;
        RECT 59.400 676.050 60.450 697.950 ;
        RECT 67.950 691.950 70.050 694.050 ;
        RECT 85.950 691.950 88.050 694.050 ;
        RECT 68.400 684.600 69.450 691.950 ;
        RECT 68.400 682.350 69.600 684.600 ;
        RECT 73.950 682.950 76.050 685.050 ;
        RECT 79.950 682.950 82.050 685.050 ;
        RECT 86.400 684.600 87.450 691.950 ;
        RECT 91.950 688.950 94.050 691.050 ;
        RECT 92.400 685.050 93.450 688.950 ;
        RECT 94.950 685.950 97.050 688.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 67.950 679.950 70.050 682.050 ;
        RECT 61.950 676.950 64.050 679.050 ;
        RECT 65.400 677.400 66.600 679.650 ;
        RECT 58.950 673.950 61.050 676.050 ;
        RECT 58.950 667.950 61.050 670.050 ;
        RECT 55.950 652.950 58.050 655.050 ;
        RECT 10.950 646.950 13.050 649.050 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 11.400 644.400 12.600 646.650 ;
        RECT 11.400 640.050 12.450 644.400 ;
        RECT 10.950 637.950 13.050 640.050 ;
        RECT 1.950 616.950 4.050 619.050 ;
        RECT 20.400 610.050 21.450 649.950 ;
        RECT 29.400 649.350 30.600 650.100 ;
        RECT 35.400 649.350 36.600 651.600 ;
        RECT 44.400 649.350 45.600 651.600 ;
        RECT 49.950 650.100 52.050 652.200 ;
        RECT 50.400 649.350 51.600 650.100 ;
        RECT 25.950 646.950 28.050 649.050 ;
        RECT 28.950 646.950 31.050 649.050 ;
        RECT 31.950 646.950 34.050 649.050 ;
        RECT 34.950 646.950 37.050 649.050 ;
        RECT 43.950 646.950 46.050 649.050 ;
        RECT 46.950 646.950 49.050 649.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 52.950 646.950 55.050 649.050 ;
        RECT 26.400 644.400 27.600 646.650 ;
        RECT 32.400 645.900 33.600 646.650 ;
        RECT 47.400 645.900 48.600 646.650 ;
        RECT 26.400 640.050 27.450 644.400 ;
        RECT 31.950 643.800 34.050 645.900 ;
        RECT 46.950 643.800 49.050 645.900 ;
        RECT 53.400 644.400 54.600 646.650 ;
        RECT 53.400 643.050 54.450 644.400 ;
        RECT 55.950 643.950 58.050 646.050 ;
        RECT 52.950 640.950 55.050 643.050 ;
        RECT 25.950 637.950 28.050 640.050 ;
        RECT 26.400 622.050 27.450 637.950 ;
        RECT 53.400 637.050 54.450 640.950 ;
        RECT 52.950 634.950 55.050 637.050 ;
        RECT 25.950 619.950 28.050 622.050 ;
        RECT 56.400 612.450 57.450 643.950 ;
        RECT 53.400 611.400 57.450 612.450 ;
        RECT 13.950 606.000 16.050 610.050 ;
        RECT 19.950 607.950 22.050 610.050 ;
        RECT 14.400 604.200 15.600 606.000 ;
        RECT 19.950 604.800 22.050 606.900 ;
        RECT 28.950 606.000 31.050 610.050 ;
        RECT 20.400 604.200 21.600 604.800 ;
        RECT 29.400 604.200 30.600 606.000 ;
        RECT 34.950 604.950 37.050 610.050 ;
        RECT 53.400 607.050 54.450 611.400 ;
        RECT 43.950 604.950 46.050 607.050 ;
        RECT 52.950 604.950 55.050 607.050 ;
        RECT 55.950 606.000 58.050 610.050 ;
        RECT 59.400 607.050 60.450 667.950 ;
        RECT 62.400 652.050 63.450 676.950 ;
        RECT 65.400 658.050 66.450 677.400 ;
        RECT 74.400 676.050 75.450 682.950 ;
        RECT 80.400 682.200 81.600 682.950 ;
        RECT 86.400 682.200 87.600 684.600 ;
        RECT 91.950 682.950 94.050 685.050 ;
        RECT 79.950 679.800 82.050 681.900 ;
        RECT 82.950 679.800 85.050 681.900 ;
        RECT 85.950 679.800 88.050 681.900 ;
        RECT 88.950 679.800 91.050 681.900 ;
        RECT 83.400 678.750 84.600 679.500 ;
        RECT 89.400 678.750 90.600 679.500 ;
        RECT 95.400 678.750 96.450 685.950 ;
        RECT 82.950 676.650 85.050 678.750 ;
        RECT 88.950 676.650 91.050 678.750 ;
        RECT 94.950 676.650 97.050 678.750 ;
        RECT 67.950 673.950 70.050 676.050 ;
        RECT 73.950 673.950 76.050 676.050 ;
        RECT 64.950 655.950 67.050 658.050 ;
        RECT 68.400 652.350 69.450 673.950 ;
        RECT 79.950 664.950 82.050 667.050 ;
        RECT 76.950 655.950 79.050 658.050 ;
        RECT 61.950 649.950 64.050 652.050 ;
        RECT 67.950 650.250 70.050 652.350 ;
        RECT 73.950 650.250 76.050 652.350 ;
        RECT 77.400 652.050 78.450 655.950 ;
        RECT 68.400 649.500 69.600 650.250 ;
        RECT 74.400 649.500 75.600 650.250 ;
        RECT 76.950 649.950 79.050 652.050 ;
        RECT 64.950 647.100 67.050 649.200 ;
        RECT 67.950 647.100 70.050 649.200 ;
        RECT 70.950 647.100 73.050 649.200 ;
        RECT 73.950 647.100 76.050 649.200 ;
        RECT 65.400 644.400 66.600 646.800 ;
        RECT 71.400 645.000 72.600 646.800 ;
        RECT 61.950 634.950 64.050 637.050 ;
        RECT 35.400 604.200 36.600 604.950 ;
        RECT 10.950 601.800 13.050 603.900 ;
        RECT 13.950 601.800 16.050 603.900 ;
        RECT 16.950 601.800 19.050 603.900 ;
        RECT 19.950 601.800 22.050 603.900 ;
        RECT 28.950 601.800 31.050 603.900 ;
        RECT 31.950 601.800 34.050 603.900 ;
        RECT 34.950 601.800 37.050 603.900 ;
        RECT 37.950 601.800 40.050 603.900 ;
        RECT 11.400 599.400 12.600 601.500 ;
        RECT 17.400 600.750 18.600 601.500 ;
        RECT 32.400 600.750 33.600 601.500 ;
        RECT 11.400 586.050 12.450 599.400 ;
        RECT 16.950 598.650 19.050 600.750 ;
        RECT 31.950 595.950 34.050 600.750 ;
        RECT 38.400 599.400 39.600 601.500 ;
        RECT 31.950 586.950 34.050 589.050 ;
        RECT 10.950 583.950 13.050 586.050 ;
        RECT 19.950 583.950 22.050 586.050 ;
        RECT 1.950 577.950 4.050 580.050 ;
        RECT 13.950 577.950 16.050 580.050 ;
        RECT 2.400 562.050 3.450 577.950 ;
        RECT 4.950 574.950 7.050 577.050 ;
        RECT 5.400 568.050 6.450 574.950 ;
        RECT 14.400 573.600 15.450 577.950 ;
        RECT 20.400 574.050 21.450 583.950 ;
        RECT 14.400 571.350 15.600 573.600 ;
        RECT 19.950 571.950 22.050 574.050 ;
        RECT 25.950 573.000 28.050 577.050 ;
        RECT 32.400 573.600 33.450 586.950 ;
        RECT 26.400 571.500 27.600 573.000 ;
        RECT 32.400 571.500 33.600 573.600 ;
        RECT 10.950 568.950 13.050 571.050 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 22.950 569.100 25.050 571.200 ;
        RECT 25.950 569.100 28.050 571.200 ;
        RECT 28.950 569.100 31.050 571.200 ;
        RECT 31.950 569.100 34.050 571.200 ;
        RECT 4.950 565.950 7.050 568.050 ;
        RECT 11.400 567.900 12.600 568.650 ;
        RECT 23.400 568.050 24.600 568.800 ;
        RECT 29.400 568.050 30.600 568.800 ;
        RECT 38.400 568.050 39.450 599.400 ;
        RECT 44.400 585.450 45.450 604.950 ;
        RECT 56.400 604.200 57.600 606.000 ;
        RECT 58.950 604.950 61.050 607.050 ;
        RECT 62.400 606.600 63.450 634.950 ;
        RECT 65.400 634.050 66.450 644.400 ;
        RECT 70.950 640.950 73.050 645.000 ;
        RECT 76.950 643.950 79.050 646.050 ;
        RECT 77.400 634.050 78.450 643.950 ;
        RECT 64.950 631.950 67.050 634.050 ;
        RECT 76.950 631.950 79.050 634.050 ;
        RECT 70.950 619.950 73.050 622.050 ;
        RECT 71.400 606.600 72.450 619.950 ;
        RECT 76.950 610.950 79.050 613.050 ;
        RECT 77.400 606.600 78.450 610.950 ;
        RECT 80.400 607.050 81.450 664.950 ;
        RECT 98.400 658.050 99.450 715.800 ;
        RECT 107.400 691.050 108.450 751.950 ;
        RECT 125.400 748.050 126.450 755.400 ;
        RECT 132.000 754.950 136.050 755.400 ;
        RECT 136.950 754.950 139.050 757.050 ;
        RECT 149.400 756.000 150.600 757.500 ;
        RECT 148.950 751.950 151.050 756.000 ;
        RECT 154.950 754.950 157.050 757.050 ;
        RECT 160.950 754.950 163.050 757.050 ;
        RECT 167.400 755.400 168.600 757.500 ;
        RECT 155.400 748.050 156.450 754.950 ;
        RECT 124.950 745.950 127.050 748.050 ;
        RECT 154.950 745.950 157.050 748.050 ;
        RECT 118.950 742.950 121.050 745.050 ;
        RECT 119.400 736.050 120.450 742.950 ;
        RECT 125.400 742.050 126.450 745.950 ;
        RECT 124.950 739.950 127.050 742.050 ;
        RECT 139.950 739.950 142.050 742.050 ;
        RECT 118.950 733.950 121.050 736.050 ;
        RECT 109.950 727.950 112.050 730.050 ;
        RECT 118.950 728.100 121.050 730.200 ;
        RECT 124.950 728.100 127.050 730.200 ;
        RECT 110.400 700.050 111.450 727.950 ;
        RECT 119.400 727.350 120.600 728.100 ;
        RECT 125.400 727.350 126.600 728.100 ;
        RECT 130.950 727.950 133.050 730.050 ;
        RECT 140.400 729.600 141.450 739.950 ;
        RECT 157.950 733.950 160.050 736.050 ;
        RECT 115.950 724.950 118.050 727.050 ;
        RECT 118.950 724.950 121.050 727.050 ;
        RECT 121.950 724.950 124.050 727.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 112.950 721.950 115.050 724.050 ;
        RECT 116.400 722.400 117.600 724.650 ;
        RECT 122.400 722.400 123.600 724.650 ;
        RECT 113.400 715.050 114.450 721.950 ;
        RECT 116.400 718.050 117.450 722.400 ;
        RECT 115.950 715.950 118.050 718.050 ;
        RECT 122.400 715.050 123.450 722.400 ;
        RECT 112.950 712.950 115.050 715.050 ;
        RECT 121.950 712.950 124.050 715.050 ;
        RECT 131.400 709.050 132.450 727.950 ;
        RECT 140.400 727.350 141.600 729.600 ;
        RECT 145.950 728.100 148.050 730.200 ;
        RECT 158.400 729.600 159.450 733.950 ;
        RECT 161.400 732.450 162.450 754.950 ;
        RECT 167.400 751.050 168.450 755.400 ;
        RECT 166.950 748.950 169.050 751.050 ;
        RECT 161.400 732.000 165.450 732.450 ;
        RECT 161.400 731.400 166.050 732.000 ;
        RECT 146.400 727.350 147.600 728.100 ;
        RECT 158.400 727.500 159.600 729.600 ;
        RECT 163.950 727.950 166.050 731.400 ;
        RECT 176.400 730.050 177.450 769.950 ;
        RECT 179.400 766.050 180.450 778.950 ;
        RECT 191.400 778.050 192.450 787.950 ;
        RECT 190.950 775.950 193.050 778.050 ;
        RECT 197.400 769.050 198.450 800.400 ;
        RECT 199.950 799.950 202.050 802.050 ;
        RECT 203.400 800.400 204.600 802.800 ;
        RECT 215.400 801.000 216.600 802.650 ;
        RECT 200.400 790.050 201.450 799.950 ;
        RECT 199.950 787.950 202.050 790.050 ;
        RECT 203.400 772.050 204.450 800.400 ;
        RECT 214.950 796.950 217.050 801.000 ;
        RECT 230.400 800.400 231.600 802.800 ;
        RECT 236.400 800.400 237.600 802.800 ;
        RECT 242.400 802.050 243.600 802.800 ;
        RECT 211.950 784.950 214.050 787.050 ;
        RECT 202.950 769.950 205.050 772.050 ;
        RECT 184.950 766.950 187.050 769.050 ;
        RECT 196.950 766.950 199.050 769.050 ;
        RECT 178.950 763.950 181.050 766.050 ;
        RECT 185.400 762.600 186.450 766.950 ;
        RECT 185.400 760.350 186.600 762.600 ;
        RECT 190.950 761.100 193.050 763.200 ;
        RECT 191.400 760.350 192.600 761.100 ;
        RECT 196.950 760.950 199.050 763.050 ;
        RECT 205.950 761.100 208.050 763.200 ;
        RECT 212.400 762.600 213.450 784.950 ;
        RECT 226.950 778.950 229.050 781.050 ;
        RECT 227.400 763.200 228.450 778.950 ;
        RECT 230.400 772.050 231.450 800.400 ;
        RECT 236.400 787.050 237.450 800.400 ;
        RECT 241.950 799.950 244.050 802.050 ;
        RECT 248.400 793.050 249.450 806.250 ;
        RECT 250.950 805.950 253.050 808.050 ;
        RECT 256.950 806.250 259.050 808.350 ;
        RECT 263.400 807.600 264.450 814.950 ;
        RECT 277.950 811.950 280.050 814.050 ;
        RECT 278.400 808.350 279.450 811.950 ;
        RECT 302.400 808.350 303.450 814.950 ;
        RECT 247.950 790.950 250.050 793.050 ;
        RECT 235.950 784.950 238.050 787.050 ;
        RECT 229.950 769.950 232.050 772.050 ;
        RECT 236.400 765.450 237.450 784.950 ;
        RECT 251.400 766.050 252.450 805.950 ;
        RECT 257.400 805.500 258.600 806.250 ;
        RECT 263.400 805.500 264.600 807.600 ;
        RECT 277.950 806.250 280.050 808.350 ;
        RECT 295.950 806.250 298.050 808.350 ;
        RECT 301.950 806.250 304.050 808.350 ;
        RECT 278.400 805.500 279.600 806.250 ;
        RECT 296.400 805.500 297.600 806.250 ;
        RECT 302.400 805.500 303.600 806.250 ;
        RECT 313.950 805.950 316.050 808.050 ;
        RECT 322.950 806.100 325.050 808.200 ;
        RECT 334.950 806.250 337.050 808.350 ;
        RECT 343.950 806.250 346.050 808.350 ;
        RECT 364.950 806.250 367.050 808.350 ;
        RECT 373.950 806.250 376.050 808.350 ;
        RECT 256.950 803.100 259.050 805.200 ;
        RECT 259.950 803.100 262.050 805.200 ;
        RECT 262.950 803.100 265.050 805.200 ;
        RECT 265.950 803.100 268.050 805.200 ;
        RECT 274.950 803.100 277.050 805.200 ;
        RECT 277.950 803.100 280.050 805.200 ;
        RECT 280.950 803.100 283.050 805.200 ;
        RECT 286.950 802.950 289.050 805.050 ;
        RECT 292.950 803.100 295.050 805.200 ;
        RECT 295.950 803.100 298.050 805.200 ;
        RECT 298.950 803.100 301.050 805.200 ;
        RECT 301.950 803.100 304.050 805.200 ;
        RECT 304.950 803.100 307.050 805.200 ;
        RECT 260.400 802.050 261.600 802.800 ;
        RECT 259.950 799.950 262.050 802.050 ;
        RECT 266.400 800.400 267.600 802.800 ;
        RECT 275.400 800.400 276.600 802.800 ;
        RECT 281.400 802.050 282.600 802.800 ;
        RECT 266.400 793.050 267.450 800.400 ;
        RECT 265.950 790.950 268.050 793.050 ;
        RECT 275.400 787.050 276.450 800.400 ;
        RECT 280.950 799.950 283.050 802.050 ;
        RECT 280.950 796.800 283.050 798.900 ;
        RECT 274.950 784.950 277.050 787.050 ;
        RECT 233.400 764.400 237.450 765.450 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 190.950 757.950 193.050 760.050 ;
        RECT 182.400 755.400 183.600 757.650 ;
        RECT 188.400 756.900 189.600 757.650 ;
        RECT 182.400 736.050 183.450 755.400 ;
        RECT 187.950 754.800 190.050 756.900 ;
        RECT 197.400 751.050 198.450 760.950 ;
        RECT 206.400 760.350 207.600 761.100 ;
        RECT 212.400 760.350 213.600 762.600 ;
        RECT 226.950 761.100 229.050 763.200 ;
        RECT 233.400 762.600 234.450 764.400 ;
        RECT 250.950 763.950 253.050 766.050 ;
        RECT 227.400 760.350 228.600 761.100 ;
        RECT 233.400 760.350 234.600 762.600 ;
        RECT 250.950 760.800 253.050 762.900 ;
        RECT 256.950 760.950 259.050 763.050 ;
        RECT 265.950 760.950 268.050 763.050 ;
        RECT 271.950 762.000 274.050 766.050 ;
        RECT 251.400 760.200 252.600 760.800 ;
        RECT 257.400 760.200 258.600 760.950 ;
        RECT 266.400 760.200 267.600 760.950 ;
        RECT 272.400 760.200 273.600 762.000 ;
        RECT 205.950 757.950 208.050 760.050 ;
        RECT 208.950 757.950 211.050 760.050 ;
        RECT 211.950 757.950 214.050 760.050 ;
        RECT 214.950 757.950 217.050 760.050 ;
        RECT 226.950 757.950 229.050 760.050 ;
        RECT 229.950 757.950 232.050 760.050 ;
        RECT 232.950 757.950 235.050 760.050 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 247.950 757.800 250.050 759.900 ;
        RECT 250.950 757.800 253.050 759.900 ;
        RECT 253.950 757.800 256.050 759.900 ;
        RECT 256.950 757.800 259.050 759.900 ;
        RECT 265.950 757.800 268.050 759.900 ;
        RECT 268.950 757.800 271.050 759.900 ;
        RECT 271.950 757.800 274.050 759.900 ;
        RECT 274.950 757.800 277.050 759.900 ;
        RECT 209.400 755.400 210.600 757.650 ;
        RECT 215.400 755.400 216.600 757.650 ;
        RECT 230.400 755.400 231.600 757.650 ;
        RECT 236.400 755.400 237.600 757.650 ;
        RECT 196.950 748.950 199.050 751.050 ;
        RECT 181.950 733.950 184.050 736.050 ;
        RECT 166.950 727.950 169.050 730.050 ;
        RECT 175.950 727.950 178.050 730.050 ;
        RECT 193.950 728.250 196.050 730.350 ;
        RECT 200.400 729.450 201.600 729.600 ;
        RECT 200.400 728.400 207.450 729.450 ;
        RECT 136.950 724.950 139.050 727.050 ;
        RECT 139.950 724.950 142.050 727.050 ;
        RECT 142.950 724.950 145.050 727.050 ;
        RECT 145.950 724.950 148.050 727.050 ;
        RECT 154.950 725.100 157.050 727.200 ;
        RECT 157.950 725.100 160.050 727.200 ;
        RECT 160.950 725.100 163.050 727.200 ;
        RECT 137.400 723.900 138.600 724.650 ;
        RECT 136.950 721.800 139.050 723.900 ;
        RECT 143.400 722.400 144.600 724.650 ;
        RECT 155.400 722.400 156.600 724.800 ;
        RECT 143.400 718.050 144.450 722.400 ;
        RECT 145.950 718.950 148.050 721.050 ;
        RECT 142.950 715.950 145.050 718.050 ;
        RECT 146.400 712.050 147.450 718.950 ;
        RECT 148.950 715.950 151.050 718.050 ;
        RECT 145.950 709.950 148.050 712.050 ;
        RECT 130.950 706.950 133.050 709.050 ;
        RECT 139.950 706.950 142.050 709.050 ;
        RECT 112.950 703.950 115.050 706.050 ;
        RECT 109.950 697.950 112.050 700.050 ;
        RECT 113.400 697.050 114.450 703.950 ;
        RECT 118.950 700.950 121.050 703.050 ;
        RECT 112.950 694.950 115.050 697.050 ;
        RECT 100.950 688.950 103.050 691.050 ;
        RECT 106.800 688.950 108.900 691.050 ;
        RECT 101.400 685.050 102.450 688.950 ;
        RECT 103.950 687.600 106.050 688.050 ;
        RECT 109.950 687.600 112.050 691.050 ;
        RECT 103.950 687.000 112.050 687.600 ;
        RECT 103.950 686.550 111.450 687.000 ;
        RECT 103.950 685.950 106.050 686.550 ;
        RECT 100.800 682.950 102.900 685.050 ;
        RECT 103.950 682.800 106.050 684.900 ;
        RECT 109.950 682.950 112.050 685.050 ;
        RECT 119.400 684.600 120.450 700.950 ;
        RECT 124.950 694.950 127.050 697.050 ;
        RECT 125.400 684.600 126.450 694.950 ;
        RECT 131.400 688.050 132.450 706.950 ;
        RECT 130.950 685.950 133.050 688.050 ;
        RECT 136.950 685.950 139.050 688.050 ;
        RECT 127.950 684.900 132.000 685.050 ;
        RECT 104.400 682.200 105.600 682.800 ;
        RECT 110.400 682.200 111.600 682.950 ;
        RECT 119.400 682.200 120.600 684.600 ;
        RECT 125.400 682.200 126.600 684.600 ;
        RECT 127.950 682.950 133.050 684.900 ;
        RECT 130.950 682.800 133.050 682.950 ;
        RECT 131.400 682.200 132.600 682.800 ;
        RECT 103.950 679.800 106.050 681.900 ;
        RECT 106.950 679.800 109.050 681.900 ;
        RECT 109.950 679.800 112.050 681.900 ;
        RECT 118.950 679.800 121.050 681.900 ;
        RECT 121.950 679.800 124.050 681.900 ;
        RECT 124.950 679.800 127.050 681.900 ;
        RECT 127.950 679.800 130.050 681.900 ;
        RECT 130.950 679.800 133.050 681.900 ;
        RECT 100.950 676.950 103.050 679.050 ;
        RECT 107.400 677.400 108.600 679.500 ;
        RECT 88.950 655.950 91.050 658.050 ;
        RECT 97.950 655.950 100.050 658.050 ;
        RECT 89.400 651.600 90.450 655.950 ;
        RECT 101.400 655.050 102.450 676.950 ;
        RECT 107.400 667.050 108.450 677.400 ;
        RECT 115.950 676.950 118.050 679.050 ;
        RECT 122.400 678.750 123.600 679.500 ;
        RECT 116.400 670.050 117.450 676.950 ;
        RECT 121.950 676.650 124.050 678.750 ;
        RECT 128.400 677.400 129.600 679.500 ;
        RECT 122.400 673.050 123.450 676.650 ;
        RECT 121.950 670.950 124.050 673.050 ;
        RECT 128.400 670.050 129.450 677.400 ;
        RECT 115.950 667.950 118.050 670.050 ;
        RECT 127.950 667.950 130.050 670.050 ;
        RECT 106.950 664.950 109.050 667.050 ;
        RECT 100.950 652.950 103.050 655.050 ;
        RECT 96.000 651.600 100.050 652.050 ;
        RECT 89.400 649.500 90.600 651.600 ;
        RECT 95.400 649.950 100.050 651.600 ;
        RECT 95.400 649.500 96.600 649.950 ;
        RECT 100.950 649.800 103.050 651.900 ;
        RECT 103.950 649.950 106.050 652.050 ;
        RECT 106.950 649.950 109.050 655.050 ;
        RECT 137.400 652.350 138.450 685.950 ;
        RECT 140.400 685.050 141.450 706.950 ;
        RECT 139.950 682.950 142.050 685.050 ;
        RECT 145.800 683.100 147.900 685.200 ;
        RECT 149.400 685.050 150.450 715.950 ;
        RECT 155.400 709.050 156.450 722.400 ;
        RECT 154.950 706.950 157.050 709.050 ;
        RECT 167.400 703.050 168.450 727.950 ;
        RECT 194.400 727.500 195.600 728.250 ;
        RECT 200.400 727.500 201.600 728.400 ;
        RECT 172.950 724.950 175.050 727.050 ;
        RECT 178.950 724.950 181.050 727.050 ;
        RECT 190.950 725.100 193.050 727.200 ;
        RECT 193.950 725.100 196.050 727.200 ;
        RECT 196.950 725.100 199.050 727.200 ;
        RECT 199.950 725.100 202.050 727.200 ;
        RECT 169.950 721.950 172.050 724.050 ;
        RECT 179.400 722.400 180.600 724.650 ;
        RECT 166.950 700.950 169.050 703.050 ;
        RECT 166.950 688.950 169.050 691.050 ;
        RECT 140.400 663.450 141.450 682.950 ;
        RECT 146.400 682.350 147.600 683.100 ;
        RECT 148.950 682.950 151.050 685.050 ;
        RECT 167.400 684.600 168.450 688.950 ;
        RECT 170.400 685.050 171.450 721.950 ;
        RECT 179.400 694.050 180.450 722.400 ;
        RECT 187.950 721.950 190.050 724.050 ;
        RECT 191.400 722.400 192.600 724.800 ;
        RECT 197.400 722.400 198.600 724.800 ;
        RECT 178.950 691.950 181.050 694.050 ;
        RECT 188.400 688.050 189.450 721.950 ;
        RECT 191.400 706.050 192.450 722.400 ;
        RECT 190.950 703.950 193.050 706.050 ;
        RECT 167.400 682.200 168.600 684.600 ;
        RECT 169.950 682.950 172.050 685.050 ;
        RECT 172.950 682.950 175.050 685.050 ;
        RECT 181.950 682.950 184.050 688.050 ;
        RECT 187.950 685.950 190.050 688.050 ;
        RECT 184.950 684.600 189.000 685.050 ;
        RECT 184.950 684.450 189.600 684.600 ;
        RECT 191.400 684.450 192.450 703.950 ;
        RECT 197.400 700.050 198.450 722.400 ;
        RECT 196.950 697.950 199.050 700.050 ;
        RECT 196.950 691.950 199.050 694.050 ;
        RECT 184.950 683.400 192.450 684.450 ;
        RECT 184.950 682.950 189.600 683.400 ;
        RECT 173.400 682.200 174.600 682.950 ;
        RECT 182.400 682.200 183.600 682.950 ;
        RECT 188.400 682.200 189.600 682.950 ;
        RECT 145.950 679.950 148.050 682.050 ;
        RECT 151.950 679.950 154.050 682.050 ;
        RECT 163.950 679.800 166.050 681.900 ;
        RECT 166.950 679.800 169.050 681.900 ;
        RECT 169.950 679.800 172.050 681.900 ;
        RECT 172.950 679.800 175.050 681.900 ;
        RECT 181.950 679.800 184.050 681.900 ;
        RECT 184.950 679.800 187.050 681.900 ;
        RECT 187.950 679.800 190.050 681.900 ;
        RECT 190.950 679.800 193.050 681.900 ;
        RECT 148.950 676.950 151.050 679.050 ;
        RECT 164.400 677.400 165.600 679.500 ;
        RECT 170.400 678.750 171.600 679.500 ;
        RECT 145.950 670.950 148.050 673.050 ;
        RECT 140.400 662.400 144.450 663.450 ;
        RECT 139.950 658.950 142.050 661.050 ;
        RECT 112.950 650.250 115.050 652.350 ;
        RECT 130.950 650.250 133.050 652.350 ;
        RECT 136.950 650.250 139.050 652.350 ;
        RECT 85.950 647.100 88.050 649.200 ;
        RECT 88.950 647.100 91.050 649.200 ;
        RECT 91.950 647.100 94.050 649.200 ;
        RECT 94.950 647.100 97.050 649.200 ;
        RECT 86.400 645.000 87.600 646.800 ;
        RECT 92.400 646.050 93.600 646.800 ;
        RECT 85.950 640.950 88.050 645.000 ;
        RECT 91.950 643.950 94.050 646.050 ;
        RECT 91.950 616.950 94.050 619.050 ;
        RECT 82.950 610.950 88.050 613.050 ;
        RECT 92.400 610.050 93.450 616.950 ;
        RECT 94.950 610.950 97.050 613.050 ;
        RECT 85.950 607.800 88.050 609.900 ;
        RECT 91.950 607.950 94.050 610.050 ;
        RECT 62.400 604.200 63.600 606.600 ;
        RECT 71.400 604.200 72.600 606.600 ;
        RECT 77.400 604.200 78.600 606.600 ;
        RECT 79.950 604.950 82.050 607.050 ;
        RECT 52.950 601.800 55.050 603.900 ;
        RECT 55.950 601.800 58.050 603.900 ;
        RECT 58.950 601.800 61.050 603.900 ;
        RECT 61.950 601.800 64.050 603.900 ;
        RECT 70.950 601.800 73.050 603.900 ;
        RECT 73.950 601.800 76.050 603.900 ;
        RECT 76.950 601.800 79.050 603.900 ;
        RECT 79.950 601.800 82.050 603.900 ;
        RECT 49.950 598.950 52.050 601.050 ;
        RECT 53.400 600.000 54.600 601.500 ;
        RECT 59.400 600.750 60.600 601.500 ;
        RECT 41.400 584.400 45.450 585.450 ;
        RECT 10.950 565.800 13.050 567.900 ;
        RECT 22.950 567.450 25.050 568.050 ;
        RECT 20.400 566.400 25.050 567.450 ;
        RECT 1.950 559.950 4.050 562.050 ;
        RECT 1.950 538.950 4.050 541.050 ;
        RECT 2.400 490.050 3.450 538.950 ;
        RECT 11.400 528.450 12.450 565.800 ;
        RECT 20.400 532.050 21.450 566.400 ;
        RECT 22.950 565.950 25.050 566.400 ;
        RECT 28.950 565.950 31.050 568.050 ;
        RECT 37.950 565.950 40.050 568.050 ;
        RECT 31.950 550.950 34.050 553.050 ;
        RECT 13.950 528.450 16.050 532.050 ;
        RECT 19.950 529.950 22.050 532.050 ;
        RECT 11.400 528.000 16.050 528.450 ;
        RECT 20.400 528.600 21.450 529.950 ;
        RECT 11.400 527.400 15.600 528.000 ;
        RECT 14.400 526.200 15.600 527.400 ;
        RECT 20.400 526.200 21.600 528.600 ;
        RECT 28.950 528.000 31.050 532.050 ;
        RECT 32.400 529.050 33.450 550.950 ;
        RECT 41.400 550.050 42.450 584.400 ;
        RECT 50.400 580.050 51.450 598.950 ;
        RECT 52.950 595.950 55.050 600.000 ;
        RECT 58.950 595.950 61.050 600.750 ;
        RECT 64.950 598.950 67.050 601.050 ;
        RECT 74.400 600.000 75.600 601.500 ;
        RECT 55.950 583.950 58.050 586.050 ;
        RECT 49.950 577.950 52.050 580.050 ;
        RECT 49.950 572.100 52.050 574.200 ;
        RECT 56.400 573.600 57.450 583.950 ;
        RECT 61.950 577.950 64.050 580.050 ;
        RECT 50.400 571.350 51.600 572.100 ;
        RECT 56.400 571.350 57.600 573.600 ;
        RECT 46.950 568.950 49.050 571.050 ;
        RECT 49.950 568.950 52.050 571.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 55.950 568.950 58.050 571.050 ;
        RECT 47.400 566.400 48.600 568.650 ;
        RECT 53.400 567.900 54.600 568.650 ;
        RECT 47.400 562.050 48.450 566.400 ;
        RECT 52.950 565.800 55.050 567.900 ;
        RECT 55.950 562.950 58.050 565.050 ;
        RECT 46.950 559.950 49.050 562.050 ;
        RECT 40.950 547.950 43.050 550.050 ;
        RECT 29.400 526.200 30.600 528.000 ;
        RECT 31.950 526.950 34.050 529.050 ;
        RECT 34.950 528.000 37.050 532.050 ;
        RECT 35.400 526.200 36.600 528.000 ;
        RECT 43.950 526.950 46.050 529.050 ;
        RECT 49.950 526.950 52.050 529.050 ;
        RECT 56.400 528.600 57.450 562.950 ;
        RECT 62.400 559.050 63.450 577.950 ;
        RECT 65.400 574.050 66.450 598.950 ;
        RECT 73.950 595.950 76.050 600.000 ;
        RECT 80.400 599.400 81.600 601.500 ;
        RECT 67.950 583.950 70.050 586.050 ;
        RECT 64.950 571.950 67.050 574.050 ;
        RECT 68.400 573.600 69.450 583.950 ;
        RECT 80.400 574.350 81.450 599.400 ;
        RECT 82.950 598.950 85.050 601.050 ;
        RECT 83.400 589.050 84.450 598.950 ;
        RECT 82.950 586.950 85.050 589.050 ;
        RECT 86.400 580.050 87.450 607.800 ;
        RECT 92.400 606.600 93.450 607.950 ;
        RECT 95.400 607.050 96.450 610.950 ;
        RECT 92.400 604.200 93.600 606.600 ;
        RECT 94.950 604.950 97.050 607.050 ;
        RECT 97.950 606.000 100.050 610.050 ;
        RECT 101.400 607.050 102.450 649.800 ;
        RECT 104.400 622.050 105.450 649.950 ;
        RECT 113.400 649.500 114.600 650.250 ;
        RECT 131.400 649.500 132.600 650.250 ;
        RECT 109.950 647.100 112.050 649.200 ;
        RECT 112.950 647.100 115.050 649.200 ;
        RECT 118.950 647.100 121.050 649.200 ;
        RECT 127.950 647.100 130.050 649.200 ;
        RECT 130.950 647.100 133.050 649.200 ;
        RECT 133.950 647.100 136.050 649.200 ;
        RECT 106.950 643.950 109.050 646.050 ;
        RECT 110.400 645.000 111.600 646.800 ;
        RECT 103.950 619.950 106.050 622.050 ;
        RECT 107.400 619.050 108.450 643.950 ;
        RECT 109.950 640.950 112.050 645.000 ;
        RECT 119.400 644.400 120.600 646.800 ;
        RECT 128.400 646.050 129.600 646.800 ;
        RECT 127.950 645.450 130.050 646.050 ;
        RECT 127.950 644.400 132.450 645.450 ;
        RECT 119.400 631.050 120.450 644.400 ;
        RECT 127.950 643.950 130.050 644.400 ;
        RECT 118.950 628.950 121.050 631.050 ;
        RECT 127.950 619.950 130.050 622.050 ;
        RECT 106.950 616.950 109.050 619.050 ;
        RECT 121.950 616.950 124.050 619.050 ;
        RECT 109.950 610.950 112.050 613.050 ;
        RECT 98.400 604.200 99.600 606.000 ;
        RECT 100.950 604.950 103.050 607.050 ;
        RECT 106.950 604.950 109.050 607.050 ;
        RECT 91.950 601.800 94.050 603.900 ;
        RECT 94.950 601.800 97.050 603.900 ;
        RECT 97.950 601.800 100.050 603.900 ;
        RECT 100.950 601.800 103.050 603.900 ;
        RECT 95.400 600.000 96.600 601.500 ;
        RECT 94.950 595.950 97.050 600.000 ;
        RECT 101.400 599.400 102.600 601.500 ;
        RECT 101.400 595.050 102.450 599.400 ;
        RECT 107.400 598.050 108.450 604.950 ;
        RECT 110.400 604.050 111.450 610.950 ;
        RECT 112.950 606.600 117.000 607.050 ;
        RECT 122.400 606.600 123.450 616.950 ;
        RECT 128.400 607.050 129.450 619.950 ;
        RECT 131.400 616.050 132.450 644.400 ;
        RECT 134.400 644.400 135.600 646.800 ;
        RECT 134.400 631.050 135.450 644.400 ;
        RECT 140.400 643.050 141.450 658.950 ;
        RECT 143.400 652.050 144.450 662.400 ;
        RECT 142.950 649.950 145.050 652.050 ;
        RECT 146.400 651.600 147.450 670.950 ;
        RECT 149.400 661.050 150.450 676.950 ;
        RECT 154.950 670.950 157.050 673.050 ;
        RECT 148.950 658.950 151.050 661.050 ;
        RECT 146.400 649.350 147.600 651.600 ;
        RECT 145.950 646.950 148.050 649.050 ;
        RECT 148.950 646.950 151.050 649.050 ;
        RECT 142.950 643.950 145.050 646.050 ;
        RECT 149.400 645.000 150.600 646.650 ;
        RECT 139.950 640.950 142.050 643.050 ;
        RECT 133.950 628.950 136.050 631.050 ;
        RECT 136.950 616.950 139.050 619.050 ;
        RECT 130.950 613.950 133.050 616.050 ;
        RECT 112.950 604.950 117.600 606.600 ;
        RECT 116.400 604.350 117.600 604.950 ;
        RECT 122.400 604.350 123.600 606.600 ;
        RECT 127.950 604.950 130.050 607.050 ;
        RECT 137.400 606.600 138.450 616.950 ;
        RECT 143.400 610.200 144.450 643.950 ;
        RECT 148.950 640.950 151.050 645.000 ;
        RECT 155.400 619.050 156.450 670.950 ;
        RECT 164.400 664.050 165.450 677.400 ;
        RECT 169.950 676.650 172.050 678.750 ;
        RECT 185.400 677.400 186.600 679.500 ;
        RECT 191.400 678.750 192.600 679.500 ;
        RECT 166.950 672.450 169.050 676.050 ;
        RECT 166.950 672.000 171.450 672.450 ;
        RECT 167.400 671.400 171.450 672.000 ;
        RECT 163.950 661.950 166.050 664.050 ;
        RECT 163.950 650.250 166.050 652.350 ;
        RECT 170.400 652.050 171.450 671.400 ;
        RECT 185.400 670.050 186.450 677.400 ;
        RECT 190.950 676.650 193.050 678.750 ;
        RECT 193.950 670.950 196.050 673.050 ;
        RECT 184.950 667.950 187.050 670.050 ;
        RECT 175.950 661.950 178.050 664.050 ;
        RECT 164.400 649.500 165.600 650.250 ;
        RECT 169.950 649.950 172.050 652.050 ;
        RECT 160.950 647.100 163.050 649.200 ;
        RECT 163.950 647.100 166.050 649.200 ;
        RECT 166.950 647.100 169.050 649.200 ;
        RECT 161.400 644.400 162.600 646.800 ;
        RECT 161.400 625.050 162.450 644.400 ;
        RECT 163.950 643.950 166.050 646.050 ;
        RECT 164.400 637.050 165.450 643.950 ;
        RECT 163.950 634.950 166.050 637.050 ;
        RECT 176.400 634.050 177.450 661.950 ;
        RECT 190.950 655.950 193.050 658.050 ;
        RECT 184.950 650.100 187.050 652.200 ;
        RECT 185.400 649.350 186.600 650.100 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 184.950 646.950 187.050 649.050 ;
        RECT 178.950 643.950 181.050 646.050 ;
        RECT 182.400 644.400 183.600 646.650 ;
        RECT 175.950 631.950 178.050 634.050 ;
        RECT 160.950 622.950 163.050 625.050 ;
        RECT 169.950 619.950 172.050 622.050 ;
        RECT 154.950 616.950 157.050 619.050 ;
        RECT 170.400 616.050 171.450 619.950 ;
        RECT 172.950 616.950 175.050 619.050 ;
        RECT 169.950 613.950 172.050 616.050 ;
        RECT 163.950 610.950 166.050 613.050 ;
        RECT 142.950 608.100 145.050 610.200 ;
        RECT 148.950 607.950 151.050 610.050 ;
        RECT 151.950 607.950 154.050 610.050 ;
        RECT 137.400 604.350 138.600 606.600 ;
        RECT 142.950 604.950 145.050 607.050 ;
        RECT 143.400 604.350 144.600 604.950 ;
        RECT 109.950 601.950 112.050 604.050 ;
        RECT 115.950 601.950 118.050 604.050 ;
        RECT 118.950 601.950 121.050 604.050 ;
        RECT 121.950 601.950 124.050 604.050 ;
        RECT 124.950 601.950 127.050 604.050 ;
        RECT 133.950 601.950 136.050 604.050 ;
        RECT 136.950 601.950 139.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 142.950 601.950 145.050 604.050 ;
        RECT 109.950 598.800 112.050 600.900 ;
        RECT 119.400 599.400 120.600 601.650 ;
        RECT 125.400 600.900 126.600 601.650 ;
        RECT 134.400 600.900 135.600 601.650 ;
        RECT 106.950 595.950 109.050 598.050 ;
        RECT 100.950 592.950 103.050 595.050 ;
        RECT 110.400 589.050 111.450 598.800 ;
        RECT 115.950 595.950 118.050 598.050 ;
        RECT 119.400 597.450 120.450 599.400 ;
        RECT 124.950 598.800 127.050 600.900 ;
        RECT 133.950 598.800 136.050 600.900 ;
        RECT 140.400 599.400 141.600 601.650 ;
        RECT 119.400 596.400 126.450 597.450 ;
        RECT 109.950 586.950 112.050 589.050 ;
        RECT 85.950 577.950 88.050 580.050 ;
        RECT 97.950 577.950 100.050 580.050 ;
        RECT 68.400 571.500 69.600 573.600 ;
        RECT 73.950 572.250 76.050 574.350 ;
        RECT 79.950 572.250 82.050 574.350 ;
        RECT 88.950 572.250 91.050 574.350 ;
        RECT 94.950 572.250 97.050 574.350 ;
        RECT 98.400 574.050 99.450 577.950 ;
        RECT 116.400 577.050 117.450 595.950 ;
        RECT 121.950 583.950 124.050 586.050 ;
        RECT 115.950 574.950 118.050 577.050 ;
        RECT 74.400 571.500 75.600 572.250 ;
        RECT 89.400 571.500 90.600 572.250 ;
        RECT 95.400 571.500 96.600 572.250 ;
        RECT 97.950 571.950 100.050 574.050 ;
        RECT 100.950 572.100 103.050 574.200 ;
        RECT 106.950 572.100 109.050 574.200 ;
        RECT 112.950 572.100 115.050 574.200 ;
        RECT 67.950 569.100 70.050 571.200 ;
        RECT 70.950 569.100 73.050 571.200 ;
        RECT 73.950 569.100 76.050 571.200 ;
        RECT 76.950 569.100 79.050 571.200 ;
        RECT 85.950 569.100 88.050 571.200 ;
        RECT 88.950 569.100 91.050 571.200 ;
        RECT 91.950 569.100 94.050 571.200 ;
        RECT 94.950 569.100 97.050 571.200 ;
        RECT 67.950 565.950 70.050 568.050 ;
        RECT 71.400 567.000 72.600 568.800 ;
        RECT 61.950 556.950 64.050 559.050 ;
        RECT 64.950 547.950 67.050 550.050 ;
        RECT 10.950 523.800 13.050 525.900 ;
        RECT 13.950 523.800 16.050 525.900 ;
        RECT 16.950 523.800 19.050 525.900 ;
        RECT 19.950 523.800 22.050 525.900 ;
        RECT 28.950 523.800 31.050 525.900 ;
        RECT 31.950 523.800 34.050 525.900 ;
        RECT 34.950 523.800 37.050 525.900 ;
        RECT 37.950 523.800 40.050 525.900 ;
        RECT 11.400 521.400 12.600 523.500 ;
        RECT 17.400 522.750 18.600 523.500 ;
        RECT 32.400 522.750 33.600 523.500 ;
        RECT 38.400 522.750 39.600 523.500 ;
        RECT 44.400 523.050 45.450 526.950 ;
        RECT 50.400 526.200 51.600 526.950 ;
        RECT 56.400 526.200 57.600 528.600 ;
        RECT 49.950 523.800 52.050 525.900 ;
        RECT 52.950 523.800 55.050 525.900 ;
        RECT 55.950 523.800 58.050 525.900 ;
        RECT 58.950 523.800 61.050 525.900 ;
        RECT 11.400 499.050 12.450 521.400 ;
        RECT 16.950 520.650 19.050 522.750 ;
        RECT 31.950 520.650 34.050 522.750 ;
        RECT 37.950 520.650 40.050 522.750 ;
        RECT 43.950 520.950 46.050 523.050 ;
        RECT 53.400 522.000 54.600 523.500 ;
        RECT 38.400 502.050 39.450 520.650 ;
        RECT 43.950 517.800 46.050 519.900 ;
        RECT 52.950 517.950 55.050 522.000 ;
        RECT 59.400 521.400 60.600 523.500 ;
        RECT 65.400 523.050 66.450 547.950 ;
        RECT 13.950 499.950 16.050 502.050 ;
        RECT 37.950 499.950 40.050 502.050 ;
        RECT 4.950 496.950 7.050 499.050 ;
        RECT 10.950 496.950 13.050 499.050 ;
        RECT 1.950 487.950 4.050 490.050 ;
        RECT 5.400 442.050 6.450 496.950 ;
        RECT 14.400 495.600 15.450 499.950 ;
        RECT 14.400 493.350 15.600 495.600 ;
        RECT 28.950 495.000 31.050 499.050 ;
        RECT 29.400 493.350 30.600 495.000 ;
        RECT 34.950 494.100 37.050 499.050 ;
        RECT 44.400 495.600 45.450 517.800 ;
        RECT 59.400 502.050 60.450 521.400 ;
        RECT 64.950 520.950 67.050 523.050 ;
        RECT 68.400 508.050 69.450 565.950 ;
        RECT 70.950 562.950 73.050 567.000 ;
        RECT 77.400 566.400 78.600 568.800 ;
        RECT 86.400 566.400 87.600 568.800 ;
        RECT 92.400 566.400 93.600 568.800 ;
        RECT 77.400 559.050 78.450 566.400 ;
        RECT 86.400 565.050 87.450 566.400 ;
        RECT 85.950 562.950 88.050 565.050 ;
        RECT 76.950 556.950 79.050 559.050 ;
        RECT 86.400 547.050 87.450 562.950 ;
        RECT 92.400 559.050 93.450 566.400 ;
        RECT 97.950 565.950 100.050 568.050 ;
        RECT 91.950 556.950 94.050 559.050 ;
        RECT 98.400 553.050 99.450 565.950 ;
        RECT 101.400 562.050 102.450 572.100 ;
        RECT 107.400 571.350 108.600 572.100 ;
        RECT 113.400 571.350 114.600 572.100 ;
        RECT 106.950 568.950 109.050 571.050 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 112.950 568.950 115.050 571.050 ;
        RECT 115.950 568.950 118.050 571.050 ;
        RECT 103.950 562.950 106.050 568.050 ;
        RECT 110.400 567.900 111.600 568.650 ;
        RECT 109.950 565.800 112.050 567.900 ;
        RECT 116.400 566.400 117.600 568.650 ;
        RECT 122.400 567.900 123.450 583.950 ;
        RECT 125.400 574.050 126.450 596.400 ;
        RECT 140.400 592.050 141.450 599.400 ;
        RECT 142.950 595.950 145.050 598.050 ;
        RECT 133.950 589.950 136.050 592.050 ;
        RECT 139.950 589.950 142.050 592.050 ;
        RECT 134.400 585.450 135.450 589.950 ;
        RECT 139.950 585.450 142.050 586.050 ;
        RECT 134.400 584.400 142.050 585.450 ;
        RECT 139.950 583.950 142.050 584.400 ;
        RECT 136.950 580.950 139.050 583.050 ;
        RECT 124.950 571.950 127.050 574.050 ;
        RECT 130.950 573.000 133.050 577.050 ;
        RECT 137.400 573.600 138.450 580.950 ;
        RECT 143.400 577.050 144.450 595.950 ;
        RECT 145.950 592.950 148.050 595.050 ;
        RECT 146.400 583.050 147.450 592.950 ;
        RECT 149.400 592.050 150.450 607.950 ;
        RECT 148.950 589.950 151.050 592.050 ;
        RECT 152.400 583.050 153.450 607.950 ;
        RECT 160.950 606.000 163.050 610.050 ;
        RECT 164.400 607.050 165.450 610.950 ;
        RECT 161.400 604.200 162.600 606.000 ;
        RECT 163.950 604.950 166.050 607.050 ;
        RECT 166.950 606.000 169.050 610.050 ;
        RECT 167.400 604.200 168.600 606.000 ;
        RECT 157.950 601.800 160.050 603.900 ;
        RECT 160.950 601.800 163.050 603.900 ;
        RECT 163.950 601.800 166.050 603.900 ;
        RECT 166.950 601.800 169.050 603.900 ;
        RECT 158.400 599.400 159.600 601.500 ;
        RECT 164.400 599.400 165.600 601.500 ;
        RECT 158.400 589.050 159.450 599.400 ;
        RECT 157.950 586.950 160.050 589.050 ;
        RECT 164.400 586.050 165.450 599.400 ;
        RECT 166.950 586.950 169.050 589.050 ;
        RECT 163.950 583.950 166.050 586.050 ;
        RECT 145.950 580.950 148.050 583.050 ;
        RECT 152.400 581.400 157.050 583.050 ;
        RECT 153.000 580.950 157.050 581.400 ;
        RECT 163.950 580.800 166.050 582.900 ;
        RECT 142.950 574.950 145.050 577.050 ;
        RECT 151.800 576.000 153.900 576.900 ;
        RECT 131.400 571.500 132.600 573.000 ;
        RECT 137.400 571.500 138.600 573.600 ;
        RECT 127.950 569.100 130.050 571.200 ;
        RECT 130.950 569.100 133.050 571.200 ;
        RECT 133.950 569.100 136.050 571.200 ;
        RECT 136.950 569.100 139.050 571.200 ;
        RECT 143.400 571.050 144.450 574.950 ;
        RECT 151.800 574.800 154.050 576.000 ;
        RECT 154.950 574.950 160.050 577.050 ;
        RECT 151.950 573.000 154.050 574.800 ;
        RECT 159.000 573.600 163.050 574.050 ;
        RECT 152.400 571.500 153.600 573.000 ;
        RECT 158.400 571.950 163.050 573.600 ;
        RECT 158.400 571.500 159.600 571.950 ;
        RECT 142.950 568.950 145.050 571.050 ;
        RECT 148.950 569.100 151.050 571.200 ;
        RECT 151.950 569.100 154.050 571.200 ;
        RECT 154.950 569.100 157.050 571.200 ;
        RECT 157.950 569.100 160.050 571.200 ;
        RECT 100.950 561.450 103.050 562.050 ;
        RECT 100.950 561.000 105.450 561.450 ;
        RECT 100.950 560.400 106.050 561.000 ;
        RECT 100.950 559.950 103.050 560.400 ;
        RECT 103.950 556.950 106.050 560.400 ;
        RECT 116.400 553.050 117.450 566.400 ;
        RECT 121.950 565.800 124.050 567.900 ;
        RECT 124.950 565.950 127.050 568.050 ;
        RECT 128.400 567.000 129.600 568.800 ;
        RECT 134.400 568.050 135.600 568.800 ;
        RECT 149.400 568.050 150.600 568.800 ;
        RECT 155.400 568.050 156.600 568.800 ;
        RECT 121.950 556.950 124.050 559.050 ;
        RECT 97.950 550.950 100.050 553.050 ;
        RECT 115.950 550.950 118.050 553.050 ;
        RECT 118.950 547.950 121.050 550.050 ;
        RECT 85.950 544.950 88.050 547.050 ;
        RECT 115.950 544.950 118.050 547.050 ;
        RECT 116.400 535.050 117.450 544.950 ;
        RECT 119.400 541.050 120.450 547.950 ;
        RECT 122.400 544.050 123.450 556.950 ;
        RECT 125.400 553.050 126.450 565.950 ;
        RECT 127.950 562.950 130.050 567.000 ;
        RECT 133.950 565.950 136.050 568.050 ;
        RECT 142.950 562.950 145.050 567.900 ;
        RECT 148.950 565.950 151.050 568.050 ;
        RECT 154.950 565.950 157.050 568.050 ;
        RECT 160.950 565.950 163.050 568.050 ;
        RECT 124.950 550.950 127.050 553.050 ;
        RECT 161.400 547.050 162.450 565.950 ;
        RECT 164.400 562.050 165.450 580.800 ;
        RECT 163.950 559.950 166.050 562.050 ;
        RECT 164.400 547.050 165.450 559.950 ;
        RECT 139.950 544.950 142.050 547.050 ;
        RECT 160.800 544.950 162.900 547.050 ;
        RECT 163.950 544.950 166.050 547.050 ;
        RECT 121.950 541.950 124.050 544.050 ;
        RECT 118.950 538.950 121.050 541.050 ;
        RECT 124.950 538.950 127.050 541.050 ;
        RECT 76.950 532.950 79.050 535.050 ;
        RECT 109.950 532.950 112.050 535.050 ;
        RECT 115.950 532.950 118.050 535.050 ;
        RECT 77.400 528.600 78.450 532.950 ;
        RECT 77.400 526.200 78.600 528.600 ;
        RECT 82.950 526.950 85.050 529.050 ;
        RECT 88.950 526.950 91.050 529.050 ;
        RECT 97.950 526.950 100.050 529.050 ;
        RECT 103.950 526.950 106.050 529.050 ;
        RECT 83.400 526.200 84.600 526.950 ;
        RECT 73.950 523.800 76.050 525.900 ;
        RECT 76.950 523.800 79.050 525.900 ;
        RECT 79.950 523.800 82.050 525.900 ;
        RECT 82.950 523.800 85.050 525.900 ;
        RECT 74.400 522.750 75.600 523.500 ;
        RECT 73.950 520.650 76.050 522.750 ;
        RECT 80.400 522.000 81.600 523.500 ;
        RECT 89.400 522.450 90.450 526.950 ;
        RECT 98.400 526.200 99.600 526.950 ;
        RECT 104.400 526.200 105.600 526.950 ;
        RECT 94.950 523.800 97.050 525.900 ;
        RECT 97.950 523.800 100.050 525.900 ;
        RECT 100.950 523.800 103.050 525.900 ;
        RECT 103.950 523.800 106.050 525.900 ;
        RECT 79.950 517.950 82.050 522.000 ;
        RECT 86.400 521.400 90.450 522.450 ;
        RECT 95.400 521.400 96.600 523.500 ;
        RECT 101.400 522.750 102.600 523.500 ;
        RECT 86.400 514.050 87.450 521.400 ;
        RECT 88.950 514.950 91.050 520.050 ;
        RECT 91.950 517.950 94.050 520.050 ;
        RECT 85.950 511.950 88.050 514.050 ;
        RECT 70.950 508.950 73.050 511.050 ;
        RECT 82.950 508.950 85.050 511.050 ;
        RECT 67.950 505.950 70.050 508.050 ;
        RECT 58.950 499.950 61.050 502.050 ;
        RECT 71.400 498.450 72.450 508.950 ;
        RECT 79.950 502.950 82.050 505.050 ;
        RECT 76.950 499.950 79.050 502.050 ;
        RECT 68.400 497.400 72.450 498.450 ;
        RECT 68.400 496.350 69.450 497.400 ;
        RECT 10.950 490.950 13.050 493.050 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 25.950 490.950 28.050 493.050 ;
        RECT 28.950 490.950 31.050 493.050 ;
        RECT 11.400 488.400 12.600 490.650 ;
        RECT 26.400 489.900 27.600 490.650 ;
        RECT 11.400 457.050 12.450 488.400 ;
        RECT 25.950 487.800 28.050 489.900 ;
        RECT 10.950 454.950 13.050 457.050 ;
        RECT 16.950 454.950 19.050 457.050 ;
        RECT 26.400 456.450 27.450 487.800 ;
        RECT 35.400 475.050 36.450 494.100 ;
        RECT 44.400 493.350 45.600 495.600 ;
        RECT 49.950 494.100 52.050 496.200 ;
        RECT 61.950 494.250 64.050 496.350 ;
        RECT 67.950 494.250 70.050 496.350 ;
        RECT 50.400 493.350 51.600 494.100 ;
        RECT 62.400 493.500 63.600 494.250 ;
        RECT 68.400 493.500 69.600 494.250 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 43.950 490.950 46.050 493.050 ;
        RECT 46.950 490.950 49.050 493.050 ;
        RECT 49.950 490.950 52.050 493.050 ;
        RECT 61.950 491.100 64.050 493.200 ;
        RECT 64.950 491.100 67.050 493.200 ;
        RECT 67.950 491.100 70.050 493.200 ;
        RECT 70.950 491.100 73.050 493.200 ;
        RECT 41.400 488.400 42.600 490.650 ;
        RECT 47.400 489.900 48.600 490.650 ;
        RECT 41.400 484.050 42.450 488.400 ;
        RECT 46.950 487.800 49.050 489.900 ;
        RECT 65.400 488.400 66.600 490.800 ;
        RECT 71.400 488.400 72.600 490.800 ;
        RECT 40.950 481.950 43.050 484.050 ;
        RECT 46.950 481.950 49.050 484.050 ;
        RECT 34.950 472.950 37.050 475.050 ;
        RECT 40.950 472.950 43.050 475.050 ;
        RECT 23.400 455.400 27.450 456.450 ;
        RECT 10.950 449.100 13.050 451.200 ;
        RECT 17.400 450.600 18.450 454.950 ;
        RECT 23.400 451.050 24.450 455.400 ;
        RECT 25.950 451.950 28.050 454.050 ;
        RECT 11.400 448.350 12.600 449.100 ;
        RECT 17.400 448.350 18.600 450.600 ;
        RECT 22.950 448.950 25.050 451.050 ;
        RECT 10.950 445.950 13.050 448.050 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 16.950 445.950 19.050 448.050 ;
        RECT 19.950 445.950 22.050 448.050 ;
        RECT 7.950 442.950 10.050 445.050 ;
        RECT 14.400 443.400 15.600 445.650 ;
        RECT 20.400 444.000 21.600 445.650 ;
        RECT 4.950 439.950 7.050 442.050 ;
        RECT 4.950 418.950 7.050 421.050 ;
        RECT 5.400 412.050 6.450 418.950 ;
        RECT 8.400 417.450 9.450 442.950 ;
        RECT 14.400 424.050 15.450 443.400 ;
        RECT 19.950 439.950 22.050 444.000 ;
        RECT 22.950 442.950 25.050 445.050 ;
        RECT 26.400 444.450 27.450 451.950 ;
        RECT 34.950 450.000 37.050 454.050 ;
        RECT 41.400 450.600 42.450 472.950 ;
        RECT 35.400 448.200 36.600 450.000 ;
        RECT 41.400 448.200 42.600 450.600 ;
        RECT 31.950 445.800 34.050 447.900 ;
        RECT 34.950 445.800 37.050 447.900 ;
        RECT 37.950 445.800 40.050 447.900 ;
        RECT 40.950 445.800 43.050 447.900 ;
        RECT 26.400 443.400 30.450 444.450 ;
        RECT 13.950 421.950 16.050 424.050 ;
        RECT 10.950 420.900 15.000 421.050 ;
        RECT 10.950 418.950 16.050 420.900 ;
        RECT 13.950 418.800 16.050 418.950 ;
        RECT 11.400 417.450 12.600 417.600 ;
        RECT 8.400 416.400 12.600 417.450 ;
        RECT 11.400 415.500 12.600 416.400 ;
        RECT 16.950 416.250 19.050 418.350 ;
        RECT 23.400 418.050 24.450 442.950 ;
        RECT 29.400 436.050 30.450 443.400 ;
        RECT 32.400 443.400 33.600 445.500 ;
        RECT 38.400 443.400 39.600 445.500 ;
        RECT 28.950 433.950 31.050 436.050 ;
        RECT 32.400 424.050 33.450 443.400 ;
        RECT 38.400 439.050 39.450 443.400 ;
        RECT 37.950 436.950 40.050 439.050 ;
        RECT 25.950 421.950 28.050 424.050 ;
        RECT 31.950 421.950 34.050 424.050 ;
        RECT 40.950 421.950 43.050 424.050 ;
        RECT 17.400 415.500 18.600 416.250 ;
        RECT 22.950 415.950 25.050 418.050 ;
        RECT 10.950 413.100 13.050 415.200 ;
        RECT 13.950 413.100 16.050 415.200 ;
        RECT 16.950 413.100 19.050 415.200 ;
        RECT 19.950 413.100 22.050 415.200 ;
        RECT 14.400 412.050 15.600 412.800 ;
        RECT 20.400 412.050 21.600 412.800 ;
        RECT 4.950 409.950 7.050 412.050 ;
        RECT 13.800 409.950 15.900 412.050 ;
        RECT 16.800 411.000 18.900 412.050 ;
        RECT 16.800 409.950 19.050 411.000 ;
        RECT 19.950 409.950 22.050 412.050 ;
        RECT 16.950 406.950 19.050 409.950 ;
        RECT 26.400 385.050 27.450 421.950 ;
        RECT 28.950 415.950 31.050 421.050 ;
        RECT 34.950 417.000 37.050 421.050 ;
        RECT 35.400 415.350 36.600 417.000 ;
        RECT 31.950 412.950 34.050 415.050 ;
        RECT 34.950 412.950 37.050 415.050 ;
        RECT 32.400 411.900 33.600 412.650 ;
        RECT 31.950 409.800 34.050 411.900 ;
        RECT 28.950 408.450 31.050 409.050 ;
        RECT 37.950 408.450 40.050 412.050 ;
        RECT 28.950 408.000 40.050 408.450 ;
        RECT 28.950 407.400 39.450 408.000 ;
        RECT 28.950 406.950 31.050 407.400 ;
        RECT 28.950 391.950 31.050 394.050 ;
        RECT 4.950 382.950 7.050 385.050 ;
        RECT 25.950 382.950 28.050 385.050 ;
        RECT 5.400 355.050 6.450 382.950 ;
        RECT 13.950 370.950 16.050 376.050 ;
        RECT 29.400 373.050 30.450 391.950 ;
        RECT 41.400 379.050 42.450 421.950 ;
        RECT 47.400 421.050 48.450 481.950 ;
        RECT 65.400 466.050 66.450 488.400 ;
        RECT 71.400 484.050 72.450 488.400 ;
        RECT 70.950 481.950 73.050 484.050 ;
        RECT 61.950 463.950 64.050 466.050 ;
        RECT 64.950 463.950 67.050 466.050 ;
        RECT 55.950 450.000 58.050 453.900 ;
        RECT 62.400 450.600 63.450 463.950 ;
        RECT 64.950 457.950 67.050 460.050 ;
        RECT 65.400 451.050 66.450 457.950 ;
        RECT 71.400 454.050 72.450 481.950 ;
        RECT 77.400 478.050 78.450 499.950 ;
        RECT 80.400 496.050 81.450 502.950 ;
        RECT 83.400 502.050 84.450 508.950 ;
        RECT 82.950 499.950 85.050 502.050 ;
        RECT 79.950 493.950 82.050 496.050 ;
        RECT 85.950 494.100 88.050 496.200 ;
        RECT 92.400 495.600 93.450 517.950 ;
        RECT 95.400 496.050 96.450 521.400 ;
        RECT 100.950 520.650 103.050 522.750 ;
        RECT 97.950 517.950 100.050 520.050 ;
        RECT 98.400 502.050 99.450 517.950 ;
        RECT 101.400 517.050 102.450 520.650 ;
        RECT 100.950 514.950 103.050 517.050 ;
        RECT 110.400 511.050 111.450 532.950 ;
        RECT 125.400 532.050 126.450 538.950 ;
        RECT 130.950 532.950 133.050 535.050 ;
        RECT 118.950 526.950 121.050 532.050 ;
        RECT 124.950 529.950 127.050 532.050 ;
        RECT 131.400 529.050 132.450 532.950 ;
        RECT 119.400 526.200 120.600 526.950 ;
        RECT 124.950 526.800 127.050 528.900 ;
        RECT 130.950 526.950 133.050 529.050 ;
        RECT 136.950 528.000 139.050 532.050 ;
        RECT 140.400 529.050 141.450 544.950 ;
        RECT 163.950 541.800 166.050 543.900 ;
        RECT 157.950 538.950 160.050 541.050 ;
        RECT 151.950 532.950 154.050 535.050 ;
        RECT 142.950 529.950 145.050 532.050 ;
        RECT 125.400 526.200 126.600 526.800 ;
        RECT 137.400 526.350 138.600 528.000 ;
        RECT 139.950 526.950 142.050 529.050 ;
        RECT 115.950 523.800 118.050 525.900 ;
        RECT 118.950 523.800 121.050 525.900 ;
        RECT 121.950 523.800 124.050 525.900 ;
        RECT 124.950 523.800 127.050 525.900 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 116.400 521.400 117.600 523.500 ;
        RECT 122.400 522.750 123.600 523.500 ;
        RECT 116.400 520.050 117.450 521.400 ;
        RECT 121.950 520.650 124.050 522.750 ;
        RECT 127.950 520.950 130.050 523.050 ;
        RECT 134.400 522.000 135.600 523.650 ;
        RECT 112.950 518.400 117.450 520.050 ;
        RECT 122.400 519.450 123.450 520.650 ;
        RECT 122.400 518.400 126.450 519.450 ;
        RECT 112.950 517.950 117.000 518.400 ;
        RECT 118.950 514.950 121.050 517.050 ;
        RECT 109.950 508.950 112.050 511.050 ;
        RECT 115.950 508.950 118.050 511.050 ;
        RECT 103.950 505.950 106.050 508.050 ;
        RECT 97.950 499.950 100.050 502.050 ;
        RECT 86.400 493.350 87.600 494.100 ;
        RECT 92.400 493.350 93.600 495.600 ;
        RECT 94.950 493.950 97.050 496.050 ;
        RECT 97.950 493.950 100.050 496.050 ;
        RECT 104.400 495.600 105.450 505.950 ;
        RECT 109.950 499.950 112.050 502.050 ;
        RECT 110.400 495.600 111.450 499.950 ;
        RECT 82.950 490.950 85.050 493.050 ;
        RECT 85.950 490.950 88.050 493.050 ;
        RECT 88.950 490.950 91.050 493.050 ;
        RECT 91.950 490.950 94.050 493.050 ;
        RECT 79.800 487.950 81.900 490.050 ;
        RECT 83.400 489.900 84.600 490.650 ;
        RECT 89.400 489.900 90.600 490.650 ;
        RECT 76.950 475.950 79.050 478.050 ;
        RECT 77.400 454.050 78.450 475.950 ;
        RECT 80.400 460.050 81.450 487.950 ;
        RECT 82.950 487.800 85.050 489.900 ;
        RECT 88.950 487.800 91.050 489.900 ;
        RECT 94.950 487.950 97.050 490.050 ;
        RECT 95.400 460.050 96.450 487.950 ;
        RECT 98.400 484.050 99.450 493.950 ;
        RECT 104.400 493.350 105.600 495.600 ;
        RECT 110.400 493.350 111.600 495.600 ;
        RECT 103.950 490.950 106.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 107.400 489.900 108.600 490.650 ;
        RECT 116.400 490.050 117.450 508.950 ;
        RECT 119.400 496.050 120.450 514.950 ;
        RECT 125.400 513.450 126.450 518.400 ;
        RECT 128.400 517.050 129.450 520.950 ;
        RECT 133.950 517.950 136.050 522.000 ;
        RECT 127.950 514.950 130.050 517.050 ;
        RECT 143.400 514.050 144.450 529.950 ;
        RECT 152.400 528.600 153.450 532.950 ;
        RECT 158.400 528.600 159.450 538.950 ;
        RECT 164.400 538.050 165.450 541.800 ;
        RECT 163.950 535.950 166.050 538.050 ;
        RECT 167.400 534.450 168.450 586.950 ;
        RECT 173.400 577.050 174.450 616.950 ;
        RECT 179.400 606.600 180.450 643.950 ;
        RECT 182.400 637.050 183.450 644.400 ;
        RECT 187.950 643.950 190.050 646.050 ;
        RECT 181.950 634.950 184.050 637.050 ;
        RECT 188.400 631.050 189.450 643.950 ;
        RECT 187.950 628.950 190.050 631.050 ;
        RECT 191.400 628.050 192.450 655.950 ;
        RECT 194.400 652.050 195.450 670.950 ;
        RECT 197.400 658.050 198.450 691.950 ;
        RECT 206.400 684.600 207.450 728.400 ;
        RECT 209.400 724.050 210.450 755.400 ;
        RECT 215.400 742.050 216.450 755.400 ;
        RECT 214.950 739.950 217.050 742.050 ;
        RECT 230.400 736.050 231.450 755.400 ;
        RECT 236.400 742.050 237.450 755.400 ;
        RECT 238.950 754.950 241.050 757.050 ;
        RECT 248.400 755.400 249.600 757.500 ;
        RECT 254.400 756.750 255.600 757.500 ;
        RECT 239.400 751.050 240.450 754.950 ;
        RECT 238.950 748.950 241.050 751.050 ;
        RECT 235.950 739.950 238.050 742.050 ;
        RECT 248.400 739.050 249.450 755.400 ;
        RECT 253.950 754.650 256.050 756.750 ;
        RECT 269.400 755.400 270.600 757.500 ;
        RECT 275.400 755.400 276.600 757.500 ;
        RECT 269.400 751.050 270.450 755.400 ;
        RECT 268.950 748.950 271.050 751.050 ;
        RECT 235.950 736.800 238.050 738.900 ;
        RECT 247.950 736.950 250.050 739.050 ;
        RECT 229.950 733.950 232.050 736.050 ;
        RECT 236.400 733.050 237.450 736.800 ;
        RECT 275.400 736.050 276.450 755.400 ;
        RECT 277.950 751.950 280.050 757.050 ;
        RECT 281.400 751.050 282.450 796.800 ;
        RECT 287.400 796.050 288.450 802.950 ;
        RECT 293.400 800.400 294.600 802.800 ;
        RECT 299.400 801.000 300.600 802.800 ;
        RECT 286.950 793.950 289.050 796.050 ;
        RECT 293.400 787.050 294.450 800.400 ;
        RECT 298.950 796.950 301.050 801.000 ;
        RECT 305.400 800.400 306.600 802.800 ;
        RECT 314.400 801.900 315.450 805.950 ;
        RECT 323.400 805.350 324.600 806.100 ;
        RECT 335.400 805.500 336.600 806.250 ;
        RECT 319.950 802.950 322.050 805.050 ;
        RECT 322.950 802.950 325.050 805.050 ;
        RECT 331.950 803.100 334.050 805.200 ;
        RECT 334.950 803.100 337.050 805.200 ;
        RECT 337.950 803.100 340.050 805.200 ;
        RECT 320.400 801.900 321.600 802.650 ;
        RECT 305.400 793.050 306.450 800.400 ;
        RECT 313.950 799.800 316.050 801.900 ;
        RECT 319.950 799.800 322.050 801.900 ;
        RECT 332.400 800.400 333.600 802.800 ;
        RECT 304.950 790.950 307.050 793.050 ;
        RECT 292.950 784.950 295.050 787.050 ;
        RECT 286.950 762.000 289.050 766.050 ;
        RECT 292.950 762.000 295.050 766.050 ;
        RECT 287.400 760.200 288.600 762.000 ;
        RECT 293.400 760.200 294.600 762.000 ;
        RECT 286.950 757.800 289.050 759.900 ;
        RECT 289.950 757.800 292.050 759.900 ;
        RECT 292.950 757.800 295.050 759.900 ;
        RECT 295.950 757.800 298.050 759.900 ;
        RECT 290.400 756.750 291.600 757.500 ;
        RECT 289.950 754.650 292.050 756.750 ;
        RECT 296.400 755.400 297.600 757.500 ;
        RECT 280.950 748.950 283.050 751.050 ;
        RECT 296.400 739.050 297.450 755.400 ;
        RECT 305.400 745.050 306.450 790.950 ;
        RECT 332.400 778.050 333.450 800.400 ;
        RECT 344.400 784.050 345.450 806.250 ;
        RECT 352.950 802.950 355.050 805.050 ;
        RECT 358.950 802.950 361.050 805.050 ;
        RECT 353.400 801.900 354.600 802.650 ;
        RECT 365.400 802.050 366.450 806.250 ;
        RECT 374.400 805.500 375.600 806.250 ;
        RECT 388.950 806.100 391.050 808.200 ;
        RECT 395.400 807.600 396.450 814.950 ;
        RECT 403.950 811.950 406.050 814.050 ;
        RECT 451.950 811.950 454.050 814.050 ;
        RECT 389.400 805.350 390.600 806.100 ;
        RECT 395.400 805.350 396.600 807.600 ;
        RECT 370.950 803.100 373.050 805.200 ;
        RECT 373.950 803.100 376.050 805.200 ;
        RECT 379.950 803.100 382.050 805.200 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 391.950 802.950 394.050 805.050 ;
        RECT 394.950 802.950 397.050 805.050 ;
        RECT 397.950 802.950 400.050 805.050 ;
        RECT 352.950 799.800 355.050 801.900 ;
        RECT 364.950 799.950 367.050 802.050 ;
        RECT 371.400 800.400 372.600 802.800 ;
        RECT 380.400 800.400 381.600 802.800 ;
        RECT 349.950 796.950 352.050 799.050 ;
        RECT 350.400 793.050 351.450 796.950 ;
        RECT 349.950 790.950 352.050 793.050 ;
        RECT 353.400 787.050 354.450 799.800 ;
        RECT 371.400 796.050 372.450 800.400 ;
        RECT 370.950 793.950 373.050 796.050 ;
        RECT 367.950 789.450 370.050 793.050 ;
        RECT 373.950 789.450 376.050 790.050 ;
        RECT 367.950 789.000 376.050 789.450 ;
        RECT 368.400 788.400 376.050 789.000 ;
        RECT 373.950 787.950 376.050 788.400 ;
        RECT 352.950 784.950 355.050 787.050 ;
        RECT 370.950 784.950 373.050 787.050 ;
        RECT 343.950 781.950 346.050 784.050 ;
        RECT 319.950 775.950 322.050 778.050 ;
        RECT 331.950 775.950 334.050 778.050 ;
        RECT 320.400 766.050 321.450 775.950 ;
        RECT 332.400 772.050 333.450 775.950 ;
        RECT 331.950 769.950 334.050 772.050 ;
        RECT 344.400 769.050 345.450 781.950 ;
        RECT 367.950 775.950 370.050 778.050 ;
        RECT 361.950 769.950 364.050 772.050 ;
        RECT 334.950 766.950 337.050 769.050 ;
        RECT 343.950 766.950 346.050 769.050 ;
        RECT 313.950 762.000 316.050 766.050 ;
        RECT 319.950 763.950 322.050 766.050 ;
        RECT 325.950 763.950 328.050 766.050 ;
        RECT 314.400 760.200 315.600 762.000 ;
        RECT 319.950 760.800 322.050 762.900 ;
        RECT 320.400 760.200 321.600 760.800 ;
        RECT 310.950 757.800 313.050 759.900 ;
        RECT 313.950 757.800 316.050 759.900 ;
        RECT 316.950 757.800 319.050 759.900 ;
        RECT 319.950 757.800 322.050 759.900 ;
        RECT 311.400 757.050 312.600 757.500 ;
        RECT 307.950 755.400 312.600 757.050 ;
        RECT 317.400 756.000 318.600 757.500 ;
        RECT 326.400 757.050 327.450 763.950 ;
        RECT 335.400 763.050 336.450 766.950 ;
        RECT 334.950 760.950 337.050 763.050 ;
        RECT 340.950 760.950 343.050 763.050 ;
        RECT 346.950 760.950 349.050 763.050 ;
        RECT 355.950 762.000 358.050 766.050 ;
        RECT 358.950 763.950 361.050 769.050 ;
        RECT 362.400 762.600 363.450 769.950 ;
        RECT 335.400 760.200 336.600 760.950 ;
        RECT 341.400 760.200 342.600 760.950 ;
        RECT 331.950 757.800 334.050 759.900 ;
        RECT 334.950 757.800 337.050 759.900 ;
        RECT 337.950 757.800 340.050 759.900 ;
        RECT 340.950 757.800 343.050 759.900 ;
        RECT 307.950 754.950 312.000 755.400 ;
        RECT 316.950 751.950 319.050 756.000 ;
        RECT 325.950 754.950 328.050 757.050 ;
        RECT 332.400 755.400 333.600 757.500 ;
        RECT 338.400 756.750 339.600 757.500 ;
        RECT 347.400 756.750 348.450 760.950 ;
        RECT 356.400 760.200 357.600 762.000 ;
        RECT 362.400 760.200 363.600 762.600 ;
        RECT 352.950 757.800 355.050 759.900 ;
        RECT 355.950 757.800 358.050 759.900 ;
        RECT 358.950 757.800 361.050 759.900 ;
        RECT 361.950 757.800 364.050 759.900 ;
        RECT 353.400 756.750 354.600 757.500 ;
        RECT 304.950 742.950 307.050 745.050 ;
        RECT 328.950 742.950 331.050 745.050 ;
        RECT 289.950 736.950 292.050 739.050 ;
        RECT 295.950 736.950 298.050 739.050 ;
        RECT 250.950 733.950 253.050 736.050 ;
        RECT 262.950 733.950 265.050 736.050 ;
        RECT 274.950 733.950 277.050 736.050 ;
        RECT 283.950 733.950 286.050 736.050 ;
        RECT 214.950 728.250 217.050 730.350 ;
        RECT 220.950 728.250 223.050 730.350 ;
        RECT 226.950 728.250 229.050 733.050 ;
        RECT 235.950 730.950 238.050 733.050 ;
        RECT 236.400 729.600 237.450 730.950 ;
        RECT 215.400 727.500 216.600 728.250 ;
        RECT 221.400 727.500 222.600 728.250 ;
        RECT 236.400 727.500 237.600 729.600 ;
        RECT 241.950 728.250 244.050 730.350 ;
        RECT 242.400 727.500 243.600 728.250 ;
        RECT 214.950 725.100 217.050 727.200 ;
        RECT 217.950 725.100 220.050 727.200 ;
        RECT 220.950 725.100 223.050 727.200 ;
        RECT 223.950 725.100 226.050 727.200 ;
        RECT 232.950 725.100 235.050 727.200 ;
        RECT 235.950 725.100 238.050 727.200 ;
        RECT 238.950 725.100 241.050 727.200 ;
        RECT 241.950 725.100 244.050 727.200 ;
        RECT 247.950 724.950 250.050 730.050 ;
        RECT 218.400 724.050 219.600 724.800 ;
        RECT 208.950 721.950 211.050 724.050 ;
        RECT 217.950 718.950 220.050 724.050 ;
        RECT 224.400 722.400 225.600 724.800 ;
        RECT 233.400 723.000 234.600 724.800 ;
        RECT 224.400 715.050 225.450 722.400 ;
        RECT 232.950 718.950 235.050 723.000 ;
        RECT 239.400 722.400 240.600 724.800 ;
        RECT 239.400 715.050 240.450 722.400 ;
        RECT 251.400 721.050 252.450 733.950 ;
        RECT 256.950 728.250 259.050 730.350 ;
        RECT 263.400 729.600 264.450 733.950 ;
        RECT 275.400 730.050 276.450 733.950 ;
        RECT 257.400 727.500 258.600 728.250 ;
        RECT 263.400 727.500 264.600 729.600 ;
        RECT 274.800 727.950 276.900 730.050 ;
        RECT 277.950 728.250 280.050 730.350 ;
        RECT 284.400 729.600 285.450 733.950 ;
        RECT 290.400 730.050 291.450 736.950 ;
        RECT 329.400 736.050 330.450 742.950 ;
        RECT 332.400 742.050 333.450 755.400 ;
        RECT 337.950 754.650 340.050 756.750 ;
        RECT 346.950 754.650 349.050 756.750 ;
        RECT 352.950 754.650 355.050 756.750 ;
        RECT 359.400 755.400 360.600 757.500 ;
        RECT 338.400 748.050 339.450 754.650 ;
        RECT 359.400 751.050 360.450 755.400 ;
        RECT 364.950 754.650 367.050 756.750 ;
        RECT 358.950 748.950 361.050 751.050 ;
        RECT 365.400 748.050 366.450 754.650 ;
        RECT 337.950 745.950 340.050 748.050 ;
        RECT 364.950 745.950 367.050 748.050 ;
        RECT 368.400 742.050 369.450 775.950 ;
        RECT 371.400 762.450 372.450 784.950 ;
        RECT 380.400 772.050 381.450 800.400 ;
        RECT 385.950 799.950 388.050 802.050 ;
        RECT 392.400 800.400 393.600 802.650 ;
        RECT 398.400 801.900 399.600 802.650 ;
        RECT 404.400 801.900 405.450 811.950 ;
        RECT 412.950 806.250 415.050 808.350 ;
        RECT 418.950 807.000 421.050 811.050 ;
        RECT 430.950 808.950 433.050 811.050 ;
        RECT 413.400 805.500 414.600 806.250 ;
        RECT 419.400 805.500 420.600 807.000 ;
        RECT 409.950 803.100 412.050 805.200 ;
        RECT 412.950 803.100 415.050 805.200 ;
        RECT 415.950 803.100 418.050 805.200 ;
        RECT 418.950 803.100 421.050 805.200 ;
        RECT 421.950 803.100 424.050 805.200 ;
        RECT 386.400 784.050 387.450 799.950 ;
        RECT 392.400 784.050 393.450 800.400 ;
        RECT 397.950 799.800 400.050 801.900 ;
        RECT 403.950 799.800 406.050 801.900 ;
        RECT 410.400 800.400 411.600 802.800 ;
        RECT 410.400 793.050 411.450 800.400 ;
        RECT 412.950 799.950 415.050 802.050 ;
        RECT 416.400 800.400 417.600 802.800 ;
        RECT 400.950 790.950 403.050 793.050 ;
        RECT 409.950 790.950 412.050 793.050 ;
        RECT 385.950 781.950 388.050 784.050 ;
        RECT 391.950 781.950 394.050 784.050 ;
        RECT 379.950 769.950 382.050 772.050 ;
        RECT 373.950 765.450 376.050 769.050 ;
        RECT 373.950 765.000 378.450 765.450 ;
        RECT 374.400 764.400 378.450 765.000 ;
        RECT 373.950 762.450 376.050 763.050 ;
        RECT 371.400 761.400 376.050 762.450 ;
        RECT 377.400 762.450 378.450 764.400 ;
        RECT 379.950 762.450 382.050 763.050 ;
        RECT 377.400 761.400 382.050 762.450 ;
        RECT 373.950 760.950 376.050 761.400 ;
        RECT 379.950 760.950 382.050 761.400 ;
        RECT 385.950 760.950 391.050 763.050 ;
        RECT 394.950 762.000 397.050 766.050 ;
        RECT 401.400 763.050 402.450 790.950 ;
        RECT 409.950 787.800 412.050 789.900 ;
        RECT 410.400 774.450 411.450 787.800 ;
        RECT 413.400 787.050 414.450 799.950 ;
        RECT 412.950 784.950 415.050 787.050 ;
        RECT 416.400 784.050 417.450 800.400 ;
        RECT 418.950 799.950 421.050 802.050 ;
        RECT 422.400 800.400 423.600 802.800 ;
        RECT 431.400 802.050 432.450 808.950 ;
        RECT 452.400 808.200 453.450 811.950 ;
        RECT 451.950 806.100 454.050 808.200 ;
        RECT 452.400 805.350 453.600 806.100 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 442.950 802.950 445.050 805.050 ;
        RECT 451.950 802.950 454.050 805.050 ;
        RECT 454.950 802.950 457.050 805.050 ;
        RECT 415.950 781.950 418.050 784.050 ;
        RECT 410.400 773.400 414.450 774.450 ;
        RECT 413.400 772.050 414.450 773.400 ;
        RECT 409.950 769.950 412.050 772.050 ;
        RECT 413.400 770.400 418.050 772.050 ;
        RECT 414.000 769.950 418.050 770.400 ;
        RECT 403.950 763.950 409.050 766.050 ;
        RECT 374.400 760.200 375.600 760.950 ;
        RECT 380.400 760.200 381.600 760.950 ;
        RECT 373.950 757.800 376.050 759.900 ;
        RECT 376.950 757.800 379.050 759.900 ;
        RECT 379.950 757.800 382.050 759.900 ;
        RECT 370.950 754.950 373.050 757.050 ;
        RECT 377.400 755.400 378.600 757.500 ;
        RECT 331.950 739.950 334.050 742.050 ;
        RECT 346.950 739.950 349.050 742.050 ;
        RECT 367.950 739.950 370.050 742.050 ;
        RECT 316.950 733.950 319.050 736.050 ;
        RECT 328.950 733.950 331.050 736.050 ;
        RECT 278.400 727.500 279.600 728.250 ;
        RECT 284.400 727.500 285.600 729.600 ;
        RECT 289.800 727.950 291.900 730.050 ;
        RECT 295.950 728.100 298.050 730.200 ;
        RECT 301.950 729.000 304.050 733.050 ;
        RECT 310.950 730.950 313.050 733.050 ;
        RECT 296.400 727.350 297.600 728.100 ;
        RECT 302.400 727.350 303.600 729.000 ;
        RECT 256.950 725.100 259.050 727.200 ;
        RECT 259.950 725.100 262.050 727.200 ;
        RECT 262.950 725.100 265.050 727.200 ;
        RECT 265.950 725.100 268.050 727.200 ;
        RECT 277.950 725.100 280.050 727.200 ;
        RECT 280.950 725.100 283.050 727.200 ;
        RECT 283.950 725.100 286.050 727.200 ;
        RECT 286.950 725.100 289.050 727.200 ;
        RECT 295.950 724.950 298.050 727.050 ;
        RECT 298.950 724.950 301.050 727.050 ;
        RECT 301.950 724.950 304.050 727.050 ;
        RECT 304.950 724.950 307.050 727.050 ;
        RECT 253.950 721.950 256.050 724.050 ;
        RECT 256.950 721.950 259.050 724.050 ;
        RECT 260.400 722.400 261.600 724.800 ;
        RECT 266.400 724.050 267.600 724.800 ;
        RECT 250.950 718.950 253.050 721.050 ;
        RECT 241.950 715.950 244.050 718.050 ;
        RECT 223.950 712.950 226.050 715.050 ;
        RECT 238.950 712.950 241.050 715.050 ;
        RECT 235.950 709.950 238.050 712.050 ;
        RECT 236.400 700.050 237.450 709.950 ;
        RECT 217.950 697.950 220.050 700.050 ;
        RECT 226.950 697.950 229.050 700.050 ;
        RECT 235.950 697.950 238.050 700.050 ;
        RECT 206.400 682.350 207.600 684.600 ;
        RECT 211.950 683.100 214.050 685.200 ;
        RECT 212.400 682.350 213.600 683.100 ;
        RECT 202.950 679.950 205.050 682.050 ;
        RECT 205.950 679.950 208.050 682.050 ;
        RECT 208.950 679.950 211.050 682.050 ;
        RECT 211.950 679.950 214.050 682.050 ;
        RECT 203.400 677.400 204.600 679.650 ;
        RECT 209.400 677.400 210.600 679.650 ;
        RECT 203.400 675.450 204.450 677.400 ;
        RECT 203.400 674.400 207.450 675.450 ;
        RECT 202.950 661.950 205.050 664.050 ;
        RECT 196.950 655.950 199.050 658.050 ;
        RECT 193.950 649.950 196.050 652.050 ;
        RECT 196.950 650.250 199.050 652.350 ;
        RECT 203.400 651.600 204.450 661.950 ;
        RECT 206.400 655.050 207.450 674.400 ;
        RECT 209.400 661.050 210.450 677.400 ;
        RECT 214.950 676.950 217.050 679.050 ;
        RECT 211.950 673.950 214.050 676.050 ;
        RECT 208.950 658.950 211.050 661.050 ;
        RECT 205.950 652.950 208.050 655.050 ;
        RECT 212.400 652.200 213.450 673.950 ;
        RECT 215.400 664.050 216.450 676.950 ;
        RECT 218.400 670.050 219.450 697.950 ;
        RECT 227.400 684.600 228.450 697.950 ;
        RECT 227.400 682.350 228.600 684.600 ;
        RECT 232.950 683.100 235.050 685.200 ;
        RECT 233.400 682.350 234.600 683.100 ;
        RECT 226.950 679.950 229.050 682.050 ;
        RECT 229.950 679.950 232.050 682.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 235.950 679.950 238.050 682.050 ;
        RECT 230.400 678.900 231.600 679.650 ;
        RECT 229.950 676.800 232.050 678.900 ;
        RECT 236.400 678.000 237.600 679.650 ;
        RECT 235.950 673.950 238.050 678.000 ;
        RECT 220.950 670.950 223.050 673.050 ;
        RECT 217.950 667.950 220.050 670.050 ;
        RECT 214.950 661.950 217.050 664.050 ;
        RECT 215.400 654.450 216.450 661.950 ;
        RECT 221.400 658.050 222.450 670.950 ;
        RECT 238.950 667.950 241.050 670.050 ;
        RECT 223.950 664.950 226.050 667.050 ;
        RECT 220.950 655.950 223.050 658.050 ;
        RECT 215.400 653.400 219.450 654.450 ;
        RECT 197.400 649.500 198.600 650.250 ;
        RECT 203.400 649.500 204.600 651.600 ;
        RECT 211.950 650.100 214.050 652.200 ;
        RECT 218.400 651.600 219.450 653.400 ;
        RECT 224.400 651.600 225.450 664.950 ;
        RECT 229.950 661.950 232.050 664.050 ;
        RECT 218.400 649.500 219.600 651.600 ;
        RECT 224.400 649.500 225.600 651.600 ;
        RECT 196.950 647.100 199.050 649.200 ;
        RECT 199.950 647.100 202.050 649.200 ;
        RECT 202.950 647.100 205.050 649.200 ;
        RECT 205.950 647.100 208.050 649.200 ;
        RECT 214.950 647.100 217.050 649.200 ;
        RECT 217.950 647.100 220.050 649.200 ;
        RECT 220.950 647.100 223.050 649.200 ;
        RECT 223.950 647.100 226.050 649.200 ;
        RECT 193.950 643.950 196.050 646.050 ;
        RECT 200.400 644.400 201.600 646.800 ;
        RECT 206.400 646.050 207.600 646.800 ;
        RECT 190.950 625.950 193.050 628.050 ;
        RECT 194.400 619.050 195.450 643.950 ;
        RECT 200.400 643.050 201.450 644.400 ;
        RECT 205.950 643.950 208.050 646.050 ;
        RECT 215.400 645.000 216.600 646.800 ;
        RECT 199.950 640.950 202.050 643.050 ;
        RECT 200.400 634.050 201.450 640.950 ;
        RECT 202.950 637.950 205.050 643.050 ;
        RECT 206.400 637.050 207.450 643.950 ;
        RECT 214.950 640.950 217.050 645.000 ;
        RECT 221.400 644.400 222.600 646.800 ;
        RECT 208.950 637.950 214.050 640.050 ;
        RECT 221.400 637.050 222.450 644.400 ;
        RECT 205.950 634.950 208.050 637.050 ;
        RECT 220.950 634.950 223.050 637.050 ;
        RECT 199.950 631.950 202.050 634.050 ;
        RECT 208.950 631.950 211.050 634.050 ;
        RECT 199.950 628.800 202.050 630.900 ;
        RECT 193.950 616.950 196.050 619.050 ;
        RECT 187.950 613.950 190.050 616.050 ;
        RECT 179.400 604.200 180.600 606.600 ;
        RECT 185.400 606.450 186.600 606.600 ;
        RECT 188.400 606.450 189.450 613.950 ;
        RECT 185.400 605.400 189.450 606.450 ;
        RECT 196.950 606.000 199.050 610.050 ;
        RECT 200.400 607.050 201.450 628.800 ;
        RECT 202.950 625.950 205.050 628.050 ;
        RECT 185.400 604.200 186.600 605.400 ;
        RECT 197.400 604.350 198.600 606.000 ;
        RECT 199.950 604.950 202.050 607.050 ;
        RECT 178.950 601.800 181.050 603.900 ;
        RECT 181.950 601.800 184.050 603.900 ;
        RECT 184.950 601.800 187.050 603.900 ;
        RECT 193.950 601.950 196.050 604.050 ;
        RECT 196.950 601.950 199.050 604.050 ;
        RECT 182.400 600.750 183.600 601.500 ;
        RECT 181.950 598.650 184.050 600.750 ;
        RECT 190.950 598.950 193.050 601.050 ;
        RECT 194.400 599.400 195.600 601.650 ;
        RECT 178.950 592.950 181.050 595.050 ;
        RECT 179.400 589.050 180.450 592.950 ;
        RECT 178.950 586.950 181.050 589.050 ;
        RECT 172.950 574.950 175.050 577.050 ;
        RECT 169.950 573.600 174.000 574.050 ;
        RECT 179.400 573.600 180.450 586.950 ;
        RECT 191.400 585.450 192.450 598.950 ;
        RECT 194.400 597.450 195.450 599.400 ;
        RECT 194.400 596.400 198.450 597.450 ;
        RECT 191.400 584.400 195.450 585.450 ;
        RECT 190.950 580.950 193.050 583.050 ;
        RECT 184.950 577.950 187.050 580.050 ;
        RECT 185.400 574.050 186.450 577.950 ;
        RECT 169.950 571.950 174.600 573.600 ;
        RECT 173.400 571.500 174.600 571.950 ;
        RECT 179.400 571.500 180.600 573.600 ;
        RECT 184.950 571.950 187.050 574.050 ;
        RECT 191.400 573.450 192.450 580.950 ;
        RECT 194.400 577.050 195.450 584.400 ;
        RECT 197.400 577.050 198.450 596.400 ;
        RECT 193.800 574.950 195.900 577.050 ;
        RECT 188.400 572.400 192.450 573.450 ;
        RECT 196.950 573.000 199.050 577.050 ;
        RECT 203.400 574.050 204.450 625.950 ;
        RECT 209.400 622.050 210.450 631.950 ;
        RECT 230.400 628.050 231.450 661.950 ;
        RECT 239.400 661.050 240.450 667.950 ;
        RECT 242.400 664.050 243.450 715.950 ;
        RECT 250.950 706.950 253.050 709.050 ;
        RECT 251.400 694.050 252.450 706.950 ;
        RECT 250.950 691.950 253.050 694.050 ;
        RECT 247.950 688.950 250.050 691.050 ;
        RECT 248.400 684.600 249.450 688.950 ;
        RECT 254.400 685.200 255.450 721.950 ;
        RECT 257.400 706.050 258.450 721.950 ;
        RECT 260.400 709.050 261.450 722.400 ;
        RECT 265.800 721.950 267.900 724.050 ;
        RECT 268.950 721.950 271.050 724.050 ;
        RECT 281.400 722.400 282.600 724.800 ;
        RECT 287.400 723.000 288.600 724.800 ;
        RECT 289.800 723.000 291.900 724.050 ;
        RECT 259.950 706.950 262.050 709.050 ;
        RECT 256.950 703.950 259.050 706.050 ;
        RECT 256.950 697.950 259.050 700.050 ;
        RECT 257.400 691.050 258.450 697.950 ;
        RECT 256.950 688.950 259.050 691.050 ;
        RECT 269.400 688.050 270.450 721.950 ;
        RECT 281.400 709.050 282.450 722.400 ;
        RECT 286.950 718.950 289.050 723.000 ;
        RECT 289.800 721.950 292.050 723.000 ;
        RECT 292.950 721.950 295.050 724.050 ;
        RECT 299.400 722.400 300.600 724.650 ;
        RECT 305.400 723.900 306.600 724.650 ;
        RECT 289.950 718.950 292.050 721.950 ;
        RECT 283.950 715.950 286.050 718.050 ;
        RECT 280.950 706.950 283.050 709.050 ;
        RECT 284.400 706.050 285.450 715.950 ;
        RECT 293.400 715.050 294.450 721.950 ;
        RECT 299.400 721.050 300.450 722.400 ;
        RECT 304.950 721.800 307.050 723.900 ;
        RECT 295.950 719.400 300.450 721.050 ;
        RECT 295.950 718.950 300.000 719.400 ;
        RECT 311.400 715.050 312.450 730.950 ;
        RECT 317.400 730.200 318.450 733.950 ;
        RECT 316.950 728.100 319.050 730.200 ;
        RECT 325.950 728.250 328.050 730.350 ;
        RECT 334.950 728.250 337.050 730.350 ;
        RECT 340.950 728.250 343.050 730.350 ;
        RECT 317.400 727.350 318.600 728.100 ;
        RECT 316.950 724.950 319.050 727.050 ;
        RECT 319.950 724.950 322.050 727.050 ;
        RECT 320.400 723.900 321.600 724.650 ;
        RECT 319.950 721.800 322.050 723.900 ;
        RECT 326.400 721.050 327.450 728.250 ;
        RECT 335.400 727.500 336.600 728.250 ;
        RECT 341.400 727.500 342.600 728.250 ;
        RECT 331.950 725.100 334.050 727.200 ;
        RECT 334.950 725.100 337.050 727.200 ;
        RECT 337.950 725.100 340.050 727.200 ;
        RECT 340.950 725.100 343.050 727.200 ;
        RECT 332.400 722.400 333.600 724.800 ;
        RECT 338.400 724.050 339.600 724.800 ;
        RECT 325.950 718.950 328.050 721.050 ;
        RECT 292.950 714.450 295.050 715.050 ;
        RECT 290.400 713.400 295.050 714.450 ;
        RECT 283.950 703.950 286.050 706.050 ;
        RECT 277.950 700.950 280.050 703.050 ;
        RECT 278.400 694.050 279.450 700.950 ;
        RECT 277.950 691.950 280.050 694.050 ;
        RECT 286.950 691.950 289.050 694.050 ;
        RECT 268.950 685.950 271.050 688.050 ;
        RECT 248.400 682.350 249.600 684.600 ;
        RECT 253.950 683.100 256.050 685.200 ;
        RECT 271.950 683.100 274.050 685.200 ;
        RECT 254.400 682.350 255.600 683.100 ;
        RECT 272.400 682.350 273.600 683.100 ;
        RECT 277.950 682.950 280.050 685.050 ;
        RECT 287.400 684.600 288.450 691.950 ;
        RECT 290.400 685.050 291.450 713.400 ;
        RECT 292.950 712.950 295.050 713.400 ;
        RECT 310.950 712.950 313.050 715.050 ;
        RECT 292.950 709.800 295.050 711.900 ;
        RECT 293.400 691.050 294.450 709.800 ;
        RECT 332.400 709.050 333.450 722.400 ;
        RECT 337.950 721.950 340.050 724.050 ;
        RECT 304.950 706.950 307.050 709.050 ;
        RECT 331.950 706.950 334.050 709.050 ;
        RECT 292.950 688.950 295.050 691.050 ;
        RECT 247.950 679.950 250.050 682.050 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 256.950 679.950 259.050 682.050 ;
        RECT 265.950 679.950 268.050 682.050 ;
        RECT 271.950 679.950 274.050 682.050 ;
        RECT 251.400 677.400 252.600 679.650 ;
        RECT 257.400 678.900 258.600 679.650 ;
        RECT 241.950 661.950 244.050 664.050 ;
        RECT 238.950 658.950 241.050 661.050 ;
        RECT 251.400 654.450 252.450 677.400 ;
        RECT 256.950 673.950 259.050 678.900 ;
        RECT 259.950 658.950 262.050 661.050 ;
        RECT 251.400 653.400 255.450 654.450 ;
        RECT 254.400 652.350 255.450 653.400 ;
        RECT 235.950 650.100 238.050 652.200 ;
        RECT 236.400 649.350 237.600 650.100 ;
        RECT 244.950 649.950 247.050 652.050 ;
        RECT 253.950 650.250 256.050 652.350 ;
        RECT 260.400 651.600 261.450 658.950 ;
        RECT 278.400 658.050 279.450 682.950 ;
        RECT 287.400 682.200 288.600 684.600 ;
        RECT 289.800 682.950 291.900 685.050 ;
        RECT 292.950 682.950 295.050 685.050 ;
        RECT 298.950 682.950 301.050 685.050 ;
        RECT 305.400 684.600 306.450 706.950 ;
        RECT 310.950 697.950 313.050 700.050 ;
        RECT 311.400 685.050 312.450 697.950 ;
        RECT 347.400 697.050 348.450 739.950 ;
        RECT 371.400 739.050 372.450 754.950 ;
        RECT 373.950 748.950 376.050 751.050 ;
        RECT 349.950 736.950 352.050 739.050 ;
        RECT 370.950 736.950 373.050 739.050 ;
        RECT 350.400 723.900 351.450 736.950 ;
        RECT 358.950 733.950 361.050 736.050 ;
        RECT 359.400 729.600 360.450 733.950 ;
        RECT 374.400 730.050 375.450 748.950 ;
        RECT 377.400 739.050 378.450 755.400 ;
        RECT 376.950 736.950 379.050 739.050 ;
        RECT 386.400 736.050 387.450 760.950 ;
        RECT 395.400 760.200 396.600 762.000 ;
        RECT 400.950 760.950 403.050 763.050 ;
        RECT 410.400 762.600 411.450 769.950 ;
        RECT 401.400 760.200 402.600 760.950 ;
        RECT 410.400 760.200 411.600 762.600 ;
        RECT 416.400 762.450 417.600 762.600 ;
        RECT 419.400 762.450 420.450 799.950 ;
        RECT 422.400 790.050 423.450 800.400 ;
        RECT 430.950 799.950 433.050 802.050 ;
        RECT 437.400 801.900 438.600 802.650 ;
        RECT 436.950 799.800 439.050 801.900 ;
        RECT 448.950 799.950 451.050 802.050 ;
        RECT 455.400 800.400 456.600 802.650 ;
        RECT 433.950 793.950 436.050 796.050 ;
        RECT 421.950 787.950 424.050 790.050 ;
        RECT 422.400 772.050 423.450 787.950 ;
        RECT 434.400 781.050 435.450 793.950 ;
        RECT 437.400 793.050 438.450 799.800 ;
        RECT 439.950 793.950 442.050 796.050 ;
        RECT 436.950 790.950 439.050 793.050 ;
        RECT 440.400 790.050 441.450 793.950 ;
        RECT 439.950 787.950 442.050 790.050 ;
        RECT 433.950 778.950 436.050 781.050 ;
        RECT 421.950 769.950 424.050 772.050 ;
        RECT 427.950 769.950 430.050 775.050 ;
        RECT 421.950 763.950 424.050 766.050 ;
        RECT 416.400 761.400 420.450 762.450 ;
        RECT 416.400 760.200 417.600 761.400 ;
        RECT 391.950 757.800 394.050 759.900 ;
        RECT 394.950 757.800 397.050 759.900 ;
        RECT 397.950 757.800 400.050 759.900 ;
        RECT 400.950 757.800 403.050 759.900 ;
        RECT 409.950 757.800 412.050 759.900 ;
        RECT 412.950 757.800 415.050 759.900 ;
        RECT 415.950 757.800 418.050 759.900 ;
        RECT 392.400 756.750 393.600 757.500 ;
        RECT 398.400 756.750 399.600 757.500 ;
        RECT 391.950 754.650 394.050 756.750 ;
        RECT 397.950 754.650 400.050 756.750 ;
        RECT 403.950 754.950 406.050 757.050 ;
        RECT 413.400 755.400 414.600 757.500 ;
        RECT 404.400 751.050 405.450 754.950 ;
        RECT 403.950 748.950 406.050 751.050 ;
        RECT 394.950 745.950 397.050 748.050 ;
        RECT 386.400 734.400 391.050 736.050 ;
        RECT 387.000 733.950 391.050 734.400 ;
        RECT 395.400 730.200 396.450 745.950 ;
        RECT 413.400 745.050 414.450 755.400 ;
        RECT 422.400 745.050 423.450 763.950 ;
        RECT 449.400 763.050 450.450 799.950 ;
        RECT 455.400 799.050 456.450 800.400 ;
        RECT 455.400 797.400 460.050 799.050 ;
        RECT 456.000 796.950 460.050 797.400 ;
        RECT 461.400 790.050 462.450 820.950 ;
        RECT 515.400 817.050 516.450 820.950 ;
        RECT 493.950 814.950 496.050 817.050 ;
        RECT 514.950 814.950 517.050 817.050 ;
        RECT 490.950 811.800 493.050 813.900 ;
        RECT 469.950 806.250 472.050 811.050 ;
        RECT 477.000 807.600 481.050 808.050 ;
        RECT 470.400 805.500 471.600 806.250 ;
        RECT 476.400 805.950 481.050 807.600 ;
        RECT 484.950 805.950 487.050 808.050 ;
        RECT 491.400 807.600 492.450 811.800 ;
        RECT 494.400 811.050 495.450 814.950 ;
        RECT 532.950 811.950 535.050 814.050 ;
        RECT 544.950 811.950 547.050 814.050 ;
        RECT 493.950 808.950 496.050 811.050 ;
        RECT 476.400 805.500 477.600 805.950 ;
        RECT 466.950 803.100 469.050 805.200 ;
        RECT 469.950 803.100 472.050 805.200 ;
        RECT 472.950 803.100 475.050 805.200 ;
        RECT 475.950 803.100 478.050 805.200 ;
        RECT 467.400 800.400 468.600 802.800 ;
        RECT 473.400 801.000 474.600 802.800 ;
        RECT 460.950 787.950 463.050 790.050 ;
        RECT 467.400 766.050 468.450 800.400 ;
        RECT 472.950 796.950 475.050 801.000 ;
        RECT 475.950 799.950 478.050 802.050 ;
        RECT 476.400 766.050 477.450 799.950 ;
        RECT 485.400 799.050 486.450 805.950 ;
        RECT 491.400 805.500 492.600 807.600 ;
        RECT 496.950 806.250 499.050 808.350 ;
        RECT 511.950 806.250 514.050 808.350 ;
        RECT 517.950 806.250 520.050 808.350 ;
        RECT 497.400 805.500 498.600 806.250 ;
        RECT 512.400 805.500 513.600 806.250 ;
        RECT 518.400 805.500 519.600 806.250 ;
        RECT 523.950 805.950 526.050 808.050 ;
        RECT 533.400 807.600 534.450 811.950 ;
        RECT 540.000 807.600 544.050 808.050 ;
        RECT 490.950 803.100 493.050 805.200 ;
        RECT 493.950 803.100 496.050 805.200 ;
        RECT 496.950 803.100 499.050 805.200 ;
        RECT 499.950 803.100 502.050 805.200 ;
        RECT 508.950 803.100 511.050 805.200 ;
        RECT 511.950 803.100 514.050 805.200 ;
        RECT 514.950 803.100 517.050 805.200 ;
        RECT 517.950 803.100 520.050 805.200 ;
        RECT 494.400 801.000 495.600 802.800 ;
        RECT 484.950 796.950 487.050 799.050 ;
        RECT 493.950 796.950 496.050 801.000 ;
        RECT 500.400 800.400 501.600 802.800 ;
        RECT 500.400 799.050 501.450 800.400 ;
        RECT 505.950 799.950 508.050 802.050 ;
        RECT 509.400 800.400 510.600 802.800 ;
        RECT 481.950 793.950 484.050 796.050 ;
        RECT 478.950 778.950 481.050 781.050 ;
        RECT 479.400 775.050 480.450 778.950 ;
        RECT 478.950 772.950 481.050 775.050 ;
        RECT 482.400 772.050 483.450 793.950 ;
        RECT 493.950 793.800 496.050 795.900 ;
        RECT 499.950 793.950 502.050 799.050 ;
        RECT 506.400 795.450 507.450 799.950 ;
        RECT 509.400 796.050 510.450 800.400 ;
        RECT 511.950 799.950 514.050 802.050 ;
        RECT 515.400 800.400 516.600 802.800 ;
        RECT 524.400 802.050 525.450 805.950 ;
        RECT 533.400 805.500 534.600 807.600 ;
        RECT 539.400 805.950 544.050 807.600 ;
        RECT 539.400 805.500 540.600 805.950 ;
        RECT 529.950 803.100 532.050 805.200 ;
        RECT 532.950 803.100 535.050 805.200 ;
        RECT 535.950 803.100 538.050 805.200 ;
        RECT 538.950 803.100 541.050 805.200 ;
        RECT 508.950 795.450 511.050 796.050 ;
        RECT 506.400 794.400 511.050 795.450 ;
        RECT 508.950 793.950 511.050 794.400 ;
        RECT 484.950 790.950 487.050 793.050 ;
        RECT 485.400 778.050 486.450 790.950 ;
        RECT 494.400 790.050 495.450 793.800 ;
        RECT 493.800 787.950 495.900 790.050 ;
        RECT 496.950 787.950 499.050 790.050 ;
        RECT 497.400 784.050 498.450 787.950 ;
        RECT 496.950 781.950 499.050 784.050 ;
        RECT 512.400 781.050 513.450 799.950 ;
        RECT 515.400 799.050 516.450 800.400 ;
        RECT 517.950 799.950 520.050 802.050 ;
        RECT 523.950 799.950 526.050 802.050 ;
        RECT 530.400 800.400 531.600 802.800 ;
        RECT 536.400 801.000 537.600 802.800 ;
        RECT 514.950 796.950 517.050 799.050 ;
        RECT 515.400 787.050 516.450 796.950 ;
        RECT 514.950 784.950 517.050 787.050 ;
        RECT 511.950 778.950 514.050 781.050 ;
        RECT 484.950 775.950 487.050 778.050 ;
        RECT 505.950 775.950 508.050 778.050 ;
        RECT 481.950 769.950 484.050 772.050 ;
        RECT 487.950 769.950 490.050 772.050 ;
        RECT 481.950 766.800 484.050 768.900 ;
        RECT 427.950 760.950 430.050 763.050 ;
        RECT 433.950 760.950 436.050 763.050 ;
        RECT 448.950 760.950 451.050 763.050 ;
        RECT 454.950 762.000 457.050 766.050 ;
        RECT 460.950 762.000 463.050 766.050 ;
        RECT 466.950 763.950 469.050 766.050 ;
        RECT 475.950 763.950 478.050 766.050 ;
        RECT 428.400 760.200 429.600 760.950 ;
        RECT 434.400 760.200 435.600 760.950 ;
        RECT 455.400 760.200 456.600 762.000 ;
        RECT 461.400 760.200 462.600 762.000 ;
        RECT 427.950 757.800 430.050 759.900 ;
        RECT 430.950 757.800 433.050 759.900 ;
        RECT 433.950 757.800 436.050 759.900 ;
        RECT 436.950 757.800 439.050 759.900 ;
        RECT 451.950 757.800 454.050 759.900 ;
        RECT 454.950 757.800 457.050 759.900 ;
        RECT 457.950 757.800 460.050 759.900 ;
        RECT 460.950 757.800 463.050 759.900 ;
        RECT 424.950 754.950 427.050 757.050 ;
        RECT 431.400 755.400 432.600 757.500 ;
        RECT 437.400 755.400 438.600 757.500 ;
        RECT 452.400 756.000 453.600 757.500 ;
        RECT 458.400 756.750 459.600 757.500 ;
        RECT 425.400 751.050 426.450 754.950 ;
        RECT 424.950 748.950 427.050 751.050 ;
        RECT 412.950 742.950 415.050 745.050 ;
        RECT 421.950 742.950 424.050 745.050 ;
        RECT 406.950 733.950 409.050 736.050 ;
        RECT 359.400 727.350 360.600 729.600 ;
        RECT 365.400 729.450 366.600 729.600 ;
        RECT 365.400 728.400 372.450 729.450 ;
        RECT 365.400 727.350 366.600 728.400 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 358.950 724.950 361.050 727.050 ;
        RECT 361.950 724.950 364.050 727.050 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 356.400 723.900 357.600 724.650 ;
        RECT 349.950 721.800 352.050 723.900 ;
        RECT 355.950 721.800 358.050 723.900 ;
        RECT 362.400 722.400 363.600 724.650 ;
        RECT 371.400 723.450 372.450 728.400 ;
        RECT 373.950 727.950 376.050 730.050 ;
        RECT 379.950 728.100 382.050 730.200 ;
        RECT 385.950 728.100 388.050 730.200 ;
        RECT 394.950 728.100 397.050 730.200 ;
        RECT 400.950 729.000 403.050 733.050 ;
        RECT 407.400 730.050 408.450 733.950 ;
        RECT 409.950 730.950 412.050 733.050 ;
        RECT 380.400 727.350 381.600 728.100 ;
        RECT 386.400 727.350 387.600 728.100 ;
        RECT 395.400 727.350 396.600 728.100 ;
        RECT 401.400 727.350 402.600 729.000 ;
        RECT 406.950 727.950 409.050 730.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 379.950 724.950 382.050 727.050 ;
        RECT 382.950 724.950 385.050 727.050 ;
        RECT 385.950 724.950 388.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 400.950 724.950 403.050 727.050 ;
        RECT 403.950 724.950 406.050 727.050 ;
        RECT 377.400 723.900 378.600 724.650 ;
        RECT 368.400 722.400 372.450 723.450 ;
        RECT 362.400 721.050 363.450 722.400 ;
        RECT 362.400 718.950 367.050 721.050 ;
        RECT 355.800 712.950 357.900 715.050 ;
        RECT 358.950 712.950 361.050 715.050 ;
        RECT 337.950 694.950 340.050 697.050 ;
        RECT 346.950 694.950 349.050 697.050 ;
        RECT 313.950 691.950 316.050 694.050 ;
        RECT 293.400 682.200 294.600 682.950 ;
        RECT 286.950 679.800 289.050 681.900 ;
        RECT 289.950 679.800 292.050 681.900 ;
        RECT 292.950 679.800 295.050 681.900 ;
        RECT 290.400 678.750 291.600 679.500 ;
        RECT 289.950 676.650 292.050 678.750 ;
        RECT 295.950 673.950 298.050 676.050 ;
        RECT 296.400 670.050 297.450 673.950 ;
        RECT 299.400 673.050 300.450 682.950 ;
        RECT 305.400 682.200 306.600 684.600 ;
        RECT 310.950 682.950 313.050 685.050 ;
        RECT 314.400 684.600 315.450 691.950 ;
        RECT 319.950 688.950 322.050 691.050 ;
        RECT 320.400 685.050 321.450 688.950 ;
        RECT 314.400 682.200 315.600 684.600 ;
        RECT 319.800 682.950 321.900 685.050 ;
        RECT 322.950 682.950 325.050 685.050 ;
        RECT 328.950 684.000 331.050 688.050 ;
        RECT 323.400 682.200 324.600 682.950 ;
        RECT 329.400 682.200 330.600 684.000 ;
        RECT 304.950 679.800 307.050 681.900 ;
        RECT 307.950 679.800 310.050 681.900 ;
        RECT 313.950 679.800 316.050 681.900 ;
        RECT 322.950 679.800 325.050 681.900 ;
        RECT 325.950 679.800 328.050 681.900 ;
        RECT 328.950 679.800 331.050 681.900 ;
        RECT 331.950 679.800 334.050 681.900 ;
        RECT 308.400 677.400 309.600 679.500 ;
        RECT 308.400 673.050 309.450 677.400 ;
        RECT 310.950 676.950 313.050 679.050 ;
        RECT 316.950 676.950 319.050 679.050 ;
        RECT 326.400 677.400 327.600 679.500 ;
        RECT 332.400 678.750 333.600 679.500 ;
        RECT 298.950 670.950 301.050 673.050 ;
        RECT 307.950 670.950 310.050 673.050 ;
        RECT 295.950 667.950 298.050 670.050 ;
        RECT 289.950 664.950 292.050 667.050 ;
        RECT 265.950 655.950 268.050 658.050 ;
        RECT 277.950 655.950 280.050 658.050 ;
        RECT 235.950 646.950 238.050 649.050 ;
        RECT 238.950 646.950 241.050 649.050 ;
        RECT 239.400 644.400 240.600 646.650 ;
        RECT 239.400 643.050 240.450 644.400 ;
        RECT 239.400 641.400 244.050 643.050 ;
        RECT 240.000 640.950 244.050 641.400 ;
        RECT 229.950 625.950 232.050 628.050 ;
        RECT 208.950 619.950 211.050 622.050 ;
        RECT 241.950 619.950 244.050 622.050 ;
        RECT 238.950 616.950 241.050 619.050 ;
        RECT 223.950 613.950 226.050 616.050 ;
        RECT 208.950 606.000 211.050 610.050 ;
        RECT 209.400 604.200 210.600 606.000 ;
        RECT 214.950 604.950 217.050 607.050 ;
        RECT 215.400 604.200 216.600 604.950 ;
        RECT 208.950 601.800 211.050 603.900 ;
        RECT 211.950 601.800 214.050 603.900 ;
        RECT 214.950 601.800 217.050 603.900 ;
        RECT 217.950 601.800 220.050 603.900 ;
        RECT 212.400 599.400 213.600 601.500 ;
        RECT 218.400 600.750 219.600 601.500 ;
        RECT 212.400 583.050 213.450 599.400 ;
        RECT 217.950 598.650 220.050 600.750 ;
        RECT 224.400 597.450 225.450 613.950 ;
        RECT 232.950 605.100 235.050 607.200 ;
        RECT 233.400 604.350 234.600 605.100 ;
        RECT 229.950 601.950 232.050 604.050 ;
        RECT 232.950 601.950 235.050 604.050 ;
        RECT 230.400 599.400 231.600 601.650 ;
        RECT 224.400 596.400 228.450 597.450 ;
        RECT 220.950 586.950 223.050 589.050 ;
        RECT 211.950 580.950 214.050 583.050 ;
        RECT 172.950 569.100 175.050 571.200 ;
        RECT 175.950 569.100 178.050 571.200 ;
        RECT 178.950 569.100 181.050 571.200 ;
        RECT 181.950 569.100 184.050 571.200 ;
        RECT 169.950 565.950 172.050 568.050 ;
        RECT 172.950 565.950 175.050 568.050 ;
        RECT 176.400 567.000 177.600 568.800 ;
        RECT 182.400 568.050 183.600 568.800 ;
        RECT 170.400 556.050 171.450 565.950 ;
        RECT 169.950 553.950 172.050 556.050 ;
        RECT 164.400 533.400 168.450 534.450 ;
        RECT 164.400 529.050 165.450 533.400 ;
        RECT 169.950 532.950 172.050 535.050 ;
        RECT 152.400 526.350 153.600 528.600 ;
        RECT 158.400 526.350 159.600 528.600 ;
        RECT 163.950 526.950 166.050 529.050 ;
        RECT 170.400 528.450 171.450 532.950 ;
        RECT 173.400 532.050 174.450 565.950 ;
        RECT 175.950 562.950 178.050 567.000 ;
        RECT 181.950 565.950 184.050 568.050 ;
        RECT 188.400 565.050 189.450 572.400 ;
        RECT 197.400 571.500 198.600 573.000 ;
        RECT 202.950 571.950 205.050 574.050 ;
        RECT 208.950 573.000 211.050 577.050 ;
        RECT 214.950 573.000 217.050 577.050 ;
        RECT 221.400 574.050 222.450 586.950 ;
        RECT 223.950 574.950 226.050 577.050 ;
        RECT 209.400 571.350 210.600 573.000 ;
        RECT 215.400 571.350 216.600 573.000 ;
        RECT 220.950 571.950 223.050 574.050 ;
        RECT 193.950 569.100 196.050 571.200 ;
        RECT 196.950 569.100 199.050 571.200 ;
        RECT 199.950 569.100 202.050 571.200 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 214.950 568.950 217.050 571.050 ;
        RECT 217.950 568.950 220.050 571.050 ;
        RECT 194.400 567.450 195.600 568.800 ;
        RECT 200.400 568.050 201.600 568.800 ;
        RECT 191.400 566.400 195.600 567.450 ;
        RECT 187.950 562.950 190.050 565.050 ;
        RECT 176.400 553.050 177.450 562.950 ;
        RECT 187.950 559.800 190.050 561.900 ;
        RECT 184.950 556.950 187.050 559.050 ;
        RECT 175.950 550.950 178.050 553.050 ;
        RECT 175.950 544.950 178.050 547.050 ;
        RECT 172.950 529.950 175.050 532.050 ;
        RECT 167.400 527.400 171.450 528.450 ;
        RECT 173.400 528.450 174.600 528.600 ;
        RECT 176.400 528.450 177.450 544.950 ;
        RECT 178.950 532.950 181.050 535.050 ;
        RECT 173.400 527.400 177.450 528.450 ;
        RECT 179.400 528.600 180.450 532.950 ;
        RECT 185.400 528.600 186.450 556.950 ;
        RECT 188.400 529.050 189.450 559.800 ;
        RECT 191.400 550.050 192.450 566.400 ;
        RECT 199.800 565.950 201.900 568.050 ;
        RECT 202.950 565.950 205.050 568.050 ;
        RECT 212.400 566.400 213.600 568.650 ;
        RECT 218.400 567.900 219.600 568.650 ;
        RECT 199.950 556.950 202.050 559.050 ;
        RECT 200.400 553.050 201.450 556.950 ;
        RECT 199.950 550.950 202.050 553.050 ;
        RECT 190.950 547.950 193.050 550.050 ;
        RECT 193.950 544.950 196.050 547.050 ;
        RECT 190.950 541.950 193.050 544.050 ;
        RECT 191.400 532.050 192.450 541.950 ;
        RECT 194.400 538.050 195.450 544.950 ;
        RECT 203.400 544.050 204.450 565.950 ;
        RECT 208.950 559.950 211.050 562.050 ;
        RECT 202.950 541.950 205.050 544.050 ;
        RECT 193.950 535.950 196.050 538.050 ;
        RECT 202.950 532.950 205.050 535.050 ;
        RECT 190.950 529.950 193.050 532.050 ;
        RECT 148.950 523.950 151.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 145.950 520.950 148.050 523.050 ;
        RECT 149.400 521.400 150.600 523.650 ;
        RECT 155.400 522.900 156.600 523.650 ;
        RECT 130.950 513.450 133.050 514.050 ;
        RECT 125.400 512.400 133.050 513.450 ;
        RECT 130.950 511.950 133.050 512.400 ;
        RECT 142.950 511.950 145.050 514.050 ;
        RECT 124.950 502.950 127.050 505.050 ;
        RECT 118.950 493.950 121.050 496.050 ;
        RECT 125.400 495.600 126.450 502.950 ;
        RECT 146.400 502.050 147.450 520.950 ;
        RECT 149.400 505.050 150.450 521.400 ;
        RECT 154.950 520.800 157.050 522.900 ;
        RECT 160.950 520.950 163.050 523.050 ;
        RECT 161.400 508.050 162.450 520.950 ;
        RECT 167.400 520.050 168.450 527.400 ;
        RECT 173.400 526.200 174.600 527.400 ;
        RECT 179.400 526.200 180.600 528.600 ;
        RECT 185.400 526.200 186.600 528.600 ;
        RECT 187.950 526.950 190.050 529.050 ;
        RECT 193.950 526.950 196.050 529.050 ;
        RECT 203.400 528.600 204.450 532.950 ;
        RECT 194.400 526.200 195.600 526.950 ;
        RECT 203.400 526.200 204.600 528.600 ;
        RECT 172.950 523.800 175.050 525.900 ;
        RECT 175.950 523.800 178.050 525.900 ;
        RECT 178.950 523.800 181.050 525.900 ;
        RECT 181.950 523.800 184.050 525.900 ;
        RECT 184.950 523.800 187.050 525.900 ;
        RECT 193.950 523.800 196.050 525.900 ;
        RECT 199.950 523.800 202.050 525.900 ;
        RECT 202.950 523.800 205.050 525.900 ;
        RECT 176.400 522.750 177.600 523.500 ;
        RECT 182.400 522.750 183.600 523.500 ;
        RECT 175.950 520.650 178.050 522.750 ;
        RECT 181.950 520.650 184.050 522.750 ;
        RECT 200.400 521.400 201.600 523.500 ;
        RECT 166.950 517.950 169.050 520.050 ;
        RECT 176.400 517.050 177.450 520.650 ;
        RECT 175.950 514.950 178.050 517.050 ;
        RECT 154.950 505.950 157.050 508.050 ;
        RECT 160.800 505.950 162.900 508.050 ;
        RECT 148.950 502.950 151.050 505.050 ;
        RECT 145.950 499.950 148.050 502.050 ;
        RECT 125.400 493.350 126.600 495.600 ;
        RECT 130.950 494.250 133.050 496.350 ;
        RECT 139.950 494.250 142.050 496.350 ;
        RECT 146.400 495.600 147.450 499.950 ;
        RECT 155.400 496.050 156.450 505.950 ;
        RECT 169.950 499.950 172.050 502.050 ;
        RECT 121.950 490.950 124.050 493.050 ;
        RECT 124.950 490.950 127.050 493.050 ;
        RECT 106.950 487.800 109.050 489.900 ;
        RECT 115.950 487.950 118.050 490.050 ;
        RECT 122.400 489.900 123.600 490.650 ;
        RECT 121.950 487.800 124.050 489.900 ;
        RECT 97.950 481.950 100.050 484.050 ;
        RECT 131.400 478.050 132.450 494.250 ;
        RECT 140.400 493.500 141.600 494.250 ;
        RECT 146.400 493.500 147.600 495.600 ;
        RECT 154.950 493.950 157.050 496.050 ;
        RECT 160.950 494.250 163.050 496.350 ;
        RECT 161.400 493.500 162.600 494.250 ;
        RECT 136.950 491.100 139.050 493.200 ;
        RECT 139.950 491.100 142.050 493.200 ;
        RECT 142.950 491.100 145.050 493.200 ;
        RECT 145.950 491.100 148.050 493.200 ;
        RECT 148.950 491.100 151.050 493.200 ;
        RECT 157.950 491.100 160.050 493.200 ;
        RECT 160.950 491.100 163.050 493.200 ;
        RECT 163.950 491.100 166.050 493.200 ;
        RECT 137.400 488.400 138.600 490.800 ;
        RECT 143.400 489.000 144.600 490.800 ;
        RECT 149.400 490.050 150.600 490.800 ;
        RECT 158.400 490.050 159.600 490.800 ;
        RECT 164.400 490.050 165.600 490.800 ;
        RECT 170.400 490.050 171.450 499.950 ;
        RECT 182.400 499.050 183.450 520.650 ;
        RECT 200.400 517.050 201.450 521.400 ;
        RECT 205.950 519.450 208.050 523.050 ;
        RECT 203.400 519.000 208.050 519.450 ;
        RECT 203.400 518.400 207.450 519.000 ;
        RECT 199.950 514.950 202.050 517.050 ;
        RECT 190.950 511.950 193.050 514.050 ;
        RECT 178.800 498.000 180.900 499.050 ;
        RECT 178.800 496.950 181.050 498.000 ;
        RECT 181.950 496.950 184.050 499.050 ;
        RECT 178.950 494.250 181.050 496.950 ;
        RECT 179.400 493.500 180.600 494.250 ;
        RECT 175.950 491.100 178.050 493.200 ;
        RECT 178.950 491.100 181.050 493.200 ;
        RECT 181.950 491.100 184.050 493.200 ;
        RECT 191.400 493.050 192.450 511.950 ;
        RECT 203.400 511.050 204.450 518.400 ;
        RECT 209.400 514.050 210.450 559.950 ;
        RECT 212.400 556.050 213.450 566.400 ;
        RECT 217.950 565.800 220.050 567.900 ;
        RECT 220.950 565.950 223.050 568.050 ;
        RECT 211.950 553.950 214.050 556.050 ;
        RECT 211.950 550.800 214.050 552.900 ;
        RECT 212.400 529.050 213.450 550.800 ;
        RECT 217.950 538.950 220.050 541.050 ;
        RECT 218.400 529.050 219.450 538.950 ;
        RECT 221.400 535.050 222.450 565.950 ;
        RECT 224.400 562.050 225.450 574.950 ;
        RECT 227.400 571.050 228.450 596.400 ;
        RECT 230.400 589.050 231.450 599.400 ;
        RECT 229.950 586.950 232.050 589.050 ;
        RECT 239.400 580.050 240.450 616.950 ;
        RECT 242.400 589.050 243.450 619.950 ;
        RECT 245.400 610.050 246.450 649.950 ;
        RECT 254.400 649.500 255.600 650.250 ;
        RECT 260.400 649.500 261.600 651.600 ;
        RECT 250.950 647.100 253.050 649.200 ;
        RECT 253.950 647.100 256.050 649.200 ;
        RECT 256.950 647.100 259.050 649.200 ;
        RECT 259.950 647.100 262.050 649.200 ;
        RECT 247.950 643.950 250.050 646.050 ;
        RECT 251.400 644.400 252.600 646.800 ;
        RECT 257.400 645.000 258.600 646.800 ;
        RECT 248.400 637.050 249.450 643.950 ;
        RECT 251.400 640.050 252.450 644.400 ;
        RECT 256.950 640.950 259.050 645.000 ;
        RECT 250.950 637.950 253.050 640.050 ;
        RECT 256.950 637.800 259.050 639.900 ;
        RECT 247.950 634.950 250.050 637.050 ;
        RECT 244.950 607.950 247.050 610.050 ;
        RECT 248.400 607.050 249.450 634.950 ;
        RECT 250.950 613.950 253.050 616.050 ;
        RECT 251.400 610.050 252.450 613.950 ;
        RECT 257.400 610.050 258.450 637.800 ;
        RECT 262.950 625.950 265.050 628.050 ;
        RECT 247.950 604.950 250.050 607.050 ;
        RECT 250.950 606.000 253.050 610.050 ;
        RECT 256.950 607.950 259.050 610.050 ;
        RECT 257.400 606.600 258.450 607.950 ;
        RECT 251.400 604.200 252.600 606.000 ;
        RECT 257.400 604.200 258.600 606.600 ;
        RECT 247.950 601.800 250.050 603.900 ;
        RECT 250.950 601.800 253.050 603.900 ;
        RECT 253.950 601.800 256.050 603.900 ;
        RECT 256.950 601.800 259.050 603.900 ;
        RECT 244.950 598.950 247.050 601.050 ;
        RECT 248.400 599.400 249.600 601.500 ;
        RECT 254.400 600.750 255.600 601.500 ;
        RECT 245.400 592.050 246.450 598.950 ;
        RECT 244.950 589.950 247.050 592.050 ;
        RECT 241.950 586.950 244.050 589.050 ;
        RECT 238.950 577.950 241.050 580.050 ;
        RECT 242.400 576.450 243.450 586.950 ;
        RECT 244.950 577.950 247.050 580.050 ;
        RECT 239.400 575.400 243.450 576.450 ;
        RECT 232.950 572.250 235.050 574.350 ;
        RECT 239.400 573.600 240.450 575.400 ;
        RECT 245.400 574.050 246.450 577.950 ;
        RECT 248.400 574.050 249.450 599.400 ;
        RECT 253.950 598.650 256.050 600.750 ;
        RECT 259.950 598.950 262.050 601.050 ;
        RECT 260.400 592.050 261.450 598.950 ;
        RECT 263.400 592.050 264.450 625.950 ;
        RECT 266.400 619.050 267.450 655.950 ;
        RECT 271.950 647.100 274.050 649.200 ;
        RECT 277.950 647.100 280.050 649.200 ;
        RECT 280.950 647.100 283.050 649.200 ;
        RECT 268.950 642.450 271.050 646.050 ;
        RECT 272.400 645.450 273.600 646.800 ;
        RECT 272.400 645.000 276.450 645.450 ;
        RECT 272.400 644.400 277.050 645.000 ;
        RECT 268.950 642.000 273.450 642.450 ;
        RECT 269.400 641.400 273.450 642.000 ;
        RECT 272.400 637.050 273.450 641.400 ;
        RECT 274.950 640.950 277.050 644.400 ;
        RECT 281.400 644.400 282.600 646.800 ;
        RECT 268.800 634.950 270.900 637.050 ;
        RECT 271.950 634.950 274.050 637.050 ;
        RECT 269.400 628.050 270.450 634.950 ;
        RECT 268.950 625.950 271.050 628.050 ;
        RECT 275.400 625.050 276.450 640.950 ;
        RECT 277.950 637.950 280.050 640.050 ;
        RECT 278.400 634.050 279.450 637.950 ;
        RECT 281.400 634.050 282.450 644.400 ;
        RECT 277.800 631.950 279.900 634.050 ;
        RECT 280.950 631.950 283.050 634.050 ;
        RECT 274.950 622.950 277.050 625.050 ;
        RECT 290.400 622.050 291.450 664.950 ;
        RECT 298.950 650.250 301.050 652.350 ;
        RECT 311.400 652.050 312.450 676.950 ;
        RECT 299.400 649.500 300.600 650.250 ;
        RECT 307.800 649.950 309.900 652.050 ;
        RECT 310.950 649.950 313.050 652.050 ;
        RECT 317.400 651.600 318.450 676.950 ;
        RECT 326.400 667.050 327.450 677.400 ;
        RECT 331.950 676.650 334.050 678.750 ;
        RECT 332.400 673.050 333.450 676.650 ;
        RECT 331.950 670.950 334.050 673.050 ;
        RECT 325.950 664.950 328.050 667.050 ;
        RECT 331.950 664.950 334.050 667.050 ;
        RECT 322.950 658.950 325.050 661.050 ;
        RECT 323.400 651.600 324.450 658.950 ;
        RECT 325.950 655.950 328.050 658.050 ;
        RECT 326.400 652.050 327.450 655.950 ;
        RECT 328.950 652.950 331.050 655.050 ;
        RECT 295.950 647.100 298.050 649.200 ;
        RECT 298.950 647.100 301.050 649.200 ;
        RECT 301.950 647.100 304.050 649.200 ;
        RECT 302.400 644.400 303.600 646.800 ;
        RECT 308.400 645.900 309.450 649.950 ;
        RECT 317.400 649.350 318.600 651.600 ;
        RECT 323.400 649.350 324.600 651.600 ;
        RECT 325.950 649.950 328.050 652.050 ;
        RECT 313.950 646.950 316.050 649.050 ;
        RECT 316.950 646.950 319.050 649.050 ;
        RECT 319.950 646.950 322.050 649.050 ;
        RECT 322.950 646.950 325.050 649.050 ;
        RECT 314.400 645.900 315.600 646.650 ;
        RECT 302.400 643.050 303.450 644.400 ;
        RECT 307.950 643.800 310.050 645.900 ;
        RECT 313.950 643.800 316.050 645.900 ;
        RECT 320.400 644.400 321.600 646.650 ;
        RECT 301.950 640.950 304.050 643.050 ;
        RECT 292.950 628.950 295.050 631.050 ;
        RECT 293.400 622.050 294.450 628.950 ;
        RECT 274.950 619.800 277.050 621.900 ;
        RECT 289.800 619.950 291.900 622.050 ;
        RECT 292.950 619.950 295.050 622.050 ;
        RECT 265.950 616.950 268.050 619.050 ;
        RECT 268.950 605.100 271.050 607.200 ;
        RECT 275.400 606.600 276.450 619.800 ;
        RECT 302.400 616.050 303.450 640.950 ;
        RECT 310.950 637.950 313.050 640.050 ;
        RECT 307.950 631.950 310.050 634.050 ;
        RECT 304.950 625.950 307.050 628.050 ;
        RECT 286.950 613.950 289.050 616.050 ;
        RECT 301.950 613.950 304.050 616.050 ;
        RECT 277.950 607.950 280.050 613.050 ;
        RECT 287.400 606.600 288.450 613.950 ;
        RECT 269.400 604.350 270.600 605.100 ;
        RECT 275.400 604.350 276.600 606.600 ;
        RECT 287.400 604.200 288.600 606.600 ;
        RECT 292.950 604.950 295.050 610.050 ;
        RECT 293.400 604.200 294.600 604.950 ;
        RECT 268.950 601.950 271.050 604.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 274.950 601.950 277.050 604.050 ;
        RECT 277.950 601.950 280.050 604.050 ;
        RECT 286.950 601.800 289.050 603.900 ;
        RECT 289.950 601.800 292.050 603.900 ;
        RECT 292.950 601.800 295.050 603.900 ;
        RECT 295.950 601.800 298.050 603.900 ;
        RECT 272.400 599.400 273.600 601.650 ;
        RECT 278.400 599.400 279.600 601.650 ;
        RECT 290.400 600.750 291.600 601.500 ;
        RECT 259.800 589.950 261.900 592.050 ;
        RECT 262.950 589.950 265.050 592.050 ;
        RECT 268.950 589.950 271.050 592.050 ;
        RECT 233.400 571.500 234.600 572.250 ;
        RECT 239.400 571.500 240.600 573.600 ;
        RECT 244.800 571.950 246.900 574.050 ;
        RECT 247.950 571.950 250.050 574.050 ;
        RECT 253.950 572.250 256.050 574.350 ;
        RECT 260.400 574.050 261.450 589.950 ;
        RECT 262.950 586.800 265.050 588.900 ;
        RECT 254.400 571.500 255.600 572.250 ;
        RECT 259.950 571.950 262.050 574.050 ;
        RECT 226.950 568.950 229.050 571.050 ;
        RECT 232.950 569.100 235.050 571.200 ;
        RECT 235.950 569.100 238.050 571.200 ;
        RECT 238.950 569.100 241.050 571.200 ;
        RECT 241.950 569.100 244.050 571.200 ;
        RECT 250.950 569.100 253.050 571.200 ;
        RECT 253.950 569.100 256.050 571.200 ;
        RECT 256.950 569.100 259.050 571.200 ;
        RECT 226.950 565.800 229.050 567.900 ;
        RECT 232.950 565.950 235.050 568.050 ;
        RECT 236.400 566.400 237.600 568.800 ;
        RECT 242.400 568.050 243.600 568.800 ;
        RECT 251.400 568.050 252.600 568.800 ;
        RECT 257.400 568.050 258.600 568.800 ;
        RECT 263.400 568.050 264.450 586.800 ;
        RECT 265.950 583.950 268.050 586.050 ;
        RECT 223.950 559.950 226.050 562.050 ;
        RECT 227.400 541.050 228.450 565.800 ;
        RECT 226.950 538.950 229.050 541.050 ;
        RECT 226.950 535.800 229.050 537.900 ;
        RECT 220.950 532.950 223.050 535.050 ;
        RECT 211.950 526.950 214.050 529.050 ;
        RECT 214.950 526.950 217.050 529.050 ;
        RECT 217.950 526.950 220.050 529.050 ;
        RECT 221.400 528.600 222.450 532.950 ;
        RECT 215.400 526.200 216.600 526.950 ;
        RECT 221.400 526.200 222.600 528.600 ;
        RECT 214.950 523.800 217.050 525.900 ;
        RECT 217.950 523.800 220.050 525.900 ;
        RECT 220.950 523.800 223.050 525.900 ;
        RECT 211.950 520.950 214.050 523.050 ;
        RECT 218.400 522.750 219.600 523.500 ;
        RECT 208.950 511.950 211.050 514.050 ;
        RECT 202.950 508.950 205.050 511.050 ;
        RECT 199.950 502.950 202.050 505.050 ;
        RECT 193.950 493.950 196.050 499.050 ;
        RECT 200.400 495.600 201.450 502.950 ;
        RECT 203.400 499.050 204.450 508.950 ;
        RECT 205.950 499.950 208.050 502.050 ;
        RECT 202.950 496.950 205.050 499.050 ;
        RECT 206.400 496.050 207.450 499.950 ;
        RECT 212.400 498.450 213.450 520.950 ;
        RECT 217.950 520.650 220.050 522.750 ;
        RECT 223.950 520.950 226.050 523.050 ;
        RECT 224.400 508.050 225.450 520.950 ;
        RECT 223.950 505.950 226.050 508.050 ;
        RECT 227.400 504.450 228.450 535.800 ;
        RECT 233.400 528.450 234.450 565.950 ;
        RECT 236.400 562.050 237.450 566.400 ;
        RECT 241.950 565.950 244.050 568.050 ;
        RECT 250.950 565.950 253.050 568.050 ;
        RECT 256.950 565.950 259.050 568.050 ;
        RECT 259.950 565.950 262.050 568.050 ;
        RECT 262.950 565.950 265.050 568.050 ;
        RECT 238.950 562.950 241.050 565.050 ;
        RECT 235.950 559.950 238.050 562.050 ;
        RECT 239.400 538.050 240.450 562.950 ;
        RECT 241.950 559.950 244.050 562.050 ;
        RECT 238.950 535.950 241.050 538.050 ;
        RECT 242.400 529.050 243.450 559.950 ;
        RECT 260.400 553.050 261.450 565.950 ;
        RECT 259.950 550.950 262.050 553.050 ;
        RECT 262.950 547.950 265.050 550.050 ;
        RECT 250.950 538.950 253.050 541.050 ;
        RECT 230.400 527.400 234.450 528.450 ;
        RECT 230.400 505.050 231.450 527.400 ;
        RECT 238.800 526.950 240.900 529.050 ;
        RECT 241.950 526.950 244.050 529.050 ;
        RECT 246.000 528.600 250.050 529.050 ;
        RECT 245.400 526.950 250.050 528.600 ;
        RECT 239.400 526.200 240.600 526.950 ;
        RECT 245.400 526.200 246.600 526.950 ;
        RECT 235.950 523.800 238.050 525.900 ;
        RECT 238.950 523.800 241.050 525.900 ;
        RECT 241.950 523.800 244.050 525.900 ;
        RECT 244.950 523.800 247.050 525.900 ;
        RECT 236.400 521.400 237.600 523.500 ;
        RECT 242.400 521.400 243.600 523.500 ;
        RECT 236.400 507.450 237.450 521.400 ;
        RECT 238.950 517.950 241.050 520.050 ;
        RECT 233.400 506.400 237.450 507.450 ;
        RECT 224.400 503.400 228.450 504.450 ;
        RECT 209.400 497.400 213.450 498.450 ;
        RECT 200.400 493.500 201.600 495.600 ;
        RECT 205.950 493.950 208.050 496.050 ;
        RECT 190.950 490.950 193.050 493.050 ;
        RECT 196.950 491.100 199.050 493.200 ;
        RECT 199.950 491.100 202.050 493.200 ;
        RECT 202.950 491.100 205.050 493.200 ;
        RECT 130.950 475.950 133.050 478.050 ;
        RECT 97.950 469.950 100.050 472.050 ;
        RECT 109.950 469.950 112.050 472.050 ;
        RECT 79.950 459.450 82.050 460.050 ;
        RECT 79.950 458.400 84.450 459.450 ;
        RECT 79.950 457.950 82.050 458.400 ;
        RECT 70.950 453.450 73.050 454.050 ;
        RECT 68.400 452.400 73.050 453.450 ;
        RECT 56.400 448.200 57.600 450.000 ;
        RECT 62.400 448.200 63.600 450.600 ;
        RECT 64.950 448.950 67.050 451.050 ;
        RECT 52.950 445.800 55.050 447.900 ;
        RECT 55.950 445.800 58.050 447.900 ;
        RECT 58.950 445.800 61.050 447.900 ;
        RECT 61.950 445.800 64.050 447.900 ;
        RECT 53.400 443.400 54.600 445.500 ;
        RECT 59.400 444.750 60.600 445.500 ;
        RECT 68.400 444.750 69.450 452.400 ;
        RECT 70.950 451.950 73.050 452.400 ;
        RECT 76.950 451.950 79.050 454.050 ;
        RECT 77.400 450.450 78.600 450.600 ;
        RECT 79.950 450.450 82.050 454.050 ;
        RECT 77.400 450.000 82.050 450.450 ;
        RECT 83.400 450.600 84.450 458.400 ;
        RECT 94.950 457.950 97.050 460.050 ;
        RECT 77.400 449.400 81.450 450.000 ;
        RECT 77.400 448.200 78.600 449.400 ;
        RECT 83.400 448.200 84.600 450.600 ;
        RECT 85.950 448.950 88.050 454.050 ;
        RECT 98.400 453.450 99.450 469.950 ;
        RECT 110.400 466.050 111.450 469.950 ;
        RECT 100.950 463.950 103.050 466.050 ;
        RECT 109.950 463.950 112.050 466.050 ;
        RECT 95.400 452.400 99.450 453.450 ;
        RECT 95.400 451.200 96.450 452.400 ;
        RECT 101.400 451.200 102.450 463.950 ;
        RECT 106.950 457.950 109.050 460.050 ;
        RECT 94.950 449.100 97.050 451.200 ;
        RECT 100.950 449.100 103.050 451.200 ;
        RECT 95.400 448.350 96.600 449.100 ;
        RECT 101.400 448.350 102.600 449.100 ;
        RECT 73.950 445.800 76.050 447.900 ;
        RECT 76.950 445.800 79.050 447.900 ;
        RECT 79.950 445.800 82.050 447.900 ;
        RECT 82.950 445.800 85.050 447.900 ;
        RECT 91.950 445.950 94.050 448.050 ;
        RECT 94.950 445.950 97.050 448.050 ;
        RECT 97.950 445.950 100.050 448.050 ;
        RECT 100.950 445.950 103.050 448.050 ;
        RECT 53.400 421.050 54.450 443.400 ;
        RECT 58.950 442.650 61.050 444.750 ;
        RECT 67.950 442.650 70.050 444.750 ;
        RECT 74.400 443.400 75.600 445.500 ;
        RECT 80.400 444.750 81.600 445.500 ;
        RECT 74.400 439.050 75.450 443.400 ;
        RECT 79.950 442.650 82.050 444.750 ;
        RECT 85.950 442.950 88.050 445.050 ;
        RECT 92.400 444.000 93.600 445.650 ;
        RECT 82.950 439.950 85.050 442.050 ;
        RECT 73.800 436.950 75.900 439.050 ;
        RECT 76.950 436.950 79.050 439.050 ;
        RECT 64.950 433.950 67.050 436.050 ;
        RECT 61.950 430.950 64.050 433.050 ;
        RECT 46.950 418.950 49.050 421.050 ;
        RECT 52.950 418.950 55.050 421.050 ;
        RECT 43.950 417.600 48.000 418.050 ;
        RECT 53.400 417.600 54.450 418.950 ;
        RECT 43.950 415.950 48.600 417.600 ;
        RECT 47.400 415.500 48.600 415.950 ;
        RECT 53.400 415.500 54.600 417.600 ;
        RECT 46.950 413.100 49.050 415.200 ;
        RECT 49.950 413.100 52.050 415.200 ;
        RECT 52.950 413.100 55.050 415.200 ;
        RECT 55.950 413.100 58.050 415.200 ;
        RECT 50.400 412.050 51.600 412.800 ;
        RECT 43.950 409.950 46.050 412.050 ;
        RECT 49.950 409.950 52.050 412.050 ;
        RECT 56.400 411.000 57.600 412.800 ;
        RECT 40.950 376.950 43.050 379.050 ;
        RECT 19.950 370.950 22.050 373.050 ;
        RECT 28.950 370.950 31.050 373.050 ;
        RECT 34.950 372.000 37.050 376.050 ;
        RECT 44.400 373.050 45.450 409.950 ;
        RECT 55.950 406.950 58.050 411.000 ;
        RECT 62.400 406.050 63.450 430.950 ;
        RECT 65.400 430.050 66.450 433.950 ;
        RECT 64.950 427.950 67.050 430.050 ;
        RECT 70.950 416.100 73.050 418.200 ;
        RECT 77.400 417.600 78.450 436.950 ;
        RECT 79.950 433.950 82.050 436.050 ;
        RECT 80.400 418.050 81.450 433.950 ;
        RECT 71.400 415.350 72.600 416.100 ;
        RECT 77.400 415.350 78.600 417.600 ;
        RECT 79.950 415.950 82.050 418.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 70.950 412.950 73.050 415.050 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 76.950 412.950 79.050 415.050 ;
        RECT 68.400 411.900 69.600 412.650 ;
        RECT 67.950 409.800 70.050 411.900 ;
        RECT 74.400 410.400 75.600 412.650 ;
        RECT 74.400 406.050 75.450 410.400 ;
        RECT 79.950 409.950 82.050 412.050 ;
        RECT 61.950 403.950 64.050 406.050 ;
        RECT 73.950 403.950 76.050 406.050 ;
        RECT 49.950 380.400 52.050 382.500 ;
        RECT 70.950 381.300 73.050 383.400 ;
        RECT 14.400 370.200 15.600 370.950 ;
        RECT 20.400 370.200 21.600 370.950 ;
        RECT 29.400 370.200 30.600 370.950 ;
        RECT 35.400 370.200 36.600 372.000 ;
        RECT 43.800 370.950 45.900 373.050 ;
        RECT 46.950 371.100 49.050 373.200 ;
        RECT 47.400 370.350 48.600 371.100 ;
        RECT 10.950 367.800 13.050 369.900 ;
        RECT 13.950 367.800 16.050 369.900 ;
        RECT 16.950 367.800 19.050 369.900 ;
        RECT 19.950 367.800 22.050 369.900 ;
        RECT 28.950 367.800 31.050 369.900 ;
        RECT 31.950 367.800 34.050 369.900 ;
        RECT 34.950 367.800 37.050 369.900 ;
        RECT 37.950 367.800 40.050 369.900 ;
        RECT 46.950 367.950 49.050 370.050 ;
        RECT 7.950 364.950 10.050 367.050 ;
        RECT 11.400 365.400 12.600 367.500 ;
        RECT 17.400 366.750 18.600 367.500 ;
        RECT 32.400 366.750 33.600 367.500 ;
        RECT 4.950 352.950 7.050 355.050 ;
        RECT 8.400 351.450 9.450 364.950 ;
        RECT 11.400 361.050 12.450 365.400 ;
        RECT 16.950 364.650 19.050 366.750 ;
        RECT 31.950 364.650 34.050 366.750 ;
        RECT 38.400 365.400 39.600 367.500 ;
        RECT 10.950 358.950 13.050 361.050 ;
        RECT 17.400 355.050 18.450 364.650 ;
        RECT 16.950 352.950 19.050 355.050 ;
        RECT 31.950 352.950 34.050 355.050 ;
        RECT 5.400 350.400 9.450 351.450 ;
        RECT 5.400 334.050 6.450 350.400 ;
        RECT 19.950 343.950 22.050 346.050 ;
        RECT 13.950 338.100 16.050 340.200 ;
        RECT 14.400 337.350 15.600 338.100 ;
        RECT 10.950 334.950 13.050 337.050 ;
        RECT 13.950 334.950 16.050 337.050 ;
        RECT 4.950 331.950 7.050 334.050 ;
        RECT 11.400 333.900 12.600 334.650 ;
        RECT 20.400 334.050 21.450 343.950 ;
        RECT 32.400 340.350 33.450 352.950 ;
        RECT 38.400 349.050 39.450 365.400 ;
        RECT 43.950 364.950 46.050 367.050 ;
        RECT 37.950 346.950 40.050 349.050 ;
        RECT 44.400 346.050 45.450 364.950 ;
        RECT 50.700 360.600 51.900 380.400 ;
        RECT 61.950 376.950 64.050 379.050 ;
        RECT 70.950 377.700 72.150 381.300 ;
        RECT 55.950 371.100 58.050 373.200 ;
        RECT 56.400 370.350 57.600 371.100 ;
        RECT 55.950 367.950 58.050 370.050 ;
        RECT 55.950 361.950 58.050 364.050 ;
        RECT 49.950 358.500 52.050 360.600 ;
        RECT 43.950 343.950 46.050 346.050 ;
        RECT 44.400 342.450 45.450 343.950 ;
        RECT 44.400 341.400 48.450 342.450 ;
        RECT 25.950 338.250 28.050 340.350 ;
        RECT 31.950 338.250 34.050 340.350 ;
        RECT 47.400 339.600 48.450 341.400 ;
        RECT 26.400 337.500 27.600 338.250 ;
        RECT 32.400 337.500 33.600 338.250 ;
        RECT 47.400 337.500 48.600 339.600 ;
        RECT 52.950 338.250 55.050 340.350 ;
        RECT 56.400 339.450 57.450 361.950 ;
        RECT 62.400 355.050 63.450 376.950 ;
        RECT 70.950 375.600 73.050 377.700 ;
        RECT 64.950 370.950 67.050 373.050 ;
        RECT 61.950 352.950 64.050 355.050 ;
        RECT 65.400 343.050 66.450 370.950 ;
        RECT 70.950 360.600 72.150 375.600 ;
        RECT 73.950 367.950 76.050 370.050 ;
        RECT 74.400 366.450 75.600 367.650 ;
        RECT 74.400 365.400 78.450 366.450 ;
        RECT 70.950 358.500 73.050 360.600 ;
        RECT 77.400 355.050 78.450 365.400 ;
        RECT 80.400 363.450 81.450 409.950 ;
        RECT 83.400 394.050 84.450 439.950 ;
        RECT 86.400 417.450 87.450 442.950 ;
        RECT 91.950 439.950 94.050 444.000 ;
        RECT 98.400 443.400 99.600 445.650 ;
        RECT 98.400 430.050 99.450 443.400 ;
        RECT 103.950 442.950 106.050 445.050 ;
        RECT 104.400 433.050 105.450 442.950 ;
        RECT 107.400 442.050 108.450 457.950 ;
        RECT 131.400 454.050 132.450 475.950 ;
        RECT 130.950 451.950 133.050 454.050 ;
        RECT 109.950 449.100 112.050 451.200 ;
        RECT 115.950 449.100 118.050 451.200 ;
        RECT 121.950 449.100 124.050 451.200 ;
        RECT 137.400 451.050 138.450 488.400 ;
        RECT 142.950 484.950 145.050 489.000 ;
        RECT 148.950 487.950 151.050 490.050 ;
        RECT 157.950 487.950 160.050 490.050 ;
        RECT 163.950 487.950 166.050 490.050 ;
        RECT 169.950 487.950 172.050 490.050 ;
        RECT 172.950 487.950 175.050 490.050 ;
        RECT 176.400 488.400 177.600 490.800 ;
        RECT 182.400 490.050 183.600 490.800 ;
        RECT 181.950 489.450 184.050 490.050 ;
        RECT 179.400 488.400 184.050 489.450 ;
        RECT 151.950 484.950 154.050 487.050 ;
        RECT 166.950 484.950 169.050 487.050 ;
        RECT 152.400 472.050 153.450 484.950 ;
        RECT 151.950 469.950 154.050 472.050 ;
        RECT 167.400 459.450 168.450 484.950 ;
        RECT 167.400 458.400 171.450 459.450 ;
        RECT 155.100 454.200 157.200 456.300 ;
        RECT 164.100 454.500 166.200 456.600 ;
        RECT 110.400 445.050 111.450 449.100 ;
        RECT 116.400 448.350 117.600 449.100 ;
        RECT 122.400 448.350 123.600 449.100 ;
        RECT 130.950 448.800 133.050 450.900 ;
        RECT 136.950 448.950 139.050 451.050 ;
        RECT 142.950 450.000 145.050 454.050 ;
        RECT 115.950 445.950 118.050 448.050 ;
        RECT 118.950 445.950 121.050 448.050 ;
        RECT 121.950 445.950 124.050 448.050 ;
        RECT 124.950 445.950 127.050 448.050 ;
        RECT 109.950 442.950 112.050 445.050 ;
        RECT 119.400 444.900 120.600 445.650 ;
        RECT 118.950 442.800 121.050 444.900 ;
        RECT 125.400 443.400 126.600 445.650 ;
        RECT 106.950 439.950 109.050 442.050 ;
        RECT 103.950 430.950 106.050 433.050 ;
        RECT 97.950 427.950 100.050 430.050 ;
        RECT 125.400 423.450 126.450 443.400 ;
        RECT 127.950 442.950 130.050 445.050 ;
        RECT 128.400 436.050 129.450 442.950 ;
        RECT 131.400 442.050 132.450 448.800 ;
        RECT 137.400 448.200 138.600 448.950 ;
        RECT 143.400 448.200 144.600 450.000 ;
        RECT 152.400 448.050 153.600 450.600 ;
        RECT 136.950 445.800 139.050 447.900 ;
        RECT 139.950 445.800 142.050 447.900 ;
        RECT 142.950 445.800 145.050 447.900 ;
        RECT 151.950 445.800 154.050 448.050 ;
        RECT 133.950 442.950 136.050 445.050 ;
        RECT 140.400 444.750 141.600 445.500 ;
        RECT 130.950 439.950 133.050 442.050 ;
        RECT 134.400 436.050 135.450 442.950 ;
        RECT 139.950 442.650 142.050 444.750 ;
        RECT 136.950 439.950 139.050 442.050 ;
        RECT 155.400 441.600 156.300 454.200 ;
        RECT 161.400 450.900 162.600 453.600 ;
        RECT 161.250 448.800 163.350 450.900 ;
        RECT 157.200 447.900 159.300 448.200 ;
        RECT 165.150 447.900 166.050 454.500 ;
        RECT 170.400 451.050 171.450 458.400 ;
        RECT 169.950 448.950 172.050 451.050 ;
        RECT 157.200 447.000 166.050 447.900 ;
        RECT 157.200 446.100 159.300 447.000 ;
        RECT 162.150 445.200 164.250 446.100 ;
        RECT 157.200 444.000 164.250 445.200 ;
        RECT 157.200 443.100 159.300 444.000 ;
        RECT 127.950 433.950 130.050 436.050 ;
        RECT 133.950 433.950 136.050 436.050 ;
        RECT 127.950 423.450 130.050 424.050 ;
        RECT 125.400 422.400 130.050 423.450 ;
        RECT 127.950 421.950 130.050 422.400 ;
        RECT 88.950 417.450 91.050 418.350 ;
        RECT 86.400 416.400 91.050 417.450 ;
        RECT 88.950 416.250 91.050 416.400 ;
        RECT 94.950 416.250 97.050 418.350 ;
        RECT 89.400 415.500 90.600 416.250 ;
        RECT 95.400 415.500 96.600 416.250 ;
        RECT 103.950 415.950 106.050 418.050 ;
        RECT 109.950 416.250 112.050 418.350 ;
        RECT 115.950 416.250 118.050 418.350 ;
        RECT 128.400 417.600 129.450 421.950 ;
        RECT 137.400 418.200 138.450 439.950 ;
        RECT 154.650 439.500 156.750 441.600 ;
        RECT 161.250 440.100 163.350 442.200 ;
        RECT 165.150 441.900 166.050 447.000 ;
        RECT 166.950 445.800 169.050 447.900 ;
        RECT 167.400 443.400 168.600 445.800 ;
        RECT 161.400 437.400 162.600 440.100 ;
        RECT 164.700 439.800 166.800 441.900 ;
        RECT 157.950 433.950 160.050 436.050 ;
        RECT 154.950 421.950 157.050 424.050 ;
        RECT 88.950 413.100 91.050 415.200 ;
        RECT 91.950 413.100 94.050 415.200 ;
        RECT 94.950 413.100 97.050 415.200 ;
        RECT 97.950 413.100 100.050 415.200 ;
        RECT 92.400 411.000 93.600 412.800 ;
        RECT 98.400 412.050 99.600 412.800 ;
        RECT 91.950 406.950 94.050 411.000 ;
        RECT 94.800 409.950 96.900 412.050 ;
        RECT 97.950 409.950 100.050 412.050 ;
        RECT 95.400 406.050 96.450 409.950 ;
        RECT 94.950 403.950 97.050 406.050 ;
        RECT 82.950 391.950 85.050 394.050 ;
        RECT 97.950 376.950 100.050 379.050 ;
        RECT 91.950 370.950 94.050 373.050 ;
        RECT 98.400 372.600 99.450 376.950 ;
        RECT 92.400 370.200 93.600 370.950 ;
        RECT 98.400 370.200 99.600 372.600 ;
        RECT 88.950 367.800 91.050 369.900 ;
        RECT 91.950 367.800 94.050 369.900 ;
        RECT 94.950 367.800 97.050 369.900 ;
        RECT 97.950 367.800 100.050 369.900 ;
        RECT 89.400 365.400 90.600 367.500 ;
        RECT 95.400 366.750 96.600 367.500 ;
        RECT 104.400 366.750 105.450 415.950 ;
        RECT 110.400 415.500 111.600 416.250 ;
        RECT 116.400 415.500 117.600 416.250 ;
        RECT 128.400 415.350 129.600 417.600 ;
        RECT 136.950 416.100 139.050 418.200 ;
        RECT 142.950 416.100 145.050 418.200 ;
        RECT 148.950 416.100 151.050 418.200 ;
        RECT 155.400 418.050 156.450 421.950 ;
        RECT 109.950 413.100 112.050 415.200 ;
        RECT 112.950 413.100 115.050 415.200 ;
        RECT 115.950 413.100 118.050 415.200 ;
        RECT 118.950 413.100 121.050 415.200 ;
        RECT 127.950 412.950 130.050 415.050 ;
        RECT 130.950 412.950 133.050 415.050 ;
        RECT 113.400 410.400 114.600 412.800 ;
        RECT 119.400 412.050 120.600 412.800 ;
        RECT 113.400 388.050 114.450 410.400 ;
        RECT 118.950 409.950 121.050 412.050 ;
        RECT 124.950 409.950 127.050 412.050 ;
        RECT 131.400 411.900 132.600 412.650 ;
        RECT 119.400 406.050 120.450 409.950 ;
        RECT 118.950 403.950 121.050 406.050 ;
        RECT 112.950 385.950 115.050 388.050 ;
        RECT 112.950 376.950 115.050 379.050 ;
        RECT 113.400 372.600 114.450 376.950 ;
        RECT 113.400 370.200 114.600 372.600 ;
        RECT 118.950 370.950 121.050 373.050 ;
        RECT 119.400 370.200 120.600 370.950 ;
        RECT 109.950 367.800 112.050 369.900 ;
        RECT 112.950 367.800 115.050 369.900 ;
        RECT 115.950 367.800 118.050 369.900 ;
        RECT 118.950 367.800 121.050 369.900 ;
        RECT 82.950 363.450 85.050 364.050 ;
        RECT 80.400 362.400 85.050 363.450 ;
        RECT 82.950 361.950 85.050 362.400 ;
        RECT 76.950 352.950 79.050 355.050 ;
        RECT 76.950 346.950 79.050 349.050 ;
        RECT 64.950 340.950 67.050 343.050 ;
        RECT 56.400 338.400 60.450 339.450 ;
        RECT 53.400 337.500 54.600 338.250 ;
        RECT 25.950 335.100 28.050 337.200 ;
        RECT 28.950 335.100 31.050 337.200 ;
        RECT 31.950 335.100 34.050 337.200 ;
        RECT 34.950 335.100 37.050 337.200 ;
        RECT 43.950 335.100 46.050 337.200 ;
        RECT 46.950 335.100 49.050 337.200 ;
        RECT 49.950 335.100 52.050 337.200 ;
        RECT 52.950 335.100 55.050 337.200 ;
        RECT 29.400 334.050 30.600 334.800 ;
        RECT 10.950 331.800 13.050 333.900 ;
        RECT 16.800 331.950 18.900 334.050 ;
        RECT 19.950 331.950 22.050 334.050 ;
        RECT 28.950 331.950 31.050 334.050 ;
        RECT 35.400 333.000 36.600 334.800 ;
        RECT 44.400 334.050 45.600 334.800 ;
        RECT 17.400 307.050 18.450 331.950 ;
        RECT 34.950 328.950 37.050 333.000 ;
        RECT 40.950 332.400 45.600 334.050 ;
        RECT 50.400 333.000 51.600 334.800 ;
        RECT 40.950 331.950 45.000 332.400 ;
        RECT 49.950 328.950 52.050 333.000 ;
        RECT 52.950 331.950 55.050 334.050 ;
        RECT 53.400 313.050 54.450 331.950 ;
        RECT 37.950 310.950 40.050 313.050 ;
        RECT 52.950 310.950 55.050 313.050 ;
        RECT 28.950 307.950 31.050 310.050 ;
        RECT 10.950 304.950 13.050 307.050 ;
        RECT 16.950 304.950 19.050 307.050 ;
        RECT 4.950 301.950 7.050 304.050 ;
        RECT 5.400 289.050 6.450 301.950 ;
        RECT 11.400 294.600 12.450 304.950 ;
        RECT 29.400 295.050 30.450 307.950 ;
        RECT 34.950 301.950 37.050 304.050 ;
        RECT 11.400 292.200 12.600 294.600 ;
        RECT 16.950 292.950 19.050 295.050 ;
        RECT 28.950 292.950 31.050 295.050 ;
        RECT 35.400 294.600 36.450 301.950 ;
        RECT 38.400 295.050 39.450 310.950 ;
        RECT 49.950 302.400 52.050 304.500 ;
        RECT 17.400 292.200 18.600 292.950 ;
        RECT 29.400 292.200 30.600 292.950 ;
        RECT 35.400 292.200 36.600 294.600 ;
        RECT 37.950 292.950 40.050 295.050 ;
        RECT 46.950 293.100 49.050 295.200 ;
        RECT 47.400 292.350 48.600 293.100 ;
        RECT 10.950 289.800 13.050 291.900 ;
        RECT 13.950 289.800 16.050 291.900 ;
        RECT 16.950 289.800 19.050 291.900 ;
        RECT 25.950 289.800 28.050 291.900 ;
        RECT 28.950 289.800 31.050 291.900 ;
        RECT 31.950 289.800 34.050 291.900 ;
        RECT 34.950 289.800 37.050 291.900 ;
        RECT 37.950 289.800 40.050 291.900 ;
        RECT 46.950 289.950 49.050 292.050 ;
        RECT 4.950 286.950 7.050 289.050 ;
        RECT 14.400 288.750 15.600 289.500 ;
        RECT 13.950 286.650 16.050 288.750 ;
        RECT 26.400 287.400 27.600 289.500 ;
        RECT 32.400 287.400 33.600 289.500 ;
        RECT 38.400 288.750 39.600 289.500 ;
        RECT 26.400 283.050 27.450 287.400 ;
        RECT 32.400 285.450 33.450 287.400 ;
        RECT 37.950 286.650 40.050 288.750 ;
        RECT 32.400 284.400 36.450 285.450 ;
        RECT 13.950 280.950 16.050 283.050 ;
        RECT 25.950 280.950 28.050 283.050 ;
        RECT 7.950 266.400 10.050 268.500 ;
        RECT 4.950 260.100 7.050 262.200 ;
        RECT 5.400 259.350 6.600 260.100 ;
        RECT 4.950 256.950 7.050 259.050 ;
        RECT 8.850 251.400 10.050 266.400 ;
        RECT 7.950 249.300 10.050 251.400 ;
        RECT 8.850 245.700 10.050 249.300 ;
        RECT 7.950 243.600 10.050 245.700 ;
        RECT 7.950 225.300 10.050 227.400 ;
        RECT 8.850 221.700 10.050 225.300 ;
        RECT 7.950 219.600 10.050 221.700 ;
        RECT 4.950 211.950 7.050 214.050 ;
        RECT 5.400 210.450 6.600 211.650 ;
        RECT 2.400 209.400 6.600 210.450 ;
        RECT 2.400 103.050 3.450 209.400 ;
        RECT 8.850 204.600 10.050 219.600 ;
        RECT 7.950 202.500 10.050 204.600 ;
        RECT 7.950 196.950 10.050 199.050 ;
        RECT 8.400 184.200 9.450 196.950 ;
        RECT 14.400 193.050 15.450 280.950 ;
        RECT 28.950 266.400 31.050 268.500 ;
        RECT 16.950 260.100 19.050 262.200 ;
        RECT 17.400 199.050 18.450 260.100 ;
        RECT 22.950 256.950 25.050 259.050 ;
        RECT 23.400 255.900 24.600 256.650 ;
        RECT 22.950 253.800 25.050 255.900 ;
        RECT 29.100 246.600 30.300 266.400 ;
        RECT 35.400 262.050 36.450 284.400 ;
        RECT 50.700 282.600 51.900 302.400 ;
        RECT 59.400 295.050 60.450 338.400 ;
        RECT 61.950 337.950 64.050 340.050 ;
        RECT 70.950 338.100 73.050 340.200 ;
        RECT 77.400 339.600 78.450 346.950 ;
        RECT 58.950 292.950 61.050 295.050 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 58.950 283.950 61.050 286.050 ;
        RECT 49.950 280.500 52.050 282.600 ;
        RECT 55.950 271.950 58.050 274.050 ;
        RECT 43.950 266.400 46.050 268.500 ;
        RECT 34.950 259.950 37.050 262.050 ;
        RECT 31.950 256.950 34.050 259.050 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 32.400 254.400 33.600 256.650 ;
        RECT 41.400 254.400 42.600 256.650 ;
        RECT 32.400 250.050 33.450 254.400 ;
        RECT 41.400 250.050 42.450 254.400 ;
        RECT 31.950 249.450 34.050 250.050 ;
        RECT 31.950 248.400 36.450 249.450 ;
        RECT 31.950 247.950 34.050 248.400 ;
        RECT 28.950 244.500 31.050 246.600 ;
        RECT 28.950 224.400 31.050 226.500 ;
        RECT 22.950 215.100 25.050 217.200 ;
        RECT 23.400 214.350 24.600 215.100 ;
        RECT 22.950 211.950 25.050 214.050 ;
        RECT 29.100 204.600 30.300 224.400 ;
        RECT 32.400 216.450 33.600 216.600 ;
        RECT 35.400 216.450 36.450 248.400 ;
        RECT 40.950 247.950 43.050 250.050 ;
        RECT 44.700 246.600 45.900 266.400 ;
        RECT 49.950 256.950 52.050 259.050 ;
        RECT 50.400 255.900 51.600 256.650 ;
        RECT 49.950 253.800 52.050 255.900 ;
        RECT 43.950 244.500 46.050 246.600 ;
        RECT 32.400 215.400 36.450 216.450 ;
        RECT 32.400 214.350 33.600 215.400 ;
        RECT 46.950 214.950 49.050 217.050 ;
        RECT 56.400 216.600 57.450 271.950 ;
        RECT 59.400 250.050 60.450 283.950 ;
        RECT 62.400 274.050 63.450 337.950 ;
        RECT 71.400 337.350 72.600 338.100 ;
        RECT 77.400 337.350 78.600 339.600 ;
        RECT 67.950 334.950 70.050 337.050 ;
        RECT 70.950 334.950 73.050 337.050 ;
        RECT 73.950 334.950 76.050 337.050 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 68.400 333.000 69.600 334.650 ;
        RECT 74.400 333.900 75.600 334.650 ;
        RECT 67.950 328.950 70.050 333.000 ;
        RECT 73.950 331.800 76.050 333.900 ;
        RECT 68.400 310.050 69.450 328.950 ;
        RECT 83.400 325.050 84.450 361.950 ;
        RECT 89.400 349.050 90.450 365.400 ;
        RECT 94.950 364.650 97.050 366.750 ;
        RECT 103.950 364.650 106.050 366.750 ;
        RECT 110.400 365.400 111.600 367.500 ;
        RECT 116.400 366.750 117.600 367.500 ;
        RECT 110.400 358.050 111.450 365.400 ;
        RECT 115.950 364.650 118.050 366.750 ;
        RECT 125.400 358.050 126.450 409.950 ;
        RECT 130.800 409.800 132.900 411.900 ;
        RECT 133.950 409.950 136.050 412.050 ;
        RECT 134.400 379.050 135.450 409.950 ;
        RECT 133.950 376.950 136.050 379.050 ;
        RECT 137.400 376.050 138.450 416.100 ;
        RECT 143.400 415.350 144.600 416.100 ;
        RECT 149.400 415.350 150.600 416.100 ;
        RECT 154.950 415.950 157.050 418.050 ;
        RECT 142.950 412.950 145.050 415.050 ;
        RECT 145.950 412.950 148.050 415.050 ;
        RECT 148.950 412.950 151.050 415.050 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 146.400 410.400 147.600 412.650 ;
        RECT 152.400 411.900 153.600 412.650 ;
        RECT 146.400 406.050 147.450 410.400 ;
        RECT 151.950 409.800 154.050 411.900 ;
        RECT 145.950 403.950 148.050 406.050 ;
        RECT 158.400 400.050 159.450 433.950 ;
        RECT 161.400 427.050 162.450 437.400 ;
        RECT 160.950 424.950 163.050 427.050 ;
        RECT 163.950 416.100 166.050 418.200 ;
        RECT 170.400 417.450 171.600 417.600 ;
        RECT 173.400 417.450 174.450 487.950 ;
        RECT 176.400 454.050 177.450 488.400 ;
        RECT 175.950 451.950 178.050 454.050 ;
        RECT 179.400 450.450 180.450 488.400 ;
        RECT 181.950 487.950 184.050 488.400 ;
        RECT 190.950 487.800 193.050 489.900 ;
        RECT 203.400 488.400 204.600 490.800 ;
        RECT 191.400 460.050 192.450 487.800 ;
        RECT 203.400 481.050 204.450 488.400 ;
        RECT 205.950 487.950 208.050 490.050 ;
        RECT 202.950 478.950 205.050 481.050 ;
        RECT 206.400 466.050 207.450 487.950 ;
        RECT 205.950 463.950 208.050 466.050 ;
        RECT 190.950 457.950 193.050 460.050 ;
        RECT 205.950 457.950 208.050 460.050 ;
        RECT 176.400 449.400 180.450 450.450 ;
        RECT 187.950 450.000 190.050 454.050 ;
        RECT 176.400 444.750 177.450 449.400 ;
        RECT 188.400 448.200 189.600 450.000 ;
        RECT 196.950 448.950 199.050 451.050 ;
        RECT 206.400 450.600 207.450 457.950 ;
        RECT 209.400 451.050 210.450 497.400 ;
        RECT 217.200 497.100 219.300 499.200 ;
        RECT 221.400 498.900 222.600 501.600 ;
        RECT 215.400 493.200 216.600 495.600 ;
        RECT 214.950 493.050 217.050 493.200 ;
        RECT 211.950 491.100 217.050 493.050 ;
        RECT 217.950 492.000 218.850 497.100 ;
        RECT 220.650 496.800 223.050 498.900 ;
        RECT 224.400 495.900 225.450 503.400 ;
        RECT 229.950 502.950 232.050 505.050 ;
        RECT 233.400 502.050 234.450 506.400 ;
        RECT 235.950 502.950 238.050 505.050 ;
        RECT 232.950 499.950 235.050 502.050 ;
        RECT 227.250 497.400 229.350 499.500 ;
        RECT 224.400 495.000 226.800 495.900 ;
        RECT 219.750 493.800 226.800 495.000 ;
        RECT 219.750 492.900 221.850 493.800 ;
        RECT 224.700 492.000 226.800 492.900 ;
        RECT 217.950 491.100 226.800 492.000 ;
        RECT 211.950 490.950 214.950 491.100 ;
        RECT 217.950 484.500 218.850 491.100 ;
        RECT 224.700 490.800 226.800 491.100 ;
        RECT 220.650 488.100 222.750 490.200 ;
        RECT 221.400 485.400 222.600 488.100 ;
        RECT 227.700 484.800 228.600 497.400 ;
        RECT 236.400 496.050 237.450 502.950 ;
        RECT 235.950 493.950 238.050 496.050 ;
        RECT 239.400 495.600 240.450 517.950 ;
        RECT 242.400 517.050 243.450 521.400 ;
        RECT 241.950 514.950 244.050 517.050 ;
        RECT 251.400 514.050 252.450 538.950 ;
        RECT 256.950 535.950 259.050 538.050 ;
        RECT 257.400 528.600 258.450 535.950 ;
        RECT 263.400 528.600 264.450 547.950 ;
        RECT 266.400 532.050 267.450 583.950 ;
        RECT 269.400 574.050 270.450 589.950 ;
        RECT 272.400 580.050 273.450 599.400 ;
        RECT 278.400 592.050 279.450 599.400 ;
        RECT 289.950 598.650 292.050 600.750 ;
        RECT 296.400 599.400 297.600 601.500 ;
        RECT 296.400 592.050 297.450 599.400 ;
        RECT 277.950 589.950 280.050 592.050 ;
        RECT 295.950 589.950 298.050 592.050 ;
        RECT 274.950 583.950 277.050 586.050 ;
        RECT 271.950 577.950 274.050 580.050 ;
        RECT 275.400 576.450 276.450 583.950 ;
        RECT 280.950 577.950 283.050 580.050 ;
        RECT 272.400 575.400 276.450 576.450 ;
        RECT 268.950 571.950 271.050 574.050 ;
        RECT 272.400 573.600 273.450 575.400 ;
        RECT 272.400 571.500 273.600 573.600 ;
        RECT 271.950 569.100 274.050 571.200 ;
        RECT 274.950 569.100 277.050 571.200 ;
        RECT 275.400 568.050 276.600 568.800 ;
        RECT 268.950 565.950 271.050 568.050 ;
        RECT 274.950 565.950 277.050 568.050 ;
        RECT 269.400 553.050 270.450 565.950 ;
        RECT 268.950 550.950 271.050 553.050 ;
        RECT 268.950 544.950 271.050 547.050 ;
        RECT 265.950 529.950 268.050 532.050 ;
        RECT 269.400 529.050 270.450 544.950 ;
        RECT 281.400 535.050 282.450 577.950 ;
        RECT 302.400 574.050 303.450 613.950 ;
        RECT 305.400 600.750 306.450 625.950 ;
        RECT 308.400 622.050 309.450 631.950 ;
        RECT 307.950 619.950 310.050 622.050 ;
        RECT 311.400 607.050 312.450 637.950 ;
        RECT 314.400 609.450 315.450 643.800 ;
        RECT 316.950 634.950 319.050 637.050 ;
        RECT 317.400 625.050 318.450 634.950 ;
        RECT 320.400 631.050 321.450 644.400 ;
        RECT 325.950 643.950 328.050 646.050 ;
        RECT 319.950 628.950 322.050 631.050 ;
        RECT 316.950 622.950 319.050 625.050 ;
        RECT 322.950 616.950 325.050 619.050 ;
        RECT 323.400 610.050 324.450 616.950 ;
        RECT 314.400 608.400 318.450 609.450 ;
        RECT 307.950 606.600 312.450 607.050 ;
        RECT 317.400 606.600 318.450 608.400 ;
        RECT 322.950 607.950 325.050 610.050 ;
        RECT 307.950 604.950 312.600 606.600 ;
        RECT 311.400 604.350 312.600 604.950 ;
        RECT 317.400 604.350 318.600 606.600 ;
        RECT 310.950 601.950 313.050 604.050 ;
        RECT 313.950 601.950 316.050 604.050 ;
        RECT 316.950 601.950 319.050 604.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 304.950 598.650 307.050 600.750 ;
        RECT 307.950 598.950 310.050 601.050 ;
        RECT 314.400 600.900 315.600 601.650 ;
        RECT 308.400 589.050 309.450 598.950 ;
        RECT 313.950 598.800 316.050 600.900 ;
        RECT 320.400 599.400 321.600 601.650 ;
        RECT 320.400 597.450 321.450 599.400 ;
        RECT 322.950 598.950 325.050 601.050 ;
        RECT 317.400 596.400 321.450 597.450 ;
        RECT 307.950 586.950 310.050 589.050 ;
        RECT 317.400 574.050 318.450 596.400 ;
        RECT 319.950 592.950 322.050 595.050 ;
        RECT 320.400 586.050 321.450 592.950 ;
        RECT 319.950 583.950 322.050 586.050 ;
        RECT 319.950 577.950 322.050 580.050 ;
        RECT 301.950 571.950 304.050 574.050 ;
        RECT 316.950 571.950 319.050 574.050 ;
        RECT 286.950 569.100 289.050 571.200 ;
        RECT 289.950 569.100 292.050 571.200 ;
        RECT 295.950 569.100 298.050 571.200 ;
        RECT 304.950 569.100 307.050 571.200 ;
        RECT 310.950 569.100 313.050 571.200 ;
        RECT 313.950 569.100 316.050 571.200 ;
        RECT 287.400 567.000 288.600 568.800 ;
        RECT 286.950 562.950 289.050 567.000 ;
        RECT 296.400 566.400 297.600 568.800 ;
        RECT 305.400 568.050 306.600 568.800 ;
        RECT 286.950 550.950 289.050 553.050 ;
        RECT 271.950 532.950 274.050 535.050 ;
        RECT 280.950 532.950 283.050 535.050 ;
        RECT 257.400 526.350 258.600 528.600 ;
        RECT 263.400 526.350 264.600 528.600 ;
        RECT 268.950 526.950 271.050 529.050 ;
        RECT 256.950 523.950 259.050 526.050 ;
        RECT 259.950 523.950 262.050 526.050 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 265.950 523.950 268.050 526.050 ;
        RECT 260.400 522.900 261.600 523.650 ;
        RECT 266.400 522.900 267.600 523.650 ;
        RECT 259.950 520.800 262.050 522.900 ;
        RECT 265.950 520.800 268.050 522.900 ;
        RECT 268.950 520.950 271.050 523.050 ;
        RECT 250.950 511.950 253.050 514.050 ;
        RECT 239.400 493.350 240.600 495.600 ;
        RECT 244.950 494.100 247.050 496.200 ;
        RECT 251.400 495.450 252.450 511.950 ;
        RECT 269.400 511.050 270.450 520.950 ;
        RECT 268.950 508.950 271.050 511.050 ;
        RECT 259.950 505.950 262.050 508.050 ;
        RECT 256.950 502.950 259.050 505.050 ;
        RECT 257.400 496.050 258.450 502.950 ;
        RECT 260.400 499.050 261.450 505.950 ;
        RECT 272.400 505.050 273.450 532.950 ;
        RECT 287.400 531.450 288.450 550.950 ;
        RECT 296.400 550.050 297.450 566.400 ;
        RECT 304.950 565.950 307.050 568.050 ;
        RECT 314.400 566.400 315.600 568.800 ;
        RECT 307.950 559.950 310.050 562.050 ;
        RECT 295.950 547.950 298.050 550.050 ;
        RECT 298.950 544.950 301.050 547.050 ;
        RECT 295.950 541.950 298.050 544.050 ;
        RECT 284.400 530.400 288.450 531.450 ;
        RECT 274.950 528.600 279.000 529.050 ;
        RECT 284.400 528.600 285.450 530.400 ;
        RECT 296.400 529.050 297.450 541.950 ;
        RECT 299.400 529.050 300.450 544.950 ;
        RECT 292.950 528.600 297.450 529.050 ;
        RECT 274.950 526.950 279.600 528.600 ;
        RECT 278.400 526.350 279.600 526.950 ;
        RECT 284.400 526.350 285.600 528.600 ;
        RECT 292.950 526.950 297.600 528.600 ;
        RECT 298.950 526.950 301.050 529.050 ;
        RECT 296.400 526.200 297.600 526.950 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 286.950 523.950 289.050 526.050 ;
        RECT 295.950 523.800 298.050 525.900 ;
        RECT 298.950 523.800 301.050 525.900 ;
        RECT 301.950 523.800 304.050 525.900 ;
        RECT 281.400 521.400 282.600 523.650 ;
        RECT 287.400 521.400 288.600 523.650 ;
        RECT 281.400 517.050 282.450 521.400 ;
        RECT 280.950 514.950 283.050 517.050 ;
        RECT 287.400 514.050 288.450 521.400 ;
        RECT 289.800 520.950 291.900 523.050 ;
        RECT 292.950 520.950 295.050 523.050 ;
        RECT 299.400 522.750 300.600 523.500 ;
        RECT 290.400 517.050 291.450 520.950 ;
        RECT 289.950 514.950 292.050 517.050 ;
        RECT 283.800 511.950 285.900 514.050 ;
        RECT 286.950 511.950 289.050 514.050 ;
        RECT 274.950 505.950 277.050 508.050 ;
        RECT 271.950 502.950 274.050 505.050 ;
        RECT 262.950 499.950 265.050 502.050 ;
        RECT 268.950 501.900 273.000 502.050 ;
        RECT 268.950 499.950 274.050 501.900 ;
        RECT 259.950 496.950 262.050 499.050 ;
        RECT 251.400 494.400 255.450 495.450 ;
        RECT 245.400 493.350 246.600 494.100 ;
        RECT 229.950 491.100 232.050 493.200 ;
        RECT 230.400 489.000 231.600 491.100 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 241.950 490.950 244.050 493.050 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 247.950 490.950 250.050 493.050 ;
        RECT 229.950 484.950 232.050 489.000 ;
        RECT 232.950 487.800 235.050 489.900 ;
        RECT 242.400 489.000 243.600 490.650 ;
        RECT 217.800 482.400 219.900 484.500 ;
        RECT 226.800 482.700 228.900 484.800 ;
        RECT 214.950 478.950 217.050 481.050 ;
        RECT 211.950 451.950 214.050 454.050 ;
        RECT 197.400 448.200 198.600 448.950 ;
        RECT 206.400 448.200 207.600 450.600 ;
        RECT 208.950 448.950 211.050 451.050 ;
        RECT 181.950 445.800 184.050 447.900 ;
        RECT 184.950 445.800 187.050 447.900 ;
        RECT 187.950 445.800 190.050 447.900 ;
        RECT 196.950 445.800 199.050 447.900 ;
        RECT 202.950 445.800 205.050 447.900 ;
        RECT 205.950 445.800 208.050 447.900 ;
        RECT 175.950 442.650 178.050 444.750 ;
        RECT 185.400 443.400 186.600 445.500 ;
        RECT 203.400 444.750 204.600 445.500 ;
        RECT 212.400 445.050 213.450 451.950 ;
        RECT 215.400 451.050 216.450 478.950 ;
        RECT 220.950 457.950 223.050 460.050 ;
        RECT 214.950 448.950 217.050 451.050 ;
        RECT 221.400 450.600 222.450 457.950 ;
        RECT 181.950 430.950 184.050 433.050 ;
        RECT 175.950 424.950 178.050 427.050 ;
        RECT 170.400 416.400 174.450 417.450 ;
        RECT 164.400 415.350 165.600 416.100 ;
        RECT 170.400 415.350 171.600 416.400 ;
        RECT 163.950 412.950 166.050 415.050 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 169.950 412.950 172.050 415.050 ;
        RECT 160.950 409.950 163.050 412.050 ;
        RECT 167.400 410.400 168.600 412.650 ;
        RECT 145.950 397.950 148.050 400.050 ;
        RECT 157.950 397.950 160.050 400.050 ;
        RECT 142.950 391.950 145.050 394.050 ;
        RECT 136.950 373.950 139.050 376.050 ;
        RECT 133.950 371.100 136.050 373.200 ;
        RECT 143.400 373.050 144.450 391.950 ;
        RECT 146.400 388.050 147.450 397.950 ;
        RECT 161.400 394.050 162.450 409.950 ;
        RECT 163.950 406.950 166.050 409.050 ;
        RECT 160.950 391.950 163.050 394.050 ;
        RECT 145.950 385.950 148.050 388.050 ;
        RECT 151.800 376.500 153.900 378.600 ;
        RECT 134.400 370.350 135.600 371.100 ;
        RECT 142.950 370.950 145.050 373.050 ;
        RECT 130.950 367.950 133.050 370.050 ;
        RECT 133.950 367.950 136.050 370.050 ;
        RECT 136.950 367.950 139.050 370.050 ;
        RECT 131.400 366.000 132.600 367.650 ;
        RECT 137.400 366.900 138.600 367.650 ;
        RECT 130.950 361.950 133.050 366.000 ;
        RECT 136.950 364.800 139.050 366.900 ;
        RECT 143.400 364.050 144.450 370.950 ;
        RECT 151.950 369.900 152.850 376.500 ;
        RECT 160.800 376.200 162.900 378.300 ;
        RECT 155.400 372.900 156.600 375.600 ;
        RECT 154.650 370.800 156.750 372.900 ;
        RECT 158.700 369.900 160.800 370.200 ;
        RECT 148.950 367.800 151.050 369.900 ;
        RECT 151.950 369.000 160.800 369.900 ;
        RECT 149.400 365.400 150.600 367.800 ;
        RECT 142.950 361.950 145.050 364.050 ;
        RECT 151.950 363.900 152.850 369.000 ;
        RECT 158.700 368.100 160.800 369.000 ;
        RECT 153.750 367.200 155.850 368.100 ;
        RECT 153.750 366.000 160.800 367.200 ;
        RECT 157.950 365.100 160.800 366.000 ;
        RECT 157.950 364.800 160.050 365.100 ;
        RECT 151.200 361.800 153.300 363.900 ;
        RECT 154.650 362.100 156.750 364.200 ;
        RECT 161.700 363.600 162.600 376.200 ;
        RECT 164.400 372.600 165.450 406.950 ;
        RECT 167.400 406.050 168.450 410.400 ;
        RECT 166.950 403.950 169.050 406.050 ;
        RECT 169.950 388.950 172.050 391.050 ;
        RECT 170.400 381.450 171.450 388.950 ;
        RECT 176.400 388.050 177.450 424.950 ;
        RECT 182.400 417.450 183.450 430.950 ;
        RECT 185.400 424.050 186.450 443.400 ;
        RECT 202.950 442.650 205.050 444.750 ;
        RECT 211.950 442.950 214.050 445.050 ;
        RECT 184.950 421.950 187.050 424.050 ;
        RECT 203.400 418.350 204.450 442.650 ;
        RECT 205.950 439.950 208.050 442.050 ;
        RECT 206.400 421.050 207.450 439.950 ;
        RECT 208.950 433.950 211.050 436.050 ;
        RECT 205.950 418.950 208.050 421.050 ;
        RECT 179.400 416.400 183.450 417.450 ;
        RECT 175.950 385.950 178.050 388.050 ;
        RECT 167.400 380.400 171.450 381.450 ;
        RECT 167.400 376.050 168.450 380.400 ;
        RECT 179.400 379.050 180.450 416.400 ;
        RECT 187.950 416.250 190.050 418.350 ;
        RECT 202.950 416.250 205.050 418.350 ;
        RECT 209.400 417.600 210.450 433.950 ;
        RECT 215.400 430.050 216.450 448.950 ;
        RECT 221.400 448.200 222.600 450.600 ;
        RECT 226.950 448.950 229.050 451.050 ;
        RECT 227.400 448.200 228.600 448.950 ;
        RECT 220.950 445.800 223.050 447.900 ;
        RECT 223.950 445.800 226.050 447.900 ;
        RECT 226.950 445.800 229.050 447.900 ;
        RECT 224.400 443.400 225.600 445.500 ;
        RECT 214.950 427.950 217.050 430.050 ;
        RECT 224.400 421.050 225.450 443.400 ;
        RECT 233.400 439.050 234.450 487.800 ;
        RECT 241.950 484.950 244.050 489.000 ;
        RECT 248.400 488.400 249.600 490.650 ;
        RECT 254.400 490.050 255.450 494.400 ;
        RECT 256.950 493.950 259.050 496.050 ;
        RECT 263.400 495.600 264.450 499.950 ;
        RECT 271.950 499.800 274.050 499.950 ;
        RECT 275.400 499.050 276.450 505.950 ;
        RECT 284.400 505.050 285.450 511.950 ;
        RECT 283.950 502.950 286.050 505.050 ;
        RECT 280.950 501.900 285.000 502.050 ;
        RECT 280.950 499.950 286.050 501.900 ;
        RECT 289.950 499.950 292.050 502.050 ;
        RECT 283.950 499.800 286.050 499.950 ;
        RECT 274.950 496.950 277.050 499.050 ;
        RECT 277.950 496.950 280.050 499.050 ;
        RECT 263.400 493.500 264.600 495.600 ;
        RECT 268.950 494.250 271.050 496.350 ;
        RECT 269.400 493.500 270.600 494.250 ;
        RECT 274.950 493.800 277.050 495.900 ;
        RECT 259.950 491.100 262.050 493.200 ;
        RECT 262.950 491.100 265.050 493.200 ;
        RECT 265.950 491.100 268.050 493.200 ;
        RECT 268.950 491.100 271.050 493.200 ;
        RECT 260.400 490.050 261.600 490.800 ;
        RECT 248.400 478.050 249.450 488.400 ;
        RECT 250.800 487.950 252.900 490.050 ;
        RECT 253.950 487.950 256.050 490.050 ;
        RECT 259.950 487.950 262.050 490.050 ;
        RECT 266.400 489.000 267.600 490.800 ;
        RECT 247.950 475.950 250.050 478.050 ;
        RECT 251.400 451.050 252.450 487.950 ;
        RECT 265.950 484.950 268.050 489.000 ;
        RECT 268.950 484.950 271.050 487.050 ;
        RECT 269.400 472.050 270.450 484.950 ;
        RECT 275.400 478.050 276.450 493.800 ;
        RECT 274.950 475.950 277.050 478.050 ;
        RECT 275.400 472.050 276.450 475.950 ;
        RECT 268.950 469.950 271.050 472.050 ;
        RECT 274.950 469.950 277.050 472.050 ;
        RECT 259.800 453.300 261.900 455.400 ;
        RECT 269.400 454.500 271.500 456.600 ;
        RECT 235.950 450.600 240.000 451.050 ;
        RECT 235.950 448.950 240.600 450.600 ;
        RECT 247.950 448.950 250.050 451.050 ;
        RECT 250.950 448.950 253.050 451.050 ;
        RECT 256.950 448.950 259.050 451.050 ;
        RECT 239.400 448.200 240.600 448.950 ;
        RECT 248.400 448.200 249.600 448.950 ;
        RECT 257.400 447.900 258.600 448.950 ;
        RECT 238.950 445.800 241.050 447.900 ;
        RECT 241.950 445.800 244.050 447.900 ;
        RECT 247.950 445.800 250.050 447.900 ;
        RECT 256.950 445.800 259.050 447.900 ;
        RECT 242.400 443.400 243.600 445.500 ;
        RECT 260.700 444.300 261.600 453.300 ;
        RECT 262.950 449.700 265.050 451.800 ;
        RECT 266.400 450.900 267.600 453.600 ;
        RECT 264.150 447.300 265.050 449.700 ;
        RECT 265.950 448.800 268.050 450.900 ;
        RECT 269.850 447.300 271.050 454.500 ;
        RECT 275.400 451.050 276.450 469.950 ;
        RECT 274.950 448.950 277.050 451.050 ;
        RECT 274.050 447.900 276.450 448.050 ;
        RECT 264.150 446.100 271.050 447.300 ;
        RECT 267.150 444.300 269.250 445.200 ;
        RECT 242.400 439.050 243.450 443.400 ;
        RECT 260.700 443.100 269.250 444.300 ;
        RECT 262.200 441.300 264.300 443.100 ;
        RECT 265.950 440.100 268.050 442.200 ;
        RECT 270.150 440.700 271.050 446.100 ;
        RECT 271.950 445.950 277.050 447.900 ;
        RECT 271.950 445.800 274.050 445.950 ;
        RECT 274.950 445.800 277.050 445.950 ;
        RECT 272.400 443.400 273.600 445.800 ;
        RECT 278.400 445.050 279.450 496.950 ;
        RECT 283.950 494.100 286.050 498.900 ;
        RECT 290.400 496.200 291.450 499.950 ;
        RECT 293.400 499.050 294.450 520.950 ;
        RECT 298.950 520.650 301.050 522.750 ;
        RECT 308.400 522.450 309.450 559.950 ;
        RECT 314.400 556.050 315.450 566.400 ;
        RECT 313.950 553.950 316.050 556.050 ;
        RECT 320.400 547.050 321.450 577.950 ;
        RECT 323.400 577.050 324.450 598.950 ;
        RECT 326.400 580.050 327.450 643.950 ;
        RECT 329.400 613.050 330.450 652.950 ;
        RECT 332.400 652.050 333.450 664.950 ;
        RECT 338.400 655.050 339.450 694.950 ;
        RECT 340.950 691.950 343.050 694.050 ;
        RECT 341.400 679.050 342.450 691.950 ;
        RECT 343.950 682.950 346.050 688.050 ;
        RECT 346.950 682.950 349.050 685.050 ;
        RECT 352.950 684.000 355.050 688.050 ;
        RECT 356.400 685.050 357.450 712.950 ;
        RECT 359.400 700.050 360.450 712.950 ;
        RECT 362.400 706.050 363.450 718.950 ;
        RECT 368.400 709.050 369.450 722.400 ;
        RECT 376.950 721.800 379.050 723.900 ;
        RECT 383.400 722.400 384.600 724.650 ;
        RECT 373.950 715.950 376.050 718.050 ;
        RECT 376.950 717.450 381.000 718.050 ;
        RECT 376.950 715.950 381.450 717.450 ;
        RECT 370.950 712.950 373.050 715.050 ;
        RECT 367.950 706.950 370.050 709.050 ;
        RECT 361.950 703.950 364.050 706.050 ;
        RECT 371.400 703.050 372.450 712.950 ;
        RECT 364.950 700.950 367.050 703.050 ;
        RECT 370.950 700.950 373.050 703.050 ;
        RECT 358.950 697.950 361.050 700.050 ;
        RECT 361.950 688.950 364.050 691.050 ;
        RECT 347.400 682.200 348.600 682.950 ;
        RECT 353.400 682.200 354.600 684.000 ;
        RECT 355.950 682.950 358.050 685.050 ;
        RECT 362.400 684.600 363.450 688.950 ;
        RECT 365.400 688.050 366.450 700.950 ;
        RECT 367.950 688.950 370.050 691.050 ;
        RECT 364.950 685.950 367.050 688.050 ;
        RECT 368.400 684.600 369.450 688.950 ;
        RECT 374.400 685.050 375.450 715.950 ;
        RECT 376.950 709.950 379.050 712.050 ;
        RECT 377.400 700.050 378.450 709.950 ;
        RECT 380.400 706.050 381.450 715.950 ;
        RECT 383.400 715.050 384.450 722.400 ;
        RECT 388.950 721.950 391.050 724.050 ;
        RECT 398.400 722.400 399.600 724.650 ;
        RECT 404.400 722.400 405.600 724.650 ;
        RECT 382.950 712.950 385.050 715.050 ;
        RECT 379.950 703.950 382.050 706.050 ;
        RECT 376.950 697.950 379.050 700.050 ;
        RECT 376.950 688.950 379.050 691.050 ;
        RECT 362.400 682.200 363.600 684.600 ;
        RECT 368.400 682.200 369.600 684.600 ;
        RECT 373.950 682.950 376.050 685.050 ;
        RECT 346.950 679.800 349.050 681.900 ;
        RECT 349.950 679.800 352.050 681.900 ;
        RECT 352.950 679.800 355.050 681.900 ;
        RECT 361.950 679.800 364.050 681.900 ;
        RECT 364.950 679.800 367.050 681.900 ;
        RECT 367.950 679.800 370.050 681.900 ;
        RECT 370.950 679.800 373.050 681.900 ;
        RECT 340.950 676.950 343.050 679.050 ;
        RECT 343.950 676.950 346.050 679.050 ;
        RECT 350.400 678.750 351.600 679.500 ;
        RECT 337.800 652.950 339.900 655.050 ;
        RECT 331.950 649.950 334.050 652.050 ;
        RECT 338.400 651.450 339.600 651.600 ;
        RECT 340.950 651.450 343.050 655.050 ;
        RECT 344.400 652.350 345.450 676.950 ;
        RECT 349.950 676.650 352.050 678.750 ;
        RECT 365.400 678.000 366.600 679.500 ;
        RECT 364.950 673.950 367.050 678.000 ;
        RECT 371.400 677.400 372.600 679.500 ;
        RECT 371.400 670.050 372.450 677.400 ;
        RECT 370.950 667.950 373.050 670.050 ;
        RECT 377.400 664.050 378.450 688.950 ;
        RECT 389.400 688.050 390.450 721.950 ;
        RECT 398.400 715.050 399.450 722.400 ;
        RECT 404.400 718.050 405.450 722.400 ;
        RECT 403.950 715.950 406.050 718.050 ;
        RECT 397.950 712.950 400.050 715.050 ;
        RECT 400.950 709.950 403.050 712.050 ;
        RECT 397.950 706.950 400.050 709.050 ;
        RECT 394.950 691.950 397.050 694.050 ;
        RECT 379.950 685.950 382.050 688.050 ;
        RECT 388.950 685.950 391.050 688.050 ;
        RECT 380.400 678.450 381.450 685.950 ;
        RECT 389.400 684.600 390.450 685.950 ;
        RECT 395.400 684.600 396.450 691.950 ;
        RECT 398.400 685.050 399.450 706.950 ;
        RECT 401.400 706.050 402.450 709.950 ;
        RECT 410.400 706.050 411.450 730.950 ;
        RECT 412.950 727.950 415.050 730.050 ;
        RECT 418.950 728.250 421.050 730.350 ;
        RECT 425.400 729.600 426.450 748.950 ;
        RECT 431.400 742.050 432.450 755.400 ;
        RECT 437.400 748.050 438.450 755.400 ;
        RECT 451.950 751.950 454.050 756.000 ;
        RECT 457.950 754.650 460.050 756.750 ;
        RECT 459.000 753.450 463.050 754.050 ;
        RECT 458.400 753.000 463.050 753.450 ;
        RECT 457.950 751.950 463.050 753.000 ;
        RECT 457.950 751.050 460.050 751.950 ;
        RECT 439.950 748.950 442.050 751.050 ;
        RECT 457.800 750.000 460.050 751.050 ;
        RECT 457.800 748.950 459.900 750.000 ;
        RECT 436.950 745.950 439.050 748.050 ;
        RECT 430.950 739.950 433.050 742.050 ;
        RECT 431.400 730.050 432.450 739.950 ;
        RECT 400.950 703.950 403.050 706.050 ;
        RECT 409.950 703.950 412.050 706.050 ;
        RECT 409.950 691.950 412.050 694.050 ;
        RECT 389.400 682.200 390.600 684.600 ;
        RECT 395.400 682.200 396.600 684.600 ;
        RECT 397.950 682.950 400.050 685.050 ;
        RECT 403.950 684.000 406.050 688.050 ;
        RECT 410.400 685.050 411.450 691.950 ;
        RECT 413.400 688.050 414.450 727.950 ;
        RECT 419.400 727.500 420.600 728.250 ;
        RECT 425.400 727.500 426.600 729.600 ;
        RECT 430.950 727.950 433.050 730.050 ;
        RECT 440.400 729.600 441.450 748.950 ;
        RECT 460.950 748.800 463.050 750.900 ;
        RECT 448.950 745.950 451.050 748.050 ;
        RECT 445.950 733.950 448.050 736.050 ;
        RECT 446.400 729.600 447.450 733.950 ;
        RECT 449.400 732.450 450.450 745.950 ;
        RECT 457.950 742.950 460.050 745.050 ;
        RECT 449.400 731.400 453.450 732.450 ;
        RECT 440.400 727.500 441.600 729.600 ;
        RECT 446.400 727.500 447.600 729.600 ;
        RECT 418.950 725.100 421.050 727.200 ;
        RECT 421.950 725.100 424.050 727.200 ;
        RECT 424.950 725.100 427.050 727.200 ;
        RECT 427.950 725.100 430.050 727.200 ;
        RECT 436.950 725.100 439.050 727.200 ;
        RECT 439.950 725.100 442.050 727.200 ;
        RECT 442.950 725.100 445.050 727.200 ;
        RECT 445.950 725.100 448.050 727.200 ;
        RECT 422.400 724.050 423.600 724.800 ;
        RECT 415.950 721.950 418.050 724.050 ;
        RECT 421.950 721.950 424.050 724.050 ;
        RECT 428.400 722.400 429.600 724.800 ;
        RECT 437.400 723.000 438.600 724.800 ;
        RECT 412.950 685.950 415.050 688.050 ;
        RECT 416.400 685.050 417.450 721.950 ;
        RECT 428.400 718.050 429.450 722.400 ;
        RECT 436.950 718.950 439.050 723.000 ;
        RECT 443.400 722.400 444.600 724.800 ;
        RECT 443.400 718.050 444.450 722.400 ;
        RECT 427.950 715.950 430.050 718.050 ;
        RECT 442.950 715.950 445.050 718.050 ;
        RECT 452.400 714.450 453.450 731.400 ;
        RECT 454.950 730.950 457.050 733.050 ;
        RECT 455.400 715.050 456.450 730.950 ;
        RECT 458.400 730.050 459.450 742.950 ;
        RECT 461.400 733.050 462.450 748.800 ;
        RECT 467.400 745.050 468.450 763.950 ;
        RECT 476.400 762.600 477.450 763.950 ;
        RECT 482.400 763.050 483.450 766.800 ;
        RECT 476.400 760.200 477.600 762.600 ;
        RECT 481.950 760.950 484.050 763.050 ;
        RECT 482.400 760.200 483.600 760.950 ;
        RECT 472.950 757.800 475.050 759.900 ;
        RECT 475.950 757.800 478.050 759.900 ;
        RECT 478.950 757.800 481.050 759.900 ;
        RECT 481.950 757.800 484.050 759.900 ;
        RECT 473.400 755.400 474.600 757.500 ;
        RECT 479.400 755.400 480.600 757.500 ;
        RECT 466.950 742.950 469.050 745.050 ;
        RECT 473.400 742.050 474.450 755.400 ;
        RECT 479.400 745.050 480.450 755.400 ;
        RECT 484.950 754.950 487.050 757.050 ;
        RECT 485.400 745.050 486.450 754.950 ;
        RECT 478.950 742.950 481.050 745.050 ;
        RECT 484.950 742.950 487.050 745.050 ;
        RECT 472.950 739.950 475.050 742.050 ;
        RECT 475.950 733.950 478.050 736.050 ;
        RECT 460.950 730.950 463.050 733.050 ;
        RECT 457.950 727.950 460.050 730.050 ;
        RECT 463.950 728.250 466.050 730.350 ;
        RECT 464.400 727.500 465.600 728.250 ;
        RECT 460.950 725.100 463.050 727.200 ;
        RECT 463.950 725.100 466.050 727.200 ;
        RECT 469.950 725.100 472.050 727.200 ;
        RECT 461.400 724.050 462.600 724.800 ;
        RECT 470.400 724.050 471.600 724.800 ;
        RECT 460.950 721.950 463.050 724.050 ;
        RECT 469.950 721.950 472.050 724.050 ;
        RECT 457.950 718.950 460.050 721.050 ;
        RECT 449.400 713.400 453.450 714.450 ;
        RECT 433.950 703.950 436.050 706.050 ;
        RECT 418.950 691.950 421.050 694.050 ;
        RECT 419.400 688.050 420.450 691.950 ;
        RECT 430.950 688.950 433.050 691.050 ;
        RECT 418.950 685.950 421.050 688.050 ;
        RECT 404.400 682.200 405.600 684.000 ;
        RECT 409.950 682.950 412.050 685.050 ;
        RECT 415.950 682.950 418.050 685.050 ;
        RECT 410.400 682.200 411.600 682.950 ;
        RECT 385.950 679.800 388.050 681.900 ;
        RECT 388.950 679.800 391.050 681.900 ;
        RECT 391.950 679.800 394.050 681.900 ;
        RECT 394.950 679.800 397.050 681.900 ;
        RECT 403.950 679.800 406.050 681.900 ;
        RECT 406.950 679.800 409.050 681.900 ;
        RECT 409.950 679.800 412.050 681.900 ;
        RECT 412.950 679.800 415.050 681.900 ;
        RECT 380.400 677.400 384.450 678.450 ;
        RECT 386.400 678.000 387.600 679.500 ;
        RECT 379.950 667.950 382.050 670.050 ;
        RECT 355.950 658.950 358.050 661.050 ;
        RECT 364.950 660.450 367.050 664.050 ;
        RECT 370.950 661.950 373.050 664.050 ;
        RECT 376.950 661.950 379.050 664.050 ;
        RECT 362.400 660.000 367.050 660.450 ;
        RECT 362.400 659.400 366.450 660.000 ;
        RECT 338.400 651.000 343.050 651.450 ;
        RECT 338.400 650.400 342.450 651.000 ;
        RECT 338.400 649.350 339.600 650.400 ;
        RECT 343.950 650.250 346.050 652.350 ;
        RECT 349.950 650.250 352.050 652.350 ;
        RECT 356.400 652.050 357.450 658.950 ;
        RECT 362.400 657.450 363.450 659.400 ;
        RECT 359.400 656.400 363.450 657.450 ;
        RECT 350.400 649.500 351.600 650.250 ;
        RECT 355.950 649.950 358.050 652.050 ;
        RECT 334.950 646.950 337.050 649.050 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 346.950 647.100 349.050 649.200 ;
        RECT 349.950 647.100 352.050 649.200 ;
        RECT 352.950 647.100 355.050 649.200 ;
        RECT 335.400 646.050 336.600 646.650 ;
        RECT 331.950 644.400 336.600 646.050 ;
        RECT 347.400 645.900 348.600 646.800 ;
        RECT 331.950 643.950 336.000 644.400 ;
        RECT 346.950 643.800 349.050 645.900 ;
        RECT 353.400 644.400 354.600 646.800 ;
        RECT 331.950 622.950 334.050 625.050 ;
        RECT 328.950 610.950 331.050 613.050 ;
        RECT 332.400 609.450 333.450 622.950 ;
        RECT 347.400 622.050 348.450 643.800 ;
        RECT 349.950 622.950 352.050 625.050 ;
        RECT 346.950 619.950 349.050 622.050 ;
        RECT 350.400 616.050 351.450 622.950 ;
        RECT 353.400 618.450 354.450 644.400 ;
        RECT 355.950 643.950 358.050 646.050 ;
        RECT 356.400 622.050 357.450 643.950 ;
        RECT 355.950 619.950 358.050 622.050 ;
        RECT 353.400 617.400 357.450 618.450 ;
        RECT 349.950 613.950 352.050 616.050 ;
        RECT 356.400 613.050 357.450 617.400 ;
        RECT 359.400 616.050 360.450 656.400 ;
        RECT 364.950 655.950 367.050 658.050 ;
        RECT 361.950 649.950 364.050 655.050 ;
        RECT 365.400 652.200 366.450 655.950 ;
        RECT 364.950 650.100 367.050 652.200 ;
        RECT 371.400 651.600 372.450 661.950 ;
        RECT 365.400 649.350 366.600 650.100 ;
        RECT 371.400 649.350 372.600 651.600 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 367.950 646.950 370.050 649.050 ;
        RECT 370.950 646.950 373.050 649.050 ;
        RECT 373.950 646.950 376.050 649.050 ;
        RECT 368.400 644.400 369.600 646.650 ;
        RECT 374.400 645.900 375.600 646.650 ;
        RECT 368.400 631.050 369.450 644.400 ;
        RECT 373.950 643.800 376.050 645.900 ;
        RECT 380.400 637.050 381.450 667.950 ;
        RECT 370.950 634.950 373.050 637.050 ;
        RECT 379.950 634.950 382.050 637.050 ;
        RECT 367.950 628.950 370.050 631.050 ;
        RECT 358.950 613.950 361.050 616.050 ;
        RECT 346.950 610.950 349.050 613.050 ;
        RECT 355.950 610.950 358.050 613.050 ;
        RECT 329.400 609.000 333.450 609.450 ;
        RECT 328.950 608.400 333.450 609.000 ;
        RECT 328.950 604.950 331.050 608.400 ;
        RECT 334.950 604.950 337.050 607.050 ;
        RECT 340.950 604.950 343.050 607.050 ;
        RECT 335.400 604.200 336.600 604.950 ;
        RECT 341.400 604.200 342.600 604.950 ;
        RECT 331.950 601.800 334.050 603.900 ;
        RECT 334.950 601.800 337.050 603.900 ;
        RECT 337.950 601.800 340.050 603.900 ;
        RECT 340.950 601.800 343.050 603.900 ;
        RECT 332.400 601.050 333.600 601.500 ;
        RECT 328.950 599.400 333.600 601.050 ;
        RECT 338.400 600.000 339.600 601.500 ;
        RECT 328.950 598.950 333.000 599.400 ;
        RECT 331.950 595.950 334.050 598.050 ;
        RECT 337.950 595.950 340.050 600.000 ;
        RECT 325.950 577.950 328.050 580.050 ;
        RECT 323.400 576.900 327.000 577.050 ;
        RECT 323.400 574.950 328.050 576.900 ;
        RECT 323.400 574.050 324.450 574.950 ;
        RECT 325.950 574.800 328.050 574.950 ;
        RECT 322.800 571.950 324.900 574.050 ;
        RECT 325.950 571.950 328.050 574.050 ;
        RECT 332.400 573.600 333.450 595.950 ;
        RECT 347.400 583.050 348.450 610.950 ;
        RECT 352.950 606.000 355.050 610.050 ;
        RECT 368.400 607.200 369.450 628.950 ;
        RECT 353.400 604.350 354.600 606.000 ;
        RECT 358.950 605.100 361.050 607.200 ;
        RECT 367.950 605.100 370.050 607.200 ;
        RECT 371.400 607.050 372.450 634.950 ;
        RECT 383.400 628.050 384.450 677.400 ;
        RECT 385.950 673.950 388.050 678.000 ;
        RECT 392.400 677.400 393.600 679.500 ;
        RECT 407.400 677.400 408.600 679.500 ;
        RECT 413.400 677.400 414.600 679.500 ;
        RECT 392.400 673.050 393.450 677.400 ;
        RECT 407.400 673.050 408.450 677.400 ;
        RECT 391.950 670.950 394.050 673.050 ;
        RECT 406.950 670.950 409.050 673.050 ;
        RECT 397.950 664.950 400.050 667.050 ;
        RECT 388.950 655.950 391.050 658.050 ;
        RECT 389.400 652.350 390.450 655.950 ;
        RECT 388.950 650.250 391.050 652.350 ;
        RECT 389.400 649.500 390.600 650.250 ;
        RECT 388.950 647.100 391.050 649.200 ;
        RECT 391.950 647.100 394.050 649.200 ;
        RECT 388.950 643.950 391.050 646.050 ;
        RECT 392.400 644.400 393.600 646.800 ;
        RECT 385.950 631.950 388.050 634.050 ;
        RECT 382.950 625.950 385.050 628.050 ;
        RECT 379.950 624.450 384.000 625.050 ;
        RECT 379.950 622.950 384.450 624.450 ;
        RECT 376.950 621.450 381.000 622.050 ;
        RECT 376.950 619.950 381.450 621.450 ;
        RECT 376.950 613.950 379.050 616.050 ;
        RECT 359.400 604.350 360.600 605.100 ;
        RECT 352.950 601.950 355.050 604.050 ;
        RECT 355.950 601.950 358.050 604.050 ;
        RECT 358.950 601.950 361.050 604.050 ;
        RECT 361.950 601.950 364.050 604.050 ;
        RECT 356.400 600.000 357.600 601.650 ;
        RECT 355.950 595.950 358.050 600.000 ;
        RECT 362.400 599.400 363.600 601.650 ;
        RECT 368.400 600.450 369.450 605.100 ;
        RECT 370.950 604.950 373.050 607.050 ;
        RECT 377.400 606.600 378.450 613.950 ;
        RECT 377.400 604.200 378.600 606.600 ;
        RECT 380.400 606.450 381.450 619.950 ;
        RECT 383.400 619.050 384.450 622.950 ;
        RECT 382.950 616.950 385.050 619.050 ;
        RECT 386.400 613.050 387.450 631.950 ;
        RECT 389.400 621.450 390.450 643.950 ;
        RECT 392.400 625.050 393.450 644.400 ;
        RECT 394.950 643.950 397.050 646.050 ;
        RECT 391.950 622.950 394.050 625.050 ;
        RECT 389.400 620.400 393.450 621.450 ;
        RECT 392.400 616.050 393.450 620.400 ;
        RECT 391.950 613.950 394.050 616.050 ;
        RECT 385.950 610.950 388.050 613.050 ;
        RECT 386.400 607.050 387.450 610.950 ;
        RECT 395.400 610.050 396.450 643.950 ;
        RECT 398.400 622.050 399.450 664.950 ;
        RECT 406.950 650.100 409.050 652.200 ;
        RECT 413.400 651.600 414.450 677.400 ;
        RECT 415.950 676.950 418.050 679.050 ;
        RECT 416.400 667.050 417.450 676.950 ;
        RECT 419.400 673.050 420.450 685.950 ;
        RECT 421.950 682.950 424.050 685.050 ;
        RECT 431.400 684.600 432.450 688.950 ;
        RECT 434.400 685.050 435.450 703.950 ;
        RECT 445.950 688.950 448.050 691.050 ;
        RECT 418.950 670.950 421.050 673.050 ;
        RECT 422.400 670.050 423.450 682.950 ;
        RECT 431.400 682.200 432.600 684.600 ;
        RECT 433.950 682.950 436.050 685.050 ;
        RECT 436.950 684.000 439.050 688.050 ;
        RECT 446.400 684.600 447.450 688.950 ;
        RECT 449.400 688.050 450.450 713.400 ;
        RECT 454.950 712.950 457.050 715.050 ;
        RECT 451.950 709.950 454.050 712.050 ;
        RECT 452.400 696.450 453.450 709.950 ;
        RECT 458.400 697.050 459.450 718.950 ;
        RECT 460.950 706.950 463.050 709.050 ;
        RECT 461.400 700.050 462.450 706.950 ;
        RECT 463.950 700.950 466.050 703.050 ;
        RECT 460.950 697.950 463.050 700.050 ;
        RECT 452.400 695.400 456.450 696.450 ;
        RECT 455.400 688.050 456.450 695.400 ;
        RECT 457.950 694.950 460.050 697.050 ;
        RECT 448.950 685.950 451.050 688.050 ;
        RECT 454.950 685.950 457.050 688.050 ;
        RECT 437.400 682.200 438.600 684.000 ;
        RECT 446.400 682.200 447.600 684.600 ;
        RECT 449.400 684.450 450.450 685.950 ;
        RECT 452.400 684.450 453.600 684.600 ;
        RECT 449.400 683.400 453.600 684.450 ;
        RECT 452.400 682.200 453.600 683.400 ;
        RECT 427.950 679.800 430.050 681.900 ;
        RECT 430.950 679.800 433.050 681.900 ;
        RECT 433.950 679.800 436.050 681.900 ;
        RECT 436.950 679.800 439.050 681.900 ;
        RECT 445.950 679.800 448.050 681.900 ;
        RECT 448.950 679.800 451.050 681.900 ;
        RECT 451.950 679.800 454.050 681.900 ;
        RECT 454.950 679.800 457.050 681.900 ;
        RECT 424.950 676.950 427.050 679.050 ;
        RECT 428.400 677.400 429.600 679.500 ;
        RECT 434.400 678.750 435.600 679.500 ;
        RECT 449.400 678.750 450.600 679.500 ;
        RECT 421.950 667.950 424.050 670.050 ;
        RECT 415.950 664.950 418.050 667.050 ;
        RECT 425.400 658.050 426.450 676.950 ;
        RECT 424.950 655.950 427.050 658.050 ;
        RECT 425.400 651.600 426.450 655.950 ;
        RECT 428.400 652.050 429.450 677.400 ;
        RECT 433.950 676.650 436.050 678.750 ;
        RECT 448.950 676.650 451.050 678.750 ;
        RECT 455.400 677.400 456.600 679.500 ;
        RECT 461.400 679.050 462.450 697.950 ;
        RECT 464.400 697.050 465.450 700.950 ;
        RECT 466.950 697.950 469.050 700.050 ;
        RECT 470.400 699.450 471.450 721.950 ;
        RECT 470.400 698.400 474.450 699.450 ;
        RECT 463.950 694.950 466.050 697.050 ;
        RECT 467.400 688.050 468.450 697.950 ;
        RECT 469.950 688.950 472.050 691.050 ;
        RECT 466.950 685.950 469.050 688.050 ;
        RECT 470.400 685.200 471.450 688.950 ;
        RECT 469.950 683.100 472.050 685.200 ;
        RECT 473.400 685.050 474.450 698.400 ;
        RECT 476.400 685.050 477.450 733.950 ;
        RECT 485.400 729.600 486.450 742.950 ;
        RECT 488.400 736.050 489.450 769.950 ;
        RECT 496.950 760.950 499.050 763.050 ;
        RECT 502.950 762.000 505.050 766.050 ;
        RECT 506.400 762.450 507.450 775.950 ;
        RECT 518.400 768.450 519.450 799.950 ;
        RECT 523.950 787.950 526.050 790.050 ;
        RECT 524.400 784.050 525.450 787.950 ;
        RECT 530.400 787.050 531.450 800.400 ;
        RECT 535.950 796.950 538.050 801.000 ;
        RECT 541.950 799.950 544.050 802.050 ;
        RECT 529.950 784.950 532.050 787.050 ;
        RECT 523.950 781.950 526.050 784.050 ;
        RECT 520.950 775.950 523.050 778.050 ;
        RECT 515.400 767.400 519.450 768.450 ;
        RECT 515.400 763.050 516.450 767.400 ;
        RECT 497.400 760.200 498.600 760.950 ;
        RECT 503.400 760.200 504.600 762.000 ;
        RECT 506.400 761.400 510.450 762.450 ;
        RECT 493.950 757.800 496.050 759.900 ;
        RECT 496.950 757.800 499.050 759.900 ;
        RECT 499.950 757.800 502.050 759.900 ;
        RECT 502.950 757.800 505.050 759.900 ;
        RECT 494.400 755.400 495.600 757.500 ;
        RECT 500.400 756.750 501.600 757.500 ;
        RECT 494.400 751.050 495.450 755.400 ;
        RECT 499.950 754.650 502.050 756.750 ;
        RECT 496.950 753.600 501.000 754.050 ;
        RECT 496.950 751.950 502.050 753.600 ;
        RECT 502.950 751.950 505.050 754.050 ;
        RECT 499.950 751.500 502.050 751.950 ;
        RECT 490.950 749.400 495.450 751.050 ;
        RECT 490.950 748.950 495.000 749.400 ;
        RECT 503.400 745.050 504.450 751.950 ;
        RECT 509.400 745.050 510.450 761.400 ;
        RECT 514.950 760.950 517.050 763.050 ;
        RECT 517.950 762.450 520.050 766.050 ;
        RECT 521.400 762.450 522.450 775.950 ;
        RECT 542.400 775.050 543.450 799.950 ;
        RECT 545.400 796.050 546.450 811.950 ;
        RECT 566.400 811.050 567.450 820.950 ;
        RECT 598.950 817.950 601.050 820.050 ;
        RECT 565.950 808.950 568.050 811.050 ;
        RECT 571.950 808.950 577.050 811.050 ;
        RECT 547.950 805.950 550.050 808.050 ;
        RECT 556.950 806.100 559.050 808.200 ;
        RECT 562.950 806.100 565.050 808.200 ;
        RECT 577.950 807.000 580.050 811.050 ;
        RECT 544.950 793.950 547.050 796.050 ;
        RECT 535.950 772.950 538.050 775.050 ;
        RECT 541.950 772.950 544.050 775.050 ;
        RECT 517.950 762.000 522.450 762.450 ;
        RECT 518.400 761.400 522.450 762.000 ;
        RECT 518.400 760.200 519.600 761.400 ;
        RECT 523.950 760.950 526.050 763.050 ;
        RECT 536.400 762.600 537.450 772.950 ;
        RECT 541.950 766.950 544.050 769.050 ;
        RECT 542.400 762.600 543.450 766.950 ;
        RECT 545.400 766.050 546.450 793.950 ;
        RECT 548.400 778.050 549.450 805.950 ;
        RECT 557.400 805.350 558.600 806.100 ;
        RECT 563.400 805.350 564.600 806.100 ;
        RECT 578.400 805.350 579.600 807.000 ;
        RECT 583.950 806.100 586.050 808.200 ;
        RECT 599.400 807.600 600.450 817.950 ;
        RECT 605.400 808.200 606.450 820.950 ;
        RECT 610.950 811.950 613.050 814.050 ;
        RECT 584.400 805.350 585.600 806.100 ;
        RECT 599.400 805.500 600.600 807.600 ;
        RECT 604.950 806.100 607.050 808.200 ;
        RECT 611.400 808.050 612.450 811.950 ;
        RECT 620.400 811.050 621.450 820.950 ;
        RECT 628.950 817.950 631.050 820.050 ;
        RECT 688.950 817.950 691.050 820.050 ;
        RECT 619.950 808.950 622.050 811.050 ;
        RECT 610.950 805.950 613.050 808.050 ;
        RECT 616.950 806.100 619.050 808.200 ;
        RECT 622.800 806.100 624.900 808.200 ;
        RECT 617.400 805.350 618.600 806.100 ;
        RECT 623.400 805.350 624.600 806.100 ;
        RECT 553.950 802.950 556.050 805.050 ;
        RECT 556.950 802.950 559.050 805.050 ;
        RECT 559.950 802.950 562.050 805.050 ;
        RECT 562.950 802.950 565.050 805.050 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 580.950 802.950 583.050 805.050 ;
        RECT 583.950 802.950 586.050 805.050 ;
        RECT 595.950 803.100 598.050 805.200 ;
        RECT 598.950 803.100 601.050 805.200 ;
        RECT 601.950 803.100 604.050 805.200 ;
        RECT 613.950 802.950 616.050 805.050 ;
        RECT 616.950 802.950 619.050 805.050 ;
        RECT 619.950 802.950 622.050 805.050 ;
        RECT 622.950 802.950 625.050 805.050 ;
        RECT 554.400 801.000 555.600 802.650 ;
        RECT 553.950 796.950 556.050 801.000 ;
        RECT 560.400 800.400 561.600 802.650 ;
        RECT 560.400 787.050 561.450 800.400 ;
        RECT 565.950 796.950 568.050 802.050 ;
        RECT 575.400 801.000 576.600 802.650 ;
        RECT 574.950 796.950 577.050 801.000 ;
        RECT 581.400 800.400 582.600 802.650 ;
        RECT 602.400 801.450 603.600 802.800 ;
        RECT 602.400 800.400 606.450 801.450 ;
        RECT 562.950 790.950 565.050 793.050 ;
        RECT 574.950 790.950 577.050 793.050 ;
        RECT 550.950 784.950 553.050 787.050 ;
        RECT 559.950 784.950 562.050 787.050 ;
        RECT 551.400 778.050 552.450 784.950 ;
        RECT 553.950 781.950 556.050 784.050 ;
        RECT 547.800 775.950 549.900 778.050 ;
        RECT 550.950 775.950 553.050 778.050 ;
        RECT 547.950 769.950 550.050 772.050 ;
        RECT 544.950 763.950 547.050 766.050 ;
        RECT 524.400 760.200 525.600 760.950 ;
        RECT 536.400 760.350 537.600 762.600 ;
        RECT 542.400 760.350 543.600 762.600 ;
        RECT 514.950 757.800 517.050 759.900 ;
        RECT 517.950 757.800 520.050 759.900 ;
        RECT 520.950 757.800 523.050 759.900 ;
        RECT 523.950 757.800 526.050 759.900 ;
        RECT 532.950 757.950 535.050 760.050 ;
        RECT 535.950 757.950 538.050 760.050 ;
        RECT 538.950 757.950 541.050 760.050 ;
        RECT 541.950 757.950 544.050 760.050 ;
        RECT 515.400 755.400 516.600 757.500 ;
        RECT 521.400 756.750 522.600 757.500 ;
        RECT 515.400 754.050 516.450 755.400 ;
        RECT 520.950 754.650 523.050 756.750 ;
        RECT 526.950 754.950 529.050 757.050 ;
        RECT 533.400 755.400 534.600 757.650 ;
        RECT 539.400 756.900 540.600 757.650 ;
        RECT 548.400 757.050 549.450 769.950 ;
        RECT 550.950 763.950 553.050 769.050 ;
        RECT 554.400 762.450 555.450 781.950 ;
        RECT 563.400 775.050 564.450 790.950 ;
        RECT 562.950 772.950 565.050 775.050 ;
        RECT 575.400 769.050 576.450 790.950 ;
        RECT 581.400 787.050 582.450 800.400 ;
        RECT 601.950 796.950 604.050 799.050 ;
        RECT 592.950 793.950 595.050 796.050 ;
        RECT 589.950 787.950 592.050 790.050 ;
        RECT 580.950 784.950 583.050 787.050 ;
        RECT 583.950 781.950 586.050 784.050 ;
        RECT 574.800 766.950 576.900 769.050 ;
        RECT 577.950 766.950 580.050 769.050 ;
        RECT 578.400 763.050 579.450 766.950 ;
        RECT 551.400 761.400 555.450 762.450 ;
        RECT 511.950 752.550 516.450 754.050 ;
        RECT 511.950 751.950 516.000 752.550 ;
        RECT 517.950 751.950 520.050 754.050 ;
        RECT 511.950 748.800 514.050 750.900 ;
        RECT 502.950 742.950 505.050 745.050 ;
        RECT 508.950 742.950 511.050 745.050 ;
        RECT 512.400 742.050 513.450 748.800 ;
        RECT 518.400 748.050 519.450 751.950 ;
        RECT 527.400 748.050 528.450 754.950 ;
        RECT 529.950 748.950 532.050 751.050 ;
        RECT 517.950 745.950 520.050 748.050 ;
        RECT 526.950 745.950 529.050 748.050 ;
        RECT 511.950 739.950 514.050 742.050 ;
        RECT 530.400 741.450 531.450 748.950 ;
        RECT 533.400 748.050 534.450 755.400 ;
        RECT 538.950 754.800 541.050 756.900 ;
        RECT 544.950 754.950 547.050 757.050 ;
        RECT 547.950 754.950 550.050 757.050 ;
        RECT 532.950 745.950 535.050 748.050 ;
        RECT 524.400 741.000 531.450 741.450 ;
        RECT 523.950 740.400 531.450 741.000 ;
        RECT 523.950 739.050 526.050 740.400 ;
        RECT 514.950 736.950 517.050 739.050 ;
        RECT 523.800 738.000 526.050 739.050 ;
        RECT 523.800 736.950 525.900 738.000 ;
        RECT 487.950 733.950 490.050 736.050 ;
        RECT 511.950 733.950 514.050 736.050 ;
        RECT 485.400 727.500 486.600 729.600 ;
        RECT 508.950 727.950 511.050 730.050 ;
        RECT 481.950 725.100 484.050 727.200 ;
        RECT 484.950 725.100 487.050 727.200 ;
        RECT 487.950 725.100 490.050 727.200 ;
        RECT 496.950 724.950 499.050 727.050 ;
        RECT 502.950 724.950 505.050 727.050 ;
        RECT 482.400 724.050 483.600 724.800 ;
        RECT 488.400 724.050 489.600 724.800 ;
        RECT 481.950 721.950 484.050 724.050 ;
        RECT 487.950 721.950 490.050 724.050 ;
        RECT 503.400 723.900 504.600 724.650 ;
        RECT 488.400 718.050 489.450 721.950 ;
        RECT 502.950 721.800 505.050 723.900 ;
        RECT 487.950 715.950 490.050 718.050 ;
        RECT 503.400 712.050 504.450 721.800 ;
        RECT 509.400 717.450 510.450 727.950 ;
        RECT 506.400 716.400 510.450 717.450 ;
        RECT 502.950 709.950 505.050 712.050 ;
        RECT 499.950 700.950 502.050 703.050 ;
        RECT 490.950 691.950 493.050 694.050 ;
        RECT 470.400 682.350 471.600 683.100 ;
        RECT 472.950 682.950 475.050 685.050 ;
        RECT 475.950 682.950 478.050 685.050 ;
        RECT 484.950 683.100 487.050 685.200 ;
        RECT 491.400 684.600 492.450 691.950 ;
        RECT 496.950 688.950 499.050 691.050 ;
        RECT 485.400 682.350 486.600 683.100 ;
        RECT 491.400 682.350 492.600 684.600 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 475.950 679.800 478.050 681.900 ;
        RECT 481.950 679.950 484.050 682.050 ;
        RECT 484.950 679.950 487.050 682.050 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 490.950 679.950 493.050 682.050 ;
        RECT 451.950 670.950 454.050 673.050 ;
        RECT 448.950 664.950 451.050 667.050 ;
        RECT 445.950 658.050 448.050 661.050 ;
        RECT 442.950 657.000 448.050 658.050 ;
        RECT 442.950 656.400 447.450 657.000 ;
        RECT 442.950 655.950 447.000 656.400 ;
        RECT 449.400 655.050 450.450 664.950 ;
        RECT 448.950 652.950 451.050 655.050 ;
        RECT 407.400 649.350 408.600 650.100 ;
        RECT 413.400 649.350 414.600 651.600 ;
        RECT 425.400 649.500 426.600 651.600 ;
        RECT 427.950 649.950 430.050 652.050 ;
        RECT 403.950 646.950 406.050 649.050 ;
        RECT 406.950 646.950 409.050 649.050 ;
        RECT 409.950 646.950 412.050 649.050 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 421.950 647.100 424.050 649.200 ;
        RECT 424.950 647.100 427.050 649.200 ;
        RECT 436.950 647.100 439.050 649.200 ;
        RECT 442.950 647.100 445.050 649.200 ;
        RECT 445.950 647.100 448.050 649.200 ;
        RECT 452.400 649.050 453.450 670.950 ;
        RECT 455.400 664.050 456.450 677.400 ;
        RECT 460.950 676.950 463.050 679.050 ;
        RECT 467.400 677.400 468.600 679.650 ;
        RECT 467.400 670.050 468.450 677.400 ;
        RECT 472.950 676.950 475.050 679.050 ;
        RECT 466.950 667.950 469.050 670.050 ;
        RECT 454.950 661.950 457.050 664.050 ;
        RECT 463.950 661.950 466.050 664.050 ;
        RECT 464.400 652.350 465.450 661.950 ;
        RECT 463.950 650.250 466.050 652.350 ;
        RECT 464.400 649.500 465.600 650.250 ;
        RECT 451.950 646.950 454.050 649.050 ;
        RECT 460.950 647.100 463.050 649.200 ;
        RECT 463.950 647.100 466.050 649.200 ;
        RECT 466.950 647.100 469.050 649.200 ;
        RECT 404.400 645.000 405.600 646.650 ;
        RECT 410.400 645.900 411.600 646.650 ;
        RECT 422.400 646.050 423.600 646.800 ;
        RECT 403.950 640.950 406.050 645.000 ;
        RECT 409.950 643.800 412.050 645.900 ;
        RECT 421.950 643.950 424.050 646.050 ;
        RECT 437.400 644.400 438.600 646.800 ;
        RECT 446.400 644.400 447.600 646.800 ;
        RECT 467.400 644.400 468.600 646.800 ;
        RECT 437.400 643.050 438.450 644.400 ;
        RECT 436.950 640.950 439.050 643.050 ;
        RECT 433.950 631.950 436.050 634.050 ;
        RECT 400.950 625.950 403.050 628.050 ;
        RECT 397.950 619.950 400.050 622.050 ;
        RECT 388.950 607.950 391.050 610.050 ;
        RECT 394.950 607.950 397.050 610.050 ;
        RECT 382.950 606.450 385.050 607.050 ;
        RECT 380.400 605.400 385.050 606.450 ;
        RECT 382.950 604.950 385.050 605.400 ;
        RECT 385.950 604.950 388.050 607.050 ;
        RECT 383.400 604.200 384.600 604.950 ;
        RECT 373.950 601.800 376.050 603.900 ;
        RECT 376.950 601.800 379.050 603.900 ;
        RECT 379.950 601.800 382.050 603.900 ;
        RECT 382.950 601.800 385.050 603.900 ;
        RECT 368.400 599.400 372.450 600.450 ;
        RECT 355.950 591.600 358.050 592.050 ;
        RECT 362.400 591.600 363.450 599.400 ;
        RECT 367.950 595.950 370.050 598.050 ;
        RECT 355.950 591.450 363.450 591.600 ;
        RECT 355.950 591.000 366.450 591.450 ;
        RECT 355.950 590.550 367.050 591.000 ;
        RECT 355.950 589.950 358.050 590.550 ;
        RECT 362.400 590.400 367.050 590.550 ;
        RECT 355.950 586.800 358.050 588.900 ;
        RECT 364.950 586.950 367.050 590.400 ;
        RECT 346.950 580.950 349.050 583.050 ;
        RECT 356.400 577.050 357.450 586.800 ;
        RECT 368.400 580.050 369.450 595.950 ;
        RECT 367.950 577.950 370.050 580.050 ;
        RECT 371.400 577.050 372.450 599.400 ;
        RECT 374.400 599.400 375.600 601.500 ;
        RECT 380.400 599.400 381.600 601.500 ;
        RECT 374.400 583.050 375.450 599.400 ;
        RECT 380.400 592.050 381.450 599.400 ;
        RECT 385.950 598.950 388.050 601.050 ;
        RECT 379.950 589.950 382.050 592.050 ;
        RECT 373.950 580.950 376.050 583.050 ;
        RECT 386.400 580.050 387.450 598.950 ;
        RECT 389.400 597.450 390.450 607.950 ;
        RECT 401.400 607.200 402.450 625.950 ;
        RECT 391.950 606.600 396.000 607.050 ;
        RECT 391.950 604.950 396.600 606.600 ;
        RECT 400.950 605.100 403.050 607.200 ;
        RECT 412.950 606.000 415.050 610.050 ;
        RECT 434.400 606.600 435.450 631.950 ;
        RECT 437.400 625.050 438.450 640.950 ;
        RECT 446.400 634.050 447.450 644.400 ;
        RECT 467.400 640.050 468.450 644.400 ;
        RECT 466.950 637.950 469.050 640.050 ;
        RECT 466.950 634.800 469.050 636.900 ;
        RECT 445.950 631.950 448.050 634.050 ;
        RECT 436.950 622.950 439.050 625.050 ;
        RECT 437.400 613.050 438.450 622.950 ;
        RECT 439.950 619.950 442.050 622.050 ;
        RECT 436.950 610.950 439.050 613.050 ;
        RECT 440.400 607.050 441.450 619.950 ;
        RECT 442.950 610.950 445.050 613.050 ;
        RECT 395.400 604.350 396.600 604.950 ;
        RECT 401.400 604.350 402.600 605.100 ;
        RECT 413.400 604.200 414.600 606.000 ;
        RECT 434.400 604.200 435.600 606.600 ;
        RECT 439.950 604.950 442.050 607.050 ;
        RECT 443.400 606.600 444.450 610.950 ;
        RECT 446.400 610.050 447.450 631.950 ;
        RECT 445.950 607.950 448.050 610.050 ;
        RECT 443.400 604.200 444.600 606.600 ;
        RECT 454.950 606.000 457.050 610.050 ;
        RECT 467.400 607.050 468.450 634.800 ;
        RECT 469.950 610.950 472.050 613.050 ;
        RECT 455.400 604.350 456.600 606.000 ;
        RECT 460.950 604.950 463.050 607.050 ;
        RECT 466.950 604.950 469.050 607.050 ;
        RECT 461.400 604.350 462.600 604.950 ;
        RECT 394.950 601.950 397.050 604.050 ;
        RECT 397.950 601.950 400.050 604.050 ;
        RECT 400.950 601.950 403.050 604.050 ;
        RECT 403.950 601.950 406.050 604.050 ;
        RECT 412.950 601.800 415.050 603.900 ;
        RECT 415.950 601.800 418.050 603.900 ;
        RECT 418.950 601.800 421.050 603.900 ;
        RECT 433.950 601.800 436.050 603.900 ;
        RECT 436.950 601.800 439.050 603.900 ;
        RECT 442.950 601.800 445.050 603.900 ;
        RECT 454.950 601.950 457.050 604.050 ;
        RECT 457.950 601.950 460.050 604.050 ;
        RECT 460.950 601.950 463.050 604.050 ;
        RECT 463.950 601.950 466.050 604.050 ;
        RECT 398.400 599.400 399.600 601.650 ;
        RECT 404.400 600.000 405.600 601.650 ;
        RECT 398.400 597.450 399.450 599.400 ;
        RECT 389.400 596.400 393.450 597.450 ;
        RECT 392.400 583.050 393.450 596.400 ;
        RECT 395.400 596.400 399.450 597.450 ;
        RECT 395.400 592.050 396.450 596.400 ;
        RECT 403.950 595.950 406.050 600.000 ;
        RECT 416.400 599.400 417.600 601.500 ;
        RECT 416.400 598.050 417.450 599.400 ;
        RECT 445.950 598.950 448.050 601.050 ;
        RECT 451.950 598.950 454.050 601.050 ;
        RECT 458.400 600.900 459.600 601.650 ;
        RECT 409.800 595.950 411.900 598.050 ;
        RECT 412.950 596.400 417.450 598.050 ;
        RECT 412.950 595.950 417.000 596.400 ;
        RECT 418.950 595.950 421.050 598.050 ;
        RECT 397.950 592.950 400.050 595.050 ;
        RECT 394.950 589.950 397.050 592.050 ;
        RECT 391.950 580.950 394.050 583.050 ;
        RECT 385.950 577.950 388.050 580.050 ;
        RECT 355.950 574.950 358.050 577.050 ;
        RECT 364.950 576.450 369.000 577.050 ;
        RECT 364.950 574.950 369.450 576.450 ;
        RECT 370.950 574.950 373.050 577.050 ;
        RECT 326.400 571.350 327.600 571.950 ;
        RECT 332.400 571.350 333.600 573.600 ;
        RECT 343.950 571.950 346.050 574.050 ;
        RECT 352.950 572.250 355.050 574.350 ;
        RECT 368.400 573.600 369.450 574.950 ;
        RECT 325.950 568.950 328.050 571.050 ;
        RECT 328.950 568.950 331.050 571.050 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 322.950 565.950 325.050 568.050 ;
        RECT 329.400 566.400 330.600 568.650 ;
        RECT 335.400 567.900 336.600 568.650 ;
        RECT 323.400 562.050 324.450 565.950 ;
        RECT 325.950 562.950 328.050 565.050 ;
        RECT 322.950 559.950 325.050 562.050 ;
        RECT 319.950 544.950 322.050 547.050 ;
        RECT 316.950 535.950 319.050 538.050 ;
        RECT 317.400 528.600 318.450 535.950 ;
        RECT 326.400 532.050 327.450 562.950 ;
        RECT 329.400 532.050 330.450 566.400 ;
        RECT 334.950 565.800 337.050 567.900 ;
        RECT 335.400 556.050 336.450 565.800 ;
        RECT 344.400 565.050 345.450 571.950 ;
        RECT 353.400 571.500 354.600 572.250 ;
        RECT 368.400 571.500 369.600 573.600 ;
        RECT 373.950 572.250 376.050 574.350 ;
        RECT 386.400 573.600 387.450 577.950 ;
        RECT 374.400 571.500 375.600 572.250 ;
        RECT 386.400 571.350 387.600 573.600 ;
        RECT 394.950 572.250 397.050 574.350 ;
        RECT 398.400 574.050 399.450 592.950 ;
        RECT 410.400 589.050 411.450 595.950 ;
        RECT 419.400 589.050 420.450 595.950 ;
        RECT 430.950 589.950 433.050 592.050 ;
        RECT 409.800 586.950 411.900 589.050 ;
        RECT 412.950 586.950 415.050 589.050 ;
        RECT 418.950 586.950 421.050 589.050 ;
        RECT 349.950 569.100 352.050 571.200 ;
        RECT 352.950 569.100 355.050 571.200 ;
        RECT 355.950 569.100 358.050 571.200 ;
        RECT 367.950 569.100 370.050 571.200 ;
        RECT 370.950 569.100 373.050 571.200 ;
        RECT 373.950 569.100 376.050 571.200 ;
        RECT 376.950 569.100 379.050 571.200 ;
        RECT 385.950 568.950 388.050 571.050 ;
        RECT 388.950 568.950 391.050 571.050 ;
        RECT 350.400 568.050 351.600 568.800 ;
        RECT 356.400 568.050 357.600 568.800 ;
        RECT 349.950 565.950 352.050 568.050 ;
        RECT 355.950 565.950 358.050 568.050 ;
        RECT 364.950 565.950 367.050 568.050 ;
        RECT 371.400 567.000 372.600 568.800 ;
        RECT 343.950 562.950 346.050 565.050 ;
        RECT 334.950 553.950 337.050 556.050 ;
        RECT 331.950 550.950 334.050 553.050 ;
        RECT 349.950 550.950 352.050 553.050 ;
        RECT 325.950 529.950 328.050 532.050 ;
        RECT 328.950 529.950 331.050 532.050 ;
        RECT 317.400 526.350 318.600 528.600 ;
        RECT 323.400 528.450 324.600 528.600 ;
        RECT 323.400 527.400 330.450 528.450 ;
        RECT 323.400 526.350 324.600 527.400 ;
        RECT 313.950 523.950 316.050 526.050 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 319.950 523.950 322.050 526.050 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 314.400 522.900 315.600 523.650 ;
        RECT 308.400 521.400 312.450 522.450 ;
        RECT 307.950 517.950 310.050 520.050 ;
        RECT 308.400 508.050 309.450 517.950 ;
        RECT 307.950 505.950 310.050 508.050 ;
        RECT 304.950 502.950 307.050 505.050 ;
        RECT 305.400 499.050 306.450 502.950 ;
        RECT 307.950 499.950 310.050 502.050 ;
        RECT 292.950 496.950 295.050 499.050 ;
        RECT 304.950 496.950 307.050 499.050 ;
        RECT 289.950 494.100 292.050 496.200 ;
        RECT 301.950 494.250 304.050 496.350 ;
        RECT 308.400 495.600 309.450 499.950 ;
        RECT 311.400 496.050 312.450 521.400 ;
        RECT 313.950 520.800 316.050 522.900 ;
        RECT 320.400 521.400 321.600 523.650 ;
        RECT 329.400 522.450 330.450 527.400 ;
        RECT 326.400 521.400 330.450 522.450 ;
        RECT 284.400 493.350 285.600 494.100 ;
        RECT 290.400 493.350 291.600 494.100 ;
        RECT 302.400 493.500 303.600 494.250 ;
        RECT 308.400 493.500 309.600 495.600 ;
        RECT 310.950 493.950 313.050 496.050 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 286.950 490.950 289.050 493.050 ;
        RECT 289.950 490.950 292.050 493.050 ;
        RECT 298.950 491.100 301.050 493.200 ;
        RECT 301.950 491.100 304.050 493.200 ;
        RECT 304.950 491.100 307.050 493.200 ;
        RECT 307.950 491.100 310.050 493.200 ;
        RECT 287.400 488.400 288.600 490.650 ;
        RECT 299.400 490.050 300.600 490.800 ;
        RECT 283.950 466.950 286.050 469.050 ;
        RECT 280.950 451.950 283.050 454.050 ;
        RECT 277.950 442.950 280.050 445.050 ;
        RECT 232.950 438.450 235.050 439.050 ;
        RECT 232.950 437.400 237.450 438.450 ;
        RECT 232.950 436.950 235.050 437.400 ;
        RECT 217.950 418.950 220.050 421.050 ;
        RECT 223.950 418.950 226.050 421.050 ;
        RECT 188.400 415.500 189.600 416.250 ;
        RECT 203.400 415.500 204.600 416.250 ;
        RECT 209.400 415.500 210.600 417.600 ;
        RECT 184.950 413.100 187.050 415.200 ;
        RECT 187.950 413.100 190.050 415.200 ;
        RECT 190.950 413.100 193.050 415.200 ;
        RECT 199.950 413.100 202.050 415.200 ;
        RECT 202.950 413.100 205.050 415.200 ;
        RECT 205.950 413.100 208.050 415.200 ;
        RECT 208.950 413.100 211.050 415.200 ;
        RECT 211.950 413.100 214.050 415.200 ;
        RECT 185.400 412.050 186.600 412.800 ;
        RECT 185.400 410.400 190.050 412.050 ;
        RECT 186.000 409.950 190.050 410.400 ;
        RECT 191.400 410.400 192.600 412.800 ;
        RECT 200.400 410.400 201.600 412.800 ;
        RECT 206.400 410.400 207.600 412.800 ;
        RECT 212.400 412.050 213.600 412.800 ;
        RECT 191.400 403.050 192.450 410.400 ;
        RECT 190.950 400.950 193.050 403.050 ;
        RECT 187.950 394.950 190.050 397.050 ;
        RECT 188.400 391.050 189.450 394.950 ;
        RECT 200.400 391.050 201.450 410.400 ;
        RECT 206.400 397.050 207.450 410.400 ;
        RECT 211.950 409.950 214.050 412.050 ;
        RECT 212.400 406.050 213.450 409.950 ;
        RECT 211.950 403.950 214.050 406.050 ;
        RECT 218.400 400.050 219.450 418.950 ;
        RECT 226.950 416.250 229.050 418.350 ;
        RECT 227.400 415.500 228.600 416.250 ;
        RECT 223.950 413.100 226.050 415.200 ;
        RECT 226.950 413.100 229.050 415.200 ;
        RECT 229.950 413.100 232.050 415.200 ;
        RECT 224.400 410.400 225.600 412.800 ;
        RECT 230.400 412.050 231.600 412.800 ;
        RECT 236.400 412.050 237.450 437.400 ;
        RECT 241.950 436.950 244.050 439.050 ;
        RECT 266.400 437.400 267.600 440.100 ;
        RECT 269.400 438.600 271.500 440.700 ;
        RECT 266.400 433.050 267.450 437.400 ;
        RECT 265.950 430.950 268.050 433.050 ;
        RECT 271.950 430.950 274.050 433.050 ;
        RECT 256.950 427.950 259.050 430.050 ;
        RECT 268.950 427.950 271.050 430.050 ;
        RECT 257.400 424.050 258.450 427.950 ;
        RECT 256.950 421.950 259.050 424.050 ;
        RECT 238.950 415.950 241.050 418.050 ;
        RECT 247.950 417.000 250.050 421.050 ;
        RECT 217.950 397.950 220.050 400.050 ;
        RECT 224.400 397.050 225.450 410.400 ;
        RECT 229.950 409.950 232.050 412.050 ;
        RECT 235.950 409.950 238.050 412.050 ;
        RECT 205.950 394.950 208.050 397.050 ;
        RECT 223.950 394.950 226.050 397.050 ;
        RECT 224.400 391.050 225.450 394.950 ;
        RECT 239.400 394.050 240.450 415.950 ;
        RECT 248.400 415.500 249.600 417.000 ;
        RECT 253.950 415.950 256.050 421.050 ;
        RECT 244.950 413.100 247.050 415.200 ;
        RECT 247.950 413.100 250.050 415.200 ;
        RECT 250.950 413.100 253.050 415.200 ;
        RECT 245.400 412.050 246.600 412.800 ;
        RECT 244.950 409.950 247.050 412.050 ;
        RECT 251.400 410.400 252.600 412.800 ;
        RECT 251.400 406.050 252.450 410.400 ;
        RECT 253.950 409.950 256.050 412.050 ;
        RECT 250.950 403.950 253.050 406.050 ;
        RECT 238.950 391.950 241.050 394.050 ;
        RECT 187.950 388.950 190.050 391.050 ;
        RECT 199.950 388.950 202.050 391.050 ;
        RECT 223.950 388.950 226.050 391.050 ;
        RECT 205.950 380.400 208.050 382.500 ;
        RECT 226.950 381.300 229.050 383.400 ;
        RECT 254.400 382.050 255.450 409.950 ;
        RECT 257.400 397.050 258.450 421.950 ;
        RECT 269.400 421.050 270.450 427.950 ;
        RECT 268.950 418.950 271.050 421.050 ;
        RECT 272.400 418.200 273.450 430.950 ;
        RECT 281.400 430.050 282.450 451.950 ;
        RECT 284.400 451.050 285.450 466.950 ;
        RECT 287.400 454.050 288.450 488.400 ;
        RECT 292.950 484.950 295.050 490.050 ;
        RECT 298.950 487.950 301.050 490.050 ;
        RECT 305.400 489.000 306.600 490.800 ;
        RECT 304.950 484.950 307.050 489.000 ;
        RECT 307.950 487.950 310.050 490.050 ;
        RECT 308.400 478.050 309.450 487.950 ;
        RECT 310.950 478.950 313.050 481.050 ;
        RECT 298.950 475.950 301.050 478.050 ;
        RECT 307.950 475.950 310.050 478.050 ;
        RECT 299.400 460.050 300.450 475.950 ;
        RECT 311.400 474.450 312.450 478.950 ;
        RECT 314.400 475.050 315.450 520.800 ;
        RECT 320.400 517.050 321.450 521.400 ;
        RECT 319.950 514.950 322.050 517.050 ;
        RECT 316.950 513.450 321.000 514.050 ;
        RECT 316.950 513.000 321.450 513.450 ;
        RECT 316.950 511.950 322.050 513.000 ;
        RECT 319.950 508.950 322.050 511.950 ;
        RECT 316.950 505.950 319.050 508.050 ;
        RECT 317.400 484.050 318.450 505.950 ;
        RECT 326.400 495.600 327.450 521.400 ;
        RECT 332.400 517.050 333.450 550.950 ;
        RECT 343.950 547.950 346.050 550.050 ;
        RECT 344.400 528.600 345.450 547.950 ;
        RECT 346.950 544.950 349.050 547.050 ;
        RECT 347.400 538.050 348.450 544.950 ;
        RECT 350.400 544.050 351.450 550.950 ;
        RECT 361.950 547.950 364.050 550.050 ;
        RECT 349.950 541.950 352.050 544.050 ;
        RECT 362.400 538.050 363.450 547.950 ;
        RECT 346.950 535.950 349.050 538.050 ;
        RECT 361.950 535.950 364.050 538.050 ;
        RECT 349.950 532.950 352.050 535.050 ;
        RECT 344.400 526.200 345.600 528.600 ;
        RECT 337.950 523.800 340.050 525.900 ;
        RECT 340.950 523.800 343.050 525.900 ;
        RECT 343.950 523.800 346.050 525.900 ;
        RECT 334.950 517.950 337.050 523.050 ;
        RECT 341.400 522.750 342.600 523.500 ;
        RECT 340.950 520.650 343.050 522.750 ;
        RECT 331.950 514.950 334.050 517.050 ;
        RECT 328.950 508.950 331.050 514.050 ;
        RECT 334.950 513.600 339.000 514.050 ;
        RECT 334.950 511.950 339.450 513.600 ;
        RECT 338.400 508.050 339.450 511.950 ;
        RECT 337.950 505.950 340.050 508.050 ;
        RECT 337.950 502.800 340.050 504.900 ;
        RECT 338.400 499.050 339.450 502.800 ;
        RECT 337.950 496.950 340.050 499.050 ;
        RECT 326.400 493.350 327.600 495.600 ;
        RECT 331.800 494.100 333.900 496.200 ;
        RECT 341.400 495.450 342.450 520.650 ;
        RECT 346.950 511.950 349.050 514.050 ;
        RECT 338.400 494.400 342.450 495.450 ;
        RECT 347.400 495.600 348.450 511.950 ;
        RECT 350.400 505.050 351.450 532.950 ;
        RECT 362.400 528.600 363.450 535.950 ;
        RECT 365.400 529.050 366.450 565.950 ;
        RECT 370.950 562.950 373.050 567.000 ;
        RECT 377.400 566.400 378.600 568.800 ;
        RECT 373.950 550.950 376.050 553.050 ;
        RECT 374.400 547.050 375.450 550.950 ;
        RECT 367.950 544.950 370.050 547.050 ;
        RECT 373.950 544.950 376.050 547.050 ;
        RECT 368.400 532.050 369.450 544.950 ;
        RECT 377.400 532.050 378.450 566.400 ;
        RECT 379.950 565.950 382.050 568.050 ;
        RECT 389.400 567.900 390.600 568.650 ;
        RECT 395.400 568.050 396.450 572.250 ;
        RECT 397.950 571.950 400.050 574.050 ;
        RECT 403.950 573.000 406.050 577.050 ;
        RECT 410.400 574.050 411.450 586.950 ;
        RECT 404.400 571.500 405.600 573.000 ;
        RECT 409.950 571.950 412.050 574.050 ;
        RECT 400.950 569.100 403.050 571.200 ;
        RECT 403.950 569.100 406.050 571.200 ;
        RECT 406.950 569.100 409.050 571.200 ;
        RECT 380.400 559.050 381.450 565.950 ;
        RECT 388.950 565.800 391.050 567.900 ;
        RECT 391.950 565.950 394.050 568.050 ;
        RECT 394.950 565.950 397.050 568.050 ;
        RECT 401.400 567.450 402.600 568.800 ;
        RECT 398.400 566.400 402.600 567.450 ;
        RECT 382.950 559.950 385.050 562.050 ;
        RECT 379.950 556.950 382.050 559.050 ;
        RECT 367.950 529.950 370.050 532.050 ;
        RECT 362.400 526.200 363.600 528.600 ;
        RECT 364.950 526.950 367.050 529.050 ;
        RECT 355.950 523.800 358.050 525.900 ;
        RECT 358.950 523.800 361.050 525.900 ;
        RECT 361.950 523.800 364.050 525.900 ;
        RECT 359.400 522.750 360.600 523.500 ;
        RECT 368.400 523.050 369.450 529.950 ;
        RECT 373.950 528.000 376.050 532.050 ;
        RECT 376.950 529.950 379.050 532.050 ;
        RECT 380.400 528.600 381.450 556.950 ;
        RECT 383.400 556.050 384.450 559.950 ;
        RECT 382.950 553.950 385.050 556.050 ;
        RECT 385.950 547.950 388.050 550.050 ;
        RECT 386.400 529.050 387.450 547.950 ;
        RECT 392.400 535.050 393.450 565.950 ;
        RECT 398.400 547.050 399.450 566.400 ;
        RECT 409.950 565.950 412.050 568.050 ;
        RECT 406.950 556.950 409.050 559.050 ;
        RECT 400.950 553.950 403.050 556.050 ;
        RECT 397.950 544.950 400.050 547.050 ;
        RECT 397.950 538.950 400.050 541.050 ;
        RECT 391.800 532.950 393.900 535.050 ;
        RECT 374.400 526.350 375.600 528.000 ;
        RECT 380.400 526.350 381.600 528.600 ;
        RECT 385.950 526.950 388.050 529.050 ;
        RECT 398.400 528.600 399.450 538.950 ;
        RECT 401.400 529.050 402.450 553.950 ;
        RECT 403.950 550.950 406.050 553.050 ;
        RECT 404.400 538.050 405.450 550.950 ;
        RECT 407.400 547.050 408.450 556.950 ;
        RECT 410.400 550.050 411.450 565.950 ;
        RECT 413.400 553.050 414.450 586.950 ;
        RECT 415.950 580.950 418.050 583.050 ;
        RECT 416.400 562.050 417.450 580.950 ;
        RECT 424.950 572.100 427.050 574.200 ;
        RECT 431.400 573.600 432.450 589.950 ;
        RECT 446.400 586.050 447.450 598.950 ;
        RECT 445.950 583.950 448.050 586.050 ;
        RECT 452.400 583.050 453.450 598.950 ;
        RECT 457.950 598.800 460.050 600.900 ;
        RECT 464.400 599.400 465.600 601.650 ;
        RECT 470.400 601.050 471.450 610.950 ;
        RECT 473.400 607.050 474.450 676.950 ;
        RECT 476.400 676.050 477.450 679.800 ;
        RECT 478.950 676.950 481.050 679.050 ;
        RECT 482.400 678.000 483.600 679.650 ;
        RECT 488.400 678.900 489.600 679.650 ;
        RECT 497.400 679.050 498.450 688.950 ;
        RECT 500.400 685.050 501.450 700.950 ;
        RECT 506.400 699.450 507.450 716.400 ;
        RECT 512.400 703.050 513.450 733.950 ;
        RECT 515.400 730.050 516.450 736.950 ;
        RECT 531.000 732.450 535.050 733.050 ;
        RECT 530.400 730.950 535.050 732.450 ;
        RECT 514.950 727.950 517.050 730.050 ;
        RECT 520.950 728.100 523.050 730.200 ;
        RECT 530.400 729.600 531.450 730.950 ;
        RECT 521.400 727.350 522.600 728.100 ;
        RECT 530.400 727.350 531.600 729.600 ;
        RECT 535.950 728.100 538.050 730.200 ;
        RECT 536.400 727.350 537.600 728.100 ;
        RECT 517.950 724.950 520.050 727.050 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 535.950 724.950 538.050 727.050 ;
        RECT 538.950 724.950 541.050 727.050 ;
        RECT 518.400 722.400 519.600 724.650 ;
        RECT 533.400 722.400 534.600 724.650 ;
        RECT 539.400 724.050 540.600 724.650 ;
        RECT 539.400 722.400 544.050 724.050 ;
        RECT 514.950 718.950 517.050 721.050 ;
        RECT 518.400 720.450 519.450 722.400 ;
        RECT 518.400 720.000 522.450 720.450 ;
        RECT 518.400 719.400 523.050 720.000 ;
        RECT 511.950 700.950 514.050 703.050 ;
        RECT 515.400 699.450 516.450 718.950 ;
        RECT 517.800 715.950 519.900 718.050 ;
        RECT 520.950 715.950 523.050 719.400 ;
        RECT 506.400 698.400 510.450 699.450 ;
        RECT 505.950 694.950 508.050 697.050 ;
        RECT 499.950 682.950 502.050 685.050 ;
        RECT 506.400 684.600 507.450 694.950 ;
        RECT 509.400 685.050 510.450 698.400 ;
        RECT 512.400 698.400 516.450 699.450 ;
        RECT 506.400 682.350 507.600 684.600 ;
        RECT 508.950 682.950 511.050 685.050 ;
        RECT 502.950 679.950 505.050 682.050 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 475.950 673.950 478.050 676.050 ;
        RECT 479.400 651.600 480.450 676.950 ;
        RECT 481.950 673.950 484.050 678.000 ;
        RECT 487.950 676.800 490.050 678.900 ;
        RECT 493.950 676.950 496.050 679.050 ;
        RECT 496.950 676.950 499.050 679.050 ;
        RECT 503.400 677.400 504.600 679.650 ;
        RECT 494.400 673.050 495.450 676.950 ;
        RECT 493.950 670.950 496.050 673.050 ;
        RECT 503.400 664.050 504.450 677.400 ;
        RECT 502.950 661.950 505.050 664.050 ;
        RECT 484.950 655.950 487.050 658.050 ;
        RECT 502.950 655.950 505.050 658.050 ;
        RECT 485.400 651.600 486.450 655.950 ;
        RECT 498.000 654.450 502.050 655.050 ;
        RECT 497.400 652.950 502.050 654.450 ;
        RECT 497.400 651.600 498.450 652.950 ;
        RECT 503.400 651.600 504.450 655.950 ;
        RECT 479.400 649.500 480.600 651.600 ;
        RECT 485.400 649.500 486.600 651.600 ;
        RECT 497.400 649.350 498.600 651.600 ;
        RECT 503.400 649.350 504.600 651.600 ;
        RECT 478.950 647.100 481.050 649.200 ;
        RECT 481.950 647.100 484.050 649.200 ;
        RECT 484.950 647.100 487.050 649.200 ;
        RECT 487.950 647.100 490.050 649.200 ;
        RECT 496.950 646.950 499.050 649.050 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 502.950 646.950 505.050 649.050 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 482.400 644.400 483.600 646.800 ;
        RECT 488.400 646.050 489.600 646.800 ;
        RECT 475.950 637.950 478.050 640.050 ;
        RECT 476.400 619.050 477.450 637.950 ;
        RECT 482.400 637.050 483.450 644.400 ;
        RECT 487.950 643.950 490.050 646.050 ;
        RECT 500.400 644.400 501.600 646.650 ;
        RECT 506.400 644.400 507.600 646.650 ;
        RECT 512.400 646.050 513.450 698.400 ;
        RECT 514.950 694.950 517.050 697.050 ;
        RECT 515.400 670.050 516.450 694.950 ;
        RECT 518.400 685.050 519.450 715.950 ;
        RECT 521.400 694.050 522.450 715.950 ;
        RECT 533.400 700.050 534.450 722.400 ;
        RECT 540.000 721.950 544.050 722.400 ;
        RECT 538.950 715.950 541.050 718.050 ;
        RECT 539.400 709.050 540.450 715.950 ;
        RECT 541.950 712.950 544.050 715.050 ;
        RECT 538.950 706.950 541.050 709.050 ;
        RECT 532.950 697.950 535.050 700.050 ;
        RECT 538.950 697.950 541.050 700.050 ;
        RECT 520.950 691.950 523.050 694.050 ;
        RECT 539.400 691.050 540.450 697.950 ;
        RECT 538.950 688.950 541.050 691.050 ;
        RECT 517.950 682.950 520.050 685.050 ;
        RECT 523.950 682.800 526.050 684.900 ;
        RECT 529.950 684.000 532.050 688.050 ;
        RECT 532.800 687.000 534.900 688.050 ;
        RECT 535.950 687.900 540.000 688.050 ;
        RECT 532.800 685.950 535.050 687.000 ;
        RECT 535.950 685.950 541.050 687.900 ;
        RECT 524.400 682.200 525.600 682.800 ;
        RECT 530.400 682.200 531.600 684.000 ;
        RECT 532.950 682.950 535.050 685.950 ;
        RECT 538.950 685.800 541.050 685.950 ;
        RECT 538.950 682.800 541.050 684.900 ;
        RECT 542.400 684.450 543.450 712.950 ;
        RECT 545.400 697.050 546.450 754.950 ;
        RECT 551.400 750.450 552.450 761.400 ;
        RECT 556.950 760.950 559.050 763.050 ;
        RECT 565.950 760.950 568.050 763.050 ;
        RECT 577.950 760.950 580.050 763.050 ;
        RECT 584.400 762.600 585.450 781.950 ;
        RECT 590.400 772.050 591.450 787.950 ;
        RECT 593.400 778.050 594.450 793.950 ;
        RECT 602.400 790.050 603.450 796.950 ;
        RECT 605.400 793.050 606.450 800.400 ;
        RECT 614.400 800.400 615.600 802.650 ;
        RECT 620.400 800.400 621.600 802.650 ;
        RECT 614.400 793.050 615.450 800.400 ;
        RECT 620.400 796.050 621.450 800.400 ;
        RECT 625.950 799.950 628.050 802.050 ;
        RECT 619.950 793.950 622.050 796.050 ;
        RECT 604.950 790.950 607.050 793.050 ;
        RECT 613.950 790.950 616.050 793.050 ;
        RECT 601.950 787.950 604.050 790.050 ;
        RECT 610.950 784.950 613.050 787.050 ;
        RECT 592.950 775.950 595.050 778.050 ;
        RECT 598.950 772.950 601.050 775.050 ;
        RECT 589.950 769.950 592.050 772.050 ;
        RECT 599.400 766.050 600.450 772.950 ;
        RECT 586.950 763.950 592.050 766.050 ;
        RECT 598.950 763.950 601.050 766.050 ;
        RECT 557.400 760.200 558.600 760.950 ;
        RECT 566.400 760.200 567.600 760.950 ;
        RECT 578.400 760.200 579.600 760.950 ;
        RECT 584.400 760.200 585.600 762.600 ;
        RECT 589.950 760.800 592.050 762.900 ;
        RECT 595.950 760.950 598.050 763.050 ;
        RECT 601.950 760.950 604.050 763.050 ;
        RECT 607.950 762.000 610.050 766.050 ;
        RECT 611.400 763.050 612.450 784.950 ;
        RECT 614.400 769.050 615.450 790.950 ;
        RECT 613.950 766.950 616.050 769.050 ;
        RECT 614.400 763.050 615.450 766.950 ;
        RECT 590.400 760.200 591.600 760.800 ;
        RECT 556.950 757.800 559.050 759.900 ;
        RECT 559.950 757.800 562.050 759.900 ;
        RECT 565.950 757.800 568.050 759.900 ;
        RECT 577.950 757.800 580.050 759.900 ;
        RECT 580.950 757.800 583.050 759.900 ;
        RECT 583.950 757.800 586.050 759.900 ;
        RECT 586.950 757.800 589.050 759.900 ;
        RECT 589.950 757.800 592.050 759.900 ;
        RECT 560.400 755.400 561.600 757.500 ;
        RECT 560.400 751.050 561.450 755.400 ;
        RECT 568.950 754.950 571.050 757.050 ;
        RECT 574.950 754.950 577.050 757.050 ;
        RECT 581.400 755.400 582.600 757.500 ;
        RECT 587.400 756.750 588.600 757.500 ;
        RECT 548.400 749.400 552.450 750.450 ;
        RECT 548.400 730.050 549.450 749.400 ;
        RECT 559.950 748.950 562.050 751.050 ;
        RECT 550.950 745.950 553.050 748.050 ;
        RECT 547.950 727.950 550.050 730.050 ;
        RECT 551.400 729.600 552.450 745.950 ;
        RECT 560.400 745.050 561.450 748.950 ;
        RECT 562.950 745.950 565.050 748.050 ;
        RECT 559.950 742.950 562.050 745.050 ;
        RECT 563.400 739.050 564.450 745.950 ;
        RECT 562.950 736.950 565.050 739.050 ;
        RECT 553.950 732.450 556.050 733.050 ;
        RECT 559.950 732.450 562.050 733.050 ;
        RECT 553.950 732.000 564.450 732.450 ;
        RECT 553.950 731.400 565.050 732.000 ;
        RECT 553.950 730.950 556.050 731.400 ;
        RECT 559.950 730.950 562.050 731.400 ;
        RECT 551.400 727.350 552.600 729.600 ;
        RECT 556.950 728.100 559.050 730.200 ;
        RECT 557.400 727.350 558.600 728.100 ;
        RECT 562.950 727.950 565.050 731.400 ;
        RECT 569.400 729.450 570.450 754.950 ;
        RECT 575.400 736.050 576.450 754.950 ;
        RECT 581.400 751.050 582.450 755.400 ;
        RECT 586.950 754.650 589.050 756.750 ;
        RECT 587.400 753.450 588.450 754.650 ;
        RECT 587.400 752.400 591.450 753.450 ;
        RECT 580.800 748.950 582.900 751.050 ;
        RECT 583.950 748.050 586.050 751.050 ;
        RECT 582.000 747.900 586.050 748.050 ;
        RECT 580.950 747.000 586.050 747.900 ;
        RECT 580.950 746.400 585.450 747.000 ;
        RECT 580.950 745.950 585.000 746.400 ;
        RECT 580.950 745.800 583.050 745.950 ;
        RECT 583.950 742.950 586.050 745.050 ;
        RECT 580.950 736.950 583.050 739.050 ;
        RECT 574.950 733.950 577.050 736.050 ;
        RECT 566.400 728.400 570.450 729.450 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 556.950 724.950 559.050 727.050 ;
        RECT 559.950 724.950 562.050 727.050 ;
        RECT 554.400 723.900 555.600 724.650 ;
        RECT 553.950 721.800 556.050 723.900 ;
        RECT 560.400 722.400 561.600 724.650 ;
        RECT 554.400 709.050 555.450 721.800 ;
        RECT 560.400 715.050 561.450 722.400 ;
        RECT 562.950 718.950 565.050 724.050 ;
        RECT 559.950 712.950 562.050 715.050 ;
        RECT 553.950 706.950 556.050 709.050 ;
        RECT 547.950 703.950 550.050 706.050 ;
        RECT 552.000 705.900 555.000 706.050 ;
        RECT 552.000 705.450 556.050 705.900 ;
        RECT 551.400 703.950 556.050 705.450 ;
        RECT 544.950 694.950 547.050 697.050 ;
        RECT 548.400 691.050 549.450 703.950 ;
        RECT 547.950 688.950 550.050 691.050 ;
        RECT 545.400 684.450 546.600 684.600 ;
        RECT 542.400 683.400 546.600 684.450 ;
        RECT 539.400 682.200 540.600 682.800 ;
        RECT 545.400 682.200 546.600 683.400 ;
        RECT 520.950 679.800 523.050 681.900 ;
        RECT 523.950 679.800 526.050 681.900 ;
        RECT 526.950 679.800 529.050 681.900 ;
        RECT 529.950 679.800 532.050 681.900 ;
        RECT 538.950 679.800 541.050 681.900 ;
        RECT 541.950 679.800 544.050 681.900 ;
        RECT 544.950 679.800 547.050 681.900 ;
        RECT 517.950 676.950 520.050 679.050 ;
        RECT 521.400 678.750 522.600 679.500 ;
        RECT 514.950 667.950 517.050 670.050 ;
        RECT 518.400 658.050 519.450 676.950 ;
        RECT 520.950 676.650 523.050 678.750 ;
        RECT 527.400 677.400 528.600 679.500 ;
        RECT 520.950 673.500 523.050 675.600 ;
        RECT 517.950 655.950 520.050 658.050 ;
        RECT 521.400 651.600 522.450 673.500 ;
        RECT 527.400 670.050 528.450 677.400 ;
        RECT 535.950 676.950 538.050 679.050 ;
        RECT 542.400 678.750 543.600 679.500 ;
        RECT 551.400 679.050 552.450 703.950 ;
        RECT 553.950 703.800 556.050 703.950 ;
        RECT 562.950 694.950 565.050 697.050 ;
        RECT 559.950 688.950 562.050 691.050 ;
        RECT 560.400 684.600 561.450 688.950 ;
        RECT 563.400 685.050 564.450 694.950 ;
        RECT 566.400 688.050 567.450 728.400 ;
        RECT 574.950 728.250 577.050 730.350 ;
        RECT 581.400 729.600 582.450 736.950 ;
        RECT 584.400 730.050 585.450 742.950 ;
        RECT 586.950 739.950 589.050 742.050 ;
        RECT 587.400 736.050 588.450 739.950 ;
        RECT 586.950 733.950 589.050 736.050 ;
        RECT 575.400 727.500 576.600 728.250 ;
        RECT 581.400 727.500 582.600 729.600 ;
        RECT 583.950 727.950 586.050 730.050 ;
        RECT 571.950 725.100 574.050 727.200 ;
        RECT 574.950 725.100 577.050 727.200 ;
        RECT 577.950 725.100 580.050 727.200 ;
        RECT 580.950 725.100 583.050 727.200 ;
        RECT 572.400 724.050 573.600 724.800 ;
        RECT 578.400 724.050 579.600 724.800 ;
        RECT 568.950 721.950 571.050 724.050 ;
        RECT 571.950 721.950 574.050 724.050 ;
        RECT 577.950 721.950 580.050 724.050 ;
        RECT 583.950 721.950 586.050 724.050 ;
        RECT 565.950 685.950 568.050 688.050 ;
        RECT 560.400 682.350 561.600 684.600 ;
        RECT 562.950 682.950 565.050 685.050 ;
        RECT 569.400 684.450 570.450 721.950 ;
        RECT 577.950 718.800 580.050 720.900 ;
        RECT 578.400 697.050 579.450 718.800 ;
        RECT 584.400 703.050 585.450 721.950 ;
        RECT 587.400 712.050 588.450 733.950 ;
        RECT 590.400 724.050 591.450 752.400 ;
        RECT 596.400 733.050 597.450 760.950 ;
        RECT 602.400 760.200 603.600 760.950 ;
        RECT 608.400 760.200 609.600 762.000 ;
        RECT 610.800 760.950 612.900 763.050 ;
        RECT 613.950 760.950 616.050 763.050 ;
        RECT 620.400 762.600 621.450 793.950 ;
        RECT 626.400 784.050 627.450 799.950 ;
        RECT 629.400 793.050 630.450 817.950 ;
        RECT 661.950 811.950 664.050 814.050 ;
        RECT 682.800 811.950 684.900 814.050 ;
        RECT 634.950 807.000 637.050 811.050 ;
        RECT 640.950 807.000 643.050 811.050 ;
        RECT 635.400 805.500 636.600 807.000 ;
        RECT 641.400 805.500 642.600 807.000 ;
        RECT 649.950 805.950 652.050 808.050 ;
        RECT 655.950 806.250 658.050 808.350 ;
        RECT 662.400 807.600 663.450 811.950 ;
        RECT 683.400 808.350 684.450 811.950 ;
        RECT 634.950 803.100 637.050 805.200 ;
        RECT 637.950 803.100 640.050 805.200 ;
        RECT 640.950 803.100 643.050 805.200 ;
        RECT 643.950 803.100 646.050 805.200 ;
        RECT 638.400 801.000 639.600 802.800 ;
        RECT 644.400 802.050 645.600 802.800 ;
        RECT 637.950 796.950 640.050 801.000 ;
        RECT 643.950 799.950 646.050 802.050 ;
        RECT 628.950 790.950 631.050 793.050 ;
        RECT 634.950 790.950 637.050 793.050 ;
        RECT 625.950 781.950 628.050 784.050 ;
        RECT 635.400 763.050 636.450 790.950 ;
        RECT 646.950 787.950 649.050 790.050 ;
        RECT 643.950 778.950 646.050 781.050 ;
        RECT 620.400 760.350 621.600 762.600 ;
        RECT 631.950 760.950 634.050 763.050 ;
        RECT 634.950 760.950 637.050 763.050 ;
        RECT 637.950 760.950 640.050 763.050 ;
        RECT 644.400 762.600 645.450 778.950 ;
        RECT 647.400 778.050 648.450 787.950 ;
        RECT 646.950 775.950 649.050 778.050 ;
        RECT 650.400 775.050 651.450 805.950 ;
        RECT 656.400 805.500 657.600 806.250 ;
        RECT 662.400 805.500 663.600 807.600 ;
        RECT 673.950 806.100 676.050 808.200 ;
        RECT 682.950 806.250 685.050 808.350 ;
        RECT 689.400 807.600 690.450 817.950 ;
        RECT 799.950 814.950 802.050 817.050 ;
        RECT 674.400 805.350 675.600 806.100 ;
        RECT 655.950 803.100 658.050 805.200 ;
        RECT 658.950 803.100 661.050 805.200 ;
        RECT 661.950 803.100 664.050 805.200 ;
        RECT 664.950 803.100 667.050 805.200 ;
        RECT 673.950 802.950 676.050 805.050 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 655.950 801.450 658.050 802.050 ;
        RECT 659.400 801.450 660.600 802.800 ;
        RECT 655.950 800.400 660.600 801.450 ;
        RECT 665.400 801.000 666.600 802.800 ;
        RECT 655.950 799.950 658.050 800.400 ;
        RECT 649.950 772.950 652.050 775.050 ;
        RECT 649.950 766.950 652.050 769.050 ;
        RECT 601.950 757.800 604.050 759.900 ;
        RECT 604.950 757.800 607.050 759.900 ;
        RECT 607.950 757.800 610.050 759.900 ;
        RECT 616.950 757.950 619.050 760.050 ;
        RECT 619.950 757.950 622.050 760.050 ;
        RECT 622.950 757.950 625.050 760.050 ;
        RECT 605.400 755.400 606.600 757.500 ;
        RECT 598.950 751.950 601.050 754.050 ;
        RECT 595.950 730.950 598.050 733.050 ;
        RECT 599.400 729.600 600.450 751.950 ;
        RECT 605.400 748.050 606.450 755.400 ;
        RECT 610.800 754.950 612.900 757.050 ;
        RECT 617.400 755.400 618.600 757.650 ;
        RECT 623.400 755.400 624.600 757.650 ;
        RECT 611.400 750.450 612.450 754.950 ;
        RECT 617.400 751.050 618.450 755.400 ;
        RECT 608.400 749.400 612.450 750.450 ;
        RECT 604.950 745.950 607.050 748.050 ;
        RECT 608.400 739.050 609.450 749.400 ;
        RECT 616.950 748.950 619.050 751.050 ;
        RECT 623.400 748.050 624.450 755.400 ;
        RECT 625.950 754.950 628.050 757.050 ;
        RECT 632.400 756.450 633.450 760.950 ;
        RECT 638.400 760.200 639.600 760.950 ;
        RECT 644.400 760.200 645.600 762.600 ;
        RECT 637.950 757.800 640.050 759.900 ;
        RECT 640.950 757.800 643.050 759.900 ;
        RECT 643.950 757.800 646.050 759.900 ;
        RECT 641.400 756.750 642.600 757.500 ;
        RECT 650.400 756.900 651.450 766.950 ;
        RECT 656.400 763.200 657.450 799.950 ;
        RECT 664.950 796.950 667.050 801.000 ;
        RECT 670.950 799.950 673.050 802.050 ;
        RECT 677.400 801.450 678.600 802.650 ;
        RECT 683.400 801.450 684.450 806.250 ;
        RECT 689.400 805.350 690.600 807.600 ;
        RECT 706.950 806.250 709.050 808.350 ;
        RECT 712.950 806.250 715.050 808.350 ;
        RECT 707.400 805.500 708.600 806.250 ;
        RECT 713.400 805.500 714.600 806.250 ;
        RECT 718.950 805.950 721.050 808.050 ;
        RECT 724.950 806.100 727.050 808.200 ;
        RECT 730.950 806.100 733.050 808.200 ;
        RECT 739.950 806.250 742.050 808.350 ;
        RECT 748.950 806.250 751.050 808.350 ;
        RECT 754.950 807.000 757.050 811.050 ;
        RECT 688.950 802.950 691.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 703.950 803.100 706.050 805.200 ;
        RECT 706.950 803.100 709.050 805.200 ;
        RECT 709.950 803.100 712.050 805.200 ;
        RECT 712.950 803.100 715.050 805.200 ;
        RECT 692.400 801.900 693.600 802.650 ;
        RECT 704.400 802.050 705.600 802.800 ;
        RECT 710.400 802.050 711.600 802.800 ;
        RECT 677.400 800.400 684.450 801.450 ;
        RECT 671.400 784.050 672.450 799.950 ;
        RECT 673.950 796.950 679.050 799.050 ;
        RECT 691.950 796.950 694.050 801.900 ;
        RECT 703.950 799.950 706.050 802.050 ;
        RECT 709.950 799.950 712.050 802.050 ;
        RECT 710.400 796.050 711.450 799.950 ;
        RECT 709.950 795.450 712.050 796.050 ;
        RECT 707.400 794.400 712.050 795.450 ;
        RECT 700.950 784.950 703.050 787.050 ;
        RECT 661.950 781.950 664.050 784.050 ;
        RECT 670.950 781.950 673.050 784.050 ;
        RECT 655.950 761.100 658.050 763.200 ;
        RECT 662.400 762.600 663.450 781.950 ;
        RECT 701.400 781.050 702.450 784.950 ;
        RECT 682.950 778.950 685.050 781.050 ;
        RECT 700.950 778.950 703.050 781.050 ;
        RECT 656.400 760.350 657.600 761.100 ;
        RECT 662.400 760.350 663.600 762.600 ;
        RECT 676.950 761.100 679.050 763.200 ;
        RECT 683.400 763.050 684.450 778.950 ;
        RECT 688.950 766.950 691.050 769.050 ;
        RECT 685.950 763.950 688.050 766.050 ;
        RECT 677.400 760.350 678.600 761.100 ;
        RECT 682.950 760.950 685.050 763.050 ;
        RECT 655.950 757.950 658.050 760.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 661.950 757.950 664.050 760.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 673.950 757.950 676.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 679.950 757.950 682.050 760.050 ;
        RECT 632.400 755.400 636.450 756.450 ;
        RECT 622.950 745.950 625.050 748.050 ;
        RECT 607.950 736.950 610.050 739.050 ;
        RECT 610.950 733.950 613.050 736.050 ;
        RECT 611.400 729.600 612.450 733.950 ;
        RECT 599.400 727.500 600.600 729.600 ;
        RECT 611.400 727.350 612.600 729.600 ;
        RECT 616.950 728.100 619.050 730.200 ;
        RECT 623.400 729.450 624.450 745.950 ;
        RECT 626.400 745.050 627.450 754.950 ;
        RECT 631.950 751.950 634.050 754.050 ;
        RECT 625.950 742.950 628.050 745.050 ;
        RECT 632.400 729.600 633.450 751.950 ;
        RECT 635.400 739.050 636.450 755.400 ;
        RECT 640.950 754.650 643.050 756.750 ;
        RECT 649.950 754.800 652.050 756.900 ;
        RECT 659.400 755.400 660.600 757.650 ;
        RECT 665.400 756.900 666.600 757.650 ;
        RECT 637.950 751.950 640.050 754.050 ;
        RECT 634.950 736.950 637.050 739.050 ;
        RECT 638.400 729.600 639.450 751.950 ;
        RECT 659.400 748.050 660.450 755.400 ;
        RECT 664.950 754.800 667.050 756.900 ;
        RECT 674.400 755.400 675.600 757.650 ;
        RECT 680.400 755.400 681.600 757.650 ;
        RECT 661.950 748.950 664.050 751.050 ;
        RECT 658.950 745.950 661.050 748.050 ;
        RECT 662.400 735.600 663.450 748.950 ;
        RECT 674.400 748.050 675.450 755.400 ;
        RECT 680.400 751.050 681.450 755.400 ;
        RECT 686.400 751.050 687.450 763.950 ;
        RECT 679.950 748.950 682.050 751.050 ;
        RECT 685.950 748.950 688.050 751.050 ;
        RECT 673.950 745.950 676.050 748.050 ;
        RECT 689.400 739.050 690.450 766.950 ;
        RECT 694.950 762.000 697.050 766.050 ;
        RECT 701.400 762.600 702.450 778.950 ;
        RECT 707.400 763.050 708.450 794.400 ;
        RECT 709.950 793.950 712.050 794.400 ;
        RECT 709.950 784.950 712.050 787.050 ;
        RECT 710.400 766.050 711.450 784.950 ;
        RECT 719.400 775.050 720.450 805.950 ;
        RECT 725.400 805.350 726.600 806.100 ;
        RECT 731.400 805.350 732.600 806.100 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 727.950 802.950 730.050 805.050 ;
        RECT 730.950 802.950 733.050 805.050 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 728.400 800.400 729.600 802.650 ;
        RECT 734.400 800.400 735.600 802.650 ;
        RECT 728.400 781.050 729.450 800.400 ;
        RECT 734.400 793.050 735.450 800.400 ;
        RECT 730.950 790.950 733.050 793.050 ;
        RECT 733.950 790.950 736.050 793.050 ;
        RECT 727.950 778.950 730.050 781.050 ;
        RECT 712.950 772.950 715.050 775.050 ;
        RECT 718.950 772.950 721.050 775.050 ;
        RECT 709.950 763.950 712.050 766.050 ;
        RECT 713.400 763.050 714.450 772.950 ;
        RECT 718.950 766.950 721.050 769.050 ;
        RECT 695.400 760.350 696.600 762.000 ;
        RECT 701.400 760.350 702.600 762.600 ;
        RECT 706.950 760.950 709.050 763.050 ;
        RECT 712.950 760.950 715.050 763.050 ;
        RECT 719.400 762.600 720.450 766.950 ;
        RECT 731.400 763.050 732.450 790.950 ;
        RECT 736.950 772.950 739.050 775.050 ;
        RECT 727.950 762.600 732.450 763.050 ;
        RECT 737.400 762.600 738.450 772.950 ;
        RECT 740.400 763.050 741.450 806.250 ;
        RECT 749.400 805.500 750.600 806.250 ;
        RECT 755.400 805.500 756.600 807.000 ;
        RECT 769.950 806.250 772.050 808.350 ;
        RECT 787.950 806.250 790.050 808.350 ;
        RECT 793.950 806.250 796.050 808.350 ;
        RECT 770.400 805.500 771.600 806.250 ;
        RECT 788.400 805.500 789.600 806.250 ;
        RECT 794.400 805.500 795.600 806.250 ;
        RECT 745.950 803.100 748.050 805.200 ;
        RECT 748.950 803.100 751.050 805.200 ;
        RECT 751.950 803.100 754.050 805.200 ;
        RECT 754.950 803.100 757.050 805.200 ;
        RECT 766.950 803.100 769.050 805.200 ;
        RECT 769.950 803.100 772.050 805.200 ;
        RECT 772.950 803.100 775.050 805.200 ;
        RECT 784.950 803.100 787.050 805.200 ;
        RECT 787.950 803.100 790.050 805.200 ;
        RECT 790.950 803.100 793.050 805.200 ;
        RECT 793.950 803.100 796.050 805.200 ;
        RECT 746.400 800.400 747.600 802.800 ;
        RECT 752.400 801.000 753.600 802.800 ;
        RECT 742.950 796.950 745.050 799.050 ;
        RECT 719.400 760.350 720.600 762.600 ;
        RECT 727.950 760.950 732.600 762.600 ;
        RECT 731.400 760.200 732.600 760.950 ;
        RECT 737.400 760.200 738.600 762.600 ;
        RECT 739.950 760.950 742.050 763.050 ;
        RECT 694.950 757.950 697.050 760.050 ;
        RECT 697.950 757.950 700.050 760.050 ;
        RECT 700.950 757.950 703.050 760.050 ;
        RECT 703.950 757.950 706.050 760.050 ;
        RECT 715.950 757.950 718.050 760.050 ;
        RECT 718.950 757.950 721.050 760.050 ;
        RECT 721.950 757.950 724.050 760.050 ;
        RECT 730.950 757.800 733.050 759.900 ;
        RECT 733.950 757.800 736.050 759.900 ;
        RECT 736.950 757.800 739.050 759.900 ;
        RECT 691.950 754.950 694.050 757.050 ;
        RECT 698.400 755.400 699.600 757.650 ;
        RECT 704.400 756.900 705.600 757.650 ;
        RECT 716.400 756.900 717.600 757.650 ;
        RECT 688.950 736.950 691.050 739.050 ;
        RECT 658.500 732.300 660.600 734.400 ;
        RECT 662.400 732.900 663.600 735.600 ;
        RECT 623.400 728.400 627.450 729.450 ;
        RECT 617.400 727.350 618.600 728.100 ;
        RECT 595.950 725.100 598.050 727.200 ;
        RECT 598.950 725.100 601.050 727.200 ;
        RECT 601.950 725.100 604.050 727.200 ;
        RECT 610.950 724.950 613.050 727.050 ;
        RECT 613.950 724.950 616.050 727.050 ;
        RECT 616.950 724.950 619.050 727.050 ;
        RECT 619.950 724.950 622.050 727.050 ;
        RECT 596.400 724.050 597.600 724.800 ;
        RECT 602.400 724.050 603.600 724.800 ;
        RECT 589.950 721.950 592.050 724.050 ;
        RECT 595.950 721.950 598.050 724.050 ;
        RECT 601.950 723.450 604.050 724.050 ;
        RECT 601.950 722.400 606.450 723.450 ;
        RECT 601.950 721.950 604.050 722.400 ;
        RECT 586.950 709.950 589.050 712.050 ;
        RECT 590.400 709.050 591.450 721.950 ;
        RECT 601.950 715.950 604.050 718.050 ;
        RECT 589.950 706.950 592.050 709.050 ;
        RECT 583.950 700.950 586.050 703.050 ;
        RECT 577.950 694.950 580.050 697.050 ;
        RECT 566.400 683.400 570.450 684.450 ;
        RECT 571.950 684.000 574.050 688.050 ;
        RECT 556.950 679.950 559.050 682.050 ;
        RECT 559.950 679.950 562.050 682.050 ;
        RECT 536.400 673.050 537.450 676.950 ;
        RECT 541.950 676.650 544.050 678.750 ;
        RECT 550.950 676.950 553.050 679.050 ;
        RECT 557.400 678.900 558.600 679.650 ;
        RECT 556.950 676.050 559.050 678.900 ;
        RECT 566.400 678.750 567.450 683.400 ;
        RECT 572.400 682.200 573.600 684.000 ;
        RECT 571.950 679.800 574.050 681.900 ;
        RECT 574.950 679.800 577.050 681.900 ;
        RECT 575.400 678.750 576.600 679.500 ;
        RECT 565.950 676.650 568.050 678.750 ;
        RECT 574.950 678.450 577.050 678.750 ;
        RECT 574.950 677.400 579.450 678.450 ;
        RECT 574.950 676.650 577.050 677.400 ;
        RECT 547.950 673.950 550.050 676.050 ;
        RECT 556.950 673.950 562.050 676.050 ;
        RECT 571.950 673.950 574.050 676.050 ;
        RECT 535.950 670.950 538.050 673.050 ;
        RECT 526.950 667.950 529.050 670.050 ;
        RECT 548.400 667.050 549.450 673.950 ;
        RECT 550.950 670.950 553.050 673.050 ;
        RECT 538.950 664.950 541.050 667.050 ;
        RECT 547.950 664.950 550.050 667.050 ;
        RECT 529.950 655.950 532.050 658.050 ;
        RECT 521.400 649.500 522.600 651.600 ;
        RECT 517.950 647.100 520.050 649.200 ;
        RECT 520.950 647.100 523.050 649.200 ;
        RECT 523.950 647.100 526.050 649.200 ;
        RECT 493.950 640.950 496.050 643.050 ;
        RECT 481.800 634.950 483.900 637.050 ;
        RECT 475.950 616.950 478.050 619.050 ;
        RECT 487.950 616.950 490.050 619.050 ;
        RECT 472.950 604.950 475.050 607.050 ;
        RECT 476.400 606.600 477.450 616.950 ;
        RECT 476.400 604.200 477.600 606.600 ;
        RECT 481.950 604.950 484.050 607.050 ;
        RECT 482.400 604.200 483.600 604.950 ;
        RECT 475.950 601.800 478.050 603.900 ;
        RECT 478.950 601.800 481.050 603.900 ;
        RECT 481.950 601.800 484.050 603.900 ;
        RECT 464.400 589.050 465.450 599.400 ;
        RECT 469.950 598.950 472.050 601.050 ;
        RECT 472.950 598.950 475.050 601.050 ;
        RECT 479.400 600.750 480.600 601.500 ;
        RECT 469.950 592.950 472.050 595.050 ;
        RECT 463.950 586.950 466.050 589.050 ;
        RECT 466.950 583.950 469.050 586.050 ;
        RECT 451.950 582.450 454.050 583.050 ;
        RECT 451.950 581.400 456.450 582.450 ;
        RECT 451.950 580.950 454.050 581.400 ;
        RECT 439.950 578.400 442.050 580.500 ;
        RECT 425.400 571.350 426.600 572.100 ;
        RECT 431.400 571.350 432.600 573.600 ;
        RECT 421.950 568.950 424.050 571.050 ;
        RECT 424.950 568.950 427.050 571.050 ;
        RECT 427.950 568.950 430.050 571.050 ;
        RECT 430.950 568.950 433.050 571.050 ;
        RECT 436.950 568.950 439.050 571.050 ;
        RECT 422.400 566.400 423.600 568.650 ;
        RECT 428.400 566.400 429.600 568.650 ;
        RECT 437.400 567.450 438.600 568.650 ;
        RECT 434.400 566.400 438.600 567.450 ;
        RECT 415.950 559.950 418.050 562.050 ;
        RECT 422.400 556.050 423.450 566.400 ;
        RECT 421.950 553.950 424.050 556.050 ;
        RECT 412.950 550.950 415.050 553.050 ;
        RECT 409.950 549.450 414.000 550.050 ;
        RECT 409.950 547.950 414.450 549.450 ;
        RECT 406.950 544.950 409.050 547.050 ;
        RECT 403.950 535.950 406.050 538.050 ;
        RECT 398.400 526.200 399.600 528.600 ;
        RECT 400.950 526.950 403.050 529.050 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 376.950 523.950 379.050 526.050 ;
        RECT 379.950 523.950 382.050 526.050 ;
        RECT 382.950 523.950 385.050 526.050 ;
        RECT 391.950 523.800 394.050 525.900 ;
        RECT 394.950 523.800 397.050 525.900 ;
        RECT 397.950 523.800 400.050 525.900 ;
        RECT 358.950 520.650 361.050 522.750 ;
        RECT 364.950 520.950 367.050 523.050 ;
        RECT 367.950 520.950 370.050 523.050 ;
        RECT 377.400 522.900 378.600 523.650 ;
        RECT 383.400 522.900 384.600 523.650 ;
        RECT 355.950 514.950 358.050 517.050 ;
        RECT 349.950 502.950 352.050 505.050 ;
        RECT 352.950 499.950 355.050 502.050 ;
        RECT 353.400 496.050 354.450 499.950 ;
        RECT 332.400 493.350 333.600 494.100 ;
        RECT 322.950 490.950 325.050 493.050 ;
        RECT 325.950 490.950 328.050 493.050 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 331.950 490.950 334.050 493.050 ;
        RECT 319.950 487.950 322.050 490.050 ;
        RECT 323.400 488.400 324.600 490.650 ;
        RECT 329.400 488.400 330.600 490.650 ;
        RECT 320.400 484.050 321.450 487.950 ;
        RECT 316.950 481.950 319.050 484.050 ;
        RECT 319.950 481.950 322.050 484.050 ;
        RECT 323.400 481.050 324.450 488.400 ;
        RECT 329.400 486.450 330.450 488.400 ;
        RECT 334.950 486.450 337.050 490.050 ;
        RECT 329.400 486.000 337.050 486.450 ;
        RECT 329.400 485.400 336.450 486.000 ;
        RECT 331.950 481.950 334.050 484.050 ;
        RECT 316.800 478.800 318.900 480.900 ;
        RECT 319.950 478.800 322.050 480.900 ;
        RECT 322.950 478.950 325.050 481.050 ;
        RECT 317.400 475.050 318.450 478.800 ;
        RECT 305.400 473.400 312.450 474.450 ;
        RECT 298.950 457.950 301.050 460.050 ;
        RECT 286.950 451.950 289.050 454.050 ;
        RECT 283.950 448.950 286.050 451.050 ;
        RECT 286.950 448.800 289.050 450.900 ;
        RECT 292.950 448.950 295.050 451.050 ;
        RECT 287.400 448.200 288.600 448.800 ;
        RECT 293.400 448.200 294.600 448.950 ;
        RECT 286.950 445.800 289.050 447.900 ;
        RECT 289.950 445.800 292.050 447.900 ;
        RECT 292.950 445.800 295.050 447.900 ;
        RECT 283.950 442.950 286.050 445.050 ;
        RECT 290.400 443.400 291.600 445.500 ;
        RECT 280.950 427.950 283.050 430.050 ;
        RECT 280.950 421.950 283.050 424.050 ;
        RECT 265.950 416.100 268.050 418.200 ;
        RECT 271.950 416.100 274.050 418.200 ;
        RECT 281.400 417.600 282.450 421.950 ;
        RECT 284.400 421.050 285.450 442.950 ;
        RECT 290.400 423.450 291.450 443.400 ;
        RECT 299.400 441.450 300.450 457.950 ;
        RECT 305.400 451.200 306.450 473.400 ;
        RECT 313.800 472.950 315.900 475.050 ;
        RECT 316.950 472.950 319.050 475.050 ;
        RECT 307.800 457.950 309.900 460.050 ;
        RECT 304.800 449.100 306.900 451.200 ;
        RECT 308.400 451.050 309.450 457.950 ;
        RECT 320.400 454.050 321.450 478.800 ;
        RECT 319.950 451.950 322.050 454.050 ;
        RECT 305.400 448.350 306.600 449.100 ;
        RECT 307.950 448.950 310.050 451.050 ;
        RECT 322.950 449.100 325.050 451.200 ;
        RECT 328.950 450.000 331.050 454.050 ;
        RECT 332.400 451.050 333.450 481.950 ;
        RECT 338.400 481.050 339.450 494.400 ;
        RECT 347.400 493.500 348.600 495.600 ;
        RECT 352.950 493.950 355.050 496.050 ;
        RECT 343.950 491.100 346.050 493.200 ;
        RECT 346.950 491.100 349.050 493.200 ;
        RECT 349.950 491.100 352.050 493.200 ;
        RECT 344.400 490.050 345.600 490.800 ;
        RECT 350.400 490.050 351.600 490.800 ;
        RECT 356.400 490.050 357.450 514.950 ;
        RECT 365.400 496.350 366.450 520.950 ;
        RECT 376.950 520.800 379.050 522.900 ;
        RECT 382.950 520.800 385.050 522.900 ;
        RECT 395.400 522.750 396.600 523.500 ;
        RECT 394.950 520.650 397.050 522.750 ;
        RECT 404.400 517.050 405.450 535.950 ;
        RECT 408.000 531.900 411.000 532.050 ;
        RECT 406.950 529.950 412.050 531.900 ;
        RECT 406.950 529.800 409.050 529.950 ;
        RECT 409.950 529.800 412.050 529.950 ;
        RECT 413.400 528.600 414.450 547.950 ;
        RECT 428.400 541.050 429.450 566.400 ;
        RECT 434.400 552.450 435.450 566.400 ;
        RECT 440.700 558.600 441.900 578.400 ;
        RECT 445.950 568.950 448.050 571.050 ;
        RECT 446.400 567.900 447.600 568.650 ;
        RECT 445.950 565.800 448.050 567.900 ;
        RECT 455.400 562.050 456.450 581.400 ;
        RECT 460.950 578.400 463.050 580.500 ;
        RECT 460.950 563.400 462.150 578.400 ;
        RECT 464.400 573.450 465.600 573.600 ;
        RECT 467.400 573.450 468.450 583.950 ;
        RECT 464.400 572.400 468.450 573.450 ;
        RECT 464.400 571.350 465.600 572.400 ;
        RECT 463.950 568.950 466.050 571.050 ;
        RECT 445.950 559.950 448.050 562.050 ;
        RECT 454.950 559.950 457.050 562.050 ;
        RECT 460.950 561.300 463.050 563.400 ;
        RECT 439.950 556.500 442.050 558.600 ;
        RECT 434.400 551.400 438.450 552.450 ;
        RECT 427.950 538.950 430.050 541.050 ;
        RECT 428.400 535.050 429.450 538.950 ;
        RECT 421.950 529.950 424.050 535.050 ;
        RECT 427.950 532.950 430.050 535.050 ;
        RECT 430.950 532.950 433.050 538.050 ;
        RECT 437.400 532.050 438.450 551.400 ;
        RECT 446.400 550.050 447.450 559.950 ;
        RECT 460.950 557.700 462.150 561.300 ;
        RECT 470.400 558.450 471.450 592.950 ;
        RECT 473.400 592.050 474.450 598.950 ;
        RECT 478.950 598.650 481.050 600.750 ;
        RECT 472.950 589.950 475.050 592.050 ;
        RECT 472.950 586.800 475.050 588.900 ;
        RECT 473.400 561.450 474.450 586.800 ;
        RECT 481.950 572.250 484.050 574.350 ;
        RECT 488.400 573.450 489.450 616.950 ;
        RECT 494.400 607.050 495.450 640.950 ;
        RECT 500.400 628.050 501.450 644.400 ;
        RECT 506.400 640.050 507.450 644.400 ;
        RECT 511.950 643.950 514.050 646.050 ;
        RECT 518.400 645.450 519.600 646.800 ;
        RECT 515.400 644.400 519.600 645.450 ;
        RECT 524.400 644.400 525.600 646.800 ;
        RECT 508.950 640.950 511.050 643.050 ;
        RECT 505.950 637.950 508.050 640.050 ;
        RECT 499.950 625.950 502.050 628.050 ;
        RECT 500.400 610.050 501.450 625.950 ;
        RECT 509.400 613.050 510.450 640.950 ;
        RECT 515.400 634.050 516.450 644.400 ;
        RECT 524.400 640.050 525.450 644.400 ;
        RECT 526.950 640.950 529.050 646.050 ;
        RECT 523.950 639.450 526.050 640.050 ;
        RECT 523.950 638.400 528.450 639.450 ;
        RECT 523.950 637.950 526.050 638.400 ;
        RECT 514.950 631.950 517.050 634.050 ;
        RECT 523.950 631.950 526.050 634.050 ;
        RECT 517.950 628.950 520.050 631.050 ;
        RECT 508.950 610.950 511.050 613.050 ;
        RECT 511.950 610.950 514.050 613.050 ;
        RECT 499.950 607.950 502.050 610.050 ;
        RECT 505.950 607.950 508.050 610.050 ;
        RECT 493.950 604.950 496.050 607.050 ;
        RECT 494.400 604.200 495.600 604.950 ;
        RECT 499.950 604.800 502.050 606.900 ;
        RECT 500.400 604.200 501.600 604.800 ;
        RECT 493.950 601.800 496.050 603.900 ;
        RECT 496.950 601.800 499.050 603.900 ;
        RECT 499.950 601.800 502.050 603.900 ;
        RECT 490.950 598.950 493.050 601.050 ;
        RECT 497.400 599.400 498.600 601.500 ;
        RECT 491.400 595.050 492.450 598.950 ;
        RECT 497.400 595.050 498.450 599.400 ;
        RECT 502.950 598.950 505.050 601.050 ;
        RECT 490.950 592.950 493.050 595.050 ;
        RECT 496.950 592.950 499.050 595.050 ;
        RECT 503.400 576.450 504.450 598.950 ;
        RECT 506.400 580.050 507.450 607.950 ;
        RECT 512.400 606.600 513.450 610.950 ;
        RECT 518.400 606.600 519.450 628.950 ;
        RECT 524.400 607.050 525.450 631.950 ;
        RECT 527.400 622.050 528.450 638.400 ;
        RECT 530.400 631.050 531.450 655.950 ;
        RECT 539.400 652.050 540.450 664.950 ;
        RECT 538.950 649.950 541.050 652.050 ;
        RECT 535.950 647.100 538.050 649.200 ;
        RECT 541.950 647.100 544.050 649.200 ;
        RECT 544.950 647.100 547.050 649.200 ;
        RECT 536.400 646.050 537.600 646.800 ;
        RECT 532.950 643.950 535.050 646.050 ;
        RECT 535.950 643.950 538.050 646.050 ;
        RECT 545.400 644.400 546.600 646.800 ;
        RECT 529.950 628.950 532.050 631.050 ;
        RECT 529.950 625.800 532.050 627.900 ;
        RECT 526.950 619.950 529.050 622.050 ;
        RECT 530.400 610.050 531.450 625.800 ;
        RECT 533.400 619.050 534.450 643.950 ;
        RECT 536.400 642.450 537.450 643.950 ;
        RECT 541.950 642.450 544.050 643.050 ;
        RECT 536.400 641.400 544.050 642.450 ;
        RECT 541.950 640.950 544.050 641.400 ;
        RECT 538.950 637.950 541.050 640.050 ;
        RECT 539.400 619.050 540.450 637.950 ;
        RECT 542.400 628.050 543.450 640.950 ;
        RECT 541.950 625.950 544.050 628.050 ;
        RECT 545.400 622.050 546.450 644.400 ;
        RECT 551.400 625.050 552.450 670.950 ;
        RECT 572.400 652.050 573.450 673.950 ;
        RECT 574.950 661.950 577.050 664.050 ;
        RECT 571.950 649.950 574.050 652.050 ;
        RECT 556.950 647.100 559.050 649.200 ;
        RECT 559.950 647.100 562.050 649.200 ;
        RECT 562.950 647.100 565.050 649.200 ;
        RECT 565.950 647.100 568.050 649.200 ;
        RECT 568.950 647.100 571.050 649.200 ;
        RECT 557.400 645.000 558.600 646.800 ;
        RECT 556.950 640.950 559.050 645.000 ;
        RECT 563.400 644.400 564.600 646.800 ;
        RECT 569.400 646.050 570.600 646.800 ;
        RECT 559.950 637.950 562.050 640.050 ;
        RECT 553.950 634.950 556.050 637.050 ;
        RECT 550.950 622.950 553.050 625.050 ;
        RECT 544.950 619.950 547.050 622.050 ;
        RECT 532.950 616.950 535.050 619.050 ;
        RECT 538.950 616.950 541.050 619.050 ;
        RECT 533.400 613.050 534.450 616.950 ;
        RECT 544.950 616.800 547.050 618.900 ;
        RECT 535.950 613.950 538.050 616.050 ;
        RECT 532.950 610.950 535.050 613.050 ;
        RECT 529.950 607.950 532.050 610.050 ;
        RECT 536.400 609.450 537.450 613.950 ;
        RECT 545.400 613.050 546.450 616.800 ;
        RECT 544.950 610.950 547.050 613.050 ;
        RECT 533.400 608.400 537.450 609.450 ;
        RECT 512.400 604.350 513.600 606.600 ;
        RECT 518.400 604.350 519.600 606.600 ;
        RECT 523.950 604.950 526.050 607.050 ;
        RECT 533.400 606.600 534.450 608.400 ;
        RECT 533.400 604.350 534.600 606.600 ;
        RECT 538.950 606.000 541.050 610.050 ;
        RECT 544.950 607.800 547.050 609.900 ;
        RECT 539.400 604.350 540.600 606.000 ;
        RECT 511.950 601.950 514.050 604.050 ;
        RECT 514.950 601.950 517.050 604.050 ;
        RECT 517.950 601.950 520.050 604.050 ;
        RECT 520.950 601.950 523.050 604.050 ;
        RECT 529.950 601.950 532.050 604.050 ;
        RECT 532.950 601.950 535.050 604.050 ;
        RECT 535.950 601.950 538.050 604.050 ;
        RECT 538.950 601.950 541.050 604.050 ;
        RECT 508.950 598.950 511.050 601.050 ;
        RECT 515.400 600.900 516.600 601.650 ;
        RECT 509.400 589.050 510.450 598.950 ;
        RECT 514.950 598.800 517.050 600.900 ;
        RECT 521.400 599.400 522.600 601.650 ;
        RECT 530.400 599.400 531.600 601.650 ;
        RECT 536.400 599.400 537.600 601.650 ;
        RECT 521.400 592.050 522.450 599.400 ;
        RECT 511.800 589.950 513.900 592.050 ;
        RECT 514.950 589.950 517.050 592.050 ;
        RECT 520.950 589.950 523.050 592.050 ;
        RECT 526.950 589.950 529.050 592.050 ;
        RECT 508.950 586.950 511.050 589.050 ;
        RECT 505.950 577.950 508.050 580.050 ;
        RECT 500.400 575.400 504.450 576.450 ;
        RECT 500.400 573.600 501.450 575.400 ;
        RECT 488.400 572.400 492.450 573.450 ;
        RECT 482.400 571.500 483.600 572.250 ;
        RECT 478.950 569.100 481.050 571.200 ;
        RECT 481.950 569.100 484.050 571.200 ;
        RECT 484.950 569.100 487.050 571.200 ;
        RECT 479.400 566.400 480.600 568.800 ;
        RECT 485.400 566.400 486.600 568.800 ;
        RECT 473.400 560.400 477.450 561.450 ;
        RECT 460.950 555.600 463.050 557.700 ;
        RECT 470.400 557.400 474.450 558.450 ;
        RECT 445.950 547.950 448.050 550.050 ;
        RECT 457.950 547.950 460.050 550.050 ;
        RECT 448.950 536.400 451.050 538.500 ;
        RECT 458.400 538.050 459.450 547.950 ;
        RECT 473.400 544.050 474.450 557.400 ;
        RECT 476.400 550.050 477.450 560.400 ;
        RECT 475.950 547.950 478.050 550.050 ;
        RECT 460.950 541.950 463.050 544.050 ;
        RECT 472.950 541.950 475.050 544.050 ;
        RECT 436.950 529.950 439.050 532.050 ;
        RECT 413.400 526.350 414.600 528.600 ;
        RECT 418.950 527.100 421.050 529.200 ;
        RECT 419.400 526.350 420.600 527.100 ;
        RECT 424.950 526.950 427.050 529.050 ;
        RECT 430.950 526.950 433.050 529.050 ;
        RECT 445.950 528.000 448.050 532.050 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 415.950 523.950 418.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 406.950 520.950 409.050 523.050 ;
        RECT 410.400 522.900 411.600 523.650 ;
        RECT 403.950 514.950 406.050 517.050 ;
        RECT 394.950 511.950 397.050 514.050 ;
        RECT 367.950 505.950 370.050 508.050 ;
        RECT 391.950 505.950 394.050 508.050 ;
        RECT 368.400 502.050 369.450 505.950 ;
        RECT 367.950 499.950 370.050 502.050 ;
        RECT 364.950 494.250 367.050 496.350 ;
        RECT 382.950 494.250 385.050 496.350 ;
        RECT 365.400 493.500 366.600 494.250 ;
        RECT 383.400 493.500 384.600 494.250 ;
        RECT 361.950 491.100 364.050 493.200 ;
        RECT 364.950 491.100 367.050 493.200 ;
        RECT 370.950 491.100 373.050 493.200 ;
        RECT 379.950 491.100 382.050 493.200 ;
        RECT 382.950 491.100 385.050 493.200 ;
        RECT 385.950 491.100 388.050 493.200 ;
        RECT 343.950 487.950 346.050 490.050 ;
        RECT 349.950 487.950 352.050 490.050 ;
        RECT 355.950 487.950 358.050 490.050 ;
        RECT 358.950 487.950 361.050 490.050 ;
        RECT 362.400 488.400 363.600 490.800 ;
        RECT 371.400 490.050 372.600 490.800 ;
        RECT 380.400 490.050 381.600 490.800 ;
        RECT 340.950 481.950 343.050 484.050 ;
        RECT 337.950 478.950 340.050 481.050 ;
        RECT 341.400 478.050 342.450 481.950 ;
        RECT 339.000 477.900 342.450 478.050 ;
        RECT 337.950 476.400 342.450 477.900 ;
        RECT 337.950 475.950 342.000 476.400 ;
        RECT 337.950 475.800 340.050 475.950 ;
        RECT 359.400 475.050 360.450 487.950 ;
        RECT 362.400 484.050 363.450 488.400 ;
        RECT 370.950 487.950 373.050 490.050 ;
        RECT 379.950 487.950 382.050 490.050 ;
        RECT 386.400 489.000 387.600 490.800 ;
        RECT 385.950 484.950 388.050 489.000 ;
        RECT 388.950 487.950 391.050 490.050 ;
        RECT 361.950 481.950 364.050 484.050 ;
        RECT 385.950 478.950 388.050 481.050 ;
        RECT 340.950 472.950 343.050 475.050 ;
        RECT 358.950 472.950 361.050 475.050 ;
        RECT 334.950 451.950 337.050 454.050 ;
        RECT 323.400 448.350 324.600 449.100 ;
        RECT 329.400 448.350 330.600 450.000 ;
        RECT 331.950 448.950 334.050 451.050 ;
        RECT 304.950 445.950 307.050 448.050 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 319.950 445.950 322.050 448.050 ;
        RECT 322.950 445.950 325.050 448.050 ;
        RECT 325.950 445.950 328.050 448.050 ;
        RECT 328.950 445.950 331.050 448.050 ;
        RECT 311.400 444.450 312.600 445.650 ;
        RECT 320.400 444.900 321.600 445.650 ;
        RECT 311.400 443.400 315.450 444.450 ;
        RECT 296.400 440.400 300.450 441.450 ;
        RECT 296.400 433.050 297.450 440.400 ;
        RECT 310.950 439.950 313.050 442.050 ;
        RECT 298.950 436.950 301.050 439.050 ;
        RECT 295.950 430.950 298.050 433.050 ;
        RECT 290.400 422.400 294.450 423.450 ;
        RECT 283.950 418.950 286.050 421.050 ;
        RECT 289.950 418.950 292.050 421.050 ;
        RECT 266.400 415.350 267.600 416.100 ;
        RECT 272.400 415.350 273.600 416.100 ;
        RECT 281.400 415.350 282.600 417.600 ;
        RECT 262.950 412.950 265.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 268.950 412.950 271.050 415.050 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 280.950 412.950 283.050 415.050 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 263.400 412.050 264.600 412.650 ;
        RECT 259.950 410.400 264.600 412.050 ;
        RECT 269.400 410.400 270.600 412.650 ;
        RECT 259.950 409.950 264.000 410.400 ;
        RECT 256.950 394.950 259.050 397.050 ;
        RECT 269.400 394.050 270.450 410.400 ;
        RECT 274.950 409.950 277.050 412.050 ;
        RECT 284.400 411.900 285.600 412.650 ;
        RECT 290.400 412.050 291.450 418.950 ;
        RECT 293.400 418.050 294.450 422.400 ;
        RECT 292.950 415.950 295.050 418.050 ;
        RECT 299.400 417.600 300.450 436.950 ;
        RECT 299.400 415.500 300.600 417.600 ;
        RECT 304.950 416.250 307.050 418.350 ;
        RECT 305.400 415.500 306.600 416.250 ;
        RECT 295.950 413.100 298.050 415.200 ;
        RECT 298.950 413.100 301.050 415.200 ;
        RECT 301.950 413.100 304.050 415.200 ;
        RECT 304.950 413.100 307.050 415.200 ;
        RECT 296.400 412.050 297.600 412.800 ;
        RECT 268.950 391.950 271.050 394.050 ;
        RECT 275.400 382.050 276.450 409.950 ;
        RECT 283.950 409.800 286.050 411.900 ;
        RECT 289.950 409.950 292.050 412.050 ;
        RECT 292.950 409.950 295.050 412.050 ;
        RECT 295.950 409.950 298.050 412.050 ;
        RECT 302.400 411.000 303.600 412.800 ;
        RECT 290.400 403.050 291.450 409.950 ;
        RECT 289.950 400.950 292.050 403.050 ;
        RECT 169.950 376.950 172.050 379.050 ;
        RECT 178.950 376.950 181.050 379.050 ;
        RECT 193.950 376.950 196.050 379.050 ;
        RECT 166.950 373.950 169.050 376.050 ;
        RECT 164.400 369.900 165.600 372.600 ;
        RECT 163.950 367.800 166.050 369.900 ;
        RECT 145.950 358.950 148.050 361.050 ;
        RECT 155.400 360.900 156.600 362.100 ;
        RECT 161.250 361.500 163.350 363.600 ;
        RECT 91.950 355.950 94.050 358.050 ;
        RECT 109.950 355.950 112.050 358.050 ;
        RECT 124.950 355.950 127.050 358.050 ;
        RECT 142.950 355.950 145.050 358.050 ;
        RECT 88.950 346.950 91.050 349.050 ;
        RECT 92.400 339.600 93.450 355.950 ;
        RECT 100.950 346.950 103.050 349.050 ;
        RECT 101.400 340.050 102.450 346.950 ;
        RECT 103.950 343.950 106.050 346.050 ;
        RECT 127.950 343.950 130.050 346.050 ;
        RECT 139.950 343.950 142.050 346.050 ;
        RECT 92.400 337.350 93.600 339.600 ;
        RECT 100.950 337.950 103.050 340.050 ;
        RECT 104.400 339.600 105.450 343.950 ;
        RECT 104.400 337.500 105.600 339.600 ;
        RECT 109.950 339.000 112.050 343.050 ;
        RECT 110.400 337.500 111.600 339.000 ;
        RECT 115.950 338.250 118.050 340.350 ;
        RECT 128.400 339.600 129.450 343.950 ;
        RECT 116.400 337.500 117.600 338.250 ;
        RECT 128.400 337.500 129.600 339.600 ;
        RECT 136.950 338.250 139.050 340.350 ;
        RECT 88.950 334.950 91.050 337.050 ;
        RECT 91.950 334.950 94.050 337.050 ;
        RECT 103.950 335.100 106.050 337.200 ;
        RECT 106.950 335.100 109.050 337.200 ;
        RECT 109.950 335.100 112.050 337.200 ;
        RECT 112.950 335.100 115.050 337.200 ;
        RECT 115.950 335.100 118.050 337.200 ;
        RECT 124.950 335.100 127.050 337.200 ;
        RECT 127.950 335.100 130.050 337.200 ;
        RECT 130.950 335.100 133.050 337.200 ;
        RECT 89.400 333.900 90.600 334.650 ;
        RECT 88.950 331.800 91.050 333.900 ;
        RECT 100.950 331.950 103.050 334.050 ;
        RECT 107.400 332.400 108.600 334.800 ;
        RECT 113.400 333.450 114.600 334.800 ;
        RECT 125.400 334.050 126.600 334.800 ;
        RECT 115.950 333.450 118.050 334.050 ;
        RECT 113.400 333.000 118.050 333.450 ;
        RECT 112.950 332.400 118.050 333.000 ;
        RECT 82.950 322.950 85.050 325.050 ;
        RECT 67.950 307.950 70.050 310.050 ;
        RECT 79.950 307.950 82.050 310.050 ;
        RECT 70.950 303.300 73.050 305.400 ;
        RECT 70.950 299.700 72.150 303.300 ;
        RECT 76.950 301.950 79.050 304.050 ;
        RECT 70.950 297.600 73.050 299.700 ;
        RECT 64.950 293.100 67.050 295.200 ;
        RECT 65.400 286.050 66.450 293.100 ;
        RECT 64.950 283.950 67.050 286.050 ;
        RECT 70.950 282.600 72.150 297.600 ;
        RECT 77.400 295.050 78.450 301.950 ;
        RECT 80.400 300.450 81.450 307.950 ;
        RECT 85.950 302.400 88.050 304.500 ;
        RECT 80.400 299.400 84.450 300.450 ;
        RECT 83.400 295.200 84.450 299.400 ;
        RECT 76.950 292.950 79.050 295.050 ;
        RECT 82.950 293.100 85.050 295.200 ;
        RECT 83.400 292.350 84.600 293.100 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 74.400 288.900 75.600 289.650 ;
        RECT 73.950 286.800 76.050 288.900 ;
        RECT 86.700 282.600 87.900 302.400 ;
        RECT 91.950 293.100 94.050 295.200 ;
        RECT 97.950 293.100 100.050 295.200 ;
        RECT 92.400 292.350 93.600 293.100 ;
        RECT 91.950 289.950 94.050 292.050 ;
        RECT 91.950 283.950 94.050 286.050 ;
        RECT 70.950 280.500 73.050 282.600 ;
        RECT 85.950 280.500 88.050 282.600 ;
        RECT 61.950 271.950 64.050 274.050 ;
        RECT 64.950 266.400 67.050 268.500 ;
        RECT 64.950 251.400 66.150 266.400 ;
        RECT 67.950 260.100 70.050 262.200 ;
        RECT 73.950 260.100 76.050 262.200 ;
        RECT 82.950 260.250 85.050 262.350 ;
        RECT 68.400 259.350 69.600 260.100 ;
        RECT 67.950 256.950 70.050 259.050 ;
        RECT 74.400 255.450 75.450 260.100 ;
        RECT 83.400 259.500 84.600 260.250 ;
        RECT 88.950 259.950 91.050 265.050 ;
        RECT 79.950 257.100 82.050 259.200 ;
        RECT 82.950 257.100 85.050 259.200 ;
        RECT 85.950 257.100 88.050 259.200 ;
        RECT 80.400 255.450 81.600 256.800 ;
        RECT 74.400 254.400 81.600 255.450 ;
        RECT 86.400 254.400 87.600 256.800 ;
        RECT 58.950 247.950 61.050 250.050 ;
        RECT 64.950 249.300 67.050 251.400 ;
        RECT 64.950 245.700 66.150 249.300 ;
        RECT 64.950 243.600 67.050 245.700 ;
        RECT 67.950 223.950 70.050 226.050 ;
        RECT 68.400 216.600 69.450 223.950 ;
        RECT 47.400 214.200 48.600 214.950 ;
        RECT 56.400 214.200 57.600 216.600 ;
        RECT 68.400 214.350 69.600 216.600 ;
        RECT 31.950 211.950 34.050 214.050 ;
        RECT 46.950 211.800 49.050 213.900 ;
        RECT 49.950 211.800 52.050 213.900 ;
        RECT 55.950 211.800 58.050 213.900 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 50.400 210.000 51.600 211.500 ;
        RECT 49.950 205.950 52.050 210.000 ;
        RECT 65.400 209.400 66.600 211.650 ;
        RECT 71.400 210.900 72.600 211.650 ;
        RECT 77.400 211.050 78.450 254.400 ;
        RECT 86.400 247.050 87.450 254.400 ;
        RECT 85.950 244.950 88.050 247.050 ;
        RECT 85.950 215.100 88.050 217.200 ;
        RECT 86.400 214.350 87.600 215.100 ;
        RECT 82.950 211.950 85.050 214.050 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 61.950 205.950 64.050 208.050 ;
        RECT 28.950 202.500 31.050 204.600 ;
        RECT 16.950 196.950 19.050 199.050 ;
        RECT 13.950 190.950 16.050 193.050 ;
        RECT 28.950 190.950 31.050 193.050 ;
        RECT 22.950 188.400 25.050 190.500 ;
        RECT 7.950 182.100 10.050 184.200 ;
        RECT 19.950 183.000 22.050 187.050 ;
        RECT 8.400 181.350 9.600 182.100 ;
        RECT 20.400 181.350 21.600 183.000 ;
        RECT 7.950 178.950 10.050 181.050 ;
        RECT 10.950 178.950 13.050 181.050 ;
        RECT 19.950 178.950 22.050 181.050 ;
        RECT 4.950 175.950 7.050 178.050 ;
        RECT 11.400 176.400 12.600 178.650 ;
        RECT 5.400 133.050 6.450 175.950 ;
        RECT 11.400 163.050 12.450 176.400 ;
        RECT 23.850 173.400 25.050 188.400 ;
        RECT 22.950 171.300 25.050 173.400 ;
        RECT 23.850 167.700 25.050 171.300 ;
        RECT 22.950 165.600 25.050 167.700 ;
        RECT 29.400 163.050 30.450 190.950 ;
        RECT 43.950 188.400 46.050 190.500 ;
        RECT 31.950 182.100 34.050 184.200 ;
        RECT 32.400 178.050 33.450 182.100 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 31.950 175.950 34.050 178.050 ;
        RECT 38.400 177.900 39.600 178.650 ;
        RECT 37.950 175.800 40.050 177.900 ;
        RECT 44.100 168.600 45.300 188.400 ;
        RECT 62.400 183.600 63.450 205.950 ;
        RECT 65.400 187.050 66.450 209.400 ;
        RECT 70.950 208.800 73.050 210.900 ;
        RECT 76.950 208.950 79.050 211.050 ;
        RECT 83.400 210.900 84.600 211.650 ;
        RECT 82.950 208.800 85.050 210.900 ;
        RECT 88.950 208.950 91.050 211.050 ;
        RECT 89.400 193.050 90.450 208.950 ;
        RECT 92.400 202.050 93.450 283.950 ;
        RECT 98.400 280.050 99.450 293.100 ;
        RECT 101.400 283.050 102.450 331.950 ;
        RECT 107.400 328.050 108.450 332.400 ;
        RECT 112.950 328.950 115.050 332.400 ;
        RECT 115.950 331.950 118.050 332.400 ;
        RECT 124.950 331.950 127.050 334.050 ;
        RECT 131.400 332.400 132.600 334.800 ;
        RECT 137.400 334.050 138.450 338.250 ;
        RECT 106.950 325.950 109.050 328.050 ;
        RECT 116.400 322.050 117.450 331.950 ;
        RECT 131.400 325.050 132.450 332.400 ;
        RECT 136.950 331.950 139.050 334.050 ;
        RECT 140.400 328.050 141.450 343.950 ;
        RECT 143.400 343.050 144.450 355.950 ;
        RECT 146.400 349.050 147.450 358.950 ;
        RECT 154.950 358.800 157.050 360.900 ;
        RECT 148.950 349.950 151.050 352.050 ;
        RECT 145.950 346.950 148.050 349.050 ;
        RECT 142.950 340.950 145.050 343.050 ;
        RECT 149.400 339.600 150.450 349.950 ;
        RECT 151.950 346.950 154.050 349.050 ;
        RECT 152.400 343.050 153.450 346.950 ;
        RECT 157.950 344.400 160.050 346.500 ;
        RECT 151.950 340.950 154.050 343.050 ;
        RECT 149.400 337.350 150.600 339.600 ;
        RECT 145.950 334.950 148.050 337.050 ;
        RECT 148.950 334.950 151.050 337.050 ;
        RECT 154.950 334.950 157.050 337.050 ;
        RECT 146.400 333.900 147.600 334.650 ;
        RECT 145.950 331.800 148.050 333.900 ;
        RECT 155.400 333.450 156.600 334.650 ;
        RECT 152.400 332.400 156.600 333.450 ;
        RECT 139.950 325.950 142.050 328.050 ;
        RECT 146.400 325.050 147.450 331.800 ;
        RECT 152.400 328.050 153.450 332.400 ;
        RECT 151.950 325.950 154.050 328.050 ;
        RECT 130.950 322.950 133.050 325.050 ;
        RECT 145.950 322.950 148.050 325.050 ;
        RECT 115.950 319.950 118.050 322.050 ;
        RECT 106.950 303.300 109.050 305.400 ;
        RECT 106.950 299.700 108.150 303.300 ;
        RECT 106.950 297.600 109.050 299.700 ;
        RECT 100.950 280.950 103.050 283.050 ;
        RECT 106.950 282.600 108.150 297.600 ;
        RECT 109.950 289.950 112.050 292.050 ;
        RECT 110.400 288.450 111.600 289.650 ;
        RECT 110.400 287.400 114.450 288.450 ;
        RECT 106.950 280.500 109.050 282.600 ;
        RECT 97.950 277.950 100.050 280.050 ;
        RECT 113.400 274.050 114.450 287.400 ;
        RECT 116.400 286.050 117.450 319.950 ;
        RECT 152.400 310.050 153.450 325.950 ;
        RECT 158.700 324.600 159.900 344.400 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 164.400 333.900 165.600 334.650 ;
        RECT 163.950 331.800 166.050 333.900 ;
        RECT 157.950 322.500 160.050 324.600 ;
        RECT 151.950 307.950 154.050 310.050 ;
        RECT 170.400 307.050 171.450 376.950 ;
        RECT 175.950 370.950 178.050 373.050 ;
        RECT 181.950 370.950 184.050 373.050 ;
        RECT 194.400 372.600 195.450 376.950 ;
        RECT 176.400 370.200 177.600 370.950 ;
        RECT 182.400 370.200 183.600 370.950 ;
        RECT 194.400 370.350 195.600 372.600 ;
        RECT 202.950 371.100 205.050 373.200 ;
        RECT 203.400 370.350 204.600 371.100 ;
        RECT 175.950 367.800 178.050 369.900 ;
        RECT 178.950 367.800 181.050 369.900 ;
        RECT 181.950 367.800 184.050 369.900 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 202.950 367.950 205.050 370.050 ;
        RECT 172.950 364.950 175.050 367.050 ;
        RECT 179.400 365.400 180.600 367.500 ;
        RECT 173.400 352.050 174.450 364.950 ;
        RECT 179.400 361.050 180.450 365.400 ;
        RECT 184.950 364.950 187.050 367.050 ;
        RECT 191.400 366.900 192.600 367.650 ;
        RECT 178.950 358.950 181.050 361.050 ;
        RECT 172.950 349.950 175.050 352.050 ;
        RECT 178.950 344.400 181.050 346.500 ;
        RECT 172.950 338.100 175.050 340.200 ;
        RECT 173.400 322.050 174.450 338.100 ;
        RECT 178.950 329.400 180.150 344.400 ;
        RECT 182.400 339.450 183.600 339.600 ;
        RECT 185.400 339.450 186.450 364.950 ;
        RECT 190.950 364.800 193.050 366.900 ;
        RECT 199.950 364.950 202.050 367.050 ;
        RECT 200.400 355.050 201.450 364.950 ;
        RECT 206.700 360.600 207.900 380.400 ;
        RECT 217.950 376.950 220.050 379.050 ;
        RECT 226.950 377.700 228.150 381.300 ;
        RECT 235.950 379.950 238.050 382.050 ;
        RECT 253.950 379.950 256.050 382.050 ;
        RECT 274.950 379.950 277.050 382.050 ;
        RECT 286.950 379.950 289.050 382.050 ;
        RECT 211.950 371.100 214.050 373.200 ;
        RECT 212.400 370.350 213.600 371.100 ;
        RECT 211.950 367.950 214.050 370.050 ;
        RECT 205.950 358.500 208.050 360.600 ;
        RECT 218.400 358.050 219.450 376.950 ;
        RECT 220.950 373.950 223.050 376.050 ;
        RECT 226.950 375.600 229.050 377.700 ;
        RECT 232.950 376.950 235.050 379.050 ;
        RECT 211.950 355.950 214.050 358.050 ;
        RECT 217.950 355.950 220.050 358.050 ;
        RECT 199.950 352.950 202.050 355.050 ;
        RECT 208.950 352.950 211.050 355.050 ;
        RECT 196.950 348.450 199.050 349.050 ;
        RECT 202.950 348.450 205.050 349.050 ;
        RECT 196.950 347.400 205.050 348.450 ;
        RECT 196.950 346.950 199.050 347.400 ;
        RECT 202.950 346.950 205.050 347.400 ;
        RECT 187.950 343.950 190.050 346.050 ;
        RECT 199.950 343.950 202.050 346.050 ;
        RECT 182.400 338.400 186.450 339.450 ;
        RECT 182.400 337.350 183.600 338.400 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 188.400 334.050 189.450 343.950 ;
        RECT 193.950 338.100 196.050 340.200 ;
        RECT 200.400 339.600 201.450 343.950 ;
        RECT 194.400 337.350 195.600 338.100 ;
        RECT 200.400 337.350 201.600 339.600 ;
        RECT 193.950 334.950 196.050 337.050 ;
        RECT 196.950 334.950 199.050 337.050 ;
        RECT 199.950 334.950 202.050 337.050 ;
        RECT 202.950 334.950 205.050 337.050 ;
        RECT 187.950 331.950 190.050 334.050 ;
        RECT 197.400 333.900 198.600 334.650 ;
        RECT 196.950 331.800 199.050 333.900 ;
        RECT 203.400 332.400 204.600 334.650 ;
        RECT 178.950 327.300 181.050 329.400 ;
        RECT 178.950 323.700 180.150 327.300 ;
        RECT 172.950 319.950 175.050 322.050 ;
        RECT 178.950 321.600 181.050 323.700 ;
        RECT 199.950 307.950 202.050 310.050 ;
        RECT 148.950 304.950 151.050 307.050 ;
        RECT 169.950 304.950 172.050 307.050 ;
        RECT 193.950 304.950 196.050 307.050 ;
        RECT 118.950 301.950 121.050 304.050 ;
        RECT 115.950 283.950 118.050 286.050 ;
        RECT 115.950 280.800 118.050 282.900 ;
        RECT 112.950 271.950 115.050 274.050 ;
        RECT 94.950 260.100 97.050 262.200 ;
        RECT 103.950 260.100 106.050 262.200 ;
        RECT 109.950 261.000 112.050 265.050 ;
        RECT 95.400 256.050 96.450 260.100 ;
        RECT 104.400 259.350 105.600 260.100 ;
        RECT 110.400 259.350 111.600 261.000 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 101.400 256.050 102.600 256.650 ;
        RECT 94.950 253.950 97.050 256.050 ;
        RECT 97.950 254.400 102.600 256.050 ;
        RECT 107.400 255.900 108.600 256.650 ;
        RECT 116.400 255.900 117.450 280.800 ;
        RECT 119.400 262.050 120.450 301.950 ;
        RECT 124.950 292.950 127.050 295.050 ;
        RECT 130.950 292.950 133.050 295.050 ;
        RECT 136.950 292.950 139.050 295.050 ;
        RECT 142.950 293.100 145.050 295.200 ;
        RECT 149.400 294.600 150.450 304.950 ;
        RECT 169.950 295.950 172.050 298.050 ;
        RECT 165.000 294.600 169.050 295.050 ;
        RECT 125.400 292.200 126.600 292.950 ;
        RECT 131.400 292.200 132.600 292.950 ;
        RECT 124.950 289.800 127.050 291.900 ;
        RECT 127.950 289.800 130.050 291.900 ;
        RECT 130.950 289.800 133.050 291.900 ;
        RECT 121.950 286.950 124.050 289.050 ;
        RECT 128.400 288.750 129.600 289.500 ;
        RECT 122.400 265.050 123.450 286.950 ;
        RECT 127.950 286.650 130.050 288.750 ;
        RECT 137.400 274.050 138.450 292.950 ;
        RECT 143.400 292.350 144.600 293.100 ;
        RECT 149.400 292.350 150.600 294.600 ;
        RECT 164.400 292.950 169.050 294.600 ;
        RECT 164.400 292.350 165.600 292.950 ;
        RECT 142.950 289.950 145.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 160.950 289.950 163.050 292.050 ;
        RECT 163.950 289.950 166.050 292.050 ;
        RECT 146.400 287.400 147.600 289.650 ;
        RECT 152.400 287.400 153.600 289.650 ;
        RECT 161.400 288.900 162.600 289.650 ;
        RECT 170.400 289.050 171.450 295.950 ;
        RECT 172.950 293.100 175.050 295.200 ;
        RECT 178.950 294.000 181.050 298.050 ;
        RECT 146.400 280.050 147.450 287.400 ;
        RECT 145.950 277.950 148.050 280.050 ;
        RECT 136.950 271.950 139.050 274.050 ;
        RECT 137.400 268.050 138.450 271.950 ;
        RECT 136.950 265.950 139.050 268.050 ;
        RECT 121.950 262.950 124.050 265.050 ;
        RECT 118.950 259.950 121.050 262.050 ;
        RECT 121.950 257.100 124.050 259.200 ;
        RECT 137.400 259.050 138.450 265.950 ;
        RECT 152.400 265.050 153.450 287.400 ;
        RECT 160.950 286.800 163.050 288.900 ;
        RECT 169.950 286.950 172.050 289.050 ;
        RECT 151.950 262.950 154.050 265.050 ;
        RECT 148.950 259.950 151.050 262.050 ;
        RECT 136.950 256.950 139.050 259.050 ;
        RECT 142.950 257.100 145.050 259.200 ;
        RECT 97.950 253.950 102.000 254.400 ;
        RECT 106.950 253.800 109.050 255.900 ;
        RECT 115.950 253.800 118.050 255.900 ;
        RECT 122.400 254.400 123.600 256.800 ;
        RECT 122.400 250.050 123.450 254.400 ;
        RECT 121.950 247.950 124.050 250.050 ;
        RECT 94.950 244.950 97.050 247.050 ;
        RECT 91.950 199.950 94.050 202.050 ;
        RECT 88.950 190.950 91.050 193.050 ;
        RECT 64.950 184.950 67.050 187.050 ;
        RECT 62.400 181.500 63.600 183.600 ;
        RECT 76.950 183.000 79.050 187.050 ;
        RECT 85.950 184.950 88.050 187.050 ;
        RECT 77.400 181.350 78.600 183.000 ;
        RECT 46.950 178.950 49.050 181.050 ;
        RECT 58.950 179.100 61.050 181.200 ;
        RECT 61.950 179.100 64.050 181.200 ;
        RECT 64.950 179.100 67.050 181.200 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 47.400 177.450 48.600 178.650 ;
        RECT 47.400 176.400 51.450 177.450 ;
        RECT 43.950 166.500 46.050 168.600 ;
        RECT 50.400 166.050 51.450 176.400 ;
        RECT 59.400 176.400 60.600 178.800 ;
        RECT 65.400 177.000 66.600 178.800 ;
        RECT 80.400 177.900 81.600 178.650 ;
        RECT 49.950 163.950 52.050 166.050 ;
        RECT 10.950 160.950 13.050 163.050 ;
        RECT 22.950 160.950 25.050 163.050 ;
        RECT 28.950 160.950 31.050 163.050 ;
        RECT 13.950 138.000 16.050 142.050 ;
        RECT 14.400 136.350 15.600 138.000 ;
        RECT 10.950 133.950 13.050 136.050 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 4.950 130.950 7.050 133.050 ;
        RECT 11.400 132.900 12.600 133.650 ;
        RECT 10.950 130.800 13.050 132.900 ;
        RECT 17.400 131.400 18.600 133.650 ;
        RECT 17.400 124.050 18.450 131.400 ;
        RECT 23.400 130.050 24.450 160.950 ;
        RECT 49.950 142.950 52.050 145.050 ;
        RECT 40.950 139.950 43.050 142.050 ;
        RECT 31.950 137.100 34.050 139.200 ;
        RECT 32.400 136.350 33.600 137.100 ;
        RECT 28.950 133.950 31.050 136.050 ;
        RECT 31.950 133.950 34.050 136.050 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 29.400 132.000 30.600 133.650 ;
        RECT 22.950 127.950 25.050 130.050 ;
        RECT 28.950 127.950 31.050 132.000 ;
        RECT 35.400 131.400 36.600 133.650 ;
        RECT 4.950 121.950 7.050 124.050 ;
        RECT 16.950 121.950 19.050 124.050 ;
        RECT 1.950 100.950 4.050 103.050 ;
        RECT 5.400 28.200 6.450 121.950 ;
        RECT 16.950 111.000 19.050 115.050 ;
        RECT 35.400 112.050 36.450 131.400 ;
        RECT 41.400 121.050 42.450 139.950 ;
        RECT 50.400 138.600 51.450 142.950 ;
        RECT 59.400 141.450 60.450 176.400 ;
        RECT 64.950 172.950 67.050 177.000 ;
        RECT 79.950 175.800 82.050 177.900 ;
        RECT 86.400 175.050 87.450 184.950 ;
        RECT 92.400 183.600 93.450 199.950 ;
        RECT 95.400 187.050 96.450 244.950 ;
        RECT 106.950 229.950 109.050 232.050 ;
        RECT 102.000 219.450 106.050 220.050 ;
        RECT 101.400 217.950 106.050 219.450 ;
        RECT 101.400 216.600 102.450 217.950 ;
        RECT 107.400 217.050 108.450 229.950 ;
        RECT 122.400 229.050 123.450 247.950 ;
        RECT 121.950 226.950 124.050 229.050 ;
        RECT 127.950 226.950 130.050 229.050 ;
        RECT 121.950 220.950 124.050 223.050 ;
        RECT 112.950 219.450 117.000 220.050 ;
        RECT 112.950 217.950 117.450 219.450 ;
        RECT 101.400 214.350 102.600 216.600 ;
        RECT 106.950 214.950 109.050 217.050 ;
        RECT 116.400 216.600 117.450 217.950 ;
        RECT 122.400 216.600 123.450 220.950 ;
        RECT 116.400 214.350 117.600 216.600 ;
        RECT 122.400 214.350 123.600 216.600 ;
        RECT 128.400 216.450 129.450 226.950 ;
        RECT 133.950 224.400 136.050 226.500 ;
        RECT 131.400 216.450 132.600 216.600 ;
        RECT 128.400 215.400 132.600 216.450 ;
        RECT 131.400 214.350 132.600 215.400 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 103.950 211.950 106.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 118.950 211.950 121.050 214.050 ;
        RECT 121.950 211.950 124.050 214.050 ;
        RECT 130.950 211.950 133.050 214.050 ;
        RECT 104.400 210.900 105.600 211.650 ;
        RECT 103.950 208.800 106.050 210.900 ;
        RECT 113.400 209.400 114.600 211.650 ;
        RECT 119.400 210.900 120.600 211.650 ;
        RECT 113.400 202.050 114.450 209.400 ;
        RECT 118.950 208.800 121.050 210.900 ;
        RECT 134.700 204.600 135.900 224.400 ;
        RECT 145.950 220.950 148.050 223.050 ;
        RECT 139.950 215.100 142.050 217.200 ;
        RECT 140.400 214.350 141.600 215.100 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 133.950 202.500 136.050 204.600 ;
        RECT 112.950 199.950 115.050 202.050 ;
        RECT 127.950 193.950 130.050 196.050 ;
        RECT 124.950 190.950 127.050 193.050 ;
        RECT 110.400 188.400 120.450 189.450 ;
        RECT 94.950 184.950 97.050 187.050 ;
        RECT 106.950 184.950 109.050 187.050 ;
        RECT 92.400 181.350 93.600 183.600 ;
        RECT 97.950 182.100 100.050 184.200 ;
        RECT 98.400 181.350 99.600 182.100 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 95.400 177.900 96.600 178.650 ;
        RECT 94.950 175.800 97.050 177.900 ;
        RECT 101.400 176.400 102.600 178.650 ;
        RECT 85.950 172.950 88.050 175.050 ;
        RECT 101.400 172.050 102.450 176.400 ;
        RECT 103.950 175.950 106.050 178.050 ;
        RECT 107.400 177.900 108.450 184.950 ;
        RECT 110.400 184.050 111.450 188.400 ;
        RECT 109.950 181.950 112.050 184.050 ;
        RECT 112.950 183.000 115.050 187.050 ;
        RECT 119.400 183.600 120.450 188.400 ;
        RECT 125.400 184.050 126.450 190.950 ;
        RECT 113.400 181.350 114.600 183.000 ;
        RECT 119.400 181.350 120.600 183.600 ;
        RECT 124.950 181.950 127.050 184.050 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 121.950 178.950 124.050 181.050 ;
        RECT 116.400 177.900 117.600 178.650 ;
        RECT 122.400 177.900 123.600 178.650 ;
        RECT 128.400 177.900 129.450 193.950 ;
        RECT 139.950 190.950 142.050 193.050 ;
        RECT 133.950 183.000 136.050 187.050 ;
        RECT 140.400 183.600 141.450 190.950 ;
        RECT 134.400 181.350 135.600 183.000 ;
        RECT 140.400 181.350 141.600 183.600 ;
        RECT 133.950 178.950 136.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 137.400 177.900 138.600 178.650 ;
        RECT 100.950 169.950 103.050 172.050 ;
        RECT 104.400 145.050 105.450 175.950 ;
        RECT 106.950 175.800 109.050 177.900 ;
        RECT 115.950 175.800 118.050 177.900 ;
        RECT 121.950 175.800 124.050 177.900 ;
        RECT 127.950 175.800 130.050 177.900 ;
        RECT 136.950 175.800 139.050 177.900 ;
        RECT 121.950 172.650 124.050 174.750 ;
        RECT 118.950 169.950 121.050 172.050 ;
        RECT 115.950 154.950 118.050 157.050 ;
        RECT 91.950 142.950 94.050 145.050 ;
        RECT 56.400 141.000 60.450 141.450 ;
        RECT 55.950 140.400 60.450 141.000 ;
        RECT 50.400 136.350 51.600 138.600 ;
        RECT 55.950 136.950 58.050 140.400 ;
        RECT 64.950 137.100 67.050 139.200 ;
        RECT 65.400 136.350 66.600 137.100 ;
        RECT 70.950 136.950 73.050 139.050 ;
        RECT 79.950 137.100 82.050 139.200 ;
        RECT 87.000 138.600 91.050 139.050 ;
        RECT 46.950 133.950 49.050 136.050 ;
        RECT 49.950 133.950 52.050 136.050 ;
        RECT 52.950 133.950 55.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 64.950 133.950 67.050 136.050 ;
        RECT 47.400 132.900 48.600 133.650 ;
        RECT 46.950 130.800 49.050 132.900 ;
        RECT 53.400 132.450 54.600 133.650 ;
        RECT 55.950 132.450 58.050 132.900 ;
        RECT 53.400 131.400 58.050 132.450 ;
        RECT 55.950 130.800 58.050 131.400 ;
        RECT 62.400 131.400 63.600 133.650 ;
        RECT 47.400 124.050 48.450 130.800 ;
        RECT 52.950 127.950 55.050 130.050 ;
        RECT 46.950 121.950 49.050 124.050 ;
        RECT 40.950 118.950 43.050 121.050 ;
        RECT 13.500 108.300 15.600 110.400 ;
        RECT 17.400 108.900 18.600 111.000 ;
        RECT 34.950 109.950 37.050 112.050 ;
        RECT 43.950 109.950 46.050 112.050 ;
        RECT 11.400 103.200 12.600 105.600 ;
        RECT 10.950 103.050 13.050 103.200 ;
        RECT 7.950 101.100 13.050 103.050 ;
        RECT 13.950 102.900 14.850 108.300 ;
        RECT 16.950 106.800 19.050 108.900 ;
        RECT 20.700 105.900 22.800 107.700 ;
        RECT 15.750 104.700 24.300 105.900 ;
        RECT 15.750 103.800 17.850 104.700 ;
        RECT 13.950 101.700 20.850 102.900 ;
        RECT 7.950 100.950 10.950 101.100 ;
        RECT 13.950 94.500 15.150 101.700 ;
        RECT 16.950 98.100 19.050 100.200 ;
        RECT 19.950 99.300 20.850 101.700 ;
        RECT 17.400 95.400 18.600 98.100 ;
        RECT 19.950 97.200 22.050 99.300 ;
        RECT 23.400 95.700 24.300 104.700 ;
        RECT 34.950 104.100 37.050 106.200 ;
        RECT 35.400 103.350 36.600 104.100 ;
        RECT 25.950 101.100 28.050 103.200 ;
        RECT 26.400 99.900 27.600 101.100 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 38.400 99.900 39.600 100.650 ;
        RECT 25.950 97.800 28.050 99.900 ;
        RECT 37.950 97.800 40.050 99.900 ;
        RECT 13.500 92.400 15.600 94.500 ;
        RECT 16.950 91.950 19.050 94.050 ;
        RECT 23.100 93.600 25.200 95.700 ;
        RECT 10.950 67.950 13.050 70.050 ;
        RECT 11.400 60.600 12.450 67.950 ;
        RECT 17.400 61.050 18.450 91.950 ;
        RECT 44.400 76.050 45.450 109.950 ;
        RECT 53.400 106.200 54.450 127.950 ;
        RECT 56.400 121.050 57.450 130.800 ;
        RECT 62.400 124.050 63.450 131.400 ;
        RECT 61.950 121.950 64.050 124.050 ;
        RECT 71.400 121.050 72.450 136.950 ;
        RECT 80.400 136.350 81.600 137.100 ;
        RECT 86.400 136.950 91.050 138.600 ;
        RECT 86.400 136.350 87.600 136.950 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 77.400 132.900 78.600 133.650 ;
        RECT 76.950 130.800 79.050 132.900 ;
        RECT 83.400 131.400 84.600 133.650 ;
        RECT 79.950 127.950 82.050 130.050 ;
        RECT 55.950 118.950 58.050 121.050 ;
        RECT 70.950 118.950 73.050 121.050 ;
        RECT 76.950 112.950 79.050 115.050 ;
        RECT 70.950 109.950 73.050 112.050 ;
        RECT 46.950 103.950 49.050 106.050 ;
        RECT 52.950 104.100 55.050 106.200 ;
        RECT 58.950 104.100 61.050 106.200 ;
        RECT 71.400 105.600 72.450 109.950 ;
        RECT 77.400 105.600 78.450 112.950 ;
        RECT 80.400 112.050 81.450 127.950 ;
        RECT 83.400 127.050 84.450 131.400 ;
        RECT 88.950 130.950 91.050 133.050 ;
        RECT 82.950 124.950 85.050 127.050 ;
        RECT 89.400 121.050 90.450 130.950 ;
        RECT 88.950 118.950 91.050 121.050 ;
        RECT 92.400 115.050 93.450 142.950 ;
        RECT 100.800 141.300 102.900 143.400 ;
        RECT 103.950 142.950 106.050 145.050 ;
        RECT 110.400 142.500 112.500 144.600 ;
        RECT 97.950 137.100 100.050 139.200 ;
        RECT 98.400 136.050 99.600 137.100 ;
        RECT 97.950 133.800 100.050 136.050 ;
        RECT 101.700 132.300 102.600 141.300 ;
        RECT 103.950 137.700 106.050 139.800 ;
        RECT 107.400 138.900 108.600 141.600 ;
        RECT 105.150 135.300 106.050 137.700 ;
        RECT 106.950 136.800 109.050 138.900 ;
        RECT 110.850 135.300 112.050 142.500 ;
        RECT 116.400 142.050 117.450 154.950 ;
        RECT 115.950 139.950 118.050 142.050 ;
        RECT 105.150 134.100 112.050 135.300 ;
        RECT 108.150 132.300 110.250 133.200 ;
        RECT 101.700 131.100 110.250 132.300 ;
        RECT 103.200 129.300 105.300 131.100 ;
        RECT 106.950 127.950 109.050 130.200 ;
        RECT 111.150 128.700 112.050 134.100 ;
        RECT 112.950 133.800 115.050 135.900 ;
        RECT 115.950 133.950 118.050 138.900 ;
        RECT 113.400 131.400 114.600 133.800 ;
        RECT 107.400 125.400 108.600 127.950 ;
        RECT 110.400 126.600 112.500 128.700 ;
        RECT 85.950 112.950 88.050 115.050 ;
        RECT 91.950 112.950 94.050 115.050 ;
        RECT 100.950 112.950 103.050 115.050 ;
        RECT 79.950 109.950 82.050 112.050 ;
        RECT 47.400 99.900 48.450 103.950 ;
        RECT 53.400 103.350 54.600 104.100 ;
        RECT 59.400 103.350 60.600 104.100 ;
        RECT 71.400 103.500 72.600 105.600 ;
        RECT 77.400 103.500 78.600 105.600 ;
        RECT 52.950 100.950 55.050 103.050 ;
        RECT 55.950 100.950 58.050 103.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 70.950 101.100 73.050 103.200 ;
        RECT 73.950 101.100 76.050 103.200 ;
        RECT 76.950 101.100 79.050 103.200 ;
        RECT 79.950 101.100 82.050 103.200 ;
        RECT 46.950 97.800 49.050 99.900 ;
        RECT 56.400 98.400 57.600 100.650 ;
        RECT 74.400 100.050 75.600 100.800 ;
        RECT 80.400 100.050 81.600 100.800 ;
        RECT 86.400 100.050 87.450 112.950 ;
        RECT 94.200 107.100 96.300 109.200 ;
        RECT 98.400 108.900 99.600 111.600 ;
        RECT 92.400 103.200 93.600 105.600 ;
        RECT 91.950 101.100 94.050 103.200 ;
        RECT 94.950 102.000 95.850 107.100 ;
        RECT 97.650 106.800 100.050 108.900 ;
        RECT 101.400 105.900 102.450 112.950 ;
        RECT 104.250 107.400 106.350 109.500 ;
        RECT 101.400 105.000 103.800 105.900 ;
        RECT 96.750 103.800 103.800 105.000 ;
        RECT 96.750 102.900 98.850 103.800 ;
        RECT 101.700 102.000 103.800 102.900 ;
        RECT 94.950 101.100 103.800 102.000 ;
        RECT 56.400 97.050 57.450 98.400 ;
        RECT 61.950 97.950 64.050 100.050 ;
        RECT 56.400 95.400 61.050 97.050 ;
        RECT 57.000 94.950 61.050 95.400 ;
        RECT 28.950 73.950 31.050 76.050 ;
        RECT 43.950 73.950 46.050 76.050 ;
        RECT 22.950 69.300 25.050 71.400 ;
        RECT 23.850 65.700 25.050 69.300 ;
        RECT 22.950 63.600 25.050 65.700 ;
        RECT 11.400 58.350 12.600 60.600 ;
        RECT 16.950 58.950 19.050 61.050 ;
        RECT 10.950 55.950 13.050 58.050 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 14.400 54.900 15.600 55.650 ;
        RECT 20.400 54.900 21.600 55.650 ;
        RECT 13.950 52.800 16.050 54.900 ;
        RECT 19.950 52.800 22.050 54.900 ;
        RECT 23.850 48.600 25.050 63.600 ;
        RECT 22.950 46.500 25.050 48.600 ;
        RECT 22.950 32.400 25.050 34.500 ;
        RECT 4.950 26.100 7.050 28.200 ;
        RECT 13.950 26.100 16.050 28.200 ;
        RECT 19.950 26.100 22.050 28.200 ;
        RECT 14.400 25.350 15.600 26.100 ;
        RECT 20.400 25.350 21.600 26.100 ;
        RECT 10.950 22.950 13.050 25.050 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 19.950 22.950 22.050 25.050 ;
        RECT 11.400 21.900 12.600 22.650 ;
        RECT 10.950 19.800 13.050 21.900 ;
        RECT 23.850 17.400 25.050 32.400 ;
        RECT 29.400 21.900 30.450 73.950 ;
        RECT 43.950 68.400 46.050 70.500 ;
        RECT 62.400 70.050 63.450 97.950 ;
        RECT 67.950 94.950 70.050 100.050 ;
        RECT 73.950 97.950 76.050 100.050 ;
        RECT 79.950 97.950 82.050 100.050 ;
        RECT 85.950 97.950 88.050 100.050 ;
        RECT 94.950 94.500 95.850 101.100 ;
        RECT 101.700 100.800 103.800 101.100 ;
        RECT 97.650 98.100 99.750 100.200 ;
        RECT 98.400 95.400 99.600 98.100 ;
        RECT 104.700 94.800 105.600 107.400 ;
        RECT 119.400 105.600 120.450 169.950 ;
        RECT 122.400 139.050 123.450 172.650 ;
        RECT 146.400 172.050 147.450 220.950 ;
        RECT 149.400 193.050 150.450 259.950 ;
        RECT 152.400 250.050 153.450 262.950 ;
        RECT 161.400 261.600 162.450 286.800 ;
        RECT 173.400 286.050 174.450 293.100 ;
        RECT 179.400 292.350 180.600 294.000 ;
        RECT 184.950 293.100 187.050 295.200 ;
        RECT 185.400 292.350 186.600 293.100 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 184.950 289.950 187.050 292.050 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 175.950 286.950 178.050 289.050 ;
        RECT 182.400 287.400 183.600 289.650 ;
        RECT 188.400 288.900 189.600 289.650 ;
        RECT 172.950 283.950 175.050 286.050 ;
        RECT 176.400 270.450 177.450 286.950 ;
        RECT 182.400 280.050 183.450 287.400 ;
        RECT 187.950 286.800 190.050 288.900 ;
        RECT 184.950 283.950 187.050 286.050 ;
        RECT 181.950 277.950 184.050 280.050 ;
        RECT 176.400 270.000 183.450 270.450 ;
        RECT 176.400 269.400 184.050 270.000 ;
        RECT 178.800 265.950 180.900 268.050 ;
        RECT 181.950 265.950 184.050 269.400 ;
        RECT 161.400 259.500 162.600 261.600 ;
        RECT 172.950 260.100 175.050 262.200 ;
        RECT 179.400 261.600 180.450 265.950 ;
        RECT 185.400 262.200 186.450 283.950 ;
        RECT 194.400 280.050 195.450 304.950 ;
        RECT 200.400 294.600 201.450 307.950 ;
        RECT 203.400 295.050 204.450 332.400 ;
        RECT 209.400 328.050 210.450 352.950 ;
        RECT 212.400 340.200 213.450 355.950 ;
        RECT 211.950 338.100 214.050 340.200 ;
        RECT 221.400 339.600 222.450 373.950 ;
        RECT 226.950 360.600 228.150 375.600 ;
        RECT 233.400 373.200 234.450 376.950 ;
        RECT 232.950 371.100 235.050 373.200 ;
        RECT 229.950 367.950 232.050 370.050 ;
        RECT 230.400 366.900 231.600 367.650 ;
        RECT 229.950 364.800 232.050 366.900 ;
        RECT 226.950 358.500 229.050 360.600 ;
        RECT 236.400 349.050 237.450 379.950 ;
        RECT 271.950 376.950 274.050 379.050 ;
        RECT 241.950 372.000 244.050 376.050 ;
        RECT 242.400 370.200 243.600 372.000 ;
        RECT 250.950 370.950 253.050 373.050 ;
        RECT 256.950 370.950 259.050 373.050 ;
        RECT 265.950 371.100 268.050 373.200 ;
        RECT 251.400 370.200 252.600 370.950 ;
        RECT 241.950 367.800 244.050 369.900 ;
        RECT 247.950 367.800 250.050 369.900 ;
        RECT 250.950 367.800 253.050 369.900 ;
        RECT 244.950 364.800 247.050 366.900 ;
        RECT 248.400 365.400 249.600 367.500 ;
        RECT 245.400 351.450 246.450 364.800 ;
        RECT 248.400 361.050 249.450 365.400 ;
        RECT 253.800 364.950 255.900 367.050 ;
        RECT 257.400 366.900 258.450 370.950 ;
        RECT 266.400 370.350 267.600 371.100 ;
        RECT 262.950 367.950 265.050 370.050 ;
        RECT 265.950 367.950 268.050 370.050 ;
        RECT 263.400 366.900 264.600 367.650 ;
        RECT 247.950 358.950 250.050 361.050 ;
        RECT 254.400 352.050 255.450 364.950 ;
        RECT 256.950 364.800 259.050 366.900 ;
        RECT 262.950 364.800 265.050 366.900 ;
        RECT 245.400 350.400 249.450 351.450 ;
        RECT 235.950 346.950 238.050 349.050 ;
        RECT 212.400 331.050 213.450 338.100 ;
        RECT 221.400 337.500 222.600 339.600 ;
        RECT 232.950 338.100 235.050 340.200 ;
        RECT 238.950 339.000 241.050 343.050 ;
        RECT 233.400 337.350 234.600 338.100 ;
        RECT 239.400 337.350 240.600 339.000 ;
        RECT 217.950 335.100 220.050 337.200 ;
        RECT 220.950 335.100 223.050 337.200 ;
        RECT 223.950 335.100 226.050 337.200 ;
        RECT 232.950 334.950 235.050 337.050 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 238.950 334.950 241.050 337.050 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 218.400 333.900 219.600 334.800 ;
        RECT 217.950 331.800 220.050 333.900 ;
        RECT 224.400 333.000 225.600 334.800 ;
        RECT 236.400 333.900 237.600 334.650 ;
        RECT 211.950 328.950 214.050 331.050 ;
        RECT 208.950 325.950 211.050 328.050 ;
        RECT 218.400 325.050 219.450 331.800 ;
        RECT 223.950 328.950 226.050 333.000 ;
        RECT 235.950 331.800 238.050 333.900 ;
        RECT 242.400 332.400 243.600 334.650 ;
        RECT 242.400 328.050 243.450 332.400 ;
        RECT 241.950 325.950 244.050 328.050 ;
        RECT 217.950 322.950 220.050 325.050 ;
        RECT 248.400 309.450 249.450 350.400 ;
        RECT 253.950 349.950 256.050 352.050 ;
        RECT 257.400 346.050 258.450 364.800 ;
        RECT 272.400 364.050 273.450 376.950 ;
        RECT 280.950 372.000 283.050 376.050 ;
        RECT 287.400 372.600 288.450 379.950 ;
        RECT 293.400 373.050 294.450 409.950 ;
        RECT 301.950 406.950 304.050 411.000 ;
        RECT 311.400 409.050 312.450 439.950 ;
        RECT 314.400 439.050 315.450 443.400 ;
        RECT 319.950 442.800 322.050 444.900 ;
        RECT 326.400 443.400 327.600 445.650 ;
        RECT 322.950 439.950 325.050 442.050 ;
        RECT 313.950 436.950 316.050 439.050 ;
        RECT 316.950 417.000 319.050 421.050 ;
        RECT 323.400 417.450 324.450 439.950 ;
        RECT 326.400 430.050 327.450 443.400 ;
        RECT 331.950 441.450 334.050 445.050 ;
        RECT 335.400 442.050 336.450 451.950 ;
        RECT 341.400 450.600 342.450 472.950 ;
        RECT 386.400 469.050 387.450 478.950 ;
        RECT 385.950 466.950 388.050 469.050 ;
        RECT 389.400 466.050 390.450 487.950 ;
        RECT 392.400 483.450 393.450 505.950 ;
        RECT 395.400 490.050 396.450 511.950 ;
        RECT 407.400 504.450 408.450 520.950 ;
        RECT 409.950 520.800 412.050 522.900 ;
        RECT 416.400 521.400 417.600 523.650 ;
        RECT 425.400 523.050 426.450 526.950 ;
        RECT 431.400 526.200 432.600 526.950 ;
        RECT 446.400 526.350 447.600 528.000 ;
        RECT 430.950 523.800 433.050 525.900 ;
        RECT 433.950 523.800 436.050 525.900 ;
        RECT 436.950 523.800 439.050 525.900 ;
        RECT 445.950 523.950 448.050 526.050 ;
        RECT 424.950 522.450 427.050 523.050 ;
        RECT 434.400 522.750 435.600 523.500 ;
        RECT 424.950 521.400 429.450 522.450 ;
        RECT 410.400 508.050 411.450 520.800 ;
        RECT 412.950 514.950 415.050 517.050 ;
        RECT 409.950 505.950 412.050 508.050 ;
        RECT 413.400 505.050 414.450 514.950 ;
        RECT 416.400 514.050 417.450 521.400 ;
        RECT 424.950 520.950 427.050 521.400 ;
        RECT 415.950 511.950 418.050 514.050 ;
        RECT 404.400 504.000 408.450 504.450 ;
        RECT 403.950 503.400 408.450 504.000 ;
        RECT 403.950 499.950 406.050 503.400 ;
        RECT 412.950 502.950 415.050 505.050 ;
        RECT 428.400 502.050 429.450 521.400 ;
        RECT 433.950 520.650 436.050 522.750 ;
        RECT 442.950 517.950 445.050 520.050 ;
        RECT 443.400 514.050 444.450 517.950 ;
        RECT 449.700 516.600 450.900 536.400 ;
        RECT 457.950 535.950 460.050 538.050 ;
        RECT 454.950 527.100 457.050 529.200 ;
        RECT 455.400 526.350 456.600 527.100 ;
        RECT 454.950 523.950 457.050 526.050 ;
        RECT 448.950 514.500 451.050 516.600 ;
        RECT 442.950 511.950 445.050 514.050 ;
        RECT 461.400 511.050 462.450 541.950 ;
        RECT 463.950 538.950 466.050 541.050 ;
        RECT 464.400 532.050 465.450 538.950 ;
        RECT 469.950 537.300 472.050 539.400 ;
        RECT 469.950 533.700 471.150 537.300 ;
        RECT 475.950 535.950 478.050 538.050 ;
        RECT 463.950 529.950 466.050 532.050 ;
        RECT 469.950 531.600 472.050 533.700 ;
        RECT 451.950 508.950 454.050 511.050 ;
        RECT 460.950 508.950 463.050 511.050 ;
        RECT 430.950 502.950 433.050 505.050 ;
        RECT 427.950 499.950 430.050 502.050 ;
        RECT 405.000 498.450 409.050 499.050 ;
        RECT 404.400 496.950 409.050 498.450 ;
        RECT 404.400 495.600 405.450 496.950 ;
        RECT 404.400 493.500 405.600 495.600 ;
        RECT 409.950 495.450 412.050 496.050 ;
        RECT 416.400 495.450 417.600 495.600 ;
        RECT 409.950 494.400 417.600 495.450 ;
        RECT 409.950 493.950 412.050 494.400 ;
        RECT 416.400 493.350 417.600 494.400 ;
        RECT 421.950 494.100 424.050 496.200 ;
        RECT 422.400 493.350 423.600 494.100 ;
        RECT 400.950 491.100 403.050 493.200 ;
        RECT 403.950 491.100 406.050 493.200 ;
        RECT 406.950 491.100 409.050 493.200 ;
        RECT 415.950 490.950 418.050 493.050 ;
        RECT 418.950 490.950 421.050 493.050 ;
        RECT 421.950 490.950 424.050 493.050 ;
        RECT 424.950 490.950 427.050 493.050 ;
        RECT 401.400 490.050 402.600 490.800 ;
        RECT 394.950 487.950 397.050 490.050 ;
        RECT 400.950 487.950 403.050 490.050 ;
        RECT 407.400 489.000 408.600 490.800 ;
        RECT 406.950 484.950 409.050 489.000 ;
        RECT 419.400 488.400 420.600 490.650 ;
        RECT 425.400 490.050 426.600 490.650 ;
        RECT 425.400 488.400 430.050 490.050 ;
        RECT 392.400 482.400 396.450 483.450 ;
        RECT 395.400 472.050 396.450 482.400 ;
        RECT 419.400 481.050 420.450 488.400 ;
        RECT 426.000 487.950 430.050 488.400 ;
        RECT 427.950 484.800 430.050 486.900 ;
        RECT 418.950 478.950 421.050 481.050 ;
        RECT 428.400 472.050 429.450 484.800 ;
        RECT 394.950 469.950 397.050 472.050 ;
        RECT 412.950 469.950 415.050 472.050 ;
        RECT 427.950 469.950 430.050 472.050 ;
        RECT 388.950 463.950 391.050 466.050 ;
        RECT 406.950 463.950 409.050 466.050 ;
        RECT 358.950 458.400 361.050 460.500 ;
        RECT 379.950 459.300 382.050 461.400 ;
        RECT 341.400 448.200 342.600 450.600 ;
        RECT 355.950 450.000 358.050 454.050 ;
        RECT 356.400 448.350 357.600 450.000 ;
        RECT 340.950 445.800 343.050 447.900 ;
        RECT 343.950 445.800 346.050 447.900 ;
        RECT 346.950 445.800 349.050 447.900 ;
        RECT 355.950 445.950 358.050 448.050 ;
        RECT 344.400 444.000 345.600 445.500 ;
        RECT 329.400 441.000 334.050 441.450 ;
        RECT 329.400 440.400 333.450 441.000 ;
        RECT 325.950 427.950 328.050 430.050 ;
        RECT 317.400 415.350 318.600 417.000 ;
        RECT 323.400 416.400 327.450 417.450 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 319.950 412.950 322.050 415.050 ;
        RECT 320.400 411.900 321.600 412.650 ;
        RECT 319.950 409.800 322.050 411.900 ;
        RECT 326.400 411.450 327.450 416.400 ;
        RECT 329.400 412.050 330.450 440.400 ;
        RECT 334.950 439.950 337.050 442.050 ;
        RECT 343.950 439.950 346.050 444.000 ;
        RECT 352.950 442.950 355.050 445.050 ;
        RECT 353.400 430.050 354.450 442.950 ;
        RECT 359.700 438.600 360.900 458.400 ;
        RECT 379.950 455.700 381.150 459.300 ;
        RECT 370.950 451.950 373.050 454.050 ;
        RECT 379.950 453.600 382.050 455.700 ;
        RECT 364.950 449.100 367.050 451.200 ;
        RECT 365.400 448.350 366.600 449.100 ;
        RECT 364.950 445.950 367.050 448.050 ;
        RECT 371.400 444.450 372.450 451.950 ;
        RECT 368.400 443.400 372.450 444.450 ;
        RECT 358.950 436.500 361.050 438.600 ;
        RECT 352.950 427.950 355.050 430.050 ;
        RECT 352.950 422.400 355.050 424.500 ;
        RECT 337.950 416.100 340.050 418.200 ;
        RECT 343.950 416.100 346.050 418.200 ;
        RECT 338.400 415.350 339.600 416.100 ;
        RECT 344.400 415.350 345.600 416.100 ;
        RECT 334.950 412.950 337.050 415.050 ;
        RECT 337.950 412.950 340.050 415.050 ;
        RECT 340.950 412.950 343.050 415.050 ;
        RECT 343.950 412.950 346.050 415.050 ;
        RECT 349.950 412.950 352.050 415.050 ;
        RECT 323.400 410.400 327.450 411.450 ;
        RECT 310.950 406.950 313.050 409.050 ;
        RECT 320.400 391.050 321.450 409.800 ;
        RECT 323.400 394.050 324.450 410.400 ;
        RECT 328.950 409.950 331.050 412.050 ;
        RECT 335.400 411.900 336.600 412.650 ;
        RECT 334.950 409.800 337.050 411.900 ;
        RECT 341.400 410.400 342.600 412.650 ;
        RECT 350.400 411.450 351.600 412.650 ;
        RECT 347.400 410.400 351.600 411.450 ;
        RECT 341.400 409.050 342.450 410.400 ;
        RECT 340.950 406.950 343.050 409.050 ;
        RECT 322.950 391.950 325.050 394.050 ;
        RECT 319.950 388.950 322.050 391.050 ;
        RECT 328.950 376.950 331.050 379.050 ;
        RECT 298.950 373.950 301.050 376.050 ;
        RECT 281.400 370.200 282.600 372.000 ;
        RECT 287.400 370.200 288.600 372.600 ;
        RECT 292.950 370.950 295.050 373.050 ;
        RECT 277.950 367.800 280.050 369.900 ;
        RECT 280.950 367.800 283.050 369.900 ;
        RECT 283.950 367.800 286.050 369.900 ;
        RECT 286.950 367.800 289.050 369.900 ;
        RECT 289.950 367.800 292.050 369.900 ;
        RECT 295.950 367.950 298.050 370.050 ;
        RECT 274.950 364.950 277.050 367.050 ;
        RECT 278.400 365.400 279.600 367.500 ;
        RECT 284.400 366.000 285.600 367.500 ;
        RECT 290.400 366.750 291.600 367.500 ;
        RECT 271.950 361.950 274.050 364.050 ;
        RECT 275.400 361.050 276.450 364.950 ;
        RECT 268.950 358.950 271.050 361.050 ;
        RECT 274.950 358.950 277.050 361.050 ;
        RECT 269.400 349.050 270.450 358.950 ;
        RECT 271.950 349.950 274.050 352.050 ;
        RECT 268.950 346.950 271.050 349.050 ;
        RECT 250.950 343.950 253.050 346.050 ;
        RECT 256.950 343.950 259.050 346.050 ;
        RECT 251.400 340.050 252.450 343.950 ;
        RECT 250.950 337.950 253.050 340.050 ;
        RECT 256.950 338.250 259.050 340.350 ;
        RECT 257.400 337.500 258.600 338.250 ;
        RECT 265.950 337.950 268.050 340.050 ;
        RECT 272.400 339.600 273.450 349.950 ;
        RECT 278.400 340.050 279.450 365.400 ;
        RECT 283.950 361.950 286.050 366.000 ;
        RECT 289.950 364.650 292.050 366.750 ;
        RECT 280.950 358.950 283.050 361.050 ;
        RECT 253.950 335.100 256.050 337.200 ;
        RECT 256.950 335.100 259.050 337.200 ;
        RECT 259.950 335.100 262.050 337.200 ;
        RECT 254.400 334.050 255.600 334.800 ;
        RECT 260.400 334.050 261.600 334.800 ;
        RECT 253.950 331.950 256.050 334.050 ;
        RECT 259.950 333.450 262.050 334.050 ;
        RECT 257.400 332.400 262.050 333.450 ;
        RECT 250.950 309.450 253.050 310.050 ;
        RECT 248.400 308.400 253.050 309.450 ;
        RECT 250.950 307.950 253.050 308.400 ;
        RECT 221.400 299.400 228.450 300.450 ;
        RECT 200.400 292.200 201.600 294.600 ;
        RECT 202.950 292.950 205.050 295.050 ;
        RECT 205.950 292.950 208.050 295.050 ;
        RECT 211.950 292.950 214.050 295.050 ;
        RECT 218.400 294.450 219.600 294.600 ;
        RECT 221.400 294.450 222.450 299.400 ;
        RECT 218.400 293.400 222.450 294.450 ;
        RECT 223.950 294.000 226.050 298.050 ;
        RECT 227.400 295.050 228.450 299.400 ;
        RECT 235.800 297.300 237.900 299.400 ;
        RECT 245.400 298.500 247.500 300.600 ;
        RECT 206.400 292.200 207.600 292.950 ;
        RECT 199.950 289.800 202.050 291.900 ;
        RECT 202.950 289.800 205.050 291.900 ;
        RECT 205.950 289.800 208.050 291.900 ;
        RECT 203.400 288.750 204.600 289.500 ;
        RECT 202.950 286.650 205.050 288.750 ;
        RECT 193.950 277.950 196.050 280.050 ;
        RECT 212.400 274.050 213.450 292.950 ;
        RECT 218.400 292.200 219.600 293.400 ;
        RECT 224.400 292.200 225.600 294.000 ;
        RECT 226.950 292.950 229.050 295.050 ;
        RECT 233.400 291.900 234.600 294.600 ;
        RECT 217.950 289.800 220.050 291.900 ;
        RECT 220.950 289.800 223.050 291.900 ;
        RECT 223.950 289.800 226.050 291.900 ;
        RECT 232.950 289.800 235.050 291.900 ;
        RECT 221.400 288.750 222.600 289.500 ;
        RECT 220.950 286.650 223.050 288.750 ;
        RECT 233.400 274.050 234.450 289.800 ;
        RECT 236.700 288.300 237.600 297.300 ;
        RECT 238.950 293.700 241.050 295.800 ;
        RECT 242.400 294.900 243.600 297.600 ;
        RECT 240.150 291.300 241.050 293.700 ;
        RECT 241.950 292.800 244.050 294.900 ;
        RECT 245.850 291.300 247.050 298.500 ;
        RECT 251.400 292.050 252.450 307.950 ;
        RECT 257.400 301.050 258.450 332.400 ;
        RECT 259.950 331.950 262.050 332.400 ;
        RECT 266.400 328.050 267.450 337.950 ;
        RECT 272.400 337.350 273.600 339.600 ;
        RECT 277.950 337.950 280.050 340.050 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 275.400 334.050 276.600 334.650 ;
        RECT 275.400 331.950 280.050 334.050 ;
        RECT 265.950 325.950 268.050 328.050 ;
        RECT 271.950 319.950 274.050 322.050 ;
        RECT 265.950 304.950 268.050 307.050 ;
        RECT 256.950 298.950 259.050 301.050 ;
        RECT 253.950 292.950 256.050 295.050 ;
        RECT 250.050 291.900 252.450 292.050 ;
        RECT 240.150 290.100 247.050 291.300 ;
        RECT 243.150 288.300 245.250 289.200 ;
        RECT 236.700 287.100 245.250 288.300 ;
        RECT 238.200 285.300 240.300 287.100 ;
        RECT 241.950 284.100 244.050 286.200 ;
        RECT 246.150 284.700 247.050 290.100 ;
        RECT 247.950 289.950 252.450 291.900 ;
        RECT 247.950 289.800 250.050 289.950 ;
        RECT 248.400 287.400 249.600 289.800 ;
        RECT 242.400 281.400 243.600 284.100 ;
        RECT 245.400 282.600 247.500 284.700 ;
        RECT 242.400 277.050 243.450 281.400 ;
        RECT 241.950 274.950 244.050 277.050 ;
        RECT 202.950 271.950 205.050 274.050 ;
        RECT 211.950 271.950 214.050 274.050 ;
        RECT 232.950 271.950 235.050 274.050 ;
        RECT 244.950 271.950 247.050 274.050 ;
        RECT 196.950 265.950 199.050 268.050 ;
        RECT 173.400 259.350 174.600 260.100 ;
        RECT 179.400 259.350 180.600 261.600 ;
        RECT 184.950 260.100 187.050 262.200 ;
        RECT 190.950 260.100 193.050 262.200 ;
        RECT 197.400 261.600 198.450 265.950 ;
        RECT 157.950 257.100 160.050 259.200 ;
        RECT 160.950 257.100 163.050 259.200 ;
        RECT 163.950 257.100 166.050 259.200 ;
        RECT 172.950 256.950 175.050 259.050 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 178.950 256.950 181.050 259.050 ;
        RECT 158.400 256.050 159.600 256.800 ;
        RECT 164.400 256.050 165.600 256.800 ;
        RECT 157.950 253.950 160.050 256.050 ;
        RECT 163.950 253.950 166.050 256.050 ;
        RECT 176.400 255.900 177.600 256.650 ;
        RECT 185.400 256.050 186.450 260.100 ;
        RECT 191.400 259.350 192.600 260.100 ;
        RECT 197.400 259.350 198.600 261.600 ;
        RECT 203.400 261.450 204.450 271.950 ;
        RECT 208.950 266.400 211.050 268.500 ;
        RECT 206.400 261.450 207.600 261.600 ;
        RECT 203.400 260.400 207.600 261.450 ;
        RECT 206.400 259.350 207.600 260.400 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 196.950 256.950 199.050 259.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 151.950 247.950 154.050 250.050 ;
        RECT 164.400 232.050 165.450 253.950 ;
        RECT 175.950 253.800 178.050 255.900 ;
        RECT 184.950 253.950 187.050 256.050 ;
        RECT 194.400 255.900 195.600 256.650 ;
        RECT 193.950 253.800 196.050 255.900 ;
        RECT 209.850 251.400 211.050 266.400 ;
        RECT 214.950 265.950 217.050 268.050 ;
        RECT 229.950 266.400 232.050 268.500 ;
        RECT 199.950 247.950 202.050 250.050 ;
        RECT 208.950 249.300 211.050 251.400 ;
        RECT 200.400 235.050 201.450 247.950 ;
        RECT 202.950 244.950 205.050 247.050 ;
        RECT 209.850 245.700 211.050 249.300 ;
        RECT 199.950 232.950 202.050 235.050 ;
        RECT 163.950 229.950 166.050 232.050 ;
        RECT 175.950 229.950 178.050 232.050 ;
        RECT 154.950 225.300 157.050 227.400 ;
        RECT 154.950 221.700 156.150 225.300 ;
        RECT 154.950 219.600 157.050 221.700 ;
        RECT 154.950 204.600 156.150 219.600 ;
        RECT 157.950 211.950 160.050 214.050 ;
        RECT 158.400 210.450 159.600 211.650 ;
        RECT 164.400 210.450 165.450 229.950 ;
        RECT 176.400 216.600 177.450 229.950 ;
        RECT 190.950 228.450 193.050 232.050 ;
        RECT 196.950 229.950 199.050 232.050 ;
        RECT 190.950 228.000 195.450 228.450 ;
        RECT 191.400 227.400 195.450 228.000 ;
        RECT 190.950 223.950 193.050 226.050 ;
        RECT 191.400 217.200 192.450 223.950 ;
        RECT 194.400 220.050 195.450 227.400 ;
        RECT 193.950 217.950 196.050 220.050 ;
        RECT 176.400 214.350 177.600 216.600 ;
        RECT 190.950 215.100 193.050 217.200 ;
        RECT 197.400 216.600 198.450 229.950 ;
        RECT 191.400 214.350 192.600 215.100 ;
        RECT 197.400 214.350 198.600 216.600 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 187.950 211.950 190.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 193.950 211.950 196.050 214.050 ;
        RECT 196.950 211.950 199.050 214.050 ;
        RECT 158.400 209.400 165.450 210.450 ;
        RECT 173.400 209.400 174.600 211.650 ;
        RECT 179.400 210.900 180.600 211.650 ;
        RECT 154.950 202.500 157.050 204.600 ;
        RECT 148.950 190.950 151.050 193.050 ;
        RECT 160.950 190.950 163.050 193.050 ;
        RECT 148.950 184.950 151.050 187.050 ;
        RECT 149.400 178.050 150.450 184.950 ;
        RECT 154.950 179.100 157.050 181.200 ;
        RECT 148.950 175.950 151.050 178.050 ;
        RECT 155.400 176.400 156.600 178.800 ;
        RECT 136.950 169.950 139.050 172.050 ;
        RECT 145.950 169.950 148.050 172.050 ;
        RECT 130.950 148.950 133.050 151.050 ;
        RECT 121.950 136.950 124.050 139.050 ;
        RECT 131.400 138.600 132.450 148.950 ;
        RECT 131.400 136.350 132.600 138.600 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 130.950 133.950 133.050 136.050 ;
        RECT 125.400 133.050 126.600 133.650 ;
        RECT 121.950 131.400 126.600 133.050 ;
        RECT 137.400 132.450 138.450 169.950 ;
        RECT 155.400 166.050 156.450 176.400 ;
        RECT 154.950 163.950 157.050 166.050 ;
        RECT 151.950 142.950 154.050 145.050 ;
        RECT 139.950 137.100 142.050 142.050 ;
        RECT 145.950 137.100 148.050 139.200 ;
        RECT 152.400 138.600 153.450 142.950 ;
        RECT 146.400 136.350 147.600 137.100 ;
        RECT 152.400 136.350 153.600 138.600 ;
        RECT 155.400 138.450 156.450 163.950 ;
        RECT 161.400 157.050 162.450 190.950 ;
        RECT 173.400 187.050 174.450 209.400 ;
        RECT 178.950 208.800 181.050 210.900 ;
        RECT 188.400 209.400 189.600 211.650 ;
        RECT 194.400 209.400 195.600 211.650 ;
        RECT 181.950 196.950 184.050 199.050 ;
        RECT 172.950 184.950 175.050 187.050 ;
        RECT 175.950 179.100 178.050 181.200 ;
        RECT 182.400 178.050 183.450 196.950 ;
        RECT 184.950 190.950 187.050 193.050 ;
        RECT 185.400 178.050 186.450 190.950 ;
        RECT 188.400 187.050 189.450 209.400 ;
        RECT 187.950 184.950 190.050 187.050 ;
        RECT 194.400 184.050 195.450 209.400 ;
        RECT 203.400 187.050 204.450 244.950 ;
        RECT 208.950 243.600 211.050 245.700 ;
        RECT 215.400 241.050 216.450 265.950 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 224.400 254.400 225.600 256.650 ;
        RECT 217.950 247.950 220.050 250.050 ;
        RECT 205.950 238.950 208.050 241.050 ;
        RECT 214.950 238.950 217.050 241.050 ;
        RECT 206.400 193.050 207.450 238.950 ;
        RECT 211.950 216.000 214.050 220.050 ;
        RECT 218.400 216.600 219.450 247.950 ;
        RECT 224.400 244.050 225.450 254.400 ;
        RECT 230.100 246.600 231.300 266.400 ;
        RECT 238.950 262.950 241.050 265.050 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 233.400 255.450 234.600 256.650 ;
        RECT 233.400 254.400 237.450 255.450 ;
        RECT 229.950 244.500 232.050 246.600 ;
        RECT 223.950 241.950 226.050 244.050 ;
        RECT 226.950 238.950 229.050 241.050 ;
        RECT 227.400 235.050 228.450 238.950 ;
        RECT 226.950 232.950 229.050 235.050 ;
        RECT 226.950 225.300 229.050 227.400 ;
        RECT 227.850 221.700 229.050 225.300 ;
        RECT 226.950 219.600 229.050 221.700 ;
        RECT 232.950 220.950 235.050 223.050 ;
        RECT 212.400 214.200 213.600 216.000 ;
        RECT 218.400 214.200 219.600 216.600 ;
        RECT 211.950 211.800 214.050 213.900 ;
        RECT 214.950 211.800 217.050 213.900 ;
        RECT 217.950 211.800 220.050 213.900 ;
        RECT 223.950 211.950 226.050 214.050 ;
        RECT 215.400 209.400 216.600 211.500 ;
        RECT 224.400 210.000 225.600 211.650 ;
        RECT 215.400 196.050 216.450 209.400 ;
        RECT 223.950 205.950 226.050 210.000 ;
        RECT 227.850 204.600 229.050 219.600 ;
        RECT 226.950 202.500 229.050 204.600 ;
        RECT 233.400 196.050 234.450 220.950 ;
        RECT 236.400 217.050 237.450 254.400 ;
        RECT 239.400 244.050 240.450 262.950 ;
        RECT 245.400 261.600 246.450 271.950 ;
        RECT 245.400 259.350 246.600 261.600 ;
        RECT 244.950 256.950 247.050 259.050 ;
        RECT 247.950 256.950 250.050 259.050 ;
        RECT 248.400 254.400 249.600 256.650 ;
        RECT 254.400 255.450 255.450 292.950 ;
        RECT 257.400 268.050 258.450 298.950 ;
        RECT 266.400 294.600 267.450 304.950 ;
        RECT 272.400 294.600 273.450 319.950 ;
        RECT 275.400 295.050 276.450 331.950 ;
        RECT 281.400 316.050 282.450 358.950 ;
        RECT 286.950 338.100 289.050 340.200 ;
        RECT 287.400 337.350 288.600 338.100 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 289.950 334.950 292.050 337.050 ;
        RECT 290.400 333.900 291.600 334.650 ;
        RECT 289.950 331.800 292.050 333.900 ;
        RECT 292.950 331.950 295.050 334.050 ;
        RECT 293.400 322.050 294.450 331.950 ;
        RECT 292.950 319.950 295.050 322.050 ;
        RECT 280.950 313.950 283.050 316.050 ;
        RECT 277.950 304.950 280.050 307.050 ;
        RECT 266.400 292.200 267.600 294.600 ;
        RECT 272.400 292.200 273.600 294.600 ;
        RECT 274.950 292.950 277.050 295.050 ;
        RECT 262.950 289.800 265.050 291.900 ;
        RECT 265.950 289.800 268.050 291.900 ;
        RECT 268.950 289.800 271.050 291.900 ;
        RECT 271.950 289.800 274.050 291.900 ;
        RECT 263.400 287.400 264.600 289.500 ;
        RECT 269.400 288.750 270.600 289.500 ;
        RECT 263.400 286.050 264.450 287.400 ;
        RECT 268.950 286.650 271.050 288.750 ;
        RECT 274.950 286.650 277.050 288.750 ;
        RECT 263.400 284.400 268.050 286.050 ;
        RECT 264.000 283.950 268.050 284.400 ;
        RECT 275.400 283.050 276.450 286.650 ;
        RECT 278.400 286.050 279.450 304.950 ;
        RECT 286.950 298.950 289.050 301.050 ;
        RECT 287.400 294.600 288.450 298.950 ;
        RECT 287.400 292.200 288.600 294.600 ;
        RECT 293.400 294.450 294.600 294.600 ;
        RECT 296.400 294.450 297.450 367.950 ;
        RECT 299.400 352.050 300.450 373.950 ;
        RECT 307.950 371.100 310.050 373.200 ;
        RECT 322.950 371.100 325.050 373.200 ;
        RECT 329.400 372.600 330.450 376.950 ;
        RECT 341.400 376.050 342.450 406.950 ;
        RECT 347.400 394.050 348.450 410.400 ;
        RECT 353.700 402.600 354.900 422.400 ;
        RECT 364.950 416.100 367.050 418.200 ;
        RECT 358.950 412.950 361.050 415.050 ;
        RECT 359.400 411.900 360.600 412.650 ;
        RECT 365.400 412.050 366.450 416.100 ;
        RECT 358.950 409.800 361.050 411.900 ;
        RECT 364.950 409.950 367.050 412.050 ;
        RECT 352.950 400.500 355.050 402.600 ;
        RECT 368.400 394.050 369.450 443.400 ;
        RECT 379.950 438.600 381.150 453.600 ;
        RECT 400.950 449.100 403.050 451.200 ;
        RECT 401.400 448.350 402.600 449.100 ;
        RECT 382.950 445.950 385.050 448.050 ;
        RECT 394.950 445.950 397.050 448.050 ;
        RECT 400.950 445.950 403.050 448.050 ;
        RECT 383.400 444.900 384.600 445.650 ;
        RECT 382.950 442.800 385.050 444.900 ;
        RECT 395.400 443.400 396.600 445.650 ;
        RECT 407.400 445.050 408.450 463.950 ;
        RECT 413.400 450.600 414.450 469.950 ;
        RECT 431.400 466.050 432.450 502.950 ;
        RECT 439.950 495.000 442.050 499.050 ;
        RECT 440.400 493.500 441.600 495.000 ;
        RECT 445.950 494.250 448.050 496.350 ;
        RECT 452.400 495.450 453.450 508.950 ;
        RECT 457.950 500.400 460.050 502.500 ;
        RECT 455.400 495.450 456.600 495.600 ;
        RECT 452.400 494.400 456.600 495.450 ;
        RECT 446.400 493.500 447.600 494.250 ;
        RECT 455.400 493.350 456.600 494.400 ;
        RECT 436.950 491.100 439.050 493.200 ;
        RECT 439.950 491.100 442.050 493.200 ;
        RECT 442.950 491.100 445.050 493.200 ;
        RECT 445.950 491.100 448.050 493.200 ;
        RECT 454.950 490.950 457.050 493.050 ;
        RECT 437.400 488.400 438.600 490.800 ;
        RECT 443.400 489.000 444.600 490.800 ;
        RECT 437.400 475.050 438.450 488.400 ;
        RECT 442.950 484.950 445.050 489.000 ;
        RECT 458.850 485.400 460.050 500.400 ;
        RECT 457.950 483.300 460.050 485.400 ;
        RECT 458.850 479.700 460.050 483.300 ;
        RECT 457.950 477.600 460.050 479.700 ;
        RECT 436.950 472.950 439.050 475.050 ;
        RECT 457.950 472.950 460.050 475.050 ;
        RECT 430.950 463.950 433.050 466.050 ;
        RECT 445.950 454.950 448.050 457.050 ;
        RECT 442.950 451.950 445.050 454.050 ;
        RECT 413.400 448.200 414.600 450.600 ;
        RECT 436.950 448.950 439.050 451.050 ;
        RECT 437.400 448.200 438.600 448.950 ;
        RECT 412.950 445.800 415.050 447.900 ;
        RECT 415.950 445.800 418.050 447.900 ;
        RECT 418.950 445.800 421.050 447.900 ;
        RECT 430.950 445.800 433.050 447.900 ;
        RECT 433.950 445.800 436.050 447.900 ;
        RECT 436.950 445.800 439.050 447.900 ;
        RECT 383.400 441.450 384.450 442.800 ;
        RECT 383.400 440.400 387.450 441.450 ;
        RECT 379.950 436.500 382.050 438.600 ;
        RECT 373.950 422.400 376.050 424.500 ;
        RECT 373.950 407.400 375.150 422.400 ;
        RECT 386.400 420.450 387.450 440.400 ;
        RECT 395.400 439.050 396.450 443.400 ;
        RECT 406.950 442.950 409.050 445.050 ;
        RECT 416.400 443.400 417.600 445.500 ;
        RECT 394.950 436.950 397.050 439.050 ;
        RECT 388.950 424.950 391.050 427.050 ;
        RECT 395.400 426.450 396.450 436.950 ;
        RECT 395.400 425.400 399.450 426.450 ;
        RECT 389.400 421.200 390.450 424.950 ;
        RECT 383.400 419.400 387.450 420.450 ;
        RECT 376.950 416.100 379.050 418.200 ;
        RECT 377.400 415.350 378.600 416.100 ;
        RECT 376.950 412.950 379.050 415.050 ;
        RECT 373.950 405.300 376.050 407.400 ;
        RECT 373.950 401.700 375.150 405.300 ;
        RECT 373.950 399.600 376.050 401.700 ;
        RECT 383.400 397.050 384.450 419.400 ;
        RECT 388.950 419.100 391.050 421.200 ;
        RECT 388.950 415.950 391.050 418.050 ;
        RECT 389.400 415.350 390.600 415.950 ;
        RECT 388.950 412.950 391.050 415.050 ;
        RECT 391.950 412.950 394.050 415.050 ;
        RECT 392.400 411.900 393.600 412.650 ;
        RECT 391.950 411.450 394.050 411.900 ;
        RECT 391.950 410.400 396.450 411.450 ;
        RECT 391.950 409.800 394.050 410.400 ;
        RECT 391.950 406.650 394.050 408.750 ;
        RECT 382.950 394.950 385.050 397.050 ;
        RECT 346.950 391.950 349.050 394.050 ;
        RECT 367.950 391.950 370.050 394.050 ;
        RECT 343.950 376.950 346.050 379.050 ;
        RECT 376.950 376.950 379.050 379.050 ;
        RECT 340.950 373.950 343.050 376.050 ;
        RECT 308.400 370.350 309.600 371.100 ;
        RECT 323.400 370.350 324.600 371.100 ;
        RECT 329.400 370.350 330.600 372.600 ;
        RECT 334.800 371.100 336.900 373.200 ;
        RECT 337.950 371.100 340.050 373.200 ;
        RECT 344.400 372.600 345.450 376.950 ;
        RECT 304.950 367.950 307.050 370.050 ;
        RECT 307.950 367.950 310.050 370.050 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 322.950 367.950 325.050 370.050 ;
        RECT 325.950 367.950 328.050 370.050 ;
        RECT 328.950 367.950 331.050 370.050 ;
        RECT 305.400 365.400 306.600 367.650 ;
        RECT 311.400 366.900 312.600 367.650 ;
        RECT 305.400 361.050 306.450 365.400 ;
        RECT 310.950 364.800 313.050 366.900 ;
        RECT 320.400 365.400 321.600 367.650 ;
        RECT 326.400 365.400 327.600 367.650 ;
        RECT 335.400 367.050 336.450 371.100 ;
        RECT 304.950 358.950 307.050 361.050 ;
        RECT 301.950 352.950 304.050 355.050 ;
        RECT 298.950 349.950 301.050 352.050 ;
        RECT 302.400 340.050 303.450 352.950 ;
        RECT 313.950 349.950 316.050 352.050 ;
        RECT 298.950 337.950 301.050 340.050 ;
        RECT 301.950 337.950 304.050 340.050 ;
        RECT 307.950 338.250 310.050 340.350 ;
        RECT 314.400 340.050 315.450 349.950 ;
        RECT 320.400 349.050 321.450 365.400 ;
        RECT 326.400 355.050 327.450 365.400 ;
        RECT 334.950 364.950 337.050 367.050 ;
        RECT 325.950 352.950 328.050 355.050 ;
        RECT 319.950 346.950 322.050 349.050 ;
        RECT 334.950 343.950 337.050 346.050 ;
        RECT 299.400 322.050 300.450 337.950 ;
        RECT 308.400 337.500 309.600 338.250 ;
        RECT 313.950 337.950 316.050 340.050 ;
        RECT 322.950 338.250 325.050 340.350 ;
        RECT 323.400 337.500 324.600 338.250 ;
        RECT 331.950 337.950 334.050 340.050 ;
        RECT 335.400 339.450 336.450 343.950 ;
        RECT 338.400 343.050 339.450 371.100 ;
        RECT 344.400 370.350 345.600 372.600 ;
        RECT 349.950 371.100 352.050 373.200 ;
        RECT 364.950 371.100 367.050 373.200 ;
        RECT 370.950 372.000 373.050 376.050 ;
        RECT 350.400 370.350 351.600 371.100 ;
        RECT 365.400 370.350 366.600 371.100 ;
        RECT 371.400 370.350 372.600 372.000 ;
        RECT 343.950 367.950 346.050 370.050 ;
        RECT 346.950 367.950 349.050 370.050 ;
        RECT 349.950 367.950 352.050 370.050 ;
        RECT 352.950 367.950 355.050 370.050 ;
        RECT 361.950 367.950 364.050 370.050 ;
        RECT 364.950 367.950 367.050 370.050 ;
        RECT 367.950 367.950 370.050 370.050 ;
        RECT 370.950 367.950 373.050 370.050 ;
        RECT 347.400 365.400 348.600 367.650 ;
        RECT 353.400 366.900 354.600 367.650 ;
        RECT 362.400 366.900 363.600 367.650 ;
        RECT 337.950 340.950 340.050 343.050 ;
        RECT 338.400 339.450 339.600 339.600 ;
        RECT 335.400 338.400 339.600 339.450 ;
        RECT 304.950 335.100 307.050 337.200 ;
        RECT 307.950 335.100 310.050 337.200 ;
        RECT 310.950 335.100 313.050 337.200 ;
        RECT 319.950 335.100 322.050 337.200 ;
        RECT 322.950 335.100 325.050 337.200 ;
        RECT 325.950 335.100 328.050 337.200 ;
        RECT 305.400 334.050 306.600 334.800 ;
        RECT 304.950 331.950 307.050 334.050 ;
        RECT 311.400 332.400 312.600 334.800 ;
        RECT 298.950 319.950 301.050 322.050 ;
        RECT 311.400 316.050 312.450 332.400 ;
        RECT 316.950 331.950 319.050 334.050 ;
        RECT 320.400 332.400 321.600 334.800 ;
        RECT 326.400 332.400 327.600 334.800 ;
        RECT 310.950 313.950 313.050 316.050 ;
        RECT 301.950 304.950 304.050 307.050 ;
        RECT 293.400 293.400 297.450 294.450 ;
        RECT 302.400 294.600 303.450 304.950 ;
        RECT 317.400 298.050 318.450 331.950 ;
        RECT 320.400 328.050 321.450 332.400 ;
        RECT 319.950 325.950 322.050 328.050 ;
        RECT 326.400 322.050 327.450 332.400 ;
        RECT 332.400 325.050 333.450 337.950 ;
        RECT 338.400 337.350 339.600 338.400 ;
        RECT 337.950 334.950 340.050 337.050 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 341.400 333.900 342.600 334.650 ;
        RECT 340.950 331.800 343.050 333.900 ;
        RECT 331.950 322.950 334.050 325.050 ;
        RECT 325.950 319.950 328.050 322.050 ;
        RECT 316.950 295.950 319.050 298.050 ;
        RECT 293.400 292.200 294.600 293.400 ;
        RECT 302.400 292.200 303.600 294.600 ;
        RECT 307.950 292.950 310.050 295.050 ;
        RECT 313.950 292.950 316.050 295.050 ;
        RECT 308.400 292.200 309.600 292.950 ;
        RECT 283.950 289.800 286.050 291.900 ;
        RECT 286.950 289.800 289.050 291.900 ;
        RECT 289.950 289.800 292.050 291.900 ;
        RECT 292.950 289.800 295.050 291.900 ;
        RECT 301.950 289.800 304.050 291.900 ;
        RECT 304.950 289.800 307.050 291.900 ;
        RECT 307.950 289.800 310.050 291.900 ;
        RECT 280.950 286.950 283.050 289.050 ;
        RECT 284.400 288.000 285.600 289.500 ;
        RECT 277.950 283.950 280.050 286.050 ;
        RECT 274.950 280.950 277.050 283.050 ;
        RECT 265.950 274.950 268.050 277.050 ;
        RECT 262.950 271.950 265.050 274.050 ;
        RECT 256.950 265.950 259.050 268.050 ;
        RECT 263.400 265.050 264.450 271.950 ;
        RECT 262.950 262.950 265.050 265.050 ;
        RECT 266.400 261.600 267.450 274.950 ;
        RECT 266.400 259.500 267.600 261.600 ;
        RECT 259.950 257.100 262.050 259.200 ;
        RECT 265.950 257.100 268.050 259.200 ;
        RECT 268.950 257.100 271.050 259.200 ;
        RECT 260.400 256.050 261.600 256.800 ;
        RECT 269.400 256.050 270.600 256.800 ;
        RECT 275.400 256.050 276.450 280.950 ;
        RECT 277.950 265.950 280.050 268.050 ;
        RECT 259.950 255.450 262.050 256.050 ;
        RECT 254.400 254.400 258.450 255.450 ;
        RECT 248.400 244.050 249.450 254.400 ;
        RECT 238.950 241.950 241.050 244.050 ;
        RECT 247.950 241.950 250.050 244.050 ;
        RECT 247.950 224.400 250.050 226.500 ;
        RECT 241.950 220.950 244.050 223.050 ;
        RECT 235.950 214.950 238.050 217.050 ;
        RECT 242.400 216.600 243.450 220.950 ;
        RECT 242.400 214.350 243.600 216.600 ;
        RECT 241.950 211.950 244.050 214.050 ;
        RECT 248.100 204.600 249.300 224.400 ;
        RECT 250.950 215.100 253.050 217.200 ;
        RECT 251.400 214.350 252.600 215.100 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 253.950 208.950 256.050 211.050 ;
        RECT 247.950 202.500 250.050 204.600 ;
        RECT 214.950 193.950 217.050 196.050 ;
        RECT 232.950 193.950 235.050 196.050 ;
        RECT 205.950 190.950 208.050 193.050 ;
        RECT 193.950 181.950 196.050 184.050 ;
        RECT 196.950 183.000 199.050 187.050 ;
        RECT 202.950 184.950 205.050 187.050 ;
        RECT 208.950 183.000 211.050 187.050 ;
        RECT 215.400 184.050 216.450 193.950 ;
        RECT 235.950 190.950 238.050 193.050 ;
        RECT 217.950 184.950 220.050 187.050 ;
        RECT 197.400 181.350 198.600 183.000 ;
        RECT 209.400 181.500 210.600 183.000 ;
        RECT 214.950 181.950 217.050 184.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 205.950 179.100 208.050 181.200 ;
        RECT 208.950 179.100 211.050 181.200 ;
        RECT 211.950 179.100 214.050 181.200 ;
        RECT 178.950 175.950 181.050 178.050 ;
        RECT 181.950 175.950 184.050 178.050 ;
        RECT 184.950 175.950 187.050 178.050 ;
        RECT 191.400 177.900 192.600 178.650 ;
        RECT 206.400 178.050 207.600 178.800 ;
        RECT 212.400 178.050 213.600 178.800 ;
        RECT 160.950 154.950 163.050 157.050 ;
        RECT 163.950 146.400 166.050 148.500 ;
        RECT 160.950 138.450 163.050 139.200 ;
        RECT 155.400 137.400 163.050 138.450 ;
        RECT 160.950 137.100 163.050 137.400 ;
        RECT 161.400 136.350 162.600 137.100 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 148.950 133.950 151.050 136.050 ;
        RECT 151.950 133.950 154.050 136.050 ;
        RECT 160.950 133.950 163.050 136.050 ;
        RECT 143.400 132.900 144.600 133.650 ;
        RECT 149.400 132.900 150.600 133.650 ;
        RECT 137.400 131.400 141.450 132.450 ;
        RECT 121.950 130.950 126.000 131.400 ;
        RECT 133.950 127.950 139.050 130.050 ;
        RECT 133.950 124.800 136.050 126.900 ;
        RECT 140.400 126.450 141.450 131.400 ;
        RECT 142.950 130.800 145.050 132.900 ;
        RECT 148.950 130.800 151.050 132.900 ;
        RECT 157.950 130.950 160.050 133.050 ;
        RECT 137.400 125.400 141.450 126.450 ;
        RECT 127.950 121.950 130.050 124.050 ;
        RECT 119.400 103.500 120.600 105.600 ;
        RECT 106.950 101.100 109.050 103.200 ;
        RECT 115.950 101.100 118.050 103.200 ;
        RECT 118.950 101.100 121.050 103.200 ;
        RECT 121.950 101.100 124.050 103.200 ;
        RECT 107.400 99.900 108.600 101.100 ;
        RECT 106.950 97.800 109.050 99.900 ;
        RECT 116.400 98.400 117.600 100.800 ;
        RECT 122.400 98.400 123.600 100.800 ;
        RECT 128.400 100.050 129.450 121.950 ;
        RECT 134.400 118.050 135.450 124.800 ;
        RECT 133.950 115.950 136.050 118.050 ;
        RECT 137.400 105.600 138.450 125.400 ;
        RECT 158.400 115.050 159.450 130.950 ;
        RECT 164.700 126.600 165.900 146.400 ;
        RECT 169.950 138.000 172.050 142.050 ;
        RECT 170.400 136.350 171.600 138.000 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 163.950 124.500 166.050 126.600 ;
        RECT 179.400 118.050 180.450 175.950 ;
        RECT 190.950 175.800 193.050 177.900 ;
        RECT 205.950 175.950 208.050 178.050 ;
        RECT 211.950 175.950 214.050 178.050 ;
        RECT 218.400 175.050 219.450 184.950 ;
        RECT 220.950 181.950 223.050 184.050 ;
        RECT 229.950 182.100 232.050 184.200 ;
        RECT 236.400 183.600 237.450 190.950 ;
        RECT 238.950 187.950 241.050 190.050 ;
        RECT 244.950 188.400 247.050 190.500 ;
        RECT 239.400 184.050 240.450 187.950 ;
        RECT 217.950 172.950 220.050 175.050 ;
        RECT 221.400 172.050 222.450 181.950 ;
        RECT 230.400 181.350 231.600 182.100 ;
        RECT 236.400 181.350 237.600 183.600 ;
        RECT 238.950 181.950 241.050 184.050 ;
        RECT 226.950 178.950 229.050 181.050 ;
        RECT 229.950 178.950 232.050 181.050 ;
        RECT 232.950 178.950 235.050 181.050 ;
        RECT 235.950 178.950 238.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 227.400 177.900 228.600 178.650 ;
        RECT 226.950 175.800 229.050 177.900 ;
        RECT 233.400 177.000 234.600 178.650 ;
        RECT 242.400 177.900 243.600 178.650 ;
        RECT 232.950 172.950 235.050 177.000 ;
        RECT 241.950 175.800 244.050 177.900 ;
        RECT 220.950 169.950 223.050 172.050 ;
        RECT 229.950 171.450 232.050 172.050 ;
        RECT 235.950 171.450 238.050 172.050 ;
        RECT 229.950 170.400 238.050 171.450 ;
        RECT 229.950 169.950 232.050 170.400 ;
        RECT 235.950 169.950 238.050 170.400 ;
        RECT 245.700 168.600 246.900 188.400 ;
        RECT 254.400 186.450 255.450 208.950 ;
        RECT 257.400 208.050 258.450 254.400 ;
        RECT 259.950 254.400 264.450 255.450 ;
        RECT 259.950 253.950 262.050 254.400 ;
        RECT 259.950 244.950 262.050 247.050 ;
        RECT 256.950 205.950 259.050 208.050 ;
        RECT 256.950 186.450 259.050 187.050 ;
        RECT 254.400 185.400 259.050 186.450 ;
        RECT 256.950 184.950 259.050 185.400 ;
        RECT 257.400 181.050 258.450 184.950 ;
        RECT 250.950 178.950 253.050 181.050 ;
        RECT 256.950 178.950 259.050 181.050 ;
        RECT 251.400 176.400 252.600 178.650 ;
        RECT 251.400 172.050 252.450 176.400 ;
        RECT 250.950 169.950 253.050 172.050 ;
        RECT 244.950 166.500 247.050 168.600 ;
        RECT 184.950 147.300 187.050 149.400 ;
        RECT 232.950 148.950 235.050 151.050 ;
        RECT 184.950 143.700 186.150 147.300 ;
        RECT 223.950 145.950 226.050 148.050 ;
        RECT 184.950 141.600 187.050 143.700 ;
        RECT 208.950 142.950 211.050 145.050 ;
        RECT 220.950 142.950 223.050 145.050 ;
        RECT 184.950 126.600 186.150 141.600 ;
        RECT 209.400 139.050 210.450 142.950 ;
        RECT 193.950 136.950 196.050 139.050 ;
        RECT 199.950 136.950 202.050 139.050 ;
        RECT 205.950 136.950 208.050 139.050 ;
        RECT 208.950 136.950 211.050 139.050 ;
        RECT 211.950 136.950 214.050 139.050 ;
        RECT 221.400 138.600 222.450 142.950 ;
        RECT 224.400 142.050 225.450 145.950 ;
        RECT 223.950 139.950 226.050 142.050 ;
        RECT 187.950 133.950 190.050 136.050 ;
        RECT 188.400 132.900 189.600 133.650 ;
        RECT 194.400 132.900 195.450 136.950 ;
        RECT 200.400 136.200 201.600 136.950 ;
        RECT 206.400 136.200 207.600 136.950 ;
        RECT 199.950 133.800 202.050 135.900 ;
        RECT 202.950 133.800 205.050 135.900 ;
        RECT 205.950 133.800 208.050 135.900 ;
        RECT 187.950 130.800 190.050 132.900 ;
        RECT 193.950 130.800 196.050 132.900 ;
        RECT 203.400 132.750 204.600 133.500 ;
        RECT 184.950 124.500 187.050 126.600 ;
        RECT 194.400 121.050 195.450 130.800 ;
        RECT 202.950 130.650 205.050 132.750 ;
        RECT 208.950 127.950 211.050 133.050 ;
        RECT 193.950 118.950 196.050 121.050 ;
        RECT 178.950 115.950 181.050 118.050 ;
        RECT 157.950 112.950 160.050 115.050 ;
        RECT 163.950 112.950 166.050 115.050 ;
        RECT 151.950 110.400 154.050 112.500 ;
        RECT 137.400 103.500 138.600 105.600 ;
        RECT 133.950 101.100 136.050 103.200 ;
        RECT 136.950 101.100 139.050 103.200 ;
        RECT 139.950 101.100 142.050 103.200 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 79.950 91.950 82.050 94.050 ;
        RECT 94.800 92.400 96.900 94.500 ;
        RECT 103.800 92.700 105.900 94.800 ;
        RECT 116.400 94.050 117.450 98.400 ;
        RECT 115.950 91.950 118.050 94.050 ;
        RECT 37.950 59.100 40.050 61.200 ;
        RECT 38.400 58.350 39.600 59.100 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 44.100 48.600 45.300 68.400 ;
        RECT 61.950 67.950 64.050 70.050 ;
        RECT 46.950 60.000 49.050 64.050 ;
        RECT 62.400 60.600 63.450 67.950 ;
        RECT 47.400 58.350 48.600 60.000 ;
        RECT 62.400 58.350 63.600 60.600 ;
        RECT 67.950 59.100 70.050 61.200 ;
        RECT 73.950 59.100 76.050 61.200 ;
        RECT 80.400 60.600 81.450 91.950 ;
        RECT 122.400 85.050 123.450 98.400 ;
        RECT 127.950 97.950 130.050 100.050 ;
        RECT 134.400 99.450 135.600 100.800 ;
        RECT 140.400 100.050 141.600 100.800 ;
        RECT 131.400 98.400 135.600 99.450 ;
        RECT 131.400 94.050 132.450 98.400 ;
        RECT 139.950 97.950 142.050 100.050 ;
        RECT 149.400 98.400 150.600 100.650 ;
        RECT 149.400 94.050 150.450 98.400 ;
        RECT 130.950 91.950 133.050 94.050 ;
        RECT 148.950 91.950 151.050 94.050 ;
        RECT 121.950 82.950 124.050 85.050 ;
        RECT 97.950 69.300 100.050 71.400 ;
        RECT 98.850 65.700 100.050 69.300 ;
        RECT 118.950 68.400 121.050 70.500 ;
        RECT 97.950 63.600 100.050 65.700 ;
        RECT 68.400 58.350 69.600 59.100 ;
        RECT 46.950 55.950 49.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 59.400 54.000 60.600 55.650 ;
        RECT 65.400 54.900 66.600 55.650 ;
        RECT 74.400 55.050 75.450 59.100 ;
        RECT 80.400 58.200 81.600 60.600 ;
        RECT 85.950 58.950 88.050 61.050 ;
        RECT 86.400 58.200 87.600 58.950 ;
        RECT 79.950 55.800 82.050 57.900 ;
        RECT 82.950 55.800 85.050 57.900 ;
        RECT 85.950 55.800 88.050 57.900 ;
        RECT 94.950 55.950 97.050 58.050 ;
        RECT 58.950 49.950 61.050 54.000 ;
        RECT 64.950 52.800 67.050 54.900 ;
        RECT 73.950 52.950 76.050 55.050 ;
        RECT 83.400 54.750 84.600 55.500 ;
        RECT 95.400 54.900 96.600 55.650 ;
        RECT 82.950 52.650 85.050 54.750 ;
        RECT 94.950 52.800 97.050 54.900 ;
        RECT 43.950 46.500 46.050 48.600 ;
        RECT 43.950 32.400 46.050 34.500 ;
        RECT 37.950 22.950 40.050 25.050 ;
        RECT 38.400 21.900 39.600 22.650 ;
        RECT 28.950 19.800 31.050 21.900 ;
        RECT 37.950 19.800 40.050 21.900 ;
        RECT 22.950 15.300 25.050 17.400 ;
        RECT 23.850 11.700 25.050 15.300 ;
        RECT 29.400 13.050 30.450 19.800 ;
        RECT 22.950 9.600 25.050 11.700 ;
        RECT 28.950 10.950 31.050 13.050 ;
        RECT 44.100 12.600 45.300 32.400 ;
        RECT 52.950 31.950 55.050 34.050 ;
        RECT 46.950 22.950 49.050 25.050 ;
        RECT 47.400 21.000 48.600 22.650 ;
        RECT 53.400 22.050 54.450 31.950 ;
        RECT 59.400 28.200 60.450 49.950 ;
        RECT 98.850 48.600 100.050 63.600 ;
        RECT 103.950 61.950 106.050 64.050 ;
        RECT 97.950 46.500 100.050 48.600 ;
        RECT 64.950 31.950 67.050 34.050 ;
        RECT 97.950 32.400 100.050 34.500 ;
        RECT 58.950 26.100 61.050 28.200 ;
        RECT 65.400 27.600 66.450 31.950 ;
        RECT 59.400 25.350 60.600 26.100 ;
        RECT 65.400 25.350 66.600 27.600 ;
        RECT 73.950 25.950 76.050 28.050 ;
        RECT 82.950 26.250 85.050 28.350 ;
        RECT 58.950 22.950 61.050 25.050 ;
        RECT 61.950 22.950 64.050 25.050 ;
        RECT 64.950 22.950 67.050 25.050 ;
        RECT 67.950 22.950 70.050 25.050 ;
        RECT 46.950 16.950 49.050 21.000 ;
        RECT 52.950 19.950 55.050 22.050 ;
        RECT 62.400 20.400 63.600 22.650 ;
        RECT 68.400 21.900 69.600 22.650 ;
        RECT 74.400 21.900 75.450 25.950 ;
        RECT 83.400 25.500 84.600 26.250 ;
        RECT 94.950 26.100 97.050 28.200 ;
        RECT 95.400 25.350 96.600 26.100 ;
        RECT 79.950 23.100 82.050 25.200 ;
        RECT 82.950 23.100 85.050 25.200 ;
        RECT 85.950 23.100 88.050 25.200 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 80.400 22.050 81.600 22.800 ;
        RECT 86.400 22.050 87.600 22.800 ;
        RECT 62.400 13.050 63.450 20.400 ;
        RECT 67.950 19.800 70.050 21.900 ;
        RECT 73.950 19.800 76.050 21.900 ;
        RECT 79.950 19.950 82.050 22.050 ;
        RECT 85.950 19.950 88.050 22.050 ;
        RECT 98.850 17.400 100.050 32.400 ;
        RECT 104.400 19.050 105.450 61.950 ;
        RECT 106.950 59.100 109.050 61.200 ;
        RECT 112.950 59.100 115.050 61.200 ;
        RECT 107.400 46.050 108.450 59.100 ;
        RECT 113.400 58.350 114.600 59.100 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 119.100 48.600 120.300 68.400 ;
        RECT 121.950 60.000 124.050 64.050 ;
        RECT 122.400 58.350 123.600 60.000 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 127.950 49.950 130.050 54.900 ;
        RECT 131.400 52.050 132.450 91.950 ;
        RECT 152.700 90.600 153.900 110.400 ;
        RECT 157.950 100.950 160.050 103.050 ;
        RECT 158.400 99.900 159.600 100.650 ;
        RECT 157.950 97.800 160.050 99.900 ;
        RECT 164.400 94.050 165.450 112.950 ;
        RECT 166.950 109.950 169.050 112.050 ;
        RECT 172.950 110.400 175.050 112.500 ;
        RECT 212.400 112.050 213.450 136.950 ;
        RECT 221.400 136.350 222.600 138.600 ;
        RECT 226.950 137.100 229.050 139.200 ;
        RECT 227.400 136.350 228.600 137.100 ;
        RECT 217.950 133.950 220.050 136.050 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 218.400 131.400 219.600 133.650 ;
        RECT 224.400 132.900 225.600 133.650 ;
        RECT 218.400 127.050 219.450 131.400 ;
        RECT 223.950 130.800 226.050 132.900 ;
        RECT 220.950 127.950 223.050 130.050 ;
        RECT 217.950 124.950 220.050 127.050 ;
        RECT 221.400 124.050 222.450 127.950 ;
        RECT 233.400 127.050 234.450 148.950 ;
        RECT 241.950 145.950 244.050 148.050 ;
        RECT 247.950 145.950 250.050 148.050 ;
        RECT 242.400 138.600 243.450 145.950 ;
        RECT 248.400 138.600 249.450 145.950 ;
        RECT 256.950 139.950 259.050 142.050 ;
        RECT 242.400 136.350 243.600 138.600 ;
        RECT 248.400 136.350 249.600 138.600 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 250.950 133.950 253.050 136.050 ;
        RECT 245.400 131.400 246.600 133.650 ;
        RECT 251.400 131.400 252.600 133.650 ;
        RECT 232.950 124.950 235.050 127.050 ;
        RECT 220.950 121.950 223.050 124.050 ;
        RECT 167.400 99.900 168.450 109.950 ;
        RECT 166.950 97.800 169.050 99.900 ;
        RECT 172.950 95.400 174.150 110.400 ;
        RECT 187.950 109.950 190.050 112.050 ;
        RECT 211.950 109.950 214.050 112.050 ;
        RECT 175.950 104.100 178.050 106.200 ;
        RECT 181.950 104.100 184.050 106.200 ;
        RECT 188.400 105.600 189.450 109.950 ;
        RECT 176.400 103.350 177.600 104.100 ;
        RECT 175.950 100.950 178.050 103.050 ;
        RECT 163.950 91.950 166.050 94.050 ;
        RECT 172.950 93.300 175.050 95.400 ;
        RECT 182.400 94.050 183.450 104.100 ;
        RECT 188.400 103.350 189.600 105.600 ;
        RECT 193.950 105.000 196.050 109.050 ;
        RECT 194.400 103.350 195.600 105.000 ;
        RECT 202.950 103.950 205.050 106.050 ;
        RECT 211.950 104.250 214.050 106.350 ;
        RECT 221.400 105.450 222.450 121.950 ;
        RECT 226.950 110.400 229.050 112.500 ;
        RECT 224.400 105.450 225.600 105.600 ;
        RECT 221.400 104.400 225.600 105.450 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 193.950 100.950 196.050 103.050 ;
        RECT 196.950 100.950 199.050 103.050 ;
        RECT 191.400 99.900 192.600 100.650 ;
        RECT 197.400 99.900 198.600 100.650 ;
        RECT 203.400 99.900 204.450 103.950 ;
        RECT 212.400 103.500 213.600 104.250 ;
        RECT 224.400 103.350 225.600 104.400 ;
        RECT 208.950 101.100 211.050 103.200 ;
        RECT 211.950 101.100 214.050 103.200 ;
        RECT 214.950 101.100 217.050 103.200 ;
        RECT 223.950 100.950 226.050 103.050 ;
        RECT 190.950 97.800 193.050 99.900 ;
        RECT 196.950 97.800 199.050 99.900 ;
        RECT 202.950 97.800 205.050 99.900 ;
        RECT 209.400 98.400 210.600 100.800 ;
        RECT 215.400 100.050 216.600 100.800 ;
        RECT 209.400 94.050 210.450 98.400 ;
        RECT 214.950 97.950 217.050 100.050 ;
        RECT 227.850 95.400 229.050 110.400 ;
        RECT 151.950 88.500 154.050 90.600 ;
        RECT 148.950 82.950 151.050 85.050 ;
        RECT 139.950 59.100 142.050 61.200 ;
        RECT 140.400 58.350 141.600 59.100 ;
        RECT 136.950 55.950 139.050 58.050 ;
        RECT 139.950 55.950 142.050 58.050 ;
        RECT 142.950 55.950 145.050 58.050 ;
        RECT 137.400 54.000 138.600 55.650 ;
        RECT 130.950 49.950 133.050 52.050 ;
        RECT 136.950 49.950 139.050 54.000 ;
        RECT 143.400 53.400 144.600 55.650 ;
        RECT 149.400 55.050 150.450 82.950 ;
        RECT 164.400 64.050 165.450 91.950 ;
        RECT 172.950 89.700 174.150 93.300 ;
        RECT 181.950 91.950 184.050 94.050 ;
        RECT 208.950 91.950 211.050 94.050 ;
        RECT 226.950 93.300 229.050 95.400 ;
        RECT 227.850 89.700 229.050 93.300 ;
        RECT 172.950 87.600 175.050 89.700 ;
        RECT 226.950 87.600 229.050 89.700 ;
        RECT 187.950 79.950 190.050 82.050 ;
        RECT 166.950 73.950 169.050 76.050 ;
        RECT 184.950 73.950 187.050 76.050 ;
        RECT 163.950 61.950 166.050 64.050 ;
        RECT 157.950 58.950 160.050 61.050 ;
        RECT 164.400 60.450 165.600 60.600 ;
        RECT 167.400 60.450 168.450 73.950 ;
        RECT 172.950 68.400 175.050 70.500 ;
        RECT 164.400 59.400 168.450 60.450 ;
        RECT 169.950 60.000 172.050 64.050 ;
        RECT 158.400 58.200 159.600 58.950 ;
        RECT 164.400 58.200 165.600 59.400 ;
        RECT 170.400 58.350 171.600 60.000 ;
        RECT 154.950 55.800 157.050 57.900 ;
        RECT 157.950 55.800 160.050 57.900 ;
        RECT 160.950 55.800 163.050 57.900 ;
        RECT 163.950 55.800 166.050 57.900 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 118.950 46.500 121.050 48.600 ;
        RECT 106.950 43.950 109.050 46.050 ;
        RECT 118.950 32.400 121.050 34.500 ;
        RECT 106.950 25.950 109.050 28.050 ;
        RECT 107.400 21.900 108.450 25.950 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 113.400 21.900 114.600 22.650 ;
        RECT 106.950 19.800 109.050 21.900 ;
        RECT 112.950 19.800 115.050 21.900 ;
        RECT 97.950 15.300 100.050 17.400 ;
        RECT 103.950 16.950 106.050 19.050 ;
        RECT 43.950 10.500 46.050 12.600 ;
        RECT 61.950 10.950 64.050 13.050 ;
        RECT 98.850 11.700 100.050 15.300 ;
        RECT 119.100 12.600 120.300 32.400 ;
        RECT 143.400 31.050 144.450 53.400 ;
        RECT 148.950 52.950 151.050 55.050 ;
        RECT 155.400 53.400 156.600 55.500 ;
        RECT 161.400 53.400 162.600 55.500 ;
        RECT 155.400 46.050 156.450 53.400 ;
        RECT 161.400 49.050 162.450 53.400 ;
        RECT 160.950 46.950 163.050 49.050 ;
        RECT 173.700 48.600 174.900 68.400 ;
        RECT 178.950 60.000 181.050 64.050 ;
        RECT 179.400 58.350 180.600 60.000 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 172.950 46.500 175.050 48.600 ;
        RECT 154.950 43.950 157.050 46.050 ;
        RECT 160.950 34.950 163.050 37.050 ;
        RECT 127.950 25.950 130.050 28.050 ;
        RECT 136.950 26.100 139.050 28.200 ;
        RECT 142.950 27.000 145.050 31.050 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 122.400 21.000 123.600 22.650 ;
        RECT 128.400 22.050 129.450 25.950 ;
        RECT 137.400 25.350 138.600 26.100 ;
        RECT 143.400 25.350 144.600 27.000 ;
        RECT 148.950 25.950 151.050 28.050 ;
        RECT 154.950 26.250 157.050 28.350 ;
        RECT 161.400 27.600 162.450 34.950 ;
        RECT 172.950 32.400 175.050 34.500 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 139.950 22.950 142.050 25.050 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 121.950 16.950 124.050 21.000 ;
        RECT 127.950 19.950 130.050 22.050 ;
        RECT 140.400 20.400 141.600 22.650 ;
        RECT 149.400 22.050 150.450 25.950 ;
        RECT 155.400 25.500 156.600 26.250 ;
        RECT 161.400 25.500 162.600 27.600 ;
        RECT 154.950 23.100 157.050 25.200 ;
        RECT 157.950 23.100 160.050 25.200 ;
        RECT 160.950 23.100 163.050 25.200 ;
        RECT 163.950 23.100 166.050 25.200 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 158.400 22.050 159.600 22.800 ;
        RECT 140.400 19.050 141.450 20.400 ;
        RECT 148.800 19.950 150.900 22.050 ;
        RECT 140.400 17.400 145.050 19.050 ;
        RECT 141.000 16.950 145.050 17.400 ;
        RECT 151.950 16.950 154.050 22.050 ;
        RECT 157.950 19.950 160.050 22.050 ;
        RECT 164.400 20.400 165.600 22.800 ;
        RECT 170.400 21.000 171.600 22.650 ;
        RECT 164.400 13.050 165.450 20.400 ;
        RECT 169.950 16.950 172.050 21.000 ;
        RECT 97.950 9.600 100.050 11.700 ;
        RECT 118.950 10.500 121.050 12.600 ;
        RECT 163.950 10.950 166.050 13.050 ;
        RECT 173.700 12.600 174.900 32.400 ;
        RECT 185.400 31.050 186.450 73.950 ;
        RECT 188.400 49.050 189.450 79.950 ;
        RECT 233.400 76.050 234.450 124.950 ;
        RECT 245.400 118.050 246.450 131.400 ;
        RECT 251.400 124.050 252.450 131.400 ;
        RECT 257.400 127.050 258.450 139.950 ;
        RECT 260.400 139.050 261.450 244.950 ;
        RECT 263.400 217.050 264.450 254.400 ;
        RECT 268.950 253.950 271.050 256.050 ;
        RECT 271.950 253.950 274.050 256.050 ;
        RECT 274.950 253.950 277.050 256.050 ;
        RECT 272.400 229.050 273.450 253.950 ;
        RECT 278.400 244.050 279.450 265.950 ;
        RECT 281.400 262.050 282.450 286.950 ;
        RECT 283.950 283.950 286.050 288.000 ;
        RECT 290.400 287.400 291.600 289.500 ;
        RECT 305.400 287.400 306.600 289.500 ;
        RECT 290.400 283.050 291.450 287.400 ;
        RECT 289.950 280.950 292.050 283.050 ;
        RECT 305.400 274.050 306.450 287.400 ;
        RECT 286.950 271.950 289.050 274.050 ;
        RECT 304.950 271.950 307.050 274.050 ;
        RECT 280.950 259.950 283.050 262.050 ;
        RECT 287.400 261.600 288.450 271.950 ;
        RECT 301.950 265.950 304.050 268.050 ;
        RECT 287.400 259.350 288.600 261.600 ;
        RECT 292.950 261.000 295.050 265.050 ;
        RECT 302.400 261.600 303.450 265.950 ;
        RECT 293.400 259.350 294.600 261.000 ;
        RECT 302.400 259.350 303.600 261.600 ;
        RECT 307.950 260.100 310.050 262.200 ;
        RECT 314.400 262.050 315.450 292.950 ;
        RECT 317.400 265.050 318.450 295.950 ;
        RECT 322.950 293.100 325.050 295.200 ;
        RECT 347.400 295.050 348.450 365.400 ;
        RECT 352.950 364.800 355.050 366.900 ;
        RECT 361.950 364.800 364.050 366.900 ;
        RECT 368.400 365.400 369.600 367.650 ;
        RECT 377.400 367.050 378.450 376.950 ;
        RECT 385.950 371.100 388.050 373.200 ;
        RECT 386.400 370.350 387.600 371.100 ;
        RECT 382.950 367.950 385.050 370.050 ;
        RECT 385.950 367.950 388.050 370.050 ;
        RECT 361.950 358.950 364.050 361.050 ;
        RECT 349.950 349.950 352.050 352.050 ;
        RECT 323.400 292.350 324.600 293.100 ;
        RECT 337.950 292.950 340.050 295.050 ;
        RECT 344.400 294.450 345.600 294.600 ;
        RECT 346.950 294.450 349.050 295.050 ;
        RECT 344.400 293.400 349.050 294.450 ;
        RECT 338.400 292.200 339.600 292.950 ;
        RECT 344.400 292.200 345.600 293.400 ;
        RECT 346.950 292.950 349.050 293.400 ;
        RECT 322.950 289.950 325.050 292.050 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 337.950 289.800 340.050 291.900 ;
        RECT 340.950 289.800 343.050 291.900 ;
        RECT 343.950 289.800 346.050 291.900 ;
        RECT 329.400 287.400 330.600 289.650 ;
        RECT 325.950 268.950 328.050 271.050 ;
        RECT 316.950 262.950 319.050 265.050 ;
        RECT 308.400 259.350 309.600 260.100 ;
        RECT 313.950 259.950 316.050 262.050 ;
        RECT 283.950 256.950 286.050 259.050 ;
        RECT 286.950 256.950 289.050 259.050 ;
        RECT 289.950 256.950 292.050 259.050 ;
        RECT 292.950 256.950 295.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 304.950 256.950 307.050 259.050 ;
        RECT 307.950 256.950 310.050 259.050 ;
        RECT 310.950 256.950 313.050 259.050 ;
        RECT 280.950 253.950 283.050 256.050 ;
        RECT 284.400 254.400 285.600 256.650 ;
        RECT 290.400 254.400 291.600 256.650 ;
        RECT 277.950 241.950 280.050 244.050 ;
        RECT 271.950 226.950 274.050 229.050 ;
        RECT 268.800 220.500 270.900 222.600 ;
        RECT 262.950 214.950 265.050 217.050 ;
        RECT 268.950 213.900 269.850 220.500 ;
        RECT 277.800 220.200 279.900 222.300 ;
        RECT 272.400 216.900 273.600 219.600 ;
        RECT 271.650 214.800 273.750 216.900 ;
        RECT 275.700 213.900 277.800 214.200 ;
        RECT 265.950 211.800 268.050 213.900 ;
        RECT 268.950 213.000 277.800 213.900 ;
        RECT 266.400 209.400 267.600 211.800 ;
        RECT 268.950 207.900 269.850 213.000 ;
        RECT 275.700 212.100 277.800 213.000 ;
        RECT 270.750 211.200 272.850 212.100 ;
        RECT 270.750 210.000 277.800 211.200 ;
        RECT 275.700 209.100 277.800 210.000 ;
        RECT 268.200 205.800 270.300 207.900 ;
        RECT 271.650 206.100 273.750 208.200 ;
        RECT 278.700 207.600 279.600 220.200 ;
        RECT 281.400 216.600 282.450 253.950 ;
        RECT 284.400 252.450 285.450 254.400 ;
        RECT 284.400 251.400 288.450 252.450 ;
        RECT 281.400 213.900 282.600 216.600 ;
        RECT 280.950 211.800 283.050 213.900 ;
        RECT 287.400 210.450 288.450 251.400 ;
        RECT 290.400 244.050 291.450 254.400 ;
        RECT 295.950 253.950 298.050 256.050 ;
        RECT 305.400 254.400 306.600 256.650 ;
        RECT 311.400 255.000 312.600 256.650 ;
        RECT 317.400 256.050 318.450 262.950 ;
        RECT 326.400 261.600 327.450 268.950 ;
        RECT 329.400 265.050 330.450 287.400 ;
        RECT 334.950 286.950 337.050 289.050 ;
        RECT 341.400 287.400 342.600 289.500 ;
        RECT 335.400 279.450 336.450 286.950 ;
        RECT 337.950 279.450 340.050 280.050 ;
        RECT 335.400 278.400 340.050 279.450 ;
        RECT 337.950 277.950 340.050 278.400 ;
        RECT 334.950 268.950 337.050 271.050 ;
        RECT 328.950 262.950 331.050 265.050 ;
        RECT 326.400 259.500 327.600 261.600 ;
        RECT 322.950 257.100 325.050 259.200 ;
        RECT 325.950 257.100 328.050 259.200 ;
        RECT 328.950 257.100 331.050 259.200 ;
        RECT 323.400 256.050 324.600 256.800 ;
        RECT 329.400 256.050 330.600 256.800 ;
        RECT 289.950 241.950 292.050 244.050 ;
        RECT 296.400 241.050 297.450 253.950 ;
        RECT 305.400 252.450 306.450 254.400 ;
        RECT 302.400 251.400 306.450 252.450 ;
        RECT 295.950 238.950 298.050 241.050 ;
        RECT 292.950 232.950 295.050 235.050 ;
        RECT 293.400 216.600 294.450 232.950 ;
        RECT 302.400 229.050 303.450 251.400 ;
        RECT 310.950 250.950 313.050 255.000 ;
        RECT 316.950 253.950 319.050 256.050 ;
        RECT 322.950 253.950 325.050 256.050 ;
        RECT 328.950 253.950 331.050 256.050 ;
        RECT 331.950 253.950 334.050 256.050 ;
        RECT 322.950 252.450 325.050 252.900 ;
        RECT 329.400 252.450 330.450 253.950 ;
        RECT 322.950 251.400 330.450 252.450 ;
        RECT 322.950 250.800 325.050 251.400 ;
        RECT 332.400 250.050 333.450 253.950 ;
        RECT 331.950 247.950 334.050 250.050 ;
        RECT 322.950 241.950 325.050 244.050 ;
        RECT 323.400 235.050 324.450 241.950 ;
        RECT 304.950 232.950 307.050 235.050 ;
        RECT 322.950 232.950 325.050 235.050 ;
        RECT 301.950 226.950 304.050 229.050 ;
        RECT 298.950 220.950 301.050 223.050 ;
        RECT 299.400 216.600 300.450 220.950 ;
        RECT 293.400 214.200 294.600 216.600 ;
        RECT 299.400 214.200 300.600 216.600 ;
        RECT 292.950 211.800 295.050 213.900 ;
        RECT 295.950 211.800 298.050 213.900 ;
        RECT 298.950 211.800 301.050 213.900 ;
        RECT 296.400 210.750 297.600 211.500 ;
        RECT 287.400 209.400 291.450 210.450 ;
        RECT 272.400 203.400 273.600 206.100 ;
        RECT 278.250 205.500 280.350 207.600 ;
        RECT 265.950 188.400 268.050 190.500 ;
        RECT 265.950 173.400 267.150 188.400 ;
        RECT 268.950 182.100 271.050 184.200 ;
        RECT 272.400 183.450 273.450 203.400 ;
        RECT 277.950 190.950 280.050 193.050 ;
        RECT 278.400 184.050 279.450 190.950 ;
        RECT 283.950 187.950 286.050 190.050 ;
        RECT 272.400 182.400 276.450 183.450 ;
        RECT 269.400 181.350 270.600 182.100 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 265.950 171.300 268.050 173.400 ;
        RECT 265.950 167.700 267.150 171.300 ;
        RECT 265.950 165.600 268.050 167.700 ;
        RECT 275.400 142.050 276.450 182.400 ;
        RECT 277.950 181.950 280.050 184.050 ;
        RECT 284.400 183.600 285.450 187.950 ;
        RECT 290.400 184.050 291.450 209.400 ;
        RECT 295.950 208.650 298.050 210.750 ;
        RECT 292.950 205.950 295.050 208.050 ;
        RECT 284.400 181.500 285.600 183.600 ;
        RECT 289.950 181.950 292.050 184.050 ;
        RECT 280.950 179.100 283.050 181.200 ;
        RECT 283.950 179.100 286.050 181.200 ;
        RECT 286.950 179.100 289.050 181.200 ;
        RECT 281.400 178.050 282.600 178.800 ;
        RECT 287.400 178.050 288.600 178.800 ;
        RECT 293.400 178.050 294.450 205.950 ;
        RECT 305.400 193.050 306.450 232.950 ;
        RECT 322.950 226.950 325.050 229.050 ;
        RECT 316.950 223.950 319.050 226.050 ;
        RECT 310.950 215.100 313.050 217.200 ;
        RECT 317.400 216.600 318.450 223.950 ;
        RECT 323.400 217.050 324.450 226.950 ;
        RECT 328.950 224.400 331.050 226.500 ;
        RECT 335.400 226.050 336.450 268.950 ;
        RECT 338.400 261.450 339.450 277.950 ;
        RECT 341.400 265.050 342.450 287.400 ;
        RECT 346.950 286.950 349.050 289.050 ;
        RECT 340.950 262.950 343.050 265.050 ;
        RECT 347.400 261.600 348.450 286.950 ;
        RECT 341.400 261.450 342.600 261.600 ;
        RECT 338.400 260.400 342.600 261.450 ;
        RECT 341.400 259.350 342.600 260.400 ;
        RECT 347.400 259.350 348.600 261.600 ;
        RECT 350.400 261.450 351.450 349.950 ;
        RECT 355.950 343.950 358.050 346.050 ;
        RECT 356.400 339.600 357.450 343.950 ;
        RECT 362.400 339.600 363.450 358.950 ;
        RECT 368.400 346.050 369.450 365.400 ;
        RECT 376.950 364.950 379.050 367.050 ;
        RECT 383.400 366.000 384.600 367.650 ;
        RECT 382.950 361.950 385.050 366.000 ;
        RECT 382.950 352.950 385.050 355.050 ;
        RECT 376.950 349.950 379.050 352.050 ;
        RECT 367.950 343.950 370.050 346.050 ;
        RECT 367.950 339.600 372.000 340.050 ;
        RECT 377.400 339.600 378.450 349.950 ;
        RECT 383.400 340.050 384.450 352.950 ;
        RECT 385.950 343.950 388.050 346.050 ;
        RECT 356.400 337.350 357.600 339.600 ;
        RECT 362.400 337.350 363.600 339.600 ;
        RECT 367.950 337.950 372.600 339.600 ;
        RECT 371.400 337.350 372.600 337.950 ;
        RECT 377.400 337.350 378.600 339.600 ;
        RECT 382.950 337.950 385.050 340.050 ;
        RECT 386.400 337.050 387.450 343.950 ;
        RECT 392.400 340.200 393.450 406.650 ;
        RECT 395.400 355.050 396.450 410.400 ;
        RECT 398.400 409.050 399.450 425.400 ;
        RECT 412.950 424.950 415.050 427.050 ;
        RECT 400.950 421.950 403.050 424.050 ;
        RECT 401.400 418.050 402.450 421.950 ;
        RECT 413.400 421.050 414.450 424.950 ;
        RECT 416.400 424.050 417.450 443.400 ;
        RECT 427.950 442.950 430.050 445.050 ;
        RECT 434.400 444.750 435.600 445.500 ;
        RECT 443.400 445.050 444.450 451.950 ;
        RECT 428.400 439.050 429.450 442.950 ;
        RECT 433.950 442.650 436.050 444.750 ;
        RECT 442.800 442.950 444.900 445.050 ;
        RECT 446.400 444.900 447.450 454.950 ;
        RECT 451.950 450.000 454.050 454.050 ;
        RECT 458.400 451.200 459.450 472.950 ;
        RECT 452.400 448.350 453.600 450.000 ;
        RECT 457.950 449.100 460.050 451.200 ;
        RECT 464.400 450.450 465.450 529.950 ;
        RECT 469.950 516.600 471.150 531.600 ;
        RECT 476.400 529.050 477.450 535.950 ;
        RECT 475.950 526.950 478.050 529.050 ;
        RECT 472.950 523.950 475.050 526.050 ;
        RECT 473.400 522.900 474.600 523.650 ;
        RECT 472.950 520.800 475.050 522.900 ;
        RECT 469.950 514.500 472.050 516.600 ;
        RECT 479.400 508.050 480.450 566.400 ;
        RECT 485.400 562.050 486.450 566.400 ;
        RECT 484.950 559.950 487.050 562.050 ;
        RECT 485.400 532.050 486.450 559.950 ;
        RECT 487.950 547.950 490.050 550.050 ;
        RECT 484.950 529.950 487.050 532.050 ;
        RECT 488.400 528.450 489.450 547.950 ;
        RECT 491.400 538.050 492.450 572.400 ;
        RECT 500.400 571.350 501.600 573.600 ;
        RECT 505.950 572.100 508.050 574.200 ;
        RECT 506.400 571.350 507.600 572.100 ;
        RECT 496.950 568.950 499.050 571.050 ;
        RECT 499.950 568.950 502.050 571.050 ;
        RECT 502.950 568.950 505.050 571.050 ;
        RECT 505.950 568.950 508.050 571.050 ;
        RECT 497.400 567.900 498.600 568.650 ;
        RECT 496.950 565.800 499.050 567.900 ;
        RECT 503.400 566.400 504.600 568.650 ;
        RECT 503.400 559.050 504.450 566.400 ;
        RECT 512.400 559.050 513.450 589.950 ;
        RECT 515.400 574.050 516.450 589.950 ;
        RECT 521.400 587.400 522.450 589.950 ;
        RECT 527.400 583.050 528.450 589.950 ;
        RECT 530.400 589.050 531.450 599.400 ;
        RECT 532.950 595.950 535.050 598.050 ;
        RECT 529.950 586.950 532.050 589.050 ;
        RECT 533.400 586.050 534.450 595.950 ;
        RECT 532.950 583.950 535.050 586.050 ;
        RECT 536.400 583.050 537.450 599.400 ;
        RECT 545.400 595.050 546.450 607.800 ;
        RECT 554.400 606.600 555.450 634.950 ;
        RECT 560.400 619.050 561.450 637.950 ;
        RECT 563.400 619.050 564.450 644.400 ;
        RECT 565.950 643.950 568.050 646.050 ;
        RECT 568.950 643.950 571.050 646.050 ;
        RECT 559.800 616.950 561.900 619.050 ;
        RECT 562.950 616.950 565.050 619.050 ;
        RECT 566.400 616.050 567.450 643.950 ;
        RECT 575.400 637.050 576.450 661.950 ;
        RECT 578.400 652.050 579.450 677.400 ;
        RECT 584.400 652.050 585.450 700.950 ;
        RECT 595.950 682.950 598.050 685.050 ;
        RECT 596.400 682.200 597.600 682.950 ;
        RECT 589.950 679.800 592.050 681.900 ;
        RECT 592.950 679.800 595.050 681.900 ;
        RECT 595.950 679.800 598.050 681.900 ;
        RECT 593.400 677.400 594.600 679.500 ;
        RECT 593.400 661.050 594.450 677.400 ;
        RECT 598.950 676.950 601.050 679.050 ;
        RECT 592.950 658.950 595.050 661.050 ;
        RECT 599.400 658.050 600.450 676.950 ;
        RECT 602.400 676.050 603.450 715.950 ;
        RECT 605.400 685.050 606.450 722.400 ;
        RECT 614.400 722.400 615.600 724.650 ;
        RECT 620.400 722.400 621.600 724.650 ;
        RECT 614.400 720.450 615.450 722.400 ;
        RECT 611.400 719.400 615.450 720.450 ;
        RECT 611.400 697.050 612.450 719.400 ;
        RECT 620.400 718.050 621.450 722.400 ;
        RECT 626.400 721.050 627.450 728.400 ;
        RECT 632.400 727.350 633.600 729.600 ;
        RECT 638.400 727.350 639.600 729.600 ;
        RECT 649.950 728.100 652.050 730.200 ;
        RECT 631.950 724.950 634.050 727.050 ;
        RECT 634.950 724.950 637.050 727.050 ;
        RECT 637.950 724.950 640.050 727.050 ;
        RECT 640.950 724.950 643.050 727.050 ;
        RECT 635.400 722.400 636.600 724.650 ;
        RECT 641.400 723.900 642.600 724.650 ;
        RECT 650.400 724.050 651.450 728.100 ;
        RECT 656.400 727.200 657.600 729.600 ;
        RECT 655.950 725.100 658.050 727.200 ;
        RECT 658.950 726.900 659.850 732.300 ;
        RECT 661.950 730.800 664.050 732.900 ;
        RECT 665.700 729.900 667.800 731.700 ;
        RECT 660.750 728.700 669.300 729.900 ;
        RECT 660.750 727.800 662.850 728.700 ;
        RECT 658.950 725.700 665.850 726.900 ;
        RECT 625.950 718.950 628.050 721.050 ;
        RECT 619.950 715.950 622.050 718.050 ;
        RECT 631.950 703.950 634.050 706.050 ;
        RECT 610.950 694.950 613.050 697.050 ;
        RECT 626.100 688.200 628.200 690.300 ;
        RECT 604.950 682.950 607.050 685.050 ;
        RECT 613.950 682.950 616.050 685.050 ;
        RECT 622.950 684.000 625.050 688.050 ;
        RECT 614.400 682.200 615.600 682.950 ;
        RECT 623.400 681.900 624.600 684.000 ;
        RECT 607.950 679.800 610.050 681.900 ;
        RECT 610.950 679.800 613.050 681.900 ;
        RECT 613.950 679.800 616.050 681.900 ;
        RECT 622.950 679.800 625.050 681.900 ;
        RECT 604.950 676.950 607.050 679.050 ;
        RECT 611.400 678.000 612.600 679.500 ;
        RECT 601.950 673.950 604.050 676.050 ;
        RECT 605.400 667.050 606.450 676.950 ;
        RECT 610.950 673.950 613.050 678.000 ;
        RECT 626.400 675.600 627.300 688.200 ;
        RECT 632.400 687.600 633.450 703.950 ;
        RECT 635.400 703.050 636.450 722.400 ;
        RECT 640.800 721.800 642.900 723.900 ;
        RECT 649.950 721.950 652.050 724.050 ;
        RECT 639.000 720.750 642.000 721.050 ;
        RECT 637.950 718.950 643.050 720.750 ;
        RECT 637.950 718.650 640.050 718.950 ;
        RECT 640.950 718.650 643.050 718.950 ;
        RECT 650.400 718.050 651.450 721.950 ;
        RECT 652.950 718.950 655.050 721.050 ;
        RECT 649.950 715.950 652.050 718.050 ;
        RECT 653.400 715.050 654.450 718.950 ;
        RECT 658.950 718.500 660.150 725.700 ;
        RECT 661.950 722.100 664.050 724.200 ;
        RECT 664.950 723.300 665.850 725.700 ;
        RECT 662.400 719.400 663.600 722.100 ;
        RECT 664.950 721.200 667.050 723.300 ;
        RECT 668.400 719.700 669.300 728.700 ;
        RECT 682.950 728.100 685.050 730.200 ;
        RECT 692.400 729.450 693.450 754.950 ;
        RECT 698.400 748.050 699.450 755.400 ;
        RECT 703.950 754.800 706.050 756.900 ;
        RECT 715.950 754.800 718.050 756.900 ;
        RECT 722.400 756.000 723.600 757.650 ;
        RECT 700.950 751.950 703.050 754.050 ;
        RECT 721.950 751.950 724.050 756.000 ;
        RECT 727.950 751.950 730.050 757.050 ;
        RECT 734.400 756.750 735.600 757.500 ;
        RECT 733.950 754.650 736.050 756.750 ;
        RECT 739.950 754.950 742.050 757.050 ;
        RECT 697.950 745.950 700.050 748.050 ;
        RECT 701.400 736.050 702.450 751.950 ;
        RECT 718.950 745.950 721.050 748.050 ;
        RECT 700.950 733.950 703.050 736.050 ;
        RECT 701.400 729.600 702.450 733.950 ;
        RECT 692.400 728.400 696.450 729.450 ;
        RECT 683.400 727.350 684.600 728.100 ;
        RECT 670.950 725.100 673.050 727.200 ;
        RECT 671.400 723.900 672.600 725.100 ;
        RECT 679.950 724.950 682.050 727.050 ;
        RECT 682.950 724.950 685.050 727.050 ;
        RECT 688.950 724.950 691.050 727.050 ;
        RECT 680.400 723.900 681.600 724.650 ;
        RECT 670.950 721.800 673.050 723.900 ;
        RECT 679.950 721.800 682.050 723.900 ;
        RECT 689.400 722.400 690.600 724.650 ;
        RECT 658.500 716.400 660.600 718.500 ;
        RECT 668.100 717.600 670.200 719.700 ;
        RECT 680.400 715.050 681.450 721.800 ;
        RECT 652.950 712.950 655.050 715.050 ;
        RECT 679.950 712.950 682.050 715.050 ;
        RECT 689.400 712.050 690.450 722.400 ;
        RECT 688.950 709.950 691.050 712.050 ;
        RECT 695.400 709.050 696.450 728.400 ;
        RECT 701.400 727.350 702.600 729.600 ;
        RECT 706.950 728.100 709.050 730.200 ;
        RECT 707.400 727.350 708.600 728.100 ;
        RECT 715.950 727.950 718.050 730.050 ;
        RECT 700.950 724.950 703.050 727.050 ;
        RECT 703.950 724.950 706.050 727.050 ;
        RECT 706.950 724.950 709.050 727.050 ;
        RECT 709.950 724.950 712.050 727.050 ;
        RECT 704.400 722.400 705.600 724.650 ;
        RECT 710.400 723.900 711.600 724.650 ;
        RECT 658.950 706.950 661.050 709.050 ;
        RECT 664.950 706.950 667.050 709.050 ;
        RECT 694.950 706.950 697.050 709.050 ;
        RECT 659.400 703.050 660.450 706.950 ;
        RECT 634.950 700.950 637.050 703.050 ;
        RECT 652.950 700.950 655.050 703.050 ;
        RECT 658.950 700.950 661.050 703.050 ;
        RECT 635.100 688.500 637.200 690.600 ;
        RECT 632.400 684.900 633.600 687.600 ;
        RECT 632.250 682.800 634.350 684.900 ;
        RECT 628.200 681.900 630.300 682.200 ;
        RECT 636.150 681.900 637.050 688.500 ;
        RECT 653.400 685.200 654.450 700.950 ;
        RECT 652.950 683.100 655.050 685.200 ;
        RECT 658.950 683.100 661.050 685.200 ;
        RECT 653.400 682.350 654.600 683.100 ;
        RECT 659.400 682.350 660.600 683.100 ;
        RECT 628.200 681.000 637.050 681.900 ;
        RECT 628.200 680.100 630.300 681.000 ;
        RECT 633.150 679.200 635.250 680.100 ;
        RECT 628.200 678.000 635.250 679.200 ;
        RECT 628.200 677.100 630.450 678.000 ;
        RECT 625.650 673.500 627.750 675.600 ;
        RECT 629.400 673.050 630.450 677.100 ;
        RECT 632.250 674.100 634.350 676.200 ;
        RECT 636.150 675.900 637.050 681.000 ;
        RECT 637.950 679.800 640.050 681.900 ;
        RECT 649.950 679.950 652.050 682.050 ;
        RECT 652.950 679.950 655.050 682.050 ;
        RECT 655.950 679.950 658.050 682.050 ;
        RECT 658.950 679.950 661.050 682.050 ;
        RECT 638.400 677.400 639.600 679.800 ;
        RECT 646.950 676.950 649.050 679.050 ;
        RECT 650.400 677.400 651.600 679.650 ;
        RECT 656.400 677.400 657.600 679.650 ;
        RECT 628.950 670.950 631.050 673.050 ;
        RECT 632.400 671.400 633.600 674.100 ;
        RECT 635.700 673.800 637.800 675.900 ;
        RECT 640.950 670.950 643.050 673.050 ;
        RECT 604.950 664.950 607.050 667.050 ;
        RECT 605.400 661.050 606.450 664.950 ;
        RECT 629.400 661.050 630.450 670.950 ;
        RECT 631.950 661.950 634.050 664.050 ;
        RECT 604.950 658.950 607.050 661.050 ;
        RECT 610.950 658.950 613.050 661.050 ;
        RECT 628.950 658.950 631.050 661.050 ;
        RECT 598.950 655.950 601.050 658.050 ;
        RECT 577.950 649.950 580.050 652.050 ;
        RECT 583.950 649.950 586.050 652.050 ;
        RECT 604.950 651.000 607.050 655.050 ;
        RECT 611.400 651.600 612.450 658.950 ;
        RECT 613.950 652.950 619.050 655.050 ;
        RECT 622.950 654.450 627.000 655.050 ;
        RECT 622.950 652.950 627.450 654.450 ;
        RECT 605.400 649.500 606.600 651.000 ;
        RECT 611.400 649.500 612.600 651.600 ;
        RECT 616.950 649.800 619.050 651.900 ;
        RECT 626.400 651.600 627.450 652.950 ;
        RECT 632.400 651.600 633.450 661.950 ;
        RECT 580.950 647.100 583.050 649.200 ;
        RECT 586.950 647.100 589.050 649.200 ;
        RECT 589.950 647.100 592.050 649.200 ;
        RECT 601.950 647.100 604.050 649.200 ;
        RECT 604.950 647.100 607.050 649.200 ;
        RECT 607.950 647.100 610.050 649.200 ;
        RECT 610.950 647.100 613.050 649.200 ;
        RECT 581.400 646.050 582.600 646.800 ;
        RECT 590.400 646.050 591.600 646.800 ;
        RECT 602.400 646.050 603.600 646.800 ;
        RECT 580.950 643.950 583.050 646.050 ;
        RECT 586.950 643.950 589.050 646.050 ;
        RECT 590.400 644.400 595.050 646.050 ;
        RECT 591.000 643.950 595.050 644.400 ;
        RECT 601.950 643.950 604.050 646.050 ;
        RECT 608.400 644.400 609.600 646.800 ;
        RECT 574.950 634.950 577.050 637.050 ;
        RECT 571.950 628.950 574.050 631.050 ;
        RECT 564.000 615.900 567.450 616.050 ;
        RECT 562.950 614.400 567.450 615.900 ;
        RECT 562.950 613.950 567.000 614.400 ;
        RECT 562.950 613.800 565.050 613.950 ;
        RECT 556.950 607.950 559.050 613.050 ;
        RECT 572.400 612.450 573.450 628.950 ;
        RECT 581.400 628.050 582.450 643.950 ;
        RECT 587.400 640.050 588.450 643.950 ;
        RECT 586.950 637.950 589.050 640.050 ;
        RECT 592.950 631.950 595.050 634.050 ;
        RECT 580.950 625.950 583.050 628.050 ;
        RECT 577.950 622.950 580.050 625.050 ;
        RECT 572.400 611.400 576.450 612.450 ;
        RECT 568.950 607.950 574.050 610.050 ;
        RECT 575.400 607.050 576.450 611.400 ;
        RECT 554.400 604.350 555.600 606.600 ;
        RECT 574.950 604.950 577.050 607.050 ;
        RECT 550.950 601.950 553.050 604.050 ;
        RECT 553.950 601.950 556.050 604.050 ;
        RECT 556.950 601.950 559.050 604.050 ;
        RECT 568.950 601.800 571.050 603.900 ;
        RECT 571.950 601.800 574.050 603.900 ;
        RECT 551.400 601.050 552.600 601.650 ;
        RECT 547.950 599.400 552.600 601.050 ;
        RECT 557.400 600.000 558.600 601.650 ;
        RECT 572.400 600.000 573.600 601.500 ;
        RECT 547.950 598.950 552.450 599.400 ;
        RECT 544.950 592.950 547.050 595.050 ;
        RECT 538.950 586.950 541.050 589.050 ;
        RECT 526.950 580.950 529.050 583.050 ;
        RECT 535.950 580.950 538.050 583.050 ;
        RECT 517.950 577.950 520.050 580.050 ;
        RECT 529.950 577.950 532.050 580.050 ;
        RECT 518.400 574.350 519.450 577.950 ;
        RECT 514.800 571.950 516.900 574.050 ;
        RECT 517.950 572.250 520.050 574.350 ;
        RECT 530.400 574.200 531.450 577.950 ;
        RECT 539.400 577.050 540.450 586.950 ;
        RECT 547.950 583.950 550.050 586.050 ;
        RECT 538.950 574.950 541.050 577.050 ;
        RECT 544.950 574.950 547.050 577.050 ;
        RECT 518.400 571.500 519.600 572.250 ;
        RECT 529.950 572.100 532.050 574.200 ;
        RECT 535.950 572.100 538.050 574.200 ;
        RECT 530.400 571.350 531.600 572.100 ;
        RECT 536.400 571.350 537.600 572.100 ;
        RECT 517.950 569.100 520.050 571.200 ;
        RECT 520.950 569.100 523.050 571.200 ;
        RECT 529.950 568.950 532.050 571.050 ;
        RECT 532.950 568.950 535.050 571.050 ;
        RECT 535.950 568.950 538.050 571.050 ;
        RECT 538.950 568.950 541.050 571.050 ;
        RECT 526.950 565.950 529.050 568.050 ;
        RECT 533.400 566.400 534.600 568.650 ;
        RECT 539.400 567.900 540.600 568.650 ;
        RECT 545.400 567.900 546.450 574.950 ;
        RECT 548.400 574.050 549.450 583.950 ;
        RECT 551.400 580.050 552.450 598.950 ;
        RECT 556.950 595.950 559.050 600.000 ;
        RECT 571.950 595.950 574.050 600.000 ;
        RECT 574.950 598.950 577.050 601.050 ;
        RECT 550.950 577.950 553.050 580.050 ;
        RECT 552.000 576.900 555.000 577.050 ;
        RECT 550.950 576.450 555.000 576.900 ;
        RECT 572.400 576.450 573.450 595.950 ;
        RECT 575.400 583.050 576.450 598.950 ;
        RECT 578.400 589.050 579.450 622.950 ;
        RECT 580.950 610.950 583.050 613.050 ;
        RECT 581.400 607.050 582.450 610.950 ;
        RECT 580.950 604.950 583.050 607.050 ;
        RECT 583.950 601.800 586.050 603.900 ;
        RECT 586.950 601.800 589.050 603.900 ;
        RECT 587.400 599.400 588.600 601.500 ;
        RECT 580.950 595.950 583.050 598.050 ;
        RECT 577.950 586.950 580.050 589.050 ;
        RECT 574.950 580.950 577.050 583.050 ;
        RECT 550.950 574.950 555.450 576.450 ;
        RECT 572.400 575.400 576.450 576.450 ;
        RECT 550.950 574.800 553.050 574.950 ;
        RECT 547.950 571.950 550.050 574.050 ;
        RECT 554.400 573.600 555.450 574.950 ;
        RECT 575.400 574.200 576.450 575.400 ;
        RECT 554.400 571.500 555.600 573.600 ;
        RECT 568.950 572.100 571.050 574.200 ;
        RECT 574.950 572.100 577.050 574.200 ;
        RECT 569.400 571.350 570.600 572.100 ;
        RECT 575.400 571.350 576.600 572.100 ;
        RECT 550.950 569.100 553.050 571.200 ;
        RECT 553.950 569.100 556.050 571.200 ;
        RECT 556.950 569.100 559.050 571.200 ;
        RECT 581.400 571.050 582.450 595.950 ;
        RECT 587.400 592.050 588.450 599.400 ;
        RECT 593.400 592.050 594.450 631.950 ;
        RECT 595.950 625.950 598.050 628.050 ;
        RECT 596.400 610.050 597.450 625.950 ;
        RECT 598.950 622.950 601.050 625.050 ;
        RECT 595.950 607.950 598.050 610.050 ;
        RECT 599.400 607.050 600.450 622.950 ;
        RECT 608.400 616.050 609.450 644.400 ;
        RECT 610.950 643.950 616.050 646.050 ;
        RECT 613.950 622.950 616.050 625.050 ;
        RECT 607.950 613.950 610.050 616.050 ;
        RECT 598.950 604.950 601.050 607.050 ;
        RECT 607.950 604.950 610.050 610.050 ;
        RECT 614.400 606.450 615.450 622.950 ;
        RECT 617.400 610.050 618.450 649.800 ;
        RECT 626.400 649.500 627.600 651.600 ;
        RECT 632.400 649.500 633.600 651.600 ;
        RECT 622.950 647.100 625.050 649.200 ;
        RECT 625.950 647.100 628.050 649.200 ;
        RECT 628.950 647.100 631.050 649.200 ;
        RECT 631.950 647.100 634.050 649.200 ;
        RECT 634.950 647.100 637.050 649.200 ;
        RECT 623.400 646.050 624.600 646.800 ;
        RECT 622.950 643.950 625.050 646.050 ;
        RECT 629.400 645.450 630.600 646.800 ;
        RECT 635.400 646.050 636.600 646.800 ;
        RECT 641.400 646.050 642.450 670.950 ;
        RECT 647.400 664.050 648.450 676.950 ;
        RECT 646.950 661.950 649.050 664.050 ;
        RECT 650.400 655.050 651.450 677.400 ;
        RECT 656.400 673.050 657.450 677.400 ;
        RECT 655.950 670.950 658.050 673.050 ;
        RECT 655.950 664.950 658.050 667.050 ;
        RECT 643.950 652.950 646.050 655.050 ;
        RECT 629.400 644.400 633.450 645.450 ;
        RECT 628.950 640.950 631.050 643.050 ;
        RECT 629.400 625.050 630.450 640.950 ;
        RECT 632.400 640.050 633.450 644.400 ;
        RECT 634.950 643.950 637.050 646.050 ;
        RECT 640.950 643.950 643.050 646.050 ;
        RECT 631.950 637.950 634.050 640.050 ;
        RECT 628.950 622.950 631.050 625.050 ;
        RECT 619.950 616.950 622.050 619.050 ;
        RECT 616.950 607.950 619.050 610.050 ;
        RECT 620.400 607.050 621.450 616.950 ;
        RECT 644.400 612.450 645.450 652.950 ;
        RECT 649.950 651.000 652.050 655.050 ;
        RECT 656.400 651.600 657.450 664.950 ;
        RECT 665.400 655.050 666.450 706.950 ;
        RECT 704.400 706.050 705.450 722.400 ;
        RECT 709.950 721.800 712.050 723.900 ;
        RECT 712.950 709.950 715.050 712.050 ;
        RECT 703.950 703.950 706.050 706.050 ;
        RECT 679.950 691.950 682.050 697.050 ;
        RECT 673.800 687.300 675.900 689.400 ;
        RECT 683.400 688.500 685.500 690.600 ;
        RECT 670.950 682.950 673.050 685.050 ;
        RECT 671.400 681.900 672.600 682.950 ;
        RECT 670.950 679.800 673.050 681.900 ;
        RECT 674.700 678.300 675.600 687.300 ;
        RECT 676.950 683.700 679.050 685.800 ;
        RECT 680.400 684.900 681.600 687.600 ;
        RECT 678.150 681.300 679.050 683.700 ;
        RECT 679.950 682.800 682.050 684.900 ;
        RECT 683.850 681.300 685.050 688.500 ;
        RECT 691.950 682.950 694.050 685.050 ;
        RECT 697.950 682.950 700.050 685.050 ;
        RECT 703.950 682.950 706.050 685.050 ;
        RECT 678.150 680.100 685.050 681.300 ;
        RECT 681.150 678.300 683.250 679.200 ;
        RECT 674.700 677.100 683.250 678.300 ;
        RECT 670.950 673.800 673.050 675.900 ;
        RECT 676.200 675.300 678.300 677.100 ;
        RECT 679.950 674.100 682.050 676.200 ;
        RECT 684.150 674.700 685.050 680.100 ;
        RECT 685.950 679.800 688.050 681.900 ;
        RECT 686.400 677.400 687.600 679.800 ;
        RECT 664.950 652.950 667.050 655.050 ;
        RECT 671.400 651.600 672.450 673.800 ;
        RECT 680.400 671.400 681.600 674.100 ;
        RECT 683.400 672.600 685.500 674.700 ;
        RECT 692.400 664.050 693.450 682.950 ;
        RECT 698.400 682.200 699.600 682.950 ;
        RECT 704.400 682.200 705.600 682.950 ;
        RECT 697.950 679.800 700.050 681.900 ;
        RECT 700.950 679.800 703.050 681.900 ;
        RECT 703.950 679.800 706.050 681.900 ;
        RECT 706.950 679.800 709.050 681.900 ;
        RECT 694.950 676.950 697.050 679.050 ;
        RECT 701.400 677.400 702.600 679.500 ;
        RECT 707.400 677.400 708.600 679.500 ;
        RECT 691.950 661.950 694.050 664.050 ;
        RECT 695.400 660.450 696.450 676.950 ;
        RECT 701.400 673.050 702.450 677.400 ;
        RECT 700.950 670.950 703.050 673.050 ;
        RECT 707.400 661.050 708.450 677.400 ;
        RECT 713.400 676.050 714.450 709.950 ;
        RECT 716.400 691.050 717.450 727.950 ;
        RECT 719.400 723.900 720.450 745.950 ;
        RECT 734.400 732.450 735.450 754.650 ;
        RECT 736.950 751.950 739.050 754.050 ;
        RECT 731.400 731.400 735.450 732.450 ;
        RECT 724.950 728.250 727.050 730.350 ;
        RECT 731.400 729.600 732.450 731.400 ;
        RECT 737.400 730.050 738.450 751.950 ;
        RECT 740.400 748.050 741.450 754.950 ;
        RECT 743.400 754.050 744.450 796.950 ;
        RECT 746.400 766.050 747.450 800.400 ;
        RECT 751.950 796.950 754.050 801.000 ;
        RECT 767.400 800.400 768.600 802.800 ;
        RECT 773.400 800.400 774.600 802.800 ;
        RECT 785.400 801.000 786.600 802.800 ;
        RECT 791.400 801.450 792.600 802.800 ;
        RECT 800.400 801.900 801.450 814.950 ;
        RECT 802.950 805.950 805.050 808.050 ;
        RECT 811.950 806.100 814.050 808.200 ;
        RECT 817.950 807.000 820.050 811.050 ;
        RECT 826.950 807.000 829.050 811.050 ;
        RECT 767.400 787.050 768.450 800.400 ;
        RECT 766.950 784.950 769.050 787.050 ;
        RECT 773.400 775.050 774.450 800.400 ;
        RECT 784.950 796.950 787.050 801.000 ;
        RECT 788.400 800.400 792.600 801.450 ;
        RECT 775.950 787.950 778.050 790.050 ;
        RECT 772.950 772.950 775.050 775.050 ;
        RECT 745.950 760.950 748.050 766.050 ;
        RECT 748.950 760.950 751.050 763.050 ;
        RECT 754.950 762.000 757.050 766.050 ;
        RECT 749.400 760.200 750.600 760.950 ;
        RECT 755.400 760.200 756.600 762.000 ;
        RECT 763.950 760.950 766.050 763.050 ;
        RECT 769.950 760.950 772.050 763.050 ;
        RECT 776.400 762.600 777.450 787.950 ;
        RECT 784.950 766.950 787.050 769.050 ;
        RECT 748.950 757.800 751.050 759.900 ;
        RECT 751.950 757.800 754.050 759.900 ;
        RECT 754.950 757.800 757.050 759.900 ;
        RECT 757.950 757.800 760.050 759.900 ;
        RECT 752.400 756.000 753.600 757.500 ;
        RECT 758.400 756.750 759.600 757.500 ;
        RECT 742.950 751.950 745.050 754.050 ;
        RECT 751.950 751.950 754.050 756.000 ;
        RECT 757.950 754.650 760.050 756.750 ;
        RECT 764.400 751.050 765.450 760.950 ;
        RECT 770.400 760.200 771.600 760.950 ;
        RECT 776.400 760.200 777.600 762.600 ;
        RECT 769.950 757.800 772.050 759.900 ;
        RECT 772.950 757.800 775.050 759.900 ;
        RECT 775.950 757.800 778.050 759.900 ;
        RECT 778.950 757.800 781.050 759.900 ;
        RECT 766.950 754.950 769.050 757.050 ;
        RECT 773.400 756.750 774.600 757.500 ;
        RECT 779.400 756.750 780.600 757.500 ;
        RECT 748.950 748.950 751.050 751.050 ;
        RECT 763.950 748.950 766.050 751.050 ;
        RECT 739.950 745.950 742.050 748.050 ;
        RECT 739.950 736.950 742.050 739.050 ;
        RECT 740.400 730.050 741.450 736.950 ;
        RECT 742.950 733.950 745.050 736.050 ;
        RECT 725.400 727.500 726.600 728.250 ;
        RECT 731.400 727.500 732.600 729.600 ;
        RECT 736.800 727.950 738.900 730.050 ;
        RECT 739.950 727.950 742.050 730.050 ;
        RECT 743.400 729.600 744.450 733.950 ;
        RECT 749.400 730.200 750.450 748.950 ;
        RECT 757.950 733.950 760.050 736.050 ;
        RECT 743.400 727.350 744.600 729.600 ;
        RECT 748.950 728.100 751.050 730.200 ;
        RECT 749.400 727.350 750.600 728.100 ;
        RECT 724.950 725.100 727.050 727.200 ;
        RECT 727.950 725.100 730.050 727.200 ;
        RECT 730.950 725.100 733.050 727.200 ;
        RECT 733.950 725.100 736.050 727.200 ;
        RECT 742.950 724.950 745.050 727.050 ;
        RECT 745.950 724.950 748.050 727.050 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 751.950 724.950 754.050 727.050 ;
        RECT 718.950 721.800 721.050 723.900 ;
        RECT 724.950 721.950 727.050 724.050 ;
        RECT 728.400 722.400 729.600 724.800 ;
        RECT 734.400 724.050 735.600 724.800 ;
        RECT 721.950 718.950 724.050 721.050 ;
        RECT 722.400 697.050 723.450 718.950 ;
        RECT 725.400 697.050 726.450 721.950 ;
        RECT 728.400 718.050 729.450 722.400 ;
        RECT 733.950 721.950 736.050 724.050 ;
        RECT 746.400 723.900 747.600 724.650 ;
        RECT 745.950 721.800 748.050 723.900 ;
        RECT 752.400 722.400 753.600 724.650 ;
        RECT 746.400 718.050 747.450 721.800 ;
        RECT 727.950 715.950 730.050 718.050 ;
        RECT 745.950 715.950 748.050 718.050 ;
        RECT 752.400 706.050 753.450 722.400 ;
        RECT 758.400 712.050 759.450 733.950 ;
        RECT 767.400 730.350 768.450 754.950 ;
        RECT 772.950 754.650 775.050 756.750 ;
        RECT 778.950 754.650 781.050 756.750 ;
        RECT 781.950 754.950 784.050 757.050 ;
        RECT 772.950 733.950 775.050 736.050 ;
        RECT 766.950 728.250 769.050 730.350 ;
        RECT 773.400 729.600 774.450 733.950 ;
        RECT 782.400 730.050 783.450 754.950 ;
        RECT 785.400 733.050 786.450 766.950 ;
        RECT 788.400 757.050 789.450 800.400 ;
        RECT 799.950 799.800 802.050 801.900 ;
        RECT 800.400 769.050 801.450 799.800 ;
        RECT 803.400 778.050 804.450 805.950 ;
        RECT 812.400 805.350 813.600 806.100 ;
        RECT 818.400 805.350 819.600 807.000 ;
        RECT 827.400 805.350 828.600 807.000 ;
        RECT 832.950 806.100 835.050 808.200 ;
        RECT 833.400 805.350 834.600 806.100 ;
        RECT 841.950 805.950 844.050 808.050 ;
        RECT 808.950 802.950 811.050 805.050 ;
        RECT 811.950 802.950 814.050 805.050 ;
        RECT 814.950 802.950 817.050 805.050 ;
        RECT 817.950 802.950 820.050 805.050 ;
        RECT 826.950 802.950 829.050 805.050 ;
        RECT 829.950 802.950 832.050 805.050 ;
        RECT 832.950 802.950 835.050 805.050 ;
        RECT 835.950 802.950 838.050 805.050 ;
        RECT 809.400 801.900 810.600 802.650 ;
        RECT 815.400 801.900 816.600 802.650 ;
        RECT 830.400 801.900 831.600 802.650 ;
        RECT 808.950 799.800 811.050 801.900 ;
        RECT 814.950 799.800 817.050 801.900 ;
        RECT 829.950 799.800 832.050 801.900 ;
        RECT 836.400 800.400 837.600 802.650 ;
        RECT 836.400 790.050 837.450 800.400 ;
        RECT 835.950 787.950 838.050 790.050 ;
        RECT 802.950 775.950 805.050 778.050 ;
        RECT 826.950 775.950 829.050 778.050 ;
        RECT 811.950 769.950 814.050 772.050 ;
        RECT 823.950 769.950 826.050 772.050 ;
        RECT 799.950 766.950 802.050 769.050 ;
        RECT 795.000 765.600 799.050 766.050 ;
        RECT 794.400 765.000 799.050 765.600 ;
        RECT 793.950 763.950 799.050 765.000 ;
        RECT 793.950 763.050 796.050 763.950 ;
        RECT 793.800 762.000 796.050 763.050 ;
        RECT 793.800 760.950 795.900 762.000 ;
        RECT 796.950 760.800 799.050 762.900 ;
        RECT 802.950 762.000 805.050 766.050 ;
        RECT 812.400 762.600 813.450 769.950 ;
        RECT 817.950 766.950 820.050 769.050 ;
        RECT 818.400 762.600 819.450 766.950 ;
        RECT 797.400 760.200 798.600 760.800 ;
        RECT 803.400 760.200 804.600 762.000 ;
        RECT 812.400 760.200 813.600 762.600 ;
        RECT 818.400 760.200 819.600 762.600 ;
        RECT 820.950 760.950 823.050 766.050 ;
        RECT 793.950 757.800 796.050 759.900 ;
        RECT 796.950 757.800 799.050 759.900 ;
        RECT 799.950 757.800 802.050 759.900 ;
        RECT 802.950 757.800 805.050 759.900 ;
        RECT 811.950 757.800 814.050 759.900 ;
        RECT 814.950 757.800 817.050 759.900 ;
        RECT 817.950 757.800 820.050 759.900 ;
        RECT 787.950 754.950 790.050 757.050 ;
        RECT 794.400 755.400 795.600 757.500 ;
        RECT 800.400 755.400 801.600 757.500 ;
        RECT 815.400 755.400 816.600 757.500 ;
        RECT 787.950 748.950 790.050 751.050 ;
        RECT 784.950 730.950 787.050 733.050 ;
        RECT 767.400 727.500 768.600 728.250 ;
        RECT 773.400 727.500 774.600 729.600 ;
        RECT 781.950 727.950 784.050 730.050 ;
        RECT 788.400 729.600 789.450 748.950 ;
        RECT 794.400 735.450 795.450 755.400 ;
        RECT 800.400 751.050 801.450 755.400 ;
        RECT 799.950 748.950 802.050 751.050 ;
        RECT 815.400 736.050 816.450 755.400 ;
        RECT 824.400 744.450 825.450 769.950 ;
        RECT 827.400 763.050 828.450 775.950 ;
        RECT 826.950 760.950 829.050 763.050 ;
        RECT 829.950 760.950 832.050 763.050 ;
        RECT 835.950 762.000 838.050 766.050 ;
        RECT 842.400 763.050 843.450 805.950 ;
        RECT 862.950 766.950 865.050 769.050 ;
        RECT 830.400 760.200 831.600 760.950 ;
        RECT 836.400 760.200 837.600 762.000 ;
        RECT 841.950 760.950 844.050 763.050 ;
        RECT 853.950 761.100 856.050 763.200 ;
        RECT 854.400 760.350 855.600 761.100 ;
        RECT 829.950 757.800 832.050 759.900 ;
        RECT 832.950 757.800 835.050 759.900 ;
        RECT 835.950 757.800 838.050 759.900 ;
        RECT 838.950 757.800 841.050 759.900 ;
        RECT 850.950 757.950 853.050 760.050 ;
        RECT 853.950 757.950 856.050 760.050 ;
        RECT 826.950 754.950 829.050 757.050 ;
        RECT 833.400 755.400 834.600 757.500 ;
        RECT 839.400 755.400 840.600 757.500 ;
        RECT 827.400 751.050 828.450 754.950 ;
        RECT 833.400 751.050 834.450 755.400 ;
        RECT 826.950 748.950 829.050 751.050 ;
        RECT 832.950 748.950 835.050 751.050 ;
        RECT 824.400 743.400 828.450 744.450 ;
        RECT 823.950 741.450 826.050 742.050 ;
        RECT 818.400 740.400 826.050 741.450 ;
        RECT 794.400 734.400 798.450 735.450 ;
        RECT 788.400 727.500 789.600 729.600 ;
        RECT 793.950 729.000 796.050 733.050 ;
        RECT 797.400 730.050 798.450 734.400 ;
        RECT 799.950 733.950 802.050 736.050 ;
        RECT 814.950 733.950 817.050 736.050 ;
        RECT 794.400 727.500 795.600 729.000 ;
        RECT 796.950 727.950 799.050 730.050 ;
        RECT 763.950 725.100 766.050 727.200 ;
        RECT 766.950 725.100 769.050 727.200 ;
        RECT 769.950 725.100 772.050 727.200 ;
        RECT 772.950 725.100 775.050 727.200 ;
        RECT 764.400 724.050 765.600 724.800 ;
        RECT 763.950 721.950 766.050 724.050 ;
        RECT 770.400 723.000 771.600 724.800 ;
        RECT 769.950 718.950 772.050 723.000 ;
        RECT 772.950 721.950 775.050 724.050 ;
        RECT 778.950 721.950 781.050 727.050 ;
        RECT 784.950 725.100 787.050 727.200 ;
        RECT 787.950 725.100 790.050 727.200 ;
        RECT 790.950 725.100 793.050 727.200 ;
        RECT 793.950 725.100 796.050 727.200 ;
        RECT 785.400 724.050 786.600 724.800 ;
        RECT 791.400 724.050 792.600 724.800 ;
        RECT 784.950 721.950 787.050 724.050 ;
        RECT 790.950 721.950 793.050 724.050 ;
        RECT 757.950 709.950 760.050 712.050 ;
        RECT 773.400 706.050 774.450 721.950 ;
        RECT 800.400 709.050 801.450 733.950 ;
        RECT 802.950 727.950 805.050 730.050 ;
        RECT 811.950 728.100 814.050 730.200 ;
        RECT 818.400 729.600 819.450 740.400 ;
        RECT 823.950 739.950 826.050 740.400 ;
        RECT 820.950 736.950 823.050 739.050 ;
        RECT 821.400 730.050 822.450 736.950 ;
        RECT 823.950 730.950 826.050 733.050 ;
        RECT 799.950 706.950 802.050 709.050 ;
        RECT 751.950 703.950 754.050 706.050 ;
        RECT 772.950 703.950 775.050 706.050 ;
        RECT 799.950 703.800 802.050 705.900 ;
        RECT 793.950 697.950 796.050 700.050 ;
        RECT 721.800 694.950 723.900 697.050 ;
        RECT 724.950 694.950 727.050 697.050 ;
        RECT 769.950 694.950 772.050 697.050 ;
        RECT 715.950 688.950 718.050 691.050 ;
        RECT 716.400 685.050 717.450 688.950 ;
        RECT 715.950 682.950 718.050 685.050 ;
        RECT 718.950 684.000 721.050 688.050 ;
        RECT 725.400 684.600 726.450 694.950 ;
        RECT 742.950 688.950 745.050 691.050 ;
        RECT 736.950 685.950 739.050 688.050 ;
        RECT 719.400 682.200 720.600 684.000 ;
        RECT 725.400 682.200 726.600 684.600 ;
        RECT 718.950 679.800 721.050 681.900 ;
        RECT 721.950 679.800 724.050 681.900 ;
        RECT 724.950 679.800 727.050 681.900 ;
        RECT 727.950 679.800 730.050 681.900 ;
        RECT 722.400 677.400 723.600 679.500 ;
        RECT 728.400 677.400 729.600 679.500 ;
        RECT 712.950 673.950 715.050 676.050 ;
        RECT 718.950 673.950 721.050 676.050 ;
        RECT 712.950 667.950 715.050 670.050 ;
        RECT 692.400 659.400 696.450 660.450 ;
        RECT 650.400 649.350 651.600 651.000 ;
        RECT 656.400 649.350 657.600 651.600 ;
        RECT 671.400 649.500 672.600 651.600 ;
        RECT 685.950 650.250 688.050 652.350 ;
        RECT 692.400 651.600 693.450 659.400 ;
        RECT 686.400 649.500 687.600 650.250 ;
        RECT 692.400 649.500 693.600 651.600 ;
        RECT 695.400 651.450 696.450 659.400 ;
        RECT 706.950 658.950 709.050 661.050 ;
        RECT 695.400 650.400 699.450 651.450 ;
        RECT 649.950 646.950 652.050 649.050 ;
        RECT 652.950 646.950 655.050 649.050 ;
        RECT 655.950 646.950 658.050 649.050 ;
        RECT 661.950 646.950 664.050 649.050 ;
        RECT 667.950 647.100 670.050 649.200 ;
        RECT 670.950 647.100 673.050 649.200 ;
        RECT 673.950 647.100 676.050 649.200 ;
        RECT 682.950 647.100 685.050 649.200 ;
        RECT 685.950 647.100 688.050 649.200 ;
        RECT 688.950 647.100 691.050 649.200 ;
        RECT 691.950 647.100 694.050 649.200 ;
        RECT 653.400 644.400 654.600 646.650 ;
        RECT 653.400 637.050 654.450 644.400 ;
        RECT 655.950 640.950 658.050 643.050 ;
        RECT 652.950 634.950 655.050 637.050 ;
        RECT 649.950 622.950 652.050 625.050 ;
        RECT 644.400 611.400 648.450 612.450 ;
        RECT 617.400 606.450 618.600 606.600 ;
        RECT 614.400 605.400 618.600 606.450 ;
        RECT 608.400 604.200 609.600 604.950 ;
        RECT 617.400 604.200 618.600 605.400 ;
        RECT 619.950 604.950 622.050 607.050 ;
        RECT 628.950 605.100 631.050 607.200 ;
        RECT 637.950 605.100 640.050 607.200 ;
        RECT 643.950 605.100 646.050 607.200 ;
        RECT 647.400 607.050 648.450 611.400 ;
        RECT 595.950 601.950 598.050 604.050 ;
        RECT 586.950 589.950 589.050 592.050 ;
        RECT 592.950 589.950 595.050 592.050 ;
        RECT 587.400 580.050 588.450 589.950 ;
        RECT 596.400 586.050 597.450 601.950 ;
        RECT 601.950 601.800 604.050 603.900 ;
        RECT 604.950 601.800 607.050 603.900 ;
        RECT 607.950 601.800 610.050 603.900 ;
        RECT 616.950 601.800 619.050 603.900 ;
        RECT 619.950 601.800 622.050 603.900 ;
        RECT 622.950 601.800 625.050 603.900 ;
        RECT 605.400 600.000 606.600 601.500 ;
        RECT 604.950 595.950 607.050 600.000 ;
        RECT 613.950 598.950 616.050 601.050 ;
        RECT 620.400 599.400 621.600 601.500 ;
        RECT 601.950 592.950 604.050 595.050 ;
        RECT 595.950 583.950 598.050 586.050 ;
        RECT 591.000 582.450 595.050 583.050 ;
        RECT 590.400 580.950 595.050 582.450 ;
        RECT 586.950 577.950 589.050 580.050 ;
        RECT 590.400 573.600 591.450 580.950 ;
        RECT 595.950 577.950 598.050 580.050 ;
        RECT 590.400 571.500 591.600 573.600 ;
        RECT 596.400 573.450 597.450 577.950 ;
        RECT 602.400 577.050 603.450 592.950 ;
        RECT 614.400 589.050 615.450 598.950 ;
        RECT 613.950 586.950 616.050 589.050 ;
        RECT 620.400 588.450 621.450 599.400 ;
        RECT 629.400 595.050 630.450 605.100 ;
        RECT 638.400 604.350 639.600 605.100 ;
        RECT 644.400 604.350 645.600 605.100 ;
        RECT 646.950 604.950 649.050 607.050 ;
        RECT 634.950 601.950 637.050 604.050 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 640.950 601.950 643.050 604.050 ;
        RECT 643.950 601.950 646.050 604.050 ;
        RECT 635.400 599.400 636.600 601.650 ;
        RECT 641.400 600.000 642.600 601.650 ;
        RECT 628.950 592.950 631.050 595.050 ;
        RECT 620.400 587.400 624.450 588.450 ;
        RECT 604.950 583.950 607.050 586.050 ;
        RECT 619.950 583.950 622.050 586.050 ;
        RECT 601.950 574.950 604.050 577.050 ;
        RECT 605.400 574.200 606.450 583.950 ;
        RECT 610.950 580.950 613.050 583.050 ;
        RECT 596.400 572.400 600.450 573.450 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 571.950 568.950 574.050 571.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 580.950 568.950 583.050 571.050 ;
        RECT 586.950 569.100 589.050 571.200 ;
        RECT 589.950 569.100 592.050 571.200 ;
        RECT 592.950 569.100 595.050 571.200 ;
        RECT 551.400 568.050 552.600 568.800 ;
        RECT 523.950 562.950 526.050 565.050 ;
        RECT 520.950 559.950 523.050 562.050 ;
        RECT 502.950 556.950 505.050 559.050 ;
        RECT 511.950 556.950 514.050 559.050 ;
        RECT 508.950 544.950 511.050 547.050 ;
        RECT 490.800 535.950 492.900 538.050 ;
        RECT 485.400 527.400 489.450 528.450 ;
        RECT 478.950 505.950 481.050 508.050 ;
        RECT 478.950 500.400 481.050 502.500 ;
        RECT 466.950 493.950 469.050 496.050 ;
        RECT 467.400 469.050 468.450 493.950 ;
        RECT 472.950 490.950 475.050 493.050 ;
        RECT 473.400 488.400 474.600 490.650 ;
        RECT 473.400 484.050 474.450 488.400 ;
        RECT 472.950 481.950 475.050 484.050 ;
        RECT 479.100 480.600 480.300 500.400 ;
        RECT 485.400 495.450 486.450 527.400 ;
        RECT 496.950 526.950 499.050 529.050 ;
        RECT 509.400 528.600 510.450 544.950 ;
        RECT 497.400 526.200 498.600 526.950 ;
        RECT 509.400 526.350 510.600 528.600 ;
        RECT 514.950 527.100 517.050 529.200 ;
        RECT 515.400 526.350 516.600 527.100 ;
        RECT 490.950 523.800 493.050 525.900 ;
        RECT 493.950 523.800 496.050 525.900 ;
        RECT 496.950 523.800 499.050 525.900 ;
        RECT 505.950 523.950 508.050 526.050 ;
        RECT 508.950 523.950 511.050 526.050 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 514.950 523.950 517.050 526.050 ;
        RECT 487.950 520.950 490.050 523.050 ;
        RECT 494.400 521.400 495.600 523.500 ;
        RECT 502.950 522.450 505.050 523.050 ;
        RECT 506.400 522.450 507.600 523.650 ;
        RECT 502.950 521.400 507.600 522.450 ;
        RECT 512.400 521.400 513.600 523.650 ;
        RECT 488.400 505.050 489.450 520.950 ;
        RECT 494.400 517.050 495.450 521.400 ;
        RECT 502.950 520.950 505.050 521.400 ;
        RECT 493.950 514.950 496.050 517.050 ;
        RECT 487.950 502.950 490.050 505.050 ;
        RECT 503.400 502.050 504.450 520.950 ;
        RECT 505.950 502.950 508.050 505.050 ;
        RECT 502.950 499.950 505.050 502.050 ;
        RECT 485.400 494.400 489.450 495.450 ;
        RECT 481.950 490.950 484.050 493.050 ;
        RECT 482.400 489.450 483.600 490.650 ;
        RECT 482.400 488.400 486.450 489.450 ;
        RECT 478.950 478.500 481.050 480.600 ;
        RECT 466.950 466.950 469.050 469.050 ;
        RECT 469.950 458.400 472.050 460.500 ;
        RECT 466.950 450.450 469.050 451.200 ;
        RECT 464.400 449.400 469.050 450.450 ;
        RECT 466.950 449.100 469.050 449.400 ;
        RECT 458.400 448.350 459.600 449.100 ;
        RECT 467.400 448.350 468.600 449.100 ;
        RECT 451.950 445.950 454.050 448.050 ;
        RECT 454.950 445.950 457.050 448.050 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 466.950 445.950 469.050 448.050 ;
        RECT 455.400 444.900 456.600 445.650 ;
        RECT 445.950 442.800 448.050 444.900 ;
        RECT 454.950 442.800 457.050 444.900 ;
        RECT 461.400 443.400 462.600 445.650 ;
        RECT 427.950 436.950 430.050 439.050 ;
        RECT 461.400 430.050 462.450 443.400 ;
        RECT 463.950 436.950 466.050 439.050 ;
        RECT 470.700 438.600 471.900 458.400 ;
        RECT 475.950 454.950 478.050 457.050 ;
        RECT 476.400 450.600 477.450 454.950 ;
        RECT 485.400 451.200 486.450 488.400 ;
        RECT 488.400 478.050 489.450 494.400 ;
        RECT 496.950 494.250 499.050 496.350 ;
        RECT 497.400 493.500 498.600 494.250 ;
        RECT 493.950 491.100 496.050 493.200 ;
        RECT 496.950 491.100 499.050 493.200 ;
        RECT 499.950 491.100 502.050 493.200 ;
        RECT 500.400 489.450 501.600 490.800 ;
        RECT 500.400 488.400 504.450 489.450 ;
        RECT 487.950 475.950 490.050 478.050 ;
        RECT 503.400 475.050 504.450 488.400 ;
        RECT 502.950 472.950 505.050 475.050 ;
        RECT 490.950 459.300 493.050 461.400 ;
        RECT 502.950 460.950 505.050 463.050 ;
        RECT 490.950 455.700 492.150 459.300 ;
        RECT 490.950 453.600 493.050 455.700 ;
        RECT 476.400 448.350 477.600 450.600 ;
        RECT 484.950 449.100 487.050 451.200 ;
        RECT 475.950 445.950 478.050 448.050 ;
        RECT 475.950 439.950 478.050 442.050 ;
        RECT 460.950 427.950 463.050 430.050 ;
        RECT 464.400 427.050 465.450 436.950 ;
        RECT 469.950 436.500 472.050 438.600 ;
        RECT 466.950 430.950 469.050 433.050 ;
        RECT 463.950 424.950 466.050 427.050 ;
        RECT 415.950 421.950 418.050 424.050 ;
        RECT 424.950 422.400 427.050 424.500 ;
        RECT 445.950 422.400 448.050 424.500 ;
        RECT 412.950 418.950 415.050 421.050 ;
        RECT 400.800 415.950 402.900 418.050 ;
        RECT 403.950 416.100 406.050 418.200 ;
        RECT 409.950 416.100 412.050 418.200 ;
        RECT 404.400 415.350 405.600 416.100 ;
        RECT 410.400 415.350 411.600 416.100 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 412.950 412.950 415.050 415.050 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 407.400 410.400 408.600 412.650 ;
        RECT 413.400 411.900 414.600 412.650 ;
        RECT 397.950 406.950 400.050 409.050 ;
        RECT 397.950 403.800 400.050 405.900 ;
        RECT 398.400 394.050 399.450 403.800 ;
        RECT 397.950 391.950 400.050 394.050 ;
        RECT 407.400 391.050 408.450 410.400 ;
        RECT 412.950 409.800 415.050 411.900 ;
        RECT 422.400 410.400 423.600 412.650 ;
        RECT 422.400 406.050 423.450 410.400 ;
        RECT 421.950 403.950 424.050 406.050 ;
        RECT 425.700 402.600 426.900 422.400 ;
        RECT 439.950 415.950 442.050 418.050 ;
        RECT 430.950 412.950 433.050 415.050 ;
        RECT 431.400 411.900 432.600 412.650 ;
        RECT 440.400 411.900 441.450 415.950 ;
        RECT 430.950 409.800 433.050 411.900 ;
        RECT 439.950 409.800 442.050 411.900 ;
        RECT 445.950 407.400 447.150 422.400 ;
        RECT 448.950 416.100 451.050 418.200 ;
        RECT 449.400 415.350 450.600 416.100 ;
        RECT 457.950 415.950 460.050 418.050 ;
        RECT 467.400 417.600 468.450 430.950 ;
        RECT 448.950 412.950 451.050 415.050 ;
        RECT 454.950 412.950 457.050 415.050 ;
        RECT 455.400 409.050 456.450 412.950 ;
        RECT 458.400 412.050 459.450 415.950 ;
        RECT 467.400 415.500 468.600 417.600 ;
        RECT 463.950 413.100 466.050 415.200 ;
        RECT 466.950 413.100 469.050 415.200 ;
        RECT 469.950 413.100 472.050 415.200 ;
        RECT 464.400 412.050 465.600 412.800 ;
        RECT 457.950 409.950 460.050 412.050 ;
        RECT 463.950 409.950 466.050 412.050 ;
        RECT 470.400 411.000 471.600 412.800 ;
        RECT 445.950 405.300 448.050 407.400 ;
        RECT 454.950 406.950 457.050 409.050 ;
        RECT 469.950 406.950 472.050 411.000 ;
        RECT 424.950 400.500 427.050 402.600 ;
        RECT 445.950 401.700 447.150 405.300 ;
        RECT 445.950 399.600 448.050 401.700 ;
        RECT 406.950 388.950 409.050 391.050 ;
        RECT 400.950 372.000 403.050 376.050 ;
        RECT 448.950 373.050 451.050 373.200 ;
        RECT 455.400 373.050 456.450 406.950 ;
        RECT 401.400 370.350 402.600 372.000 ;
        RECT 412.950 370.950 415.050 373.050 ;
        RECT 418.950 370.950 421.050 373.050 ;
        RECT 427.950 370.950 430.050 373.050 ;
        RECT 436.950 372.600 441.000 373.050 ;
        RECT 436.950 370.950 441.600 372.600 ;
        RECT 448.950 371.100 454.050 373.050 ;
        RECT 400.950 367.950 403.050 370.050 ;
        RECT 406.950 367.950 409.050 370.050 ;
        RECT 407.400 365.400 408.600 367.650 ;
        RECT 394.950 352.950 397.050 355.050 ;
        RECT 407.400 352.050 408.450 365.400 ;
        RECT 413.400 364.050 414.450 370.950 ;
        RECT 419.400 370.200 420.600 370.950 ;
        RECT 428.400 370.200 429.600 370.950 ;
        RECT 440.400 370.350 441.600 370.950 ;
        RECT 449.400 370.950 454.050 371.100 ;
        RECT 454.950 370.950 457.050 373.050 ;
        RECT 457.950 370.950 460.050 373.050 ;
        RECT 463.950 370.950 466.050 373.050 ;
        RECT 469.800 370.950 471.900 373.050 ;
        RECT 472.950 371.100 475.050 373.200 ;
        RECT 476.400 373.050 477.450 439.950 ;
        RECT 485.400 432.450 486.450 449.100 ;
        RECT 490.950 438.600 492.150 453.600 ;
        RECT 499.950 448.950 502.050 451.050 ;
        RECT 493.950 445.950 496.050 448.050 ;
        RECT 494.400 444.900 495.600 445.650 ;
        RECT 493.950 442.800 496.050 444.900 ;
        RECT 490.950 436.500 493.050 438.600 ;
        RECT 500.400 433.050 501.450 448.950 ;
        RECT 503.400 444.900 504.450 460.950 ;
        RECT 506.400 454.050 507.450 502.950 ;
        RECT 512.400 495.450 513.450 521.400 ;
        RECT 517.950 520.950 520.050 523.050 ;
        RECT 518.400 517.050 519.450 520.950 ;
        RECT 517.950 514.950 520.050 517.050 ;
        RECT 517.950 508.950 520.050 511.050 ;
        RECT 509.400 494.400 513.450 495.450 ;
        RECT 518.400 495.600 519.450 508.950 ;
        RECT 521.400 499.050 522.450 559.950 ;
        RECT 524.400 547.050 525.450 562.950 ;
        RECT 527.400 562.050 528.450 565.950 ;
        RECT 533.400 562.050 534.450 566.400 ;
        RECT 538.950 565.800 541.050 567.900 ;
        RECT 544.950 565.800 547.050 567.900 ;
        RECT 550.950 565.950 553.050 568.050 ;
        RECT 559.950 565.950 562.050 568.050 ;
        RECT 572.400 567.900 573.600 568.650 ;
        RECT 587.400 568.050 588.600 568.800 ;
        RECT 526.950 559.950 529.050 562.050 ;
        RECT 532.950 559.950 535.050 562.050 ;
        RECT 551.400 550.050 552.450 565.950 ;
        RECT 560.400 559.050 561.450 565.950 ;
        RECT 571.950 565.800 574.050 567.900 ;
        RECT 580.950 565.800 583.050 567.900 ;
        RECT 586.950 565.950 589.050 568.050 ;
        RECT 589.950 565.950 592.050 568.050 ;
        RECT 595.800 565.950 597.900 568.050 ;
        RECT 599.400 567.900 600.450 572.400 ;
        RECT 604.950 572.100 607.050 574.200 ;
        RECT 611.400 573.600 612.450 580.950 ;
        RECT 605.400 571.350 606.600 572.100 ;
        RECT 611.400 571.350 612.600 573.600 ;
        RECT 604.950 568.950 607.050 571.050 ;
        RECT 607.950 568.950 610.050 571.050 ;
        RECT 610.950 568.950 613.050 571.050 ;
        RECT 613.950 568.950 616.050 571.050 ;
        RECT 608.400 567.900 609.600 568.650 ;
        RECT 614.400 567.900 615.600 568.650 ;
        RECT 559.950 556.950 562.050 559.050 ;
        RECT 550.950 547.950 553.050 550.050 ;
        RECT 577.950 547.950 580.050 550.050 ;
        RECT 523.950 544.950 526.050 547.050 ;
        RECT 529.950 541.950 532.050 544.050 ;
        RECT 547.950 541.950 550.050 544.050 ;
        RECT 530.400 529.050 531.450 541.950 ;
        RECT 532.950 532.950 535.050 535.050 ;
        RECT 533.400 529.050 534.450 532.950 ;
        RECT 529.950 526.950 532.050 529.050 ;
        RECT 532.950 526.950 535.050 529.050 ;
        RECT 538.950 526.950 541.050 529.200 ;
        RECT 548.400 528.600 549.450 541.950 ;
        RECT 559.950 538.950 562.050 541.050 ;
        RECT 533.400 526.200 534.600 526.950 ;
        RECT 526.950 523.800 529.050 525.900 ;
        RECT 529.950 523.800 532.050 525.900 ;
        RECT 532.950 523.800 535.050 525.900 ;
        RECT 530.400 522.750 531.600 523.500 ;
        RECT 539.400 523.050 540.450 526.950 ;
        RECT 548.400 526.350 549.600 528.600 ;
        RECT 553.950 527.100 556.050 529.200 ;
        RECT 560.400 528.450 561.450 538.950 ;
        RECT 565.950 536.400 568.050 538.500 ;
        RECT 563.400 528.450 564.600 528.600 ;
        RECT 560.400 527.400 564.600 528.450 ;
        RECT 554.400 526.350 555.600 527.100 ;
        RECT 563.400 526.350 564.600 527.400 ;
        RECT 541.950 523.950 544.050 526.050 ;
        RECT 547.950 523.950 550.050 526.050 ;
        RECT 550.950 523.950 553.050 526.050 ;
        RECT 553.950 523.950 556.050 526.050 ;
        RECT 556.950 523.950 559.050 526.050 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 529.950 520.650 532.050 522.750 ;
        RECT 538.950 520.950 541.050 523.050 ;
        RECT 538.950 517.800 541.050 519.900 ;
        RECT 523.950 505.950 526.050 508.050 ;
        RECT 520.950 496.950 523.050 499.050 ;
        RECT 524.400 495.600 525.450 505.950 ;
        RECT 532.950 499.950 535.050 502.050 ;
        RECT 533.400 495.600 534.450 499.950 ;
        RECT 539.400 495.600 540.450 517.800 ;
        RECT 542.400 511.050 543.450 523.950 ;
        RECT 544.950 520.950 547.050 523.050 ;
        RECT 551.400 521.400 552.600 523.650 ;
        RECT 557.400 522.450 558.600 523.650 ;
        RECT 557.400 522.000 561.450 522.450 ;
        RECT 557.400 521.400 562.050 522.000 ;
        RECT 541.950 508.950 544.050 511.050 ;
        RECT 545.400 496.050 546.450 520.950 ;
        RECT 551.400 511.050 552.450 521.400 ;
        RECT 553.950 511.950 556.050 514.050 ;
        RECT 550.950 508.950 553.050 511.050 ;
        RECT 547.950 496.950 550.050 499.050 ;
        RECT 509.400 484.050 510.450 494.400 ;
        RECT 518.400 493.350 519.600 495.600 ;
        RECT 524.400 493.350 525.600 495.600 ;
        RECT 533.400 493.350 534.600 495.600 ;
        RECT 539.400 493.350 540.600 495.600 ;
        RECT 544.950 493.950 547.050 496.050 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 520.950 490.950 523.050 493.050 ;
        RECT 523.950 490.950 526.050 493.050 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 535.950 490.950 538.050 493.050 ;
        RECT 538.950 490.950 541.050 493.050 ;
        RECT 541.950 490.950 544.050 493.050 ;
        RECT 515.400 489.900 516.600 490.650 ;
        RECT 514.950 487.800 517.050 489.900 ;
        RECT 521.400 488.400 522.600 490.650 ;
        RECT 517.950 484.950 520.050 487.050 ;
        RECT 508.950 481.950 511.050 484.050 ;
        RECT 518.400 481.050 519.450 484.950 ;
        RECT 517.950 478.950 520.050 481.050 ;
        RECT 514.950 475.950 517.050 478.050 ;
        RECT 505.950 451.950 508.050 454.050 ;
        RECT 515.400 451.200 516.450 475.950 ;
        RECT 521.400 475.050 522.450 488.400 ;
        RECT 529.950 487.950 532.050 490.050 ;
        RECT 536.400 489.900 537.600 490.650 ;
        RECT 530.400 475.050 531.450 487.950 ;
        RECT 535.950 487.800 538.050 489.900 ;
        RECT 542.400 489.000 543.600 490.650 ;
        RECT 548.400 489.900 549.450 496.950 ;
        RECT 550.950 494.100 553.050 496.200 ;
        RECT 554.400 496.050 555.450 511.950 ;
        RECT 557.400 502.050 558.450 521.400 ;
        RECT 559.950 517.950 562.050 521.400 ;
        RECT 566.700 516.600 567.900 536.400 ;
        RECT 571.950 527.100 574.050 529.200 ;
        RECT 572.400 526.350 573.600 527.100 ;
        RECT 571.950 523.950 574.050 526.050 ;
        RECT 574.950 520.950 577.050 523.050 ;
        RECT 565.950 514.500 568.050 516.600 ;
        RECT 562.950 508.950 565.050 511.050 ;
        RECT 575.400 510.450 576.450 520.950 ;
        RECT 578.400 514.050 579.450 547.950 ;
        RECT 581.400 544.050 582.450 565.800 ;
        RECT 590.400 556.050 591.450 565.950 ;
        RECT 589.950 553.950 592.050 556.050 ;
        RECT 580.950 541.950 583.050 544.050 ;
        RECT 580.950 535.950 583.050 538.050 ;
        RECT 586.950 537.300 589.050 539.400 ;
        RECT 577.950 511.950 580.050 514.050 ;
        RECT 575.400 509.400 579.450 510.450 ;
        RECT 556.950 499.950 559.050 502.050 ;
        RECT 541.950 484.950 544.050 489.000 ;
        RECT 547.950 487.800 550.050 489.900 ;
        RECT 551.400 487.050 552.450 494.100 ;
        RECT 553.950 493.950 556.050 496.050 ;
        RECT 559.800 494.100 561.900 496.200 ;
        RECT 563.400 496.050 564.450 508.950 ;
        RECT 568.950 505.950 571.050 508.050 ;
        RECT 574.950 505.950 577.050 508.050 ;
        RECT 560.400 493.350 561.600 494.100 ;
        RECT 562.950 493.950 565.050 496.050 ;
        RECT 569.400 495.600 570.450 505.950 ;
        RECT 575.400 502.050 576.450 505.950 ;
        RECT 574.950 499.950 577.050 502.050 ;
        RECT 578.400 496.200 579.450 509.400 ;
        RECT 581.400 508.050 582.450 535.950 ;
        RECT 586.950 533.700 588.150 537.300 ;
        RECT 586.950 531.600 589.050 533.700 ;
        RECT 586.950 516.600 588.150 531.600 ;
        RECT 589.950 523.950 592.050 526.050 ;
        RECT 590.400 522.900 591.600 523.650 ;
        RECT 589.950 520.800 592.050 522.900 ;
        RECT 596.400 520.050 597.450 565.950 ;
        RECT 598.950 565.800 601.050 567.900 ;
        RECT 607.950 565.800 610.050 567.900 ;
        RECT 613.950 565.800 616.050 567.900 ;
        RECT 598.950 559.950 601.050 562.050 ;
        RECT 595.950 517.950 598.050 520.050 ;
        RECT 586.950 514.500 589.050 516.600 ;
        RECT 583.950 508.950 586.050 511.050 ;
        RECT 580.950 505.950 583.050 508.050 ;
        RECT 580.950 502.800 583.050 504.900 ;
        RECT 569.400 493.350 570.600 495.600 ;
        RECT 574.800 494.100 576.900 496.200 ;
        RECT 577.950 494.100 580.050 496.200 ;
        RECT 575.400 493.350 576.600 494.100 ;
        RECT 556.950 490.950 559.050 493.050 ;
        RECT 559.950 490.950 562.050 493.050 ;
        RECT 568.950 490.950 571.050 493.050 ;
        RECT 571.950 490.950 574.050 493.050 ;
        RECT 574.950 490.950 577.050 493.050 ;
        RECT 553.950 487.950 556.050 490.050 ;
        RECT 557.400 488.400 558.600 490.650 ;
        RECT 572.400 489.000 573.600 490.650 ;
        RECT 550.950 484.950 553.050 487.050 ;
        RECT 520.950 472.950 523.050 475.050 ;
        RECT 529.950 472.950 532.050 475.050 ;
        RECT 544.950 472.950 547.050 475.050 ;
        RECT 532.950 460.950 535.050 463.050 ;
        RECT 507.000 450.900 510.000 451.050 ;
        RECT 505.950 450.600 510.000 450.900 ;
        RECT 505.950 448.950 510.600 450.600 ;
        RECT 514.950 449.100 517.050 451.200 ;
        RECT 505.950 448.800 508.050 448.950 ;
        RECT 509.400 448.350 510.600 448.950 ;
        RECT 515.400 448.350 516.600 449.100 ;
        RECT 523.950 448.950 526.050 451.050 ;
        RECT 533.400 450.600 534.450 460.950 ;
        RECT 545.400 450.600 546.450 472.950 ;
        RECT 554.400 463.050 555.450 487.950 ;
        RECT 553.950 460.950 556.050 463.050 ;
        RECT 550.950 457.950 553.050 460.050 ;
        RECT 551.400 450.600 552.450 457.950 ;
        RECT 557.400 451.200 558.450 488.400 ;
        RECT 571.950 484.950 574.050 489.000 ;
        RECT 577.950 475.950 580.050 481.050 ;
        RECT 581.400 478.050 582.450 502.800 ;
        RECT 584.400 502.050 585.450 508.950 ;
        RECT 583.950 499.950 586.050 502.050 ;
        RECT 596.400 499.050 597.450 517.950 ;
        RECT 599.400 505.050 600.450 559.950 ;
        RECT 604.950 550.950 607.050 553.050 ;
        RECT 605.400 544.050 606.450 550.950 ;
        RECT 608.400 550.050 609.450 565.800 ;
        RECT 620.400 562.050 621.450 583.950 ;
        RECT 623.400 574.050 624.450 587.400 ;
        RECT 622.950 571.950 625.050 574.050 ;
        RECT 629.400 573.600 630.450 592.950 ;
        RECT 635.400 586.050 636.450 599.400 ;
        RECT 640.950 595.950 643.050 600.000 ;
        RECT 646.950 598.950 649.050 601.050 ;
        RECT 634.950 583.950 637.050 586.050 ;
        RECT 635.400 573.600 636.450 583.950 ;
        RECT 647.400 577.200 648.450 598.950 ;
        RECT 646.950 575.100 649.050 577.200 ;
        RECT 650.400 574.050 651.450 622.950 ;
        RECT 652.950 605.100 655.050 607.200 ;
        RECT 656.400 607.050 657.450 640.950 ;
        RECT 662.400 637.050 663.450 646.950 ;
        RECT 668.400 645.000 669.600 646.800 ;
        RECT 674.400 646.050 675.600 646.800 ;
        RECT 683.400 646.050 684.600 646.800 ;
        RECT 667.950 640.950 670.050 645.000 ;
        RECT 673.950 643.950 676.050 646.050 ;
        RECT 682.950 643.950 688.050 646.050 ;
        RECT 689.400 644.400 690.600 646.800 ;
        RECT 661.950 634.950 664.050 637.050 ;
        RECT 668.400 634.050 669.450 640.950 ;
        RECT 667.950 631.950 670.050 634.050 ;
        RECT 664.950 616.950 667.050 619.050 ;
        RECT 653.400 583.050 654.450 605.100 ;
        RECT 655.950 604.950 658.050 607.050 ;
        RECT 658.950 605.100 661.050 607.200 ;
        RECT 665.400 606.600 666.450 616.950 ;
        RECT 674.400 613.050 675.450 643.950 ;
        RECT 689.400 634.050 690.450 644.400 ;
        RECT 688.950 631.950 691.050 634.050 ;
        RECT 698.400 619.050 699.450 650.400 ;
        RECT 706.950 650.250 709.050 652.350 ;
        RECT 713.400 651.600 714.450 667.950 ;
        RECT 707.400 649.500 708.600 650.250 ;
        RECT 713.400 649.500 714.600 651.600 ;
        RECT 703.950 647.100 706.050 649.200 ;
        RECT 706.950 647.100 709.050 649.200 ;
        RECT 709.950 647.100 712.050 649.200 ;
        RECT 712.950 647.100 715.050 649.200 ;
        RECT 704.400 644.400 705.600 646.800 ;
        RECT 710.400 644.400 711.600 646.800 ;
        RECT 704.400 634.050 705.450 644.400 ;
        RECT 710.400 637.050 711.450 644.400 ;
        RECT 709.950 634.950 712.050 637.050 ;
        RECT 703.950 631.950 706.050 634.050 ;
        RECT 679.950 616.950 682.050 619.050 ;
        RECT 691.950 616.950 694.050 619.050 ;
        RECT 697.950 616.950 700.050 619.050 ;
        RECT 712.950 616.950 715.050 619.050 ;
        RECT 673.950 610.950 676.050 613.050 ;
        RECT 674.400 607.050 675.450 610.950 ;
        RECT 659.400 604.350 660.600 605.100 ;
        RECT 665.400 604.350 666.600 606.600 ;
        RECT 673.950 604.950 676.050 607.050 ;
        RECT 680.400 606.600 681.450 616.950 ;
        RECT 685.950 610.950 688.050 613.050 ;
        RECT 686.400 606.600 687.450 610.950 ;
        RECT 680.400 604.350 681.600 606.600 ;
        RECT 686.400 604.350 687.600 606.600 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 661.950 601.950 664.050 604.050 ;
        RECT 664.950 601.950 667.050 604.050 ;
        RECT 667.950 601.950 670.050 604.050 ;
        RECT 676.950 601.950 679.050 604.050 ;
        RECT 679.950 601.950 682.050 604.050 ;
        RECT 682.950 601.950 685.050 604.050 ;
        RECT 685.950 601.950 688.050 604.050 ;
        RECT 655.950 595.950 658.050 601.050 ;
        RECT 662.400 600.900 663.600 601.650 ;
        RECT 661.950 598.800 664.050 600.900 ;
        RECT 668.400 599.400 669.600 601.650 ;
        RECT 668.400 595.050 669.450 599.400 ;
        RECT 673.950 598.950 676.050 601.050 ;
        RECT 677.400 599.400 678.600 601.650 ;
        RECT 683.400 599.400 684.600 601.650 ;
        RECT 667.950 592.950 670.050 595.050 ;
        RECT 658.950 586.950 661.050 589.050 ;
        RECT 652.950 580.950 655.050 583.050 ;
        RECT 659.400 577.050 660.450 586.950 ;
        RECT 664.950 580.950 667.050 583.050 ;
        RECT 658.950 574.950 661.050 577.050 ;
        RECT 665.400 576.450 666.450 580.950 ;
        RECT 665.400 575.400 669.450 576.450 ;
        RECT 629.400 571.350 630.600 573.600 ;
        RECT 635.400 571.350 636.600 573.600 ;
        RECT 646.800 571.950 648.900 574.050 ;
        RECT 649.950 571.950 652.050 574.050 ;
        RECT 647.400 571.350 648.600 571.950 ;
        RECT 658.950 571.800 661.050 573.900 ;
        RECT 668.400 573.600 669.450 575.400 ;
        RECT 674.400 573.600 675.450 598.950 ;
        RECT 677.400 595.050 678.450 599.400 ;
        RECT 676.950 592.950 679.050 595.050 ;
        RECT 677.400 574.050 678.450 592.950 ;
        RECT 683.400 577.050 684.450 599.400 ;
        RECT 692.400 598.050 693.450 616.950 ;
        RECT 697.950 606.000 700.050 610.050 ;
        RECT 698.400 604.200 699.600 606.000 ;
        RECT 703.950 604.950 706.050 607.050 ;
        RECT 704.400 604.200 705.600 604.950 ;
        RECT 697.950 601.800 700.050 603.900 ;
        RECT 700.950 601.800 703.050 603.900 ;
        RECT 703.950 601.800 706.050 603.900 ;
        RECT 706.950 601.800 709.050 603.900 ;
        RECT 701.400 600.750 702.600 601.500 ;
        RECT 700.950 598.650 703.050 600.750 ;
        RECT 707.400 599.400 708.600 601.500 ;
        RECT 713.400 600.750 714.450 616.950 ;
        RECT 719.400 610.050 720.450 673.950 ;
        RECT 722.400 673.050 723.450 677.400 ;
        RECT 721.950 670.950 724.050 673.050 ;
        RECT 728.400 658.050 729.450 677.400 ;
        RECT 737.400 667.050 738.450 685.950 ;
        RECT 743.400 684.600 744.450 688.950 ;
        RECT 743.400 682.350 744.600 684.600 ;
        RECT 748.950 683.100 751.050 685.200 ;
        RECT 763.950 683.100 766.050 685.200 ;
        RECT 770.400 684.600 771.450 694.950 ;
        RECT 749.400 682.350 750.600 683.100 ;
        RECT 764.400 682.350 765.600 683.100 ;
        RECT 770.400 682.350 771.600 684.600 ;
        RECT 784.950 683.100 787.050 685.200 ;
        RECT 785.400 682.350 786.600 683.100 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 748.950 679.950 751.050 682.050 ;
        RECT 751.950 679.950 754.050 682.050 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 769.950 679.950 772.050 682.050 ;
        RECT 781.950 679.950 784.050 682.050 ;
        RECT 784.950 679.950 787.050 682.050 ;
        RECT 746.400 677.400 747.600 679.650 ;
        RECT 752.400 677.400 753.600 679.650 ;
        RECT 761.400 677.400 762.600 679.650 ;
        RECT 767.400 678.000 768.600 679.650 ;
        RECT 736.950 664.950 739.050 667.050 ;
        RECT 746.400 658.050 747.450 677.400 ;
        RECT 752.400 670.050 753.450 677.400 ;
        RECT 757.950 673.950 760.050 676.050 ;
        RECT 751.950 667.950 754.050 670.050 ;
        RECT 727.950 655.950 730.050 658.050 ;
        RECT 742.800 655.950 744.900 658.050 ;
        RECT 745.950 655.950 748.050 658.050 ;
        RECT 751.950 655.950 754.050 658.050 ;
        RECT 730.950 650.100 733.050 652.200 ;
        RECT 743.400 651.600 744.450 655.950 ;
        RECT 731.400 649.350 732.600 650.100 ;
        RECT 743.400 649.500 744.600 651.600 ;
        RECT 748.950 650.250 751.050 652.350 ;
        RECT 752.400 652.050 753.450 655.950 ;
        RECT 758.400 652.050 759.450 673.950 ;
        RECT 761.400 670.050 762.450 677.400 ;
        RECT 766.950 673.950 769.050 678.000 ;
        RECT 782.400 677.400 783.600 679.650 ;
        RECT 794.400 678.900 795.450 697.950 ;
        RECT 800.400 684.600 801.450 703.800 ;
        RECT 803.400 687.450 804.450 727.950 ;
        RECT 812.400 727.350 813.600 728.100 ;
        RECT 818.400 727.350 819.600 729.600 ;
        RECT 820.950 727.950 823.050 730.050 ;
        RECT 808.950 724.950 811.050 727.050 ;
        RECT 811.950 724.950 814.050 727.050 ;
        RECT 814.950 724.950 817.050 727.050 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 809.400 722.400 810.600 724.650 ;
        RECT 815.400 723.000 816.600 724.650 ;
        RECT 809.400 706.050 810.450 722.400 ;
        RECT 814.950 718.950 817.050 723.000 ;
        RECT 820.950 721.950 823.050 724.050 ;
        RECT 808.950 703.950 811.050 706.050 ;
        RECT 811.950 697.950 814.050 700.050 ;
        RECT 803.400 687.000 807.450 687.450 ;
        RECT 803.400 686.400 808.050 687.000 ;
        RECT 800.400 682.350 801.600 684.600 ;
        RECT 805.950 682.950 808.050 686.400 ;
        RECT 812.400 684.600 813.450 697.950 ;
        RECT 812.400 682.200 813.600 684.600 ;
        RECT 818.400 684.450 819.600 684.600 ;
        RECT 821.400 684.450 822.450 721.950 ;
        RECT 824.400 721.050 825.450 730.950 ;
        RECT 827.400 730.050 828.450 743.400 ;
        RECT 829.950 739.950 832.050 742.050 ;
        RECT 826.950 727.950 829.050 730.050 ;
        RECT 830.400 729.600 831.450 739.950 ;
        RECT 839.400 739.050 840.450 755.400 ;
        RECT 841.950 754.950 844.050 757.050 ;
        RECT 847.950 754.950 850.050 757.050 ;
        RECT 851.400 755.400 852.600 757.650 ;
        RECT 838.950 736.950 841.050 739.050 ;
        RECT 830.400 727.500 831.600 729.600 ;
        RECT 835.950 729.000 838.050 733.050 ;
        RECT 842.400 730.050 843.450 754.950 ;
        RECT 836.400 727.500 837.600 729.000 ;
        RECT 841.950 727.950 844.050 730.050 ;
        RECT 848.400 729.600 849.450 754.950 ;
        RECT 851.400 733.050 852.450 755.400 ;
        RECT 850.950 730.950 853.050 733.050 ;
        RECT 848.400 727.350 849.600 729.600 ;
        RECT 853.950 728.100 856.050 730.200 ;
        RECT 854.400 727.350 855.600 728.100 ;
        RECT 829.950 725.100 832.050 727.200 ;
        RECT 832.950 725.100 835.050 727.200 ;
        RECT 835.950 725.100 838.050 727.200 ;
        RECT 838.950 725.100 841.050 727.200 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 853.950 724.950 856.050 727.050 ;
        RECT 856.950 724.950 859.050 727.050 ;
        RECT 833.400 722.400 834.600 724.800 ;
        RECT 839.400 724.050 840.600 724.800 ;
        RECT 833.400 721.050 834.450 722.400 ;
        RECT 835.800 721.950 837.900 724.050 ;
        RECT 838.950 721.950 841.050 724.050 ;
        RECT 823.950 718.950 826.050 721.050 ;
        RECT 832.950 718.950 835.050 721.050 ;
        RECT 826.950 706.950 829.050 709.050 ;
        RECT 818.400 683.400 822.450 684.450 ;
        RECT 818.400 682.200 819.600 683.400 ;
        RECT 799.950 679.950 802.050 682.050 ;
        RECT 802.950 679.950 805.050 682.050 ;
        RECT 811.950 679.800 814.050 681.900 ;
        RECT 814.950 679.800 817.050 681.900 ;
        RECT 817.950 679.800 820.050 681.900 ;
        RECT 820.950 679.800 823.050 681.900 ;
        RECT 803.400 678.900 804.600 679.650 ;
        RECT 760.950 667.950 763.050 670.050 ;
        RECT 766.950 667.950 769.050 670.050 ;
        RECT 763.950 658.950 766.050 661.050 ;
        RECT 749.400 649.500 750.600 650.250 ;
        RECT 751.950 649.950 754.050 652.050 ;
        RECT 754.800 649.950 756.900 652.050 ;
        RECT 757.950 649.950 760.050 652.050 ;
        RECT 764.400 651.600 765.450 658.950 ;
        RECT 767.400 655.050 768.450 667.950 ;
        RECT 782.400 667.050 783.450 677.400 ;
        RECT 793.950 676.800 796.050 678.900 ;
        RECT 802.950 676.800 805.050 678.900 ;
        RECT 808.950 676.950 811.050 679.050 ;
        RECT 815.400 677.400 816.600 679.500 ;
        RECT 821.400 677.400 822.600 679.500 ;
        RECT 784.950 667.950 787.050 670.050 ;
        RECT 781.950 664.950 784.050 667.050 ;
        RECT 772.950 658.950 775.050 661.050 ;
        RECT 766.950 652.950 769.050 655.050 ;
        RECT 721.950 646.950 724.050 649.050 ;
        RECT 727.950 646.950 730.050 649.050 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 739.950 647.100 742.050 649.200 ;
        RECT 742.950 647.100 745.050 649.200 ;
        RECT 745.950 647.100 748.050 649.200 ;
        RECT 748.950 647.100 751.050 649.200 ;
        RECT 722.400 640.050 723.450 646.950 ;
        RECT 728.400 644.400 729.600 646.650 ;
        RECT 740.400 644.400 741.600 646.800 ;
        RECT 746.400 646.050 747.600 646.800 ;
        RECT 721.950 637.950 724.050 640.050 ;
        RECT 728.400 634.050 729.450 644.400 ;
        RECT 740.400 640.050 741.450 644.400 ;
        RECT 745.950 643.950 748.050 646.050 ;
        RECT 751.950 640.950 754.050 646.050 ;
        RECT 739.950 637.950 742.050 640.050 ;
        RECT 755.400 637.050 756.450 649.950 ;
        RECT 764.400 649.500 765.600 651.600 ;
        RECT 769.950 650.250 772.050 652.350 ;
        RECT 773.400 652.050 774.450 658.950 ;
        RECT 770.400 649.500 771.600 650.250 ;
        RECT 772.950 649.950 775.050 652.050 ;
        RECT 775.950 649.950 778.050 652.050 ;
        RECT 785.400 651.600 786.450 667.950 ;
        RECT 796.950 661.950 799.050 664.050 ;
        RECT 760.950 647.100 763.050 649.200 ;
        RECT 763.950 647.100 766.050 649.200 ;
        RECT 766.950 647.100 769.050 649.200 ;
        RECT 769.950 647.100 772.050 649.200 ;
        RECT 757.950 640.950 760.050 646.050 ;
        RECT 761.400 644.400 762.600 646.800 ;
        RECT 754.950 634.950 757.050 637.050 ;
        RECT 761.400 634.050 762.450 644.400 ;
        RECT 763.950 643.950 766.050 646.050 ;
        RECT 767.400 645.000 768.600 646.800 ;
        RECT 776.400 646.050 777.450 649.950 ;
        RECT 785.400 649.500 786.600 651.600 ;
        RECT 793.950 649.950 796.050 652.050 ;
        RECT 781.950 647.100 784.050 649.200 ;
        RECT 784.950 647.100 787.050 649.200 ;
        RECT 787.950 647.100 790.050 649.200 ;
        RECT 782.400 646.050 783.600 646.800 ;
        RECT 788.400 646.050 789.600 646.800 ;
        RECT 727.950 631.950 730.050 634.050 ;
        RECT 760.950 631.950 763.050 634.050 ;
        RECT 751.950 619.950 754.050 622.050 ;
        RECT 752.400 616.050 753.450 619.950 ;
        RECT 764.400 616.050 765.450 643.950 ;
        RECT 766.950 640.950 769.050 645.000 ;
        RECT 775.950 643.950 778.050 646.050 ;
        RECT 781.950 643.950 784.050 646.050 ;
        RECT 787.950 643.950 790.050 646.050 ;
        RECT 788.400 640.050 789.450 643.950 ;
        RECT 794.400 640.050 795.450 649.950 ;
        RECT 787.950 637.950 790.050 640.050 ;
        RECT 793.950 637.950 796.050 640.050 ;
        RECT 797.400 637.050 798.450 661.950 ;
        RECT 809.400 655.050 810.450 676.950 ;
        RECT 815.400 673.050 816.450 677.400 ;
        RECT 821.400 675.450 822.450 677.400 ;
        RECT 818.400 674.400 822.450 675.450 ;
        RECT 814.950 670.950 817.050 673.050 ;
        RECT 818.400 655.050 819.450 674.400 ;
        RECT 820.950 670.950 823.050 673.050 ;
        RECT 805.800 654.000 807.900 655.050 ;
        RECT 805.800 652.950 808.050 654.000 ;
        RECT 808.950 652.950 811.050 655.050 ;
        RECT 817.950 652.950 820.050 655.050 ;
        RECT 805.950 651.000 808.050 652.950 ;
        RECT 821.400 651.600 822.450 670.950 ;
        RECT 827.400 661.050 828.450 706.950 ;
        RECT 833.400 703.050 834.450 718.950 ;
        RECT 832.950 700.950 835.050 703.050 ;
        RECT 833.400 684.600 834.450 700.950 ;
        RECT 836.400 685.050 837.450 721.950 ;
        RECT 833.400 682.200 834.600 684.600 ;
        RECT 835.950 682.950 838.050 685.050 ;
        RECT 839.400 684.600 840.450 721.950 ;
        RECT 844.950 718.950 847.050 724.050 ;
        RECT 851.400 722.400 852.600 724.650 ;
        RECT 857.400 723.000 858.600 724.650 ;
        RECT 851.400 712.050 852.450 722.400 ;
        RECT 856.950 718.950 859.050 723.000 ;
        RECT 859.950 721.950 862.050 724.050 ;
        RECT 850.950 709.950 853.050 712.050 ;
        RECT 839.400 682.200 840.600 684.600 ;
        RECT 853.950 682.950 856.050 685.050 ;
        RECT 832.950 679.800 835.050 681.900 ;
        RECT 835.950 679.800 838.050 681.900 ;
        RECT 838.950 679.800 841.050 681.900 ;
        RECT 841.950 679.800 844.050 681.900 ;
        RECT 829.950 676.950 832.050 679.050 ;
        RECT 836.400 678.750 837.600 679.500 ;
        RECT 826.950 658.950 829.050 661.050 ;
        RECT 806.400 649.500 807.600 651.000 ;
        RECT 821.400 649.500 822.600 651.600 ;
        RECT 826.950 651.000 829.050 655.050 ;
        RECT 830.400 652.050 831.450 676.950 ;
        RECT 835.950 676.650 838.050 678.750 ;
        RECT 842.400 677.400 843.600 679.500 ;
        RECT 842.400 673.050 843.450 677.400 ;
        RECT 841.950 670.950 844.050 673.050 ;
        RECT 841.950 661.950 844.050 664.050 ;
        RECT 835.950 658.950 838.050 661.050 ;
        RECT 832.950 652.950 835.050 655.050 ;
        RECT 827.400 649.500 828.600 651.000 ;
        RECT 829.950 649.950 832.050 652.050 ;
        RECT 802.950 647.100 805.050 649.200 ;
        RECT 805.950 647.100 808.050 649.200 ;
        RECT 808.950 647.100 811.050 649.200 ;
        RECT 817.950 647.100 820.050 649.200 ;
        RECT 820.950 647.100 823.050 649.200 ;
        RECT 823.950 647.100 826.050 649.200 ;
        RECT 826.950 647.100 829.050 649.200 ;
        RECT 803.400 644.400 804.600 646.800 ;
        RECT 786.000 636.900 789.000 637.050 ;
        RECT 784.950 634.950 790.050 636.900 ;
        RECT 796.950 634.950 799.050 637.050 ;
        RECT 799.950 634.950 802.050 640.050 ;
        RECT 803.400 637.050 804.450 644.400 ;
        RECT 805.950 643.950 808.050 646.050 ;
        RECT 809.400 644.400 810.600 646.800 ;
        RECT 818.400 646.050 819.600 646.800 ;
        RECT 802.950 634.950 805.050 637.050 ;
        RECT 784.950 634.800 787.050 634.950 ;
        RECT 787.950 634.800 790.050 634.950 ;
        RECT 769.950 628.950 772.050 631.050 ;
        RECT 751.950 613.950 754.050 616.050 ;
        RECT 763.950 613.950 766.050 616.050 ;
        RECT 718.950 607.950 721.050 610.050 ;
        RECT 719.400 606.600 720.450 607.950 ;
        RECT 719.400 604.200 720.600 606.600 ;
        RECT 724.950 604.950 727.050 607.050 ;
        RECT 733.950 604.950 736.050 607.050 ;
        RECT 742.950 606.000 745.050 610.050 ;
        RECT 725.400 604.200 726.600 604.950 ;
        RECT 718.950 601.800 721.050 603.900 ;
        RECT 721.950 601.800 724.050 603.900 ;
        RECT 724.950 601.800 727.050 603.900 ;
        RECT 727.950 601.800 730.050 603.900 ;
        RECT 685.950 595.950 688.050 598.050 ;
        RECT 688.950 595.950 691.050 598.050 ;
        RECT 691.950 595.950 694.050 598.050 ;
        RECT 694.950 595.950 697.050 598.050 ;
        RECT 682.950 574.950 685.050 577.050 ;
        RECT 622.950 568.800 625.050 570.900 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 631.950 568.950 634.050 571.050 ;
        RECT 634.950 568.950 637.050 571.050 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 646.950 568.950 649.050 571.050 ;
        RECT 652.950 568.950 655.050 571.050 ;
        RECT 619.950 559.950 622.050 562.050 ;
        RECT 607.950 547.950 610.050 550.050 ;
        RECT 623.400 544.050 624.450 568.800 ;
        RECT 625.950 565.950 628.050 568.050 ;
        RECT 632.400 566.400 633.600 568.650 ;
        RECT 626.400 547.050 627.450 565.950 ;
        RECT 632.400 559.050 633.450 566.400 ;
        RECT 637.950 565.950 640.050 568.050 ;
        RECT 644.400 566.400 645.600 568.650 ;
        RECT 638.400 562.050 639.450 565.950 ;
        RECT 644.400 562.050 645.450 566.400 ;
        RECT 649.950 565.950 652.050 568.050 ;
        RECT 653.400 567.000 654.600 568.650 ;
        RECT 637.950 559.950 640.050 562.050 ;
        RECT 643.950 559.950 646.050 562.050 ;
        RECT 631.950 556.950 634.050 559.050 ;
        RECT 634.950 553.950 637.050 556.050 ;
        RECT 631.950 550.950 634.050 553.050 ;
        RECT 625.950 544.950 628.050 547.050 ;
        RECT 604.950 541.950 607.050 544.050 ;
        RECT 610.950 541.950 613.050 544.050 ;
        RECT 622.950 541.950 625.050 544.050 ;
        RECT 611.400 529.050 612.450 541.950 ;
        RECT 632.400 541.050 633.450 550.950 ;
        RECT 631.950 538.950 634.050 541.050 ;
        RECT 619.950 536.400 622.050 538.500 ;
        RECT 610.950 526.950 613.050 529.050 ;
        RECT 616.950 527.100 619.050 529.200 ;
        RECT 611.400 526.200 612.600 526.950 ;
        RECT 617.400 526.350 618.600 527.100 ;
        RECT 604.950 523.800 607.050 525.900 ;
        RECT 607.950 523.800 610.050 525.900 ;
        RECT 610.950 523.800 613.050 525.900 ;
        RECT 616.950 523.950 619.050 526.050 ;
        RECT 608.400 521.400 609.600 523.500 ;
        RECT 604.950 517.950 607.050 520.050 ;
        RECT 605.400 508.050 606.450 517.950 ;
        RECT 608.400 511.050 609.450 521.400 ;
        RECT 620.700 516.600 621.900 536.400 ;
        RECT 626.400 528.450 627.600 528.600 ;
        RECT 626.400 527.400 633.450 528.450 ;
        RECT 626.400 526.350 627.600 527.400 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 619.950 514.500 622.050 516.600 ;
        RECT 607.950 508.950 610.050 511.050 ;
        RECT 604.950 505.950 607.050 508.050 ;
        RECT 598.950 502.950 601.050 505.050 ;
        RECT 608.400 499.200 609.450 508.950 ;
        RECT 632.400 508.050 633.450 527.400 ;
        RECT 622.950 505.950 625.050 508.050 ;
        RECT 631.950 505.950 634.050 508.050 ;
        RECT 613.950 499.950 616.050 502.050 ;
        RECT 595.950 496.950 598.050 499.050 ;
        RECT 601.950 496.950 604.050 499.050 ;
        RECT 607.950 497.100 610.050 499.200 ;
        RECT 589.950 494.100 592.050 496.200 ;
        RECT 590.400 493.350 591.600 494.100 ;
        RECT 586.950 490.950 589.050 493.050 ;
        RECT 589.950 490.950 592.050 493.050 ;
        RECT 595.950 490.950 598.050 493.050 ;
        RECT 583.950 487.950 586.050 490.050 ;
        RECT 587.400 488.400 588.600 490.650 ;
        RECT 596.400 488.400 597.600 490.650 ;
        RECT 584.400 484.050 585.450 487.950 ;
        RECT 583.950 481.950 586.050 484.050 ;
        RECT 583.950 478.800 586.050 480.900 ;
        RECT 580.950 475.950 583.050 478.050 ;
        RECT 584.400 471.450 585.450 478.800 ;
        RECT 587.400 478.050 588.450 488.400 ;
        RECT 586.950 475.950 589.050 478.050 ;
        RECT 584.400 470.400 588.450 471.450 ;
        RECT 571.950 463.950 574.050 466.050 ;
        RECT 572.400 451.200 573.450 463.950 ;
        RECT 587.400 463.050 588.450 470.400 ;
        RECT 586.950 460.950 589.050 463.050 ;
        RECT 582.000 459.450 586.050 460.050 ;
        RECT 581.400 457.950 586.050 459.450 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 511.950 445.950 514.050 448.050 ;
        RECT 514.950 445.950 517.050 448.050 ;
        RECT 517.950 445.950 520.050 448.050 ;
        RECT 502.950 442.800 505.050 444.900 ;
        RECT 512.400 443.400 513.600 445.650 ;
        RECT 518.400 444.900 519.600 445.650 ;
        RECT 512.400 439.050 513.450 443.400 ;
        RECT 517.950 442.800 520.050 444.900 ;
        RECT 524.400 444.750 525.450 448.950 ;
        RECT 533.400 448.200 534.600 450.600 ;
        RECT 545.400 448.350 546.600 450.600 ;
        RECT 551.400 448.350 552.600 450.600 ;
        RECT 556.950 449.100 559.050 451.200 ;
        RECT 562.950 449.100 565.050 451.200 ;
        RECT 571.950 449.100 574.050 451.200 ;
        RECT 563.400 448.350 564.600 449.100 ;
        RECT 572.400 448.350 573.600 449.100 ;
        RECT 529.950 445.800 532.050 447.900 ;
        RECT 532.950 445.800 535.050 447.900 ;
        RECT 544.950 445.950 547.050 448.050 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 550.950 445.950 553.050 448.050 ;
        RECT 553.950 445.950 556.050 448.050 ;
        RECT 562.950 445.950 565.050 448.050 ;
        RECT 565.950 445.950 568.050 448.050 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 530.400 444.750 531.600 445.500 ;
        RECT 511.950 436.950 514.050 439.050 ;
        RECT 485.400 431.400 489.450 432.450 ;
        RECT 481.950 413.100 484.050 415.200 ;
        RECT 482.400 410.400 483.600 412.800 ;
        RECT 482.400 406.050 483.450 410.400 ;
        RECT 488.400 406.050 489.450 431.400 ;
        RECT 499.950 430.950 502.050 433.050 ;
        RECT 518.400 427.050 519.450 442.800 ;
        RECT 523.950 442.650 526.050 444.750 ;
        RECT 529.950 442.650 532.050 444.750 ;
        RECT 548.400 443.400 549.600 445.650 ;
        RECT 554.400 444.900 555.600 445.650 ;
        RECT 566.400 444.900 567.600 445.650 ;
        RECT 581.400 444.900 582.450 457.950 ;
        RECT 586.950 450.000 589.050 454.050 ;
        RECT 587.400 448.350 588.600 450.000 ;
        RECT 586.950 445.950 589.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 590.400 444.900 591.600 445.650 ;
        RECT 524.400 430.050 525.450 442.650 ;
        RECT 523.950 427.950 526.050 430.050 ;
        RECT 517.950 424.950 520.050 427.050 ;
        RECT 548.400 418.350 549.450 443.400 ;
        RECT 553.950 442.800 556.050 444.900 ;
        RECT 565.950 442.800 568.050 444.900 ;
        RECT 580.950 442.800 583.050 444.900 ;
        RECT 589.950 442.800 592.050 444.900 ;
        RECT 565.950 421.950 568.050 424.050 ;
        RECT 589.950 421.950 592.050 424.050 ;
        RECT 547.950 416.250 550.050 418.350 ;
        RECT 556.950 416.250 559.050 418.350 ;
        RECT 566.400 418.050 567.450 421.950 ;
        RECT 557.400 415.500 558.600 416.250 ;
        RECT 565.950 415.950 568.050 418.050 ;
        RECT 571.950 416.100 574.050 418.200 ;
        RECT 590.400 417.600 591.450 421.950 ;
        RECT 572.400 415.350 573.600 416.100 ;
        RECT 590.400 415.350 591.600 417.600 ;
        RECT 596.400 417.450 597.450 488.400 ;
        RECT 602.400 481.050 603.450 496.950 ;
        RECT 607.950 493.950 610.050 496.050 ;
        RECT 614.400 495.600 615.450 499.950 ;
        RECT 608.400 493.350 609.600 493.950 ;
        RECT 614.400 493.350 615.600 495.600 ;
        RECT 607.950 490.950 610.050 493.050 ;
        RECT 610.950 490.950 613.050 493.050 ;
        RECT 613.950 490.950 616.050 493.050 ;
        RECT 616.950 490.950 619.050 493.050 ;
        RECT 611.400 489.900 612.600 490.650 ;
        RECT 610.950 487.800 613.050 489.900 ;
        RECT 617.400 488.400 618.600 490.650 ;
        RECT 617.400 481.050 618.450 488.400 ;
        RECT 623.400 484.050 624.450 505.950 ;
        RECT 635.400 504.450 636.450 553.950 ;
        RECT 640.950 537.300 643.050 539.400 ;
        RECT 640.950 533.700 642.150 537.300 ;
        RECT 640.950 531.600 643.050 533.700 ;
        RECT 650.400 532.050 651.450 565.950 ;
        RECT 652.950 562.950 655.050 567.000 ;
        RECT 655.950 565.950 658.050 568.050 ;
        RECT 640.950 516.600 642.150 531.600 ;
        RECT 649.950 529.950 652.050 532.050 ;
        RECT 656.400 529.050 657.450 565.950 ;
        RECT 659.400 562.050 660.450 571.800 ;
        RECT 668.400 571.500 669.600 573.600 ;
        RECT 674.400 571.500 675.600 573.600 ;
        RECT 676.950 571.950 679.050 574.050 ;
        RECT 686.400 573.450 687.450 595.950 ;
        RECT 689.400 592.050 690.450 595.950 ;
        RECT 695.400 592.050 696.450 595.950 ;
        RECT 688.950 589.950 691.050 592.050 ;
        RECT 694.950 589.950 697.050 592.050 ;
        RECT 707.400 586.050 708.450 599.400 ;
        RECT 712.950 598.650 715.050 600.750 ;
        RECT 722.400 600.000 723.600 601.500 ;
        RECT 721.950 595.950 724.050 600.000 ;
        RECT 728.400 599.400 729.600 601.500 ;
        RECT 728.400 586.050 729.450 599.400 ;
        RECT 706.950 583.950 709.050 586.050 ;
        RECT 712.950 583.950 715.050 586.050 ;
        RECT 727.950 583.950 730.050 586.050 ;
        RECT 691.950 580.950 694.050 583.050 ;
        RECT 692.400 577.050 693.450 580.950 ;
        RECT 713.400 577.050 714.450 583.950 ;
        RECT 718.950 577.950 721.050 580.050 ;
        RECT 683.400 572.400 687.450 573.450 ;
        RECT 691.950 573.000 694.050 577.050 ;
        RECT 712.950 574.950 715.050 577.050 ;
        RECT 664.950 569.100 667.050 571.200 ;
        RECT 667.950 569.100 670.050 571.200 ;
        RECT 670.950 569.100 673.050 571.200 ;
        RECT 673.950 569.100 676.050 571.200 ;
        RECT 665.400 566.400 666.600 568.800 ;
        RECT 671.400 567.000 672.600 568.800 ;
        RECT 658.950 559.950 661.050 562.050 ;
        RECT 665.400 559.050 666.450 566.400 ;
        RECT 670.950 562.950 673.050 567.000 ;
        RECT 676.950 565.950 679.050 568.050 ;
        RECT 670.950 559.800 673.050 561.900 ;
        RECT 664.950 556.950 667.050 559.050 ;
        RECT 664.950 547.950 667.050 550.050 ;
        RECT 665.400 529.200 666.450 547.950 ;
        RECT 667.950 529.950 670.050 532.050 ;
        RECT 649.950 526.800 652.050 528.900 ;
        RECT 655.950 526.950 658.050 529.050 ;
        RECT 664.950 527.100 667.050 529.200 ;
        RECT 643.950 523.950 646.050 526.050 ;
        RECT 644.400 522.450 645.600 523.650 ;
        RECT 650.400 522.450 651.450 526.800 ;
        RECT 656.400 526.200 657.600 526.950 ;
        RECT 655.950 523.800 658.050 525.900 ;
        RECT 658.950 523.800 661.050 525.900 ;
        RECT 661.950 523.800 664.050 525.900 ;
        RECT 644.400 521.400 651.450 522.450 ;
        RECT 652.950 517.950 655.050 523.050 ;
        RECT 659.400 522.750 660.600 523.500 ;
        RECT 658.950 520.650 661.050 522.750 ;
        RECT 640.950 514.500 643.050 516.600 ;
        RECT 668.400 511.050 669.450 529.950 ;
        RECT 671.400 529.050 672.450 559.800 ;
        RECT 677.400 547.050 678.450 565.950 ;
        RECT 676.950 544.950 679.050 547.050 ;
        RECT 683.400 529.200 684.450 572.400 ;
        RECT 692.400 571.350 693.600 573.000 ;
        RECT 697.950 571.950 700.050 574.050 ;
        RECT 706.950 572.100 709.050 574.200 ;
        RECT 713.400 573.600 714.450 574.950 ;
        RECT 688.950 568.950 691.050 571.050 ;
        RECT 691.950 568.950 694.050 571.050 ;
        RECT 689.400 567.900 690.600 568.650 ;
        RECT 688.950 565.800 691.050 567.900 ;
        RECT 698.400 562.050 699.450 571.950 ;
        RECT 707.400 571.350 708.600 572.100 ;
        RECT 713.400 571.350 714.600 573.600 ;
        RECT 703.950 568.950 706.050 571.050 ;
        RECT 706.950 568.950 709.050 571.050 ;
        RECT 709.950 568.950 712.050 571.050 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 704.400 567.900 705.600 568.650 ;
        RECT 710.400 567.900 711.600 568.650 ;
        RECT 703.950 565.800 706.050 567.900 ;
        RECT 709.950 565.800 712.050 567.900 ;
        RECT 697.950 559.950 700.050 562.050 ;
        RECT 719.400 559.050 720.450 577.950 ;
        RECT 728.400 573.600 729.450 583.950 ;
        RECT 734.400 580.050 735.450 604.950 ;
        RECT 743.400 604.350 744.600 606.000 ;
        RECT 748.950 604.950 751.050 607.050 ;
        RECT 754.950 604.950 757.050 607.050 ;
        RECT 760.950 606.000 763.050 610.050 ;
        RECT 739.950 601.950 742.050 604.050 ;
        RECT 742.950 601.950 745.050 604.050 ;
        RECT 740.400 599.400 741.600 601.650 ;
        RECT 733.950 577.950 736.050 580.050 ;
        RECT 740.400 577.050 741.450 599.400 ;
        RECT 745.950 583.950 748.050 586.050 ;
        RECT 739.950 574.950 742.050 577.050 ;
        RECT 746.400 573.600 747.450 583.950 ;
        RECT 749.400 583.050 750.450 604.950 ;
        RECT 755.400 604.200 756.600 604.950 ;
        RECT 761.400 604.200 762.600 606.000 ;
        RECT 754.950 601.800 757.050 603.900 ;
        RECT 757.950 601.800 760.050 603.900 ;
        RECT 760.950 601.800 763.050 603.900 ;
        RECT 763.950 601.800 766.050 603.900 ;
        RECT 758.400 599.400 759.600 601.500 ;
        RECT 764.400 599.400 765.600 601.500 ;
        RECT 758.400 589.050 759.450 599.400 ;
        RECT 757.950 586.950 760.050 589.050 ;
        RECT 748.950 582.450 751.050 583.050 ;
        RECT 748.950 581.400 753.450 582.450 ;
        RECT 748.950 580.950 751.050 581.400 ;
        RECT 752.400 574.050 753.450 581.400 ;
        RECT 728.400 571.350 729.600 573.600 ;
        RECT 740.400 573.450 741.600 573.600 ;
        RECT 734.400 572.400 741.600 573.450 ;
        RECT 724.950 568.950 727.050 571.050 ;
        RECT 727.950 568.950 730.050 571.050 ;
        RECT 725.400 567.900 726.600 568.650 ;
        RECT 724.950 565.800 727.050 567.900 ;
        RECT 718.950 556.950 721.050 559.050 ;
        RECT 727.950 550.950 730.050 553.050 ;
        RECT 728.400 541.050 729.450 550.950 ;
        RECT 734.400 547.050 735.450 572.400 ;
        RECT 740.400 571.500 741.600 572.400 ;
        RECT 746.400 571.500 747.600 573.600 ;
        RECT 751.950 571.950 754.050 574.050 ;
        RECT 764.400 573.600 765.450 599.400 ;
        RECT 770.400 598.050 771.450 628.950 ;
        RECT 802.950 625.950 805.050 628.050 ;
        RECT 772.950 619.950 775.050 622.050 ;
        RECT 784.950 619.950 787.050 622.050 ;
        RECT 769.950 595.950 772.050 598.050 ;
        RECT 773.400 595.050 774.450 619.950 ;
        RECT 785.400 607.050 786.450 619.950 ;
        RECT 790.950 613.950 793.050 616.050 ;
        RECT 778.950 604.950 781.050 607.050 ;
        RECT 784.950 604.950 787.050 607.050 ;
        RECT 779.400 604.200 780.600 604.950 ;
        RECT 785.400 604.200 786.600 604.950 ;
        RECT 778.950 601.800 781.050 603.900 ;
        RECT 781.950 601.800 784.050 603.900 ;
        RECT 784.950 601.800 787.050 603.900 ;
        RECT 782.400 599.400 783.600 601.500 ;
        RECT 772.950 592.950 775.050 595.050 ;
        RECT 775.950 577.950 778.050 580.050 ;
        RECT 772.950 574.950 775.050 577.050 ;
        RECT 764.400 571.500 765.600 573.600 ;
        RECT 739.950 569.100 742.050 571.200 ;
        RECT 742.950 569.100 745.050 571.200 ;
        RECT 745.950 569.100 748.050 571.200 ;
        RECT 748.950 569.100 751.050 571.200 ;
        RECT 757.950 569.100 760.050 571.200 ;
        RECT 763.950 569.100 766.050 571.200 ;
        RECT 766.950 569.100 769.050 571.200 ;
        RECT 743.400 568.050 744.600 568.800 ;
        RECT 749.400 568.050 750.600 568.800 ;
        RECT 742.950 565.950 745.050 568.050 ;
        RECT 749.400 566.400 754.050 568.050 ;
        RECT 750.000 565.950 754.050 566.400 ;
        RECT 758.400 566.400 759.600 568.800 ;
        RECT 767.400 566.400 768.600 568.800 ;
        RECT 758.400 562.050 759.450 566.400 ;
        RECT 767.400 562.050 768.450 566.400 ;
        RECT 757.950 559.950 760.050 562.050 ;
        RECT 766.950 559.950 769.050 562.050 ;
        RECT 748.950 556.950 751.050 559.050 ;
        RECT 733.950 544.950 736.050 547.050 ;
        RECT 727.950 538.950 730.050 541.050 ;
        RECT 670.950 526.950 673.050 529.050 ;
        RECT 676.950 527.100 679.050 529.200 ;
        RECT 682.950 527.100 685.050 529.200 ;
        RECT 677.400 526.350 678.600 527.100 ;
        RECT 683.400 526.350 684.600 527.100 ;
        RECT 688.800 526.950 690.900 529.050 ;
        RECT 691.950 527.100 694.050 529.200 ;
        RECT 697.950 527.100 700.050 529.200 ;
        RECT 703.950 528.000 706.050 532.050 ;
        RECT 718.950 528.000 721.050 532.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 679.950 523.950 682.050 526.050 ;
        RECT 682.950 523.950 685.050 526.050 ;
        RECT 674.400 523.050 675.600 523.650 ;
        RECT 670.950 521.400 675.600 523.050 ;
        RECT 680.400 522.900 681.600 523.650 ;
        RECT 670.950 520.950 675.000 521.400 ;
        RECT 671.400 514.050 672.450 520.950 ;
        RECT 679.950 520.800 682.050 522.900 ;
        RECT 682.950 517.950 688.050 520.050 ;
        RECT 670.950 511.950 673.050 514.050 ;
        RECT 667.950 508.950 670.050 511.050 ;
        RECT 676.950 505.950 679.050 508.050 ;
        RECT 632.400 503.400 636.450 504.450 ;
        RECT 632.400 496.050 633.450 503.400 ;
        RECT 634.950 499.950 637.050 502.050 ;
        RECT 677.400 501.600 678.450 505.950 ;
        RECT 631.950 493.950 634.050 496.050 ;
        RECT 635.400 495.600 636.450 499.950 ;
        RECT 670.650 497.400 672.750 499.500 ;
        RECT 677.400 498.900 678.600 501.600 ;
        RECT 635.400 493.500 636.600 495.600 ;
        RECT 643.950 493.950 646.050 496.050 ;
        RECT 655.950 494.250 658.050 496.350 ;
        RECT 628.950 491.100 631.050 493.200 ;
        RECT 634.950 491.100 637.050 493.200 ;
        RECT 637.950 491.100 640.050 493.200 ;
        RECT 629.400 488.400 630.600 490.800 ;
        RECT 638.400 490.050 639.600 490.800 ;
        RECT 622.950 481.950 625.050 484.050 ;
        RECT 601.950 478.950 604.050 481.050 ;
        RECT 616.950 478.950 619.050 481.050 ;
        RECT 629.400 466.050 630.450 488.400 ;
        RECT 637.950 487.950 640.050 490.050 ;
        RECT 634.950 481.950 637.050 484.050 ;
        RECT 631.950 478.950 634.050 481.050 ;
        RECT 632.400 469.050 633.450 478.950 ;
        RECT 631.950 466.950 634.050 469.050 ;
        RECT 628.950 463.950 631.050 466.050 ;
        RECT 604.950 454.950 607.050 457.050 ;
        RECT 605.400 450.600 606.450 454.950 ;
        RECT 605.400 448.200 606.600 450.600 ;
        RECT 610.950 448.950 613.050 451.050 ;
        RECT 616.950 448.950 619.050 451.050 ;
        RECT 625.950 450.000 628.050 454.050 ;
        RECT 632.400 450.600 633.450 466.950 ;
        RECT 635.400 463.050 636.450 481.950 ;
        RECT 644.400 478.050 645.450 493.950 ;
        RECT 656.400 493.500 657.600 494.250 ;
        RECT 652.950 491.100 655.050 493.200 ;
        RECT 655.950 491.100 658.050 493.200 ;
        RECT 658.950 491.100 661.050 493.200 ;
        RECT 667.950 491.100 670.050 493.200 ;
        RECT 653.400 490.050 654.600 490.800 ;
        RECT 659.400 490.050 660.600 490.800 ;
        RECT 652.950 487.950 655.050 490.050 ;
        RECT 658.950 487.950 661.050 490.050 ;
        RECT 668.400 489.000 669.600 491.100 ;
        RECT 653.400 486.450 654.450 487.950 ;
        RECT 658.950 486.450 661.050 486.900 ;
        RECT 653.400 485.400 661.050 486.450 ;
        RECT 658.950 484.800 661.050 485.400 ;
        RECT 667.950 484.950 670.050 489.000 ;
        RECT 671.400 484.800 672.300 497.400 ;
        RECT 677.250 496.800 679.350 498.900 ;
        RECT 680.700 497.100 682.800 499.200 ;
        RECT 673.200 495.000 675.300 495.900 ;
        RECT 673.200 493.800 680.250 495.000 ;
        RECT 678.150 492.900 680.250 493.800 ;
        RECT 673.200 492.000 675.300 492.900 ;
        RECT 681.150 492.000 682.050 497.100 ;
        RECT 683.400 493.200 684.600 495.600 ;
        RECT 673.200 491.100 682.050 492.000 ;
        RECT 682.950 493.050 685.050 493.200 ;
        RECT 682.950 491.100 688.050 493.050 ;
        RECT 673.200 490.800 675.300 491.100 ;
        RECT 677.250 488.100 679.350 490.200 ;
        RECT 677.400 485.400 678.600 488.100 ;
        RECT 671.100 482.700 673.200 484.800 ;
        RECT 681.150 484.500 682.050 491.100 ;
        RECT 685.050 490.950 688.050 491.100 ;
        RECT 680.100 482.400 682.200 484.500 ;
        RECT 643.950 475.950 646.050 478.050 ;
        RECT 673.950 475.950 676.050 478.050 ;
        RECT 643.950 466.950 646.050 469.050 ;
        RECT 634.950 460.950 637.050 463.050 ;
        RECT 644.400 460.050 645.450 466.950 ;
        RECT 670.950 460.950 673.050 463.050 ;
        RECT 643.950 457.950 646.050 460.050 ;
        RECT 658.950 454.950 661.050 457.050 ;
        RECT 637.950 451.950 640.050 454.050 ;
        RECT 611.400 448.200 612.600 448.950 ;
        RECT 601.950 445.800 604.050 447.900 ;
        RECT 604.950 445.800 607.050 447.900 ;
        RECT 607.950 445.800 610.050 447.900 ;
        RECT 610.950 445.800 613.050 447.900 ;
        RECT 602.400 443.400 603.600 445.500 ;
        RECT 608.400 443.400 609.600 445.500 ;
        RECT 602.400 418.050 603.450 443.400 ;
        RECT 604.950 423.450 607.050 424.050 ;
        RECT 608.400 423.450 609.450 443.400 ;
        RECT 617.400 433.050 618.450 448.950 ;
        RECT 626.400 448.200 627.600 450.000 ;
        RECT 632.400 448.200 633.600 450.600 ;
        RECT 622.950 445.800 625.050 447.900 ;
        RECT 625.950 445.800 628.050 447.900 ;
        RECT 628.950 445.800 631.050 447.900 ;
        RECT 631.950 445.800 634.050 447.900 ;
        RECT 623.400 443.400 624.600 445.500 ;
        RECT 629.400 444.750 630.600 445.500 ;
        RECT 619.950 436.950 622.050 439.050 ;
        RECT 610.950 430.950 613.050 433.050 ;
        RECT 616.950 430.950 619.050 433.050 ;
        RECT 604.950 422.400 609.450 423.450 ;
        RECT 604.950 421.950 607.050 422.400 ;
        RECT 596.400 416.400 600.450 417.450 ;
        RECT 502.950 413.100 505.050 415.200 ;
        RECT 517.950 413.100 520.050 415.200 ;
        RECT 538.950 413.100 541.050 415.200 ;
        RECT 553.950 413.100 556.050 415.200 ;
        RECT 556.950 413.100 559.050 415.200 ;
        RECT 562.950 413.100 565.050 415.200 ;
        RECT 571.950 412.950 574.050 415.050 ;
        RECT 577.950 412.950 580.050 415.050 ;
        RECT 589.950 412.950 592.050 415.050 ;
        RECT 592.950 412.950 595.050 415.050 ;
        RECT 539.400 410.400 540.600 412.800 ;
        RECT 554.400 412.050 555.600 412.800 ;
        RECT 481.950 403.950 484.050 406.050 ;
        RECT 487.950 403.950 490.050 406.050 ;
        RECT 484.950 385.950 487.050 388.050 ;
        RECT 539.400 387.450 540.450 410.400 ;
        RECT 553.950 409.950 556.050 412.050 ;
        RECT 563.400 410.400 564.600 412.800 ;
        RECT 563.400 406.050 564.450 410.400 ;
        RECT 565.950 409.950 568.050 412.050 ;
        RECT 578.400 411.000 579.600 412.650 ;
        RECT 593.400 411.900 594.600 412.650 ;
        RECT 562.950 403.950 565.050 406.050 ;
        RECT 541.950 387.450 544.050 388.050 ;
        RECT 539.400 386.400 544.050 387.450 ;
        RECT 541.950 385.950 544.050 386.400 ;
        RECT 449.400 370.350 450.600 370.950 ;
        RECT 458.400 370.200 459.600 370.950 ;
        RECT 464.400 370.200 465.600 370.950 ;
        RECT 418.950 367.800 421.050 369.900 ;
        RECT 421.950 367.800 424.050 369.900 ;
        RECT 427.950 367.800 430.050 369.900 ;
        RECT 439.950 367.950 442.050 370.050 ;
        RECT 445.950 367.950 448.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 457.950 367.800 460.050 369.900 ;
        RECT 460.950 367.800 463.050 369.900 ;
        RECT 463.950 367.800 466.050 369.900 ;
        RECT 422.400 366.750 423.600 367.500 ;
        RECT 421.950 364.650 424.050 366.750 ;
        RECT 436.950 364.950 439.050 367.050 ;
        RECT 446.400 366.000 447.600 367.650 ;
        RECT 412.950 361.950 415.050 364.050 ;
        RECT 422.400 358.050 423.450 364.650 ;
        RECT 421.950 355.950 424.050 358.050 ;
        RECT 406.950 349.950 409.050 352.050 ;
        RECT 430.950 349.950 433.050 352.050 ;
        RECT 391.950 338.100 394.050 340.200 ;
        RECT 392.400 337.350 393.600 338.100 ;
        RECT 355.950 334.950 358.050 337.050 ;
        RECT 358.950 334.950 361.050 337.050 ;
        RECT 361.950 334.950 364.050 337.050 ;
        RECT 370.950 334.950 373.050 337.050 ;
        RECT 373.950 334.950 376.050 337.050 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 379.950 334.950 382.050 337.050 ;
        RECT 385.950 334.950 388.050 337.050 ;
        RECT 391.950 334.950 394.050 337.050 ;
        RECT 397.950 334.950 400.050 337.050 ;
        RECT 359.400 333.900 360.600 334.650 ;
        RECT 358.950 331.800 361.050 333.900 ;
        RECT 367.950 331.950 370.050 334.050 ;
        RECT 374.400 333.900 375.600 334.650 ;
        RECT 352.950 292.950 355.050 295.050 ;
        RECT 355.950 292.950 358.050 298.050 ;
        RECT 361.950 294.000 364.050 298.050 ;
        RECT 368.400 295.050 369.450 331.950 ;
        RECT 373.950 331.800 376.050 333.900 ;
        RECT 380.400 333.000 381.600 334.650 ;
        RECT 379.950 328.950 382.050 333.000 ;
        RECT 388.950 331.950 391.050 334.050 ;
        RECT 398.400 332.400 399.600 334.650 ;
        RECT 385.950 328.950 388.050 331.050 ;
        RECT 370.950 298.950 373.050 301.050 ;
        RECT 353.400 289.050 354.450 292.950 ;
        RECT 362.400 292.350 363.600 294.000 ;
        RECT 367.950 292.950 370.050 295.050 ;
        RECT 358.950 289.950 361.050 292.050 ;
        RECT 361.950 289.950 364.050 292.050 ;
        RECT 364.950 289.950 367.050 292.050 ;
        RECT 352.950 286.950 355.050 289.050 ;
        RECT 355.950 286.950 358.050 289.050 ;
        RECT 359.400 288.900 360.600 289.650 ;
        RECT 365.400 288.900 366.600 289.650 ;
        RECT 356.400 262.050 357.450 286.950 ;
        RECT 358.950 286.800 361.050 288.900 ;
        RECT 364.950 286.800 367.050 288.900 ;
        RECT 365.400 280.050 366.450 286.800 ;
        RECT 364.950 277.950 367.050 280.050 ;
        RECT 367.950 262.950 370.050 265.050 ;
        RECT 355.950 261.450 358.050 262.050 ;
        RECT 359.400 261.450 360.600 261.600 ;
        RECT 350.400 260.400 354.450 261.450 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 344.400 254.400 345.600 256.650 ;
        RECT 340.950 235.950 343.050 238.050 ;
        RECT 337.950 232.950 340.050 235.050 ;
        RECT 311.400 214.350 312.600 215.100 ;
        RECT 317.400 214.350 318.600 216.600 ;
        RECT 322.800 214.950 324.900 217.050 ;
        RECT 325.950 215.100 328.050 217.200 ;
        RECT 326.400 214.350 327.600 215.100 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 319.950 211.950 322.050 214.050 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 314.400 209.400 315.600 211.650 ;
        RECT 320.400 210.900 321.600 211.650 ;
        RECT 307.950 199.950 310.050 202.050 ;
        RECT 304.950 190.950 307.050 193.050 ;
        RECT 308.400 187.050 309.450 199.950 ;
        RECT 307.950 184.950 310.050 187.050 ;
        RECT 295.950 181.950 298.050 184.050 ;
        RECT 304.950 182.100 307.050 184.200 ;
        RECT 310.950 182.100 313.050 184.200 ;
        RECT 314.400 183.450 315.450 209.400 ;
        RECT 319.950 208.800 322.050 210.900 ;
        RECT 329.700 204.600 330.900 224.400 ;
        RECT 334.950 223.950 337.050 226.050 ;
        RECT 335.400 216.450 336.600 216.600 ;
        RECT 338.400 216.450 339.450 232.950 ;
        RECT 341.400 220.050 342.450 235.950 ;
        RECT 344.400 229.050 345.450 254.400 ;
        RECT 353.400 235.050 354.450 260.400 ;
        RECT 355.950 260.400 360.600 261.450 ;
        RECT 355.950 259.950 358.050 260.400 ;
        RECT 359.400 259.350 360.600 260.400 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 362.400 255.900 363.600 256.650 ;
        RECT 361.950 253.800 364.050 255.900 ;
        RECT 358.950 235.950 361.050 238.050 ;
        RECT 352.950 232.950 355.050 235.050 ;
        RECT 343.950 226.950 346.050 229.050 ;
        RECT 349.950 225.300 352.050 227.400 ;
        RECT 343.950 220.950 346.050 223.050 ;
        RECT 349.950 221.700 351.150 225.300 ;
        RECT 355.950 223.950 358.050 226.050 ;
        RECT 340.950 217.950 343.050 220.050 ;
        RECT 335.400 215.400 339.450 216.450 ;
        RECT 335.400 214.350 336.600 215.400 ;
        RECT 334.950 211.950 337.050 214.050 ;
        RECT 328.950 202.500 331.050 204.600 ;
        RECT 341.400 202.050 342.450 217.950 ;
        RECT 340.950 199.950 343.050 202.050 ;
        RECT 344.400 196.050 345.450 220.950 ;
        RECT 349.950 219.600 352.050 221.700 ;
        RECT 349.950 204.600 351.150 219.600 ;
        RECT 356.400 217.050 357.450 223.950 ;
        RECT 355.950 214.950 358.050 217.050 ;
        RECT 359.400 216.450 360.450 235.950 ;
        RECT 362.400 232.050 363.450 253.800 ;
        RECT 368.400 232.050 369.450 262.950 ;
        RECT 361.950 229.950 364.050 232.050 ;
        RECT 367.950 229.950 370.050 232.050 ;
        RECT 364.950 224.400 367.050 226.500 ;
        RECT 362.400 216.450 363.600 216.600 ;
        RECT 359.400 215.400 363.600 216.450 ;
        RECT 362.400 214.350 363.600 215.400 ;
        RECT 352.950 211.950 355.050 214.050 ;
        RECT 361.950 211.950 364.050 214.050 ;
        RECT 353.400 210.900 354.600 211.650 ;
        RECT 352.950 208.800 355.050 210.900 ;
        RECT 365.700 204.600 366.900 224.400 ;
        RECT 371.400 220.050 372.450 298.950 ;
        RECT 386.400 295.050 387.450 328.950 ;
        RECT 389.400 301.050 390.450 331.950 ;
        RECT 398.400 322.050 399.450 332.400 ;
        RECT 403.950 331.800 406.050 333.900 ;
        RECT 397.950 319.950 400.050 322.050 ;
        RECT 400.950 310.950 403.050 313.050 ;
        RECT 388.950 298.950 391.050 301.050 ;
        RECT 376.950 292.950 379.050 295.050 ;
        RECT 382.950 292.950 385.050 295.050 ;
        RECT 385.950 292.950 388.050 295.050 ;
        RECT 388.950 292.950 391.050 295.050 ;
        RECT 394.950 292.950 397.050 295.050 ;
        RECT 401.400 294.600 402.450 310.950 ;
        RECT 404.400 295.050 405.450 331.800 ;
        RECT 377.400 292.200 378.600 292.950 ;
        RECT 383.400 292.200 384.600 292.950 ;
        RECT 376.950 289.800 379.050 291.900 ;
        RECT 379.950 289.800 382.050 291.900 ;
        RECT 382.950 289.800 385.050 291.900 ;
        RECT 380.400 287.400 381.600 289.500 ;
        RECT 380.400 268.050 381.450 287.400 ;
        RECT 373.950 265.950 376.050 268.050 ;
        RECT 379.800 265.950 381.900 268.050 ;
        RECT 374.400 262.050 375.450 265.950 ;
        RECT 382.950 264.450 385.050 268.050 ;
        RECT 380.400 264.000 385.050 264.450 ;
        RECT 380.400 263.400 384.450 264.000 ;
        RECT 373.950 259.950 376.050 262.050 ;
        RECT 380.400 261.600 381.450 263.400 ;
        RECT 389.400 262.050 390.450 292.950 ;
        RECT 395.400 292.200 396.600 292.950 ;
        RECT 401.400 292.200 402.600 294.600 ;
        RECT 403.950 292.950 406.050 295.050 ;
        RECT 394.950 289.800 397.050 291.900 ;
        RECT 397.950 289.800 400.050 291.900 ;
        RECT 400.950 289.800 403.050 291.900 ;
        RECT 391.950 285.450 394.050 289.050 ;
        RECT 398.400 288.750 399.600 289.500 ;
        RECT 397.950 286.650 400.050 288.750 ;
        RECT 391.950 285.000 396.450 285.450 ;
        RECT 392.400 284.400 396.450 285.000 ;
        RECT 380.400 259.500 381.600 261.600 ;
        RECT 388.950 259.950 391.050 262.050 ;
        RECT 395.400 261.600 396.450 284.400 ;
        RECT 395.400 259.500 396.600 261.600 ;
        RECT 407.400 261.450 408.450 349.950 ;
        RECT 415.950 343.950 418.050 346.050 ;
        RECT 427.950 343.950 430.050 346.050 ;
        RECT 416.400 339.600 417.450 343.950 ;
        RECT 416.400 337.350 417.600 339.600 ;
        RECT 421.950 338.100 424.050 340.200 ;
        RECT 422.400 337.350 423.600 338.100 ;
        RECT 412.950 334.950 415.050 337.050 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 418.950 334.950 421.050 337.050 ;
        RECT 421.950 334.950 424.050 337.050 ;
        RECT 413.400 333.900 414.600 334.650 ;
        RECT 412.950 331.800 415.050 333.900 ;
        RECT 419.400 333.000 420.600 334.650 ;
        RECT 428.400 334.050 429.450 343.950 ;
        RECT 431.400 340.050 432.450 349.950 ;
        RECT 437.400 343.050 438.450 364.950 ;
        RECT 445.950 361.950 448.050 366.000 ;
        RECT 454.950 364.950 457.050 367.050 ;
        RECT 461.400 365.400 462.600 367.500 ;
        RECT 445.950 344.400 448.050 346.500 ;
        RECT 436.950 340.950 439.050 343.050 ;
        RECT 430.950 337.950 433.050 340.050 ;
        RECT 437.400 339.600 438.450 340.950 ;
        RECT 437.400 337.350 438.600 339.600 ;
        RECT 442.950 339.000 445.050 343.050 ;
        RECT 443.400 337.350 444.600 339.000 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 436.950 334.950 439.050 337.050 ;
        RECT 442.950 334.950 445.050 337.050 ;
        RECT 418.950 328.950 421.050 333.000 ;
        RECT 424.800 331.950 426.900 334.050 ;
        RECT 427.950 331.950 430.050 334.050 ;
        RECT 434.400 333.000 435.600 334.650 ;
        RECT 425.400 313.050 426.450 331.950 ;
        RECT 433.950 328.950 436.050 333.000 ;
        RECT 446.850 329.400 448.050 344.400 ;
        RECT 445.950 327.300 448.050 329.400 ;
        RECT 446.850 323.700 448.050 327.300 ;
        RECT 445.950 321.600 448.050 323.700 ;
        RECT 455.400 322.050 456.450 364.950 ;
        RECT 461.400 358.050 462.450 365.400 ;
        RECT 470.400 364.050 471.450 370.950 ;
        RECT 469.950 361.950 472.050 364.050 ;
        RECT 473.400 358.050 474.450 371.100 ;
        RECT 475.950 370.950 478.050 373.050 ;
        RECT 478.950 371.100 481.050 373.200 ;
        RECT 485.400 372.600 486.450 385.950 ;
        RECT 514.950 381.300 517.050 383.400 ;
        RECT 508.950 378.450 511.050 379.050 ;
        RECT 494.400 377.400 511.050 378.450 ;
        RECT 515.850 377.700 517.050 381.300 ;
        RECT 535.950 380.400 538.050 382.500 ;
        RECT 494.400 373.050 495.450 377.400 ;
        RECT 508.950 376.950 511.050 377.400 ;
        RECT 496.950 375.450 499.050 376.050 ;
        RECT 505.950 375.450 508.050 376.050 ;
        RECT 514.950 375.600 517.050 377.700 ;
        RECT 529.950 376.950 532.050 379.050 ;
        RECT 496.950 374.400 508.050 375.450 ;
        RECT 479.400 370.350 480.600 371.100 ;
        RECT 485.400 370.350 486.600 372.600 ;
        RECT 493.950 370.950 496.050 373.050 ;
        RECT 496.950 372.000 499.050 374.400 ;
        RECT 505.950 373.950 508.050 374.400 ;
        RECT 497.400 370.200 498.600 372.000 ;
        RECT 502.950 370.950 505.050 373.050 ;
        RECT 503.400 370.200 504.600 370.950 ;
        RECT 478.950 367.950 481.050 370.050 ;
        RECT 481.950 367.950 484.050 370.050 ;
        RECT 484.950 367.950 487.050 370.050 ;
        RECT 487.950 367.950 490.050 370.050 ;
        RECT 496.950 367.800 499.050 369.900 ;
        RECT 499.950 367.800 502.050 369.900 ;
        RECT 502.950 367.800 505.050 369.900 ;
        RECT 511.950 367.950 514.050 370.050 ;
        RECT 475.950 364.950 478.050 367.050 ;
        RECT 482.400 366.900 483.600 367.650 ;
        RECT 488.400 366.900 489.600 367.650 ;
        RECT 460.950 355.950 463.050 358.050 ;
        RECT 472.950 355.950 475.050 358.050 ;
        RECT 466.950 344.400 469.050 346.500 ;
        RECT 460.950 334.950 463.050 337.050 ;
        RECT 461.400 333.900 462.600 334.650 ;
        RECT 460.950 331.800 463.050 333.900 ;
        RECT 467.100 324.600 468.300 344.400 ;
        RECT 469.950 334.950 472.050 337.050 ;
        RECT 470.400 333.450 471.600 334.650 ;
        RECT 470.400 332.400 474.450 333.450 ;
        RECT 466.950 322.500 469.050 324.600 ;
        RECT 454.950 319.950 457.050 322.050 ;
        RECT 424.950 310.950 427.050 313.050 ;
        RECT 412.950 293.100 415.050 295.200 ;
        RECT 418.950 294.000 421.050 298.050 ;
        RECT 425.400 295.050 426.450 310.950 ;
        RECT 473.400 310.050 474.450 332.400 ;
        RECT 472.950 307.950 475.050 310.050 ;
        RECT 430.950 301.950 433.050 304.050 ;
        RECT 445.950 303.300 448.050 305.400 ;
        RECT 431.400 295.050 432.450 301.950 ;
        RECT 446.850 299.700 448.050 303.300 ;
        RECT 460.950 301.950 463.050 304.050 ;
        RECT 466.950 302.400 469.050 304.500 ;
        RECT 413.400 292.350 414.600 293.100 ;
        RECT 419.400 292.350 420.600 294.000 ;
        RECT 424.950 292.950 427.050 295.050 ;
        RECT 430.950 292.950 433.050 295.050 ;
        RECT 433.950 294.000 436.050 298.050 ;
        RECT 445.950 297.600 448.050 299.700 ;
        RECT 434.400 292.350 435.600 294.000 ;
        RECT 412.950 289.950 415.050 292.050 ;
        RECT 415.950 289.950 418.050 292.050 ;
        RECT 418.950 289.950 421.050 292.050 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 433.950 289.950 436.050 292.050 ;
        RECT 436.950 289.950 439.050 292.050 ;
        RECT 442.950 289.950 445.050 292.050 ;
        RECT 416.400 287.400 417.600 289.650 ;
        RECT 422.400 288.900 423.600 289.650 ;
        RECT 421.950 288.450 424.050 288.900 ;
        RECT 421.950 287.400 426.450 288.450 ;
        RECT 412.950 283.950 415.050 286.050 ;
        RECT 404.400 260.400 408.450 261.450 ;
        RECT 413.400 261.600 414.450 283.950 ;
        RECT 416.400 283.050 417.450 287.400 ;
        RECT 421.950 286.800 424.050 287.400 ;
        RECT 415.950 280.950 418.050 283.050 ;
        RECT 418.950 265.950 421.050 268.050 ;
        RECT 419.400 262.050 420.450 265.950 ;
        RECT 425.400 265.050 426.450 287.400 ;
        RECT 430.950 286.950 433.050 289.050 ;
        RECT 437.400 287.400 438.600 289.650 ;
        RECT 431.400 283.050 432.450 286.950 ;
        RECT 430.950 280.950 433.050 283.050 ;
        RECT 437.400 277.050 438.450 287.400 ;
        RECT 439.950 286.950 442.050 289.050 ;
        RECT 443.400 288.000 444.600 289.650 ;
        RECT 440.400 280.050 441.450 286.950 ;
        RECT 442.950 283.950 445.050 288.000 ;
        RECT 446.850 282.600 448.050 297.600 ;
        RECT 461.400 294.600 462.450 301.950 ;
        RECT 461.400 292.350 462.600 294.600 ;
        RECT 460.950 289.950 463.050 292.050 ;
        RECT 451.950 283.950 454.050 286.050 ;
        RECT 445.950 280.500 448.050 282.600 ;
        RECT 439.950 277.950 442.050 280.050 ;
        RECT 452.400 277.050 453.450 283.950 ;
        RECT 467.100 282.600 468.300 302.400 ;
        RECT 473.400 297.450 474.450 307.950 ;
        RECT 470.400 296.400 474.450 297.450 ;
        RECT 470.400 294.600 471.450 296.400 ;
        RECT 470.400 292.350 471.600 294.600 ;
        RECT 469.950 289.950 472.050 292.050 ;
        RECT 466.950 280.500 469.050 282.600 ;
        RECT 436.950 274.950 439.050 277.050 ;
        RECT 451.950 274.950 454.050 277.050 ;
        RECT 427.950 271.950 430.050 274.050 ;
        RECT 428.400 265.050 429.450 271.950 ;
        RECT 439.950 265.950 442.050 268.050 ;
        RECT 451.950 265.950 454.050 268.050 ;
        RECT 463.950 265.950 466.050 268.050 ;
        RECT 424.950 262.950 427.050 265.050 ;
        RECT 376.950 257.100 379.050 259.200 ;
        RECT 379.950 257.100 382.050 259.200 ;
        RECT 382.950 257.100 385.050 259.200 ;
        RECT 391.950 257.100 394.050 259.200 ;
        RECT 394.950 257.100 397.050 259.200 ;
        RECT 397.950 257.100 400.050 259.200 ;
        RECT 377.400 256.050 378.600 256.800 ;
        RECT 383.400 256.050 384.600 256.800 ;
        RECT 376.950 253.950 379.050 256.050 ;
        RECT 382.950 253.950 385.050 256.050 ;
        RECT 392.400 254.400 393.600 256.800 ;
        RECT 392.400 232.050 393.450 254.400 ;
        RECT 394.950 253.950 397.050 256.050 ;
        RECT 398.400 254.400 399.600 256.800 ;
        RECT 376.950 229.950 379.050 232.050 ;
        RECT 391.950 229.950 394.050 232.050 ;
        RECT 370.950 217.950 373.050 220.050 ;
        RECT 372.000 216.600 376.050 217.050 ;
        RECT 371.400 214.950 376.050 216.600 ;
        RECT 371.400 214.350 372.600 214.950 ;
        RECT 370.950 211.950 373.050 214.050 ;
        RECT 373.950 208.950 376.050 211.050 ;
        RECT 349.950 202.500 352.050 204.600 ;
        RECT 364.950 202.500 367.050 204.600 ;
        RECT 355.950 199.950 358.050 202.050 ;
        RECT 325.950 193.950 328.050 196.050 ;
        RECT 343.950 193.950 346.050 196.050 ;
        RECT 352.950 193.950 355.050 196.050 ;
        RECT 326.400 183.600 327.450 193.950 ;
        RECT 331.950 190.950 334.050 193.050 ;
        RECT 332.400 183.600 333.450 190.950 ;
        RECT 340.950 188.400 343.050 190.500 ;
        RECT 314.400 182.400 318.450 183.450 ;
        RECT 280.950 175.950 283.050 178.050 ;
        RECT 286.950 175.950 289.050 178.050 ;
        RECT 289.950 175.950 292.050 178.050 ;
        RECT 292.950 175.950 295.050 178.050 ;
        RECT 281.400 169.050 282.450 175.950 ;
        RECT 286.950 169.950 289.050 172.050 ;
        RECT 280.950 166.950 283.050 169.050 ;
        RECT 280.950 146.400 283.050 148.500 ;
        RECT 287.400 148.050 288.450 169.950 ;
        RECT 259.950 136.950 262.050 139.050 ;
        RECT 262.950 138.000 265.050 142.050 ;
        RECT 268.950 138.000 271.050 142.050 ;
        RECT 274.950 139.950 277.050 142.050 ;
        RECT 263.400 136.350 264.600 138.000 ;
        RECT 269.400 136.350 270.600 138.000 ;
        RECT 277.950 137.100 280.050 139.200 ;
        RECT 278.400 136.350 279.600 137.100 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 259.950 130.950 262.050 133.050 ;
        RECT 266.400 132.000 267.600 133.650 ;
        RECT 256.950 124.950 259.050 127.050 ;
        RECT 250.950 121.950 253.050 124.050 ;
        RECT 256.950 121.800 259.050 123.900 ;
        RECT 238.950 115.950 241.050 118.050 ;
        RECT 244.950 115.950 247.050 118.050 ;
        RECT 235.950 109.950 238.050 112.050 ;
        RECT 236.400 103.050 237.450 109.950 ;
        RECT 239.400 106.050 240.450 115.950 ;
        RECT 247.950 110.400 250.050 112.500 ;
        RECT 238.950 103.950 241.050 106.050 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 241.950 100.950 244.050 103.050 ;
        RECT 242.400 99.900 243.600 100.650 ;
        RECT 241.950 97.800 244.050 99.900 ;
        RECT 248.100 90.600 249.300 110.400 ;
        RECT 250.950 100.950 253.050 103.050 ;
        RECT 251.400 98.400 252.600 100.650 ;
        RECT 257.400 99.450 258.450 121.800 ;
        RECT 260.400 105.450 261.450 130.950 ;
        RECT 265.950 127.950 268.050 132.000 ;
        RECT 272.400 131.400 273.600 133.650 ;
        RECT 272.400 118.050 273.450 131.400 ;
        RECT 274.950 130.950 277.050 133.050 ;
        RECT 271.950 115.950 274.050 118.050 ;
        RECT 272.400 112.050 273.450 115.950 ;
        RECT 271.950 109.950 274.050 112.050 ;
        RECT 263.400 105.450 264.600 105.600 ;
        RECT 260.400 104.400 264.600 105.450 ;
        RECT 263.400 103.350 264.600 104.400 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 269.400 99.900 270.600 100.650 ;
        RECT 254.400 98.400 258.450 99.450 ;
        RECT 251.400 94.050 252.450 98.400 ;
        RECT 250.950 91.950 253.050 94.050 ;
        RECT 247.950 88.500 250.050 90.600 ;
        RECT 235.950 76.950 238.050 79.050 ;
        RECT 220.950 73.950 223.050 76.050 ;
        RECT 232.950 73.950 235.050 76.050 ;
        RECT 193.950 69.300 196.050 71.400 ;
        RECT 193.950 65.700 195.150 69.300 ;
        RECT 193.950 63.600 196.050 65.700 ;
        RECT 187.950 46.950 190.050 49.050 ;
        RECT 193.950 48.600 195.150 63.600 ;
        RECT 202.950 61.950 205.050 64.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 197.400 54.900 198.600 55.650 ;
        RECT 203.400 55.050 204.450 61.950 ;
        RECT 205.950 58.950 208.050 61.050 ;
        RECT 214.950 58.950 217.050 61.050 ;
        RECT 221.400 60.600 222.450 73.950 ;
        RECT 229.950 69.300 232.050 71.400 ;
        RECT 230.850 65.700 232.050 69.300 ;
        RECT 229.950 63.600 232.050 65.700 ;
        RECT 196.950 54.450 199.050 54.900 ;
        RECT 196.950 53.400 201.450 54.450 ;
        RECT 196.950 52.800 199.050 53.400 ;
        RECT 200.400 49.050 201.450 53.400 ;
        RECT 202.950 52.950 205.050 55.050 ;
        RECT 193.950 46.500 196.050 48.600 ;
        RECT 199.950 46.950 202.050 49.050 ;
        RECT 193.950 32.400 196.050 34.500 ;
        RECT 184.950 28.950 187.050 31.050 ;
        RECT 178.950 22.950 181.050 25.050 ;
        RECT 179.400 21.900 180.600 22.650 ;
        RECT 178.950 19.800 181.050 21.900 ;
        RECT 185.400 13.050 186.450 28.950 ;
        RECT 193.950 17.400 195.150 32.400 ;
        RECT 196.950 26.100 199.050 28.200 ;
        RECT 202.950 26.100 205.050 28.200 ;
        RECT 197.400 25.350 198.600 26.100 ;
        RECT 196.950 22.950 199.050 25.050 ;
        RECT 193.950 15.300 196.050 17.400 ;
        RECT 203.400 16.050 204.450 26.100 ;
        RECT 206.400 19.050 207.450 58.950 ;
        RECT 215.400 58.200 216.600 58.950 ;
        RECT 221.400 58.200 222.600 60.600 ;
        RECT 211.950 55.800 214.050 57.900 ;
        RECT 214.950 55.800 217.050 57.900 ;
        RECT 217.950 55.800 220.050 57.900 ;
        RECT 220.950 55.800 223.050 57.900 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 212.400 54.750 213.600 55.500 ;
        RECT 218.400 54.750 219.600 55.500 ;
        RECT 227.400 54.900 228.600 55.650 ;
        RECT 211.950 52.650 214.050 54.750 ;
        RECT 217.950 52.650 220.050 54.750 ;
        RECT 226.950 52.800 229.050 54.900 ;
        RECT 211.950 46.950 214.050 49.050 ;
        RECT 230.850 48.600 232.050 63.600 ;
        RECT 236.400 58.050 237.450 76.950 ;
        RECT 254.400 76.050 255.450 98.400 ;
        RECT 268.950 97.800 271.050 99.900 ;
        RECT 275.400 94.050 276.450 130.950 ;
        RECT 281.700 126.600 282.900 146.400 ;
        RECT 286.950 145.950 289.050 148.050 ;
        RECT 286.950 138.000 289.050 142.050 ;
        RECT 290.400 139.050 291.450 175.950 ;
        RECT 296.400 166.050 297.450 181.950 ;
        RECT 305.400 181.350 306.600 182.100 ;
        RECT 311.400 181.350 312.600 182.100 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 304.950 178.950 307.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 310.950 178.950 313.050 181.050 ;
        RECT 302.400 177.900 303.600 178.650 ;
        RECT 301.950 175.800 304.050 177.900 ;
        RECT 308.400 176.400 309.600 178.650 ;
        RECT 295.950 163.950 298.050 166.050 ;
        RECT 301.950 147.300 304.050 149.400 ;
        RECT 301.950 143.700 303.150 147.300 ;
        RECT 308.400 145.050 309.450 176.400 ;
        RECT 313.950 175.950 316.050 178.050 ;
        RECT 310.950 169.950 313.050 175.050 ;
        RECT 314.400 172.050 315.450 175.950 ;
        RECT 317.400 175.050 318.450 182.400 ;
        RECT 326.400 181.350 327.600 183.600 ;
        RECT 332.400 181.350 333.600 183.600 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 325.950 178.950 328.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 337.950 178.950 340.050 181.050 ;
        RECT 316.950 172.950 319.050 175.050 ;
        RECT 319.950 172.950 322.050 178.050 ;
        RECT 323.400 176.400 324.600 178.650 ;
        RECT 329.400 177.900 330.600 178.650 ;
        RECT 313.950 169.950 316.050 172.050 ;
        RECT 319.950 169.800 322.050 171.900 ;
        RECT 320.400 163.050 321.450 169.800 ;
        RECT 323.400 166.050 324.450 176.400 ;
        RECT 328.950 175.800 331.050 177.900 ;
        RECT 338.400 177.450 339.600 178.650 ;
        RECT 335.400 176.400 339.600 177.450 ;
        RECT 335.400 166.050 336.450 176.400 ;
        RECT 341.700 168.600 342.900 188.400 ;
        RECT 353.400 184.200 354.450 193.950 ;
        RECT 352.950 182.100 355.050 184.200 ;
        RECT 346.950 178.950 349.050 181.050 ;
        RECT 347.400 177.000 348.600 178.650 ;
        RECT 346.950 172.950 349.050 177.000 ;
        RECT 340.950 166.500 343.050 168.600 ;
        RECT 322.950 163.950 325.050 166.050 ;
        RECT 334.950 163.950 337.050 166.050 ;
        RECT 319.950 160.950 322.050 163.050 ;
        RECT 334.950 160.800 337.050 162.900 ;
        RECT 292.950 139.950 295.050 142.050 ;
        RECT 301.950 141.600 304.050 143.700 ;
        RECT 307.950 142.950 310.050 145.050 ;
        RECT 287.400 136.350 288.600 138.000 ;
        RECT 289.950 136.950 292.050 139.050 ;
        RECT 286.950 133.950 289.050 136.050 ;
        RECT 289.950 130.950 292.050 133.050 ;
        RECT 280.950 124.500 283.050 126.600 ;
        RECT 290.400 118.050 291.450 130.950 ;
        RECT 293.400 130.050 294.450 139.950 ;
        RECT 292.950 127.950 295.050 130.050 ;
        RECT 301.950 126.600 303.150 141.600 ;
        RECT 310.950 136.950 313.050 139.050 ;
        RECT 316.950 136.950 319.050 139.050 ;
        RECT 322.950 136.950 325.050 139.050 ;
        RECT 328.950 136.950 331.050 139.050 ;
        RECT 335.400 138.600 336.450 160.800 ;
        RECT 340.950 154.950 343.050 157.050 ;
        RECT 341.400 138.600 342.450 154.950 ;
        RECT 346.950 151.950 349.050 154.050 ;
        RECT 347.400 139.050 348.450 151.950 ;
        RECT 353.400 148.050 354.450 182.100 ;
        RECT 352.950 145.950 355.050 148.050 ;
        RECT 349.950 142.950 352.050 145.050 ;
        RECT 350.400 139.050 351.450 142.950 ;
        RECT 356.400 141.450 357.450 199.950 ;
        RECT 374.400 199.050 375.450 208.950 ;
        RECT 373.950 196.950 376.050 199.050 ;
        RECT 361.950 188.400 364.050 190.500 ;
        RECT 377.400 190.050 378.450 229.950 ;
        RECT 385.950 225.300 388.050 227.400 ;
        RECT 392.400 226.050 393.450 229.950 ;
        RECT 385.950 221.700 387.150 225.300 ;
        RECT 391.950 223.950 394.050 226.050 ;
        RECT 379.950 217.950 382.050 220.050 ;
        RECT 385.950 219.600 388.050 221.700 ;
        RECT 380.400 202.050 381.450 217.950 ;
        RECT 385.950 204.600 387.150 219.600 ;
        RECT 388.950 211.950 391.050 214.050 ;
        RECT 389.400 210.900 390.600 211.650 ;
        RECT 388.950 208.800 391.050 210.900 ;
        RECT 395.400 210.450 396.450 253.950 ;
        RECT 398.400 244.050 399.450 254.400 ;
        RECT 404.400 247.050 405.450 260.400 ;
        RECT 413.400 259.500 414.600 261.600 ;
        RECT 418.950 259.950 421.050 262.050 ;
        RECT 427.950 261.000 430.050 265.050 ;
        RECT 428.400 259.350 429.600 261.000 ;
        RECT 409.950 257.100 412.050 259.200 ;
        RECT 412.950 257.100 415.050 259.200 ;
        RECT 415.950 257.100 418.050 259.200 ;
        RECT 427.950 256.950 430.050 259.050 ;
        RECT 433.950 256.950 436.050 259.050 ;
        RECT 410.400 254.400 411.600 256.800 ;
        RECT 416.400 256.050 417.600 256.800 ;
        RECT 403.950 244.950 406.050 247.050 ;
        RECT 397.950 241.950 400.050 244.050 ;
        RECT 406.950 220.950 409.050 223.050 ;
        RECT 407.400 216.600 408.450 220.950 ;
        RECT 410.400 220.050 411.450 254.400 ;
        RECT 415.950 253.950 418.050 256.050 ;
        RECT 434.400 254.400 435.600 256.650 ;
        RECT 434.400 250.050 435.450 254.400 ;
        RECT 433.950 247.950 436.050 250.050 ;
        RECT 434.400 244.050 435.450 247.950 ;
        RECT 440.400 244.050 441.450 265.950 ;
        RECT 445.950 260.100 448.050 262.200 ;
        RECT 452.400 261.600 453.450 265.950 ;
        RECT 446.400 259.350 447.600 260.100 ;
        RECT 452.400 259.350 453.600 261.600 ;
        RECT 460.950 260.100 463.050 262.200 ;
        RECT 445.950 256.950 448.050 259.050 ;
        RECT 448.950 256.950 451.050 259.050 ;
        RECT 451.950 256.950 454.050 259.050 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 449.400 255.900 450.600 256.650 ;
        RECT 455.400 255.900 456.600 256.650 ;
        RECT 448.950 253.800 451.050 255.900 ;
        RECT 454.950 253.800 457.050 255.900 ;
        RECT 461.400 250.050 462.450 260.100 ;
        RECT 460.950 247.950 463.050 250.050 ;
        RECT 448.950 244.950 451.050 247.050 ;
        RECT 433.950 241.950 436.050 244.050 ;
        RECT 439.950 241.950 442.050 244.050 ;
        RECT 445.950 229.950 448.050 232.050 ;
        RECT 418.950 223.950 421.050 226.050 ;
        RECT 439.950 225.300 442.050 227.400 ;
        RECT 409.950 217.950 412.050 220.050 ;
        RECT 419.400 217.050 420.450 223.950 ;
        RECT 424.950 220.950 427.050 223.050 ;
        RECT 440.850 221.700 442.050 225.300 ;
        RECT 407.400 214.350 408.600 216.600 ;
        RECT 418.950 214.950 421.050 217.050 ;
        RECT 425.400 216.600 426.450 220.950 ;
        RECT 439.950 219.600 442.050 221.700 ;
        RECT 419.400 214.200 420.600 214.950 ;
        RECT 425.400 214.200 426.600 216.600 ;
        RECT 403.950 211.950 406.050 214.050 ;
        RECT 406.950 211.950 409.050 214.050 ;
        RECT 409.950 211.950 412.050 214.050 ;
        RECT 418.950 211.800 421.050 213.900 ;
        RECT 421.950 211.800 424.050 213.900 ;
        RECT 424.950 211.800 427.050 213.900 ;
        RECT 427.950 211.800 430.050 213.900 ;
        RECT 436.950 211.950 439.050 214.050 ;
        RECT 404.400 210.900 405.600 211.650 ;
        RECT 410.400 210.900 411.600 211.650 ;
        RECT 397.950 210.450 400.050 210.900 ;
        RECT 395.400 209.400 400.050 210.450 ;
        RECT 397.950 208.800 400.050 209.400 ;
        RECT 403.950 208.800 406.050 210.900 ;
        RECT 409.950 208.800 412.050 210.900 ;
        RECT 422.400 209.400 423.600 211.500 ;
        RECT 428.400 210.750 429.600 211.500 ;
        RECT 385.950 202.500 388.050 204.600 ;
        RECT 379.950 199.950 382.050 202.050 ;
        RECT 382.950 196.950 385.050 199.050 ;
        RECT 361.950 173.400 363.150 188.400 ;
        RECT 370.950 187.950 373.050 190.050 ;
        RECT 376.950 187.950 379.050 190.050 ;
        RECT 364.950 182.100 367.050 184.200 ;
        RECT 365.400 181.350 366.600 182.100 ;
        RECT 364.950 178.950 367.050 181.050 ;
        RECT 361.950 171.300 364.050 173.400 ;
        RECT 361.950 167.700 363.150 171.300 ;
        RECT 361.950 165.600 364.050 167.700 ;
        RECT 361.950 160.950 364.050 163.050 ;
        RECT 362.400 148.050 363.450 160.950 ;
        RECT 358.800 145.950 360.900 148.050 ;
        RECT 361.950 145.950 364.050 148.050 ;
        RECT 353.400 140.400 357.450 141.450 ;
        RECT 304.950 133.950 307.050 136.050 ;
        RECT 305.400 132.900 306.600 133.650 ;
        RECT 311.400 132.900 312.450 136.950 ;
        RECT 317.400 136.200 318.600 136.950 ;
        RECT 323.400 136.200 324.600 136.950 ;
        RECT 316.950 133.800 319.050 135.900 ;
        RECT 319.950 133.800 322.050 135.900 ;
        RECT 322.950 133.800 325.050 135.900 ;
        RECT 304.950 130.800 307.050 132.900 ;
        RECT 310.950 130.800 313.050 132.900 ;
        RECT 320.400 131.400 321.600 133.500 ;
        RECT 311.400 127.050 312.450 130.800 ;
        RECT 301.950 124.500 304.050 126.600 ;
        RECT 310.950 124.950 313.050 127.050 ;
        RECT 320.400 124.050 321.450 131.400 ;
        RECT 307.950 123.450 310.050 124.050 ;
        RECT 313.950 123.450 316.050 124.050 ;
        RECT 307.950 122.400 316.050 123.450 ;
        RECT 307.950 121.950 310.050 122.400 ;
        RECT 313.950 121.950 316.050 122.400 ;
        RECT 319.950 121.950 322.050 124.050 ;
        RECT 292.950 118.950 295.050 121.050 ;
        RECT 283.950 115.950 286.050 118.050 ;
        RECT 289.950 115.950 292.050 118.050 ;
        RECT 284.400 105.600 285.450 115.950 ;
        RECT 293.400 109.050 294.450 118.950 ;
        RECT 307.950 115.950 310.050 118.050 ;
        RECT 298.950 110.400 301.050 112.500 ;
        RECT 292.950 106.950 295.050 109.050 ;
        RECT 284.400 103.500 285.600 105.600 ;
        RECT 295.950 104.100 298.050 106.200 ;
        RECT 296.400 103.350 297.600 104.100 ;
        RECT 280.950 101.100 283.050 103.200 ;
        RECT 283.950 101.100 286.050 103.200 ;
        RECT 286.950 101.100 289.050 103.200 ;
        RECT 295.950 100.950 298.050 103.050 ;
        RECT 281.400 100.050 282.600 100.800 ;
        RECT 287.400 100.050 288.600 100.800 ;
        RECT 280.950 97.950 283.050 100.050 ;
        RECT 286.950 97.950 289.050 100.050 ;
        RECT 256.950 91.950 259.050 94.050 ;
        RECT 274.950 91.950 277.050 94.050 ;
        RECT 253.950 73.950 256.050 76.050 ;
        RECT 238.950 70.950 241.050 73.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 212.400 27.600 213.450 46.950 ;
        RECT 229.950 46.500 232.050 48.600 ;
        RECT 239.400 37.050 240.450 70.950 ;
        RECT 250.950 68.400 253.050 70.500 ;
        RECT 244.950 64.950 247.050 67.050 ;
        RECT 245.400 60.600 246.450 64.950 ;
        RECT 245.400 58.350 246.600 60.600 ;
        RECT 244.950 55.950 247.050 58.050 ;
        RECT 251.100 48.600 252.300 68.400 ;
        RECT 257.400 63.450 258.450 91.950 ;
        RECT 262.950 85.950 265.050 88.050 ;
        RECT 263.400 82.050 264.450 85.950 ;
        RECT 262.950 79.950 265.050 82.050 ;
        RECT 259.950 73.950 262.050 76.050 ;
        RECT 260.400 67.050 261.450 73.950 ;
        RECT 259.950 64.950 262.050 67.050 ;
        RECT 254.400 62.400 258.450 63.450 ;
        RECT 254.400 60.600 255.450 62.400 ;
        RECT 259.950 61.800 262.050 63.900 ;
        RECT 254.400 58.350 255.600 60.600 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 260.400 54.900 261.450 61.800 ;
        RECT 263.400 61.050 264.450 79.950 ;
        RECT 277.950 73.950 280.050 76.050 ;
        RECT 271.950 69.450 274.050 70.050 ;
        RECT 266.400 68.400 274.050 69.450 ;
        RECT 266.400 64.050 267.450 68.400 ;
        RECT 271.950 67.950 274.050 68.400 ;
        RECT 268.950 64.950 271.050 67.050 ;
        RECT 265.950 61.950 268.050 64.050 ;
        RECT 262.950 58.950 265.050 61.050 ;
        RECT 269.400 60.600 270.450 64.950 ;
        RECT 269.400 58.350 270.600 60.600 ;
        RECT 274.950 59.100 277.050 61.200 ;
        RECT 278.400 61.050 279.450 73.950 ;
        RECT 275.400 58.350 276.600 59.100 ;
        RECT 277.950 58.950 280.050 61.050 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 274.950 55.950 277.050 58.050 ;
        RECT 266.400 54.900 267.600 55.650 ;
        RECT 259.950 52.800 262.050 54.900 ;
        RECT 265.950 52.800 268.050 54.900 ;
        RECT 272.400 53.400 273.600 55.650 ;
        RECT 272.400 49.050 273.450 53.400 ;
        RECT 277.950 52.950 280.050 55.050 ;
        RECT 278.400 49.050 279.450 52.950 ;
        RECT 281.400 52.050 282.450 97.950 ;
        RECT 287.400 85.050 288.450 97.950 ;
        RECT 299.850 95.400 301.050 110.400 ;
        RECT 308.400 99.900 309.450 115.950 ;
        RECT 319.950 110.400 322.050 112.500 ;
        RECT 329.400 112.050 330.450 136.950 ;
        RECT 335.400 136.200 336.600 138.600 ;
        RECT 341.400 136.200 342.600 138.600 ;
        RECT 346.950 136.950 349.050 139.050 ;
        RECT 349.950 136.950 352.050 139.050 ;
        RECT 347.400 136.200 348.600 136.950 ;
        RECT 334.950 133.800 337.050 135.900 ;
        RECT 337.950 133.800 340.050 135.900 ;
        RECT 340.950 133.800 343.050 135.900 ;
        RECT 343.950 133.800 346.050 135.900 ;
        RECT 346.950 133.800 349.050 135.900 ;
        RECT 338.400 131.400 339.600 133.500 ;
        RECT 344.400 131.400 345.600 133.500 ;
        RECT 353.400 133.050 354.450 140.400 ;
        RECT 359.400 138.450 360.450 145.950 ;
        RECT 356.400 137.400 360.450 138.450 ;
        RECT 362.400 138.600 363.450 145.950 ;
        RECT 371.400 139.050 372.450 187.950 ;
        RECT 376.950 182.100 379.050 184.200 ;
        RECT 383.400 183.600 384.450 196.950 ;
        RECT 394.950 187.950 397.050 190.050 ;
        RECT 377.400 181.350 378.600 182.100 ;
        RECT 383.400 181.350 384.600 183.600 ;
        RECT 391.950 182.100 394.050 184.200 ;
        RECT 376.950 178.950 379.050 181.050 ;
        RECT 379.950 178.950 382.050 181.050 ;
        RECT 382.950 178.950 385.050 181.050 ;
        RECT 385.950 178.950 388.050 181.050 ;
        RECT 380.400 177.900 381.600 178.650 ;
        RECT 379.950 175.800 382.050 177.900 ;
        RECT 386.400 177.000 387.600 178.650 ;
        RECT 380.400 174.450 381.450 175.800 ;
        RECT 380.400 173.400 384.450 174.450 ;
        RECT 313.950 100.950 316.050 103.050 ;
        RECT 314.400 99.900 315.600 100.650 ;
        RECT 307.950 97.800 310.050 99.900 ;
        RECT 313.950 97.800 316.050 99.900 ;
        RECT 298.950 93.300 301.050 95.400 ;
        RECT 299.850 89.700 301.050 93.300 ;
        RECT 320.100 90.600 321.300 110.400 ;
        RECT 328.950 109.950 331.050 112.050 ;
        RECT 338.400 109.050 339.450 131.400 ;
        RECT 344.400 127.050 345.450 131.400 ;
        RECT 352.950 130.950 355.050 133.050 ;
        RECT 352.950 127.800 355.050 129.900 ;
        RECT 343.950 124.950 346.050 127.050 ;
        RECT 340.950 115.950 343.050 118.050 ;
        RECT 337.950 106.950 340.050 109.050 ;
        RECT 341.400 105.600 342.450 115.950 ;
        RECT 349.950 112.950 352.050 115.050 ;
        RECT 335.400 105.450 336.600 105.600 ;
        RECT 329.400 104.400 336.600 105.450 ;
        RECT 322.950 100.950 325.050 103.050 ;
        RECT 323.400 98.400 324.600 100.650 ;
        RECT 323.400 94.050 324.450 98.400 ;
        RECT 322.950 91.950 325.050 94.050 ;
        RECT 298.950 87.600 301.050 89.700 ;
        RECT 319.950 88.500 322.050 90.600 ;
        RECT 329.400 88.050 330.450 104.400 ;
        RECT 335.400 103.350 336.600 104.400 ;
        RECT 341.400 103.350 342.600 105.600 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 337.950 100.950 340.050 103.050 ;
        RECT 340.950 100.950 343.050 103.050 ;
        RECT 343.950 100.950 346.050 103.050 ;
        RECT 338.400 99.900 339.600 100.650 ;
        RECT 344.400 100.050 345.600 100.650 ;
        RECT 337.950 97.800 340.050 99.900 ;
        RECT 344.400 98.400 349.050 100.050 ;
        RECT 345.000 97.950 349.050 98.400 ;
        RECT 337.950 91.950 340.050 94.050 ;
        RECT 328.950 85.950 331.050 88.050 ;
        RECT 286.950 82.950 289.050 85.050 ;
        RECT 338.400 70.050 339.450 91.950 ;
        RECT 350.400 91.050 351.450 112.950 ;
        RECT 353.400 97.050 354.450 127.800 ;
        RECT 356.400 124.050 357.450 137.400 ;
        RECT 362.400 136.350 363.600 138.600 ;
        RECT 370.950 136.950 373.050 139.050 ;
        RECT 373.950 136.950 376.050 139.050 ;
        RECT 379.800 137.100 381.900 139.200 ;
        RECT 383.400 139.050 384.450 173.400 ;
        RECT 385.950 172.950 388.050 177.000 ;
        RECT 392.400 172.050 393.450 182.100 ;
        RECT 391.950 169.950 394.050 172.050 ;
        RECT 395.400 169.050 396.450 187.950 ;
        RECT 398.400 184.050 399.450 208.800 ;
        RECT 404.400 205.050 405.450 208.800 ;
        RECT 403.950 202.950 406.050 205.050 ;
        RECT 410.400 184.200 411.450 208.800 ;
        RECT 422.400 202.050 423.450 209.400 ;
        RECT 427.950 208.650 430.050 210.750 ;
        RECT 437.400 210.450 438.600 211.650 ;
        RECT 434.400 209.400 438.600 210.450 ;
        RECT 434.400 205.050 435.450 209.400 ;
        RECT 433.950 202.950 436.050 205.050 ;
        RECT 440.850 204.600 442.050 219.600 ;
        RECT 439.950 202.500 442.050 204.600 ;
        RECT 421.950 199.950 424.050 202.050 ;
        RECT 430.950 199.950 433.050 202.050 ;
        RECT 422.400 196.050 423.450 199.950 ;
        RECT 421.950 193.950 424.050 196.050 ;
        RECT 397.950 181.950 400.050 184.050 ;
        RECT 403.950 182.100 406.050 184.200 ;
        RECT 409.950 182.100 412.050 184.200 ;
        RECT 418.950 182.100 421.050 184.200 ;
        RECT 424.950 182.100 427.050 184.200 ;
        RECT 404.400 181.350 405.600 182.100 ;
        RECT 410.400 181.350 411.600 182.100 ;
        RECT 419.400 181.350 420.600 182.100 ;
        RECT 425.400 181.350 426.600 182.100 ;
        RECT 400.950 178.950 403.050 181.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 406.950 178.950 409.050 181.050 ;
        RECT 409.950 178.950 412.050 181.050 ;
        RECT 418.950 178.950 421.050 181.050 ;
        RECT 421.950 178.950 424.050 181.050 ;
        RECT 424.950 178.950 427.050 181.050 ;
        RECT 401.400 177.900 402.600 178.650 ;
        RECT 400.950 175.800 403.050 177.900 ;
        RECT 407.400 176.400 408.600 178.650 ;
        RECT 422.400 176.400 423.600 178.650 ;
        RECT 403.950 169.950 406.050 172.050 ;
        RECT 394.950 166.950 397.050 169.050 ;
        RECT 400.950 163.950 403.050 166.050 ;
        RECT 388.950 157.950 391.050 160.050 ;
        RECT 361.950 133.950 364.050 136.050 ;
        RECT 367.950 133.950 370.050 136.050 ;
        RECT 368.400 132.900 369.600 133.650 ;
        RECT 367.950 130.800 370.050 132.900 ;
        RECT 370.950 130.950 373.050 133.050 ;
        RECT 355.950 121.950 358.050 124.050 ;
        RECT 371.400 121.050 372.450 130.950 ;
        RECT 374.400 129.450 375.450 136.950 ;
        RECT 380.400 136.350 381.600 137.100 ;
        RECT 382.950 136.950 385.050 139.050 ;
        RECT 389.400 138.450 390.450 157.950 ;
        RECT 394.950 146.400 397.050 148.500 ;
        RECT 401.400 148.050 402.450 163.950 ;
        RECT 392.400 138.450 393.600 138.600 ;
        RECT 389.400 137.400 393.600 138.450 ;
        RECT 392.400 136.350 393.600 137.400 ;
        RECT 379.950 133.950 382.050 136.050 ;
        RECT 385.950 133.950 388.050 136.050 ;
        RECT 391.950 133.950 394.050 136.050 ;
        RECT 382.950 130.950 385.050 133.050 ;
        RECT 386.400 131.400 387.600 133.650 ;
        RECT 374.400 128.400 378.450 129.450 ;
        RECT 373.950 124.950 376.050 127.050 ;
        RECT 370.950 118.950 373.050 121.050 ;
        RECT 355.950 103.950 358.050 109.050 ;
        RECT 361.950 104.100 364.050 106.200 ;
        RECT 367.950 104.100 370.050 106.200 ;
        RECT 362.400 103.350 363.600 104.100 ;
        RECT 368.400 103.350 369.600 104.100 ;
        RECT 358.950 100.950 361.050 103.050 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 359.400 98.400 360.600 100.650 ;
        RECT 365.400 99.000 366.600 100.650 ;
        RECT 374.400 100.050 375.450 124.950 ;
        RECT 377.400 112.050 378.450 128.400 ;
        RECT 383.400 118.050 384.450 130.950 ;
        RECT 386.400 121.050 387.450 131.400 ;
        RECT 388.950 130.950 391.050 133.050 ;
        RECT 389.400 127.050 390.450 130.950 ;
        RECT 388.950 124.950 391.050 127.050 ;
        RECT 395.700 126.600 396.900 146.400 ;
        RECT 400.950 145.950 403.050 148.050 ;
        RECT 401.400 139.200 402.450 145.950 ;
        RECT 404.400 141.450 405.450 169.950 ;
        RECT 407.400 145.050 408.450 176.400 ;
        RECT 422.400 175.050 423.450 176.400 ;
        RECT 421.950 172.950 424.050 175.050 ;
        RECT 427.950 174.450 430.050 178.050 ;
        RECT 425.400 174.000 430.050 174.450 ;
        RECT 425.400 173.400 429.450 174.000 ;
        RECT 422.400 154.050 423.450 172.950 ;
        RECT 421.950 151.950 424.050 154.050 ;
        RECT 415.950 147.300 418.050 149.400 ;
        RECT 406.950 142.950 409.050 145.050 ;
        RECT 415.950 143.700 417.150 147.300 ;
        RECT 425.400 145.050 426.450 173.400 ;
        RECT 431.400 171.450 432.450 199.950 ;
        RECT 439.950 183.000 442.050 187.050 ;
        RECT 446.400 183.600 447.450 229.950 ;
        RECT 449.400 187.050 450.450 244.950 ;
        RECT 464.400 231.450 465.450 265.950 ;
        RECT 476.400 265.050 477.450 364.950 ;
        RECT 481.950 364.800 484.050 366.900 ;
        RECT 487.950 364.800 490.050 366.900 ;
        RECT 500.400 365.400 501.600 367.500 ;
        RECT 512.400 366.900 513.600 367.650 ;
        RECT 488.400 352.050 489.450 364.800 ;
        RECT 500.400 358.050 501.450 365.400 ;
        RECT 511.950 364.800 514.050 366.900 ;
        RECT 515.850 360.600 517.050 375.600 ;
        RECT 530.400 372.600 531.450 376.950 ;
        RECT 530.400 370.350 531.600 372.600 ;
        RECT 529.950 367.950 532.050 370.050 ;
        RECT 536.100 360.600 537.300 380.400 ;
        RECT 542.400 373.200 543.450 385.950 ;
        RECT 550.950 380.400 553.050 382.500 ;
        RECT 539.400 372.450 540.600 372.600 ;
        RECT 541.950 372.450 544.050 373.200 ;
        RECT 539.400 371.400 544.050 372.450 ;
        RECT 539.400 370.350 540.600 371.400 ;
        RECT 541.950 371.100 544.050 371.400 ;
        RECT 547.950 371.100 550.050 373.200 ;
        RECT 548.400 370.350 549.600 371.100 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 547.950 367.950 550.050 370.050 ;
        RECT 551.700 360.600 552.900 380.400 ;
        RECT 556.950 371.100 559.050 373.200 ;
        RECT 562.950 371.100 565.050 373.200 ;
        RECT 557.400 370.350 558.600 371.100 ;
        RECT 556.950 367.950 559.050 370.050 ;
        RECT 563.400 361.050 564.450 371.100 ;
        RECT 514.950 358.500 517.050 360.600 ;
        RECT 535.950 358.500 538.050 360.600 ;
        RECT 550.950 358.500 553.050 360.600 ;
        RECT 562.950 358.950 565.050 361.050 ;
        RECT 499.950 355.950 502.050 358.050 ;
        RECT 487.950 349.950 490.050 352.050 ;
        RECT 499.950 349.950 502.050 352.050 ;
        RECT 490.950 343.950 493.050 346.050 ;
        RECT 491.400 340.200 492.450 343.950 ;
        RECT 500.400 340.200 501.450 349.950 ;
        RECT 566.400 349.050 567.450 409.950 ;
        RECT 577.950 406.950 580.050 411.000 ;
        RECT 592.950 409.800 595.050 411.900 ;
        RECT 599.400 406.050 600.450 416.400 ;
        RECT 601.950 415.950 604.050 418.050 ;
        RECT 605.400 417.600 606.450 421.950 ;
        RECT 611.400 417.600 612.450 430.950 ;
        RECT 620.400 430.050 621.450 436.950 ;
        RECT 619.950 427.950 622.050 430.050 ;
        RECT 616.950 421.950 619.050 424.050 ;
        RECT 605.400 415.350 606.600 417.600 ;
        RECT 611.400 415.350 612.600 417.600 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 601.950 409.950 604.050 412.050 ;
        RECT 608.400 410.400 609.600 412.650 ;
        RECT 598.950 403.950 601.050 406.050 ;
        RECT 571.950 381.300 574.050 383.400 ;
        RECT 571.950 377.700 573.150 381.300 ;
        RECT 599.400 379.050 600.450 403.950 ;
        RECT 602.400 397.050 603.450 409.950 ;
        RECT 604.950 406.950 607.050 409.050 ;
        RECT 601.950 394.950 604.050 397.050 ;
        RECT 571.950 375.600 574.050 377.700 ;
        RECT 598.950 376.950 601.050 379.050 ;
        RECT 571.950 360.600 573.150 375.600 ;
        RECT 589.950 371.100 592.050 373.200 ;
        RECT 605.400 373.050 606.450 406.950 ;
        RECT 608.400 376.050 609.450 410.400 ;
        RECT 617.400 382.050 618.450 421.950 ;
        RECT 623.400 421.200 624.450 443.400 ;
        RECT 628.950 442.650 631.050 444.750 ;
        RECT 638.400 442.050 639.450 451.950 ;
        RECT 659.400 451.200 660.450 454.950 ;
        RECT 643.950 449.100 646.050 451.200 ;
        RECT 658.950 449.100 661.050 451.200 ;
        RECT 664.950 449.100 667.050 451.200 ;
        RECT 644.400 448.350 645.600 449.100 ;
        RECT 659.400 448.350 660.600 449.100 ;
        RECT 665.400 448.350 666.600 449.100 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 646.950 445.950 649.050 448.050 ;
        RECT 655.950 445.950 658.050 448.050 ;
        RECT 658.950 445.950 661.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 647.400 444.900 648.600 445.650 ;
        RECT 646.950 442.800 649.050 444.900 ;
        RECT 656.400 443.400 657.600 445.650 ;
        RECT 662.400 444.000 663.600 445.650 ;
        RECT 637.950 439.950 640.050 442.050 ;
        RECT 656.400 439.050 657.450 443.400 ;
        RECT 661.950 439.950 664.050 444.000 ;
        RECT 671.400 439.050 672.450 460.950 ;
        RECT 655.950 436.950 658.050 439.050 ;
        RECT 670.950 436.950 673.050 439.050 ;
        RECT 628.950 421.950 631.050 424.050 ;
        RECT 643.950 422.400 646.050 424.500 ;
        RECT 622.950 419.100 625.050 421.200 ;
        RECT 622.950 415.950 625.050 418.050 ;
        RECT 629.400 417.600 630.450 421.950 ;
        RECT 623.400 415.350 624.600 415.950 ;
        RECT 629.400 415.350 630.600 417.600 ;
        RECT 640.950 416.100 643.050 418.200 ;
        RECT 641.400 415.350 642.600 416.100 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 631.950 412.950 634.050 415.050 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 626.400 411.900 627.600 412.650 ;
        RECT 625.950 409.800 628.050 411.900 ;
        RECT 632.400 411.000 633.600 412.650 ;
        RECT 631.950 406.950 634.050 411.000 ;
        RECT 644.850 407.400 646.050 422.400 ;
        RECT 652.950 421.950 655.050 424.050 ;
        RECT 664.950 422.400 667.050 424.500 ;
        RECT 649.950 416.100 652.050 418.200 ;
        RECT 650.400 412.050 651.450 416.100 ;
        RECT 649.950 409.950 652.050 412.050 ;
        RECT 653.400 411.450 654.450 421.950 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 659.400 411.450 660.600 412.650 ;
        RECT 653.400 410.400 660.600 411.450 ;
        RECT 643.950 405.300 646.050 407.400 ;
        RECT 644.850 401.700 646.050 405.300 ;
        RECT 643.950 399.600 646.050 401.700 ;
        RECT 646.950 394.950 649.050 397.050 ;
        RECT 640.950 385.950 643.050 388.050 ;
        RECT 610.950 379.950 613.050 382.050 ;
        RECT 616.950 379.950 619.050 382.050 ;
        RECT 607.950 373.950 610.050 376.050 ;
        RECT 590.400 370.350 591.600 371.100 ;
        RECT 595.950 370.950 598.050 373.050 ;
        RECT 604.950 370.950 607.050 373.050 ;
        RECT 611.400 372.600 612.450 379.950 ;
        RECT 625.950 376.950 628.050 379.050 ;
        RECT 619.950 373.950 622.050 376.050 ;
        RECT 574.950 367.950 577.050 370.050 ;
        RECT 586.950 367.950 589.050 370.050 ;
        RECT 589.950 367.950 592.050 370.050 ;
        RECT 575.400 366.900 576.600 367.650 ;
        RECT 587.400 366.900 588.600 367.650 ;
        RECT 574.950 364.800 577.050 366.900 ;
        RECT 586.950 364.800 589.050 366.900 ;
        RECT 596.400 366.750 597.450 370.950 ;
        RECT 605.400 370.200 606.600 370.950 ;
        RECT 611.400 370.200 612.600 372.600 ;
        RECT 601.950 367.800 604.050 369.900 ;
        RECT 604.950 367.800 607.050 369.900 ;
        RECT 607.950 367.800 610.050 369.900 ;
        RECT 610.950 367.800 613.050 369.900 ;
        RECT 613.950 367.800 616.050 369.900 ;
        RECT 602.400 366.750 603.600 367.500 ;
        RECT 595.950 366.450 598.050 366.750 ;
        RECT 593.400 365.400 598.050 366.450 ;
        RECT 571.950 358.500 574.050 360.600 ;
        RECT 565.950 346.950 568.050 349.050 ;
        RECT 538.950 344.400 541.050 346.500 ;
        RECT 559.950 344.400 562.050 346.500 ;
        RECT 490.950 338.100 493.050 340.200 ;
        RECT 499.950 338.100 502.050 340.200 ;
        RECT 505.950 338.100 508.050 340.200 ;
        RECT 491.400 337.350 492.600 338.100 ;
        RECT 500.400 337.350 501.600 338.100 ;
        RECT 506.400 337.350 507.600 338.100 ;
        RECT 511.950 337.950 514.050 343.050 ;
        RECT 514.950 337.950 517.050 340.050 ;
        RECT 517.950 337.950 520.050 340.050 ;
        RECT 526.950 338.250 529.050 340.350 ;
        RECT 484.950 334.950 487.050 337.050 ;
        RECT 490.950 334.950 493.050 337.050 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 505.950 334.950 508.050 337.050 ;
        RECT 508.950 334.950 511.050 337.050 ;
        RECT 485.400 332.400 486.600 334.650 ;
        RECT 503.400 332.400 504.600 334.650 ;
        RECT 509.400 333.900 510.600 334.650 ;
        RECT 515.400 333.900 516.450 337.950 ;
        RECT 485.400 313.050 486.450 332.400 ;
        RECT 503.400 325.050 504.450 332.400 ;
        RECT 508.950 331.800 511.050 333.900 ;
        RECT 514.950 331.800 517.050 333.900 ;
        RECT 518.400 328.050 519.450 337.950 ;
        RECT 527.400 337.500 528.600 338.250 ;
        RECT 535.950 338.100 538.050 340.200 ;
        RECT 536.400 337.350 537.600 338.100 ;
        RECT 523.950 335.100 526.050 337.200 ;
        RECT 526.950 335.100 529.050 337.200 ;
        RECT 529.950 335.100 532.050 337.200 ;
        RECT 535.950 334.950 538.050 337.050 ;
        RECT 524.400 334.050 525.600 334.800 ;
        RECT 530.400 334.050 531.600 334.800 ;
        RECT 523.950 331.950 526.050 334.050 ;
        RECT 529.950 331.950 532.050 334.050 ;
        RECT 517.950 325.950 520.050 328.050 ;
        RECT 502.950 322.950 505.050 325.050 ;
        RECT 514.950 316.950 517.050 319.050 ;
        RECT 484.950 310.950 487.050 313.050 ;
        RECT 485.400 295.050 486.450 310.950 ;
        RECT 478.950 292.950 481.050 295.050 ;
        RECT 484.950 292.950 487.050 295.050 ;
        RECT 490.950 292.950 493.050 295.050 ;
        RECT 496.950 292.950 499.050 295.050 ;
        RECT 479.400 288.750 480.450 292.950 ;
        RECT 491.400 292.200 492.600 292.950 ;
        RECT 484.950 289.800 487.050 291.900 ;
        RECT 490.950 289.800 493.050 291.900 ;
        RECT 485.400 288.750 486.600 289.500 ;
        RECT 478.950 286.650 481.050 288.750 ;
        RECT 484.950 286.650 487.050 288.750 ;
        RECT 485.400 280.050 486.450 286.650 ;
        RECT 484.950 277.950 487.050 280.050 ;
        RECT 497.400 274.050 498.450 292.950 ;
        RECT 508.950 289.800 511.050 291.900 ;
        RECT 496.950 271.950 499.050 274.050 ;
        RECT 484.950 266.400 487.050 268.500 ;
        RECT 505.950 266.400 508.050 268.500 ;
        RECT 475.950 262.950 478.050 265.050 ;
        RECT 472.950 260.250 475.050 262.350 ;
        RECT 473.400 259.500 474.600 260.250 ;
        RECT 469.950 257.100 472.050 259.200 ;
        RECT 472.950 257.100 475.050 259.200 ;
        RECT 475.950 257.100 478.050 259.200 ;
        RECT 481.950 256.950 484.050 259.050 ;
        RECT 470.400 254.400 471.600 256.800 ;
        RECT 476.400 255.000 477.600 256.800 ;
        RECT 470.400 250.050 471.450 254.400 ;
        RECT 475.950 250.950 478.050 255.000 ;
        RECT 482.400 254.400 483.600 256.650 ;
        RECT 482.400 250.050 483.450 254.400 ;
        RECT 469.950 247.950 472.050 250.050 ;
        RECT 481.950 247.950 484.050 250.050 ;
        RECT 485.700 246.600 486.900 266.400 ;
        RECT 496.950 262.950 499.050 265.050 ;
        RECT 490.950 256.950 493.050 259.050 ;
        RECT 491.400 254.400 492.600 256.650 ;
        RECT 484.950 244.500 487.050 246.600 ;
        RECT 491.400 244.050 492.450 254.400 ;
        RECT 490.950 241.950 493.050 244.050 ;
        RECT 464.400 230.400 468.450 231.450 ;
        RECT 460.950 224.400 463.050 226.500 ;
        RECT 454.950 215.100 457.050 217.200 ;
        RECT 455.400 214.350 456.600 215.100 ;
        RECT 454.950 211.950 457.050 214.050 ;
        RECT 461.100 204.600 462.300 224.400 ;
        RECT 464.400 216.450 465.600 216.600 ;
        RECT 467.400 216.450 468.450 230.400 ;
        RECT 497.400 229.050 498.450 262.950 ;
        RECT 499.950 260.100 502.050 262.200 ;
        RECT 500.400 253.050 501.450 260.100 ;
        RECT 499.950 250.950 502.050 253.050 ;
        RECT 505.950 251.400 507.150 266.400 ;
        RECT 508.950 260.100 511.050 262.200 ;
        RECT 509.400 259.350 510.600 260.100 ;
        RECT 508.950 256.950 511.050 259.050 ;
        RECT 515.400 256.050 516.450 316.950 ;
        RECT 524.400 298.050 525.450 331.950 ;
        RECT 530.400 304.050 531.450 331.950 ;
        RECT 532.950 328.950 535.050 331.050 ;
        RECT 539.850 329.400 541.050 344.400 ;
        RECT 553.950 334.950 556.050 337.050 ;
        RECT 533.400 310.050 534.450 328.950 ;
        RECT 538.950 327.300 541.050 329.400 ;
        RECT 554.400 332.400 555.600 334.650 ;
        RECT 554.400 328.050 555.450 332.400 ;
        RECT 539.850 323.700 541.050 327.300 ;
        RECT 553.950 325.950 556.050 328.050 ;
        RECT 560.100 324.600 561.300 344.400 ;
        RECT 575.400 339.450 576.600 339.600 ;
        RECT 569.400 338.400 576.600 339.450 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 563.400 333.900 564.600 334.650 ;
        RECT 562.950 330.450 565.050 333.900 ;
        RECT 562.950 329.400 567.450 330.450 ;
        RECT 562.950 328.950 565.050 329.400 ;
        RECT 538.950 321.600 541.050 323.700 ;
        RECT 559.950 322.500 562.050 324.600 ;
        RECT 532.950 307.950 535.050 310.050 ;
        RECT 529.950 301.950 532.050 304.050 ;
        RECT 533.400 300.450 534.450 307.950 ;
        RECT 547.950 304.950 550.050 307.050 ;
        RECT 535.950 301.950 538.050 304.050 ;
        RECT 530.400 299.400 534.450 300.450 ;
        RECT 523.950 295.950 526.050 298.050 ;
        RECT 530.400 294.600 531.450 299.400 ;
        RECT 530.400 292.200 531.600 294.600 ;
        RECT 529.950 289.800 532.050 291.900 ;
        RECT 536.400 262.350 537.450 301.950 ;
        RECT 544.950 294.000 547.050 298.050 ;
        RECT 548.400 295.050 549.450 304.950 ;
        RECT 559.950 303.300 562.050 305.400 ;
        RECT 560.850 299.700 562.050 303.300 ;
        RECT 559.950 297.600 562.050 299.700 ;
        RECT 545.400 292.200 546.600 294.000 ;
        RECT 547.800 292.950 549.900 295.050 ;
        RECT 550.950 292.950 553.050 295.050 ;
        RECT 551.400 292.200 552.600 292.950 ;
        RECT 544.950 289.800 547.050 291.900 ;
        RECT 547.950 289.800 550.050 291.900 ;
        RECT 550.950 289.800 553.050 291.900 ;
        RECT 556.950 289.950 559.050 292.050 ;
        RECT 548.400 288.750 549.600 289.500 ;
        RECT 557.400 288.900 558.600 289.650 ;
        RECT 547.800 286.650 549.900 288.750 ;
        RECT 556.950 286.800 559.050 288.900 ;
        RECT 560.850 282.600 562.050 297.600 ;
        RECT 566.400 295.200 567.450 329.400 ;
        RECT 569.400 313.050 570.450 338.400 ;
        RECT 575.400 337.350 576.600 338.400 ;
        RECT 580.950 338.100 583.050 340.200 ;
        RECT 589.950 338.100 592.050 340.200 ;
        RECT 581.400 337.350 582.600 338.100 ;
        RECT 574.950 334.950 577.050 337.050 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 578.400 333.900 579.600 334.650 ;
        RECT 577.950 331.800 580.050 333.900 ;
        RECT 584.400 332.400 585.600 334.650 ;
        RECT 584.400 325.050 585.450 332.400 ;
        RECT 590.400 328.050 591.450 338.100 ;
        RECT 589.950 325.950 592.050 328.050 ;
        RECT 583.950 322.950 586.050 325.050 ;
        RECT 589.950 322.800 592.050 324.900 ;
        RECT 568.950 310.950 571.050 313.050 ;
        RECT 580.950 302.400 583.050 304.500 ;
        RECT 574.950 298.950 577.050 301.050 ;
        RECT 568.950 295.950 571.050 298.050 ;
        RECT 565.950 293.100 568.050 295.200 ;
        RECT 559.950 280.500 562.050 282.600 ;
        RECT 566.400 277.050 567.450 293.100 ;
        RECT 569.400 283.050 570.450 295.950 ;
        RECT 575.400 294.600 576.450 298.950 ;
        RECT 575.400 292.350 576.600 294.600 ;
        RECT 574.950 289.950 577.050 292.050 ;
        RECT 571.950 286.950 574.050 289.050 ;
        RECT 568.950 280.950 571.050 283.050 ;
        RECT 556.950 274.950 559.050 277.050 ;
        RECT 565.950 274.950 568.050 277.050 ;
        RECT 544.950 266.400 547.050 268.500 ;
        RECT 557.400 268.050 558.450 274.950 ;
        RECT 523.950 260.250 526.050 262.350 ;
        RECT 529.950 260.250 532.050 262.350 ;
        RECT 535.950 260.250 538.050 262.350 ;
        RECT 524.400 259.500 525.600 260.250 ;
        RECT 530.400 259.500 531.600 260.250 ;
        RECT 520.950 257.100 523.050 259.200 ;
        RECT 523.950 257.100 526.050 259.200 ;
        RECT 526.950 257.100 529.050 259.200 ;
        RECT 529.950 257.100 532.050 259.200 ;
        RECT 532.950 257.100 535.050 259.200 ;
        RECT 541.950 256.950 544.050 259.050 ;
        RECT 521.400 256.050 522.600 256.800 ;
        RECT 514.950 253.950 517.050 256.050 ;
        RECT 520.950 253.950 523.050 256.050 ;
        RECT 527.400 254.400 528.600 256.800 ;
        RECT 533.400 254.400 534.600 256.800 ;
        RECT 542.400 255.900 543.600 256.650 ;
        RECT 505.950 249.300 508.050 251.400 ;
        RECT 499.950 244.950 502.050 247.050 ;
        RECT 505.950 245.700 507.150 249.300 ;
        RECT 500.400 238.050 501.450 244.950 ;
        RECT 505.950 243.600 508.050 245.700 ;
        RECT 499.950 235.950 502.050 238.050 ;
        RECT 472.950 226.950 475.050 229.050 ;
        RECT 496.950 226.950 499.050 229.050 ;
        RECT 464.400 215.400 468.450 216.450 ;
        RECT 464.400 214.350 465.600 215.400 ;
        RECT 463.950 211.950 466.050 214.050 ;
        RECT 460.950 202.500 463.050 204.600 ;
        RECT 448.950 184.950 451.050 187.050 ;
        RECT 440.400 181.500 441.600 183.000 ;
        RECT 446.400 181.500 447.600 183.600 ;
        RECT 436.950 179.100 439.050 181.200 ;
        RECT 439.950 179.100 442.050 181.200 ;
        RECT 442.950 179.100 445.050 181.200 ;
        RECT 445.950 179.100 448.050 181.200 ;
        RECT 448.950 179.100 451.050 181.200 ;
        RECT 463.950 179.100 466.050 181.200 ;
        RECT 428.400 170.400 432.450 171.450 ;
        RECT 437.400 176.400 438.600 178.800 ;
        RECT 443.400 176.400 444.600 178.800 ;
        RECT 449.400 177.000 450.600 178.800 ;
        RECT 415.950 141.600 418.050 143.700 ;
        RECT 424.950 142.950 427.050 145.050 ;
        RECT 404.400 140.400 408.450 141.450 ;
        RECT 400.950 137.100 403.050 139.200 ;
        RECT 401.400 136.350 402.600 137.100 ;
        RECT 400.950 133.950 403.050 136.050 ;
        RECT 394.950 124.500 397.050 126.600 ;
        RECT 400.950 121.950 403.050 124.050 ;
        RECT 385.950 118.950 388.050 121.050 ;
        RECT 382.950 115.950 385.050 118.050 ;
        RECT 376.950 109.950 379.050 112.050 ;
        RECT 383.400 105.600 384.450 115.950 ;
        RECT 394.950 112.950 397.050 115.050 ;
        RECT 395.400 105.600 396.450 112.950 ;
        RECT 401.400 105.600 402.450 121.950 ;
        RECT 403.950 115.950 406.050 118.050 ;
        RECT 404.400 109.050 405.450 115.950 ;
        RECT 403.950 106.950 406.050 109.050 ;
        RECT 383.400 103.350 384.600 105.600 ;
        RECT 395.400 103.500 396.600 105.600 ;
        RECT 401.400 103.500 402.600 105.600 ;
        RECT 407.400 105.450 408.450 140.400 ;
        RECT 409.950 136.950 412.050 139.050 ;
        RECT 410.400 124.050 411.450 136.950 ;
        RECT 415.950 126.600 417.150 141.600 ;
        RECT 418.950 133.950 421.050 136.050 ;
        RECT 419.400 131.400 420.600 133.650 ;
        RECT 419.400 129.450 420.450 131.400 ;
        RECT 419.400 128.400 423.450 129.450 ;
        RECT 415.950 124.500 418.050 126.600 ;
        RECT 409.950 121.950 412.050 124.050 ;
        RECT 410.400 109.050 411.450 121.950 ;
        RECT 422.400 115.050 423.450 128.400 ;
        RECT 412.950 112.950 415.050 115.050 ;
        RECT 421.950 112.950 424.050 115.050 ;
        RECT 409.950 106.950 412.050 109.050 ;
        RECT 407.400 104.400 411.450 105.450 ;
        RECT 379.950 100.950 382.050 103.050 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 391.950 101.100 394.050 103.200 ;
        RECT 394.950 101.100 397.050 103.200 ;
        RECT 397.950 101.100 400.050 103.200 ;
        RECT 400.950 101.100 403.050 103.200 ;
        RECT 403.950 101.100 406.050 103.200 ;
        RECT 352.950 94.950 355.050 97.050 ;
        RECT 349.950 88.950 352.050 91.050 ;
        RECT 359.400 85.050 360.450 98.400 ;
        RECT 364.950 94.950 367.050 99.000 ;
        RECT 373.950 97.950 376.050 100.050 ;
        RECT 380.400 99.900 381.600 100.650 ;
        RECT 392.400 100.050 393.600 100.800 ;
        RECT 379.950 97.800 382.050 99.900 ;
        RECT 391.950 97.950 394.050 100.050 ;
        RECT 398.400 98.400 399.600 100.800 ;
        RECT 404.400 100.050 405.600 100.800 ;
        RECT 376.950 88.950 379.050 91.050 ;
        RECT 377.400 85.050 378.450 88.950 ;
        RECT 382.950 85.950 385.050 88.050 ;
        RECT 358.950 82.950 361.050 85.050 ;
        RECT 376.950 82.950 379.050 85.050 ;
        RECT 355.950 76.950 358.050 79.050 ;
        RECT 286.950 67.950 289.050 70.050 ;
        RECT 301.950 67.950 304.050 70.050 ;
        RECT 337.950 67.950 340.050 70.050 ;
        RECT 343.950 68.400 346.050 70.500 ;
        RECT 356.400 70.050 357.450 76.950 ;
        RECT 287.400 61.050 288.450 67.950 ;
        RECT 292.950 64.950 295.050 67.050 ;
        RECT 298.950 64.950 301.050 67.050 ;
        RECT 286.950 58.950 289.050 61.050 ;
        RECT 293.400 60.600 294.450 64.950 ;
        RECT 287.400 58.200 288.600 58.950 ;
        RECT 293.400 58.200 294.600 60.600 ;
        RECT 286.950 55.800 289.050 57.900 ;
        RECT 289.950 55.800 292.050 57.900 ;
        RECT 292.950 55.800 295.050 57.900 ;
        RECT 290.400 54.750 291.600 55.500 ;
        RECT 289.950 52.650 292.050 54.750 ;
        RECT 295.950 52.950 298.050 55.050 ;
        RECT 280.950 49.950 283.050 52.050 ;
        RECT 250.950 46.500 253.050 48.600 ;
        RECT 271.950 46.950 274.050 49.050 ;
        RECT 277.950 46.950 280.050 49.050 ;
        RECT 238.950 34.950 241.050 37.050 ;
        RECT 212.400 25.350 213.600 27.600 ;
        RECT 217.950 27.000 220.050 31.050 ;
        RECT 218.400 25.350 219.600 27.000 ;
        RECT 223.950 25.950 226.050 28.050 ;
        RECT 232.950 26.100 235.050 28.200 ;
        RECT 239.400 27.600 240.450 34.950 ;
        RECT 259.950 31.950 262.050 34.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 215.400 21.000 216.600 22.650 ;
        RECT 224.400 21.900 225.450 25.950 ;
        RECT 233.400 25.350 234.600 26.100 ;
        RECT 239.400 25.350 240.600 27.600 ;
        RECT 250.950 26.250 253.050 28.350 ;
        RECT 251.400 25.500 252.600 26.250 ;
        RECT 229.950 22.950 232.050 25.050 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 247.950 23.100 250.050 25.200 ;
        RECT 250.950 23.100 253.050 25.200 ;
        RECT 253.950 23.100 256.050 25.200 ;
        RECT 230.400 21.900 231.600 22.650 ;
        RECT 205.950 16.950 208.050 19.050 ;
        RECT 214.950 16.950 217.050 21.000 ;
        RECT 223.950 19.800 226.050 21.900 ;
        RECT 229.950 19.800 232.050 21.900 ;
        RECT 236.400 21.000 237.600 22.650 ;
        RECT 248.400 22.050 249.600 22.800 ;
        RECT 254.400 22.050 255.600 22.800 ;
        RECT 260.400 22.050 261.450 31.950 ;
        RECT 281.400 31.050 282.450 49.950 ;
        RECT 296.400 37.050 297.450 52.950 ;
        RECT 295.950 34.950 298.050 37.050 ;
        RECT 272.400 29.400 279.450 30.450 ;
        RECT 272.400 27.600 273.450 29.400 ;
        RECT 272.400 25.500 273.600 27.600 ;
        RECT 278.400 27.450 279.450 29.400 ;
        RECT 280.950 28.950 283.050 31.050 ;
        RECT 278.400 26.400 282.450 27.450 ;
        RECT 268.950 23.100 271.050 25.200 ;
        RECT 271.950 23.100 274.050 25.200 ;
        RECT 274.950 23.100 277.050 25.200 ;
        RECT 269.400 22.050 270.600 22.800 ;
        RECT 275.400 22.050 276.600 22.800 ;
        RECT 235.950 16.950 238.050 21.000 ;
        RECT 247.950 19.950 250.050 22.050 ;
        RECT 248.400 16.050 249.450 19.950 ;
        RECT 253.950 16.950 256.050 22.050 ;
        RECT 259.950 19.950 262.050 22.050 ;
        RECT 268.950 19.950 271.050 22.050 ;
        RECT 274.950 19.950 277.050 22.050 ;
        RECT 281.400 21.900 282.450 26.400 ;
        RECT 289.950 26.100 292.050 28.200 ;
        RECT 296.400 27.600 297.450 34.950 ;
        RECT 299.400 34.050 300.450 64.950 ;
        RECT 302.400 46.050 303.450 67.950 ;
        RECT 328.950 63.450 331.050 64.050 ;
        RECT 334.950 63.450 337.050 64.050 ;
        RECT 328.950 62.400 337.050 63.450 ;
        RECT 328.950 61.950 331.050 62.400 ;
        RECT 334.950 61.950 337.050 62.400 ;
        RECT 307.950 58.950 310.050 61.050 ;
        RECT 313.950 58.950 316.050 61.050 ;
        RECT 319.950 59.100 322.050 61.200 ;
        RECT 325.950 59.100 328.050 61.200 ;
        RECT 331.950 59.100 334.050 61.200 ;
        RECT 338.400 60.450 339.450 67.950 ;
        RECT 341.400 60.450 342.600 60.600 ;
        RECT 338.400 59.400 342.600 60.450 ;
        RECT 308.400 58.200 309.600 58.950 ;
        RECT 314.400 58.200 315.600 58.950 ;
        RECT 307.950 55.800 310.050 57.900 ;
        RECT 310.950 55.800 313.050 57.900 ;
        RECT 313.950 55.800 316.050 57.900 ;
        RECT 311.400 53.400 312.600 55.500 ;
        RECT 311.400 52.050 312.450 53.400 ;
        RECT 320.400 52.050 321.450 59.100 ;
        RECT 326.400 58.350 327.600 59.100 ;
        RECT 332.400 58.350 333.600 59.100 ;
        RECT 341.400 58.350 342.600 59.400 ;
        RECT 325.950 55.950 328.050 58.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 340.950 55.950 343.050 58.050 ;
        RECT 329.400 54.900 330.600 55.650 ;
        RECT 328.950 52.800 331.050 54.900 ;
        RECT 335.400 53.400 336.600 55.650 ;
        RECT 311.400 50.400 316.050 52.050 ;
        RECT 312.000 49.950 316.050 50.400 ;
        RECT 319.950 49.950 322.050 52.050 ;
        RECT 301.950 43.950 304.050 46.050 ;
        RECT 319.950 43.950 322.050 46.050 ;
        RECT 298.950 31.950 301.050 34.050 ;
        RECT 304.950 32.400 307.050 34.500 ;
        RECT 290.400 25.350 291.600 26.100 ;
        RECT 296.400 25.350 297.600 27.600 ;
        RECT 286.950 22.950 289.050 25.050 ;
        RECT 289.950 22.950 292.050 25.050 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 287.400 21.900 288.600 22.650 ;
        RECT 280.950 19.800 283.050 21.900 ;
        RECT 286.950 19.800 289.050 21.900 ;
        RECT 293.400 20.400 294.600 22.650 ;
        RECT 293.400 16.050 294.450 20.400 ;
        RECT 298.800 19.950 300.900 22.050 ;
        RECT 302.400 21.900 303.600 22.650 ;
        RECT 172.950 10.500 175.050 12.600 ;
        RECT 184.950 10.950 187.050 13.050 ;
        RECT 193.950 11.700 195.150 15.300 ;
        RECT 202.950 13.950 205.050 16.050 ;
        RECT 232.950 15.450 235.050 16.050 ;
        RECT 238.950 15.450 241.050 16.050 ;
        RECT 232.950 14.400 241.050 15.450 ;
        RECT 232.950 13.950 235.050 14.400 ;
        RECT 238.950 13.950 241.050 14.400 ;
        RECT 247.950 13.950 250.050 16.050 ;
        RECT 292.950 13.950 295.050 16.050 ;
        RECT 299.400 13.050 300.450 19.950 ;
        RECT 301.950 19.800 304.050 21.900 ;
        RECT 193.950 9.600 196.050 11.700 ;
        RECT 298.950 10.950 301.050 13.050 ;
        RECT 305.700 12.600 306.900 32.400 ;
        RECT 310.950 22.950 313.050 25.050 ;
        RECT 311.400 20.400 312.600 22.650 ;
        RECT 320.400 21.900 321.450 43.950 ;
        RECT 335.400 40.050 336.450 53.400 ;
        RECT 344.700 48.600 345.900 68.400 ;
        RECT 355.950 67.950 358.050 70.050 ;
        RECT 364.950 69.300 367.050 71.400 ;
        RECT 349.950 60.000 352.050 64.050 ;
        RECT 350.400 58.350 351.600 60.000 ;
        RECT 349.950 55.950 352.050 58.050 ;
        RECT 343.950 46.500 346.050 48.600 ;
        RECT 356.400 43.050 357.450 67.950 ;
        RECT 364.950 65.700 366.150 69.300 ;
        RECT 383.400 67.050 384.450 85.950 ;
        RECT 398.400 79.050 399.450 98.400 ;
        RECT 403.950 97.950 406.050 100.050 ;
        RECT 397.950 76.950 400.050 79.050 ;
        RECT 410.400 70.050 411.450 104.400 ;
        RECT 413.400 100.050 414.450 112.950 ;
        RECT 425.400 106.350 426.450 142.950 ;
        RECT 428.400 121.050 429.450 170.400 ;
        RECT 437.400 166.050 438.450 176.400 ;
        RECT 436.950 163.950 439.050 166.050 ;
        RECT 443.400 148.050 444.450 176.400 ;
        RECT 448.950 172.950 451.050 177.000 ;
        RECT 473.400 175.050 474.450 226.950 ;
        RECT 500.400 217.050 501.450 235.950 ;
        RECT 515.400 226.050 516.450 253.950 ;
        RECT 527.400 247.050 528.450 254.400 ;
        RECT 529.950 247.950 532.050 250.050 ;
        RECT 526.950 244.950 529.050 247.050 ;
        RECT 514.950 223.950 517.050 226.050 ;
        RECT 490.950 214.950 493.050 217.050 ;
        RECT 499.950 214.950 502.050 217.050 ;
        RECT 505.950 214.950 508.050 217.050 ;
        RECT 511.950 214.950 514.050 217.050 ;
        RECT 517.950 214.950 520.050 217.050 ;
        RECT 478.950 211.800 481.050 213.900 ;
        RECT 475.950 184.950 478.050 187.050 ;
        RECT 472.950 172.950 475.050 175.050 ;
        RECT 476.400 151.050 477.450 184.950 ;
        RECT 484.950 179.100 487.050 181.200 ;
        RECT 478.950 175.950 481.050 178.050 ;
        RECT 485.400 176.400 486.600 178.800 ;
        RECT 491.400 177.900 492.450 214.950 ;
        RECT 500.400 214.200 501.600 214.950 ;
        RECT 499.950 211.800 502.050 213.900 ;
        RECT 499.950 205.950 502.050 208.050 ;
        RECT 500.400 183.600 501.450 205.950 ;
        RECT 506.400 202.050 507.450 214.950 ;
        RECT 512.400 214.200 513.600 214.950 ;
        RECT 518.400 214.200 519.600 214.950 ;
        RECT 511.950 211.800 514.050 213.900 ;
        RECT 514.950 211.800 517.050 213.900 ;
        RECT 517.950 211.800 520.050 213.900 ;
        RECT 520.950 211.800 523.050 213.900 ;
        RECT 515.400 210.000 516.600 211.500 ;
        RECT 521.400 210.750 522.600 211.500 ;
        RECT 530.400 211.050 531.450 247.950 ;
        RECT 533.400 229.050 534.450 254.400 ;
        RECT 541.950 253.800 544.050 255.900 ;
        RECT 545.700 246.600 546.900 266.400 ;
        RECT 556.950 265.950 559.050 268.050 ;
        RECT 565.950 266.400 568.050 268.500 ;
        RECT 550.950 256.950 553.050 259.050 ;
        RECT 551.400 254.400 552.600 256.650 ;
        RECT 557.400 255.900 558.450 265.950 ;
        RECT 559.950 260.100 562.050 262.200 ;
        RECT 551.400 250.050 552.450 254.400 ;
        RECT 556.950 253.800 559.050 255.900 ;
        RECT 550.950 247.950 553.050 250.050 ;
        RECT 544.950 244.500 547.050 246.600 ;
        RECT 544.950 238.950 547.050 241.050 ;
        RECT 532.950 226.950 535.050 229.050 ;
        RECT 538.950 215.100 541.050 217.200 ;
        RECT 545.400 217.050 546.450 238.950 ;
        RECT 557.400 228.450 558.450 253.800 ;
        RECT 560.400 241.050 561.450 260.100 ;
        RECT 565.950 251.400 567.150 266.400 ;
        RECT 568.950 260.100 571.050 262.200 ;
        RECT 572.400 261.450 573.450 286.950 ;
        RECT 581.100 282.600 582.300 302.400 ;
        RECT 583.950 293.100 586.050 295.200 ;
        RECT 584.400 292.350 585.600 293.100 ;
        RECT 583.950 289.950 586.050 292.050 ;
        RECT 590.400 288.450 591.450 322.800 ;
        RECT 593.400 316.050 594.450 365.400 ;
        RECT 595.950 364.650 598.050 365.400 ;
        RECT 601.950 364.650 604.050 366.750 ;
        RECT 608.400 365.400 609.600 367.500 ;
        RECT 614.400 366.750 615.600 367.500 ;
        RECT 620.400 366.750 621.450 373.950 ;
        RECT 626.400 372.600 627.450 376.950 ;
        RECT 626.400 370.200 627.600 372.600 ;
        RECT 634.950 370.950 637.050 373.050 ;
        RECT 635.400 370.200 636.600 370.950 ;
        RECT 625.950 367.800 628.050 369.900 ;
        RECT 631.950 367.800 634.050 369.900 ;
        RECT 634.950 367.800 637.050 369.900 ;
        RECT 632.400 366.750 633.600 367.500 ;
        RECT 608.400 361.050 609.450 365.400 ;
        RECT 613.950 364.650 616.050 366.750 ;
        RECT 619.950 364.650 622.050 366.750 ;
        RECT 631.950 364.650 634.050 366.750 ;
        RECT 607.950 358.950 610.050 361.050 ;
        RECT 641.400 352.050 642.450 385.950 ;
        RECT 643.950 376.950 646.050 379.050 ;
        RECT 625.950 349.950 628.050 352.050 ;
        RECT 640.950 349.950 643.050 352.050 ;
        RECT 610.950 344.400 613.050 346.500 ;
        RECT 601.950 339.000 604.050 343.050 ;
        RECT 602.400 337.350 603.600 339.000 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 601.950 334.950 604.050 337.050 ;
        RECT 607.950 334.950 610.050 337.050 ;
        RECT 599.400 333.900 600.600 334.650 ;
        RECT 598.950 331.800 601.050 333.900 ;
        RECT 608.400 333.000 609.600 334.650 ;
        RECT 607.950 328.950 610.050 333.000 ;
        RECT 611.700 324.600 612.900 344.400 ;
        RECT 616.950 334.950 619.050 337.050 ;
        RECT 617.400 332.400 618.600 334.650 ;
        RECT 617.400 328.050 618.450 332.400 ;
        RECT 616.950 325.950 619.050 328.050 ;
        RECT 610.950 322.500 613.050 324.600 ;
        RECT 592.950 313.950 595.050 316.050 ;
        RECT 613.950 313.950 616.050 316.050 ;
        RECT 604.950 307.950 607.050 310.050 ;
        RECT 598.950 304.950 601.050 307.050 ;
        RECT 592.950 298.950 595.050 301.050 ;
        RECT 593.400 289.050 594.450 298.950 ;
        RECT 599.400 294.600 600.450 304.950 ;
        RECT 605.400 294.600 606.450 307.950 ;
        RECT 599.400 292.350 600.600 294.600 ;
        RECT 605.400 292.350 606.600 294.600 ;
        RECT 598.950 289.950 601.050 292.050 ;
        RECT 601.950 289.950 604.050 292.050 ;
        RECT 604.950 289.950 607.050 292.050 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 587.400 287.400 591.450 288.450 ;
        RECT 580.950 280.500 583.050 282.600 ;
        RECT 587.400 261.600 588.450 287.400 ;
        RECT 592.950 286.950 595.050 289.050 ;
        RECT 602.400 288.900 603.600 289.650 ;
        RECT 608.400 288.900 609.600 289.650 ;
        RECT 601.950 286.800 604.050 288.900 ;
        RECT 607.950 286.800 610.050 288.900 ;
        RECT 608.400 283.050 609.450 286.800 ;
        RECT 607.950 280.950 610.050 283.050 ;
        RECT 598.950 277.950 601.050 280.050 ;
        RECT 599.400 262.200 600.450 277.950 ;
        RECT 572.400 260.400 576.450 261.450 ;
        RECT 569.400 259.350 570.600 260.100 ;
        RECT 568.950 256.950 571.050 259.050 ;
        RECT 565.950 249.300 568.050 251.400 ;
        RECT 565.950 245.700 567.150 249.300 ;
        RECT 565.950 243.600 568.050 245.700 ;
        RECT 559.950 238.950 562.050 241.050 ;
        RECT 575.400 232.050 576.450 260.400 ;
        RECT 587.400 259.500 588.600 261.600 ;
        RECT 598.950 260.100 601.050 262.200 ;
        RECT 604.950 260.100 607.050 262.200 ;
        RECT 599.400 259.350 600.600 260.100 ;
        RECT 605.400 259.350 606.600 260.100 ;
        RECT 583.950 257.100 586.050 259.200 ;
        RECT 586.950 257.100 589.050 259.200 ;
        RECT 589.950 257.100 592.050 259.200 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 604.950 256.950 607.050 259.050 ;
        RECT 607.950 256.950 610.050 259.050 ;
        RECT 584.400 254.400 585.600 256.800 ;
        RECT 590.400 256.050 591.600 256.800 ;
        RECT 580.950 244.950 583.050 247.050 ;
        RECT 574.950 229.950 577.050 232.050 ;
        RECT 557.400 227.400 561.450 228.450 ;
        RECT 556.950 223.950 559.050 226.050 ;
        RECT 539.400 214.350 540.600 215.100 ;
        RECT 544.950 214.950 547.050 217.050 ;
        RECT 550.950 214.950 553.050 217.050 ;
        RECT 557.400 216.600 558.450 223.950 ;
        RECT 560.400 217.200 561.450 227.400 ;
        RECT 571.950 224.400 574.050 226.500 ;
        RECT 551.400 214.200 552.600 214.950 ;
        RECT 557.400 214.200 558.600 216.600 ;
        RECT 559.950 215.100 562.050 217.200 ;
        RECT 568.950 215.100 571.050 220.050 ;
        RECT 569.400 214.350 570.600 215.100 ;
        RECT 535.950 211.950 538.050 214.050 ;
        RECT 538.950 211.950 541.050 214.050 ;
        RECT 541.950 211.950 544.050 214.050 ;
        RECT 550.950 211.800 553.050 213.900 ;
        RECT 553.950 211.800 556.050 213.900 ;
        RECT 556.950 211.800 559.050 213.900 ;
        RECT 559.950 211.800 562.050 213.900 ;
        RECT 568.950 211.950 571.050 214.050 ;
        RECT 514.950 205.950 517.050 210.000 ;
        RECT 520.950 208.650 523.050 210.750 ;
        RECT 529.950 208.950 532.050 211.050 ;
        RECT 536.400 210.000 537.600 211.650 ;
        RECT 542.400 210.900 543.600 211.650 ;
        RECT 535.950 205.950 538.050 210.000 ;
        RECT 541.950 208.800 544.050 210.900 ;
        RECT 547.950 208.950 550.050 211.050 ;
        RECT 554.400 209.400 555.600 211.500 ;
        RECT 560.400 210.750 561.600 211.500 ;
        RECT 505.950 199.950 508.050 202.050 ;
        RECT 544.950 190.950 547.050 193.050 ;
        RECT 517.950 188.400 520.050 190.500 ;
        RECT 538.950 188.400 541.050 190.500 ;
        RECT 500.400 181.500 501.600 183.600 ;
        RECT 505.950 182.250 508.050 184.350 ;
        RECT 506.400 181.500 507.600 182.250 ;
        RECT 496.950 179.100 499.050 181.200 ;
        RECT 499.950 179.100 502.050 181.200 ;
        RECT 502.950 179.100 505.050 181.200 ;
        RECT 505.950 179.100 508.050 181.200 ;
        RECT 514.950 178.950 517.050 181.050 ;
        RECT 479.400 160.050 480.450 175.950 ;
        RECT 485.400 166.050 486.450 176.400 ;
        RECT 490.950 175.800 493.050 177.900 ;
        RECT 497.400 176.400 498.600 178.800 ;
        RECT 503.400 176.400 504.600 178.800 ;
        RECT 484.950 163.950 487.050 166.050 ;
        RECT 478.950 157.950 481.050 160.050 ;
        RECT 442.950 145.950 445.050 148.050 ;
        RECT 448.950 146.400 451.050 148.500 ;
        RECT 469.950 147.300 472.050 149.400 ;
        RECT 475.950 148.950 478.050 151.050 ;
        RECT 433.950 136.950 436.050 139.050 ;
        RECT 439.950 136.950 442.050 139.050 ;
        RECT 445.950 138.000 448.050 142.050 ;
        RECT 434.400 136.200 435.600 136.950 ;
        RECT 440.400 136.200 441.600 136.950 ;
        RECT 446.400 136.350 447.600 138.000 ;
        RECT 433.950 133.800 436.050 135.900 ;
        RECT 436.950 133.800 439.050 135.900 ;
        RECT 439.950 133.800 442.050 135.900 ;
        RECT 445.950 133.950 448.050 136.050 ;
        RECT 430.950 130.950 433.050 133.050 ;
        RECT 437.400 131.400 438.600 133.500 ;
        RECT 427.950 118.950 430.050 121.050 ;
        RECT 431.400 112.050 432.450 130.950 ;
        RECT 437.400 112.050 438.450 131.400 ;
        RECT 449.700 126.600 450.900 146.400 ;
        RECT 469.950 143.700 471.150 147.300 ;
        RECT 469.950 141.600 472.050 143.700 ;
        RECT 479.400 142.050 480.450 157.950 ;
        RECT 454.950 137.100 457.050 139.200 ;
        RECT 460.950 137.100 463.050 139.200 ;
        RECT 455.400 136.350 456.600 137.100 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 448.950 124.500 451.050 126.600 ;
        RECT 454.950 121.950 457.050 124.050 ;
        RECT 448.950 118.950 451.050 121.050 ;
        RECT 430.950 109.950 433.050 112.050 ;
        RECT 436.950 109.950 439.050 112.050 ;
        RECT 418.950 104.250 421.050 106.350 ;
        RECT 424.950 104.250 427.050 106.350 ;
        RECT 431.400 105.600 432.450 109.950 ;
        RECT 438.000 108.450 442.050 109.050 ;
        RECT 437.400 106.950 442.050 108.450 ;
        RECT 445.950 106.950 448.050 109.050 ;
        RECT 437.400 105.600 438.450 106.950 ;
        RECT 419.400 103.500 420.600 104.250 ;
        RECT 431.400 103.350 432.600 105.600 ;
        RECT 437.400 103.350 438.600 105.600 ;
        RECT 418.950 101.100 421.050 103.200 ;
        RECT 421.950 101.100 424.050 103.200 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 436.950 100.950 439.050 103.050 ;
        RECT 439.950 100.950 442.050 103.050 ;
        RECT 422.400 100.050 423.600 100.800 ;
        RECT 412.950 97.950 415.050 100.050 ;
        RECT 421.950 97.950 424.050 100.050 ;
        RECT 434.400 98.400 435.600 100.650 ;
        RECT 440.400 99.900 441.600 100.650 ;
        RECT 434.400 91.050 435.450 98.400 ;
        RECT 439.950 97.800 442.050 99.900 ;
        RECT 446.400 97.050 447.450 106.950 ;
        RECT 445.950 94.950 448.050 97.050 ;
        RECT 445.950 91.800 448.050 93.900 ;
        RECT 415.950 88.950 418.050 91.050 ;
        RECT 433.950 88.950 436.050 91.050 ;
        RECT 409.950 67.950 412.050 70.050 ;
        RECT 364.950 63.600 367.050 65.700 ;
        RECT 382.950 64.950 385.050 67.050 ;
        RECT 416.400 64.050 417.450 88.950 ;
        RECT 436.950 64.950 439.050 67.050 ;
        RECT 358.950 55.950 361.050 58.050 ;
        RECT 359.400 49.050 360.450 55.950 ;
        RECT 358.950 46.950 361.050 49.050 ;
        RECT 364.950 48.600 366.150 63.600 ;
        RECT 415.950 61.950 418.050 64.050 ;
        RECT 379.950 58.950 382.050 61.050 ;
        RECT 385.950 58.950 388.050 61.050 ;
        RECT 394.950 58.950 397.050 61.050 ;
        RECT 400.950 58.950 403.050 61.050 ;
        RECT 406.950 58.950 409.050 61.050 ;
        RECT 412.950 58.950 415.050 61.050 ;
        RECT 380.400 58.200 381.600 58.950 ;
        RECT 386.400 58.200 387.600 58.950 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 379.950 55.800 382.050 57.900 ;
        RECT 382.950 55.800 385.050 57.900 ;
        RECT 385.950 55.800 388.050 57.900 ;
        RECT 388.950 55.800 391.050 57.900 ;
        RECT 368.400 54.900 369.600 55.650 ;
        RECT 367.950 52.800 370.050 54.900 ;
        RECT 383.400 53.400 384.600 55.500 ;
        RECT 389.400 54.750 390.600 55.500 ;
        RECT 364.950 46.500 367.050 48.600 ;
        RECT 355.950 40.950 358.050 43.050 ;
        RECT 367.950 40.950 370.050 43.050 ;
        RECT 334.950 37.950 337.050 40.050 ;
        RECT 364.950 37.950 367.050 40.050 ;
        RECT 325.950 32.400 328.050 34.500 ;
        RECT 311.400 13.050 312.450 20.400 ;
        RECT 319.950 19.800 322.050 21.900 ;
        RECT 325.950 17.400 327.150 32.400 ;
        RECT 328.950 26.100 331.050 28.200 ;
        RECT 340.950 26.100 343.050 31.050 ;
        RECT 329.400 25.350 330.600 26.100 ;
        RECT 341.400 25.350 342.600 26.100 ;
        RECT 365.400 25.050 366.450 37.950 ;
        RECT 328.950 22.950 331.050 25.050 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 344.400 20.400 345.600 22.650 ;
        RECT 359.400 20.400 360.600 22.650 ;
        RECT 368.400 22.050 369.450 40.950 ;
        RECT 383.400 31.050 384.450 53.400 ;
        RECT 388.950 52.650 391.050 54.750 ;
        RECT 391.950 52.950 394.050 55.050 ;
        RECT 382.950 28.950 385.050 31.050 ;
        RECT 392.400 27.600 393.450 52.950 ;
        RECT 395.400 43.050 396.450 58.950 ;
        RECT 401.400 58.200 402.600 58.950 ;
        RECT 407.400 58.200 408.600 58.950 ;
        RECT 400.950 55.800 403.050 57.900 ;
        RECT 403.950 55.800 406.050 57.900 ;
        RECT 406.950 55.800 409.050 57.900 ;
        RECT 404.400 54.000 405.600 55.500 ;
        RECT 413.400 55.050 414.450 58.950 ;
        RECT 415.950 58.800 418.050 60.900 ;
        RECT 421.950 59.100 424.050 61.200 ;
        RECT 437.400 60.600 438.450 64.950 ;
        RECT 403.950 49.950 406.050 54.000 ;
        RECT 409.950 49.950 412.050 55.050 ;
        RECT 412.950 52.950 415.050 55.050 ;
        RECT 416.400 49.050 417.450 58.800 ;
        RECT 422.400 58.350 423.600 59.100 ;
        RECT 437.400 58.350 438.600 60.600 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 424.950 55.950 427.050 58.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 446.400 57.450 447.450 91.800 ;
        RECT 449.400 61.050 450.450 118.950 ;
        RECT 455.400 105.600 456.450 121.950 ;
        RECT 461.400 115.050 462.450 137.100 ;
        RECT 463.950 130.950 466.050 133.050 ;
        RECT 464.400 127.050 465.450 130.950 ;
        RECT 463.950 124.950 466.050 127.050 ;
        RECT 469.950 126.600 471.150 141.600 ;
        RECT 478.950 139.950 481.050 142.050 ;
        RECT 485.400 138.450 486.450 163.950 ;
        RECT 482.400 137.400 486.450 138.450 ;
        RECT 490.950 138.000 493.050 142.050 ;
        RECT 497.400 139.050 498.450 176.400 ;
        RECT 503.400 166.050 504.450 176.400 ;
        RECT 508.950 175.950 511.050 178.050 ;
        RECT 515.400 177.900 516.600 178.650 ;
        RECT 502.950 163.950 505.050 166.050 ;
        RECT 509.400 145.050 510.450 175.950 ;
        RECT 514.950 175.800 517.050 177.900 ;
        RECT 518.700 168.600 519.900 188.400 ;
        RECT 529.950 181.950 532.050 184.050 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 524.400 177.450 525.600 178.650 ;
        RECT 530.400 177.450 531.450 181.950 ;
        RECT 524.400 176.400 531.450 177.450 ;
        RECT 538.950 173.400 540.150 188.400 ;
        RECT 542.400 183.450 543.600 183.600 ;
        RECT 545.400 183.450 546.450 190.950 ;
        RECT 542.400 182.400 546.450 183.450 ;
        RECT 542.400 181.350 543.600 182.400 ;
        RECT 541.950 178.950 544.050 181.050 ;
        RECT 548.400 175.050 549.450 208.950 ;
        RECT 554.400 208.050 555.450 209.400 ;
        RECT 559.950 208.650 562.050 210.750 ;
        RECT 553.950 205.950 556.050 208.050 ;
        RECT 554.400 202.050 555.450 205.950 ;
        RECT 572.700 204.600 573.900 224.400 ;
        RECT 577.950 215.100 580.050 217.200 ;
        RECT 581.400 216.450 582.450 244.950 ;
        RECT 584.400 241.050 585.450 254.400 ;
        RECT 589.950 253.950 592.050 256.050 ;
        RECT 602.400 255.000 603.600 256.650 ;
        RECT 601.950 250.950 604.050 255.000 ;
        RECT 608.400 254.400 609.600 256.650 ;
        RECT 608.400 247.050 609.450 254.400 ;
        RECT 601.950 244.950 604.050 247.050 ;
        RECT 607.950 244.950 610.050 247.050 ;
        RECT 583.950 238.950 586.050 241.050 ;
        RECT 586.950 229.950 589.050 232.050 ;
        RECT 581.400 215.400 585.450 216.450 ;
        RECT 578.400 214.350 579.600 215.100 ;
        RECT 577.950 211.950 580.050 214.050 ;
        RECT 571.950 202.500 574.050 204.600 ;
        RECT 553.950 199.950 556.050 202.050 ;
        RECT 559.950 199.950 562.050 202.050 ;
        RECT 553.950 190.950 556.050 193.050 ;
        RECT 554.400 183.600 555.450 190.950 ;
        RECT 560.400 184.200 561.450 199.950 ;
        RECT 568.950 190.950 571.050 193.050 ;
        RECT 577.950 190.950 580.050 193.050 ;
        RECT 554.400 181.350 555.600 183.600 ;
        RECT 559.950 182.100 562.050 184.200 ;
        RECT 560.400 181.350 561.600 182.100 ;
        RECT 553.950 178.950 556.050 181.050 ;
        RECT 556.950 178.950 559.050 181.050 ;
        RECT 559.950 178.950 562.050 181.050 ;
        RECT 557.400 176.400 558.600 178.650 ;
        RECT 569.400 178.050 570.450 190.950 ;
        RECT 578.400 184.200 579.450 190.950 ;
        RECT 577.950 182.100 580.050 184.200 ;
        RECT 574.950 179.100 577.050 181.200 ;
        RECT 538.950 171.300 541.050 173.400 ;
        RECT 547.950 172.950 550.050 175.050 ;
        RECT 553.950 172.950 556.050 175.050 ;
        RECT 517.950 166.500 520.050 168.600 ;
        RECT 538.950 167.700 540.150 171.300 ;
        RECT 538.950 165.600 541.050 167.700 ;
        RECT 511.950 154.950 514.050 157.050 ;
        RECT 532.950 154.950 535.050 157.050 ;
        RECT 508.950 142.950 511.050 145.050 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 473.400 132.000 474.600 133.650 ;
        RECT 472.950 127.950 475.050 132.000 ;
        RECT 460.950 112.950 463.050 115.050 ;
        RECT 461.400 105.600 462.450 112.950 ;
        RECT 464.400 109.050 465.450 124.950 ;
        RECT 469.950 124.500 472.050 126.600 ;
        RECT 478.950 118.950 481.050 121.050 ;
        RECT 469.950 110.400 472.050 112.500 ;
        RECT 463.950 106.950 466.050 109.050 ;
        RECT 455.400 103.350 456.600 105.600 ;
        RECT 461.400 103.350 462.600 105.600 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 457.950 100.950 460.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 458.400 99.900 459.600 100.650 ;
        RECT 457.950 97.800 460.050 99.900 ;
        RECT 467.400 99.000 468.600 100.650 ;
        RECT 454.950 96.450 457.050 97.050 ;
        RECT 460.950 96.450 463.050 97.050 ;
        RECT 454.950 95.400 463.050 96.450 ;
        RECT 454.950 94.950 457.050 95.400 ;
        RECT 460.950 94.950 463.050 95.400 ;
        RECT 466.950 94.950 469.050 99.000 ;
        RECT 470.700 90.600 471.900 110.400 ;
        RECT 479.400 106.050 480.450 118.950 ;
        RECT 478.950 103.950 481.050 106.050 ;
        RECT 475.950 100.950 478.050 103.050 ;
        RECT 476.400 99.900 477.600 100.650 ;
        RECT 482.400 99.900 483.450 137.400 ;
        RECT 491.400 136.350 492.600 138.000 ;
        RECT 496.950 136.950 499.050 139.050 ;
        RECT 505.950 138.000 508.050 142.050 ;
        RECT 512.400 138.600 513.450 154.950 ;
        RECT 517.950 148.950 520.050 151.050 ;
        RECT 518.400 139.050 519.450 148.950 ;
        RECT 523.950 146.400 526.050 148.500 ;
        RECT 533.400 148.050 534.450 154.950 ;
        RECT 520.950 142.950 523.050 145.050 ;
        RECT 506.400 136.350 507.600 138.000 ;
        RECT 512.400 136.350 513.600 138.600 ;
        RECT 517.950 136.950 520.050 139.050 ;
        RECT 521.400 138.600 522.450 142.950 ;
        RECT 521.400 136.350 522.600 138.600 ;
        RECT 487.950 133.950 490.050 136.050 ;
        RECT 490.950 133.950 493.050 136.050 ;
        RECT 493.950 133.950 496.050 136.050 ;
        RECT 502.950 133.950 505.050 136.050 ;
        RECT 505.950 133.950 508.050 136.050 ;
        RECT 508.950 133.950 511.050 136.050 ;
        RECT 511.950 133.950 514.050 136.050 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 484.950 130.950 487.050 133.050 ;
        RECT 488.400 131.400 489.600 133.650 ;
        RECT 494.400 132.000 495.600 133.650 ;
        RECT 503.400 132.900 504.600 133.650 ;
        RECT 475.950 97.800 478.050 99.900 ;
        RECT 481.950 97.800 484.050 99.900 ;
        RECT 469.950 88.500 472.050 90.600 ;
        RECT 463.950 79.950 466.050 82.050 ;
        RECT 457.950 64.950 460.050 67.050 ;
        RECT 448.950 58.950 451.050 61.050 ;
        RECT 458.400 60.600 459.450 64.950 ;
        RECT 464.400 60.600 465.450 79.950 ;
        RECT 485.400 73.050 486.450 130.950 ;
        RECT 488.400 127.050 489.450 131.400 ;
        RECT 493.950 127.950 496.050 132.000 ;
        RECT 502.950 130.800 505.050 132.900 ;
        RECT 509.400 132.000 510.600 133.650 ;
        RECT 508.950 127.950 511.050 132.000 ;
        RECT 517.950 130.950 520.050 133.050 ;
        RECT 514.950 127.950 517.050 130.050 ;
        RECT 487.950 124.950 490.050 127.050 ;
        RECT 494.400 118.050 495.450 127.950 ;
        RECT 493.950 115.950 496.050 118.050 ;
        RECT 490.950 110.400 493.050 112.500 ;
        RECT 505.950 110.400 508.050 112.500 ;
        RECT 490.950 95.400 492.150 110.400 ;
        RECT 493.950 105.000 496.050 109.050 ;
        RECT 494.400 103.350 495.600 105.000 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 503.400 99.900 504.600 100.650 ;
        RECT 502.950 97.800 505.050 99.900 ;
        RECT 490.950 93.300 493.050 95.400 ;
        RECT 490.950 89.700 492.150 93.300 ;
        RECT 506.700 90.600 507.900 110.400 ;
        RECT 515.400 106.050 516.450 127.950 ;
        RECT 514.950 103.950 517.050 106.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 512.400 99.000 513.600 100.650 ;
        RECT 511.950 94.950 514.050 99.000 ;
        RECT 514.950 97.950 517.050 100.050 ;
        RECT 515.400 94.050 516.450 97.950 ;
        RECT 514.950 91.950 517.050 94.050 ;
        RECT 490.950 87.600 493.050 89.700 ;
        RECT 505.950 88.500 508.050 90.600 ;
        RECT 511.950 82.950 514.050 85.050 ;
        RECT 487.950 79.950 490.050 82.050 ;
        RECT 493.950 79.950 496.050 82.050 ;
        RECT 484.950 70.950 487.050 73.050 ;
        RECT 478.950 67.950 481.050 70.050 ;
        RECT 479.400 61.200 480.450 67.950 ;
        RECT 458.400 58.200 459.600 60.600 ;
        RECT 464.400 58.200 465.600 60.600 ;
        RECT 478.950 59.100 481.050 61.200 ;
        RECT 479.400 58.350 480.600 59.100 ;
        RECT 446.400 56.400 450.450 57.450 ;
        RECT 425.400 54.900 426.600 55.650 ;
        RECT 424.950 49.950 427.050 54.900 ;
        RECT 434.400 54.000 435.600 55.650 ;
        RECT 433.950 49.950 436.050 54.000 ;
        RECT 440.400 53.400 441.600 55.650 ;
        RECT 415.950 46.950 418.050 49.050 ;
        RECT 394.950 40.950 397.050 43.050 ;
        RECT 406.950 40.950 409.050 43.050 ;
        RECT 403.950 34.950 406.050 37.050 ;
        RECT 392.400 25.350 393.600 27.600 ;
        RECT 397.950 26.100 400.050 28.200 ;
        RECT 398.400 25.350 399.600 26.100 ;
        RECT 373.950 22.950 376.050 25.050 ;
        RECT 376.950 22.950 379.050 25.050 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 391.950 22.950 394.050 25.050 ;
        RECT 394.950 22.950 397.050 25.050 ;
        RECT 397.950 22.950 400.050 25.050 ;
        RECT 325.950 15.300 328.050 17.400 ;
        RECT 344.400 16.050 345.450 20.400 ;
        RECT 304.950 10.500 307.050 12.600 ;
        RECT 310.950 10.950 313.050 13.050 ;
        RECT 325.950 11.700 327.150 15.300 ;
        RECT 343.950 13.950 346.050 16.050 ;
        RECT 325.950 9.600 328.050 11.700 ;
        RECT 359.400 10.050 360.450 20.400 ;
        RECT 367.950 19.950 370.050 22.050 ;
        RECT 374.400 21.900 375.600 22.650 ;
        RECT 373.950 19.800 376.050 21.900 ;
        RECT 389.400 20.400 390.600 22.650 ;
        RECT 395.400 21.900 396.600 22.650 ;
        RECT 404.400 21.900 405.450 34.950 ;
        RECT 407.400 28.050 408.450 40.950 ;
        RECT 412.950 34.950 415.050 37.050 ;
        RECT 406.950 25.950 409.050 28.050 ;
        RECT 413.400 27.600 414.450 34.950 ;
        RECT 416.400 28.050 417.450 46.950 ;
        RECT 440.400 43.050 441.450 53.400 ;
        RECT 445.950 52.650 448.050 54.750 ;
        RECT 449.400 54.450 450.450 56.400 ;
        RECT 454.950 55.800 457.050 57.900 ;
        RECT 457.950 55.800 460.050 57.900 ;
        RECT 460.950 55.800 463.050 57.900 ;
        RECT 463.950 55.800 466.050 57.900 ;
        RECT 466.950 55.800 469.050 57.900 ;
        RECT 475.950 55.950 478.050 58.050 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 455.400 54.750 456.600 55.500 ;
        RECT 449.400 53.400 453.450 54.450 ;
        RECT 442.950 43.950 445.050 49.050 ;
        RECT 439.950 40.950 442.050 43.050 ;
        RECT 446.400 42.450 447.450 52.650 ;
        RECT 448.950 43.950 451.050 49.050 ;
        RECT 446.400 41.400 450.450 42.450 ;
        RECT 427.950 31.950 430.050 34.050 ;
        RECT 442.950 32.400 445.050 34.500 ;
        RECT 449.400 34.050 450.450 41.400 ;
        RECT 413.400 25.350 414.600 27.600 ;
        RECT 415.950 25.950 418.050 28.050 ;
        RECT 421.950 26.100 424.050 28.200 ;
        RECT 428.400 27.600 429.450 31.950 ;
        RECT 422.400 25.350 423.600 26.100 ;
        RECT 428.400 25.350 429.600 27.600 ;
        RECT 409.950 22.950 412.050 25.050 ;
        RECT 412.950 22.950 415.050 25.050 ;
        RECT 421.950 22.950 424.050 25.050 ;
        RECT 424.950 22.950 427.050 25.050 ;
        RECT 427.950 22.950 430.050 25.050 ;
        RECT 430.950 22.950 433.050 25.050 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 410.400 22.050 411.600 22.650 ;
        RECT 389.400 16.050 390.450 20.400 ;
        RECT 394.950 19.800 397.050 21.900 ;
        RECT 403.950 19.800 406.050 21.900 ;
        RECT 406.950 20.400 411.600 22.050 ;
        RECT 425.400 21.000 426.600 22.650 ;
        RECT 431.400 21.900 432.600 22.650 ;
        RECT 440.400 21.900 441.600 22.650 ;
        RECT 406.950 19.950 411.000 20.400 ;
        RECT 424.950 16.950 427.050 21.000 ;
        RECT 430.950 19.800 433.050 21.900 ;
        RECT 439.950 19.800 442.050 21.900 ;
        RECT 361.950 13.950 367.050 16.050 ;
        RECT 370.950 13.950 376.050 16.050 ;
        RECT 388.950 13.950 391.050 16.050 ;
        RECT 358.950 7.950 361.050 10.050 ;
        RECT 431.400 7.050 432.450 19.800 ;
        RECT 443.700 12.600 444.900 32.400 ;
        RECT 448.950 31.950 451.050 34.050 ;
        RECT 452.400 28.050 453.450 53.400 ;
        RECT 454.950 52.650 457.050 54.750 ;
        RECT 461.400 53.400 462.600 55.500 ;
        RECT 467.400 54.750 468.600 55.500 ;
        RECT 461.400 43.050 462.450 53.400 ;
        RECT 466.950 52.650 469.050 54.750 ;
        RECT 476.400 53.400 477.600 55.650 ;
        RECT 472.950 46.950 475.050 49.050 ;
        RECT 454.950 40.950 457.050 43.050 ;
        RECT 460.950 40.950 463.050 43.050 ;
        RECT 451.950 25.950 454.050 28.050 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 449.400 21.450 450.600 22.650 ;
        RECT 455.400 21.450 456.450 40.950 ;
        RECT 457.950 37.950 460.050 40.050 ;
        RECT 449.400 20.400 456.450 21.450 ;
        RECT 442.950 10.500 445.050 12.600 ;
        RECT 458.400 7.050 459.450 37.950 ;
        RECT 463.950 32.400 466.050 34.500 ;
        RECT 463.950 17.400 465.150 32.400 ;
        RECT 466.950 27.000 469.050 31.050 ;
        RECT 467.400 25.350 468.600 27.000 ;
        RECT 466.950 22.950 469.050 25.050 ;
        RECT 463.950 15.300 466.050 17.400 ;
        RECT 463.950 11.700 465.150 15.300 ;
        RECT 473.400 13.050 474.450 46.950 ;
        RECT 476.400 31.050 477.450 53.400 ;
        RECT 485.400 31.050 486.450 70.950 ;
        RECT 488.400 40.050 489.450 79.950 ;
        RECT 494.400 73.050 495.450 79.950 ;
        RECT 493.950 70.950 496.050 73.050 ;
        RECT 494.400 60.600 495.450 70.950 ;
        RECT 494.400 58.350 495.600 60.600 ;
        RECT 505.950 58.950 508.050 61.050 ;
        RECT 512.400 60.600 513.450 82.950 ;
        RECT 518.400 61.050 519.450 130.950 ;
        RECT 524.700 126.600 525.900 146.400 ;
        RECT 532.950 145.950 535.050 148.050 ;
        RECT 544.950 147.300 547.050 149.400 ;
        RECT 529.950 144.450 532.050 145.050 ;
        RECT 535.950 144.450 538.050 145.050 ;
        RECT 529.950 143.400 538.050 144.450 ;
        RECT 529.950 142.950 532.050 143.400 ;
        RECT 535.950 142.950 538.050 143.400 ;
        RECT 544.950 143.700 546.150 147.300 ;
        RECT 544.950 141.600 547.050 143.700 ;
        RECT 550.950 142.950 553.050 145.050 ;
        RECT 529.950 137.100 532.050 139.200 ;
        RECT 535.950 137.100 538.050 139.200 ;
        RECT 530.400 136.350 531.600 137.100 ;
        RECT 529.950 133.950 532.050 136.050 ;
        RECT 523.950 124.500 526.050 126.600 ;
        RECT 520.950 115.950 523.050 118.050 ;
        RECT 521.400 97.050 522.450 115.950 ;
        RECT 526.950 110.400 529.050 112.500 ;
        RECT 520.950 94.950 523.050 97.050 ;
        RECT 526.950 95.400 528.150 110.400 ;
        RECT 536.400 106.200 537.450 137.100 ;
        RECT 544.950 126.600 546.150 141.600 ;
        RECT 551.400 139.050 552.450 142.950 ;
        RECT 550.950 136.950 553.050 139.050 ;
        RECT 547.950 133.950 550.050 136.050 ;
        RECT 548.400 132.900 549.600 133.650 ;
        RECT 547.950 127.950 550.050 132.900 ;
        RECT 544.950 124.500 547.050 126.600 ;
        RECT 547.950 118.950 550.050 121.050 ;
        RECT 544.950 112.950 547.050 115.050 ;
        RECT 529.950 104.100 532.050 106.200 ;
        RECT 535.950 104.100 538.050 106.200 ;
        RECT 545.400 105.600 546.450 112.950 ;
        RECT 548.400 109.050 549.450 118.950 ;
        RECT 547.950 106.950 550.050 109.050 ;
        RECT 530.400 103.350 531.600 104.100 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 536.400 100.050 537.450 104.100 ;
        RECT 545.400 103.500 546.600 105.600 ;
        RECT 550.950 104.250 553.050 106.350 ;
        RECT 554.400 106.050 555.450 172.950 ;
        RECT 557.400 166.050 558.450 176.400 ;
        RECT 568.950 175.950 571.050 178.050 ;
        RECT 556.950 163.950 559.050 166.050 ;
        RECT 562.950 148.950 565.050 151.050 ;
        RECT 563.400 138.600 564.450 148.950 ;
        RECT 584.400 145.050 585.450 215.400 ;
        RECT 587.400 151.050 588.450 229.950 ;
        RECT 592.950 225.300 595.050 227.400 ;
        RECT 592.950 221.700 594.150 225.300 ;
        RECT 592.950 219.600 595.050 221.700 ;
        RECT 592.950 204.600 594.150 219.600 ;
        RECT 595.950 211.950 598.050 214.050 ;
        RECT 596.400 210.900 597.600 211.650 ;
        RECT 595.950 208.800 598.050 210.900 ;
        RECT 592.950 202.500 595.050 204.600 ;
        RECT 589.950 196.950 592.050 199.050 ;
        RECT 586.950 148.950 589.050 151.050 ;
        RECT 583.950 142.950 586.050 145.050 ;
        RECT 585.000 141.450 589.050 142.050 ;
        RECT 584.400 139.950 589.050 141.450 ;
        RECT 563.400 136.350 564.600 138.600 ;
        RECT 568.950 137.100 571.050 139.200 ;
        RECT 584.400 138.600 585.450 139.950 ;
        RECT 590.400 139.050 591.450 196.950 ;
        RECT 602.400 184.050 603.450 244.950 ;
        RECT 614.400 229.050 615.450 313.950 ;
        RECT 626.400 298.050 627.450 349.950 ;
        RECT 631.950 344.400 634.050 346.500 ;
        RECT 631.950 329.400 633.150 344.400 ;
        RECT 644.400 343.050 645.450 376.950 ;
        RECT 647.400 372.450 648.450 394.950 ;
        RECT 650.400 376.050 651.450 409.950 ;
        RECT 665.100 402.600 666.300 422.400 ;
        RECT 667.950 412.950 670.050 415.050 ;
        RECT 668.400 411.450 669.600 412.650 ;
        RECT 668.400 410.400 672.450 411.450 ;
        RECT 664.950 400.500 667.050 402.600 ;
        RECT 671.400 388.050 672.450 410.400 ;
        RECT 674.400 400.050 675.450 475.950 ;
        RECT 689.400 469.050 690.450 526.950 ;
        RECT 692.400 523.050 693.450 527.100 ;
        RECT 698.400 526.350 699.600 527.100 ;
        RECT 704.400 526.350 705.600 528.000 ;
        RECT 719.400 526.200 720.600 528.000 ;
        RECT 724.950 526.950 727.050 529.050 ;
        RECT 725.400 526.200 726.600 526.950 ;
        RECT 697.950 523.950 700.050 526.050 ;
        RECT 700.950 523.950 703.050 526.050 ;
        RECT 703.950 523.950 706.050 526.050 ;
        RECT 706.950 523.950 709.050 526.050 ;
        RECT 715.950 523.800 718.050 525.900 ;
        RECT 718.950 523.800 721.050 525.900 ;
        RECT 721.950 523.800 724.050 525.900 ;
        RECT 724.950 523.800 727.050 525.900 ;
        RECT 727.950 523.800 730.050 525.900 ;
        RECT 691.950 520.950 694.050 523.050 ;
        RECT 701.400 521.400 702.600 523.650 ;
        RECT 707.400 522.900 708.600 523.650 ;
        RECT 693.000 519.900 697.050 520.050 ;
        RECT 691.950 517.950 697.050 519.900 ;
        RECT 691.950 517.800 694.050 517.950 ;
        RECT 701.400 517.050 702.450 521.400 ;
        RECT 706.950 520.800 709.050 522.900 ;
        RECT 716.400 522.750 717.600 523.500 ;
        RECT 715.950 520.650 718.050 522.750 ;
        RECT 722.400 521.400 723.600 523.500 ;
        RECT 728.400 522.750 729.600 523.500 ;
        RECT 700.950 514.950 703.050 517.050 ;
        RECT 722.400 511.050 723.450 521.400 ;
        RECT 727.950 520.650 730.050 522.750 ;
        RECT 730.950 520.950 733.050 523.050 ;
        RECT 694.950 508.950 697.050 511.050 ;
        RECT 721.950 508.950 724.050 511.050 ;
        RECT 691.950 494.100 694.050 496.200 ;
        RECT 695.400 496.050 696.450 508.950 ;
        RECT 697.950 505.950 700.050 508.050 ;
        RECT 715.950 505.950 718.050 508.050 ;
        RECT 692.400 487.050 693.450 494.100 ;
        RECT 694.950 493.950 697.050 496.050 ;
        RECT 698.400 495.600 699.450 505.950 ;
        RECT 712.950 502.950 715.050 505.050 ;
        RECT 709.950 496.950 712.050 499.050 ;
        RECT 698.400 493.350 699.600 495.600 ;
        RECT 703.950 494.100 706.050 496.200 ;
        RECT 704.400 493.350 705.600 494.100 ;
        RECT 697.950 490.950 700.050 493.050 ;
        RECT 700.950 490.950 703.050 493.050 ;
        RECT 703.950 490.950 706.050 493.050 ;
        RECT 701.400 488.400 702.600 490.650 ;
        RECT 691.950 484.950 694.050 487.050 ;
        RECT 688.950 466.950 691.050 469.050 ;
        RECT 701.400 466.050 702.450 488.400 ;
        RECT 679.950 463.950 682.050 466.050 ;
        RECT 700.950 463.950 703.050 466.050 ;
        RECT 680.400 451.200 681.450 463.950 ;
        RECT 694.950 454.950 697.050 457.050 ;
        RECT 679.950 449.100 682.050 451.200 ;
        RECT 685.950 449.100 688.050 451.200 ;
        RECT 680.400 448.350 681.600 449.100 ;
        RECT 686.400 448.350 687.600 449.100 ;
        RECT 679.950 445.950 682.050 448.050 ;
        RECT 682.950 445.950 685.050 448.050 ;
        RECT 685.950 445.950 688.050 448.050 ;
        RECT 688.950 445.950 691.050 448.050 ;
        RECT 683.400 443.400 684.600 445.650 ;
        RECT 689.400 444.900 690.600 445.650 ;
        RECT 695.400 445.050 696.450 454.950 ;
        RECT 710.400 454.050 711.450 496.950 ;
        RECT 713.400 496.050 714.450 502.950 ;
        RECT 712.950 493.950 715.050 496.050 ;
        RECT 716.400 495.600 717.450 505.950 ;
        RECT 721.950 499.050 724.050 499.350 ;
        RECT 731.400 499.050 732.450 520.950 ;
        RECT 718.950 497.250 724.050 499.050 ;
        RECT 718.950 496.950 723.000 497.250 ;
        RECT 730.950 496.950 733.050 499.050 ;
        RECT 734.400 496.200 735.450 544.950 ;
        RECT 749.400 544.050 750.450 556.950 ;
        RECT 757.950 550.950 760.050 553.050 ;
        RECT 748.950 541.950 751.050 544.050 ;
        RECT 736.950 535.950 739.050 538.050 ;
        RECT 737.400 529.050 738.450 535.950 ;
        RECT 742.800 531.300 744.900 533.400 ;
        RECT 752.400 532.500 754.500 534.600 ;
        RECT 736.950 526.950 739.050 529.050 ;
        RECT 740.400 526.050 741.600 528.600 ;
        RECT 739.950 523.800 742.050 526.050 ;
        RECT 743.700 522.300 744.600 531.300 ;
        RECT 745.950 527.700 748.050 529.800 ;
        RECT 749.400 528.900 750.600 531.600 ;
        RECT 747.150 525.300 748.050 527.700 ;
        RECT 748.950 526.800 751.050 528.900 ;
        RECT 752.850 525.300 754.050 532.500 ;
        RECT 758.400 529.050 759.450 550.950 ;
        RECT 757.950 526.950 760.050 529.050 ;
        RECT 760.950 526.950 763.050 529.050 ;
        RECT 769.950 528.000 772.050 532.050 ;
        RECT 773.400 529.050 774.450 574.950 ;
        RECT 757.050 525.900 760.050 526.050 ;
        RECT 747.150 524.100 754.050 525.300 ;
        RECT 750.150 522.300 752.250 523.200 ;
        RECT 743.700 521.100 752.250 522.300 ;
        RECT 745.200 519.300 747.300 521.100 ;
        RECT 748.950 518.100 751.050 520.200 ;
        RECT 753.150 518.700 754.050 524.100 ;
        RECT 754.950 523.950 760.050 525.900 ;
        RECT 754.950 523.800 757.050 523.950 ;
        RECT 755.400 521.400 756.600 523.800 ;
        RECT 761.400 520.050 762.450 526.950 ;
        RECT 770.400 526.350 771.600 528.000 ;
        RECT 772.950 526.950 775.050 529.050 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 769.950 523.950 772.050 526.050 ;
        RECT 767.400 522.900 768.600 523.650 ;
        RECT 766.950 520.800 769.050 522.900 ;
        RECT 749.400 515.400 750.600 518.100 ;
        RECT 752.400 516.600 754.500 518.700 ;
        RECT 760.950 517.950 763.050 520.050 ;
        RECT 742.950 508.950 745.050 511.050 ;
        RECT 739.950 502.950 742.050 505.050 ;
        RECT 716.400 493.500 717.600 495.600 ;
        RECT 721.950 494.100 724.050 496.200 ;
        RECT 733.950 494.100 736.050 496.200 ;
        RECT 740.400 495.600 741.450 502.950 ;
        RECT 743.400 496.050 744.450 508.950 ;
        RECT 761.400 508.050 762.450 517.950 ;
        RECT 745.950 505.950 748.050 508.050 ;
        RECT 760.950 505.950 763.050 508.050 ;
        RECT 722.400 493.500 723.600 494.100 ;
        RECT 734.400 493.350 735.600 494.100 ;
        RECT 740.400 493.350 741.600 495.600 ;
        RECT 742.950 493.950 745.050 496.050 ;
        RECT 715.950 491.100 718.050 493.200 ;
        RECT 718.950 491.100 721.050 493.200 ;
        RECT 721.950 491.100 724.050 493.200 ;
        RECT 724.950 491.100 727.050 493.200 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 739.950 490.950 742.050 493.050 ;
        RECT 719.400 488.400 720.600 490.800 ;
        RECT 725.400 490.050 726.600 490.800 ;
        RECT 719.400 469.050 720.450 488.400 ;
        RECT 724.950 487.950 727.050 490.050 ;
        RECT 737.400 489.000 738.600 490.650 ;
        RECT 736.950 484.950 739.050 489.000 ;
        RECT 742.950 487.950 745.050 490.050 ;
        RECT 739.950 484.950 742.050 487.050 ;
        RECT 740.400 469.050 741.450 484.950 ;
        RECT 743.400 484.050 744.450 487.950 ;
        RECT 742.950 481.950 745.050 484.050 ;
        RECT 718.950 466.950 721.050 469.050 ;
        RECT 739.950 466.950 742.050 469.050 ;
        RECT 703.950 450.000 706.050 454.050 ;
        RECT 709.950 451.950 712.050 454.050 ;
        RECT 719.400 451.050 720.450 466.950 ;
        RECT 740.400 454.050 741.450 466.950 ;
        RECT 746.400 463.050 747.450 505.950 ;
        RECT 748.950 496.950 751.050 502.050 ;
        RECT 761.400 498.900 762.600 501.600 ;
        RECT 757.200 495.900 759.300 497.700 ;
        RECT 760.950 496.800 763.050 498.900 ;
        RECT 764.400 498.300 766.500 500.400 ;
        RECT 755.700 494.700 764.250 495.900 ;
        RECT 751.950 491.100 754.050 493.200 ;
        RECT 752.400 489.450 753.600 491.100 ;
        RECT 749.400 488.400 753.600 489.450 ;
        RECT 749.400 472.050 750.450 488.400 ;
        RECT 755.700 485.700 756.600 494.700 ;
        RECT 762.150 493.800 764.250 494.700 ;
        RECT 765.150 492.900 766.050 498.300 ;
        RECT 767.400 493.200 768.600 495.600 ;
        RECT 772.950 493.950 775.050 496.050 ;
        RECT 776.400 495.450 777.450 577.950 ;
        RECT 782.400 577.050 783.450 599.400 ;
        RECT 781.950 574.950 784.050 577.050 ;
        RECT 791.400 576.450 792.450 613.950 ;
        RECT 796.950 606.000 799.050 610.050 ;
        RECT 803.400 606.600 804.450 625.950 ;
        RECT 806.400 613.050 807.450 643.950 ;
        RECT 809.400 640.050 810.450 644.400 ;
        RECT 811.950 643.950 814.050 646.050 ;
        RECT 817.950 643.950 820.050 646.050 ;
        RECT 824.400 644.400 825.600 646.800 ;
        RECT 808.950 637.950 811.050 640.050 ;
        RECT 805.950 610.950 808.050 613.050 ;
        RECT 812.400 610.050 813.450 643.950 ;
        RECT 824.400 637.050 825.450 644.400 ;
        RECT 823.950 634.950 826.050 637.050 ;
        RECT 833.400 622.050 834.450 652.950 ;
        RECT 836.400 652.050 837.450 658.950 ;
        RECT 835.950 649.950 838.050 652.050 ;
        RECT 842.400 651.600 843.450 661.950 ;
        RECT 854.400 654.450 855.450 682.950 ;
        RECT 857.400 678.750 858.450 718.950 ;
        RECT 856.950 676.650 859.050 678.750 ;
        RECT 854.400 653.400 858.450 654.450 ;
        RECT 842.400 649.500 843.600 651.600 ;
        RECT 847.950 650.250 850.050 652.350 ;
        RECT 848.400 649.500 849.600 650.250 ;
        RECT 853.950 649.950 856.050 652.050 ;
        RECT 838.950 647.100 841.050 649.200 ;
        RECT 841.950 647.100 844.050 649.200 ;
        RECT 844.950 647.100 847.050 649.200 ;
        RECT 847.950 647.100 850.050 649.200 ;
        RECT 839.400 644.400 840.600 646.800 ;
        RECT 845.400 646.050 846.600 646.800 ;
        RECT 839.400 640.050 840.450 644.400 ;
        RECT 841.800 643.950 843.900 646.050 ;
        RECT 844.950 643.950 847.050 646.050 ;
        RECT 838.950 637.950 841.050 640.050 ;
        RECT 838.950 625.950 841.050 628.050 ;
        RECT 832.950 619.950 835.050 622.050 ;
        RECT 823.950 610.950 826.050 613.050 ;
        RECT 811.950 607.950 814.050 610.050 ;
        RECT 797.400 604.200 798.600 606.000 ;
        RECT 803.400 604.200 804.600 606.600 ;
        RECT 796.950 601.800 799.050 603.900 ;
        RECT 799.950 601.800 802.050 603.900 ;
        RECT 802.950 601.800 805.050 603.900 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 817.950 601.950 820.050 604.050 ;
        RECT 793.950 598.950 796.050 601.050 ;
        RECT 800.400 600.750 801.600 601.500 ;
        RECT 788.400 575.400 792.450 576.450 ;
        RECT 788.400 574.200 789.450 575.400 ;
        RECT 787.950 572.100 790.050 574.200 ;
        RECT 794.400 574.050 795.450 598.950 ;
        RECT 799.950 598.650 802.050 600.750 ;
        RECT 812.400 599.400 813.600 601.650 ;
        RECT 812.400 595.050 813.450 599.400 ;
        RECT 820.950 598.950 823.050 601.050 ;
        RECT 817.950 595.950 820.050 598.050 ;
        RECT 811.950 592.950 814.050 595.050 ;
        RECT 802.950 577.950 805.050 580.050 ;
        RECT 788.400 571.350 789.600 572.100 ;
        RECT 793.950 571.950 796.050 574.050 ;
        RECT 803.400 573.600 804.450 577.950 ;
        RECT 811.950 574.950 814.050 577.050 ;
        RECT 803.400 571.500 804.600 573.600 ;
        RECT 781.950 568.950 784.050 571.050 ;
        RECT 787.950 568.950 790.050 571.050 ;
        RECT 790.950 568.950 793.050 571.050 ;
        RECT 799.950 569.100 802.050 571.200 ;
        RECT 802.950 569.100 805.050 571.200 ;
        RECT 805.950 569.100 808.050 571.200 ;
        RECT 782.400 566.400 783.600 568.650 ;
        RECT 782.400 538.050 783.450 566.400 ;
        RECT 784.950 565.950 787.050 568.050 ;
        RECT 791.400 566.400 792.600 568.650 ;
        RECT 800.400 566.400 801.600 568.800 ;
        RECT 806.400 568.050 807.600 568.800 ;
        RECT 781.950 535.950 784.050 538.050 ;
        RECT 782.400 528.450 783.600 528.600 ;
        RECT 785.400 528.450 786.450 565.950 ;
        RECT 791.400 562.050 792.450 566.400 ;
        RECT 787.950 559.950 790.050 562.050 ;
        RECT 790.950 559.950 793.050 562.050 ;
        RECT 782.400 527.400 786.450 528.450 ;
        RECT 788.400 528.600 789.450 559.950 ;
        RECT 800.400 559.050 801.450 566.400 ;
        RECT 805.950 565.950 808.050 568.050 ;
        RECT 806.400 562.050 807.450 565.950 ;
        RECT 805.950 559.950 808.050 562.050 ;
        RECT 799.950 556.950 802.050 559.050 ;
        RECT 782.400 526.200 783.600 527.400 ;
        RECT 788.400 526.200 789.600 528.600 ;
        RECT 793.950 526.950 796.050 529.050 ;
        RECT 802.950 527.100 805.050 529.200 ;
        RECT 812.400 528.450 813.450 574.950 ;
        RECT 818.400 573.600 819.450 595.950 ;
        RECT 821.400 574.050 822.450 598.950 ;
        RECT 824.400 577.050 825.450 610.950 ;
        RECT 832.950 605.100 835.050 607.200 ;
        RECT 839.400 607.050 840.450 625.950 ;
        RECT 833.400 604.350 834.600 605.100 ;
        RECT 838.950 604.950 841.050 607.050 ;
        RECT 829.950 601.950 832.050 604.050 ;
        RECT 832.950 601.950 835.050 604.050 ;
        RECT 835.950 601.950 838.050 604.050 ;
        RECT 830.400 599.400 831.600 601.650 ;
        RECT 836.400 599.400 837.600 601.650 ;
        RECT 830.400 586.050 831.450 599.400 ;
        RECT 832.950 595.950 835.050 598.050 ;
        RECT 829.950 583.950 832.050 586.050 ;
        RECT 829.950 577.950 832.050 580.050 ;
        RECT 823.950 574.950 826.050 577.050 ;
        RECT 818.400 571.350 819.600 573.600 ;
        RECT 820.950 571.950 823.050 574.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 823.950 568.950 826.050 571.050 ;
        RECT 820.950 565.950 823.050 568.050 ;
        RECT 821.400 544.050 822.450 565.950 ;
        RECT 820.950 541.950 823.050 544.050 ;
        RECT 830.400 538.050 831.450 577.950 ;
        RECT 833.400 574.050 834.450 595.950 ;
        RECT 836.400 595.050 837.450 599.400 ;
        RECT 838.950 598.950 841.050 601.050 ;
        RECT 835.950 592.950 838.050 595.050 ;
        RECT 832.950 571.950 835.050 574.050 ;
        RECT 839.400 573.450 840.450 598.950 ;
        RECT 842.400 580.050 843.450 643.950 ;
        RECT 854.400 628.050 855.450 649.950 ;
        RECT 853.950 625.950 856.050 628.050 ;
        RECT 857.400 610.050 858.450 653.400 ;
        RECT 860.400 646.050 861.450 721.950 ;
        RECT 859.950 643.950 862.050 646.050 ;
        RECT 863.400 642.450 864.450 766.950 ;
        RECT 860.400 641.400 864.450 642.450 ;
        RECT 856.950 607.950 859.050 610.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 853.950 601.950 856.050 604.050 ;
        RECT 848.400 599.400 849.600 601.650 ;
        RECT 848.400 592.050 849.450 599.400 ;
        RECT 853.950 592.950 856.050 595.050 ;
        RECT 847.950 589.950 850.050 592.050 ;
        RECT 841.950 577.950 844.050 580.050 ;
        RECT 841.950 573.450 844.050 574.350 ;
        RECT 839.400 572.400 844.050 573.450 ;
        RECT 841.950 572.250 844.050 572.400 ;
        RECT 842.400 571.500 843.600 572.250 ;
        RECT 850.950 571.950 853.050 574.050 ;
        RECT 835.950 569.100 838.050 571.200 ;
        RECT 841.950 569.100 844.050 571.200 ;
        RECT 844.950 569.100 847.050 571.200 ;
        RECT 832.950 565.950 835.050 568.050 ;
        RECT 836.400 566.400 837.600 568.800 ;
        RECT 845.400 566.400 846.600 568.800 ;
        RECT 829.950 535.950 832.050 538.050 ;
        RECT 817.800 531.300 819.900 533.400 ;
        RECT 827.400 532.500 829.500 534.600 ;
        RECT 809.400 527.400 813.450 528.450 ;
        RECT 781.950 523.800 784.050 525.900 ;
        RECT 784.950 523.800 787.050 525.900 ;
        RECT 787.950 523.800 790.050 525.900 ;
        RECT 785.400 521.400 786.600 523.500 ;
        RECT 785.400 502.050 786.450 521.400 ;
        RECT 784.950 499.950 787.050 502.050 ;
        RECT 779.400 495.450 780.600 495.600 ;
        RECT 776.400 494.400 780.600 495.450 ;
        RECT 759.150 491.700 766.050 492.900 ;
        RECT 759.150 489.300 760.050 491.700 ;
        RECT 757.950 487.200 760.050 489.300 ;
        RECT 760.950 488.100 763.050 490.200 ;
        RECT 754.800 483.600 756.900 485.700 ;
        RECT 761.400 485.400 762.600 488.100 ;
        RECT 764.850 484.500 766.050 491.700 ;
        RECT 766.950 491.100 769.050 493.200 ;
        RECT 773.400 490.050 774.450 493.950 ;
        RECT 779.400 493.350 780.600 494.400 ;
        RECT 784.950 494.100 787.050 496.200 ;
        RECT 794.400 495.450 795.450 526.950 ;
        RECT 803.400 526.350 804.600 527.100 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 800.400 522.000 801.600 523.650 ;
        RECT 799.950 517.950 802.050 522.000 ;
        RECT 805.950 520.950 808.050 523.050 ;
        RECT 806.400 505.050 807.450 520.950 ;
        RECT 809.400 514.050 810.450 527.400 ;
        RECT 815.400 526.050 816.600 528.600 ;
        RECT 814.950 523.800 817.050 526.050 ;
        RECT 818.700 522.300 819.600 531.300 ;
        RECT 820.950 527.700 823.050 529.800 ;
        RECT 824.400 528.900 825.600 531.600 ;
        RECT 822.150 525.300 823.050 527.700 ;
        RECT 823.950 526.800 826.050 528.900 ;
        RECT 827.850 525.300 829.050 532.500 ;
        RECT 833.400 529.050 834.450 565.950 ;
        RECT 836.400 562.050 837.450 566.400 ;
        RECT 835.950 559.950 838.050 562.050 ;
        RECT 838.950 547.950 841.050 550.050 ;
        RECT 835.950 535.950 838.050 538.050 ;
        RECT 832.950 526.950 835.050 529.050 ;
        RECT 822.150 524.100 829.050 525.300 ;
        RECT 825.150 522.300 827.250 523.200 ;
        RECT 818.700 521.100 827.250 522.300 ;
        RECT 811.950 517.950 814.050 520.050 ;
        RECT 820.200 519.300 822.300 521.100 ;
        RECT 823.950 518.100 826.050 520.200 ;
        RECT 828.150 518.700 829.050 524.100 ;
        RECT 829.950 523.800 832.050 525.900 ;
        RECT 830.400 521.400 831.600 523.800 ;
        RECT 808.950 511.950 811.050 514.050 ;
        RECT 805.950 502.950 808.050 505.050 ;
        RECT 791.400 494.400 795.450 495.450 ;
        RECT 785.400 493.350 786.600 494.100 ;
        RECT 778.950 490.950 781.050 493.050 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 772.950 487.950 775.050 490.050 ;
        RECT 782.400 488.400 783.600 490.650 ;
        RECT 764.400 482.400 766.500 484.500 ;
        RECT 778.950 478.950 781.050 481.050 ;
        RECT 760.950 472.950 763.050 478.050 ;
        RECT 748.950 469.950 751.050 472.050 ;
        RECT 745.950 460.950 748.050 463.050 ;
        RECT 766.950 460.950 769.050 463.050 ;
        RECT 704.400 448.200 705.600 450.000 ;
        RECT 709.950 448.800 712.050 450.900 ;
        RECT 718.950 450.450 721.050 451.050 ;
        RECT 716.400 449.400 721.050 450.450 ;
        RECT 721.950 450.000 724.050 454.050 ;
        RECT 727.950 450.000 730.050 454.050 ;
        RECT 739.950 451.950 742.050 454.050 ;
        RECT 710.400 448.200 711.600 448.800 ;
        RECT 700.950 445.800 703.050 447.900 ;
        RECT 703.950 445.800 706.050 447.900 ;
        RECT 706.950 445.800 709.050 447.900 ;
        RECT 709.950 445.800 712.050 447.900 ;
        RECT 683.400 433.050 684.450 443.400 ;
        RECT 688.950 442.800 691.050 444.900 ;
        RECT 694.950 442.950 697.050 445.050 ;
        RECT 701.400 444.750 702.600 445.500 ;
        RECT 700.950 442.650 703.050 444.750 ;
        RECT 707.400 443.400 708.600 445.500 ;
        RECT 685.950 439.950 688.050 442.050 ;
        RECT 686.400 436.050 687.450 439.950 ;
        RECT 707.400 439.050 708.450 443.400 ;
        RECT 706.950 436.950 709.050 439.050 ;
        RECT 716.400 438.450 717.450 449.400 ;
        RECT 718.950 448.950 721.050 449.400 ;
        RECT 722.400 448.200 723.600 450.000 ;
        RECT 728.400 448.200 729.600 450.000 ;
        RECT 739.950 448.800 742.050 450.900 ;
        RECT 745.950 450.000 748.050 454.050 ;
        RECT 759.000 453.450 763.050 454.050 ;
        RECT 758.400 451.950 763.050 453.450 ;
        RECT 763.950 451.950 766.050 454.050 ;
        RECT 758.400 450.600 759.450 451.950 ;
        RECT 740.400 448.200 741.600 448.800 ;
        RECT 746.400 448.200 747.600 450.000 ;
        RECT 758.400 448.350 759.600 450.600 ;
        RECT 721.950 445.800 724.050 447.900 ;
        RECT 724.950 445.800 727.050 447.900 ;
        RECT 727.950 445.800 730.050 447.900 ;
        RECT 739.950 445.800 742.050 447.900 ;
        RECT 742.950 445.800 745.050 447.900 ;
        RECT 745.950 445.800 748.050 447.900 ;
        RECT 754.950 445.950 757.050 448.050 ;
        RECT 757.950 445.950 760.050 448.050 ;
        RECT 725.400 444.750 726.600 445.500 ;
        RECT 724.950 442.650 727.050 444.750 ;
        RECT 730.950 442.950 733.050 445.050 ;
        RECT 736.950 442.950 739.050 445.050 ;
        RECT 743.400 443.400 744.600 445.500 ;
        RECT 755.400 444.900 756.600 445.650 ;
        RECT 764.400 445.050 765.450 451.950 ;
        RECT 716.400 437.400 720.450 438.450 ;
        RECT 685.950 433.950 688.050 436.050 ;
        RECT 715.950 433.950 718.050 436.050 ;
        RECT 682.950 430.950 685.050 433.050 ;
        RECT 703.950 421.950 706.050 424.050 ;
        RECT 682.950 416.250 685.050 418.350 ;
        RECT 683.400 415.500 684.600 416.250 ;
        RECT 691.950 415.950 694.050 418.050 ;
        RECT 697.950 416.100 700.050 418.200 ;
        RECT 704.400 417.600 705.450 421.950 ;
        RECT 679.950 413.100 682.050 415.200 ;
        RECT 682.950 413.100 685.050 415.200 ;
        RECT 685.950 413.100 688.050 415.200 ;
        RECT 680.400 412.050 681.600 412.800 ;
        RECT 686.400 412.050 687.600 412.800 ;
        RECT 679.950 409.950 682.050 412.050 ;
        RECT 685.950 409.950 688.050 412.050 ;
        RECT 673.950 397.950 676.050 400.050 ;
        RECT 686.400 388.050 687.450 409.950 ;
        RECT 692.400 406.050 693.450 415.950 ;
        RECT 698.400 415.350 699.600 416.100 ;
        RECT 704.400 415.350 705.600 417.600 ;
        RECT 712.950 415.950 715.050 418.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 700.950 412.950 703.050 415.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 706.950 412.950 709.050 415.050 ;
        RECT 701.400 410.400 702.600 412.650 ;
        RECT 707.400 410.400 708.600 412.650 ;
        RECT 691.950 403.950 694.050 406.050 ;
        RECT 701.400 400.050 702.450 410.400 ;
        RECT 707.400 406.050 708.450 410.400 ;
        RECT 706.950 403.950 709.050 406.050 ;
        RECT 713.400 400.050 714.450 415.950 ;
        RECT 716.400 406.050 717.450 433.950 ;
        RECT 719.400 418.050 720.450 437.400 ;
        RECT 718.950 415.950 721.050 418.050 ;
        RECT 724.950 416.100 727.050 418.200 ;
        RECT 731.400 417.600 732.450 442.950 ;
        RECT 737.400 436.050 738.450 442.950 ;
        RECT 736.950 433.950 739.050 436.050 ;
        RECT 743.400 421.050 744.450 443.400 ;
        RECT 754.950 442.800 757.050 444.900 ;
        RECT 763.950 442.950 766.050 445.050 ;
        RECT 767.400 439.050 768.450 460.950 ;
        RECT 772.950 450.000 775.050 454.050 ;
        RECT 779.400 450.600 780.450 478.950 ;
        RECT 782.400 454.050 783.450 488.400 ;
        RECT 791.400 478.050 792.450 494.400 ;
        RECT 799.950 494.250 802.050 496.350 ;
        RECT 800.400 493.500 801.600 494.250 ;
        RECT 796.950 491.100 799.050 493.200 ;
        RECT 799.950 491.100 802.050 493.200 ;
        RECT 802.950 491.100 805.050 493.200 ;
        RECT 797.400 489.450 798.600 490.800 ;
        RECT 803.400 490.050 804.600 490.800 ;
        RECT 809.400 490.050 810.450 511.950 ;
        RECT 812.400 496.050 813.450 517.950 ;
        RECT 824.400 515.400 825.600 518.100 ;
        RECT 827.400 516.600 829.500 518.700 ;
        RECT 817.950 511.950 820.050 514.050 ;
        RECT 811.950 493.950 814.050 496.050 ;
        RECT 818.400 495.600 819.450 511.950 ;
        RECT 824.400 498.450 825.450 515.400 ;
        RECT 824.400 498.000 828.450 498.450 ;
        RECT 824.400 497.400 829.050 498.000 ;
        RECT 818.400 493.500 819.600 495.600 ;
        RECT 823.950 494.250 826.050 496.350 ;
        RECT 824.400 493.500 825.600 494.250 ;
        RECT 826.950 493.950 829.050 497.400 ;
        RECT 829.950 496.950 832.050 499.050 ;
        RECT 814.950 491.100 817.050 493.200 ;
        RECT 817.950 491.100 820.050 493.200 ;
        RECT 820.950 491.100 823.050 493.200 ;
        RECT 823.950 491.100 826.050 493.200 ;
        RECT 797.400 488.400 801.450 489.450 ;
        RECT 800.400 481.050 801.450 488.400 ;
        RECT 802.950 487.950 805.050 490.050 ;
        RECT 805.950 487.950 808.050 490.050 ;
        RECT 808.950 487.950 811.050 490.050 ;
        RECT 815.400 488.400 816.600 490.800 ;
        RECT 821.400 489.000 822.600 490.800 ;
        RECT 799.950 478.950 802.050 481.050 ;
        RECT 790.950 475.950 793.050 478.050 ;
        RECT 796.950 475.950 799.050 478.050 ;
        RECT 790.950 469.950 793.050 472.050 ;
        RECT 781.950 451.950 784.050 454.050 ;
        RECT 791.400 450.600 792.450 469.950 ;
        RECT 797.400 451.050 798.450 475.950 ;
        RECT 773.400 448.350 774.600 450.000 ;
        RECT 779.400 448.350 780.600 450.600 ;
        RECT 791.400 448.200 792.600 450.600 ;
        RECT 796.950 448.950 799.050 451.050 ;
        RECT 797.400 448.200 798.600 448.950 ;
        RECT 772.950 445.950 775.050 448.050 ;
        RECT 775.950 445.950 778.050 448.050 ;
        RECT 778.950 445.950 781.050 448.050 ;
        RECT 781.950 445.950 784.050 448.050 ;
        RECT 790.950 445.800 793.050 447.900 ;
        RECT 793.950 445.800 796.050 447.900 ;
        RECT 796.950 445.800 799.050 447.900 ;
        RECT 799.950 445.800 802.050 447.900 ;
        RECT 776.400 443.400 777.600 445.650 ;
        RECT 782.400 444.900 783.600 445.650 ;
        RECT 766.950 436.950 769.050 439.050 ;
        RECT 772.950 436.950 775.050 439.050 ;
        RECT 766.950 424.950 769.050 427.050 ;
        RECT 742.950 418.950 745.050 421.050 ;
        RECT 725.400 415.350 726.600 416.100 ;
        RECT 731.400 415.350 732.600 417.600 ;
        RECT 736.950 415.950 739.050 418.050 ;
        RECT 745.950 416.250 748.050 418.350 ;
        RECT 760.950 417.000 763.050 421.050 ;
        RECT 767.400 417.600 768.450 424.950 ;
        RECT 721.950 412.950 724.050 415.050 ;
        RECT 724.950 412.950 727.050 415.050 ;
        RECT 727.950 412.950 730.050 415.050 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 722.400 412.050 723.600 412.650 ;
        RECT 718.950 411.900 723.600 412.050 ;
        RECT 718.950 409.950 724.050 411.900 ;
        RECT 721.950 409.800 724.050 409.950 ;
        RECT 728.400 410.400 729.600 412.650 ;
        RECT 718.950 406.800 721.050 408.900 ;
        RECT 715.950 403.950 718.050 406.050 ;
        RECT 700.950 397.950 703.050 400.050 ;
        RECT 712.950 397.950 715.050 400.050 ;
        RECT 664.950 385.950 667.050 388.050 ;
        RECT 670.950 385.950 673.050 388.050 ;
        RECT 685.950 385.950 688.050 388.050 ;
        RECT 661.950 382.950 664.050 385.050 ;
        RECT 655.950 376.950 658.050 379.050 ;
        RECT 649.950 373.950 652.050 376.050 ;
        RECT 656.400 372.600 657.450 376.950 ;
        RECT 662.400 372.600 663.450 382.950 ;
        RECT 665.400 379.050 666.450 385.950 ;
        RECT 682.950 382.950 685.050 385.050 ;
        RECT 670.950 380.400 673.050 382.500 ;
        RECT 664.950 376.950 667.050 379.050 ;
        RECT 650.400 372.450 651.600 372.600 ;
        RECT 647.400 371.400 651.600 372.450 ;
        RECT 650.400 370.200 651.600 371.400 ;
        RECT 656.400 370.200 657.600 372.600 ;
        RECT 662.400 370.200 663.600 372.600 ;
        RECT 665.400 372.450 666.450 376.950 ;
        RECT 668.400 372.450 669.600 372.600 ;
        RECT 665.400 371.400 669.600 372.450 ;
        RECT 668.400 370.350 669.600 371.400 ;
        RECT 649.950 367.800 652.050 369.900 ;
        RECT 652.950 367.800 655.050 369.900 ;
        RECT 655.950 367.800 658.050 369.900 ;
        RECT 658.950 367.800 661.050 369.900 ;
        RECT 661.950 367.800 664.050 369.900 ;
        RECT 667.950 367.950 670.050 370.050 ;
        RECT 653.400 366.750 654.600 367.500 ;
        RECT 652.950 364.650 655.050 366.750 ;
        RECT 659.400 365.400 660.600 367.500 ;
        RECT 659.400 361.050 660.450 365.400 ;
        RECT 664.950 364.950 667.050 367.050 ;
        RECT 658.950 358.950 661.050 361.050 ;
        RECT 634.950 339.000 637.050 343.050 ;
        RECT 640.950 340.950 643.050 343.050 ;
        RECT 643.950 340.950 646.050 343.050 ;
        RECT 665.400 342.450 666.450 364.950 ;
        RECT 671.700 360.600 672.900 380.400 ;
        RECT 676.950 371.100 679.050 373.200 ;
        RECT 677.400 370.350 678.600 371.100 ;
        RECT 676.950 367.950 679.050 370.050 ;
        RECT 683.400 366.450 684.450 382.950 ;
        RECT 680.400 365.400 684.450 366.450 ;
        RECT 670.950 358.500 673.050 360.600 ;
        RECT 665.400 341.400 669.450 342.450 ;
        RECT 635.400 337.350 636.600 339.000 ;
        RECT 634.950 334.950 637.050 337.050 ;
        RECT 631.950 327.300 634.050 329.400 ;
        RECT 631.950 323.700 633.150 327.300 ;
        RECT 641.400 325.050 642.450 340.950 ;
        RECT 643.950 337.800 646.050 339.900 ;
        RECT 652.950 338.250 655.050 340.350 ;
        RECT 668.400 340.200 669.450 341.400 ;
        RECT 631.950 321.600 634.050 323.700 ;
        RECT 640.950 322.950 643.050 325.050 ;
        RECT 644.400 319.050 645.450 337.800 ;
        RECT 653.400 337.500 654.600 338.250 ;
        RECT 667.950 338.100 670.050 340.200 ;
        RECT 668.400 337.350 669.600 338.100 ;
        RECT 649.950 335.100 652.050 337.200 ;
        RECT 652.950 335.100 655.050 337.200 ;
        RECT 655.950 335.100 658.050 337.200 ;
        RECT 664.950 334.950 667.050 337.050 ;
        RECT 667.950 334.950 670.050 337.050 ;
        RECT 673.950 334.950 676.050 337.050 ;
        RECT 650.400 334.050 651.600 334.800 ;
        RECT 656.400 334.050 657.600 334.800 ;
        RECT 646.950 331.950 649.050 334.050 ;
        RECT 649.950 331.950 652.050 334.050 ;
        RECT 655.950 331.950 658.050 334.050 ;
        RECT 665.400 333.900 666.600 334.650 ;
        RECT 674.400 333.900 675.600 334.650 ;
        RECT 643.950 316.950 646.050 319.050 ;
        RECT 634.950 302.400 637.050 304.500 ;
        RECT 647.400 304.050 648.450 331.950 ;
        RECT 656.400 325.050 657.450 331.950 ;
        RECT 664.950 331.800 667.050 333.900 ;
        RECT 673.950 331.800 676.050 333.900 ;
        RECT 680.400 328.050 681.450 365.400 ;
        RECT 686.400 361.050 687.450 385.950 ;
        RECT 691.950 381.300 694.050 383.400 ;
        RECT 691.950 377.700 693.150 381.300 ;
        RECT 706.950 380.400 709.050 382.500 ;
        RECT 691.950 375.600 694.050 377.700 ;
        RECT 703.950 376.950 706.050 379.050 ;
        RECT 685.950 358.950 688.050 361.050 ;
        RECT 691.950 360.600 693.150 375.600 ;
        RECT 704.400 372.600 705.450 376.950 ;
        RECT 704.400 370.350 705.600 372.600 ;
        RECT 694.950 367.950 697.050 370.050 ;
        RECT 703.950 367.950 706.050 370.050 ;
        RECT 695.400 366.450 696.600 367.650 ;
        RECT 695.400 365.400 699.450 366.450 ;
        RECT 691.950 358.500 694.050 360.600 ;
        RECT 698.400 343.050 699.450 365.400 ;
        RECT 707.700 360.600 708.900 380.400 ;
        RECT 712.950 371.100 715.050 373.200 ;
        RECT 713.400 370.350 714.600 371.100 ;
        RECT 712.950 367.950 715.050 370.050 ;
        RECT 709.950 363.450 712.050 367.050 ;
        RECT 709.950 363.000 714.450 363.450 ;
        RECT 710.400 362.400 714.450 363.000 ;
        RECT 706.950 358.500 709.050 360.600 ;
        RECT 697.950 340.950 700.050 343.050 ;
        RECT 691.950 338.250 694.050 340.350 ;
        RECT 713.400 339.600 714.450 362.400 ;
        RECT 719.400 339.600 720.450 406.800 ;
        RECT 728.400 406.050 729.450 410.400 ;
        RECT 727.950 403.950 730.050 406.050 ;
        RECT 737.400 397.050 738.450 415.950 ;
        RECT 746.400 415.500 747.600 416.250 ;
        RECT 761.400 415.500 762.600 417.000 ;
        RECT 767.400 415.500 768.600 417.600 ;
        RECT 742.950 413.100 745.050 415.200 ;
        RECT 745.950 413.100 748.050 415.200 ;
        RECT 748.950 413.100 751.050 415.200 ;
        RECT 757.950 413.100 760.050 415.200 ;
        RECT 760.950 413.100 763.050 415.200 ;
        RECT 763.950 413.100 766.050 415.200 ;
        RECT 766.950 413.100 769.050 415.200 ;
        RECT 743.400 410.400 744.600 412.800 ;
        RECT 749.400 410.400 750.600 412.800 ;
        RECT 743.400 403.050 744.450 410.400 ;
        RECT 749.400 406.050 750.450 410.400 ;
        RECT 754.950 409.950 757.050 412.050 ;
        RECT 758.400 411.000 759.600 412.800 ;
        RECT 764.400 412.050 765.600 412.800 ;
        RECT 748.950 403.950 751.050 406.050 ;
        RECT 742.950 400.950 745.050 403.050 ;
        RECT 755.400 400.050 756.450 409.950 ;
        RECT 757.950 408.450 760.050 411.000 ;
        RECT 763.950 409.950 766.050 412.050 ;
        RECT 757.950 407.400 762.450 408.450 ;
        RECT 757.950 406.950 760.050 407.400 ;
        RECT 754.950 397.950 757.050 400.050 ;
        RECT 736.950 394.950 739.050 397.050 ;
        RECT 727.950 381.300 730.050 383.400 ;
        RECT 727.950 377.700 729.150 381.300 ;
        RECT 727.950 375.600 730.050 377.700 ;
        RECT 721.950 371.100 724.050 373.200 ;
        RECT 722.400 361.050 723.450 371.100 ;
        RECT 721.950 358.950 724.050 361.050 ;
        RECT 727.950 360.600 729.150 375.600 ;
        RECT 739.950 370.950 742.050 373.050 ;
        RECT 745.950 371.100 748.050 373.200 ;
        RECT 761.400 372.600 762.450 407.400 ;
        RECT 769.950 406.950 772.050 412.050 ;
        RECT 773.400 406.050 774.450 436.950 ;
        RECT 776.400 418.050 777.450 443.400 ;
        RECT 781.950 442.800 784.050 444.900 ;
        RECT 794.400 443.400 795.600 445.500 ;
        RECT 800.400 443.400 801.600 445.500 ;
        RECT 784.950 439.950 787.050 442.050 ;
        RECT 794.400 441.450 795.450 443.400 ;
        RECT 791.400 441.000 795.450 441.450 ;
        RECT 790.950 440.400 795.450 441.000 ;
        RECT 781.950 430.950 784.050 433.050 ;
        RECT 775.950 415.950 778.050 418.050 ;
        RECT 782.400 417.600 783.450 430.950 ;
        RECT 785.400 430.050 786.450 439.950 ;
        RECT 790.950 439.050 793.050 440.400 ;
        RECT 790.800 438.000 793.050 439.050 ;
        RECT 790.800 436.950 792.900 438.000 ;
        RECT 793.950 436.950 796.050 439.050 ;
        RECT 784.950 427.950 787.050 430.050 ;
        RECT 790.950 424.950 793.050 427.050 ;
        RECT 782.400 415.500 783.600 417.600 ;
        RECT 787.950 417.000 790.050 421.050 ;
        RECT 791.400 418.050 792.450 424.950 ;
        RECT 788.400 415.500 789.600 417.000 ;
        RECT 790.950 415.950 793.050 418.050 ;
        RECT 778.950 413.100 781.050 415.200 ;
        RECT 781.950 413.100 784.050 415.200 ;
        RECT 784.950 413.100 787.050 415.200 ;
        RECT 787.950 413.100 790.050 415.200 ;
        RECT 775.950 409.950 778.050 412.050 ;
        RECT 779.400 410.400 780.600 412.800 ;
        RECT 785.400 411.000 786.600 412.800 ;
        RECT 776.400 406.050 777.450 409.950 ;
        RECT 772.800 403.950 774.900 406.050 ;
        RECT 775.950 403.950 778.050 406.050 ;
        RECT 779.400 400.050 780.450 410.400 ;
        RECT 784.950 406.950 787.050 411.000 ;
        RECT 787.950 409.950 790.050 412.050 ;
        RECT 778.950 397.950 781.050 400.050 ;
        RECT 766.950 379.950 769.050 382.050 ;
        RECT 778.950 380.400 781.050 382.500 ;
        RECT 788.400 382.050 789.450 409.950 ;
        RECT 767.400 372.600 768.450 379.950 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 731.400 366.000 732.600 367.650 ;
        RECT 740.400 366.900 741.450 370.950 ;
        RECT 746.400 370.350 747.600 371.100 ;
        RECT 761.400 370.350 762.600 372.600 ;
        RECT 767.400 370.350 768.600 372.600 ;
        RECT 775.950 372.000 778.050 376.050 ;
        RECT 776.400 370.350 777.600 372.000 ;
        RECT 745.950 367.950 748.050 370.050 ;
        RECT 748.950 367.950 751.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 763.950 367.950 766.050 370.050 ;
        RECT 766.950 367.950 769.050 370.050 ;
        RECT 775.950 367.950 778.050 370.050 ;
        RECT 730.950 361.950 733.050 366.000 ;
        RECT 739.950 364.800 742.050 366.900 ;
        RECT 749.400 366.000 750.600 367.650 ;
        RECT 758.400 366.900 759.600 367.650 ;
        RECT 748.950 361.950 751.050 366.000 ;
        RECT 757.950 364.800 760.050 366.900 ;
        RECT 764.400 365.400 765.600 367.650 ;
        RECT 727.950 358.500 730.050 360.600 ;
        RECT 749.400 349.050 750.450 361.950 ;
        RECT 748.950 346.950 751.050 349.050 ;
        RECT 754.950 343.950 757.050 346.050 ;
        RECT 692.400 337.500 693.600 338.250 ;
        RECT 713.400 337.350 714.600 339.600 ;
        RECT 719.400 337.350 720.600 339.600 ;
        RECT 724.950 337.950 727.050 340.050 ;
        RECT 733.950 339.000 736.050 343.050 ;
        RECT 685.950 335.100 688.050 337.200 ;
        RECT 691.950 335.100 694.050 337.200 ;
        RECT 694.950 335.100 697.050 337.200 ;
        RECT 700.950 334.950 703.050 337.050 ;
        RECT 709.950 334.950 712.050 337.050 ;
        RECT 712.950 334.950 715.050 337.050 ;
        RECT 715.950 334.950 718.050 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 686.400 334.050 687.600 334.800 ;
        RECT 685.950 331.950 688.050 334.050 ;
        RECT 695.400 332.400 696.600 334.800 ;
        RECT 664.950 325.950 667.050 328.050 ;
        RECT 679.950 325.950 682.050 328.050 ;
        RECT 655.950 322.950 658.050 325.050 ;
        RECT 625.950 295.950 628.050 298.050 ;
        RECT 619.950 293.100 622.050 295.200 ;
        RECT 631.950 294.000 634.050 298.050 ;
        RECT 620.400 292.350 621.600 293.100 ;
        RECT 632.400 292.350 633.600 294.000 ;
        RECT 619.950 289.950 622.050 292.050 ;
        RECT 625.950 289.950 628.050 292.050 ;
        RECT 631.950 289.950 634.050 292.050 ;
        RECT 626.400 287.400 627.600 289.650 ;
        RECT 626.400 274.050 627.450 287.400 ;
        RECT 635.700 282.600 636.900 302.400 ;
        RECT 640.950 301.950 643.050 304.050 ;
        RECT 646.950 301.950 649.050 304.050 ;
        RECT 655.950 303.300 658.050 305.400 ;
        RECT 641.400 294.600 642.450 301.950 ;
        RECT 655.950 299.700 657.150 303.300 ;
        RECT 646.950 295.950 649.050 298.050 ;
        RECT 655.950 297.600 658.050 299.700 ;
        RECT 641.400 292.350 642.600 294.600 ;
        RECT 640.950 289.950 643.050 292.050 ;
        RECT 634.950 280.500 637.050 282.600 ;
        RECT 625.950 271.950 628.050 274.050 ;
        RECT 634.950 266.400 637.050 268.500 ;
        RECT 616.950 260.100 619.050 262.200 ;
        RECT 625.950 260.100 628.050 262.200 ;
        RECT 617.400 250.050 618.450 260.100 ;
        RECT 626.400 259.350 627.600 260.100 ;
        RECT 622.950 256.950 625.050 259.050 ;
        RECT 625.950 256.950 628.050 259.050 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 623.400 255.900 624.600 256.650 ;
        RECT 632.400 255.900 633.600 256.650 ;
        RECT 622.950 253.800 625.050 255.900 ;
        RECT 631.950 253.800 634.050 255.900 ;
        RECT 616.950 247.950 619.050 250.050 ;
        RECT 635.700 246.600 636.900 266.400 ;
        RECT 640.950 256.950 643.050 259.050 ;
        RECT 641.400 254.400 642.600 256.650 ;
        RECT 647.400 255.900 648.450 295.950 ;
        RECT 655.950 282.600 657.150 297.600 ;
        RECT 658.950 289.950 661.050 292.050 ;
        RECT 659.400 288.450 660.600 289.650 ;
        RECT 659.400 287.400 663.450 288.450 ;
        RECT 662.400 283.050 663.450 287.400 ;
        RECT 655.950 280.500 658.050 282.600 ;
        RECT 661.950 280.950 664.050 283.050 ;
        RECT 661.950 277.800 664.050 279.900 ;
        RECT 649.950 271.950 652.050 274.050 ;
        RECT 641.400 250.050 642.450 254.400 ;
        RECT 646.950 253.800 649.050 255.900 ;
        RECT 640.950 247.950 643.050 250.050 ;
        RECT 634.950 244.500 637.050 246.600 ;
        RECT 650.400 235.050 651.450 271.950 ;
        RECT 655.950 266.400 658.050 268.500 ;
        RECT 655.950 251.400 657.150 266.400 ;
        RECT 658.950 261.450 661.050 262.200 ;
        RECT 662.400 261.450 663.450 277.800 ;
        RECT 658.950 260.400 663.450 261.450 ;
        RECT 658.950 260.100 661.050 260.400 ;
        RECT 659.400 259.350 660.600 260.100 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 655.950 249.300 658.050 251.400 ;
        RECT 665.400 250.050 666.450 325.950 ;
        RECT 679.950 304.950 682.050 310.050 ;
        RECT 691.950 301.950 694.050 304.050 ;
        RECT 676.500 298.500 678.600 300.600 ;
        RECT 670.950 292.950 673.050 298.050 ;
        RECT 673.950 289.800 676.050 291.900 ;
        RECT 676.950 291.300 678.150 298.500 ;
        RECT 680.400 294.900 681.600 297.600 ;
        RECT 686.100 297.300 688.200 299.400 ;
        RECT 679.950 292.800 682.050 294.900 ;
        RECT 682.950 293.700 685.050 295.800 ;
        RECT 682.950 291.300 683.850 293.700 ;
        RECT 676.950 290.100 683.850 291.300 ;
        RECT 674.400 287.400 675.600 289.800 ;
        RECT 676.950 284.700 677.850 290.100 ;
        RECT 678.750 288.300 680.850 289.200 ;
        RECT 686.400 288.300 687.300 297.300 ;
        RECT 689.400 294.450 690.600 294.600 ;
        RECT 692.400 294.450 693.450 301.950 ;
        RECT 695.400 295.050 696.450 332.400 ;
        RECT 701.400 319.050 702.450 334.950 ;
        RECT 710.400 333.900 711.600 334.650 ;
        RECT 716.400 333.900 717.600 334.650 ;
        RECT 725.400 333.900 726.450 337.950 ;
        RECT 734.400 337.350 735.600 339.000 ;
        RECT 742.950 338.100 745.050 340.200 ;
        RECT 748.950 339.000 751.050 343.050 ;
        RECT 743.400 337.350 744.600 338.100 ;
        RECT 749.400 337.350 750.600 339.000 ;
        RECT 730.950 334.950 733.050 337.050 ;
        RECT 733.950 334.950 736.050 337.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 731.400 333.900 732.600 334.650 ;
        RECT 703.950 331.800 706.050 333.900 ;
        RECT 709.950 331.800 712.050 333.900 ;
        RECT 715.950 331.800 718.050 333.900 ;
        RECT 724.950 331.800 727.050 333.900 ;
        RECT 730.950 331.800 733.050 333.900 ;
        RECT 746.400 333.000 747.600 334.650 ;
        RECT 700.950 316.950 703.050 319.050 ;
        RECT 697.950 304.950 700.050 307.050 ;
        RECT 698.400 298.050 699.450 304.950 ;
        RECT 697.950 295.950 700.050 298.050 ;
        RECT 689.400 293.400 693.450 294.450 ;
        RECT 689.400 291.900 690.600 293.400 ;
        RECT 694.950 292.950 697.050 295.050 ;
        RECT 700.950 293.100 703.050 295.200 ;
        RECT 704.400 295.050 705.450 331.800 ;
        RECT 745.950 328.950 748.050 333.000 ;
        RECT 755.400 331.050 756.450 343.950 ;
        RECT 758.400 343.050 759.450 364.800 ;
        RECT 764.400 361.050 765.450 365.400 ;
        RECT 763.950 358.950 766.050 361.050 ;
        RECT 779.700 360.600 780.900 380.400 ;
        RECT 787.950 379.950 790.050 382.050 ;
        RECT 784.950 371.100 787.050 373.200 ;
        RECT 790.950 371.100 793.050 373.200 ;
        RECT 785.400 370.350 786.600 371.100 ;
        RECT 784.950 367.950 787.050 370.050 ;
        RECT 778.950 358.500 781.050 360.600 ;
        RECT 791.400 352.050 792.450 371.100 ;
        RECT 790.950 349.950 793.050 352.050 ;
        RECT 766.950 346.950 769.050 349.050 ;
        RECT 757.950 340.950 760.050 343.050 ;
        RECT 760.950 339.000 763.050 343.050 ;
        RECT 767.400 339.600 768.450 346.950 ;
        RECT 784.950 343.950 787.050 346.050 ;
        RECT 761.400 337.350 762.600 339.000 ;
        RECT 767.400 337.350 768.600 339.600 ;
        RECT 772.950 338.100 775.050 340.200 ;
        RECT 778.950 338.100 781.050 340.200 ;
        RECT 785.400 339.600 786.450 343.950 ;
        RECT 760.950 334.950 763.050 337.050 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 764.400 333.900 765.600 334.650 ;
        RECT 773.400 334.050 774.450 338.100 ;
        RECT 779.400 337.350 780.600 338.100 ;
        RECT 785.400 337.350 786.600 339.600 ;
        RECT 794.400 339.450 795.450 436.950 ;
        RECT 800.400 436.050 801.450 443.400 ;
        RECT 799.950 433.950 802.050 436.050 ;
        RECT 796.950 430.950 799.050 433.050 ;
        RECT 797.400 418.050 798.450 430.950 ;
        RECT 802.950 424.950 805.050 427.050 ;
        RECT 796.950 415.950 799.050 418.050 ;
        RECT 803.400 417.600 804.450 424.950 ;
        RECT 806.400 424.050 807.450 487.950 ;
        RECT 815.400 472.050 816.450 488.400 ;
        RECT 820.950 484.950 823.050 489.000 ;
        RECT 826.950 487.950 829.050 490.050 ;
        RECT 814.950 469.950 817.050 472.050 ;
        RECT 823.950 462.450 826.050 463.050 ;
        RECT 827.400 462.450 828.450 487.950 ;
        RECT 830.400 481.050 831.450 496.950 ;
        RECT 836.400 495.450 837.450 535.950 ;
        RECT 839.400 529.050 840.450 547.950 ;
        RECT 841.950 541.950 844.050 544.050 ;
        RECT 842.400 529.050 843.450 541.950 ;
        RECT 838.950 526.950 841.050 529.050 ;
        RECT 841.950 526.950 844.050 529.050 ;
        RECT 845.400 528.450 846.450 566.400 ;
        RECT 851.400 559.050 852.450 571.950 ;
        RECT 850.950 556.950 853.050 559.050 ;
        RECT 854.400 535.050 855.450 592.950 ;
        RECT 860.400 567.450 861.450 641.400 ;
        RECT 862.950 607.950 865.050 610.050 ;
        RECT 863.400 595.050 864.450 607.950 ;
        RECT 862.950 592.950 865.050 595.050 ;
        RECT 862.950 583.950 865.050 586.050 ;
        RECT 857.400 566.400 861.450 567.450 ;
        RECT 853.950 532.950 856.050 535.050 ;
        RECT 857.400 532.050 858.450 566.400 ;
        RECT 859.950 532.950 862.050 535.050 ;
        RECT 856.950 529.950 859.050 532.050 ;
        RECT 847.950 528.450 850.050 529.050 ;
        RECT 845.400 527.400 850.050 528.450 ;
        RECT 847.950 526.950 850.050 527.400 ;
        RECT 842.400 526.200 843.600 526.950 ;
        RECT 848.400 526.200 849.600 526.950 ;
        RECT 856.950 526.800 859.050 528.900 ;
        RECT 841.950 523.800 844.050 525.900 ;
        RECT 844.950 523.800 847.050 525.900 ;
        RECT 847.950 523.800 850.050 525.900 ;
        RECT 850.950 523.800 853.050 525.900 ;
        RECT 845.400 521.400 846.600 523.500 ;
        RECT 851.400 522.450 852.600 523.500 ;
        RECT 851.400 521.400 855.450 522.450 ;
        RECT 841.950 517.950 844.050 520.050 ;
        RECT 842.400 499.050 843.450 517.950 ;
        RECT 845.400 514.050 846.450 521.400 ;
        RECT 850.950 517.950 853.050 520.050 ;
        RECT 844.950 511.950 847.050 514.050 ;
        RECT 841.950 496.950 844.050 499.050 ;
        RECT 833.400 494.400 837.450 495.450 ;
        RECT 842.400 495.600 843.450 496.950 ;
        RECT 829.950 478.950 832.050 481.050 ;
        RECT 823.950 461.400 828.450 462.450 ;
        RECT 823.950 460.950 826.050 461.400 ;
        RECT 811.950 445.950 814.050 448.050 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 812.400 444.000 813.600 445.650 ;
        RECT 811.950 439.950 814.050 444.000 ;
        RECT 805.950 421.950 808.050 424.050 ;
        RECT 824.400 420.450 825.450 460.950 ;
        RECT 833.400 460.050 834.450 494.400 ;
        RECT 842.400 493.350 843.600 495.600 ;
        RECT 838.950 490.950 841.050 493.050 ;
        RECT 841.950 490.950 844.050 493.050 ;
        RECT 839.400 489.000 840.600 490.650 ;
        RECT 838.950 484.950 841.050 489.000 ;
        RECT 826.950 457.950 829.050 460.050 ;
        RECT 832.950 457.950 835.050 460.050 ;
        RECT 827.400 439.050 828.450 457.950 ;
        RECT 835.500 454.500 837.600 456.600 ;
        RECT 829.950 448.950 832.050 454.050 ;
        RECT 832.950 445.800 835.050 447.900 ;
        RECT 835.950 447.300 837.150 454.500 ;
        RECT 839.400 450.900 840.600 453.600 ;
        RECT 845.100 453.300 847.200 455.400 ;
        RECT 851.400 454.050 852.450 517.950 ;
        RECT 854.400 511.050 855.450 521.400 ;
        RECT 857.400 520.050 858.450 526.800 ;
        RECT 856.950 517.950 859.050 520.050 ;
        RECT 856.950 514.800 859.050 516.900 ;
        RECT 853.950 508.950 856.050 511.050 ;
        RECT 853.950 493.950 856.050 496.050 ;
        RECT 838.950 448.800 841.050 450.900 ;
        RECT 841.950 449.700 844.050 451.800 ;
        RECT 841.950 447.300 842.850 449.700 ;
        RECT 835.950 446.100 842.850 447.300 ;
        RECT 833.400 443.400 834.600 445.800 ;
        RECT 835.950 440.700 836.850 446.100 ;
        RECT 837.750 444.300 839.850 445.200 ;
        RECT 845.400 444.300 846.300 453.300 ;
        RECT 850.950 451.950 853.050 454.050 ;
        RECT 854.400 451.050 855.450 493.950 ;
        RECT 847.950 448.950 850.050 451.050 ;
        RECT 853.950 448.950 856.050 451.050 ;
        RECT 848.400 447.900 849.600 448.950 ;
        RECT 847.950 445.800 850.050 447.900 ;
        RECT 837.750 443.100 846.300 444.300 ;
        RECT 826.950 436.950 829.050 439.050 ;
        RECT 835.500 438.600 837.600 440.700 ;
        RECT 838.950 440.100 841.050 442.200 ;
        RECT 842.700 441.300 844.800 443.100 ;
        RECT 839.400 437.400 840.600 440.100 ;
        RECT 829.950 424.950 832.050 427.050 ;
        RECT 826.950 421.950 829.050 424.050 ;
        RECT 821.400 419.400 825.450 420.450 ;
        RECT 810.000 417.600 814.050 418.050 ;
        RECT 803.400 415.500 804.600 417.600 ;
        RECT 809.400 415.950 814.050 417.600 ;
        RECT 814.950 416.100 817.050 418.200 ;
        RECT 821.400 417.600 822.450 419.400 ;
        RECT 827.400 418.050 828.450 421.950 ;
        RECT 809.400 415.500 810.600 415.950 ;
        RECT 799.950 413.100 802.050 415.200 ;
        RECT 802.950 413.100 805.050 415.200 ;
        RECT 805.950 413.100 808.050 415.200 ;
        RECT 808.950 413.100 811.050 415.200 ;
        RECT 800.400 411.000 801.600 412.800 ;
        RECT 799.950 406.950 802.050 411.000 ;
        RECT 806.400 410.400 807.600 412.800 ;
        RECT 806.400 406.050 807.450 410.400 ;
        RECT 815.400 409.050 816.450 416.100 ;
        RECT 821.400 415.350 822.600 417.600 ;
        RECT 826.950 415.950 829.050 418.050 ;
        RECT 820.950 412.950 823.050 415.050 ;
        RECT 823.950 412.950 826.050 415.050 ;
        RECT 817.950 409.950 820.050 412.050 ;
        RECT 824.400 411.900 825.600 412.650 ;
        RECT 814.950 406.950 817.050 409.050 ;
        RECT 805.950 403.950 808.050 406.050 ;
        RECT 799.950 381.300 802.050 383.400 ;
        RECT 799.950 377.700 801.150 381.300 ;
        RECT 811.950 379.950 814.050 382.050 ;
        RECT 799.950 375.600 802.050 377.700 ;
        RECT 799.950 360.600 801.150 375.600 ;
        RECT 808.950 370.950 811.050 373.050 ;
        RECT 802.950 367.950 805.050 370.050 ;
        RECT 803.400 366.900 804.600 367.650 ;
        RECT 802.950 366.450 805.050 366.900 ;
        RECT 802.950 365.400 807.450 366.450 ;
        RECT 802.950 364.800 805.050 365.400 ;
        RECT 799.950 358.500 802.050 360.600 ;
        RECT 791.400 338.400 795.450 339.450 ;
        RECT 778.950 334.950 781.050 337.050 ;
        RECT 781.950 334.950 784.050 337.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 763.950 331.800 766.050 333.900 ;
        RECT 772.950 331.950 775.050 334.050 ;
        RECT 782.400 332.400 783.600 334.650 ;
        RECT 754.950 328.950 757.050 331.050 ;
        RECT 721.950 316.950 724.050 319.050 ;
        RECT 701.400 292.350 702.600 293.100 ;
        RECT 703.950 292.950 706.050 295.050 ;
        RECT 706.950 292.950 709.050 295.050 ;
        RECT 715.950 293.100 718.050 295.200 ;
        RECT 722.400 294.600 723.450 316.950 ;
        RECT 739.950 301.950 742.050 304.050 ;
        RECT 727.950 298.950 730.050 301.050 ;
        RECT 688.950 289.800 691.050 291.900 ;
        RECT 697.950 289.950 700.050 292.050 ;
        RECT 700.950 289.950 703.050 292.050 ;
        RECT 698.400 288.900 699.600 289.650 ;
        RECT 707.400 288.900 708.450 292.950 ;
        RECT 716.400 292.350 717.600 293.100 ;
        RECT 722.400 292.350 723.600 294.600 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 715.950 289.950 718.050 292.050 ;
        RECT 718.950 289.950 721.050 292.050 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 678.750 287.100 687.300 288.300 ;
        RECT 667.950 280.950 670.050 283.050 ;
        RECT 676.500 282.600 678.600 284.700 ;
        RECT 679.950 284.100 682.050 286.200 ;
        RECT 683.700 285.300 685.800 287.100 ;
        RECT 697.950 286.800 700.050 288.900 ;
        RECT 706.950 286.800 709.050 288.900 ;
        RECT 709.950 286.950 712.050 289.050 ;
        RECT 713.400 288.900 714.600 289.650 ;
        RECT 680.400 281.400 681.600 284.100 ;
        RECT 668.400 253.050 669.450 280.950 ;
        RECT 673.950 268.950 676.050 271.050 ;
        RECT 674.400 265.050 675.450 268.950 ;
        RECT 698.400 268.050 699.450 286.800 ;
        RECT 679.950 265.950 682.050 268.050 ;
        RECT 697.950 265.950 700.050 268.050 ;
        RECT 673.950 262.950 676.050 265.050 ;
        RECT 674.400 261.600 675.450 262.950 ;
        RECT 680.400 261.600 681.450 265.950 ;
        RECT 674.400 259.350 675.600 261.600 ;
        RECT 680.400 259.350 681.600 261.600 ;
        RECT 694.950 260.100 697.050 262.200 ;
        RECT 700.950 260.100 703.050 262.200 ;
        RECT 707.400 262.050 708.450 286.800 ;
        RECT 710.400 262.050 711.450 286.950 ;
        RECT 712.950 286.800 715.050 288.900 ;
        RECT 719.400 287.400 720.600 289.650 ;
        RECT 695.400 259.350 696.600 260.100 ;
        RECT 701.400 259.350 702.600 260.100 ;
        RECT 706.950 259.950 709.050 262.050 ;
        RECT 709.950 259.950 712.050 262.050 ;
        RECT 715.950 261.000 718.050 265.050 ;
        RECT 719.400 262.050 720.450 287.400 ;
        RECT 721.950 283.950 724.050 286.050 ;
        RECT 716.400 259.350 717.600 261.000 ;
        RECT 718.950 259.950 721.050 262.050 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 679.950 256.950 682.050 259.050 ;
        RECT 691.950 256.950 694.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 700.950 256.950 703.050 259.050 ;
        RECT 706.950 256.800 709.050 258.900 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 677.400 254.400 678.600 256.650 ;
        RECT 667.950 250.950 670.050 253.050 ;
        RECT 673.950 250.950 676.050 253.050 ;
        RECT 677.400 252.450 678.450 254.400 ;
        RECT 688.950 253.950 691.050 256.050 ;
        RECT 692.400 254.400 693.600 256.650 ;
        RECT 698.400 255.900 699.600 256.650 ;
        RECT 677.400 251.400 681.450 252.450 ;
        RECT 655.950 245.700 657.150 249.300 ;
        RECT 664.950 247.950 667.050 250.050 ;
        RECT 655.950 243.600 658.050 245.700 ;
        RECT 649.950 232.950 652.050 235.050 ;
        RECT 613.950 226.950 616.050 229.050 ;
        RECT 637.950 226.950 640.050 229.050 ;
        RECT 610.950 223.950 613.050 226.050 ;
        RECT 625.950 224.400 628.050 226.500 ;
        RECT 611.400 216.600 612.450 223.950 ;
        RECT 611.400 214.350 612.600 216.600 ;
        RECT 622.950 216.000 625.050 220.050 ;
        RECT 623.400 214.350 624.600 216.000 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 613.950 211.950 616.050 214.050 ;
        RECT 622.950 211.950 625.050 214.050 ;
        RECT 608.400 210.900 609.600 211.650 ;
        RECT 607.950 208.800 610.050 210.900 ;
        RECT 614.400 209.400 615.600 211.650 ;
        RECT 608.400 205.050 609.450 208.800 ;
        RECT 607.950 202.950 610.050 205.050 ;
        RECT 604.950 199.950 607.050 202.050 ;
        RECT 601.950 181.950 604.050 184.050 ;
        RECT 595.950 179.100 598.050 181.200 ;
        RECT 596.400 176.400 597.600 178.800 ;
        RECT 596.400 166.050 597.450 176.400 ;
        RECT 595.950 165.450 598.050 166.050 ;
        RECT 593.400 164.400 598.050 165.450 ;
        RECT 569.400 136.350 570.600 137.100 ;
        RECT 584.400 136.350 585.600 138.600 ;
        RECT 589.950 136.950 592.050 139.050 ;
        RECT 559.950 133.950 562.050 136.050 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 565.950 133.950 568.050 136.050 ;
        RECT 568.950 133.950 571.050 136.050 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 583.950 133.950 586.050 136.050 ;
        RECT 586.950 133.950 589.050 136.050 ;
        RECT 560.400 131.400 561.600 133.650 ;
        RECT 566.400 132.900 567.600 133.650 ;
        RECT 560.400 115.050 561.450 131.400 ;
        RECT 565.950 130.800 568.050 132.900 ;
        RECT 571.950 130.950 574.050 133.050 ;
        RECT 581.400 131.400 582.600 133.650 ;
        RECT 587.400 132.900 588.600 133.650 ;
        RECT 572.400 121.050 573.450 130.950 ;
        RECT 571.950 118.950 574.050 121.050 ;
        RECT 581.400 118.050 582.450 131.400 ;
        RECT 586.950 130.800 589.050 132.900 ;
        RECT 574.950 115.950 577.050 118.050 ;
        RECT 580.950 115.950 583.050 118.050 ;
        RECT 559.950 112.950 562.050 115.050 ;
        RECT 565.950 112.950 568.050 115.050 ;
        RECT 571.950 112.950 574.050 115.050 ;
        RECT 556.950 106.950 559.050 109.050 ;
        RECT 551.400 103.500 552.600 104.250 ;
        RECT 553.950 103.950 556.050 106.050 ;
        RECT 541.950 101.100 544.050 103.200 ;
        RECT 544.950 101.100 547.050 103.200 ;
        RECT 547.950 101.100 550.050 103.200 ;
        RECT 550.950 101.100 553.050 103.200 ;
        RECT 542.400 100.050 543.600 100.800 ;
        RECT 548.400 100.050 549.600 100.800 ;
        RECT 535.950 97.950 538.050 100.050 ;
        RECT 541.950 97.950 544.050 100.050 ;
        RECT 544.950 98.400 549.600 100.050 ;
        RECT 544.950 97.950 549.000 98.400 ;
        RECT 550.950 97.950 553.050 100.050 ;
        RECT 553.950 97.950 556.050 100.050 ;
        RECT 526.950 93.300 529.050 95.400 ;
        RECT 526.950 89.700 528.150 93.300 ;
        RECT 538.950 91.950 541.050 97.050 ;
        RECT 526.950 87.600 529.050 89.700 ;
        RECT 547.950 88.950 550.050 94.050 ;
        RECT 526.950 82.950 529.050 85.050 ;
        RECT 541.950 82.950 544.050 85.050 ;
        RECT 527.400 61.200 528.450 82.950 ;
        RECT 493.950 55.950 496.050 58.050 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 500.400 54.900 501.600 55.650 ;
        RECT 506.400 54.900 507.450 58.950 ;
        RECT 512.400 58.350 513.600 60.600 ;
        RECT 517.950 58.950 520.050 61.050 ;
        RECT 526.950 59.100 529.050 61.200 ;
        RECT 532.950 60.000 535.050 64.050 ;
        RECT 538.950 61.950 541.050 64.050 ;
        RECT 527.400 58.350 528.600 59.100 ;
        RECT 533.400 58.350 534.600 60.000 ;
        RECT 511.950 55.950 514.050 58.050 ;
        RECT 514.950 55.950 517.050 58.050 ;
        RECT 523.950 55.950 526.050 58.050 ;
        RECT 526.950 55.950 529.050 58.050 ;
        RECT 529.950 55.950 532.050 58.050 ;
        RECT 532.950 55.950 535.050 58.050 ;
        RECT 499.950 52.800 502.050 54.900 ;
        RECT 505.950 52.800 508.050 54.900 ;
        RECT 524.400 54.450 525.600 55.650 ;
        RECT 521.400 53.400 525.600 54.450 ;
        RECT 530.400 53.400 531.600 55.650 ;
        RECT 521.400 49.050 522.450 53.400 ;
        RECT 523.950 49.950 526.050 52.050 ;
        RECT 520.950 46.950 523.050 49.050 ;
        RECT 524.400 46.050 525.450 49.950 ;
        RECT 530.400 46.050 531.450 53.400 ;
        RECT 535.950 52.950 538.050 55.050 ;
        RECT 523.950 43.950 526.050 46.050 ;
        RECT 529.950 43.950 532.050 46.050 ;
        RECT 487.950 37.950 490.050 40.050 ;
        RECT 520.950 37.950 523.050 40.050 ;
        RECT 508.950 34.950 511.050 37.050 ;
        RECT 490.950 31.950 493.050 34.050 ;
        RECT 475.950 28.950 478.050 31.050 ;
        RECT 484.950 28.950 487.050 31.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 484.950 22.950 487.050 25.050 ;
        RECT 482.400 21.900 483.600 22.650 ;
        RECT 481.950 19.800 484.050 21.900 ;
        RECT 463.950 9.600 466.050 11.700 ;
        RECT 472.950 10.950 475.050 13.050 ;
        RECT 491.400 10.050 492.450 31.950 ;
        RECT 499.950 26.250 502.050 28.350 ;
        RECT 500.400 25.500 501.600 26.250 ;
        RECT 496.950 23.100 499.050 25.200 ;
        RECT 499.950 23.100 502.050 25.200 ;
        RECT 502.950 23.100 505.050 25.200 ;
        RECT 497.400 21.000 498.600 22.800 ;
        RECT 496.950 16.950 499.050 21.000 ;
        RECT 503.400 20.400 504.600 22.800 ;
        RECT 503.400 13.050 504.450 20.400 ;
        RECT 509.400 16.050 510.450 34.950 ;
        RECT 517.950 31.950 520.050 34.050 ;
        RECT 518.400 27.600 519.450 31.950 ;
        RECT 521.400 31.050 522.450 37.950 ;
        RECT 520.950 28.950 523.050 31.050 ;
        RECT 524.400 27.600 525.450 43.950 ;
        RECT 536.400 40.050 537.450 52.950 ;
        RECT 539.400 49.050 540.450 61.950 ;
        RECT 542.400 52.050 543.450 82.950 ;
        RECT 547.950 60.450 550.050 61.200 ;
        RECT 551.400 60.450 552.450 97.950 ;
        RECT 554.400 82.050 555.450 97.950 ;
        RECT 553.950 79.950 556.050 82.050 ;
        RECT 553.950 64.950 556.050 67.050 ;
        RECT 547.950 59.400 552.450 60.450 ;
        RECT 554.400 60.600 555.450 64.950 ;
        RECT 557.400 61.050 558.450 106.950 ;
        RECT 566.400 105.600 567.450 112.950 ;
        RECT 566.400 103.500 567.600 105.600 ;
        RECT 562.950 101.100 565.050 103.200 ;
        RECT 565.950 101.100 568.050 103.200 ;
        RECT 563.400 100.050 564.600 100.800 ;
        RECT 572.400 100.050 573.450 112.950 ;
        RECT 575.400 106.050 576.450 115.950 ;
        RECT 593.400 109.050 594.450 164.400 ;
        RECT 595.950 163.950 598.050 164.400 ;
        RECT 605.400 151.050 606.450 199.950 ;
        RECT 614.400 193.050 615.450 209.400 ;
        RECT 626.700 204.600 627.900 224.400 ;
        RECT 631.950 215.100 634.050 217.200 ;
        RECT 632.400 214.350 633.600 215.100 ;
        RECT 631.950 211.950 634.050 214.050 ;
        RECT 634.950 208.950 637.050 211.050 ;
        RECT 625.950 202.500 628.050 204.600 ;
        RECT 613.950 190.950 616.050 193.050 ;
        RECT 628.950 190.950 631.050 193.050 ;
        RECT 629.400 184.350 630.450 190.950 ;
        RECT 613.950 182.250 616.050 184.350 ;
        RECT 628.950 182.250 631.050 184.350 ;
        RECT 635.400 183.600 636.450 208.950 ;
        RECT 638.400 202.050 639.450 226.950 ;
        RECT 646.950 225.300 649.050 227.400 ;
        RECT 646.950 221.700 648.150 225.300 ;
        RECT 667.950 223.950 670.050 226.050 ;
        RECT 646.950 219.600 649.050 221.700 ;
        RECT 646.950 204.600 648.150 219.600 ;
        RECT 661.950 214.950 664.050 217.050 ;
        RECT 668.400 216.600 669.450 223.950 ;
        RECT 662.400 214.200 663.600 214.950 ;
        RECT 668.400 214.200 669.600 216.600 ;
        RECT 649.950 211.950 652.050 214.050 ;
        RECT 661.950 211.800 664.050 213.900 ;
        RECT 664.950 211.800 667.050 213.900 ;
        RECT 667.950 211.800 670.050 213.900 ;
        RECT 650.400 210.000 651.600 211.650 ;
        RECT 649.950 205.950 652.050 210.000 ;
        RECT 658.950 208.950 661.050 211.050 ;
        RECT 665.400 210.750 666.600 211.500 ;
        RECT 655.950 205.950 658.050 208.050 ;
        RECT 646.950 202.500 649.050 204.600 ;
        RECT 637.950 199.950 640.050 202.050 ;
        RECT 656.400 187.050 657.450 205.950 ;
        RECT 655.950 184.950 658.050 187.050 ;
        RECT 614.400 181.500 615.600 182.250 ;
        RECT 629.400 181.500 630.600 182.250 ;
        RECT 635.400 181.500 636.600 183.600 ;
        RECT 649.950 182.100 652.050 184.200 ;
        RECT 656.400 183.600 657.450 184.950 ;
        RECT 659.400 184.050 660.450 208.950 ;
        RECT 664.950 208.650 667.050 210.750 ;
        RECT 670.950 208.950 673.050 211.050 ;
        RECT 664.950 188.400 667.050 190.500 ;
        RECT 650.400 181.350 651.600 182.100 ;
        RECT 656.400 181.350 657.600 183.600 ;
        RECT 658.950 183.450 661.050 184.050 ;
        RECT 662.400 183.450 663.600 183.600 ;
        RECT 658.950 182.400 663.600 183.450 ;
        RECT 658.950 181.950 661.050 182.400 ;
        RECT 662.400 181.350 663.600 182.400 ;
        RECT 610.950 179.100 613.050 181.200 ;
        RECT 613.950 179.100 616.050 181.200 ;
        RECT 616.950 179.100 619.050 181.200 ;
        RECT 625.950 179.100 628.050 181.200 ;
        RECT 628.950 179.100 631.050 181.200 ;
        RECT 631.950 179.100 634.050 181.200 ;
        RECT 634.950 179.100 637.050 181.200 ;
        RECT 649.950 178.950 652.050 181.050 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 655.950 178.950 658.050 181.050 ;
        RECT 661.950 178.950 664.050 181.050 ;
        RECT 611.400 178.050 612.600 178.800 ;
        RECT 610.950 175.950 613.050 178.050 ;
        RECT 617.400 176.400 618.600 178.800 ;
        RECT 617.400 172.050 618.450 176.400 ;
        RECT 622.950 175.950 625.050 178.050 ;
        RECT 626.400 177.450 627.600 178.800 ;
        RECT 632.400 178.050 633.600 178.800 ;
        RECT 626.400 176.400 630.450 177.450 ;
        RECT 616.950 169.950 619.050 172.050 ;
        RECT 604.950 148.950 607.050 151.050 ;
        RECT 613.950 148.950 616.050 151.050 ;
        RECT 607.950 142.950 610.050 145.050 ;
        RECT 595.950 136.950 598.050 142.050 ;
        RECT 601.950 138.000 604.050 142.050 ;
        RECT 608.400 138.600 609.450 142.950 ;
        RECT 602.400 136.350 603.600 138.000 ;
        RECT 608.400 136.350 609.600 138.600 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 604.950 133.950 607.050 136.050 ;
        RECT 607.950 133.950 610.050 136.050 ;
        RECT 599.400 132.900 600.600 133.650 ;
        RECT 598.950 130.800 601.050 132.900 ;
        RECT 605.400 131.400 606.600 133.650 ;
        RECT 595.950 127.950 598.050 130.050 ;
        RECT 592.950 106.950 595.050 109.050 ;
        RECT 574.950 103.950 577.050 106.050 ;
        RECT 580.950 104.250 583.050 106.350 ;
        RECT 581.400 103.500 582.600 104.250 ;
        RECT 589.950 103.950 592.050 106.050 ;
        RECT 596.400 105.600 597.450 127.950 ;
        RECT 605.400 106.050 606.450 131.400 ;
        RECT 614.400 112.050 615.450 148.950 ;
        RECT 623.400 138.600 624.450 175.950 ;
        RECT 629.400 139.050 630.450 176.400 ;
        RECT 631.950 175.950 634.050 178.050 ;
        RECT 653.400 177.900 654.600 178.650 ;
        RECT 652.950 175.800 655.050 177.900 ;
        RECT 658.950 175.950 661.050 178.050 ;
        RECT 640.950 154.950 643.050 157.050 ;
        RECT 631.950 139.950 634.050 142.050 ;
        RECT 623.400 136.350 624.600 138.600 ;
        RECT 628.950 136.950 631.050 139.050 ;
        RECT 619.950 133.950 622.050 136.050 ;
        RECT 622.950 133.950 625.050 136.050 ;
        RECT 625.950 133.950 628.050 136.050 ;
        RECT 620.400 131.400 621.600 133.650 ;
        RECT 626.400 132.450 627.600 133.650 ;
        RECT 632.400 133.050 633.450 139.950 ;
        RECT 634.950 136.950 637.050 139.050 ;
        RECT 641.400 138.600 642.450 154.950 ;
        RECT 646.950 142.950 649.050 145.050 ;
        RECT 647.400 138.600 648.450 142.950 ;
        RECT 659.400 141.450 660.450 175.950 ;
        RECT 665.850 173.400 667.050 188.400 ;
        RECT 664.950 171.300 667.050 173.400 ;
        RECT 665.850 167.700 667.050 171.300 ;
        RECT 664.950 165.600 667.050 167.700 ;
        RECT 671.400 148.050 672.450 208.950 ;
        RECT 670.950 145.950 673.050 148.050 ;
        RECT 667.950 144.900 672.000 145.050 ;
        RECT 667.950 142.950 673.050 144.900 ;
        RECT 670.950 142.800 673.050 142.950 ;
        RECT 659.400 140.400 663.450 141.450 ;
        RECT 662.400 138.600 663.450 140.400 ;
        RECT 626.400 131.400 630.450 132.450 ;
        RECT 620.400 115.050 621.450 131.400 ;
        RECT 625.950 127.950 628.050 130.050 ;
        RECT 619.950 112.950 622.050 115.050 ;
        RECT 607.950 109.950 610.050 112.050 ;
        RECT 613.950 109.950 616.050 112.050 ;
        RECT 577.950 101.100 580.050 103.200 ;
        RECT 580.950 101.100 583.050 103.200 ;
        RECT 583.950 101.100 586.050 103.200 ;
        RECT 578.400 100.050 579.600 100.800 ;
        RECT 562.950 97.950 565.050 100.050 ;
        RECT 571.950 97.950 574.050 100.050 ;
        RECT 577.950 97.950 580.050 100.050 ;
        RECT 584.400 98.400 585.600 100.800 ;
        RECT 563.400 91.050 564.450 97.950 ;
        RECT 584.400 91.050 585.450 98.400 ;
        RECT 562.950 88.950 565.050 91.050 ;
        RECT 574.950 88.950 577.050 91.050 ;
        RECT 583.950 88.950 586.050 91.050 ;
        RECT 562.950 68.400 565.050 70.500 ;
        RECT 575.400 70.050 576.450 88.950 ;
        RECT 590.400 85.050 591.450 103.950 ;
        RECT 596.400 103.350 597.600 105.600 ;
        RECT 604.950 103.950 607.050 106.050 ;
        RECT 595.950 100.950 598.050 103.050 ;
        RECT 601.950 100.950 604.050 103.050 ;
        RECT 602.400 99.900 603.600 100.650 ;
        RECT 601.950 97.800 604.050 99.900 ;
        RECT 589.950 82.950 592.050 85.050 ;
        RECT 547.950 59.100 550.050 59.400 ;
        RECT 548.400 58.200 549.600 59.100 ;
        RECT 554.400 58.200 555.600 60.600 ;
        RECT 556.950 60.450 559.050 61.050 ;
        RECT 560.400 60.450 561.600 60.600 ;
        RECT 556.950 59.400 561.600 60.450 ;
        RECT 556.950 58.950 559.050 59.400 ;
        RECT 560.400 58.350 561.600 59.400 ;
        RECT 547.950 55.800 550.050 57.900 ;
        RECT 550.950 55.800 553.050 57.900 ;
        RECT 553.950 55.800 556.050 57.900 ;
        RECT 559.950 55.950 562.050 58.050 ;
        RECT 551.400 53.400 552.600 55.500 ;
        RECT 541.950 49.950 544.050 52.050 ;
        RECT 551.400 49.050 552.450 53.400 ;
        RECT 556.950 52.950 559.050 55.050 ;
        RECT 538.950 46.950 541.050 49.050 ;
        RECT 550.950 46.950 553.050 49.050 ;
        RECT 557.400 40.050 558.450 52.950 ;
        RECT 563.700 48.600 564.900 68.400 ;
        RECT 574.950 67.950 577.050 70.050 ;
        RECT 583.950 69.300 586.050 71.400 ;
        RECT 592.950 70.950 595.050 73.050 ;
        RECT 598.950 70.950 601.050 73.050 ;
        RECT 577.950 64.950 580.050 67.050 ;
        RECT 583.950 65.700 585.150 69.300 ;
        RECT 568.950 59.100 571.050 61.200 ;
        RECT 574.950 59.100 577.050 61.200 ;
        RECT 569.400 58.350 570.600 59.100 ;
        RECT 568.950 55.950 571.050 58.050 ;
        RECT 562.950 46.500 565.050 48.600 ;
        RECT 575.400 46.050 576.450 59.100 ;
        RECT 578.400 54.900 579.450 64.950 ;
        RECT 583.950 63.600 586.050 65.700 ;
        RECT 577.950 52.800 580.050 54.900 ;
        RECT 583.950 48.600 585.150 63.600 ;
        RECT 586.950 55.950 589.050 58.050 ;
        RECT 587.400 54.900 588.600 55.650 ;
        RECT 586.950 52.800 589.050 54.900 ;
        RECT 583.950 46.500 586.050 48.600 ;
        RECT 574.950 43.950 577.050 46.050 ;
        RECT 535.950 37.950 538.050 40.050 ;
        RECT 556.950 37.950 559.050 40.050 ;
        RECT 562.950 37.950 565.050 40.050 ;
        RECT 532.950 32.400 535.050 34.500 ;
        RECT 518.400 25.350 519.600 27.600 ;
        RECT 524.400 25.350 525.600 27.600 ;
        RECT 529.950 26.100 532.050 28.200 ;
        RECT 530.400 25.350 531.600 26.100 ;
        RECT 514.950 22.950 517.050 25.050 ;
        RECT 517.950 22.950 520.050 25.050 ;
        RECT 520.950 22.950 523.050 25.050 ;
        RECT 523.950 22.950 526.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 515.400 21.900 516.600 22.650 ;
        RECT 521.400 21.900 522.600 22.650 ;
        RECT 514.950 19.800 517.050 21.900 ;
        RECT 520.950 16.950 523.050 21.900 ;
        RECT 526.950 19.950 529.050 22.050 ;
        RECT 508.950 13.950 511.050 16.050 ;
        RECT 517.950 15.450 520.050 16.050 ;
        RECT 523.950 15.450 526.050 16.050 ;
        RECT 517.950 14.400 526.050 15.450 ;
        RECT 517.950 13.950 520.050 14.400 ;
        RECT 523.950 13.950 526.050 14.400 ;
        RECT 502.950 10.950 505.050 13.050 ;
        RECT 514.950 12.450 517.050 13.050 ;
        RECT 527.400 12.450 528.450 19.950 ;
        RECT 533.850 17.400 535.050 32.400 ;
        RECT 538.950 31.950 541.050 34.050 ;
        RECT 553.950 32.400 556.050 34.500 ;
        RECT 532.950 15.300 535.050 17.400 ;
        RECT 539.400 16.050 540.450 31.950 ;
        RECT 547.950 22.950 550.050 25.050 ;
        RECT 548.400 20.400 549.600 22.650 ;
        RECT 514.950 11.400 528.450 12.450 ;
        RECT 533.850 11.700 535.050 15.300 ;
        RECT 538.950 13.950 541.050 16.050 ;
        RECT 514.950 10.950 517.050 11.400 ;
        RECT 490.950 7.950 493.050 10.050 ;
        RECT 532.950 9.600 535.050 11.700 ;
        RECT 548.400 10.050 549.450 20.400 ;
        RECT 554.100 12.600 555.300 32.400 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 557.400 21.900 558.600 22.650 ;
        RECT 563.400 21.900 564.450 37.950 ;
        RECT 593.400 37.050 594.450 70.950 ;
        RECT 599.400 60.600 600.450 70.950 ;
        RECT 604.950 64.950 607.050 67.050 ;
        RECT 605.400 60.600 606.450 64.950 ;
        RECT 608.400 61.050 609.450 109.950 ;
        RECT 613.950 104.100 616.050 106.200 ;
        RECT 614.400 103.350 615.600 104.100 ;
        RECT 613.950 100.950 616.050 103.050 ;
        RECT 619.950 100.950 622.050 103.050 ;
        RECT 610.950 97.950 613.050 100.050 ;
        RECT 611.400 94.050 612.450 97.950 ;
        RECT 613.950 94.950 616.050 97.050 ;
        RECT 610.950 91.950 613.050 94.050 ;
        RECT 614.400 90.450 615.450 94.950 ;
        RECT 622.950 91.950 625.050 94.050 ;
        RECT 611.400 89.400 615.450 90.450 ;
        RECT 599.400 58.200 600.600 60.600 ;
        RECT 605.400 58.200 606.600 60.600 ;
        RECT 607.950 58.950 610.050 61.050 ;
        RECT 598.950 55.800 601.050 57.900 ;
        RECT 601.950 55.800 604.050 57.900 ;
        RECT 604.950 55.800 607.050 57.900 ;
        RECT 602.400 54.750 603.600 55.500 ;
        RECT 611.400 55.050 612.450 89.400 ;
        RECT 623.400 85.050 624.450 91.950 ;
        RECT 626.400 88.050 627.450 127.950 ;
        RECT 629.400 127.050 630.450 131.400 ;
        RECT 631.950 130.950 634.050 133.050 ;
        RECT 635.400 130.050 636.450 136.950 ;
        RECT 641.400 136.350 642.600 138.600 ;
        RECT 647.400 136.350 648.600 138.600 ;
        RECT 662.400 136.350 663.600 138.600 ;
        RECT 667.950 137.100 670.050 139.200 ;
        RECT 668.400 136.350 669.600 137.100 ;
        RECT 640.950 133.950 643.050 136.050 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 646.950 133.950 649.050 136.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 658.950 133.950 661.050 136.050 ;
        RECT 661.950 133.950 664.050 136.050 ;
        RECT 664.950 133.950 667.050 136.050 ;
        RECT 667.950 133.950 670.050 136.050 ;
        RECT 644.400 131.400 645.600 133.650 ;
        RECT 650.400 131.400 651.600 133.650 ;
        RECT 659.400 131.400 660.600 133.650 ;
        RECT 665.400 132.900 666.600 133.650 ;
        RECT 634.950 127.950 637.050 130.050 ;
        RECT 628.950 124.950 631.050 127.050 ;
        RECT 628.950 109.950 631.050 112.050 ;
        RECT 629.400 106.050 630.450 109.950 ;
        RECT 628.950 103.950 631.050 106.050 ;
        RECT 631.950 104.100 634.050 106.200 ;
        RECT 632.400 103.350 633.600 104.100 ;
        RECT 631.950 100.950 634.050 103.050 ;
        RECT 637.950 100.950 640.050 103.050 ;
        RECT 628.950 97.050 631.050 100.050 ;
        RECT 628.800 96.000 631.050 97.050 ;
        RECT 628.800 94.950 630.900 96.000 ;
        RECT 631.950 94.950 634.050 97.050 ;
        RECT 628.950 88.950 631.050 91.050 ;
        RECT 625.950 85.950 628.050 88.050 ;
        RECT 622.950 82.950 625.050 85.050 ;
        RECT 629.400 84.450 630.450 88.950 ;
        RECT 626.400 83.400 630.450 84.450 ;
        RECT 626.400 81.450 627.450 83.400 ;
        RECT 623.400 81.000 627.450 81.450 ;
        RECT 622.950 80.400 627.450 81.000 ;
        RECT 622.950 76.950 625.050 80.400 ;
        RECT 613.950 58.950 616.050 61.050 ;
        RECT 601.950 52.650 604.050 54.750 ;
        RECT 610.950 52.950 613.050 55.050 ;
        RECT 614.400 52.050 615.450 58.950 ;
        RECT 619.950 58.800 622.050 60.900 ;
        RECT 625.950 60.000 628.050 64.050 ;
        RECT 620.400 58.200 621.600 58.800 ;
        RECT 626.400 58.200 627.600 60.000 ;
        RECT 619.950 55.800 622.050 57.900 ;
        RECT 622.950 55.800 625.050 57.900 ;
        RECT 625.950 55.800 628.050 57.900 ;
        RECT 623.400 53.400 624.600 55.500 ;
        RECT 613.950 49.950 616.050 52.050 ;
        RECT 623.400 43.050 624.450 53.400 ;
        RECT 622.950 40.950 625.050 43.050 ;
        RECT 632.400 40.050 633.450 94.950 ;
        RECT 644.400 79.050 645.450 131.400 ;
        RECT 650.400 127.050 651.450 131.400 ;
        RECT 649.950 124.950 652.050 127.050 ;
        RECT 659.400 115.050 660.450 131.400 ;
        RECT 664.950 130.800 667.050 132.900 ;
        RECT 670.950 130.950 673.050 133.050 ;
        RECT 661.950 124.950 664.050 127.050 ;
        RECT 658.950 112.950 661.050 115.050 ;
        RECT 649.950 109.950 652.050 112.050 ;
        RECT 646.950 104.100 649.050 106.200 ;
        RECT 650.400 106.050 651.450 109.950 ;
        RECT 647.400 97.050 648.450 104.100 ;
        RECT 649.950 103.950 652.050 106.050 ;
        RECT 655.950 104.100 658.050 106.200 ;
        RECT 662.400 105.600 663.450 124.950 ;
        RECT 671.400 121.050 672.450 130.950 ;
        RECT 674.400 130.050 675.450 250.950 ;
        RECT 676.950 247.950 679.050 250.050 ;
        RECT 677.400 211.050 678.450 247.950 ;
        RECT 680.400 217.050 681.450 251.400 ;
        RECT 679.950 214.950 682.050 217.050 ;
        RECT 682.950 215.100 685.050 217.200 ;
        RECT 689.400 216.600 690.450 253.950 ;
        RECT 692.400 247.050 693.450 254.400 ;
        RECT 697.950 253.800 700.050 255.900 ;
        RECT 691.950 244.950 694.050 247.050 ;
        RECT 707.400 220.050 708.450 256.800 ;
        RECT 713.400 255.900 714.600 256.650 ;
        RECT 722.400 256.050 723.450 283.950 ;
        RECT 728.400 283.050 729.450 298.950 ;
        RECT 740.400 294.600 741.450 301.950 ;
        RECT 746.400 295.050 747.450 328.950 ;
        RECT 757.950 319.950 760.050 322.050 ;
        RECT 769.950 319.950 772.050 322.050 ;
        RECT 751.950 304.950 754.050 307.050 ;
        RECT 752.400 298.050 753.450 304.950 ;
        RECT 740.400 292.350 741.600 294.600 ;
        RECT 745.950 292.950 748.050 295.050 ;
        RECT 751.950 294.000 754.050 298.050 ;
        RECT 758.400 294.600 759.450 319.950 ;
        RECT 752.400 292.200 753.600 294.000 ;
        RECT 758.400 292.200 759.600 294.600 ;
        RECT 736.950 289.950 739.050 292.050 ;
        RECT 739.950 289.950 742.050 292.050 ;
        RECT 742.950 289.950 745.050 292.050 ;
        RECT 751.950 289.800 754.050 291.900 ;
        RECT 754.950 289.800 757.050 291.900 ;
        RECT 757.950 289.800 760.050 291.900 ;
        RECT 760.950 289.800 763.050 291.900 ;
        RECT 737.400 287.400 738.600 289.650 ;
        RECT 743.400 288.900 744.600 289.650 ;
        RECT 727.950 280.950 730.050 283.050 ;
        RECT 737.400 271.050 738.450 287.400 ;
        RECT 742.950 283.950 745.050 288.900 ;
        RECT 755.400 288.000 756.600 289.500 ;
        RECT 754.950 283.950 757.050 288.000 ;
        RECT 761.400 287.400 762.600 289.500 ;
        RECT 770.400 288.900 771.450 319.950 ;
        RECT 782.400 316.050 783.450 332.400 ;
        RECT 791.400 328.050 792.450 338.400 ;
        RECT 796.950 338.100 799.050 340.200 ;
        RECT 803.400 339.450 804.600 339.600 ;
        RECT 806.400 339.450 807.450 365.400 ;
        RECT 803.400 338.400 807.450 339.450 ;
        RECT 797.400 337.350 798.600 338.100 ;
        RECT 803.400 337.350 804.600 338.400 ;
        RECT 796.950 334.950 799.050 337.050 ;
        RECT 799.950 334.950 802.050 337.050 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 800.400 332.400 801.600 334.650 ;
        RECT 790.950 325.950 793.050 328.050 ;
        RECT 781.950 313.950 784.050 316.050 ;
        RECT 796.950 313.950 799.050 316.050 ;
        RECT 793.950 307.950 796.050 310.050 ;
        RECT 794.400 301.050 795.450 307.950 ;
        RECT 793.950 298.950 796.050 301.050 ;
        RECT 778.950 294.000 781.050 298.050 ;
        RECT 790.950 294.000 793.050 298.050 ;
        RECT 797.400 295.050 798.450 313.950 ;
        RECT 800.400 295.050 801.450 332.400 ;
        RECT 805.950 316.950 808.050 319.050 ;
        RECT 802.950 301.950 805.050 304.050 ;
        RECT 779.400 292.350 780.600 294.000 ;
        RECT 791.400 292.200 792.600 294.000 ;
        RECT 796.950 292.950 799.050 295.050 ;
        RECT 799.950 292.950 802.050 295.050 ;
        RECT 797.400 292.200 798.600 292.950 ;
        RECT 775.950 289.950 778.050 292.050 ;
        RECT 778.950 289.950 781.050 292.050 ;
        RECT 781.950 289.950 784.050 292.050 ;
        RECT 790.950 289.800 793.050 291.900 ;
        RECT 793.950 289.800 796.050 291.900 ;
        RECT 796.950 289.800 799.050 291.900 ;
        RECT 776.400 288.900 777.600 289.650 ;
        RECT 754.950 277.950 757.050 280.050 ;
        RECT 736.950 268.950 739.050 271.050 ;
        RECT 727.950 260.100 730.050 262.200 ;
        RECT 733.950 260.100 736.050 262.200 ;
        RECT 745.950 260.250 748.050 262.350 ;
        RECT 751.950 261.000 754.050 265.050 ;
        RECT 755.400 262.050 756.450 277.950 ;
        RECT 761.400 277.050 762.450 287.400 ;
        RECT 769.950 286.800 772.050 288.900 ;
        RECT 775.950 286.800 778.050 288.900 ;
        RECT 782.400 288.000 783.600 289.650 ;
        RECT 781.950 283.950 784.050 288.000 ;
        RECT 794.400 287.400 795.600 289.500 ;
        RECT 760.950 274.950 763.050 277.050 ;
        RECT 778.950 274.950 781.050 277.050 ;
        RECT 775.950 268.950 778.050 271.050 ;
        RECT 728.400 259.350 729.600 260.100 ;
        RECT 734.400 259.350 735.600 260.100 ;
        RECT 746.400 259.500 747.600 260.250 ;
        RECT 752.400 259.500 753.600 261.000 ;
        RECT 754.950 259.950 757.050 262.050 ;
        RECT 757.950 260.100 760.050 262.200 ;
        RECT 763.950 260.100 766.050 262.200 ;
        RECT 769.950 260.100 772.050 265.050 ;
        RECT 727.950 256.950 730.050 259.050 ;
        RECT 730.950 256.950 733.050 259.050 ;
        RECT 733.950 256.950 736.050 259.050 ;
        RECT 742.950 257.100 745.050 259.200 ;
        RECT 745.950 257.100 748.050 259.200 ;
        RECT 748.950 257.100 751.050 259.200 ;
        RECT 751.950 257.100 754.050 259.200 ;
        RECT 712.950 253.800 715.050 255.900 ;
        RECT 718.950 253.950 721.050 256.050 ;
        RECT 721.950 253.950 724.050 256.050 ;
        RECT 731.400 254.400 732.600 256.650 ;
        RECT 743.400 256.050 744.600 256.800 ;
        RECT 709.950 244.950 712.050 247.050 ;
        RECT 706.950 217.950 709.050 220.050 ;
        RECT 710.400 217.050 711.450 244.950 ;
        RECT 719.400 225.450 720.450 253.950 ;
        RECT 731.400 247.050 732.450 254.400 ;
        RECT 736.950 253.950 739.050 256.050 ;
        RECT 742.800 253.950 744.900 256.050 ;
        RECT 745.950 253.950 748.050 256.050 ;
        RECT 749.400 255.450 750.600 256.800 ;
        RECT 754.950 255.450 757.050 256.050 ;
        RECT 749.400 254.400 757.050 255.450 ;
        RECT 754.950 253.950 757.050 254.400 ;
        RECT 730.950 244.950 733.050 247.050 ;
        RECT 737.400 232.050 738.450 253.950 ;
        RECT 746.400 247.050 747.450 253.950 ;
        RECT 758.400 250.050 759.450 260.100 ;
        RECT 764.400 259.350 765.600 260.100 ;
        RECT 770.400 259.350 771.600 260.100 ;
        RECT 763.950 256.950 766.050 259.050 ;
        RECT 766.950 256.950 769.050 259.050 ;
        RECT 769.950 256.950 772.050 259.050 ;
        RECT 767.400 255.900 768.600 256.650 ;
        RECT 776.400 256.050 777.450 268.950 ;
        RECT 766.950 253.800 769.050 255.900 ;
        RECT 775.950 253.950 778.050 256.050 ;
        RECT 779.400 253.050 780.450 274.950 ;
        RECT 787.950 260.100 790.050 262.200 ;
        RECT 794.400 261.600 795.450 287.400 ;
        RECT 799.950 286.950 802.050 289.050 ;
        RECT 788.400 259.350 789.600 260.100 ;
        RECT 794.400 259.350 795.600 261.600 ;
        RECT 800.400 261.450 801.450 286.950 ;
        RECT 803.400 265.050 804.450 301.950 ;
        RECT 806.400 295.050 807.450 316.950 ;
        RECT 809.400 298.050 810.450 370.950 ;
        RECT 812.400 364.050 813.450 379.950 ;
        RECT 814.950 376.950 817.050 379.050 ;
        RECT 815.400 373.050 816.450 376.950 ;
        RECT 814.950 370.950 817.050 373.050 ;
        RECT 818.400 372.600 819.450 409.950 ;
        RECT 823.950 409.800 826.050 411.900 ;
        RECT 826.950 409.950 829.050 412.050 ;
        RECT 823.950 382.950 826.050 385.050 ;
        RECT 824.400 372.600 825.450 382.950 ;
        RECT 827.400 373.050 828.450 409.950 ;
        RECT 830.400 397.050 831.450 424.950 ;
        RECT 839.400 421.050 840.450 437.400 ;
        RECT 838.950 418.950 841.050 421.050 ;
        RECT 835.950 416.100 838.050 418.200 ;
        RECT 836.400 415.350 837.600 416.100 ;
        RECT 847.950 415.950 850.050 418.050 ;
        RECT 835.950 412.950 838.050 415.050 ;
        RECT 841.950 412.950 844.050 415.050 ;
        RECT 844.950 409.950 847.050 412.050 ;
        RECT 829.950 394.950 832.050 397.050 ;
        RECT 838.950 388.950 841.050 391.050 ;
        RECT 832.950 376.950 835.050 379.050 ;
        RECT 818.400 370.200 819.600 372.600 ;
        RECT 824.400 370.200 825.600 372.600 ;
        RECT 826.950 370.950 829.050 373.050 ;
        RECT 833.400 372.600 834.450 376.950 ;
        RECT 839.400 373.050 840.450 388.950 ;
        RECT 833.400 370.200 834.600 372.600 ;
        RECT 838.950 370.950 841.050 373.050 ;
        RECT 839.400 370.200 840.600 370.950 ;
        RECT 817.950 367.800 820.050 369.900 ;
        RECT 820.950 367.800 823.050 369.900 ;
        RECT 823.950 367.800 826.050 369.900 ;
        RECT 832.950 367.800 835.050 369.900 ;
        RECT 835.950 367.800 838.050 369.900 ;
        RECT 838.950 367.800 841.050 369.900 ;
        RECT 814.950 364.950 817.050 367.050 ;
        RECT 821.400 365.400 822.600 367.500 ;
        RECT 836.400 366.000 837.600 367.500 ;
        RECT 811.950 361.950 814.050 364.050 ;
        RECT 815.400 339.450 816.450 364.950 ;
        RECT 821.400 352.050 822.450 365.400 ;
        RECT 835.950 361.950 838.050 366.000 ;
        RECT 820.950 349.950 823.050 352.050 ;
        RECT 829.950 346.950 832.050 349.050 ;
        RECT 826.950 343.950 829.050 346.050 ;
        RECT 812.400 338.400 816.450 339.450 ;
        RECT 812.400 304.050 813.450 338.400 ;
        RECT 820.950 338.100 823.050 340.200 ;
        RECT 821.400 337.350 822.600 338.100 ;
        RECT 817.950 334.950 820.050 337.050 ;
        RECT 820.950 334.950 823.050 337.050 ;
        RECT 814.950 331.950 817.050 334.050 ;
        RECT 818.400 332.400 819.600 334.650 ;
        RECT 815.400 319.050 816.450 331.950 ;
        RECT 818.400 322.050 819.450 332.400 ;
        RECT 823.950 331.950 826.050 334.050 ;
        RECT 817.950 319.950 820.050 322.050 ;
        RECT 814.950 316.950 817.050 319.050 ;
        RECT 815.400 310.050 816.450 316.950 ;
        RECT 814.950 307.950 817.050 310.050 ;
        RECT 811.950 301.950 814.050 304.050 ;
        RECT 808.950 295.950 811.050 298.050 ;
        RECT 805.950 292.950 808.050 295.050 ;
        RECT 812.400 294.600 813.450 301.950 ;
        RECT 812.400 292.350 813.600 294.600 ;
        RECT 817.950 293.100 820.050 295.200 ;
        RECT 818.400 292.350 819.600 293.100 ;
        RECT 808.950 289.950 811.050 292.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 814.950 289.950 817.050 292.050 ;
        RECT 817.950 289.950 820.050 292.050 ;
        RECT 805.950 286.950 808.050 289.050 ;
        RECT 809.400 288.900 810.600 289.650 ;
        RECT 806.400 283.050 807.450 286.950 ;
        RECT 808.950 286.800 811.050 288.900 ;
        RECT 815.400 287.400 816.600 289.650 ;
        RECT 811.950 283.950 814.050 286.050 ;
        RECT 805.950 280.950 808.050 283.050 ;
        RECT 802.950 262.950 805.050 265.050 ;
        RECT 812.400 262.050 813.450 283.950 ;
        RECT 815.400 280.050 816.450 287.400 ;
        RECT 820.950 286.950 823.050 289.050 ;
        RECT 814.950 277.950 817.050 280.050 ;
        RECT 821.400 274.050 822.450 286.950 ;
        RECT 820.950 271.950 823.050 274.050 ;
        RECT 817.950 266.400 820.050 268.500 ;
        RECT 803.400 261.450 804.600 261.600 ;
        RECT 800.400 260.400 804.600 261.450 ;
        RECT 803.400 259.350 804.600 260.400 ;
        RECT 811.950 259.950 814.050 262.050 ;
        RECT 784.950 256.950 787.050 259.050 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 802.950 256.950 805.050 259.050 ;
        RECT 805.950 256.950 808.050 259.050 ;
        RECT 814.950 256.950 817.050 259.050 ;
        RECT 785.400 255.000 786.600 256.650 ;
        RECT 791.400 255.900 792.600 256.650 ;
        RECT 778.950 250.950 781.050 253.050 ;
        RECT 784.950 250.950 787.050 255.000 ;
        RECT 790.950 253.800 793.050 255.900 ;
        RECT 796.950 253.950 799.050 256.050 ;
        RECT 806.400 254.400 807.600 256.650 ;
        RECT 757.950 249.450 760.050 250.050 ;
        RECT 757.950 248.400 762.450 249.450 ;
        RECT 757.950 247.950 760.050 248.400 ;
        RECT 745.950 244.950 748.050 247.050 ;
        RECT 751.950 238.950 754.050 241.050 ;
        RECT 739.950 232.950 742.050 235.050 ;
        RECT 736.950 229.950 739.050 232.050 ;
        RECT 716.400 224.400 720.450 225.450 ;
        RECT 683.400 214.350 684.600 215.100 ;
        RECT 689.400 214.350 690.600 216.600 ;
        RECT 697.950 214.950 700.050 217.050 ;
        RECT 703.950 214.950 706.050 217.050 ;
        RECT 709.950 214.950 712.050 217.050 ;
        RECT 716.400 216.450 717.450 224.400 ;
        RECT 721.800 219.300 723.900 221.400 ;
        RECT 731.400 220.500 733.500 222.600 ;
        RECT 719.400 216.450 720.600 216.600 ;
        RECT 716.400 215.400 720.600 216.450 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 688.950 211.950 691.050 214.050 ;
        RECT 691.950 211.950 694.050 214.050 ;
        RECT 676.950 208.950 679.050 211.050 ;
        RECT 679.950 205.950 682.050 211.050 ;
        RECT 686.400 209.400 687.600 211.650 ;
        RECT 692.400 210.000 693.600 211.650 ;
        RECT 686.400 196.050 687.450 209.400 ;
        RECT 691.950 205.950 694.050 210.000 ;
        RECT 694.950 208.950 697.050 211.050 ;
        RECT 676.950 193.950 679.050 196.050 ;
        RECT 685.950 193.950 688.050 196.050 ;
        RECT 677.400 184.050 678.450 193.950 ;
        RECT 685.950 188.400 688.050 190.500 ;
        RECT 676.950 181.950 679.050 184.050 ;
        RECT 679.950 178.950 682.050 181.050 ;
        RECT 680.400 177.900 681.600 178.650 ;
        RECT 679.950 175.800 682.050 177.900 ;
        RECT 686.100 168.600 687.300 188.400 ;
        RECT 688.950 178.950 691.050 181.050 ;
        RECT 689.400 177.450 690.600 178.650 ;
        RECT 689.400 176.400 693.450 177.450 ;
        RECT 685.950 166.500 688.050 168.600 ;
        RECT 692.400 166.050 693.450 176.400 ;
        RECT 695.400 172.050 696.450 208.950 ;
        RECT 698.400 205.050 699.450 214.950 ;
        RECT 704.400 214.200 705.600 214.950 ;
        RECT 710.400 214.200 711.600 214.950 ;
        RECT 719.400 213.900 720.600 215.400 ;
        RECT 703.950 211.800 706.050 213.900 ;
        RECT 706.950 211.800 709.050 213.900 ;
        RECT 709.950 211.800 712.050 213.900 ;
        RECT 718.950 211.800 721.050 213.900 ;
        RECT 707.400 210.750 708.600 211.500 ;
        RECT 706.950 208.650 709.050 210.750 ;
        RECT 722.700 210.300 723.600 219.300 ;
        RECT 724.950 215.700 727.050 217.800 ;
        RECT 728.400 216.900 729.600 219.600 ;
        RECT 726.150 213.300 727.050 215.700 ;
        RECT 727.950 214.800 730.050 216.900 ;
        RECT 731.850 213.300 733.050 220.500 ;
        RECT 737.400 217.050 738.450 229.950 ;
        RECT 736.950 214.950 739.050 217.050 ;
        RECT 726.150 212.100 733.050 213.300 ;
        RECT 729.150 210.300 731.250 211.200 ;
        RECT 722.700 209.100 731.250 210.300 ;
        RECT 724.200 207.300 726.300 209.100 ;
        RECT 727.950 206.100 730.050 208.200 ;
        RECT 732.150 206.700 733.050 212.100 ;
        RECT 733.950 211.800 736.050 213.900 ;
        RECT 734.400 209.400 735.600 211.800 ;
        RECT 740.400 210.900 741.450 232.950 ;
        RECT 752.400 226.050 753.450 238.950 ;
        RECT 757.950 232.950 760.050 235.050 ;
        RECT 751.950 223.950 754.050 226.050 ;
        RECT 752.400 216.600 753.450 223.950 ;
        RECT 752.400 214.350 753.600 216.600 ;
        RECT 745.950 211.950 748.050 214.050 ;
        RECT 751.950 211.950 754.050 214.050 ;
        RECT 746.400 210.900 747.600 211.650 ;
        RECT 739.950 208.800 742.050 210.900 ;
        RECT 745.950 208.800 748.050 210.900 ;
        RECT 697.950 202.950 700.050 205.050 ;
        RECT 728.400 203.400 729.600 206.100 ;
        RECT 731.400 204.600 733.500 206.700 ;
        RECT 697.950 190.950 700.050 193.050 ;
        RECT 706.950 190.950 709.050 193.050 ;
        RECT 694.950 169.950 697.050 172.050 ;
        RECT 698.400 166.050 699.450 190.950 ;
        RECT 700.950 181.950 703.050 187.050 ;
        RECT 707.400 183.600 708.450 190.950 ;
        RECT 728.400 187.050 729.450 203.400 ;
        RECT 730.950 187.950 733.050 190.050 ;
        RECT 727.950 184.950 730.050 187.050 ;
        RECT 707.400 181.500 708.600 183.600 ;
        RECT 703.950 179.100 706.050 181.200 ;
        RECT 706.950 179.100 709.050 181.200 ;
        RECT 709.950 179.100 712.050 181.200 ;
        RECT 715.950 178.950 718.050 184.050 ;
        RECT 724.950 182.100 727.050 184.200 ;
        RECT 731.400 183.600 732.450 187.950 ;
        RECT 725.400 181.350 726.600 182.100 ;
        RECT 731.400 181.350 732.600 183.600 ;
        RECT 740.400 183.450 741.450 208.800 ;
        RECT 745.950 187.950 748.050 190.050 ;
        RECT 751.950 187.950 754.050 190.050 ;
        RECT 737.400 182.400 741.450 183.450 ;
        RECT 746.400 183.600 747.450 187.950 ;
        RECT 752.400 183.600 753.450 187.950 ;
        RECT 758.400 184.050 759.450 232.950 ;
        RECT 761.400 190.050 762.450 248.400 ;
        RECT 791.400 235.050 792.450 253.800 ;
        RECT 793.950 241.950 796.050 244.050 ;
        RECT 790.950 232.950 793.050 235.050 ;
        RECT 766.950 229.950 769.050 232.050 ;
        RECT 767.400 216.600 768.450 229.950 ;
        RECT 790.950 223.950 793.050 226.050 ;
        RECT 767.400 214.350 768.600 216.600 ;
        RECT 781.950 215.100 784.050 217.200 ;
        RECT 782.400 214.350 783.600 215.100 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 769.950 211.950 772.050 214.050 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 781.950 211.950 784.050 214.050 ;
        RECT 784.950 211.950 787.050 214.050 ;
        RECT 770.400 210.900 771.600 211.650 ;
        RECT 769.950 208.800 772.050 210.900 ;
        RECT 779.400 209.400 780.600 211.650 ;
        RECT 785.400 210.900 786.600 211.650 ;
        RECT 779.400 205.050 780.450 209.400 ;
        RECT 784.950 208.800 787.050 210.900 ;
        RECT 778.950 202.950 781.050 205.050 ;
        RECT 763.950 196.950 766.050 199.050 ;
        RECT 760.950 187.950 763.050 190.050 ;
        RECT 764.400 184.050 765.450 196.950 ;
        RECT 766.950 187.950 769.050 190.050 ;
        RECT 775.950 187.950 778.050 190.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 727.950 178.950 730.050 181.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 704.400 178.050 705.600 178.800 ;
        RECT 703.950 175.950 706.050 178.050 ;
        RECT 710.400 176.400 711.600 178.800 ;
        RECT 710.400 172.050 711.450 176.400 ;
        RECT 715.950 175.800 718.050 177.900 ;
        RECT 718.950 175.950 721.050 178.050 ;
        RECT 722.400 177.900 723.600 178.650 ;
        RECT 709.950 169.950 712.050 172.050 ;
        RECT 691.950 163.950 694.050 166.050 ;
        RECT 697.950 163.950 700.050 166.050 ;
        RECT 692.400 160.050 693.450 163.950 ;
        RECT 691.950 157.950 694.050 160.050 ;
        RECT 710.400 157.050 711.450 169.950 ;
        RECT 688.950 154.950 691.050 157.050 ;
        RECT 709.950 154.950 712.050 157.050 ;
        RECT 676.950 145.950 679.050 148.050 ;
        RECT 677.400 139.050 678.450 145.950 ;
        RECT 679.950 142.950 685.050 145.050 ;
        RECT 676.950 136.950 679.050 139.050 ;
        RECT 682.950 137.100 685.050 139.200 ;
        RECT 683.400 136.350 684.600 137.100 ;
        RECT 679.950 133.950 682.050 136.050 ;
        RECT 682.950 133.950 685.050 136.050 ;
        RECT 676.950 130.950 679.050 133.050 ;
        RECT 680.400 131.400 681.600 133.650 ;
        RECT 673.950 127.950 676.050 130.050 ;
        RECT 670.950 118.950 673.050 121.050 ;
        RECT 677.400 112.050 678.450 130.950 ;
        RECT 680.400 121.050 681.450 131.400 ;
        RECT 685.950 130.950 688.050 133.050 ;
        RECT 682.950 127.950 685.050 130.050 ;
        RECT 683.400 123.450 684.450 127.950 ;
        RECT 686.400 127.050 687.450 130.950 ;
        RECT 685.950 124.950 688.050 127.050 ;
        RECT 683.400 122.400 687.450 123.450 ;
        RECT 679.950 118.950 682.050 121.050 ;
        RECT 686.400 118.050 687.450 122.400 ;
        RECT 685.950 115.950 688.050 118.050 ;
        RECT 682.950 112.950 685.050 115.050 ;
        RECT 667.950 109.950 670.050 112.050 ;
        RECT 676.950 109.950 679.050 112.050 ;
        RECT 656.400 103.350 657.600 104.100 ;
        RECT 662.400 103.350 663.600 105.600 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 661.950 100.950 664.050 103.050 ;
        RECT 649.950 97.950 652.050 100.050 ;
        RECT 653.400 98.400 654.600 100.650 ;
        RECT 659.400 99.900 660.600 100.650 ;
        RECT 646.950 94.950 649.050 97.050 ;
        RECT 650.400 79.050 651.450 97.950 ;
        RECT 653.400 91.050 654.450 98.400 ;
        RECT 658.950 97.800 661.050 99.900 ;
        RECT 652.950 88.950 655.050 91.050 ;
        RECT 634.950 76.950 637.050 79.050 ;
        RECT 643.950 76.950 646.050 79.050 ;
        RECT 649.950 76.950 652.050 79.050 ;
        RECT 635.400 61.050 636.450 76.950 ;
        RECT 668.400 67.050 669.450 109.950 ;
        RECT 676.950 104.100 679.050 106.200 ;
        RECT 683.400 105.600 684.450 112.950 ;
        RECT 686.400 106.050 687.450 115.950 ;
        RECT 689.400 109.050 690.450 154.950 ;
        RECT 697.950 145.950 700.050 148.050 ;
        RECT 709.950 147.300 712.050 149.400 ;
        RECT 691.950 142.950 694.050 145.050 ;
        RECT 692.400 139.050 693.450 142.950 ;
        RECT 691.950 136.950 694.050 139.050 ;
        RECT 698.400 138.600 699.450 145.950 ;
        RECT 710.850 143.700 712.050 147.300 ;
        RECT 709.950 141.600 712.050 143.700 ;
        RECT 698.400 136.350 699.600 138.600 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 697.950 133.950 700.050 136.050 ;
        RECT 706.950 133.950 709.050 136.050 ;
        RECT 691.950 130.950 694.050 133.050 ;
        RECT 695.400 131.400 696.600 133.650 ;
        RECT 707.400 133.050 708.600 133.650 ;
        RECT 703.950 131.400 708.600 133.050 ;
        RECT 688.950 106.950 691.050 109.050 ;
        RECT 677.400 103.350 678.600 104.100 ;
        RECT 683.400 103.350 684.600 105.600 ;
        RECT 685.950 103.950 688.050 106.050 ;
        RECT 692.400 105.450 693.450 130.950 ;
        RECT 695.400 118.050 696.450 131.400 ;
        RECT 703.950 130.950 708.000 131.400 ;
        RECT 710.850 126.600 712.050 141.600 ;
        RECT 709.950 124.500 712.050 126.600 ;
        RECT 694.950 115.950 697.050 118.050 ;
        RECT 697.950 109.950 700.050 112.050 ;
        RECT 689.400 104.400 693.450 105.450 ;
        RECT 698.400 105.600 699.450 109.950 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 676.950 100.950 679.050 103.050 ;
        RECT 679.950 100.950 682.050 103.050 ;
        RECT 682.950 100.950 685.050 103.050 ;
        RECT 674.400 99.450 675.600 100.650 ;
        RECT 671.400 98.400 675.600 99.450 ;
        RECT 680.400 98.400 681.600 100.650 ;
        RECT 671.400 94.050 672.450 98.400 ;
        RECT 670.950 91.950 673.050 94.050 ;
        RECT 680.400 85.050 681.450 98.400 ;
        RECT 685.950 97.950 688.050 100.050 ;
        RECT 679.950 82.950 682.050 85.050 ;
        RECT 667.950 64.950 670.050 67.050 ;
        RECT 679.950 64.950 682.050 67.050 ;
        RECT 686.400 66.450 687.450 97.950 ;
        RECT 689.400 85.050 690.450 104.400 ;
        RECT 698.400 103.350 699.600 105.600 ;
        RECT 703.950 105.000 706.050 109.050 ;
        RECT 716.400 105.600 717.450 175.800 ;
        RECT 719.400 139.200 720.450 175.950 ;
        RECT 721.950 175.800 724.050 177.900 ;
        RECT 728.400 176.400 729.600 178.650 ;
        RECT 728.400 172.050 729.450 176.400 ;
        RECT 733.950 175.950 736.050 178.050 ;
        RECT 737.400 177.450 738.450 182.400 ;
        RECT 746.400 181.350 747.600 183.600 ;
        RECT 752.400 181.350 753.600 183.600 ;
        RECT 757.950 181.950 760.050 184.050 ;
        RECT 763.950 181.950 766.050 184.050 ;
        RECT 767.400 183.600 768.450 187.950 ;
        RECT 767.400 181.500 768.600 183.600 ;
        RECT 742.950 178.950 745.050 181.050 ;
        RECT 745.950 178.950 748.050 181.050 ;
        RECT 748.950 178.950 751.050 181.050 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 760.950 179.100 763.050 181.200 ;
        RECT 766.950 179.100 769.050 181.200 ;
        RECT 769.950 179.100 772.050 181.200 ;
        RECT 737.400 176.400 741.450 177.450 ;
        RECT 743.400 177.000 744.600 178.650 ;
        RECT 749.400 177.900 750.600 178.650 ;
        RECT 761.400 178.050 762.600 178.800 ;
        RECT 727.950 169.950 730.050 172.050 ;
        RECT 734.400 154.050 735.450 175.950 ;
        RECT 736.950 169.950 739.050 175.050 ;
        RECT 736.950 157.950 739.050 160.050 ;
        RECT 733.950 151.950 736.050 154.050 ;
        RECT 730.950 146.400 733.050 148.500 ;
        RECT 718.950 137.100 721.050 139.200 ;
        RECT 724.950 137.100 727.050 139.200 ;
        RECT 725.400 136.350 726.600 137.100 ;
        RECT 724.950 133.950 727.050 136.050 ;
        RECT 721.950 130.950 724.050 133.050 ;
        RECT 722.400 127.050 723.450 130.950 ;
        RECT 721.950 124.950 724.050 127.050 ;
        RECT 731.100 126.600 732.300 146.400 ;
        RECT 734.400 138.450 735.600 138.600 ;
        RECT 737.400 138.450 738.450 157.950 ;
        RECT 734.400 137.400 738.450 138.450 ;
        RECT 734.400 136.350 735.600 137.400 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 740.400 130.050 741.450 176.400 ;
        RECT 742.950 172.950 745.050 177.000 ;
        RECT 748.950 175.800 751.050 177.900 ;
        RECT 760.950 175.950 763.050 178.050 ;
        RECT 770.400 176.400 771.600 178.800 ;
        RECT 770.400 172.050 771.450 176.400 ;
        RECT 776.400 175.050 777.450 187.950 ;
        RECT 791.400 187.050 792.450 223.950 ;
        RECT 794.400 199.050 795.450 241.950 ;
        RECT 797.400 226.050 798.450 253.950 ;
        RECT 806.400 250.050 807.450 254.400 ;
        RECT 808.950 253.950 811.050 256.050 ;
        RECT 815.400 255.900 816.600 256.650 ;
        RECT 805.950 247.950 808.050 250.050 ;
        RECT 796.950 223.950 799.050 226.050 ;
        RECT 799.950 215.100 802.050 217.200 ;
        RECT 800.400 214.350 801.600 215.100 ;
        RECT 799.950 211.950 802.050 214.050 ;
        RECT 802.950 211.950 805.050 214.050 ;
        RECT 803.400 210.900 804.600 211.650 ;
        RECT 802.950 208.800 805.050 210.900 ;
        RECT 809.400 205.050 810.450 253.950 ;
        RECT 814.950 253.800 817.050 255.900 ;
        RECT 811.950 247.950 814.050 250.050 ;
        RECT 812.400 217.050 813.450 247.950 ;
        RECT 818.700 246.600 819.900 266.400 ;
        RECT 824.400 264.450 825.450 331.950 ;
        RECT 827.400 268.050 828.450 343.950 ;
        RECT 830.400 340.200 831.450 346.950 ;
        RECT 835.950 343.950 838.050 346.050 ;
        RECT 829.950 338.100 832.050 340.200 ;
        RECT 836.400 339.600 837.450 343.950 ;
        RECT 845.400 340.050 846.450 409.950 ;
        RECT 848.400 343.050 849.450 415.950 ;
        RECT 853.950 376.950 856.050 379.050 ;
        RECT 850.950 346.950 853.050 349.050 ;
        RECT 847.950 340.950 850.050 343.050 ;
        RECT 836.400 337.500 837.600 339.600 ;
        RECT 844.950 337.950 847.050 340.050 ;
        RECT 851.400 339.600 852.450 346.950 ;
        RECT 854.400 343.050 855.450 376.950 ;
        RECT 857.400 373.050 858.450 514.800 ;
        RECT 860.400 418.050 861.450 532.950 ;
        RECT 859.950 415.950 862.050 418.050 ;
        RECT 863.400 375.450 864.450 583.950 ;
        RECT 860.400 374.400 864.450 375.450 ;
        RECT 856.950 370.950 859.050 373.050 ;
        RECT 853.950 340.950 856.050 343.050 ;
        RECT 851.400 337.500 852.600 339.600 ;
        RECT 832.950 335.100 835.050 337.200 ;
        RECT 835.950 335.100 838.050 337.200 ;
        RECT 838.950 335.100 841.050 337.200 ;
        RECT 847.950 335.100 850.050 337.200 ;
        RECT 850.950 335.100 853.050 337.200 ;
        RECT 853.950 335.100 856.050 337.200 ;
        RECT 833.400 334.050 834.600 334.800 ;
        RECT 832.950 331.950 835.050 334.050 ;
        RECT 839.400 332.400 840.600 334.800 ;
        RECT 832.950 325.950 835.050 328.050 ;
        RECT 833.400 294.600 834.450 325.950 ;
        RECT 839.400 301.050 840.450 332.400 ;
        RECT 841.950 331.950 844.050 334.050 ;
        RECT 848.400 332.400 849.600 334.800 ;
        RECT 854.400 334.050 855.600 334.800 ;
        RECT 838.950 298.950 841.050 301.050 ;
        RECT 842.400 297.450 843.450 331.950 ;
        RECT 848.400 319.050 849.450 332.400 ;
        RECT 853.950 331.950 856.050 334.050 ;
        RECT 850.950 328.950 853.050 331.050 ;
        RECT 847.950 316.950 850.050 319.050 ;
        RECT 839.400 296.400 843.450 297.450 ;
        RECT 839.400 294.600 840.450 296.400 ;
        RECT 833.400 292.350 834.600 294.600 ;
        RECT 839.400 292.350 840.600 294.600 ;
        RECT 832.950 289.950 835.050 292.050 ;
        RECT 835.950 289.950 838.050 292.050 ;
        RECT 838.950 289.950 841.050 292.050 ;
        RECT 841.950 289.950 844.050 292.050 ;
        RECT 829.950 286.800 832.050 288.900 ;
        RECT 836.400 287.400 837.600 289.650 ;
        RECT 842.400 288.900 843.600 289.650 ;
        RECT 826.950 265.950 829.050 268.050 ;
        RECT 824.400 264.000 828.450 264.450 ;
        RECT 824.400 263.400 829.050 264.000 ;
        RECT 826.950 259.950 829.050 263.400 ;
        RECT 823.950 256.950 826.050 259.050 ;
        RECT 820.950 253.950 823.050 256.050 ;
        RECT 824.400 255.000 825.600 256.650 ;
        RECT 821.400 250.050 822.450 253.950 ;
        RECT 823.950 250.950 826.050 255.000 ;
        RECT 826.950 253.950 829.050 256.050 ;
        RECT 820.950 247.950 823.050 250.050 ;
        RECT 817.950 244.500 820.050 246.600 ;
        RECT 827.400 244.050 828.450 253.950 ;
        RECT 826.950 241.950 829.050 244.050 ;
        RECT 830.400 241.050 831.450 286.800 ;
        RECT 836.400 273.450 837.450 287.400 ;
        RECT 841.950 286.800 844.050 288.900 ;
        RECT 833.400 272.400 837.450 273.450 ;
        RECT 833.400 253.050 834.450 272.400 ;
        RECT 838.950 266.400 841.050 268.500 ;
        RECT 832.950 250.950 835.050 253.050 ;
        RECT 838.950 251.400 840.150 266.400 ;
        RECT 847.950 265.950 850.050 268.050 ;
        RECT 841.950 260.100 844.050 262.200 ;
        RECT 842.400 259.350 843.600 260.100 ;
        RECT 841.950 256.950 844.050 259.050 ;
        RECT 838.950 249.300 841.050 251.400 ;
        RECT 838.950 245.700 840.150 249.300 ;
        RECT 838.950 243.600 841.050 245.700 ;
        RECT 829.950 238.950 832.050 241.050 ;
        RECT 820.950 229.950 823.050 232.050 ;
        RECT 826.950 229.950 829.050 232.050 ;
        RECT 814.950 223.950 817.050 226.050 ;
        RECT 811.950 214.950 814.050 217.050 ;
        RECT 815.400 216.600 816.450 223.950 ;
        RECT 821.400 216.600 822.450 229.950 ;
        RECT 815.400 214.200 816.600 216.600 ;
        RECT 821.400 214.200 822.600 216.600 ;
        RECT 814.950 211.800 817.050 213.900 ;
        RECT 817.950 211.800 820.050 213.900 ;
        RECT 820.950 211.800 823.050 213.900 ;
        RECT 818.400 210.750 819.600 211.500 ;
        RECT 817.950 208.650 820.050 210.750 ;
        RECT 808.950 202.950 811.050 205.050 ;
        RECT 793.950 196.950 796.050 199.050 ;
        RECT 814.950 196.950 817.050 199.050 ;
        RECT 793.950 187.950 796.050 190.050 ;
        RECT 802.950 188.400 805.050 190.500 ;
        RECT 778.950 182.100 781.050 184.200 ;
        RECT 772.950 172.950 775.050 175.050 ;
        RECT 775.950 172.950 778.050 175.050 ;
        RECT 744.000 171.900 747.000 172.050 ;
        RECT 742.950 169.950 748.050 171.900 ;
        RECT 769.950 169.950 772.050 172.050 ;
        RECT 742.950 169.800 745.050 169.950 ;
        RECT 745.950 169.800 748.050 169.950 ;
        RECT 773.400 166.050 774.450 172.950 ;
        RECT 779.400 169.050 780.450 182.100 ;
        RECT 781.950 181.950 784.050 187.050 ;
        RECT 790.950 184.950 793.050 187.050 ;
        RECT 787.950 182.100 790.050 184.200 ;
        RECT 794.400 183.600 795.450 187.950 ;
        RECT 788.400 181.350 789.600 182.100 ;
        RECT 794.400 181.350 795.600 183.600 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 793.950 178.950 796.050 181.050 ;
        RECT 799.950 178.950 802.050 181.050 ;
        RECT 781.950 175.950 784.050 178.050 ;
        RECT 785.400 177.000 786.600 178.650 ;
        RECT 778.950 166.950 781.050 169.050 ;
        RECT 772.950 163.950 775.050 166.050 ;
        RECT 766.950 151.950 769.050 154.050 ;
        RECT 751.950 138.000 754.050 142.050 ;
        RECT 757.950 139.950 760.050 142.050 ;
        RECT 752.400 136.350 753.600 138.000 ;
        RECT 745.950 133.950 748.050 136.050 ;
        RECT 751.950 133.950 754.050 136.050 ;
        RECT 746.400 132.000 747.600 133.650 ;
        RECT 739.950 127.950 742.050 130.050 ;
        RECT 745.950 127.950 748.050 132.000 ;
        RECT 758.400 130.050 759.450 139.950 ;
        RECT 767.400 138.600 768.450 151.950 ;
        RECT 767.400 136.350 768.600 138.600 ;
        RECT 772.950 137.100 775.050 139.200 ;
        RECT 778.950 137.100 781.050 139.200 ;
        RECT 773.400 136.350 774.600 137.100 ;
        RECT 763.950 133.950 766.050 136.050 ;
        RECT 766.950 133.950 769.050 136.050 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 764.400 132.000 765.600 133.650 ;
        RECT 751.950 127.950 754.050 130.050 ;
        RECT 757.950 127.950 760.050 130.050 ;
        RECT 763.950 127.950 766.050 132.000 ;
        RECT 770.400 131.400 771.600 133.650 ;
        RECT 779.400 133.050 780.450 137.100 ;
        RECT 730.950 124.500 733.050 126.600 ;
        RECT 745.950 110.400 748.050 112.500 ;
        RECT 704.400 103.350 705.600 105.000 ;
        RECT 716.400 103.500 717.600 105.600 ;
        RECT 737.400 105.450 738.600 105.600 ;
        RECT 743.400 105.450 744.600 105.600 ;
        RECT 737.400 104.400 744.600 105.450 ;
        RECT 737.400 103.350 738.600 104.400 ;
        RECT 743.400 103.350 744.600 104.400 ;
        RECT 694.950 100.950 697.050 103.050 ;
        RECT 697.950 100.950 700.050 103.050 ;
        RECT 700.950 100.950 703.050 103.050 ;
        RECT 703.950 100.950 706.050 103.050 ;
        RECT 712.950 101.100 715.050 103.200 ;
        RECT 715.950 101.100 718.050 103.200 ;
        RECT 718.950 101.100 721.050 103.200 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 742.950 100.950 745.050 103.050 ;
        RECT 695.400 98.400 696.600 100.650 ;
        RECT 701.400 98.400 702.600 100.650 ;
        RECT 713.400 98.400 714.600 100.800 ;
        RECT 719.400 100.050 720.600 100.800 ;
        RECT 688.950 82.950 691.050 85.050 ;
        RECT 695.400 79.050 696.450 98.400 ;
        RECT 701.400 88.050 702.450 98.400 ;
        RECT 700.950 85.950 703.050 88.050 ;
        RECT 694.950 76.950 697.050 79.050 ;
        RECT 691.950 67.950 694.050 70.050 ;
        RECT 697.950 67.950 700.050 70.050 ;
        RECT 683.400 65.400 687.450 66.450 ;
        RECT 676.950 63.450 679.050 64.050 ;
        RECT 641.400 63.000 648.450 63.450 ;
        RECT 668.400 63.000 679.050 63.450 ;
        RECT 641.400 62.400 649.050 63.000 ;
        RECT 634.950 58.950 637.050 61.050 ;
        RECT 641.400 60.600 642.450 62.400 ;
        RECT 641.400 58.350 642.600 60.600 ;
        RECT 646.950 58.950 649.050 62.400 ;
        RECT 667.950 62.400 679.050 63.000 ;
        RECT 667.950 58.950 670.050 62.400 ;
        RECT 676.950 61.950 679.050 62.400 ;
        RECT 673.950 59.100 676.050 61.200 ;
        RECT 680.400 61.050 681.450 64.950 ;
        RECT 674.400 58.350 675.600 59.100 ;
        RECT 679.950 58.950 682.050 61.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 652.950 55.950 655.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 670.950 55.950 673.050 58.050 ;
        RECT 673.950 55.950 676.050 58.050 ;
        RECT 676.950 55.950 679.050 58.050 ;
        RECT 634.950 52.950 637.050 55.050 ;
        RECT 638.400 54.000 639.600 55.650 ;
        RECT 644.400 54.900 645.600 55.650 ;
        RECT 635.400 49.050 636.450 52.950 ;
        RECT 637.950 49.950 640.050 54.000 ;
        RECT 643.950 52.800 646.050 54.900 ;
        RECT 653.400 53.400 654.600 55.650 ;
        RECT 634.950 46.950 637.050 49.050 ;
        RECT 643.950 46.950 646.050 49.050 ;
        RECT 631.950 37.950 634.050 40.050 ;
        RECT 592.950 34.950 595.050 37.050 ;
        RECT 598.950 34.950 601.050 37.050 ;
        RECT 565.950 25.950 568.050 28.050 ;
        RECT 574.950 26.250 577.050 28.350 ;
        RECT 566.400 22.050 567.450 25.950 ;
        RECT 575.400 25.500 576.600 26.250 ;
        RECT 580.950 25.950 583.050 31.050 ;
        RECT 599.400 28.200 600.450 34.950 ;
        RECT 607.950 32.400 610.050 34.500 ;
        RECT 628.950 32.400 631.050 34.500 ;
        RECT 583.950 26.100 586.050 28.200 ;
        RECT 592.950 26.100 595.050 28.200 ;
        RECT 598.950 26.100 601.050 28.200 ;
        RECT 571.950 23.100 574.050 25.200 ;
        RECT 574.950 23.100 577.050 25.200 ;
        RECT 577.950 23.100 580.050 25.200 ;
        RECT 572.400 22.050 573.600 22.800 ;
        RECT 578.400 22.050 579.600 22.800 ;
        RECT 556.950 19.800 559.050 21.900 ;
        RECT 562.950 19.800 565.050 21.900 ;
        RECT 565.950 19.950 568.050 22.050 ;
        RECT 571.950 19.950 574.050 22.050 ;
        RECT 577.950 19.950 580.050 22.050 ;
        RECT 584.400 13.050 585.450 26.100 ;
        RECT 593.400 25.350 594.600 26.100 ;
        RECT 599.400 25.350 600.600 26.100 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 592.950 22.950 595.050 25.050 ;
        RECT 595.950 22.950 598.050 25.050 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 590.400 22.050 591.600 22.650 ;
        RECT 586.950 20.400 591.600 22.050 ;
        RECT 596.400 21.900 597.600 22.650 ;
        RECT 586.950 19.950 591.000 20.400 ;
        RECT 595.950 19.800 598.050 21.900 ;
        RECT 605.400 21.000 606.600 22.650 ;
        RECT 604.950 16.950 607.050 21.000 ;
        RECT 553.950 10.500 556.050 12.600 ;
        RECT 583.950 10.950 586.050 13.050 ;
        RECT 608.700 12.600 609.900 32.400 ;
        RECT 613.950 22.950 616.050 25.050 ;
        RECT 614.400 20.400 615.600 22.650 ;
        RECT 614.400 13.050 615.450 20.400 ;
        RECT 628.950 17.400 630.150 32.400 ;
        RECT 631.950 26.100 634.050 28.200 ;
        RECT 644.400 27.600 645.450 46.950 ;
        RECT 653.400 40.050 654.450 53.400 ;
        RECT 667.950 52.950 670.050 55.050 ;
        RECT 671.400 53.400 672.600 55.650 ;
        RECT 677.400 54.900 678.600 55.650 ;
        RECT 668.400 49.050 669.450 52.950 ;
        RECT 667.950 46.950 670.050 49.050 ;
        RECT 652.950 37.950 655.050 40.050 ;
        RECT 632.400 25.350 633.600 26.100 ;
        RECT 644.400 25.350 645.600 27.600 ;
        RECT 661.950 26.100 664.050 28.200 ;
        RECT 662.400 25.350 663.600 26.100 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 649.950 22.950 652.050 25.050 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 664.950 22.950 667.050 25.050 ;
        RECT 665.400 21.900 666.600 22.650 ;
        RECT 671.400 21.900 672.450 53.400 ;
        RECT 676.950 52.800 679.050 54.900 ;
        RECT 676.950 26.100 679.050 28.200 ;
        RECT 683.400 27.600 684.450 65.400 ;
        RECT 685.950 58.950 688.050 64.050 ;
        RECT 692.400 60.600 693.450 67.950 ;
        RECT 692.400 58.350 693.600 60.600 ;
        RECT 698.400 60.450 699.450 67.950 ;
        RECT 701.400 64.050 702.450 85.950 ;
        RECT 713.400 85.050 714.450 98.400 ;
        RECT 718.950 97.950 721.050 100.050 ;
        RECT 734.400 98.400 735.600 100.650 ;
        RECT 734.400 88.050 735.450 98.400 ;
        RECT 746.850 95.400 748.050 110.400 ;
        RECT 752.400 100.050 753.450 127.950 ;
        RECT 770.400 121.050 771.450 131.400 ;
        RECT 778.950 130.950 781.050 133.050 ;
        RECT 757.950 118.950 760.050 121.050 ;
        RECT 769.950 118.950 772.050 121.050 ;
        RECT 758.400 106.050 759.450 118.950 ;
        RECT 760.950 108.450 763.050 112.050 ;
        RECT 766.950 110.400 769.050 112.500 ;
        RECT 760.950 108.000 765.450 108.450 ;
        RECT 761.400 107.400 766.050 108.000 ;
        RECT 757.950 103.950 760.050 106.050 ;
        RECT 763.950 103.950 766.050 107.400 ;
        RECT 760.950 100.950 763.050 103.050 ;
        RECT 761.400 100.050 762.600 100.650 ;
        RECT 751.950 97.950 754.050 100.050 ;
        RECT 757.950 97.950 760.050 100.050 ;
        RECT 761.400 98.400 766.050 100.050 ;
        RECT 762.000 97.950 766.050 98.400 ;
        RECT 745.950 93.300 748.050 95.400 ;
        RECT 746.850 89.700 748.050 93.300 ;
        RECT 733.950 85.950 736.050 88.050 ;
        RECT 745.950 87.600 748.050 89.700 ;
        RECT 712.950 82.950 715.050 85.050 ;
        RECT 752.400 76.050 753.450 97.950 ;
        RECT 758.400 88.050 759.450 97.950 ;
        RECT 760.950 94.950 763.050 97.050 ;
        RECT 757.950 85.950 760.050 88.050 ;
        RECT 751.950 73.950 754.050 76.050 ;
        RECT 718.950 67.950 721.050 70.050 ;
        RECT 700.950 61.950 703.050 64.050 ;
        RECT 698.400 59.400 702.450 60.450 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 691.950 55.950 694.050 58.050 ;
        RECT 694.950 55.950 697.050 58.050 ;
        RECT 689.400 53.400 690.600 55.650 ;
        RECT 695.400 53.400 696.600 55.650 ;
        RECT 677.400 25.350 678.600 26.100 ;
        RECT 683.400 25.350 684.600 27.600 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 680.400 21.900 681.600 22.650 ;
        RECT 689.400 22.050 690.450 53.400 ;
        RECT 695.400 49.050 696.450 53.400 ;
        RECT 694.950 46.950 697.050 49.050 ;
        RECT 701.400 40.050 702.450 59.400 ;
        RECT 703.950 58.950 706.050 61.050 ;
        RECT 712.950 58.950 715.050 61.050 ;
        RECT 719.400 60.600 720.450 67.950 ;
        RECT 761.400 67.050 762.450 94.950 ;
        RECT 767.100 90.600 768.300 110.400 ;
        RECT 782.400 109.200 783.450 175.950 ;
        RECT 784.950 172.950 787.050 177.000 ;
        RECT 791.400 176.400 792.600 178.650 ;
        RECT 800.400 176.400 801.600 178.650 ;
        RECT 787.950 172.950 790.050 175.050 ;
        RECT 791.400 174.450 792.450 176.400 ;
        RECT 791.400 173.400 795.450 174.450 ;
        RECT 788.400 142.050 789.450 172.950 ;
        RECT 790.950 169.950 793.050 172.050 ;
        RECT 791.400 160.050 792.450 169.950 ;
        RECT 794.400 163.050 795.450 173.400 ;
        RECT 800.400 172.050 801.450 176.400 ;
        RECT 799.950 169.950 802.050 172.050 ;
        RECT 803.700 168.600 804.900 188.400 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 809.400 176.400 810.600 178.650 ;
        RECT 809.400 169.050 810.450 176.400 ;
        RECT 815.400 175.050 816.450 196.950 ;
        RECT 827.400 196.050 828.450 229.950 ;
        RECT 848.400 220.050 849.450 265.950 ;
        RECT 851.400 262.200 852.450 328.950 ;
        RECT 860.400 303.450 861.450 374.400 ;
        RECT 862.950 370.950 865.050 373.050 ;
        RECT 857.400 302.400 861.450 303.450 ;
        RECT 850.950 260.100 853.050 262.200 ;
        RECT 851.400 226.050 852.450 260.100 ;
        RECT 857.400 232.050 858.450 302.400 ;
        RECT 859.950 298.950 862.050 301.050 ;
        RECT 856.950 229.950 859.050 232.050 ;
        RECT 850.950 223.950 853.050 226.050 ;
        RECT 832.950 216.000 835.050 220.050 ;
        RECT 847.950 217.950 850.050 220.050 ;
        RECT 833.400 214.350 834.600 216.000 ;
        RECT 838.950 215.100 841.050 217.200 ;
        RECT 856.950 215.100 859.050 217.200 ;
        RECT 839.400 214.350 840.600 215.100 ;
        RECT 832.950 211.950 835.050 214.050 ;
        RECT 835.950 211.950 838.050 214.050 ;
        RECT 838.950 211.950 841.050 214.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 836.400 209.400 837.600 211.650 ;
        RECT 842.400 210.900 843.600 211.650 ;
        RECT 826.950 193.950 829.050 196.050 ;
        RECT 823.950 188.400 826.050 190.500 ;
        RECT 817.950 178.950 820.050 181.050 ;
        RECT 814.950 172.950 817.050 175.050 ;
        RECT 802.950 166.500 805.050 168.600 ;
        RECT 808.950 166.950 811.050 169.050 ;
        RECT 793.950 160.950 796.050 163.050 ;
        RECT 790.950 157.950 793.050 160.050 ;
        RECT 791.400 148.050 792.450 157.950 ;
        RECT 818.400 151.050 819.450 178.950 ;
        RECT 823.950 173.400 825.150 188.400 ;
        RECT 826.950 182.100 829.050 184.200 ;
        RECT 836.400 183.450 837.450 209.400 ;
        RECT 841.950 208.800 844.050 210.900 ;
        RECT 853.950 208.800 856.050 210.900 ;
        RECT 838.950 193.950 841.050 196.050 ;
        RECT 839.400 184.200 840.450 193.950 ;
        RECT 833.400 182.400 837.450 183.450 ;
        RECT 827.400 181.350 828.600 182.100 ;
        RECT 826.950 178.950 829.050 181.050 ;
        RECT 823.950 171.300 826.050 173.400 ;
        RECT 823.950 167.700 825.150 171.300 ;
        RECT 823.950 165.600 826.050 167.700 ;
        RECT 817.950 148.950 820.050 151.050 ;
        RECT 790.950 145.950 793.050 148.050 ;
        RECT 787.950 138.000 790.050 142.050 ;
        RECT 796.950 139.050 799.050 139.200 ;
        RECT 795.000 138.600 799.050 139.050 ;
        RECT 788.400 136.200 789.600 138.000 ;
        RECT 794.400 137.100 799.050 138.600 ;
        RECT 805.950 137.100 808.050 139.200 ;
        RECT 811.950 138.000 814.050 142.050 ;
        RECT 818.400 139.050 819.450 148.950 ;
        RECT 823.950 147.300 826.050 149.400 ;
        RECT 824.850 143.700 826.050 147.300 ;
        RECT 823.950 141.600 826.050 143.700 ;
        RECT 794.400 136.950 798.000 137.100 ;
        RECT 794.400 136.200 795.600 136.950 ;
        RECT 806.400 136.350 807.600 137.100 ;
        RECT 812.400 136.350 813.600 138.000 ;
        RECT 817.950 136.950 820.050 139.050 ;
        RECT 787.950 133.800 790.050 135.900 ;
        RECT 790.950 133.800 793.050 135.900 ;
        RECT 793.950 133.800 796.050 135.900 ;
        RECT 802.950 133.950 805.050 136.050 ;
        RECT 805.950 133.950 808.050 136.050 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 820.950 133.950 823.050 136.050 ;
        RECT 791.400 132.750 792.600 133.500 ;
        RECT 790.950 130.650 793.050 132.750 ;
        RECT 803.400 131.400 804.600 133.650 ;
        RECT 809.400 132.000 810.600 133.650 ;
        RECT 787.950 129.450 790.050 130.050 ;
        RECT 793.950 129.450 796.050 130.050 ;
        RECT 787.950 128.400 796.050 129.450 ;
        RECT 787.950 127.950 790.050 128.400 ;
        RECT 793.950 127.950 796.050 128.400 ;
        RECT 787.950 121.950 790.050 124.050 ;
        RECT 775.950 106.950 778.050 109.050 ;
        RECT 781.950 107.100 784.050 109.200 ;
        RECT 769.950 100.950 772.050 103.050 ;
        RECT 770.400 99.000 771.600 100.650 ;
        RECT 769.950 94.950 772.050 99.000 ;
        RECT 776.400 91.050 777.450 106.950 ;
        RECT 781.950 103.950 784.050 106.050 ;
        RECT 788.400 105.600 789.450 121.950 ;
        RECT 803.400 115.050 804.450 131.400 ;
        RECT 808.950 127.950 811.050 132.000 ;
        RECT 814.950 130.950 817.050 133.050 ;
        RECT 821.400 132.900 822.600 133.650 ;
        RECT 805.950 121.950 808.050 124.050 ;
        RECT 802.950 114.450 805.050 115.050 ;
        RECT 800.400 113.400 805.050 114.450 ;
        RECT 796.950 106.950 799.050 109.050 ;
        RECT 782.400 103.350 783.600 103.950 ;
        RECT 788.400 103.350 789.600 105.600 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 784.950 100.950 787.050 103.050 ;
        RECT 787.950 100.950 790.050 103.050 ;
        RECT 790.950 100.950 793.050 103.050 ;
        RECT 778.950 97.950 781.050 100.050 ;
        RECT 785.400 98.400 786.600 100.650 ;
        RECT 791.400 98.400 792.600 100.650 ;
        RECT 766.950 88.500 769.050 90.600 ;
        RECT 775.950 88.950 778.050 91.050 ;
        RECT 779.400 82.050 780.450 97.950 ;
        RECT 785.400 96.450 786.450 98.400 ;
        RECT 782.400 95.400 786.450 96.450 ;
        RECT 766.950 79.950 769.050 82.050 ;
        RECT 778.950 79.950 781.050 82.050 ;
        RECT 760.950 64.950 763.050 67.050 ;
        RECT 767.400 61.200 768.450 79.950 ;
        RECT 772.950 73.950 775.050 76.050 ;
        RECT 704.400 49.050 705.450 58.950 ;
        RECT 713.400 58.200 714.600 58.950 ;
        RECT 719.400 58.200 720.600 60.600 ;
        RECT 730.950 59.100 733.050 61.200 ;
        RECT 731.400 58.350 732.600 59.100 ;
        RECT 736.950 58.950 739.050 61.050 ;
        RECT 742.950 58.950 745.050 61.050 ;
        RECT 751.950 58.950 754.050 61.050 ;
        RECT 757.950 58.950 760.050 61.050 ;
        RECT 766.950 59.100 769.050 61.200 ;
        RECT 709.950 55.800 712.050 57.900 ;
        RECT 712.950 55.800 715.050 57.900 ;
        RECT 715.950 55.800 718.050 57.900 ;
        RECT 718.950 55.800 721.050 57.900 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 730.950 55.950 733.050 58.050 ;
        RECT 710.400 53.400 711.600 55.500 ;
        RECT 716.400 54.750 717.600 55.500 ;
        RECT 728.400 54.900 729.600 55.650 ;
        RECT 703.950 46.950 706.050 49.050 ;
        RECT 700.950 37.950 703.050 40.050 ;
        RECT 710.400 28.200 711.450 53.400 ;
        RECT 715.950 52.650 718.050 54.750 ;
        RECT 727.950 52.800 730.050 54.900 ;
        RECT 730.950 37.950 733.050 40.050 ;
        RECT 712.950 31.950 715.050 34.050 ;
        RECT 718.950 31.950 721.050 34.050 ;
        RECT 700.950 26.100 703.050 28.200 ;
        RECT 709.950 26.100 712.050 28.200 ;
        RECT 713.400 27.600 714.450 31.950 ;
        RECT 719.400 27.600 720.450 31.950 ;
        RECT 731.400 27.600 732.450 37.950 ;
        RECT 737.400 28.050 738.450 58.950 ;
        RECT 743.400 58.200 744.600 58.950 ;
        RECT 752.400 58.200 753.600 58.950 ;
        RECT 742.950 55.800 745.050 57.900 ;
        RECT 748.950 55.800 751.050 57.900 ;
        RECT 751.950 55.800 754.050 57.900 ;
        RECT 749.400 53.400 750.600 55.500 ;
        RECT 749.400 43.050 750.450 53.400 ;
        RECT 748.950 40.950 751.050 43.050 ;
        RECT 758.400 36.450 759.450 58.950 ;
        RECT 767.400 58.350 768.600 59.100 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 764.400 54.900 765.600 55.650 ;
        RECT 763.950 52.800 766.050 54.900 ;
        RECT 764.400 43.050 765.450 52.800 ;
        RECT 766.950 49.950 769.050 52.050 ;
        RECT 763.950 40.950 766.050 43.050 ;
        RECT 758.400 35.400 762.450 36.450 ;
        RECT 748.950 31.950 754.050 34.050 ;
        RECT 757.950 31.950 760.050 34.050 ;
        RECT 701.400 25.350 702.600 26.100 ;
        RECT 713.400 25.500 714.600 27.600 ;
        RECT 719.400 25.500 720.600 27.600 ;
        RECT 731.400 25.350 732.600 27.600 ;
        RECT 736.950 25.950 739.050 28.050 ;
        RECT 739.950 26.100 742.050 28.200 ;
        RECT 745.950 26.100 748.050 28.200 ;
        RECT 751.950 27.000 754.050 30.900 ;
        RECT 697.950 22.950 700.050 25.050 ;
        RECT 700.950 22.950 703.050 25.050 ;
        RECT 712.950 23.100 715.050 25.200 ;
        RECT 715.950 23.100 718.050 25.200 ;
        RECT 718.950 23.100 721.050 25.200 ;
        RECT 721.950 23.100 724.050 25.200 ;
        RECT 730.950 22.950 733.050 25.050 ;
        RECT 733.950 22.950 736.050 25.050 ;
        RECT 664.950 19.800 667.050 21.900 ;
        RECT 670.950 19.800 673.050 21.900 ;
        RECT 679.950 19.800 682.050 21.900 ;
        RECT 688.950 19.950 691.050 22.050 ;
        RECT 698.400 21.900 699.600 22.650 ;
        RECT 716.400 22.050 717.600 22.800 ;
        RECT 722.400 22.050 723.600 22.800 ;
        RECT 697.950 19.800 700.050 21.900 ;
        RECT 715.950 19.950 718.050 22.050 ;
        RECT 721.950 19.950 724.050 22.050 ;
        RECT 734.400 21.900 735.600 22.650 ;
        RECT 740.400 22.050 741.450 26.100 ;
        RECT 746.400 25.350 747.600 26.100 ;
        RECT 752.400 25.350 753.600 27.000 ;
        RECT 745.950 22.950 748.050 25.050 ;
        RECT 748.950 22.950 751.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 733.950 19.800 736.050 21.900 ;
        RECT 739.950 19.950 742.050 22.050 ;
        RECT 742.950 19.950 745.050 22.050 ;
        RECT 749.400 21.900 750.600 22.650 ;
        RECT 758.400 22.050 759.450 31.950 ;
        RECT 761.400 31.050 762.450 35.400 ;
        RECT 767.400 34.050 768.450 49.950 ;
        RECT 773.400 34.050 774.450 73.950 ;
        RECT 782.400 61.200 783.450 95.400 ;
        RECT 791.400 91.050 792.450 98.400 ;
        RECT 790.950 88.950 793.050 91.050 ;
        RECT 797.400 76.050 798.450 106.950 ;
        RECT 800.400 106.050 801.450 113.400 ;
        RECT 802.950 112.950 805.050 113.400 ;
        RECT 799.950 103.950 802.050 106.050 ;
        RECT 806.400 105.600 807.450 121.950 ;
        RECT 806.400 103.500 807.600 105.600 ;
        RECT 815.400 105.450 816.450 130.950 ;
        RECT 820.950 130.800 823.050 132.900 ;
        RECT 824.850 126.600 826.050 141.600 ;
        RECT 829.950 139.950 832.050 142.050 ;
        RECT 823.950 124.500 826.050 126.600 ;
        RECT 830.400 124.050 831.450 139.950 ;
        RECT 833.400 139.200 834.450 182.400 ;
        RECT 838.950 182.100 841.050 184.200 ;
        RECT 839.400 181.350 840.600 182.100 ;
        RECT 838.950 178.950 841.050 181.050 ;
        RECT 841.950 178.950 844.050 181.050 ;
        RECT 842.400 176.400 843.600 178.650 ;
        RECT 842.400 163.050 843.450 176.400 ;
        RECT 841.950 160.950 844.050 163.050 ;
        RECT 844.950 146.400 847.050 148.500 ;
        RECT 832.950 137.100 835.050 139.200 ;
        RECT 838.950 137.100 841.050 139.200 ;
        RECT 839.400 136.350 840.600 137.100 ;
        RECT 838.950 133.950 841.050 136.050 ;
        RECT 845.100 126.600 846.300 146.400 ;
        RECT 847.950 142.950 850.050 145.050 ;
        RECT 848.400 139.200 849.450 142.950 ;
        RECT 847.950 137.100 850.050 139.200 ;
        RECT 848.400 136.350 849.600 137.100 ;
        RECT 847.950 133.950 850.050 136.050 ;
        RECT 850.950 130.950 853.050 133.050 ;
        RECT 844.950 124.500 847.050 126.600 ;
        RECT 829.950 121.950 832.050 124.050 ;
        RECT 820.950 110.400 823.050 112.500 ;
        RECT 841.950 110.400 844.050 112.500 ;
        RECT 818.400 105.450 819.600 105.600 ;
        RECT 815.400 104.400 819.600 105.450 ;
        RECT 818.400 103.350 819.600 104.400 ;
        RECT 802.950 101.100 805.050 103.200 ;
        RECT 805.950 101.100 808.050 103.200 ;
        RECT 808.950 101.100 811.050 103.200 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 803.400 100.050 804.600 100.800 ;
        RECT 802.950 97.950 805.050 100.050 ;
        RECT 809.400 98.400 810.600 100.800 ;
        RECT 809.400 85.050 810.450 98.400 ;
        RECT 814.950 97.800 817.050 99.900 ;
        RECT 815.400 88.050 816.450 97.800 ;
        RECT 821.850 95.400 823.050 110.400 ;
        RECT 835.950 100.950 838.050 103.050 ;
        RECT 836.400 99.900 837.600 100.650 ;
        RECT 835.950 97.800 838.050 99.900 ;
        RECT 820.950 93.300 823.050 95.400 ;
        RECT 821.850 89.700 823.050 93.300 ;
        RECT 842.100 90.600 843.300 110.400 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 845.400 99.450 846.600 100.650 ;
        RECT 851.400 99.450 852.450 130.950 ;
        RECT 845.400 98.400 852.450 99.450 ;
        RECT 847.950 94.950 850.050 97.050 ;
        RECT 814.950 85.950 817.050 88.050 ;
        RECT 820.950 87.600 823.050 89.700 ;
        RECT 841.950 88.500 844.050 90.600 ;
        RECT 808.950 82.950 811.050 85.050 ;
        RECT 823.950 82.950 826.050 85.050 ;
        RECT 796.950 73.950 799.050 76.050 ;
        RECT 808.950 73.950 811.050 76.050 ;
        RECT 793.950 68.400 796.050 70.500 ;
        RECT 790.950 64.950 793.050 67.050 ;
        RECT 775.950 58.950 778.050 61.050 ;
        RECT 781.950 59.100 784.050 61.200 ;
        RECT 791.400 60.600 792.450 64.950 ;
        RECT 766.950 31.950 769.050 34.050 ;
        RECT 772.950 31.950 775.050 34.050 ;
        RECT 776.400 33.450 777.450 58.950 ;
        RECT 782.400 58.350 783.600 59.100 ;
        RECT 791.400 58.350 792.600 60.600 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 790.950 55.950 793.050 58.050 ;
        RECT 785.400 54.000 786.600 55.650 ;
        RECT 784.950 49.950 787.050 54.000 ;
        RECT 794.700 48.600 795.900 68.400 ;
        RECT 799.950 59.100 802.050 61.200 ;
        RECT 805.950 59.100 808.050 61.200 ;
        RECT 800.400 58.350 801.600 59.100 ;
        RECT 799.950 55.950 802.050 58.050 ;
        RECT 793.950 46.500 796.050 48.600 ;
        RECT 806.400 40.050 807.450 59.100 ;
        RECT 809.400 52.050 810.450 73.950 ;
        RECT 814.950 69.300 817.050 71.400 ;
        RECT 814.950 65.700 816.150 69.300 ;
        RECT 814.950 63.600 817.050 65.700 ;
        RECT 808.950 49.950 811.050 52.050 ;
        RECT 814.950 48.600 816.150 63.600 ;
        RECT 824.400 61.200 825.450 82.950 ;
        RECT 823.950 59.100 826.050 61.200 ;
        RECT 832.950 59.100 835.050 61.200 ;
        RECT 848.400 60.600 849.450 94.950 ;
        RECT 851.400 67.050 852.450 98.400 ;
        RECT 854.400 97.050 855.450 208.800 ;
        RECT 857.400 127.050 858.450 215.100 ;
        RECT 860.400 151.050 861.450 298.950 ;
        RECT 863.400 289.050 864.450 370.950 ;
        RECT 862.950 286.950 865.050 289.050 ;
        RECT 859.950 148.950 862.050 151.050 ;
        RECT 856.950 124.950 859.050 127.050 ;
        RECT 853.950 94.950 856.050 97.050 ;
        RECT 850.950 64.950 853.050 67.050 ;
        RECT 817.950 55.950 820.050 58.050 ;
        RECT 818.400 54.900 819.600 55.650 ;
        RECT 817.950 52.800 820.050 54.900 ;
        RECT 824.400 54.450 825.450 59.100 ;
        RECT 833.400 58.350 834.600 59.100 ;
        RECT 848.400 58.350 849.600 60.600 ;
        RECT 829.950 55.950 832.050 58.050 ;
        RECT 832.950 55.950 835.050 58.050 ;
        RECT 844.950 55.950 847.050 58.050 ;
        RECT 847.950 55.950 850.050 58.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 830.400 54.900 831.600 55.650 ;
        RECT 821.400 53.400 825.450 54.450 ;
        RECT 814.950 46.500 817.050 48.600 ;
        RECT 805.950 37.950 808.050 40.050 ;
        RECT 817.950 37.950 820.050 40.050 ;
        RECT 776.400 32.400 780.450 33.450 ;
        RECT 760.950 30.450 763.050 31.050 ;
        RECT 760.950 29.400 777.450 30.450 ;
        RECT 760.950 28.950 763.050 29.400 ;
        RECT 760.950 25.800 763.050 27.900 ;
        RECT 769.950 26.100 772.050 28.200 ;
        RECT 776.400 27.600 777.450 29.400 ;
        RECT 779.400 28.050 780.450 32.400 ;
        RECT 814.950 31.950 817.050 34.050 ;
        RECT 628.950 15.300 631.050 17.400 ;
        RECT 743.400 16.050 744.450 19.950 ;
        RECT 748.950 19.800 751.050 21.900 ;
        RECT 757.950 19.950 760.050 22.050 ;
        RECT 607.950 10.500 610.050 12.600 ;
        RECT 613.950 10.950 616.050 13.050 ;
        RECT 628.950 11.700 630.150 15.300 ;
        RECT 742.950 13.950 745.050 16.050 ;
        RECT 547.950 7.950 550.050 10.050 ;
        RECT 628.950 9.600 631.050 11.700 ;
        RECT 761.400 10.050 762.450 25.800 ;
        RECT 770.400 25.350 771.600 26.100 ;
        RECT 776.400 25.350 777.600 27.600 ;
        RECT 778.950 25.950 781.050 28.050 ;
        RECT 787.950 26.100 790.050 28.200 ;
        RECT 799.950 26.250 802.050 28.350 ;
        RECT 808.950 26.250 811.050 28.350 ;
        RECT 815.400 27.600 816.450 31.950 ;
        RECT 818.400 28.050 819.450 37.950 ;
        RECT 788.400 25.350 789.600 26.100 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 784.950 22.950 787.050 25.050 ;
        RECT 787.950 22.950 790.050 25.050 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 767.400 20.400 768.600 22.650 ;
        RECT 773.400 21.900 774.600 22.650 ;
        RECT 767.400 16.050 768.450 20.400 ;
        RECT 772.950 19.800 775.050 21.900 ;
        RECT 785.400 20.400 786.600 22.650 ;
        RECT 794.400 20.400 795.600 22.650 ;
        RECT 766.950 13.950 769.050 16.050 ;
        RECT 785.400 10.050 786.450 20.400 ;
        RECT 794.400 16.050 795.450 20.400 ;
        RECT 800.400 19.050 801.450 26.250 ;
        RECT 809.400 25.500 810.600 26.250 ;
        RECT 815.400 25.500 816.600 27.600 ;
        RECT 817.950 25.950 820.050 28.050 ;
        RECT 805.950 23.100 808.050 25.200 ;
        RECT 808.950 23.100 811.050 25.200 ;
        RECT 811.950 23.100 814.050 25.200 ;
        RECT 814.950 23.100 817.050 25.200 ;
        RECT 806.400 20.400 807.600 22.800 ;
        RECT 812.400 22.050 813.600 22.800 ;
        RECT 821.400 22.050 822.450 53.400 ;
        RECT 829.950 52.800 832.050 54.900 ;
        RECT 845.400 53.400 846.600 55.650 ;
        RECT 851.400 53.400 852.600 55.650 ;
        RECT 845.400 43.050 846.450 53.400 ;
        RECT 851.400 49.050 852.450 53.400 ;
        RECT 850.950 46.950 853.050 49.050 ;
        RECT 844.950 40.950 847.050 43.050 ;
        RECT 826.950 33.450 829.050 34.050 ;
        RECT 826.950 32.400 834.450 33.450 ;
        RECT 826.950 31.950 829.050 32.400 ;
        RECT 829.950 27.000 832.050 31.050 ;
        RECT 833.400 30.450 834.450 32.400 ;
        RECT 833.400 29.400 837.450 30.450 ;
        RECT 836.400 27.600 837.450 29.400 ;
        RECT 830.400 25.500 831.600 27.000 ;
        RECT 836.400 25.500 837.600 27.600 ;
        RECT 826.950 23.100 829.050 25.200 ;
        RECT 829.950 23.100 832.050 25.200 ;
        RECT 832.950 23.100 835.050 25.200 ;
        RECT 835.950 23.100 838.050 25.200 ;
        RECT 838.950 23.100 841.050 25.200 ;
        RECT 827.400 22.050 828.600 22.800 ;
        RECT 812.400 20.400 817.050 22.050 ;
        RECT 799.950 16.950 802.050 19.050 ;
        RECT 793.950 13.950 796.050 16.050 ;
        RECT 806.400 10.050 807.450 20.400 ;
        RECT 813.000 19.950 817.050 20.400 ;
        RECT 820.950 19.950 823.050 22.050 ;
        RECT 823.950 16.950 826.050 22.050 ;
        RECT 826.950 19.950 829.050 22.050 ;
        RECT 833.400 21.000 834.600 22.800 ;
        RECT 832.950 16.950 835.050 21.000 ;
        RECT 839.400 20.400 840.600 22.800 ;
        RECT 839.400 16.050 840.450 20.400 ;
        RECT 808.950 15.450 811.050 16.050 ;
        RECT 814.950 15.450 817.050 16.050 ;
        RECT 808.950 14.400 817.050 15.450 ;
        RECT 808.950 13.950 811.050 14.400 ;
        RECT 814.950 13.950 817.050 14.400 ;
        RECT 838.950 13.950 841.050 16.050 ;
        RECT 760.950 7.950 763.050 10.050 ;
        RECT 784.950 7.950 787.050 10.050 ;
        RECT 805.950 7.950 808.050 10.050 ;
        RECT 430.950 4.950 433.050 7.050 ;
        RECT 457.950 4.950 460.050 7.050 ;
      LAYER metal3 ;
        RECT 46.950 822.600 49.050 823.050 ;
        RECT 88.950 822.600 91.050 823.050 ;
        RECT 46.950 821.400 91.050 822.600 ;
        RECT 46.950 820.950 49.050 821.400 ;
        RECT 88.950 820.950 91.050 821.400 ;
        RECT 439.950 822.600 442.050 823.050 ;
        RECT 460.800 822.600 462.900 823.050 ;
        RECT 439.950 821.400 462.900 822.600 ;
        RECT 439.950 820.950 442.050 821.400 ;
        RECT 460.800 820.950 462.900 821.400 ;
        RECT 514.950 822.600 517.050 823.050 ;
        RECT 565.800 822.600 567.900 823.050 ;
        RECT 514.950 821.400 567.900 822.600 ;
        RECT 514.950 820.950 517.050 821.400 ;
        RECT 565.800 820.950 567.900 821.400 ;
        RECT 604.950 822.600 607.050 823.050 ;
        RECT 619.950 822.600 622.050 823.050 ;
        RECT 604.950 821.400 622.050 822.600 ;
        RECT 604.950 820.950 607.050 821.400 ;
        RECT 619.950 820.950 622.050 821.400 ;
        RECT 49.950 819.600 52.050 820.050 ;
        RECT 91.950 819.600 94.050 820.050 ;
        RECT 49.950 818.400 94.050 819.600 ;
        RECT 49.950 817.950 52.050 818.400 ;
        RECT 91.950 817.950 94.050 818.400 ;
        RECT 112.950 819.600 115.050 820.050 ;
        RECT 133.950 819.600 136.050 820.050 ;
        RECT 112.950 818.400 136.050 819.600 ;
        RECT 112.950 817.950 115.050 818.400 ;
        RECT 133.950 817.950 136.050 818.400 ;
        RECT 598.950 819.600 601.050 820.050 ;
        RECT 628.950 819.600 631.050 820.050 ;
        RECT 688.950 819.600 691.050 820.050 ;
        RECT 598.950 818.400 691.050 819.600 ;
        RECT 598.950 817.950 601.050 818.400 ;
        RECT 628.950 817.950 631.050 818.400 ;
        RECT 688.950 817.950 691.050 818.400 ;
        RECT 262.950 816.600 265.050 817.050 ;
        RECT 301.950 816.600 304.050 817.050 ;
        RECT 262.950 815.400 304.050 816.600 ;
        RECT 262.950 814.950 265.050 815.400 ;
        RECT 301.950 814.950 304.050 815.400 ;
        RECT 394.950 816.600 397.050 817.050 ;
        RECT 439.800 816.600 441.900 817.050 ;
        RECT 394.950 815.400 441.900 816.600 ;
        RECT 394.950 814.950 397.050 815.400 ;
        RECT 439.800 814.950 441.900 815.400 ;
        RECT 493.950 816.600 496.050 817.050 ;
        RECT 514.950 816.600 517.050 817.050 ;
        RECT 799.950 816.600 802.050 817.050 ;
        RECT 493.950 815.400 517.050 816.600 ;
        RECT 493.950 814.950 496.050 815.400 ;
        RECT 514.950 814.950 517.050 815.400 ;
        RECT 659.400 815.400 802.050 816.600 ;
        RECT 31.950 813.600 34.050 814.050 ;
        RECT 49.950 813.600 52.050 814.050 ;
        RECT 31.950 812.400 52.050 813.600 ;
        RECT 31.950 811.950 34.050 812.400 ;
        RECT 49.950 811.950 52.050 812.400 ;
        RECT 58.950 813.600 61.050 814.050 ;
        RECT 85.950 813.600 88.050 814.050 ;
        RECT 58.950 812.400 88.050 813.600 ;
        RECT 58.950 811.950 61.050 812.400 ;
        RECT 85.950 811.950 88.050 812.400 ;
        RECT 172.950 813.600 175.050 814.050 ;
        RECT 184.950 813.600 187.050 814.050 ;
        RECT 172.950 812.400 187.050 813.600 ;
        RECT 172.950 811.950 175.050 812.400 ;
        RECT 184.950 811.950 187.050 812.400 ;
        RECT 277.950 813.600 280.050 814.050 ;
        RECT 403.950 813.600 406.050 814.050 ;
        RECT 277.950 812.400 406.050 813.600 ;
        RECT 277.950 811.950 280.050 812.400 ;
        RECT 403.950 811.950 406.050 812.400 ;
        RECT 451.950 813.600 454.050 814.050 ;
        RECT 490.950 813.600 493.050 813.900 ;
        RECT 451.950 812.400 493.050 813.600 ;
        RECT 451.950 811.950 454.050 812.400 ;
        RECT 490.950 811.800 493.050 812.400 ;
        RECT 532.950 813.600 535.050 814.050 ;
        RECT 544.950 813.600 547.050 814.050 ;
        RECT 532.950 812.400 547.050 813.600 ;
        RECT 532.950 811.950 535.050 812.400 ;
        RECT 544.950 811.950 547.050 812.400 ;
        RECT 610.950 813.600 613.050 814.050 ;
        RECT 659.400 813.600 660.600 815.400 ;
        RECT 799.950 814.950 802.050 815.400 ;
        RECT 610.950 812.400 660.600 813.600 ;
        RECT 661.950 813.600 664.050 814.050 ;
        RECT 682.800 813.600 684.900 814.050 ;
        RECT 661.950 812.400 684.900 813.600 ;
        RECT 610.950 811.950 613.050 812.400 ;
        RECT 661.950 811.950 664.050 812.400 ;
        RECT 682.800 811.950 684.900 812.400 ;
        RECT 97.950 810.600 100.050 811.050 ;
        RECT 121.950 810.600 124.050 811.050 ;
        RECT 97.950 809.400 124.050 810.600 ;
        RECT 97.950 808.950 100.050 809.400 ;
        RECT 121.950 808.950 124.050 809.400 ;
        RECT 469.950 810.600 472.050 811.050 ;
        RECT 493.950 810.600 496.050 811.050 ;
        RECT 469.950 809.400 496.050 810.600 ;
        RECT 469.950 808.950 472.050 809.400 ;
        RECT 493.950 808.950 496.050 809.400 ;
        RECT 574.950 808.950 580.050 811.050 ;
        RECT 619.950 810.600 622.050 811.050 ;
        RECT 634.950 810.600 637.050 811.050 ;
        RECT 619.950 809.400 637.050 810.600 ;
        RECT 619.950 808.950 622.050 809.400 ;
        RECT 634.950 808.950 637.050 809.400 ;
        RECT 640.950 810.600 643.050 811.050 ;
        RECT 662.400 810.600 663.600 811.950 ;
        RECT 640.950 809.400 663.600 810.600 ;
        RECT 754.950 810.600 757.050 811.050 ;
        RECT 817.950 810.600 820.050 811.050 ;
        RECT 826.950 810.600 829.050 811.050 ;
        RECT 754.950 809.400 829.050 810.600 ;
        RECT 640.950 808.950 643.050 809.400 ;
        RECT 754.950 808.950 757.050 809.400 ;
        RECT 817.950 808.950 820.050 809.400 ;
        RECT 826.950 808.950 829.050 809.400 ;
        RECT 4.950 807.600 7.050 808.050 ;
        RECT 10.950 807.600 13.050 808.350 ;
        RECT 4.950 806.400 13.050 807.600 ;
        RECT 4.950 805.950 7.050 806.400 ;
        RECT 10.950 806.250 13.050 806.400 ;
        RECT 16.950 806.250 19.050 808.350 ;
        RECT 31.950 807.600 34.050 808.350 ;
        RECT 20.400 806.400 34.050 807.600 ;
        RECT 17.400 802.050 18.600 806.250 ;
        RECT 20.400 802.050 21.600 806.400 ;
        RECT 31.950 806.250 34.050 806.400 ;
        RECT 37.950 807.900 40.050 808.350 ;
        RECT 43.950 807.900 46.050 808.350 ;
        RECT 37.950 806.700 46.050 807.900 ;
        RECT 37.950 806.250 40.050 806.700 ;
        RECT 43.950 806.250 46.050 806.700 ;
        RECT 73.950 807.600 76.050 808.350 ;
        RECT 82.950 807.600 85.050 808.050 ;
        RECT 73.950 806.400 85.050 807.600 ;
        RECT 73.950 806.250 76.050 806.400 ;
        RECT 82.950 805.950 85.050 806.400 ;
        RECT 88.950 807.600 91.050 808.050 ;
        RECT 112.950 807.600 115.050 808.350 ;
        RECT 88.950 806.400 115.050 807.600 ;
        RECT 88.950 805.950 91.050 806.400 ;
        RECT 112.950 806.250 115.050 806.400 ;
        RECT 127.950 806.100 130.050 808.200 ;
        RECT 184.950 807.900 187.050 808.350 ;
        RECT 193.950 807.900 196.050 808.350 ;
        RECT 184.950 806.700 196.050 807.900 ;
        RECT 184.950 806.250 187.050 806.700 ;
        RECT 193.950 806.250 196.050 806.700 ;
        RECT 199.950 806.250 202.050 808.350 ;
        RECT 238.950 807.900 241.050 808.350 ;
        RECT 247.800 807.900 249.900 808.350 ;
        RECT 238.950 806.700 249.900 807.900 ;
        RECT 238.950 806.250 241.050 806.700 ;
        RECT 247.800 806.250 249.900 806.700 ;
        RECT 250.950 807.600 253.050 808.050 ;
        RECT 256.950 807.600 259.050 808.350 ;
        RECT 250.950 806.400 259.050 807.600 ;
        RECT 128.400 804.600 129.600 806.100 ;
        RECT 98.400 803.400 129.600 804.600 ;
        RECT 16.800 799.950 18.900 802.050 ;
        RECT 19.950 799.950 22.050 802.050 ;
        RECT 34.950 801.600 37.050 802.050 ;
        RECT 40.950 801.600 43.050 802.050 ;
        RECT 34.950 800.400 43.050 801.600 ;
        RECT 34.950 799.950 37.050 800.400 ;
        RECT 40.950 799.950 43.050 800.400 ;
        RECT 46.950 801.600 49.050 802.050 ;
        RECT 55.950 801.600 58.050 802.050 ;
        RECT 46.950 800.400 58.050 801.600 ;
        RECT 46.950 799.950 49.050 800.400 ;
        RECT 55.950 799.950 58.050 800.400 ;
        RECT 61.950 801.600 64.050 802.050 ;
        RECT 70.950 801.600 73.050 802.050 ;
        RECT 61.950 800.400 73.050 801.600 ;
        RECT 61.950 799.950 64.050 800.400 ;
        RECT 70.950 799.950 73.050 800.400 ;
        RECT 82.950 801.600 85.050 802.050 ;
        RECT 94.950 801.600 97.050 802.050 ;
        RECT 98.400 801.600 99.600 803.400 ;
        RECT 200.400 802.050 201.600 806.250 ;
        RECT 250.950 805.950 253.050 806.400 ;
        RECT 256.950 806.250 259.050 806.400 ;
        RECT 277.950 806.250 280.050 808.350 ;
        RECT 295.950 807.600 298.050 808.350 ;
        RECT 290.400 806.400 298.050 807.600 ;
        RECT 151.950 801.600 154.050 801.900 ;
        RECT 82.950 800.400 99.600 801.600 ;
        RECT 113.400 800.400 154.050 801.600 ;
        RECT 82.950 799.950 85.050 800.400 ;
        RECT 94.950 799.950 97.050 800.400 ;
        RECT 113.400 799.050 114.600 800.400 ;
        RECT 151.950 799.800 154.050 800.400 ;
        RECT 199.950 799.950 202.050 802.050 ;
        RECT 241.950 801.600 244.050 802.050 ;
        RECT 259.950 801.600 262.050 802.050 ;
        RECT 278.400 801.600 279.600 806.250 ;
        RECT 286.950 804.600 289.050 805.050 ;
        RECT 290.400 804.600 291.600 806.400 ;
        RECT 295.950 806.250 298.050 806.400 ;
        RECT 301.950 807.600 304.050 808.350 ;
        RECT 313.950 807.600 316.050 808.050 ;
        RECT 301.950 806.400 316.050 807.600 ;
        RECT 301.950 806.250 304.050 806.400 ;
        RECT 313.950 805.950 316.050 806.400 ;
        RECT 322.950 807.600 325.050 808.200 ;
        RECT 334.950 807.900 337.050 808.350 ;
        RECT 343.950 807.900 346.050 808.350 ;
        RECT 334.950 807.600 346.050 807.900 ;
        RECT 322.950 806.700 346.050 807.600 ;
        RECT 322.950 806.400 337.050 806.700 ;
        RECT 322.950 806.100 325.050 806.400 ;
        RECT 334.950 806.250 337.050 806.400 ;
        RECT 343.950 806.250 346.050 806.700 ;
        RECT 364.950 807.900 367.050 808.350 ;
        RECT 373.950 807.900 376.050 808.350 ;
        RECT 364.950 806.700 376.050 807.900 ;
        RECT 364.950 806.250 367.050 806.700 ;
        RECT 373.950 806.250 376.050 806.700 ;
        RECT 388.950 806.100 391.050 808.200 ;
        RECT 412.950 806.250 415.050 808.350 ;
        RECT 451.950 807.600 454.050 808.200 ;
        RECT 449.400 806.400 454.050 807.600 ;
        RECT 281.400 804.000 291.600 804.600 ;
        RECT 241.950 800.400 279.600 801.600 ;
        RECT 280.950 803.400 291.600 804.000 ;
        RECT 241.950 799.950 244.050 800.400 ;
        RECT 259.950 799.950 262.050 800.400 ;
        RECT 280.950 799.950 283.050 803.400 ;
        RECT 286.950 802.950 289.050 803.400 ;
        RECT 389.400 802.050 390.600 806.100 ;
        RECT 413.400 802.050 414.600 806.250 ;
        RECT 449.400 802.050 450.600 806.400 ;
        RECT 451.950 806.100 454.050 806.400 ;
        RECT 469.950 807.600 472.050 808.350 ;
        RECT 478.950 807.600 481.050 808.050 ;
        RECT 484.950 807.600 487.050 808.050 ;
        RECT 469.950 806.400 477.600 807.600 ;
        RECT 469.950 806.250 472.050 806.400 ;
        RECT 476.400 802.050 477.600 806.400 ;
        RECT 478.950 806.400 487.050 807.600 ;
        RECT 478.950 805.950 481.050 806.400 ;
        RECT 484.950 805.950 487.050 806.400 ;
        RECT 496.950 806.250 499.050 808.350 ;
        RECT 511.950 806.250 514.050 808.350 ;
        RECT 517.950 807.600 520.050 808.350 ;
        RECT 523.950 807.600 526.050 808.050 ;
        RECT 517.950 806.400 526.050 807.600 ;
        RECT 517.950 806.250 520.050 806.400 ;
        RECT 313.950 801.450 316.050 801.900 ;
        RECT 319.950 801.450 322.050 801.900 ;
        RECT 313.950 800.250 322.050 801.450 ;
        RECT 313.950 799.800 316.050 800.250 ;
        RECT 319.950 799.800 322.050 800.250 ;
        RECT 352.950 801.600 355.050 801.900 ;
        RECT 364.950 801.600 367.050 802.050 ;
        RECT 352.950 800.400 367.050 801.600 ;
        RECT 352.950 799.800 355.050 800.400 ;
        RECT 364.950 799.950 367.050 800.400 ;
        RECT 385.950 800.400 390.600 802.050 ;
        RECT 397.950 801.450 400.050 801.900 ;
        RECT 403.950 801.450 406.050 801.900 ;
        RECT 385.950 799.950 390.000 800.400 ;
        RECT 397.950 800.250 406.050 801.450 ;
        RECT 397.950 799.800 400.050 800.250 ;
        RECT 403.950 799.800 406.050 800.250 ;
        RECT 412.950 799.950 415.050 802.050 ;
        RECT 418.950 801.600 421.050 802.050 ;
        RECT 430.950 801.600 433.050 802.050 ;
        RECT 436.950 801.600 439.050 801.900 ;
        RECT 418.950 800.400 439.050 801.600 ;
        RECT 418.950 799.950 421.050 800.400 ;
        RECT 430.950 799.950 433.050 800.400 ;
        RECT 436.950 799.800 439.050 800.400 ;
        RECT 448.950 799.950 451.050 802.050 ;
        RECT 475.950 799.950 478.050 802.050 ;
        RECT 497.400 801.600 498.600 806.250 ;
        RECT 512.400 804.600 513.600 806.250 ;
        RECT 523.950 805.950 526.050 806.400 ;
        RECT 547.950 807.600 550.050 808.050 ;
        RECT 556.950 807.600 559.050 808.200 ;
        RECT 547.950 806.400 559.050 807.600 ;
        RECT 547.950 805.950 550.050 806.400 ;
        RECT 556.950 806.100 559.050 806.400 ;
        RECT 562.950 807.600 565.050 808.200 ;
        RECT 583.950 807.750 586.050 808.200 ;
        RECT 604.950 807.750 607.050 808.200 ;
        RECT 583.950 807.600 607.050 807.750 ;
        RECT 562.950 806.550 607.050 807.600 ;
        RECT 562.950 806.400 586.050 806.550 ;
        RECT 562.950 806.100 565.050 806.400 ;
        RECT 583.950 806.100 586.050 806.400 ;
        RECT 604.950 806.100 607.050 806.550 ;
        RECT 610.950 805.950 613.050 808.050 ;
        RECT 616.950 806.100 619.050 808.200 ;
        RECT 622.800 806.100 624.900 808.200 ;
        RECT 649.950 807.600 652.050 808.050 ;
        RECT 655.950 807.600 658.050 808.350 ;
        RECT 649.950 806.400 658.050 807.600 ;
        RECT 512.400 803.400 558.600 804.600 ;
        RECT 512.400 802.050 513.600 803.400 ;
        RECT 505.950 801.600 508.050 802.050 ;
        RECT 497.400 800.400 508.050 801.600 ;
        RECT 505.950 799.950 508.050 800.400 ;
        RECT 511.950 799.950 514.050 802.050 ;
        RECT 517.950 801.600 520.050 802.050 ;
        RECT 523.950 801.600 526.050 802.050 ;
        RECT 517.950 800.400 526.050 801.600 ;
        RECT 557.400 801.600 558.600 803.400 ;
        RECT 565.950 801.600 568.050 802.050 ;
        RECT 557.400 800.400 568.050 801.600 ;
        RECT 517.950 799.950 520.050 800.400 ;
        RECT 523.950 799.950 526.050 800.400 ;
        RECT 565.950 799.950 568.050 800.400 ;
        RECT 13.950 798.600 16.050 799.050 ;
        RECT 28.950 798.600 31.050 799.050 ;
        RECT 13.950 797.400 31.050 798.600 ;
        RECT 13.950 796.950 16.050 797.400 ;
        RECT 28.950 796.950 31.050 797.400 ;
        RECT 85.950 798.600 88.050 799.050 ;
        RECT 112.950 798.600 115.050 799.050 ;
        RECT 85.950 797.400 115.050 798.600 ;
        RECT 85.950 796.950 88.050 797.400 ;
        RECT 112.950 796.950 115.050 797.400 ;
        RECT 118.950 798.600 121.050 799.050 ;
        RECT 166.950 798.600 169.050 799.050 ;
        RECT 118.950 797.400 169.050 798.600 ;
        RECT 118.950 796.950 121.050 797.400 ;
        RECT 166.950 796.950 169.050 797.400 ;
        RECT 184.950 798.600 187.050 799.050 ;
        RECT 214.950 798.600 217.050 799.050 ;
        RECT 280.950 798.600 283.050 798.900 ;
        RECT 184.950 797.400 283.050 798.600 ;
        RECT 184.950 796.950 187.050 797.400 ;
        RECT 214.950 796.950 217.050 797.400 ;
        RECT 76.950 795.600 79.050 796.050 ;
        RECT 86.400 795.600 87.600 796.950 ;
        RECT 76.950 794.400 87.600 795.600 ;
        RECT 115.950 795.600 118.050 796.050 ;
        RECT 121.950 795.600 124.050 796.050 ;
        RECT 185.400 795.600 186.600 796.950 ;
        RECT 280.950 796.800 283.050 797.400 ;
        RECT 298.950 798.600 301.050 799.050 ;
        RECT 349.950 798.600 352.050 799.050 ;
        RECT 298.950 797.400 352.050 798.600 ;
        RECT 298.950 796.950 301.050 797.400 ;
        RECT 349.950 796.950 352.050 797.400 ;
        RECT 484.950 798.600 487.050 799.050 ;
        RECT 499.950 798.600 502.050 799.050 ;
        RECT 535.950 798.600 538.050 799.050 ;
        RECT 553.950 798.600 556.050 799.050 ;
        RECT 484.950 797.400 498.600 798.600 ;
        RECT 484.950 796.950 487.050 797.400 ;
        RECT 115.950 794.400 186.600 795.600 ;
        RECT 286.950 795.600 289.050 796.050 ;
        RECT 370.950 795.600 373.050 796.050 ;
        RECT 433.950 795.600 436.050 796.050 ;
        RECT 286.950 794.400 436.050 795.600 ;
        RECT 76.950 793.950 79.050 794.400 ;
        RECT 115.950 793.950 118.050 794.400 ;
        RECT 121.950 793.950 124.050 794.400 ;
        RECT 286.950 793.950 289.050 794.400 ;
        RECT 370.950 793.950 373.050 794.400 ;
        RECT 433.950 793.950 436.050 794.400 ;
        RECT 439.950 795.600 442.050 796.050 ;
        RECT 481.950 795.600 484.050 796.050 ;
        RECT 439.950 794.400 484.050 795.600 ;
        RECT 497.400 795.600 498.600 797.400 ;
        RECT 499.950 797.400 556.050 798.600 ;
        RECT 499.950 796.950 502.050 797.400 ;
        RECT 535.950 796.950 538.050 797.400 ;
        RECT 553.950 796.950 556.050 797.400 ;
        RECT 601.950 798.600 604.050 799.050 ;
        RECT 611.400 798.600 612.600 805.950 ;
        RECT 617.400 804.600 618.600 806.100 ;
        RECT 601.950 797.400 612.600 798.600 ;
        RECT 614.400 803.400 618.600 804.600 ;
        RECT 601.950 796.950 604.050 797.400 ;
        RECT 508.950 795.600 511.050 796.050 ;
        RECT 544.950 795.600 547.050 796.050 ;
        RECT 497.400 794.400 504.600 795.600 ;
        RECT 439.950 793.950 442.050 794.400 ;
        RECT 481.950 793.950 484.050 794.400 ;
        RECT 247.950 792.600 250.050 793.050 ;
        RECT 265.950 792.600 268.050 793.050 ;
        RECT 304.950 792.600 307.050 793.050 ;
        RECT 247.950 791.400 307.050 792.600 ;
        RECT 247.950 790.950 250.050 791.400 ;
        RECT 265.950 790.950 268.050 791.400 ;
        RECT 304.950 790.950 307.050 791.400 ;
        RECT 349.950 792.600 352.050 793.050 ;
        RECT 367.950 792.600 370.050 793.050 ;
        RECT 349.950 791.400 370.050 792.600 ;
        RECT 349.950 790.950 352.050 791.400 ;
        RECT 367.950 790.950 370.050 791.400 ;
        RECT 400.950 792.600 403.050 793.050 ;
        RECT 409.950 792.600 412.050 793.050 ;
        RECT 400.950 791.400 412.050 792.600 ;
        RECT 400.950 790.950 403.050 791.400 ;
        RECT 409.950 790.950 412.050 791.400 ;
        RECT 436.950 792.600 439.050 793.050 ;
        RECT 484.950 792.600 487.050 793.050 ;
        RECT 436.950 791.400 487.050 792.600 ;
        RECT 503.400 792.600 504.600 794.400 ;
        RECT 508.950 794.400 547.050 795.600 ;
        RECT 508.950 793.950 511.050 794.400 ;
        RECT 544.950 793.950 547.050 794.400 ;
        RECT 592.950 795.600 595.050 796.050 ;
        RECT 614.400 795.600 615.600 803.400 ;
        RECT 623.400 802.050 624.600 806.100 ;
        RECT 649.950 805.950 652.050 806.400 ;
        RECT 655.950 806.250 658.050 806.400 ;
        RECT 673.950 806.100 676.050 808.200 ;
        RECT 682.950 807.900 685.050 808.350 ;
        RECT 706.950 807.900 709.050 808.350 ;
        RECT 682.950 806.700 709.050 807.900 ;
        RECT 682.950 806.250 685.050 806.700 ;
        RECT 706.950 806.250 709.050 806.700 ;
        RECT 712.950 807.600 715.050 808.350 ;
        RECT 718.950 807.600 721.050 808.050 ;
        RECT 712.950 806.400 721.050 807.600 ;
        RECT 712.950 806.250 715.050 806.400 ;
        RECT 674.400 802.050 675.600 806.100 ;
        RECT 718.950 805.950 721.050 806.400 ;
        RECT 724.950 806.100 727.050 808.200 ;
        RECT 730.950 807.600 733.050 808.200 ;
        RECT 739.950 807.900 742.050 808.350 ;
        RECT 748.950 807.900 751.050 808.350 ;
        RECT 730.950 806.400 738.600 807.600 ;
        RECT 730.950 806.100 733.050 806.400 ;
        RECT 623.400 800.400 628.050 802.050 ;
        RECT 624.000 799.950 628.050 800.400 ;
        RECT 643.950 801.600 646.050 802.050 ;
        RECT 655.950 801.600 658.050 802.050 ;
        RECT 643.950 800.400 658.050 801.600 ;
        RECT 643.950 799.950 646.050 800.400 ;
        RECT 655.950 799.950 658.050 800.400 ;
        RECT 670.950 800.400 675.600 802.050 ;
        RECT 691.950 801.600 694.050 801.900 ;
        RECT 703.950 801.600 706.050 802.050 ;
        RECT 691.950 800.400 706.050 801.600 ;
        RECT 670.950 799.950 675.000 800.400 ;
        RECT 691.950 799.800 694.050 800.400 ;
        RECT 703.950 799.950 706.050 800.400 ;
        RECT 709.950 801.600 712.050 802.050 ;
        RECT 725.400 801.600 726.600 806.100 ;
        RECT 737.400 804.600 738.600 806.400 ;
        RECT 739.950 806.700 751.050 807.900 ;
        RECT 739.950 806.250 742.050 806.700 ;
        RECT 748.950 806.250 751.050 806.700 ;
        RECT 769.950 807.600 772.050 808.350 ;
        RECT 787.950 807.600 790.050 808.350 ;
        RECT 769.950 806.400 790.050 807.600 ;
        RECT 769.950 806.250 772.050 806.400 ;
        RECT 787.950 806.250 790.050 806.400 ;
        RECT 793.950 807.600 796.050 808.350 ;
        RECT 802.950 807.600 805.050 808.050 ;
        RECT 811.950 807.600 814.050 808.200 ;
        RECT 793.950 806.400 801.600 807.600 ;
        RECT 793.950 806.250 796.050 806.400 ;
        RECT 800.400 804.600 801.600 806.400 ;
        RECT 802.950 806.400 814.050 807.600 ;
        RECT 802.950 805.950 805.050 806.400 ;
        RECT 811.950 806.100 814.050 806.400 ;
        RECT 832.950 807.600 835.050 808.200 ;
        RECT 841.950 807.600 844.050 808.050 ;
        RECT 832.950 806.400 844.050 807.600 ;
        RECT 832.950 806.100 835.050 806.400 ;
        RECT 841.950 805.950 844.050 806.400 ;
        RECT 737.400 803.400 747.600 804.600 ;
        RECT 800.400 803.400 816.600 804.600 ;
        RECT 709.950 800.400 726.600 801.600 ;
        RECT 746.400 801.600 747.600 803.400 ;
        RECT 815.400 801.900 816.600 803.400 ;
        RECT 746.400 800.400 750.600 801.600 ;
        RECT 709.950 799.950 712.050 800.400 ;
        RECT 637.950 798.600 640.050 799.050 ;
        RECT 664.950 798.600 667.050 799.050 ;
        RECT 637.950 797.400 667.050 798.600 ;
        RECT 637.950 796.950 640.050 797.400 ;
        RECT 664.950 796.950 667.050 797.400 ;
        RECT 676.950 798.600 679.050 799.050 ;
        RECT 691.950 798.600 694.050 799.050 ;
        RECT 676.950 797.400 694.050 798.600 ;
        RECT 749.400 798.600 750.600 800.400 ;
        RECT 799.950 801.450 802.050 801.900 ;
        RECT 808.950 801.450 811.050 801.900 ;
        RECT 799.950 800.250 811.050 801.450 ;
        RECT 799.950 799.800 802.050 800.250 ;
        RECT 808.950 799.800 811.050 800.250 ;
        RECT 814.950 801.600 817.050 801.900 ;
        RECT 829.950 801.600 832.050 801.900 ;
        RECT 814.950 800.400 832.050 801.600 ;
        RECT 814.950 799.800 817.050 800.400 ;
        RECT 829.950 799.800 832.050 800.400 ;
        RECT 784.950 798.600 787.050 799.050 ;
        RECT 749.400 797.400 787.050 798.600 ;
        RECT 676.950 796.950 679.050 797.400 ;
        RECT 691.950 796.950 694.050 797.400 ;
        RECT 784.950 796.950 787.050 797.400 ;
        RECT 592.950 794.400 615.600 795.600 ;
        RECT 619.950 795.600 622.050 796.050 ;
        RECT 709.950 795.600 712.050 796.050 ;
        RECT 619.950 794.400 712.050 795.600 ;
        RECT 592.950 793.950 595.050 794.400 ;
        RECT 619.950 793.950 622.050 794.400 ;
        RECT 709.950 793.950 712.050 794.400 ;
        RECT 562.950 792.600 565.050 793.050 ;
        RECT 503.400 791.400 565.050 792.600 ;
        RECT 436.950 790.950 439.050 791.400 ;
        RECT 484.950 790.950 487.050 791.400 ;
        RECT 562.950 790.950 565.050 791.400 ;
        RECT 574.950 792.600 577.050 793.050 ;
        RECT 604.950 792.600 607.050 793.050 ;
        RECT 574.950 791.400 607.050 792.600 ;
        RECT 574.950 790.950 577.050 791.400 ;
        RECT 604.950 790.950 607.050 791.400 ;
        RECT 613.950 792.600 616.050 793.050 ;
        RECT 628.950 792.600 631.050 793.050 ;
        RECT 613.950 791.400 631.050 792.600 ;
        RECT 613.950 790.950 616.050 791.400 ;
        RECT 628.950 790.950 631.050 791.400 ;
        RECT 634.950 792.600 637.050 793.050 ;
        RECT 730.950 792.600 733.050 793.050 ;
        RECT 733.950 792.600 736.050 793.050 ;
        RECT 634.950 791.400 736.050 792.600 ;
        RECT 634.950 790.950 637.050 791.400 ;
        RECT 730.950 790.950 733.050 791.400 ;
        RECT 733.950 790.950 736.050 791.400 ;
        RECT 61.950 789.600 64.050 790.050 ;
        RECT 82.950 789.600 85.050 790.050 ;
        RECT 61.950 788.400 85.050 789.600 ;
        RECT 61.950 787.950 64.050 788.400 ;
        RECT 82.950 787.950 85.050 788.400 ;
        RECT 109.950 789.600 112.050 790.050 ;
        RECT 118.950 789.600 121.050 790.050 ;
        RECT 109.950 788.400 121.050 789.600 ;
        RECT 109.950 787.950 112.050 788.400 ;
        RECT 118.950 787.950 121.050 788.400 ;
        RECT 166.950 789.600 169.050 790.050 ;
        RECT 190.950 789.600 193.050 790.050 ;
        RECT 166.950 788.400 193.050 789.600 ;
        RECT 166.950 787.950 169.050 788.400 ;
        RECT 190.950 787.950 193.050 788.400 ;
        RECT 199.950 789.600 202.050 790.050 ;
        RECT 373.950 789.600 376.050 790.050 ;
        RECT 409.950 789.600 412.050 789.900 ;
        RECT 199.950 788.400 354.600 789.600 ;
        RECT 199.950 787.950 202.050 788.400 ;
        RECT 353.400 787.050 354.600 788.400 ;
        RECT 373.950 788.400 412.050 789.600 ;
        RECT 373.950 787.950 376.050 788.400 ;
        RECT 409.950 787.800 412.050 788.400 ;
        RECT 421.950 789.600 424.050 790.050 ;
        RECT 439.950 789.600 442.050 790.050 ;
        RECT 421.950 788.400 442.050 789.600 ;
        RECT 421.950 787.950 424.050 788.400 ;
        RECT 439.950 787.950 442.050 788.400 ;
        RECT 460.950 789.600 463.050 790.050 ;
        RECT 493.800 789.600 495.900 790.050 ;
        RECT 460.950 788.400 495.900 789.600 ;
        RECT 460.950 787.950 463.050 788.400 ;
        RECT 493.800 787.950 495.900 788.400 ;
        RECT 496.950 789.600 499.050 790.050 ;
        RECT 523.950 789.600 526.050 790.050 ;
        RECT 496.950 788.400 526.050 789.600 ;
        RECT 496.950 787.950 499.050 788.400 ;
        RECT 523.950 787.950 526.050 788.400 ;
        RECT 589.950 789.600 592.050 790.050 ;
        RECT 601.950 789.600 604.050 790.050 ;
        RECT 589.950 788.400 604.050 789.600 ;
        RECT 589.950 787.950 592.050 788.400 ;
        RECT 601.950 787.950 604.050 788.400 ;
        RECT 646.950 789.600 649.050 790.050 ;
        RECT 775.950 789.600 778.050 790.050 ;
        RECT 835.950 789.600 838.050 790.050 ;
        RECT 646.950 788.400 838.050 789.600 ;
        RECT 646.950 787.950 649.050 788.400 ;
        RECT 775.950 787.950 778.050 788.400 ;
        RECT 835.950 787.950 838.050 788.400 ;
        RECT 211.950 786.600 214.050 787.050 ;
        RECT 235.950 786.600 238.050 787.050 ;
        RECT 211.950 785.400 238.050 786.600 ;
        RECT 211.950 784.950 214.050 785.400 ;
        RECT 235.950 784.950 238.050 785.400 ;
        RECT 274.950 786.600 277.050 787.050 ;
        RECT 292.950 786.600 295.050 787.050 ;
        RECT 274.950 785.400 295.050 786.600 ;
        RECT 274.950 784.950 277.050 785.400 ;
        RECT 292.950 784.950 295.050 785.400 ;
        RECT 352.950 786.600 355.050 787.050 ;
        RECT 370.950 786.600 373.050 787.050 ;
        RECT 412.950 786.600 415.050 787.050 ;
        RECT 352.950 785.400 415.050 786.600 ;
        RECT 352.950 784.950 355.050 785.400 ;
        RECT 370.950 784.950 373.050 785.400 ;
        RECT 412.950 784.950 415.050 785.400 ;
        RECT 514.950 786.600 517.050 787.050 ;
        RECT 529.950 786.600 532.050 787.050 ;
        RECT 550.950 786.600 553.050 787.050 ;
        RECT 514.950 785.400 553.050 786.600 ;
        RECT 514.950 784.950 517.050 785.400 ;
        RECT 529.950 784.950 532.050 785.400 ;
        RECT 550.950 784.950 553.050 785.400 ;
        RECT 559.950 786.600 562.050 787.050 ;
        RECT 580.950 786.600 583.050 787.050 ;
        RECT 610.950 786.600 613.050 787.050 ;
        RECT 700.950 786.600 703.050 787.050 ;
        RECT 559.950 785.400 703.050 786.600 ;
        RECT 559.950 784.950 562.050 785.400 ;
        RECT 580.950 784.950 583.050 785.400 ;
        RECT 610.950 784.950 613.050 785.400 ;
        RECT 700.950 784.950 703.050 785.400 ;
        RECT 709.950 786.600 712.050 787.050 ;
        RECT 766.950 786.600 769.050 787.050 ;
        RECT 709.950 785.400 769.050 786.600 ;
        RECT 709.950 784.950 712.050 785.400 ;
        RECT 766.950 784.950 769.050 785.400 ;
        RECT 28.950 783.600 31.050 784.050 ;
        RECT 82.950 783.600 85.050 784.050 ;
        RECT 28.950 782.400 85.050 783.600 ;
        RECT 28.950 781.950 31.050 782.400 ;
        RECT 82.950 781.950 85.050 782.400 ;
        RECT 169.950 783.600 172.050 784.050 ;
        RECT 175.950 783.600 178.050 784.050 ;
        RECT 275.400 783.600 276.600 784.950 ;
        RECT 169.950 782.400 276.600 783.600 ;
        RECT 343.950 783.600 346.050 784.050 ;
        RECT 385.950 783.600 388.050 784.050 ;
        RECT 343.950 782.400 388.050 783.600 ;
        RECT 169.950 781.950 172.050 782.400 ;
        RECT 175.950 781.950 178.050 782.400 ;
        RECT 343.950 781.950 346.050 782.400 ;
        RECT 385.950 781.950 388.050 782.400 ;
        RECT 391.950 783.600 394.050 784.050 ;
        RECT 415.950 783.600 418.050 784.050 ;
        RECT 496.950 783.600 499.050 784.050 ;
        RECT 391.950 782.400 418.050 783.600 ;
        RECT 391.950 781.950 394.050 782.400 ;
        RECT 415.950 781.950 418.050 782.400 ;
        RECT 458.400 782.400 499.050 783.600 ;
        RECT 178.950 780.600 181.050 781.050 ;
        RECT 226.950 780.600 229.050 781.050 ;
        RECT 178.950 779.400 229.050 780.600 ;
        RECT 178.950 778.950 181.050 779.400 ;
        RECT 226.950 778.950 229.050 779.400 ;
        RECT 433.950 780.600 436.050 781.050 ;
        RECT 458.400 780.600 459.600 782.400 ;
        RECT 496.950 781.950 499.050 782.400 ;
        RECT 523.950 783.600 526.050 784.050 ;
        RECT 553.950 783.600 556.050 784.050 ;
        RECT 583.950 783.600 586.050 784.050 ;
        RECT 625.950 783.600 628.050 784.050 ;
        RECT 661.950 783.600 664.050 784.050 ;
        RECT 670.950 783.600 673.050 784.050 ;
        RECT 523.950 782.400 582.600 783.600 ;
        RECT 523.950 781.950 526.050 782.400 ;
        RECT 553.950 781.950 556.050 782.400 ;
        RECT 433.950 779.400 459.600 780.600 ;
        RECT 478.950 780.600 481.050 781.050 ;
        RECT 511.950 780.600 514.050 781.050 ;
        RECT 478.950 779.400 514.050 780.600 ;
        RECT 581.400 780.600 582.600 782.400 ;
        RECT 583.950 782.400 673.050 783.600 ;
        RECT 583.950 781.950 586.050 782.400 ;
        RECT 625.950 781.950 628.050 782.400 ;
        RECT 661.950 781.950 664.050 782.400 ;
        RECT 670.950 781.950 673.050 782.400 ;
        RECT 643.950 780.600 646.050 781.050 ;
        RECT 682.950 780.600 685.050 781.050 ;
        RECT 581.400 779.400 685.050 780.600 ;
        RECT 433.950 778.950 436.050 779.400 ;
        RECT 478.950 778.950 481.050 779.400 ;
        RECT 511.950 778.950 514.050 779.400 ;
        RECT 643.950 778.950 646.050 779.400 ;
        RECT 682.950 778.950 685.050 779.400 ;
        RECT 700.950 780.600 703.050 781.050 ;
        RECT 727.950 780.600 730.050 781.050 ;
        RECT 700.950 779.400 730.050 780.600 ;
        RECT 700.950 778.950 703.050 779.400 ;
        RECT 727.950 778.950 730.050 779.400 ;
        RECT 70.950 777.600 73.050 778.050 ;
        RECT 145.950 777.600 148.050 778.050 ;
        RECT 70.950 776.400 148.050 777.600 ;
        RECT 70.950 775.950 73.050 776.400 ;
        RECT 145.950 775.950 148.050 776.400 ;
        RECT 190.950 777.600 193.050 778.050 ;
        RECT 319.950 777.600 322.050 778.050 ;
        RECT 190.950 776.400 322.050 777.600 ;
        RECT 190.950 775.950 193.050 776.400 ;
        RECT 319.950 775.950 322.050 776.400 ;
        RECT 331.950 777.600 334.050 778.050 ;
        RECT 367.950 777.600 370.050 778.050 ;
        RECT 331.950 776.400 370.050 777.600 ;
        RECT 331.950 775.950 334.050 776.400 ;
        RECT 367.950 775.950 370.050 776.400 ;
        RECT 484.950 777.600 487.050 778.050 ;
        RECT 505.950 777.600 508.050 778.050 ;
        RECT 484.950 776.400 508.050 777.600 ;
        RECT 484.950 775.950 487.050 776.400 ;
        RECT 505.950 775.950 508.050 776.400 ;
        RECT 520.950 777.600 523.050 778.050 ;
        RECT 547.800 777.600 549.900 778.050 ;
        RECT 520.950 776.400 549.900 777.600 ;
        RECT 520.950 775.950 523.050 776.400 ;
        RECT 547.800 775.950 549.900 776.400 ;
        RECT 550.950 777.600 553.050 778.050 ;
        RECT 592.950 777.600 595.050 778.050 ;
        RECT 646.950 777.600 649.050 778.050 ;
        RECT 550.950 776.400 595.050 777.600 ;
        RECT 550.950 775.950 553.050 776.400 ;
        RECT 592.950 775.950 595.050 776.400 ;
        RECT 596.400 776.400 649.050 777.600 ;
        RECT 43.950 774.600 46.050 775.050 ;
        RECT 79.950 774.600 82.050 775.050 ;
        RECT 43.950 773.400 82.050 774.600 ;
        RECT 43.950 772.950 46.050 773.400 ;
        RECT 79.950 772.950 82.050 773.400 ;
        RECT 427.950 774.600 430.050 775.050 ;
        RECT 478.950 774.600 481.050 775.050 ;
        RECT 427.950 773.400 481.050 774.600 ;
        RECT 427.950 772.950 430.050 773.400 ;
        RECT 478.950 772.950 481.050 773.400 ;
        RECT 535.950 774.600 538.050 775.050 ;
        RECT 541.950 774.600 544.050 775.050 ;
        RECT 535.950 773.400 544.050 774.600 ;
        RECT 535.950 772.950 538.050 773.400 ;
        RECT 541.950 772.950 544.050 773.400 ;
        RECT 562.950 774.600 565.050 775.050 ;
        RECT 596.400 774.600 597.600 776.400 ;
        RECT 646.950 775.950 649.050 776.400 ;
        RECT 802.950 777.600 805.050 778.050 ;
        RECT 826.950 777.600 829.050 778.050 ;
        RECT 802.950 776.400 829.050 777.600 ;
        RECT 802.950 775.950 805.050 776.400 ;
        RECT 826.950 775.950 829.050 776.400 ;
        RECT 562.950 773.400 597.600 774.600 ;
        RECT 598.950 774.600 601.050 775.050 ;
        RECT 649.950 774.600 652.050 775.050 ;
        RECT 598.950 773.400 652.050 774.600 ;
        RECT 562.950 772.950 565.050 773.400 ;
        RECT 598.950 772.950 601.050 773.400 ;
        RECT 649.950 772.950 652.050 773.400 ;
        RECT 712.950 774.600 715.050 775.050 ;
        RECT 718.950 774.600 721.050 775.050 ;
        RECT 736.950 774.600 739.050 775.050 ;
        RECT 772.950 774.600 775.050 775.050 ;
        RECT 712.950 773.400 775.050 774.600 ;
        RECT 712.950 772.950 715.050 773.400 ;
        RECT 718.950 772.950 721.050 773.400 ;
        RECT 736.950 772.950 739.050 773.400 ;
        RECT 772.950 772.950 775.050 773.400 ;
        RECT 175.950 771.600 178.050 772.050 ;
        RECT 202.950 771.600 205.050 772.050 ;
        RECT 229.950 771.600 232.050 772.050 ;
        RECT 331.950 771.600 334.050 772.050 ;
        RECT 161.400 770.400 334.050 771.600 ;
        RECT 16.950 768.600 19.050 769.050 ;
        RECT 31.950 768.600 34.050 769.050 ;
        RECT 46.950 768.600 49.050 769.050 ;
        RECT 16.950 767.400 49.050 768.600 ;
        RECT 16.950 766.950 19.050 767.400 ;
        RECT 31.950 766.950 34.050 767.400 ;
        RECT 46.950 766.950 49.050 767.400 ;
        RECT 70.950 768.600 73.050 769.050 ;
        RECT 97.950 768.600 100.050 769.050 ;
        RECT 70.950 767.400 100.050 768.600 ;
        RECT 70.950 766.950 73.050 767.400 ;
        RECT 97.950 766.950 100.050 767.400 ;
        RECT 145.950 768.600 148.050 769.050 ;
        RECT 161.400 768.600 162.600 770.400 ;
        RECT 175.950 769.950 178.050 770.400 ;
        RECT 202.950 769.950 205.050 770.400 ;
        RECT 229.950 769.950 232.050 770.400 ;
        RECT 331.950 769.950 334.050 770.400 ;
        RECT 361.950 771.600 364.050 772.050 ;
        RECT 379.950 771.600 382.050 772.050 ;
        RECT 409.950 771.600 412.050 772.050 ;
        RECT 421.950 771.600 424.050 772.050 ;
        RECT 361.950 770.400 424.050 771.600 ;
        RECT 361.950 769.950 364.050 770.400 ;
        RECT 379.950 769.950 382.050 770.400 ;
        RECT 409.950 769.950 412.050 770.400 ;
        RECT 421.950 769.950 424.050 770.400 ;
        RECT 547.950 771.600 550.050 772.050 ;
        RECT 589.950 771.600 592.050 772.050 ;
        RECT 547.950 770.400 592.050 771.600 ;
        RECT 547.950 769.950 550.050 770.400 ;
        RECT 589.950 769.950 592.050 770.400 ;
        RECT 811.950 771.600 814.050 772.050 ;
        RECT 823.950 771.600 826.050 772.050 ;
        RECT 811.950 770.400 826.050 771.600 ;
        RECT 811.950 769.950 814.050 770.400 ;
        RECT 823.950 769.950 826.050 770.400 ;
        RECT 145.950 767.400 162.600 768.600 ;
        RECT 184.950 768.600 187.050 769.050 ;
        RECT 196.950 768.600 199.050 769.050 ;
        RECT 184.950 767.400 199.050 768.600 ;
        RECT 145.950 766.950 148.050 767.400 ;
        RECT 184.950 766.950 187.050 767.400 ;
        RECT 196.950 766.950 199.050 767.400 ;
        RECT 334.950 768.600 337.050 769.050 ;
        RECT 343.950 768.600 346.050 769.050 ;
        RECT 334.950 767.400 346.050 768.600 ;
        RECT 334.950 766.950 337.050 767.400 ;
        RECT 343.950 766.950 346.050 767.400 ;
        RECT 481.950 768.600 484.050 768.900 ;
        RECT 541.950 768.600 544.050 769.050 ;
        RECT 481.950 767.400 544.050 768.600 ;
        RECT 481.950 766.800 484.050 767.400 ;
        RECT 541.950 766.950 544.050 767.400 ;
        RECT 550.950 768.600 553.050 769.050 ;
        RECT 574.800 768.600 576.900 769.050 ;
        RECT 550.950 767.400 576.900 768.600 ;
        RECT 550.950 766.950 553.050 767.400 ;
        RECT 574.800 766.950 576.900 767.400 ;
        RECT 577.950 768.600 580.050 769.050 ;
        RECT 613.950 768.600 616.050 769.050 ;
        RECT 649.950 768.600 652.050 769.050 ;
        RECT 577.950 767.400 591.600 768.600 ;
        RECT 577.950 766.950 580.050 767.400 ;
        RECT 103.950 765.600 106.050 766.050 ;
        RECT 136.800 765.600 138.900 766.050 ;
        RECT 103.950 764.400 138.900 765.600 ;
        RECT 103.950 763.950 106.050 764.400 ;
        RECT 136.800 763.950 138.900 764.400 ;
        RECT 139.950 765.600 142.050 766.050 ;
        RECT 178.950 765.600 181.050 766.050 ;
        RECT 139.950 764.400 181.050 765.600 ;
        RECT 139.950 763.950 142.050 764.400 ;
        RECT 178.950 763.950 181.050 764.400 ;
        RECT 250.950 765.600 253.050 766.050 ;
        RECT 271.950 765.600 274.050 766.050 ;
        RECT 286.950 765.600 289.050 766.050 ;
        RECT 250.950 764.400 289.050 765.600 ;
        RECT 250.950 763.950 253.050 764.400 ;
        RECT 10.950 761.100 13.050 763.200 ;
        RECT 37.950 762.600 40.050 763.200 ;
        RECT 43.950 762.600 46.050 763.050 ;
        RECT 52.950 762.600 55.050 763.200 ;
        RECT 37.950 761.400 55.050 762.600 ;
        RECT 37.950 761.100 40.050 761.400 ;
        RECT 11.400 759.600 12.600 761.100 ;
        RECT 43.950 760.950 46.050 761.400 ;
        RECT 52.950 761.100 55.050 761.400 ;
        RECT 76.950 762.600 79.050 763.050 ;
        RECT 91.950 762.600 94.050 763.050 ;
        RECT 76.950 761.400 94.050 762.600 ;
        RECT 76.950 760.950 79.050 761.400 ;
        RECT 91.950 760.950 94.050 761.400 ;
        RECT 109.950 762.600 112.050 763.200 ;
        RECT 121.950 762.600 124.050 763.050 ;
        RECT 109.950 761.400 124.050 762.600 ;
        RECT 109.950 761.100 112.050 761.400 ;
        RECT 121.950 760.950 124.050 761.400 ;
        RECT 151.950 762.600 154.050 763.050 ;
        RECT 163.950 762.600 166.050 763.050 ;
        RECT 151.950 761.400 166.050 762.600 ;
        RECT 151.950 760.950 154.050 761.400 ;
        RECT 11.400 758.400 15.600 759.600 ;
        RECT 14.400 756.600 15.600 758.400 ;
        RECT 161.400 757.050 162.600 761.400 ;
        RECT 163.950 760.950 166.050 761.400 ;
        RECT 190.950 762.600 193.050 763.200 ;
        RECT 196.950 762.600 199.050 763.050 ;
        RECT 190.950 761.400 199.050 762.600 ;
        RECT 190.950 761.100 193.050 761.400 ;
        RECT 196.950 760.950 199.050 761.400 ;
        RECT 205.950 761.100 208.050 763.200 ;
        RECT 226.950 762.750 229.050 763.200 ;
        RECT 250.950 762.750 253.050 762.900 ;
        RECT 226.950 761.550 253.050 762.750 ;
        RECT 226.950 761.100 229.050 761.550 ;
        RECT 40.950 756.600 43.050 757.050 ;
        RECT 14.400 755.400 43.050 756.600 ;
        RECT 40.950 754.950 43.050 755.400 ;
        RECT 46.950 756.600 49.050 757.050 ;
        RECT 67.950 756.600 70.050 756.750 ;
        RECT 46.950 755.400 70.050 756.600 ;
        RECT 46.950 754.950 49.050 755.400 ;
        RECT 67.950 754.650 70.050 755.400 ;
        RECT 82.950 756.600 85.050 757.050 ;
        RECT 103.950 756.600 106.050 757.050 ;
        RECT 82.950 755.400 106.050 756.600 ;
        RECT 82.950 754.950 85.050 755.400 ;
        RECT 103.950 754.950 106.050 755.400 ;
        RECT 136.950 756.600 139.050 757.050 ;
        RECT 154.950 756.600 157.050 757.050 ;
        RECT 136.950 755.400 157.050 756.600 ;
        RECT 136.950 754.950 139.050 755.400 ;
        RECT 154.950 754.950 157.050 755.400 ;
        RECT 160.950 754.950 163.050 757.050 ;
        RECT 187.950 756.600 190.050 756.900 ;
        RECT 206.400 756.600 207.600 761.100 ;
        RECT 250.950 760.800 253.050 761.550 ;
        RECT 238.950 756.600 241.050 757.050 ;
        RECT 254.400 756.750 255.600 764.400 ;
        RECT 271.950 763.950 274.050 764.400 ;
        RECT 286.950 763.950 289.050 764.400 ;
        RECT 319.950 765.600 322.050 766.050 ;
        RECT 358.950 765.600 361.050 766.050 ;
        RECT 319.950 764.400 361.050 765.600 ;
        RECT 319.950 763.950 322.050 764.400 ;
        RECT 358.950 763.950 361.050 764.400 ;
        RECT 406.950 765.600 409.050 766.050 ;
        RECT 421.950 765.600 424.050 766.050 ;
        RECT 406.950 764.400 424.050 765.600 ;
        RECT 406.950 763.950 409.050 764.400 ;
        RECT 421.950 763.950 424.050 764.400 ;
        RECT 460.950 765.600 463.050 766.050 ;
        RECT 475.950 765.600 478.050 766.050 ;
        RECT 460.950 764.400 478.050 765.600 ;
        RECT 460.950 763.950 463.050 764.400 ;
        RECT 475.950 763.950 478.050 764.400 ;
        RECT 502.950 765.600 505.050 766.050 ;
        RECT 517.950 765.600 520.050 766.050 ;
        RECT 502.950 764.400 520.050 765.600 ;
        RECT 502.950 763.950 505.050 764.400 ;
        RECT 517.950 763.950 520.050 764.400 ;
        RECT 544.950 765.600 547.050 766.050 ;
        RECT 586.950 765.600 589.050 766.050 ;
        RECT 544.950 764.400 589.050 765.600 ;
        RECT 590.400 765.600 591.600 767.400 ;
        RECT 613.950 767.400 652.050 768.600 ;
        RECT 613.950 766.950 616.050 767.400 ;
        RECT 649.950 766.950 652.050 767.400 ;
        RECT 688.950 768.600 691.050 769.050 ;
        RECT 718.950 768.600 721.050 769.050 ;
        RECT 688.950 767.400 721.050 768.600 ;
        RECT 688.950 766.950 691.050 767.400 ;
        RECT 718.950 766.950 721.050 767.400 ;
        RECT 784.950 768.600 787.050 769.050 ;
        RECT 799.950 768.600 802.050 769.050 ;
        RECT 784.950 767.400 802.050 768.600 ;
        RECT 784.950 766.950 787.050 767.400 ;
        RECT 799.950 766.950 802.050 767.400 ;
        RECT 817.950 768.600 820.050 769.050 ;
        RECT 862.950 768.600 865.050 769.050 ;
        RECT 817.950 767.400 865.050 768.600 ;
        RECT 817.950 766.950 820.050 767.400 ;
        RECT 862.950 766.950 865.050 767.400 ;
        RECT 607.950 765.600 610.050 766.050 ;
        RECT 590.400 764.400 610.050 765.600 ;
        RECT 544.950 763.950 547.050 764.400 ;
        RECT 586.950 763.950 589.050 764.400 ;
        RECT 607.950 763.950 610.050 764.400 ;
        RECT 685.950 765.600 688.050 766.050 ;
        RECT 694.950 765.600 697.050 766.050 ;
        RECT 709.950 765.600 712.050 766.050 ;
        RECT 685.950 764.400 712.050 765.600 ;
        RECT 685.950 763.950 688.050 764.400 ;
        RECT 694.950 763.950 697.050 764.400 ;
        RECT 709.950 763.950 712.050 764.400 ;
        RECT 745.950 765.600 748.050 766.050 ;
        RECT 754.950 765.600 757.050 766.050 ;
        RECT 745.950 764.400 757.050 765.600 ;
        RECT 745.950 763.950 748.050 764.400 ;
        RECT 754.950 763.950 757.050 764.400 ;
        RECT 802.950 765.600 805.050 766.050 ;
        RECT 802.950 765.000 822.600 765.600 ;
        RECT 802.950 764.400 823.050 765.000 ;
        RECT 802.950 763.950 805.050 764.400 ;
        RECT 256.950 762.600 259.050 763.050 ;
        RECT 265.950 762.600 268.050 763.050 ;
        RECT 319.950 762.600 322.050 762.900 ;
        RECT 334.950 762.600 337.050 763.050 ;
        RECT 256.950 761.400 270.600 762.600 ;
        RECT 256.950 760.950 259.050 761.400 ;
        RECT 265.950 760.950 268.050 761.400 ;
        RECT 269.400 759.600 270.600 761.400 ;
        RECT 319.950 761.400 337.050 762.600 ;
        RECT 319.950 760.800 322.050 761.400 ;
        RECT 334.950 760.950 337.050 761.400 ;
        RECT 340.950 762.600 343.050 763.050 ;
        RECT 346.950 762.600 349.050 763.050 ;
        RECT 340.950 761.400 349.050 762.600 ;
        RECT 340.950 760.950 343.050 761.400 ;
        RECT 346.950 760.950 349.050 761.400 ;
        RECT 373.950 762.600 376.050 763.050 ;
        RECT 388.950 762.600 391.050 763.050 ;
        RECT 400.950 762.600 403.050 763.050 ;
        RECT 373.950 761.400 387.600 762.600 ;
        RECT 373.950 760.950 376.050 761.400 ;
        RECT 386.400 759.600 387.600 761.400 ;
        RECT 388.950 761.400 403.050 762.600 ;
        RECT 388.950 760.950 391.050 761.400 ;
        RECT 400.950 760.950 403.050 761.400 ;
        RECT 433.950 759.600 436.050 763.050 ;
        RECT 448.950 762.600 451.050 763.050 ;
        RECT 448.950 761.400 459.600 762.600 ;
        RECT 448.950 760.950 451.050 761.400 ;
        RECT 269.400 758.400 288.600 759.600 ;
        RECT 386.400 758.400 399.600 759.600 ;
        RECT 404.400 759.000 436.050 759.600 ;
        RECT 458.400 759.600 459.600 761.400 ;
        RECT 481.950 759.600 484.050 763.050 ;
        RECT 496.950 760.950 499.050 763.050 ;
        RECT 514.950 762.600 517.050 763.050 ;
        RECT 514.950 761.400 522.600 762.600 ;
        RECT 514.950 760.950 517.050 761.400 ;
        RECT 187.950 755.400 241.050 756.600 ;
        RECT 187.950 754.800 190.050 755.400 ;
        RECT 238.950 754.950 241.050 755.400 ;
        RECT 253.950 754.650 256.050 756.750 ;
        RECT 287.400 756.600 288.600 758.400 ;
        RECT 289.950 756.600 292.050 756.750 ;
        RECT 307.950 756.600 310.050 757.050 ;
        RECT 287.400 755.400 310.050 756.600 ;
        RECT 289.950 754.650 292.050 755.400 ;
        RECT 307.950 754.950 310.050 755.400 ;
        RECT 325.950 756.600 328.050 757.050 ;
        RECT 398.400 756.750 399.600 758.400 ;
        RECT 403.950 758.400 435.600 759.000 ;
        RECT 458.400 758.400 468.600 759.600 ;
        RECT 337.950 756.600 340.050 756.750 ;
        RECT 325.950 755.400 340.050 756.600 ;
        RECT 325.950 754.950 328.050 755.400 ;
        RECT 337.950 754.650 340.050 755.400 ;
        RECT 346.950 756.300 349.050 756.750 ;
        RECT 352.950 756.300 355.050 756.750 ;
        RECT 346.950 755.100 355.050 756.300 ;
        RECT 346.950 754.650 349.050 755.100 ;
        RECT 352.950 754.650 355.050 755.100 ;
        RECT 364.950 756.300 367.050 756.750 ;
        RECT 391.950 756.300 394.050 756.750 ;
        RECT 364.950 755.100 394.050 756.300 ;
        RECT 364.950 754.650 367.050 755.100 ;
        RECT 391.950 754.650 394.050 755.100 ;
        RECT 397.950 754.650 400.050 756.750 ;
        RECT 403.950 754.950 406.050 758.400 ;
        RECT 458.400 756.750 459.600 758.400 ;
        RECT 457.950 754.650 460.050 756.750 ;
        RECT 467.400 756.600 468.600 758.400 ;
        RECT 479.400 759.000 484.050 759.600 ;
        RECT 479.400 758.400 483.600 759.000 ;
        RECT 479.400 756.600 480.600 758.400 ;
        RECT 467.400 755.400 480.600 756.600 ;
        RECT 484.950 756.600 487.050 757.050 ;
        RECT 497.400 756.600 498.600 760.950 ;
        RECT 521.400 756.750 522.600 761.400 ;
        RECT 523.950 760.950 526.050 763.050 ;
        RECT 556.950 762.600 559.050 763.050 ;
        RECT 565.950 762.600 568.050 763.050 ;
        RECT 577.950 762.600 580.050 763.050 ;
        RECT 600.000 762.600 604.050 763.050 ;
        RECT 556.950 761.400 564.600 762.600 ;
        RECT 556.950 760.950 559.050 761.400 ;
        RECT 524.400 757.050 525.600 760.950 ;
        RECT 563.400 759.600 564.600 761.400 ;
        RECT 565.950 761.400 580.050 762.600 ;
        RECT 565.950 760.950 568.050 761.400 ;
        RECT 577.950 760.950 580.050 761.400 ;
        RECT 599.400 760.950 604.050 762.600 ;
        RECT 610.800 760.950 612.900 763.050 ;
        RECT 613.950 762.600 616.050 763.050 ;
        RECT 613.950 761.400 627.600 762.600 ;
        RECT 613.950 760.950 616.050 761.400 ;
        RECT 563.400 759.000 576.600 759.600 ;
        RECT 563.400 758.400 577.050 759.000 ;
        RECT 484.950 755.400 498.600 756.600 ;
        RECT 499.950 756.600 502.050 756.750 ;
        RECT 520.950 756.600 523.050 756.750 ;
        RECT 499.950 755.400 523.050 756.600 ;
        RECT 524.400 755.400 529.050 757.050 ;
        RECT 484.950 754.950 487.050 755.400 ;
        RECT 499.950 754.650 502.050 755.400 ;
        RECT 520.950 754.650 523.050 755.400 ;
        RECT 525.000 754.950 529.050 755.400 ;
        RECT 538.950 756.600 541.050 756.900 ;
        RECT 547.950 756.600 550.050 757.050 ;
        RECT 538.950 755.400 550.050 756.600 ;
        RECT 538.950 754.800 541.050 755.400 ;
        RECT 547.950 754.950 550.050 755.400 ;
        RECT 574.950 754.950 577.050 758.400 ;
        RECT 586.950 756.600 589.050 756.750 ;
        RECT 599.400 756.600 600.600 760.950 ;
        RECT 611.250 757.050 612.450 760.950 ;
        RECT 626.400 757.050 627.600 761.400 ;
        RECT 634.950 760.950 637.050 763.050 ;
        RECT 655.950 762.600 658.050 763.200 ;
        RECT 653.400 761.400 658.050 762.600 ;
        RECT 586.950 755.400 600.600 756.600 ;
        RECT 586.950 754.650 589.050 755.400 ;
        RECT 610.800 754.950 612.900 757.050 ;
        RECT 625.950 754.950 628.050 757.050 ;
        RECT 4.950 753.600 7.050 754.050 ;
        RECT 19.950 753.600 22.050 754.050 ;
        RECT 28.950 753.600 31.050 754.050 ;
        RECT 4.950 752.400 31.050 753.600 ;
        RECT 4.950 751.950 7.050 752.400 ;
        RECT 19.950 751.950 22.050 752.400 ;
        RECT 28.950 751.950 31.050 752.400 ;
        RECT 106.950 753.600 109.050 754.050 ;
        RECT 115.950 753.600 118.050 754.050 ;
        RECT 148.950 753.600 151.050 754.050 ;
        RECT 277.950 753.600 280.050 754.050 ;
        RECT 106.950 752.400 151.050 753.600 ;
        RECT 106.950 751.950 109.050 752.400 ;
        RECT 115.950 751.950 118.050 752.400 ;
        RECT 148.950 751.950 151.050 752.400 ;
        RECT 269.400 752.400 280.050 753.600 ;
        RECT 269.400 751.050 270.600 752.400 ;
        RECT 277.950 751.950 280.050 752.400 ;
        RECT 316.950 753.600 319.050 754.050 ;
        RECT 347.400 753.600 348.600 754.650 ;
        RECT 635.400 754.050 636.600 760.950 ;
        RECT 653.400 759.600 654.600 761.400 ;
        RECT 655.950 761.100 658.050 761.400 ;
        RECT 676.950 762.600 679.050 763.200 ;
        RECT 705.000 762.600 709.050 763.050 ;
        RECT 676.950 761.400 684.600 762.600 ;
        RECT 676.950 761.100 679.050 761.400 ;
        RECT 647.400 758.400 654.600 759.600 ;
        RECT 683.400 759.600 684.600 761.400 ;
        RECT 704.400 760.950 709.050 762.600 ;
        RECT 712.950 762.600 717.000 763.050 ;
        RECT 712.950 760.950 717.600 762.600 ;
        RECT 727.950 760.950 730.050 763.050 ;
        RECT 739.950 762.600 742.050 763.050 ;
        RECT 748.950 762.600 751.050 763.050 ;
        RECT 737.400 761.400 751.050 762.600 ;
        RECT 683.400 758.400 696.600 759.600 ;
        RECT 640.950 756.600 643.050 756.750 ;
        RECT 647.400 756.600 648.600 758.400 ;
        RECT 640.950 755.400 648.600 756.600 ;
        RECT 649.950 756.450 652.050 756.900 ;
        RECT 664.950 756.450 667.050 756.900 ;
        RECT 640.950 754.650 643.050 755.400 ;
        RECT 649.950 755.250 667.050 756.450 ;
        RECT 695.400 756.600 696.600 758.400 ;
        RECT 704.400 756.900 705.600 760.950 ;
        RECT 716.400 756.900 717.600 760.950 ;
        RECT 728.400 757.050 729.600 760.950 ;
        RECT 695.400 756.000 702.600 756.600 ;
        RECT 695.400 755.400 703.050 756.000 ;
        RECT 649.950 754.800 652.050 755.250 ;
        RECT 664.950 754.800 667.050 755.250 ;
        RECT 451.950 753.600 454.050 754.050 ;
        RECT 316.950 752.400 348.600 753.600 ;
        RECT 416.400 752.400 454.050 753.600 ;
        RECT 316.950 751.950 319.050 752.400 ;
        RECT 40.950 750.600 43.050 751.050 ;
        RECT 55.950 750.600 58.050 751.050 ;
        RECT 40.950 749.400 58.050 750.600 ;
        RECT 40.950 748.950 43.050 749.400 ;
        RECT 55.950 748.950 58.050 749.400 ;
        RECT 166.950 750.600 169.050 751.050 ;
        RECT 196.950 750.600 199.050 751.050 ;
        RECT 166.950 749.400 199.050 750.600 ;
        RECT 166.950 748.950 169.050 749.400 ;
        RECT 196.950 748.950 199.050 749.400 ;
        RECT 238.950 750.600 241.050 751.050 ;
        RECT 268.950 750.600 271.050 751.050 ;
        RECT 238.950 749.400 271.050 750.600 ;
        RECT 238.950 748.950 241.050 749.400 ;
        RECT 268.950 748.950 271.050 749.400 ;
        RECT 280.950 750.600 283.050 751.050 ;
        RECT 358.950 750.600 361.050 751.050 ;
        RECT 280.950 749.400 361.050 750.600 ;
        RECT 280.950 748.950 283.050 749.400 ;
        RECT 358.950 748.950 361.050 749.400 ;
        RECT 373.950 750.600 376.050 751.050 ;
        RECT 403.950 750.600 406.050 751.050 ;
        RECT 416.400 750.600 417.600 752.400 ;
        RECT 451.950 751.950 454.050 752.400 ;
        RECT 460.950 753.600 463.050 754.050 ;
        RECT 496.950 753.600 499.050 754.050 ;
        RECT 460.950 752.400 499.050 753.600 ;
        RECT 460.950 751.950 463.050 752.400 ;
        RECT 496.950 751.950 499.050 752.400 ;
        RECT 502.950 753.600 505.050 754.050 ;
        RECT 517.950 753.600 520.050 754.050 ;
        RECT 502.950 752.400 520.050 753.600 ;
        RECT 502.950 751.950 505.050 752.400 ;
        RECT 517.950 751.950 520.050 752.400 ;
        RECT 598.950 753.600 601.050 754.050 ;
        RECT 631.950 753.600 634.050 754.050 ;
        RECT 598.950 752.400 634.050 753.600 ;
        RECT 635.400 752.400 640.050 754.050 ;
        RECT 598.950 751.950 601.050 752.400 ;
        RECT 631.950 751.950 634.050 752.400 ;
        RECT 636.000 751.950 640.050 752.400 ;
        RECT 700.950 751.950 703.050 755.400 ;
        RECT 703.950 754.800 706.050 756.900 ;
        RECT 715.950 754.800 718.050 756.900 ;
        RECT 727.950 754.950 730.050 757.050 ;
        RECT 733.950 756.600 736.050 756.750 ;
        RECT 737.400 756.600 738.600 761.400 ;
        RECT 739.950 760.950 742.050 761.400 ;
        RECT 748.950 760.950 751.050 761.400 ;
        RECT 763.950 762.600 766.050 763.050 ;
        RECT 769.950 762.600 772.050 763.050 ;
        RECT 793.800 762.600 795.900 763.050 ;
        RECT 763.950 761.400 772.050 762.600 ;
        RECT 763.950 760.950 766.050 761.400 ;
        RECT 769.950 760.950 772.050 761.400 ;
        RECT 788.400 761.400 795.900 762.600 ;
        RECT 733.950 755.400 738.600 756.600 ;
        RECT 757.950 756.600 760.050 756.750 ;
        RECT 766.950 756.600 769.050 757.050 ;
        RECT 772.950 756.600 775.050 756.750 ;
        RECT 757.950 755.400 775.050 756.600 ;
        RECT 733.950 754.650 736.050 755.400 ;
        RECT 757.950 754.650 760.050 755.400 ;
        RECT 766.950 754.950 769.050 755.400 ;
        RECT 772.950 754.650 775.050 755.400 ;
        RECT 778.950 756.600 781.050 756.750 ;
        RECT 788.400 756.600 789.600 761.400 ;
        RECT 793.800 760.950 795.900 761.400 ;
        RECT 796.950 759.600 799.050 762.900 ;
        RECT 820.950 760.950 823.050 764.400 ;
        RECT 829.950 759.600 832.050 763.050 ;
        RECT 841.950 760.950 844.050 763.050 ;
        RECT 853.950 762.600 856.050 763.200 ;
        RECT 848.400 761.400 856.050 762.600 ;
        RECT 796.950 759.000 834.600 759.600 ;
        RECT 797.400 758.400 834.600 759.000 ;
        RECT 778.950 755.400 789.600 756.600 ;
        RECT 778.950 754.650 781.050 755.400 ;
        RECT 736.950 753.600 739.050 754.050 ;
        RECT 742.950 753.600 745.050 754.050 ;
        RECT 751.950 753.600 754.050 754.050 ;
        RECT 736.950 752.400 754.050 753.600 ;
        RECT 833.400 753.600 834.600 758.400 ;
        RECT 842.400 757.050 843.600 760.950 ;
        RECT 848.400 757.050 849.600 761.400 ;
        RECT 853.950 761.100 856.050 761.400 ;
        RECT 841.950 754.950 844.050 757.050 ;
        RECT 847.950 754.950 850.050 757.050 ;
        RECT 848.400 753.600 849.600 754.950 ;
        RECT 833.400 752.400 849.600 753.600 ;
        RECT 736.950 751.950 739.050 752.400 ;
        RECT 742.950 751.950 745.050 752.400 ;
        RECT 751.950 751.950 754.050 752.400 ;
        RECT 373.950 749.400 406.050 750.600 ;
        RECT 373.950 748.950 376.050 749.400 ;
        RECT 403.950 748.950 406.050 749.400 ;
        RECT 407.400 749.400 417.600 750.600 ;
        RECT 424.950 750.600 427.050 751.050 ;
        RECT 439.950 750.600 442.050 751.050 ;
        RECT 457.800 750.600 459.900 751.050 ;
        RECT 424.950 749.400 459.900 750.600 ;
        RECT 73.950 747.600 76.050 748.050 ;
        RECT 94.950 747.600 97.050 748.050 ;
        RECT 124.950 747.600 127.050 748.050 ;
        RECT 73.950 746.400 127.050 747.600 ;
        RECT 73.950 745.950 76.050 746.400 ;
        RECT 94.950 745.950 97.050 746.400 ;
        RECT 124.950 745.950 127.050 746.400 ;
        RECT 154.950 747.600 157.050 748.050 ;
        RECT 167.400 747.600 168.600 748.950 ;
        RECT 154.950 746.400 168.600 747.600 ;
        RECT 337.950 747.600 340.050 748.050 ;
        RECT 364.950 747.600 367.050 748.050 ;
        RECT 337.950 746.400 367.050 747.600 ;
        RECT 154.950 745.950 157.050 746.400 ;
        RECT 337.950 745.950 340.050 746.400 ;
        RECT 364.950 745.950 367.050 746.400 ;
        RECT 394.950 747.600 397.050 748.050 ;
        RECT 407.400 747.600 408.600 749.400 ;
        RECT 424.950 748.950 427.050 749.400 ;
        RECT 439.950 748.950 442.050 749.400 ;
        RECT 457.800 748.950 459.900 749.400 ;
        RECT 460.950 750.600 463.050 750.900 ;
        RECT 490.950 750.600 493.050 751.050 ;
        RECT 511.950 750.600 514.050 750.900 ;
        RECT 460.950 749.400 493.050 750.600 ;
        RECT 460.950 748.800 463.050 749.400 ;
        RECT 490.950 748.950 493.050 749.400 ;
        RECT 494.400 749.400 514.050 750.600 ;
        RECT 394.950 746.400 408.600 747.600 ;
        RECT 436.950 747.600 439.050 748.050 ;
        RECT 448.950 747.600 451.050 748.050 ;
        RECT 494.400 747.600 495.600 749.400 ;
        RECT 511.950 748.800 514.050 749.400 ;
        RECT 529.950 750.600 532.050 751.050 ;
        RECT 559.950 750.600 562.050 751.050 ;
        RECT 580.800 750.600 582.900 751.050 ;
        RECT 529.950 749.400 537.600 750.600 ;
        RECT 529.950 748.950 532.050 749.400 ;
        RECT 436.950 746.400 451.050 747.600 ;
        RECT 394.950 745.950 397.050 746.400 ;
        RECT 436.950 745.950 439.050 746.400 ;
        RECT 448.950 745.950 451.050 746.400 ;
        RECT 452.400 746.400 495.600 747.600 ;
        RECT 517.950 747.600 520.050 748.050 ;
        RECT 526.950 747.600 529.050 748.050 ;
        RECT 532.950 747.600 535.050 748.050 ;
        RECT 517.950 746.400 535.050 747.600 ;
        RECT 536.400 747.600 537.600 749.400 ;
        RECT 559.950 749.400 582.900 750.600 ;
        RECT 559.950 748.950 562.050 749.400 ;
        RECT 580.800 748.950 582.900 749.400 ;
        RECT 583.950 750.600 586.050 751.050 ;
        RECT 616.950 750.600 619.050 751.050 ;
        RECT 583.950 749.400 619.050 750.600 ;
        RECT 583.950 748.950 586.050 749.400 ;
        RECT 616.950 748.950 619.050 749.400 ;
        RECT 661.950 750.600 664.050 751.050 ;
        RECT 679.950 750.600 682.050 751.050 ;
        RECT 685.950 750.600 688.050 751.050 ;
        RECT 661.950 749.400 688.050 750.600 ;
        RECT 661.950 748.950 664.050 749.400 ;
        RECT 679.950 748.950 682.050 749.400 ;
        RECT 685.950 748.950 688.050 749.400 ;
        RECT 748.950 750.600 751.050 751.050 ;
        RECT 763.950 750.600 766.050 751.050 ;
        RECT 787.950 750.600 790.050 751.050 ;
        RECT 748.950 749.400 790.050 750.600 ;
        RECT 748.950 748.950 751.050 749.400 ;
        RECT 763.950 748.950 766.050 749.400 ;
        RECT 787.950 748.950 790.050 749.400 ;
        RECT 799.950 750.600 802.050 751.050 ;
        RECT 826.950 750.600 829.050 751.050 ;
        RECT 832.950 750.600 835.050 751.050 ;
        RECT 799.950 749.400 835.050 750.600 ;
        RECT 799.950 748.950 802.050 749.400 ;
        RECT 826.950 748.950 829.050 749.400 ;
        RECT 832.950 748.950 835.050 749.400 ;
        RECT 550.950 747.600 553.050 748.050 ;
        RECT 536.400 746.400 553.050 747.600 ;
        RECT 34.950 744.600 37.050 745.050 ;
        RECT 49.950 744.600 52.050 745.050 ;
        RECT 34.950 743.400 52.050 744.600 ;
        RECT 34.950 742.950 37.050 743.400 ;
        RECT 49.950 742.950 52.050 743.400 ;
        RECT 103.950 744.600 106.050 745.050 ;
        RECT 118.950 744.600 121.050 745.050 ;
        RECT 103.950 743.400 121.050 744.600 ;
        RECT 103.950 742.950 106.050 743.400 ;
        RECT 118.950 742.950 121.050 743.400 ;
        RECT 304.950 744.600 307.050 745.050 ;
        RECT 328.950 744.600 331.050 745.050 ;
        RECT 304.950 743.400 331.050 744.600 ;
        RECT 304.950 742.950 307.050 743.400 ;
        RECT 328.950 742.950 331.050 743.400 ;
        RECT 412.950 744.600 415.050 745.050 ;
        RECT 421.950 744.600 424.050 745.050 ;
        RECT 452.400 744.600 453.600 746.400 ;
        RECT 517.950 745.950 520.050 746.400 ;
        RECT 526.950 745.950 529.050 746.400 ;
        RECT 532.950 745.950 535.050 746.400 ;
        RECT 550.950 745.950 553.050 746.400 ;
        RECT 562.950 747.600 565.050 748.050 ;
        RECT 580.950 747.600 583.050 747.900 ;
        RECT 562.950 746.400 583.050 747.600 ;
        RECT 562.950 745.950 565.050 746.400 ;
        RECT 580.950 745.800 583.050 746.400 ;
        RECT 604.950 747.600 607.050 748.050 ;
        RECT 622.950 747.600 625.050 748.050 ;
        RECT 604.950 746.400 625.050 747.600 ;
        RECT 604.950 745.950 607.050 746.400 ;
        RECT 622.950 745.950 625.050 746.400 ;
        RECT 658.950 747.600 661.050 748.050 ;
        RECT 673.950 747.600 676.050 748.050 ;
        RECT 658.950 746.400 676.050 747.600 ;
        RECT 658.950 745.950 661.050 746.400 ;
        RECT 673.950 745.950 676.050 746.400 ;
        RECT 697.950 747.600 700.050 748.050 ;
        RECT 718.950 747.600 721.050 748.050 ;
        RECT 739.950 747.600 742.050 748.050 ;
        RECT 697.950 746.400 742.050 747.600 ;
        RECT 697.950 745.950 700.050 746.400 ;
        RECT 718.950 745.950 721.050 746.400 ;
        RECT 739.950 745.950 742.050 746.400 ;
        RECT 412.950 743.400 453.600 744.600 ;
        RECT 457.950 744.600 460.050 745.050 ;
        RECT 466.950 744.600 469.050 745.050 ;
        RECT 478.950 744.600 481.050 745.050 ;
        RECT 457.950 743.400 481.050 744.600 ;
        RECT 412.950 742.950 415.050 743.400 ;
        RECT 421.950 742.950 424.050 743.400 ;
        RECT 457.950 742.950 460.050 743.400 ;
        RECT 466.950 742.950 469.050 743.400 ;
        RECT 478.950 742.950 481.050 743.400 ;
        RECT 484.950 744.600 487.050 745.050 ;
        RECT 502.950 744.600 505.050 745.050 ;
        RECT 484.950 743.400 505.050 744.600 ;
        RECT 484.950 742.950 487.050 743.400 ;
        RECT 502.950 742.950 505.050 743.400 ;
        RECT 508.950 744.600 511.050 745.050 ;
        RECT 559.950 744.600 562.050 745.050 ;
        RECT 508.950 743.400 562.050 744.600 ;
        RECT 508.950 742.950 511.050 743.400 ;
        RECT 559.950 742.950 562.050 743.400 ;
        RECT 583.950 744.600 586.050 745.050 ;
        RECT 625.950 744.600 628.050 745.050 ;
        RECT 583.950 743.400 628.050 744.600 ;
        RECT 583.950 742.950 586.050 743.400 ;
        RECT 625.950 742.950 628.050 743.400 ;
        RECT 1.950 741.600 4.050 742.050 ;
        RECT 10.950 741.600 13.050 742.050 ;
        RECT 1.950 740.400 13.050 741.600 ;
        RECT 1.950 739.950 4.050 740.400 ;
        RECT 10.950 739.950 13.050 740.400 ;
        RECT 16.950 741.600 19.050 742.050 ;
        RECT 31.950 741.600 34.050 742.050 ;
        RECT 52.950 741.600 55.050 742.050 ;
        RECT 16.950 740.400 55.050 741.600 ;
        RECT 16.950 739.950 19.050 740.400 ;
        RECT 31.950 739.950 34.050 740.400 ;
        RECT 52.950 739.950 55.050 740.400 ;
        RECT 124.950 741.600 127.050 742.050 ;
        RECT 139.950 741.600 142.050 742.050 ;
        RECT 124.950 740.400 142.050 741.600 ;
        RECT 124.950 739.950 127.050 740.400 ;
        RECT 139.950 739.950 142.050 740.400 ;
        RECT 214.950 741.600 217.050 742.050 ;
        RECT 235.950 741.600 238.050 742.050 ;
        RECT 331.950 741.600 334.050 742.050 ;
        RECT 214.950 740.400 334.050 741.600 ;
        RECT 214.950 739.950 217.050 740.400 ;
        RECT 235.950 739.950 238.050 740.400 ;
        RECT 331.950 739.950 334.050 740.400 ;
        RECT 346.950 741.600 349.050 742.050 ;
        RECT 367.950 741.600 370.050 742.050 ;
        RECT 346.950 740.400 370.050 741.600 ;
        RECT 346.950 739.950 349.050 740.400 ;
        RECT 367.950 739.950 370.050 740.400 ;
        RECT 430.950 741.600 433.050 742.050 ;
        RECT 472.950 741.600 475.050 742.050 ;
        RECT 430.950 740.400 475.050 741.600 ;
        RECT 430.950 739.950 433.050 740.400 ;
        RECT 472.950 739.950 475.050 740.400 ;
        RECT 511.950 741.600 514.050 742.050 ;
        RECT 586.950 741.600 589.050 742.050 ;
        RECT 823.950 741.600 826.050 742.050 ;
        RECT 829.950 741.600 832.050 742.050 ;
        RECT 511.950 740.400 549.600 741.600 ;
        RECT 511.950 739.950 514.050 740.400 ;
        RECT 88.950 738.600 91.050 739.050 ;
        RECT 59.400 737.400 91.050 738.600 ;
        RECT 59.400 736.050 60.600 737.400 ;
        RECT 88.950 736.950 91.050 737.400 ;
        RECT 235.950 738.600 238.050 738.900 ;
        RECT 247.950 738.600 250.050 739.050 ;
        RECT 235.950 737.400 250.050 738.600 ;
        RECT 235.950 736.800 238.050 737.400 ;
        RECT 247.950 736.950 250.050 737.400 ;
        RECT 289.950 738.600 292.050 739.050 ;
        RECT 295.950 738.600 298.050 739.050 ;
        RECT 289.950 737.400 298.050 738.600 ;
        RECT 289.950 736.950 292.050 737.400 ;
        RECT 295.950 736.950 298.050 737.400 ;
        RECT 349.950 738.600 352.050 739.050 ;
        RECT 370.950 738.600 373.050 739.050 ;
        RECT 376.950 738.600 379.050 739.050 ;
        RECT 349.950 737.400 379.050 738.600 ;
        RECT 349.950 736.950 352.050 737.400 ;
        RECT 370.950 736.950 373.050 737.400 ;
        RECT 376.950 736.950 379.050 737.400 ;
        RECT 514.950 738.600 517.050 739.050 ;
        RECT 523.800 738.600 525.900 739.050 ;
        RECT 514.950 737.400 525.900 738.600 ;
        RECT 548.400 738.600 549.600 740.400 ;
        RECT 586.950 740.400 624.600 741.600 ;
        RECT 586.950 739.950 589.050 740.400 ;
        RECT 562.950 738.600 565.050 739.050 ;
        RECT 548.400 737.400 565.050 738.600 ;
        RECT 514.950 736.950 517.050 737.400 ;
        RECT 523.800 736.950 525.900 737.400 ;
        RECT 562.950 736.950 565.050 737.400 ;
        RECT 580.950 738.600 583.050 739.050 ;
        RECT 607.950 738.600 610.050 739.050 ;
        RECT 580.950 737.400 610.050 738.600 ;
        RECT 623.400 738.600 624.600 740.400 ;
        RECT 823.950 740.400 832.050 741.600 ;
        RECT 823.950 739.950 826.050 740.400 ;
        RECT 829.950 739.950 832.050 740.400 ;
        RECT 634.950 738.600 637.050 739.050 ;
        RECT 623.400 737.400 637.050 738.600 ;
        RECT 580.950 736.950 583.050 737.400 ;
        RECT 607.950 736.950 610.050 737.400 ;
        RECT 634.950 736.950 637.050 737.400 ;
        RECT 688.950 738.600 691.050 739.050 ;
        RECT 739.950 738.600 742.050 739.050 ;
        RECT 688.950 737.400 742.050 738.600 ;
        RECT 688.950 736.950 691.050 737.400 ;
        RECT 739.950 736.950 742.050 737.400 ;
        RECT 820.950 738.600 823.050 739.050 ;
        RECT 838.950 738.600 841.050 739.050 ;
        RECT 820.950 737.400 841.050 738.600 ;
        RECT 820.950 736.950 823.050 737.400 ;
        RECT 838.950 736.950 841.050 737.400 ;
        RECT 46.950 735.600 49.050 736.050 ;
        RECT 58.950 735.600 61.050 736.050 ;
        RECT 46.950 734.400 61.050 735.600 ;
        RECT 46.950 733.950 49.050 734.400 ;
        RECT 58.950 733.950 61.050 734.400 ;
        RECT 70.950 735.600 73.050 736.050 ;
        RECT 79.950 735.600 82.050 736.050 ;
        RECT 70.950 734.400 82.050 735.600 ;
        RECT 70.950 733.950 73.050 734.400 ;
        RECT 79.950 733.950 82.050 734.400 ;
        RECT 118.950 735.600 121.050 736.050 ;
        RECT 157.950 735.600 160.050 736.050 ;
        RECT 181.950 735.600 184.050 736.050 ;
        RECT 118.950 734.400 184.050 735.600 ;
        RECT 118.950 733.950 121.050 734.400 ;
        RECT 157.950 733.950 160.050 734.400 ;
        RECT 181.950 733.950 184.050 734.400 ;
        RECT 229.950 735.600 232.050 736.050 ;
        RECT 250.950 735.600 253.050 736.050 ;
        RECT 262.950 735.600 265.050 736.050 ;
        RECT 229.950 734.400 265.050 735.600 ;
        RECT 229.950 733.950 232.050 734.400 ;
        RECT 250.950 733.950 253.050 734.400 ;
        RECT 262.950 733.950 265.050 734.400 ;
        RECT 274.950 735.600 277.050 736.050 ;
        RECT 283.950 735.600 286.050 736.050 ;
        RECT 316.950 735.600 319.050 736.050 ;
        RECT 274.950 734.400 319.050 735.600 ;
        RECT 274.950 733.950 277.050 734.400 ;
        RECT 283.950 733.950 286.050 734.400 ;
        RECT 316.950 733.950 319.050 734.400 ;
        RECT 328.950 735.600 331.050 736.050 ;
        RECT 358.950 735.600 361.050 736.050 ;
        RECT 328.950 734.400 361.050 735.600 ;
        RECT 328.950 733.950 331.050 734.400 ;
        RECT 358.950 733.950 361.050 734.400 ;
        RECT 388.950 735.600 391.050 736.050 ;
        RECT 406.950 735.600 409.050 736.050 ;
        RECT 388.950 734.400 409.050 735.600 ;
        RECT 388.950 733.950 391.050 734.400 ;
        RECT 406.950 733.950 409.050 734.400 ;
        RECT 445.950 735.600 448.050 736.050 ;
        RECT 475.950 735.600 478.050 736.050 ;
        RECT 445.950 734.400 478.050 735.600 ;
        RECT 445.950 733.950 448.050 734.400 ;
        RECT 475.950 733.950 478.050 734.400 ;
        RECT 487.950 735.600 490.050 736.050 ;
        RECT 511.950 735.600 514.050 736.050 ;
        RECT 487.950 734.400 514.050 735.600 ;
        RECT 487.950 733.950 490.050 734.400 ;
        RECT 511.950 733.950 514.050 734.400 ;
        RECT 574.950 735.600 577.050 736.050 ;
        RECT 586.950 735.600 589.050 736.050 ;
        RECT 610.950 735.600 613.050 736.050 ;
        RECT 574.950 734.400 589.050 735.600 ;
        RECT 574.950 733.950 577.050 734.400 ;
        RECT 586.950 733.950 589.050 734.400 ;
        RECT 593.400 734.400 613.050 735.600 ;
        RECT 4.950 732.600 7.050 733.050 ;
        RECT 13.950 732.600 16.050 733.050 ;
        RECT 4.950 731.400 16.050 732.600 ;
        RECT 4.950 730.950 7.050 731.400 ;
        RECT 13.950 730.950 16.050 731.400 ;
        RECT 55.950 730.950 58.050 733.050 ;
        RECT 61.950 732.600 64.050 733.050 ;
        RECT 67.950 732.600 70.050 733.050 ;
        RECT 61.950 731.400 70.050 732.600 ;
        RECT 61.950 730.950 64.050 731.400 ;
        RECT 67.950 730.950 70.050 731.400 ;
        RECT 301.950 732.600 304.050 733.050 ;
        RECT 310.950 732.600 313.050 733.050 ;
        RECT 301.950 731.400 313.050 732.600 ;
        RECT 301.950 730.950 304.050 731.400 ;
        RECT 310.950 730.950 313.050 731.400 ;
        RECT 400.950 732.600 403.050 733.050 ;
        RECT 409.950 732.600 412.050 733.050 ;
        RECT 400.950 731.400 412.050 732.600 ;
        RECT 400.950 730.950 403.050 731.400 ;
        RECT 409.950 730.950 412.050 731.400 ;
        RECT 454.950 732.600 457.050 733.050 ;
        RECT 460.950 732.600 463.050 733.050 ;
        RECT 454.950 731.400 463.050 732.600 ;
        RECT 454.950 730.950 457.050 731.400 ;
        RECT 460.950 730.950 463.050 731.400 ;
        RECT 532.950 732.600 535.050 733.050 ;
        RECT 553.950 732.600 556.050 733.050 ;
        RECT 532.950 731.400 556.050 732.600 ;
        RECT 532.950 730.950 535.050 731.400 ;
        RECT 553.950 730.950 556.050 731.400 ;
        RECT 559.950 732.600 562.050 733.050 ;
        RECT 593.400 732.600 594.600 734.400 ;
        RECT 610.950 733.950 613.050 734.400 ;
        RECT 700.950 735.600 703.050 736.050 ;
        RECT 742.950 735.600 745.050 736.050 ;
        RECT 700.950 734.400 745.050 735.600 ;
        RECT 700.950 733.950 703.050 734.400 ;
        RECT 742.950 733.950 745.050 734.400 ;
        RECT 757.950 735.600 760.050 736.050 ;
        RECT 772.950 735.600 775.050 736.050 ;
        RECT 757.950 734.400 775.050 735.600 ;
        RECT 757.950 733.950 760.050 734.400 ;
        RECT 772.950 733.950 775.050 734.400 ;
        RECT 799.950 735.600 802.050 736.050 ;
        RECT 814.950 735.600 817.050 736.050 ;
        RECT 799.950 734.400 817.050 735.600 ;
        RECT 799.950 733.950 802.050 734.400 ;
        RECT 814.950 733.950 817.050 734.400 ;
        RECT 559.950 731.400 594.600 732.600 ;
        RECT 595.950 732.600 598.050 733.050 ;
        RECT 784.950 732.600 787.050 733.050 ;
        RECT 793.950 732.600 796.050 733.050 ;
        RECT 823.950 732.600 826.050 733.050 ;
        RECT 835.950 732.600 838.050 733.050 ;
        RECT 595.950 731.400 603.600 732.600 ;
        RECT 559.950 730.950 562.050 731.400 ;
        RECT 595.950 730.950 598.050 731.400 ;
        RECT 37.950 729.600 40.050 730.350 ;
        RECT 49.950 729.600 54.000 730.050 ;
        RECT 37.950 728.400 42.600 729.600 ;
        RECT 37.950 728.250 40.050 728.400 ;
        RECT 41.400 724.050 42.600 728.400 ;
        RECT 49.950 727.950 54.600 729.600 ;
        RECT 53.400 724.050 54.600 727.950 ;
        RECT 4.950 723.600 7.050 724.050 ;
        RECT 13.950 723.600 16.050 724.050 ;
        RECT 28.950 723.600 31.050 724.050 ;
        RECT 4.950 722.400 31.050 723.600 ;
        RECT 4.950 721.950 7.050 722.400 ;
        RECT 13.950 721.950 16.050 722.400 ;
        RECT 28.950 721.950 31.050 722.400 ;
        RECT 40.950 721.950 43.050 724.050 ;
        RECT 52.950 721.950 55.050 724.050 ;
        RECT 31.950 720.600 34.050 721.050 ;
        RECT 56.400 720.600 57.600 730.950 ;
        RECT 73.950 728.250 76.050 730.350 ;
        RECT 79.950 729.600 82.050 730.350 ;
        RECT 94.950 729.600 97.050 730.350 ;
        RECT 79.950 728.400 97.050 729.600 ;
        RECT 79.950 728.250 82.050 728.400 ;
        RECT 94.950 728.250 97.050 728.400 ;
        RECT 109.950 729.600 112.050 730.050 ;
        RECT 118.950 729.600 121.050 730.200 ;
        RECT 109.950 728.400 121.050 729.600 ;
        RECT 74.400 724.050 75.600 728.250 ;
        RECT 109.950 727.950 112.050 728.400 ;
        RECT 118.950 728.100 121.050 728.400 ;
        RECT 124.950 729.600 127.050 730.200 ;
        RECT 130.950 729.600 133.050 730.050 ;
        RECT 124.950 728.400 133.050 729.600 ;
        RECT 124.950 728.100 127.050 728.400 ;
        RECT 130.950 727.950 133.050 728.400 ;
        RECT 145.950 728.100 148.050 730.200 ;
        RECT 166.950 729.600 169.050 730.050 ;
        RECT 175.950 729.600 178.050 730.050 ;
        RECT 193.950 729.600 196.050 730.350 ;
        RECT 214.950 729.600 217.050 730.350 ;
        RECT 166.950 728.400 178.050 729.600 ;
        RECT 73.950 721.950 76.050 724.050 ;
        RECT 88.950 723.450 91.050 723.900 ;
        RECT 136.950 723.450 139.050 723.900 ;
        RECT 88.950 722.250 139.050 723.450 ;
        RECT 88.950 721.800 91.050 722.250 ;
        RECT 136.950 721.800 139.050 722.250 ;
        RECT 146.400 721.050 147.600 728.100 ;
        RECT 166.950 727.950 169.050 728.400 ;
        RECT 175.950 727.950 178.050 728.400 ;
        RECT 188.400 728.400 217.050 729.600 ;
        RECT 188.400 724.050 189.600 728.400 ;
        RECT 193.950 728.250 196.050 728.400 ;
        RECT 214.950 728.250 217.050 728.400 ;
        RECT 220.950 729.900 223.050 730.350 ;
        RECT 226.950 729.900 229.050 730.350 ;
        RECT 220.950 728.700 229.050 729.900 ;
        RECT 220.950 728.250 223.050 728.700 ;
        RECT 226.950 728.250 229.050 728.700 ;
        RECT 241.950 729.600 244.050 730.350 ;
        RECT 247.950 729.600 250.050 730.050 ;
        RECT 241.950 728.400 250.050 729.600 ;
        RECT 241.950 728.250 244.050 728.400 ;
        RECT 247.950 727.950 250.050 728.400 ;
        RECT 256.950 728.250 259.050 730.350 ;
        RECT 274.800 729.600 276.900 730.050 ;
        RECT 266.250 728.400 276.900 729.600 ;
        RECT 257.400 724.050 258.600 728.250 ;
        RECT 266.250 724.050 267.450 728.400 ;
        RECT 274.800 727.950 276.900 728.400 ;
        RECT 277.950 728.250 280.050 730.350 ;
        RECT 278.400 726.600 279.600 728.250 ;
        RECT 289.800 727.950 291.900 730.050 ;
        RECT 295.950 728.100 298.050 730.200 ;
        RECT 316.950 729.600 319.050 730.200 ;
        RECT 305.400 728.400 319.050 729.600 ;
        RECT 269.400 726.000 279.600 726.600 ;
        RECT 268.950 725.400 279.600 726.000 ;
        RECT 187.950 721.950 190.050 724.050 ;
        RECT 208.950 723.600 211.050 724.050 ;
        RECT 217.950 723.600 220.050 724.050 ;
        RECT 208.950 722.400 220.050 723.600 ;
        RECT 208.950 721.950 211.050 722.400 ;
        RECT 217.950 721.950 220.050 722.400 ;
        RECT 256.950 721.950 259.050 724.050 ;
        RECT 265.800 721.950 267.900 724.050 ;
        RECT 268.950 721.950 271.050 725.400 ;
        RECT 290.250 724.050 291.450 727.950 ;
        RECT 296.400 724.050 297.600 728.100 ;
        RECT 289.800 721.950 291.900 724.050 ;
        RECT 292.950 722.400 297.600 724.050 ;
        RECT 305.400 723.900 306.600 728.400 ;
        RECT 316.950 728.100 319.050 728.400 ;
        RECT 325.950 729.900 328.050 730.350 ;
        RECT 334.950 729.900 337.050 730.350 ;
        RECT 325.950 728.700 337.050 729.900 ;
        RECT 325.950 728.250 328.050 728.700 ;
        RECT 334.950 728.250 337.050 728.700 ;
        RECT 340.950 729.600 343.050 730.350 ;
        RECT 373.950 729.600 376.050 730.050 ;
        RECT 379.950 729.600 382.050 730.200 ;
        RECT 385.950 729.600 388.050 730.200 ;
        RECT 394.950 729.600 397.050 730.200 ;
        RECT 340.950 728.400 378.600 729.600 ;
        RECT 340.950 728.250 343.050 728.400 ;
        RECT 373.950 727.950 376.050 728.400 ;
        RECT 292.950 721.950 297.000 722.400 ;
        RECT 304.950 721.800 307.050 723.900 ;
        RECT 319.950 723.600 322.050 723.900 ;
        RECT 337.950 723.600 340.050 724.050 ;
        RECT 377.400 723.900 378.600 728.400 ;
        RECT 379.950 728.400 384.600 729.600 ;
        RECT 379.950 728.100 382.050 728.400 ;
        RECT 383.400 726.600 384.600 728.400 ;
        RECT 385.950 728.400 397.050 729.600 ;
        RECT 385.950 728.100 388.050 728.400 ;
        RECT 394.950 728.100 397.050 728.400 ;
        RECT 412.950 729.600 415.050 730.050 ;
        RECT 418.950 729.600 421.050 730.350 ;
        RECT 430.950 729.600 433.050 730.050 ;
        RECT 412.950 728.400 421.050 729.600 ;
        RECT 412.950 727.950 415.050 728.400 ;
        RECT 418.950 728.250 421.050 728.400 ;
        RECT 422.400 728.400 433.050 729.600 ;
        RECT 383.400 726.000 390.600 726.600 ;
        RECT 383.400 725.400 391.050 726.000 ;
        RECT 319.950 722.400 340.050 723.600 ;
        RECT 319.950 721.800 322.050 722.400 ;
        RECT 337.950 721.950 340.050 722.400 ;
        RECT 349.950 723.450 352.050 723.900 ;
        RECT 355.950 723.450 358.050 723.900 ;
        RECT 349.950 722.250 358.050 723.450 ;
        RECT 349.950 721.800 352.050 722.250 ;
        RECT 355.950 721.800 358.050 722.250 ;
        RECT 376.950 721.800 379.050 723.900 ;
        RECT 388.950 721.950 391.050 725.400 ;
        RECT 422.400 724.050 423.600 728.400 ;
        RECT 430.950 727.950 433.050 728.400 ;
        RECT 457.950 727.950 460.050 730.050 ;
        RECT 463.950 728.250 466.050 730.350 ;
        RECT 520.950 729.600 523.050 730.200 ;
        RECT 503.400 728.400 523.050 729.600 ;
        RECT 458.400 724.050 459.600 727.950 ;
        RECT 421.950 721.950 424.050 724.050 ;
        RECT 458.400 722.400 463.050 724.050 ;
        RECT 464.400 723.600 465.600 728.250 ;
        RECT 487.950 723.600 490.050 724.050 ;
        RECT 503.400 723.900 504.600 728.400 ;
        RECT 520.950 728.100 523.050 728.400 ;
        RECT 535.950 729.600 538.050 730.200 ;
        RECT 547.950 729.600 550.050 730.050 ;
        RECT 535.950 728.400 540.600 729.600 ;
        RECT 535.950 728.100 538.050 728.400 ;
        RECT 464.400 722.400 490.050 723.600 ;
        RECT 459.000 721.950 463.050 722.400 ;
        RECT 487.950 721.950 490.050 722.400 ;
        RECT 82.950 720.600 85.050 721.050 ;
        RECT 31.950 719.400 85.050 720.600 ;
        RECT 31.950 718.950 34.050 719.400 ;
        RECT 82.950 718.950 85.050 719.400 ;
        RECT 145.950 718.950 148.050 721.050 ;
        RECT 250.950 720.600 253.050 721.050 ;
        RECT 286.950 720.600 289.050 721.050 ;
        RECT 325.950 720.600 328.050 721.050 ;
        RECT 152.400 719.400 237.600 720.600 ;
        RECT 46.950 717.600 49.050 718.050 ;
        RECT 70.950 717.600 73.050 718.050 ;
        RECT 46.950 716.400 73.050 717.600 ;
        RECT 46.950 715.950 49.050 716.400 ;
        RECT 70.950 715.950 73.050 716.400 ;
        RECT 76.950 717.600 79.050 718.050 ;
        RECT 91.950 717.600 94.050 718.050 ;
        RECT 76.950 716.400 94.050 717.600 ;
        RECT 76.950 715.950 79.050 716.400 ;
        RECT 91.950 715.950 94.050 716.400 ;
        RECT 97.950 717.600 100.050 717.900 ;
        RECT 115.950 717.600 118.050 718.050 ;
        RECT 97.950 716.400 118.050 717.600 ;
        RECT 97.950 715.800 100.050 716.400 ;
        RECT 115.950 715.950 118.050 716.400 ;
        RECT 142.950 717.600 145.050 718.050 ;
        RECT 148.950 717.600 151.050 718.050 ;
        RECT 152.400 717.600 153.600 719.400 ;
        RECT 142.950 716.400 153.600 717.600 ;
        RECT 236.400 717.600 237.600 719.400 ;
        RECT 250.950 719.400 328.050 720.600 ;
        RECT 422.400 720.600 423.600 721.950 ;
        RECT 502.950 721.800 505.050 723.900 ;
        RECT 436.950 720.600 439.050 721.050 ;
        RECT 422.400 719.400 439.050 720.600 ;
        RECT 250.950 718.950 253.050 719.400 ;
        RECT 286.950 718.950 289.050 719.400 ;
        RECT 325.950 718.950 328.050 719.400 ;
        RECT 436.950 718.950 439.050 719.400 ;
        RECT 457.950 720.600 460.050 721.050 ;
        RECT 514.950 720.600 517.050 721.050 ;
        RECT 457.950 719.400 517.050 720.600 ;
        RECT 539.400 720.600 540.600 728.400 ;
        RECT 542.400 728.400 550.050 729.600 ;
        RECT 542.400 724.050 543.600 728.400 ;
        RECT 547.950 727.950 550.050 728.400 ;
        RECT 556.950 728.100 559.050 730.200 ;
        RECT 574.950 728.250 577.050 730.350 ;
        RECT 583.950 729.600 586.050 730.050 ;
        RECT 578.400 728.400 586.050 729.600 ;
        RECT 557.400 726.600 558.600 728.100 ;
        RECT 557.400 726.000 573.600 726.600 ;
        RECT 557.400 725.400 574.050 726.000 ;
        RECT 541.950 721.950 544.050 724.050 ;
        RECT 553.950 723.600 556.050 723.900 ;
        RECT 562.950 723.600 565.050 724.050 ;
        RECT 553.950 722.400 565.050 723.600 ;
        RECT 553.950 721.800 556.050 722.400 ;
        RECT 562.950 721.950 565.050 722.400 ;
        RECT 571.950 721.950 574.050 725.400 ;
        RECT 575.400 720.600 576.600 728.250 ;
        RECT 578.400 724.050 579.600 728.400 ;
        RECT 583.950 727.950 586.050 728.400 ;
        RECT 602.400 724.050 603.600 731.400 ;
        RECT 784.950 731.400 792.600 732.600 ;
        RECT 784.950 730.950 787.050 731.400 ;
        RECT 616.950 729.600 619.050 730.200 ;
        RECT 649.950 729.750 652.050 730.200 ;
        RECT 682.950 729.750 685.050 730.200 ;
        RECT 616.950 728.400 621.600 729.600 ;
        RECT 616.950 728.100 619.050 728.400 ;
        RECT 577.950 721.950 580.050 724.050 ;
        RECT 583.950 723.600 586.050 724.050 ;
        RECT 601.950 723.600 604.050 724.050 ;
        RECT 583.950 722.400 604.050 723.600 ;
        RECT 620.400 723.600 621.600 728.400 ;
        RECT 649.950 728.550 685.050 729.750 ;
        RECT 649.950 728.100 652.050 728.550 ;
        RECT 682.950 728.100 685.050 728.550 ;
        RECT 706.950 729.600 709.050 730.200 ;
        RECT 715.950 729.600 718.050 730.050 ;
        RECT 706.950 728.400 718.050 729.600 ;
        RECT 706.950 728.100 709.050 728.400 ;
        RECT 715.950 727.950 718.050 728.400 ;
        RECT 724.950 728.250 727.050 730.350 ;
        RECT 725.400 724.050 726.600 728.250 ;
        RECT 736.800 727.950 738.900 730.050 ;
        RECT 739.950 729.600 742.050 730.050 ;
        RECT 748.950 729.600 751.050 730.200 ;
        RECT 766.950 729.600 769.050 730.350 ;
        RECT 739.950 728.400 747.600 729.600 ;
        RECT 739.950 727.950 742.050 728.400 ;
        RECT 737.250 724.050 738.450 727.950 ;
        RECT 640.800 723.600 642.900 723.900 ;
        RECT 620.400 722.400 642.900 723.600 ;
        RECT 583.950 721.950 586.050 722.400 ;
        RECT 601.950 721.950 604.050 722.400 ;
        RECT 640.800 721.800 642.900 722.400 ;
        RECT 670.950 723.600 673.050 723.900 ;
        RECT 679.950 723.600 682.050 723.900 ;
        RECT 670.950 722.400 682.050 723.600 ;
        RECT 670.950 721.800 673.050 722.400 ;
        RECT 679.950 721.800 682.050 722.400 ;
        RECT 709.950 723.450 712.050 723.900 ;
        RECT 718.950 723.450 721.050 723.900 ;
        RECT 709.950 722.250 721.050 723.450 ;
        RECT 709.950 721.800 712.050 722.250 ;
        RECT 718.950 721.800 721.050 722.250 ;
        RECT 724.950 721.950 727.050 724.050 ;
        RECT 733.950 722.400 738.450 724.050 ;
        RECT 746.400 723.900 747.600 728.400 ;
        RECT 748.950 728.400 756.600 729.600 ;
        RECT 748.950 728.100 751.050 728.400 ;
        RECT 733.950 721.950 738.000 722.400 ;
        RECT 539.400 719.400 576.600 720.600 ;
        RECT 625.950 720.600 628.050 721.050 ;
        RECT 637.950 720.600 640.050 720.750 ;
        RECT 625.950 719.400 640.050 720.600 ;
        RECT 457.950 718.950 460.050 719.400 ;
        RECT 514.950 718.950 517.050 719.400 ;
        RECT 625.950 718.950 628.050 719.400 ;
        RECT 637.950 718.650 640.050 719.400 ;
        RECT 721.950 720.600 724.050 721.050 ;
        RECT 734.400 720.600 735.600 721.950 ;
        RECT 745.950 721.800 748.050 723.900 ;
        RECT 755.400 723.600 756.600 728.400 ;
        RECT 766.950 728.400 777.600 729.600 ;
        RECT 766.950 728.250 769.050 728.400 ;
        RECT 776.400 727.050 777.600 728.400 ;
        RECT 781.950 727.950 784.050 730.050 ;
        RECT 776.400 725.400 781.050 727.050 ;
        RECT 777.000 724.950 781.050 725.400 ;
        RECT 763.950 723.600 766.050 724.050 ;
        RECT 755.400 722.400 766.050 723.600 ;
        RECT 763.950 721.950 766.050 722.400 ;
        RECT 772.950 723.600 775.050 724.050 ;
        RECT 782.400 723.600 783.600 727.950 ;
        RECT 791.400 724.050 792.600 731.400 ;
        RECT 793.950 731.400 838.050 732.600 ;
        RECT 793.950 730.950 796.050 731.400 ;
        RECT 823.950 730.950 826.050 731.400 ;
        RECT 835.950 730.950 838.050 731.400 ;
        RECT 850.950 730.950 853.050 733.050 ;
        RECT 796.950 729.600 801.000 730.050 ;
        RECT 802.950 729.600 805.050 730.050 ;
        RECT 811.950 729.600 814.050 730.200 ;
        RECT 796.950 727.950 801.600 729.600 ;
        RECT 802.950 728.400 814.050 729.600 ;
        RECT 802.950 727.950 805.050 728.400 ;
        RECT 811.950 728.100 814.050 728.400 ;
        RECT 820.950 727.950 823.050 730.050 ;
        RECT 826.950 729.600 829.050 730.050 ;
        RECT 840.000 729.600 844.050 730.050 ;
        RECT 826.950 728.400 837.450 729.600 ;
        RECT 826.950 727.950 829.050 728.400 ;
        RECT 772.950 722.400 783.600 723.600 ;
        RECT 772.950 721.950 775.050 722.400 ;
        RECT 790.950 721.950 793.050 724.050 ;
        RECT 721.950 719.400 735.600 720.600 ;
        RECT 769.950 720.600 772.050 721.050 ;
        RECT 791.400 720.600 792.600 721.950 ;
        RECT 769.950 719.400 792.600 720.600 ;
        RECT 800.400 720.600 801.600 727.950 ;
        RECT 821.400 724.050 822.600 727.950 ;
        RECT 836.250 724.050 837.450 728.400 ;
        RECT 839.400 727.950 844.050 729.600 ;
        RECT 839.400 724.050 840.600 727.950 ;
        RECT 851.400 726.600 852.600 730.950 ;
        RECT 853.950 729.600 856.050 730.200 ;
        RECT 853.950 728.400 861.600 729.600 ;
        RECT 853.950 728.100 856.050 728.400 ;
        RECT 848.400 725.400 852.600 726.600 ;
        RECT 848.400 724.050 849.600 725.400 ;
        RECT 860.400 724.050 861.600 728.400 ;
        RECT 820.950 721.950 823.050 724.050 ;
        RECT 835.800 721.950 837.900 724.050 ;
        RECT 838.950 721.950 841.050 724.050 ;
        RECT 844.950 722.400 849.600 724.050 ;
        RECT 844.950 721.950 849.000 722.400 ;
        RECT 859.950 721.950 862.050 724.050 ;
        RECT 814.950 720.600 817.050 721.050 ;
        RECT 800.400 719.400 817.050 720.600 ;
        RECT 721.950 718.950 724.050 719.400 ;
        RECT 769.950 718.950 772.050 719.400 ;
        RECT 814.950 718.950 817.050 719.400 ;
        RECT 823.950 720.600 826.050 721.050 ;
        RECT 856.950 720.600 859.050 721.050 ;
        RECT 823.950 719.400 859.050 720.600 ;
        RECT 823.950 718.950 826.050 719.400 ;
        RECT 856.950 718.950 859.050 719.400 ;
        RECT 241.950 717.600 244.050 718.050 ;
        RECT 283.950 717.600 286.050 718.050 ;
        RECT 236.400 716.400 286.050 717.600 ;
        RECT 142.950 715.950 145.050 716.400 ;
        RECT 148.950 715.950 151.050 716.400 ;
        RECT 241.950 715.950 244.050 716.400 ;
        RECT 283.950 715.950 286.050 716.400 ;
        RECT 373.950 717.600 376.050 718.050 ;
        RECT 403.950 717.600 406.050 718.050 ;
        RECT 427.950 717.600 430.050 718.050 ;
        RECT 442.950 717.600 445.050 718.050 ;
        RECT 373.950 716.400 445.050 717.600 ;
        RECT 373.950 715.950 376.050 716.400 ;
        RECT 403.950 715.950 406.050 716.400 ;
        RECT 427.950 715.950 430.050 716.400 ;
        RECT 442.950 715.950 445.050 716.400 ;
        RECT 487.950 717.600 490.050 718.050 ;
        RECT 517.800 717.600 519.900 718.050 ;
        RECT 487.950 716.400 519.900 717.600 ;
        RECT 487.950 715.950 490.050 716.400 ;
        RECT 517.800 715.950 519.900 716.400 ;
        RECT 520.950 717.600 523.050 718.050 ;
        RECT 538.950 717.600 541.050 718.050 ;
        RECT 520.950 716.400 541.050 717.600 ;
        RECT 520.950 715.950 523.050 716.400 ;
        RECT 538.950 715.950 541.050 716.400 ;
        RECT 601.950 717.600 604.050 718.050 ;
        RECT 619.950 717.600 622.050 718.050 ;
        RECT 649.950 717.600 652.050 718.050 ;
        RECT 601.950 716.400 652.050 717.600 ;
        RECT 601.950 715.950 604.050 716.400 ;
        RECT 619.950 715.950 622.050 716.400 ;
        RECT 649.950 715.950 652.050 716.400 ;
        RECT 727.950 717.600 730.050 718.050 ;
        RECT 745.950 717.600 748.050 718.050 ;
        RECT 727.950 716.400 748.050 717.600 ;
        RECT 727.950 715.950 730.050 716.400 ;
        RECT 745.950 715.950 748.050 716.400 ;
        RECT 43.950 714.600 46.050 715.050 ;
        RECT 55.950 714.600 58.050 715.050 ;
        RECT 43.950 713.400 58.050 714.600 ;
        RECT 43.950 712.950 46.050 713.400 ;
        RECT 55.950 712.950 58.050 713.400 ;
        RECT 73.950 714.600 76.050 715.050 ;
        RECT 98.400 714.600 99.600 715.800 ;
        RECT 73.950 713.400 99.600 714.600 ;
        RECT 112.950 714.600 115.050 715.050 ;
        RECT 121.950 714.600 124.050 715.050 ;
        RECT 112.950 713.400 124.050 714.600 ;
        RECT 73.950 712.950 76.050 713.400 ;
        RECT 112.950 712.950 115.050 713.400 ;
        RECT 121.950 712.950 124.050 713.400 ;
        RECT 223.950 714.600 226.050 715.050 ;
        RECT 238.950 714.600 241.050 715.050 ;
        RECT 292.950 714.600 295.050 715.050 ;
        RECT 223.950 713.400 295.050 714.600 ;
        RECT 223.950 712.950 226.050 713.400 ;
        RECT 238.950 712.950 241.050 713.400 ;
        RECT 292.950 712.950 295.050 713.400 ;
        RECT 310.950 714.600 313.050 715.050 ;
        RECT 355.800 714.600 357.900 715.050 ;
        RECT 310.950 713.400 357.900 714.600 ;
        RECT 310.950 712.950 313.050 713.400 ;
        RECT 355.800 712.950 357.900 713.400 ;
        RECT 358.950 714.600 361.050 715.050 ;
        RECT 370.950 714.600 373.050 715.050 ;
        RECT 358.950 713.400 373.050 714.600 ;
        RECT 358.950 712.950 361.050 713.400 ;
        RECT 370.950 712.950 373.050 713.400 ;
        RECT 382.950 714.600 385.050 715.050 ;
        RECT 397.950 714.600 400.050 715.050 ;
        RECT 454.950 714.600 457.050 715.050 ;
        RECT 382.950 713.400 457.050 714.600 ;
        RECT 518.400 714.600 519.600 715.950 ;
        RECT 541.950 714.600 544.050 715.050 ;
        RECT 518.400 713.400 544.050 714.600 ;
        RECT 382.950 712.950 385.050 713.400 ;
        RECT 397.950 712.950 400.050 713.400 ;
        RECT 454.950 712.950 457.050 713.400 ;
        RECT 541.950 712.950 544.050 713.400 ;
        RECT 559.950 714.600 562.050 715.050 ;
        RECT 652.950 714.600 655.050 715.050 ;
        RECT 679.950 714.600 682.050 715.050 ;
        RECT 559.950 713.400 567.600 714.600 ;
        RECT 559.950 712.950 562.050 713.400 ;
        RECT 145.950 711.600 148.050 712.050 ;
        RECT 235.950 711.600 238.050 712.050 ;
        RECT 145.950 710.400 238.050 711.600 ;
        RECT 145.950 709.950 148.050 710.400 ;
        RECT 235.950 709.950 238.050 710.400 ;
        RECT 292.950 711.600 295.050 711.900 ;
        RECT 376.950 711.600 379.050 712.050 ;
        RECT 292.950 710.400 379.050 711.600 ;
        RECT 292.950 709.800 295.050 710.400 ;
        RECT 376.950 709.950 379.050 710.400 ;
        RECT 400.950 711.600 403.050 712.050 ;
        RECT 451.950 711.600 454.050 712.050 ;
        RECT 400.950 710.400 454.050 711.600 ;
        RECT 400.950 709.950 403.050 710.400 ;
        RECT 451.950 709.950 454.050 710.400 ;
        RECT 502.950 711.600 505.050 712.050 ;
        RECT 566.400 711.600 567.600 713.400 ;
        RECT 652.950 713.400 682.050 714.600 ;
        RECT 652.950 712.950 655.050 713.400 ;
        RECT 679.950 712.950 682.050 713.400 ;
        RECT 586.950 711.600 589.050 712.050 ;
        RECT 502.950 710.400 564.600 711.600 ;
        RECT 566.400 710.400 589.050 711.600 ;
        RECT 502.950 709.950 505.050 710.400 ;
        RECT 19.950 708.600 22.050 709.050 ;
        RECT 34.950 708.600 37.050 709.050 ;
        RECT 130.950 708.600 133.050 709.050 ;
        RECT 19.950 707.400 133.050 708.600 ;
        RECT 19.950 706.950 22.050 707.400 ;
        RECT 34.950 706.950 37.050 707.400 ;
        RECT 130.950 706.950 133.050 707.400 ;
        RECT 139.950 708.600 142.050 709.050 ;
        RECT 154.950 708.600 157.050 709.050 ;
        RECT 250.950 708.600 253.050 709.050 ;
        RECT 139.950 707.400 253.050 708.600 ;
        RECT 139.950 706.950 142.050 707.400 ;
        RECT 154.950 706.950 157.050 707.400 ;
        RECT 250.950 706.950 253.050 707.400 ;
        RECT 259.950 708.600 262.050 709.050 ;
        RECT 280.950 708.600 283.050 709.050 ;
        RECT 304.950 708.600 307.050 709.050 ;
        RECT 331.950 708.600 334.050 709.050 ;
        RECT 259.950 707.400 334.050 708.600 ;
        RECT 259.950 706.950 262.050 707.400 ;
        RECT 280.950 706.950 283.050 707.400 ;
        RECT 304.950 706.950 307.050 707.400 ;
        RECT 331.950 706.950 334.050 707.400 ;
        RECT 367.950 708.600 370.050 709.050 ;
        RECT 397.950 708.600 400.050 709.050 ;
        RECT 367.950 707.400 400.050 708.600 ;
        RECT 367.950 706.950 370.050 707.400 ;
        RECT 397.950 706.950 400.050 707.400 ;
        RECT 460.950 708.600 463.050 709.050 ;
        RECT 538.950 708.600 541.050 709.050 ;
        RECT 553.950 708.600 556.050 709.050 ;
        RECT 460.950 707.400 537.600 708.600 ;
        RECT 460.950 706.950 463.050 707.400 ;
        RECT 37.950 705.600 40.050 706.050 ;
        RECT 112.950 705.600 115.050 706.050 ;
        RECT 37.950 704.400 115.050 705.600 ;
        RECT 37.950 703.950 40.050 704.400 ;
        RECT 112.950 703.950 115.050 704.400 ;
        RECT 190.950 705.600 193.050 706.050 ;
        RECT 256.950 705.600 259.050 706.050 ;
        RECT 190.950 704.400 259.050 705.600 ;
        RECT 190.950 703.950 193.050 704.400 ;
        RECT 256.950 703.950 259.050 704.400 ;
        RECT 283.950 705.600 286.050 706.050 ;
        RECT 361.950 705.600 364.050 706.050 ;
        RECT 283.950 704.400 364.050 705.600 ;
        RECT 283.950 703.950 286.050 704.400 ;
        RECT 361.950 703.950 364.050 704.400 ;
        RECT 379.950 705.600 382.050 706.050 ;
        RECT 400.950 705.600 403.050 706.050 ;
        RECT 379.950 704.400 403.050 705.600 ;
        RECT 379.950 703.950 382.050 704.400 ;
        RECT 400.950 703.950 403.050 704.400 ;
        RECT 409.950 705.600 412.050 706.050 ;
        RECT 433.950 705.600 436.050 706.050 ;
        RECT 409.950 704.400 436.050 705.600 ;
        RECT 536.400 705.600 537.600 707.400 ;
        RECT 538.950 707.400 556.050 708.600 ;
        RECT 563.400 708.600 564.600 710.400 ;
        RECT 586.950 709.950 589.050 710.400 ;
        RECT 688.950 711.600 691.050 712.050 ;
        RECT 712.950 711.600 715.050 712.050 ;
        RECT 688.950 710.400 715.050 711.600 ;
        RECT 688.950 709.950 691.050 710.400 ;
        RECT 712.950 709.950 715.050 710.400 ;
        RECT 757.950 711.600 760.050 712.050 ;
        RECT 850.950 711.600 853.050 712.050 ;
        RECT 757.950 710.400 853.050 711.600 ;
        RECT 757.950 709.950 760.050 710.400 ;
        RECT 850.950 709.950 853.050 710.400 ;
        RECT 589.950 708.600 592.050 709.050 ;
        RECT 658.950 708.600 661.050 709.050 ;
        RECT 563.400 707.400 592.050 708.600 ;
        RECT 538.950 706.950 541.050 707.400 ;
        RECT 553.950 706.950 556.050 707.400 ;
        RECT 589.950 706.950 592.050 707.400 ;
        RECT 629.400 707.400 661.050 708.600 ;
        RECT 547.950 705.600 550.050 706.050 ;
        RECT 536.400 704.400 550.050 705.600 ;
        RECT 409.950 703.950 412.050 704.400 ;
        RECT 433.950 703.950 436.050 704.400 ;
        RECT 547.950 703.950 550.050 704.400 ;
        RECT 553.950 705.600 556.050 705.900 ;
        RECT 629.400 705.600 630.600 707.400 ;
        RECT 658.950 706.950 661.050 707.400 ;
        RECT 664.950 708.600 667.050 709.050 ;
        RECT 694.950 708.600 697.050 709.050 ;
        RECT 664.950 707.400 697.050 708.600 ;
        RECT 664.950 706.950 667.050 707.400 ;
        RECT 694.950 706.950 697.050 707.400 ;
        RECT 799.950 708.600 802.050 709.050 ;
        RECT 826.950 708.600 829.050 709.050 ;
        RECT 799.950 707.400 829.050 708.600 ;
        RECT 799.950 706.950 802.050 707.400 ;
        RECT 826.950 706.950 829.050 707.400 ;
        RECT 553.950 704.400 630.600 705.600 ;
        RECT 631.950 705.600 634.050 706.050 ;
        RECT 703.950 705.600 706.050 706.050 ;
        RECT 751.950 705.600 754.050 706.050 ;
        RECT 772.950 705.600 775.050 706.050 ;
        RECT 631.950 704.400 775.050 705.600 ;
        RECT 553.950 703.800 556.050 704.400 ;
        RECT 631.950 703.950 634.050 704.400 ;
        RECT 703.950 703.950 706.050 704.400 ;
        RECT 751.950 703.950 754.050 704.400 ;
        RECT 772.950 703.950 775.050 704.400 ;
        RECT 799.950 705.600 802.050 705.900 ;
        RECT 808.950 705.600 811.050 706.050 ;
        RECT 799.950 704.400 811.050 705.600 ;
        RECT 799.950 703.800 802.050 704.400 ;
        RECT 808.950 703.950 811.050 704.400 ;
        RECT 118.950 702.600 121.050 703.050 ;
        RECT 166.950 702.600 169.050 703.050 ;
        RECT 118.950 701.400 169.050 702.600 ;
        RECT 118.950 700.950 121.050 701.400 ;
        RECT 166.950 700.950 169.050 701.400 ;
        RECT 277.950 702.600 280.050 703.050 ;
        RECT 364.950 702.600 367.050 703.050 ;
        RECT 277.950 701.400 367.050 702.600 ;
        RECT 277.950 700.950 280.050 701.400 ;
        RECT 364.950 700.950 367.050 701.400 ;
        RECT 370.950 702.600 373.050 703.050 ;
        RECT 463.950 702.600 466.050 703.050 ;
        RECT 370.950 701.400 466.050 702.600 ;
        RECT 370.950 700.950 373.050 701.400 ;
        RECT 463.950 700.950 466.050 701.400 ;
        RECT 499.950 702.600 502.050 703.050 ;
        RECT 511.950 702.600 514.050 703.050 ;
        RECT 583.950 702.600 586.050 703.050 ;
        RECT 499.950 701.400 586.050 702.600 ;
        RECT 499.950 700.950 502.050 701.400 ;
        RECT 511.950 700.950 514.050 701.400 ;
        RECT 583.950 700.950 586.050 701.400 ;
        RECT 634.950 702.600 637.050 703.050 ;
        RECT 652.950 702.600 655.050 703.050 ;
        RECT 634.950 701.400 655.050 702.600 ;
        RECT 634.950 700.950 637.050 701.400 ;
        RECT 652.950 700.950 655.050 701.400 ;
        RECT 658.950 702.600 661.050 703.050 ;
        RECT 832.950 702.600 835.050 703.050 ;
        RECT 658.950 701.400 835.050 702.600 ;
        RECT 658.950 700.950 661.050 701.400 ;
        RECT 832.950 700.950 835.050 701.400 ;
        RECT 34.950 699.600 37.050 700.050 ;
        RECT 58.950 699.600 61.050 700.050 ;
        RECT 67.950 699.600 70.050 700.050 ;
        RECT 88.950 699.600 91.050 700.050 ;
        RECT 34.950 698.400 91.050 699.600 ;
        RECT 34.950 697.950 37.050 698.400 ;
        RECT 58.950 697.950 61.050 698.400 ;
        RECT 67.950 697.950 70.050 698.400 ;
        RECT 88.950 697.950 91.050 698.400 ;
        RECT 109.950 699.600 112.050 700.050 ;
        RECT 196.950 699.600 199.050 700.050 ;
        RECT 217.950 699.600 220.050 700.050 ;
        RECT 226.950 699.600 229.050 700.050 ;
        RECT 109.950 698.400 229.050 699.600 ;
        RECT 109.950 697.950 112.050 698.400 ;
        RECT 196.950 697.950 199.050 698.400 ;
        RECT 217.950 697.950 220.050 698.400 ;
        RECT 226.950 697.950 229.050 698.400 ;
        RECT 235.950 699.600 238.050 700.050 ;
        RECT 256.950 699.600 259.050 700.050 ;
        RECT 235.950 698.400 259.050 699.600 ;
        RECT 235.950 697.950 238.050 698.400 ;
        RECT 256.950 697.950 259.050 698.400 ;
        RECT 310.950 699.600 313.050 700.050 ;
        RECT 358.950 699.600 361.050 700.050 ;
        RECT 310.950 698.400 361.050 699.600 ;
        RECT 310.950 697.950 313.050 698.400 ;
        RECT 358.950 697.950 361.050 698.400 ;
        RECT 376.950 699.600 379.050 700.050 ;
        RECT 460.950 699.600 463.050 700.050 ;
        RECT 376.950 698.400 463.050 699.600 ;
        RECT 376.950 697.950 379.050 698.400 ;
        RECT 460.950 697.950 463.050 698.400 ;
        RECT 466.950 699.600 469.050 700.050 ;
        RECT 532.950 699.600 535.050 700.050 ;
        RECT 466.950 698.400 535.050 699.600 ;
        RECT 466.950 697.950 469.050 698.400 ;
        RECT 532.950 697.950 535.050 698.400 ;
        RECT 538.950 699.600 541.050 700.050 ;
        RECT 793.950 699.600 796.050 700.050 ;
        RECT 811.950 699.600 814.050 700.050 ;
        RECT 538.950 698.400 814.050 699.600 ;
        RECT 538.950 697.950 541.050 698.400 ;
        RECT 793.950 697.950 796.050 698.400 ;
        RECT 811.950 697.950 814.050 698.400 ;
        RECT 112.950 696.600 115.050 697.050 ;
        RECT 124.950 696.600 127.050 697.050 ;
        RECT 337.950 696.600 340.050 697.050 ;
        RECT 112.950 695.400 127.050 696.600 ;
        RECT 112.950 694.950 115.050 695.400 ;
        RECT 124.950 694.950 127.050 695.400 ;
        RECT 314.400 695.400 340.050 696.600 ;
        RECT 314.400 694.050 315.600 695.400 ;
        RECT 337.950 694.950 340.050 695.400 ;
        RECT 346.950 696.600 349.050 697.050 ;
        RECT 457.950 696.600 460.050 697.050 ;
        RECT 346.950 695.400 460.050 696.600 ;
        RECT 346.950 694.950 349.050 695.400 ;
        RECT 457.950 694.950 460.050 695.400 ;
        RECT 463.950 696.600 466.050 697.050 ;
        RECT 505.950 696.600 508.050 697.050 ;
        RECT 514.950 696.600 517.050 697.050 ;
        RECT 463.950 695.400 495.600 696.600 ;
        RECT 463.950 694.950 466.050 695.400 ;
        RECT 4.950 693.600 7.050 694.050 ;
        RECT 28.950 693.600 31.050 694.050 ;
        RECT 37.950 693.600 40.050 694.050 ;
        RECT 4.950 692.400 40.050 693.600 ;
        RECT 4.950 691.950 7.050 692.400 ;
        RECT 28.950 691.950 31.050 692.400 ;
        RECT 37.950 691.950 40.050 692.400 ;
        RECT 67.950 693.600 70.050 694.050 ;
        RECT 85.950 693.600 88.050 694.050 ;
        RECT 67.950 692.400 88.050 693.600 ;
        RECT 67.950 691.950 70.050 692.400 ;
        RECT 85.950 691.950 88.050 692.400 ;
        RECT 178.950 693.600 181.050 694.050 ;
        RECT 196.950 693.600 199.050 694.050 ;
        RECT 178.950 692.400 199.050 693.600 ;
        RECT 178.950 691.950 181.050 692.400 ;
        RECT 196.950 691.950 199.050 692.400 ;
        RECT 250.950 693.600 253.050 694.050 ;
        RECT 277.950 693.600 280.050 694.050 ;
        RECT 250.950 692.400 280.050 693.600 ;
        RECT 250.950 691.950 253.050 692.400 ;
        RECT 277.950 691.950 280.050 692.400 ;
        RECT 286.950 693.600 289.050 694.050 ;
        RECT 313.950 693.600 316.050 694.050 ;
        RECT 286.950 692.400 316.050 693.600 ;
        RECT 286.950 691.950 289.050 692.400 ;
        RECT 313.950 691.950 316.050 692.400 ;
        RECT 340.950 693.600 343.050 694.050 ;
        RECT 394.950 693.600 397.050 694.050 ;
        RECT 409.950 693.600 412.050 694.050 ;
        RECT 340.950 692.400 412.050 693.600 ;
        RECT 340.950 691.950 343.050 692.400 ;
        RECT 394.950 691.950 397.050 692.400 ;
        RECT 409.950 691.950 412.050 692.400 ;
        RECT 418.950 693.600 421.050 694.050 ;
        RECT 490.950 693.600 493.050 694.050 ;
        RECT 418.950 692.400 493.050 693.600 ;
        RECT 494.400 693.600 495.600 695.400 ;
        RECT 505.950 695.400 517.050 696.600 ;
        RECT 505.950 694.950 508.050 695.400 ;
        RECT 514.950 694.950 517.050 695.400 ;
        RECT 544.950 696.600 547.050 697.050 ;
        RECT 562.950 696.600 565.050 697.050 ;
        RECT 544.950 695.400 565.050 696.600 ;
        RECT 544.950 694.950 547.050 695.400 ;
        RECT 562.950 694.950 565.050 695.400 ;
        RECT 577.950 696.600 580.050 697.050 ;
        RECT 610.950 696.600 613.050 697.050 ;
        RECT 721.800 696.600 723.900 697.050 ;
        RECT 577.950 695.400 613.050 696.600 ;
        RECT 680.400 696.000 723.900 696.600 ;
        RECT 577.950 694.950 580.050 695.400 ;
        RECT 610.950 694.950 613.050 695.400 ;
        RECT 679.950 695.400 723.900 696.000 ;
        RECT 520.950 693.600 523.050 694.050 ;
        RECT 494.400 692.400 523.050 693.600 ;
        RECT 418.950 691.950 421.050 692.400 ;
        RECT 490.950 691.950 493.050 692.400 ;
        RECT 520.950 691.950 523.050 692.400 ;
        RECT 679.950 691.950 682.050 695.400 ;
        RECT 721.800 694.950 723.900 695.400 ;
        RECT 724.950 696.600 727.050 697.050 ;
        RECT 769.950 696.600 772.050 697.050 ;
        RECT 724.950 695.400 772.050 696.600 ;
        RECT 724.950 694.950 727.050 695.400 ;
        RECT 769.950 694.950 772.050 695.400 ;
        RECT 40.950 690.600 43.050 691.050 ;
        RECT 91.950 690.600 94.050 691.050 ;
        RECT 40.950 689.400 94.050 690.600 ;
        RECT 40.950 688.950 43.050 689.400 ;
        RECT 91.950 688.950 94.050 689.400 ;
        RECT 100.950 690.600 103.050 691.050 ;
        RECT 106.800 690.600 108.900 691.050 ;
        RECT 100.950 689.400 108.900 690.600 ;
        RECT 100.950 688.950 103.050 689.400 ;
        RECT 106.800 688.950 108.900 689.400 ;
        RECT 109.950 690.600 112.050 691.050 ;
        RECT 166.950 690.600 169.050 691.050 ;
        RECT 247.950 690.600 250.050 691.050 ;
        RECT 109.950 689.400 250.050 690.600 ;
        RECT 109.950 688.950 112.050 689.400 ;
        RECT 166.950 688.950 169.050 689.400 ;
        RECT 247.950 688.950 250.050 689.400 ;
        RECT 256.950 690.600 259.050 691.050 ;
        RECT 292.950 690.600 295.050 691.050 ;
        RECT 256.950 689.400 295.050 690.600 ;
        RECT 256.950 688.950 259.050 689.400 ;
        RECT 292.950 688.950 295.050 689.400 ;
        RECT 319.950 690.600 322.050 691.050 ;
        RECT 361.950 690.600 364.050 691.050 ;
        RECT 319.950 689.400 364.050 690.600 ;
        RECT 319.950 688.950 322.050 689.400 ;
        RECT 361.950 688.950 364.050 689.400 ;
        RECT 367.950 690.600 370.050 691.050 ;
        RECT 376.950 690.600 379.050 691.050 ;
        RECT 367.950 689.400 379.050 690.600 ;
        RECT 367.950 688.950 370.050 689.400 ;
        RECT 376.950 688.950 379.050 689.400 ;
        RECT 430.950 690.600 433.050 691.050 ;
        RECT 445.950 690.600 448.050 691.050 ;
        RECT 469.950 690.600 472.050 691.050 ;
        RECT 430.950 689.400 472.050 690.600 ;
        RECT 430.950 688.950 433.050 689.400 ;
        RECT 445.950 688.950 448.050 689.400 ;
        RECT 469.950 688.950 472.050 689.400 ;
        RECT 496.950 690.600 499.050 691.050 ;
        RECT 538.950 690.600 541.050 691.050 ;
        RECT 496.950 689.400 541.050 690.600 ;
        RECT 496.950 688.950 499.050 689.400 ;
        RECT 538.950 688.950 541.050 689.400 ;
        RECT 547.950 690.600 550.050 691.050 ;
        RECT 559.950 690.600 562.050 691.050 ;
        RECT 547.950 689.400 562.050 690.600 ;
        RECT 547.950 688.950 550.050 689.400 ;
        RECT 559.950 688.950 562.050 689.400 ;
        RECT 715.950 690.600 718.050 691.050 ;
        RECT 742.950 690.600 745.050 691.050 ;
        RECT 715.950 689.400 745.050 690.600 ;
        RECT 715.950 688.950 718.050 689.400 ;
        RECT 742.950 688.950 745.050 689.400 ;
        RECT 52.950 687.600 55.050 688.050 ;
        RECT 130.950 687.600 133.050 688.050 ;
        RECT 136.950 687.600 139.050 688.050 ;
        RECT 52.950 686.400 63.600 687.600 ;
        RECT 52.950 685.950 55.050 686.400 ;
        RECT 10.950 684.600 13.050 685.200 ;
        RECT 19.950 684.600 22.050 685.050 ;
        RECT 10.950 683.400 22.050 684.600 ;
        RECT 10.950 683.100 13.050 683.400 ;
        RECT 19.950 682.950 22.050 683.400 ;
        RECT 31.950 682.950 34.050 685.050 ;
        RECT 49.950 683.100 52.050 685.200 ;
        RECT 4.950 678.450 7.050 678.900 ;
        RECT 13.950 678.450 16.050 678.900 ;
        RECT 32.400 678.750 33.600 682.950 ;
        RECT 50.400 681.600 51.600 683.100 ;
        RECT 50.400 681.000 57.600 681.600 ;
        RECT 50.400 680.400 58.050 681.000 ;
        RECT 4.950 677.250 16.050 678.450 ;
        RECT 4.950 676.800 7.050 677.250 ;
        RECT 13.950 676.800 16.050 677.250 ;
        RECT 31.950 676.650 34.050 678.750 ;
        RECT 37.950 678.600 40.050 678.750 ;
        RECT 46.950 678.600 49.050 678.900 ;
        RECT 37.950 677.400 49.050 678.600 ;
        RECT 37.950 676.650 40.050 677.400 ;
        RECT 46.950 676.800 49.050 677.400 ;
        RECT 55.950 676.950 58.050 680.400 ;
        RECT 62.400 679.050 63.600 686.400 ;
        RECT 130.950 686.400 139.050 687.600 ;
        RECT 130.950 685.950 133.050 686.400 ;
        RECT 136.950 685.950 139.050 686.400 ;
        RECT 181.950 687.600 184.050 688.050 ;
        RECT 187.950 687.600 190.050 688.050 ;
        RECT 268.950 687.600 271.050 688.050 ;
        RECT 181.950 686.400 190.050 687.600 ;
        RECT 181.950 685.950 184.050 686.400 ;
        RECT 187.950 685.950 190.050 686.400 ;
        RECT 257.400 686.400 271.050 687.600 ;
        RECT 73.950 684.600 76.050 685.050 ;
        RECT 79.950 684.600 82.050 685.050 ;
        RECT 73.950 683.400 82.050 684.600 ;
        RECT 73.950 682.950 76.050 683.400 ;
        RECT 79.950 682.950 82.050 683.400 ;
        RECT 100.800 682.950 102.900 685.050 ;
        RECT 61.950 678.600 64.050 679.050 ;
        RECT 82.950 678.600 85.050 678.750 ;
        RECT 61.950 677.400 85.050 678.600 ;
        RECT 61.950 676.950 64.050 677.400 ;
        RECT 82.950 676.650 85.050 677.400 ;
        RECT 88.950 678.300 91.050 678.750 ;
        RECT 94.950 678.300 97.050 678.750 ;
        RECT 88.950 677.100 97.050 678.300 ;
        RECT 101.400 678.600 102.600 682.950 ;
        RECT 103.950 681.600 106.050 684.900 ;
        RECT 109.950 684.600 112.050 685.050 ;
        RECT 127.950 684.600 130.050 685.050 ;
        RECT 145.800 684.600 147.900 685.200 ;
        RECT 109.950 683.400 130.050 684.600 ;
        RECT 109.950 682.950 112.050 683.400 ;
        RECT 127.950 682.950 130.050 683.400 ;
        RECT 131.400 683.400 147.900 684.600 ;
        RECT 131.400 681.600 132.600 683.400 ;
        RECT 145.800 683.100 147.900 683.400 ;
        RECT 148.950 682.950 151.050 685.050 ;
        RECT 168.000 684.600 172.050 685.050 ;
        RECT 167.400 682.950 172.050 684.600 ;
        RECT 103.950 681.000 132.600 681.600 ;
        RECT 104.400 680.400 132.600 681.000 ;
        RECT 115.950 678.600 118.050 679.050 ;
        RECT 122.400 678.750 123.600 680.400 ;
        RECT 149.400 679.050 150.600 682.950 ;
        RECT 167.400 681.600 168.600 682.950 ;
        RECT 184.950 681.600 187.050 685.050 ;
        RECT 211.950 683.100 214.050 685.200 ;
        RECT 232.950 684.600 235.050 685.200 ;
        RECT 253.950 684.600 256.050 685.200 ;
        RECT 232.950 683.400 256.050 684.600 ;
        RECT 232.950 683.100 235.050 683.400 ;
        RECT 253.950 683.100 256.050 683.400 ;
        RECT 164.400 680.400 168.600 681.600 ;
        RECT 170.400 681.000 187.050 681.600 ;
        RECT 170.400 680.400 186.600 681.000 ;
        RECT 101.400 677.400 118.050 678.600 ;
        RECT 88.950 676.650 91.050 677.100 ;
        RECT 94.950 676.650 97.050 677.100 ;
        RECT 115.950 676.950 118.050 677.400 ;
        RECT 121.950 676.650 124.050 678.750 ;
        RECT 148.950 676.950 151.050 679.050 ;
        RECT 164.400 676.050 165.600 680.400 ;
        RECT 170.400 678.750 171.600 680.400 ;
        RECT 169.950 676.650 172.050 678.750 ;
        RECT 190.950 678.600 193.050 678.750 ;
        RECT 212.400 678.600 213.600 683.100 ;
        RECT 190.950 678.000 213.600 678.600 ;
        RECT 214.950 678.600 217.050 679.050 ;
        RECT 257.400 678.900 258.600 686.400 ;
        RECT 268.950 685.950 271.050 686.400 ;
        RECT 328.950 687.600 331.050 688.050 ;
        RECT 343.950 687.600 346.050 688.050 ;
        RECT 352.950 687.600 355.050 688.050 ;
        RECT 328.950 686.400 355.050 687.600 ;
        RECT 328.950 685.950 331.050 686.400 ;
        RECT 343.950 685.950 346.050 686.400 ;
        RECT 352.950 685.950 355.050 686.400 ;
        RECT 364.950 687.600 367.050 688.050 ;
        RECT 379.950 687.600 382.050 688.050 ;
        RECT 364.950 686.400 382.050 687.600 ;
        RECT 364.950 685.950 367.050 686.400 ;
        RECT 379.950 685.950 382.050 686.400 ;
        RECT 412.950 687.600 415.050 688.050 ;
        RECT 418.950 687.600 421.050 688.050 ;
        RECT 412.950 686.400 421.050 687.600 ;
        RECT 412.950 685.950 415.050 686.400 ;
        RECT 418.950 685.950 421.050 686.400 ;
        RECT 436.950 687.600 439.050 688.050 ;
        RECT 448.950 687.600 451.050 688.050 ;
        RECT 436.950 686.400 451.050 687.600 ;
        RECT 436.950 685.950 439.050 686.400 ;
        RECT 448.950 685.950 451.050 686.400 ;
        RECT 454.950 687.600 457.050 688.050 ;
        RECT 466.950 687.600 469.050 688.050 ;
        RECT 454.950 686.400 469.050 687.600 ;
        RECT 454.950 685.950 457.050 686.400 ;
        RECT 466.950 685.950 469.050 686.400 ;
        RECT 532.800 687.000 534.900 688.050 ;
        RECT 537.000 687.900 540.000 688.050 ;
        RECT 537.000 687.600 541.050 687.900 ;
        RECT 532.800 685.950 535.050 687.000 ;
        RECT 271.950 684.600 274.050 685.200 ;
        RECT 277.950 684.600 280.050 685.050 ;
        RECT 271.950 683.400 280.050 684.600 ;
        RECT 271.950 683.100 274.050 683.400 ;
        RECT 277.950 682.950 280.050 683.400 ;
        RECT 289.800 682.950 291.900 685.050 ;
        RECT 292.950 684.600 295.050 685.050 ;
        RECT 298.950 684.600 301.050 685.050 ;
        RECT 292.950 683.400 301.050 684.600 ;
        RECT 292.950 682.950 295.050 683.400 ;
        RECT 298.950 682.950 301.050 683.400 ;
        RECT 310.950 682.950 313.050 685.050 ;
        RECT 319.800 684.000 321.900 685.050 ;
        RECT 319.800 682.950 322.050 684.000 ;
        RECT 322.950 682.950 325.050 685.050 ;
        RECT 229.950 678.600 232.050 678.900 ;
        RECT 190.950 677.400 214.050 678.000 ;
        RECT 190.950 676.650 193.050 677.400 ;
        RECT 67.950 675.600 70.050 676.050 ;
        RECT 73.950 675.600 76.050 676.050 ;
        RECT 67.950 674.400 76.050 675.600 ;
        RECT 164.400 674.400 169.050 676.050 ;
        RECT 67.950 673.950 70.050 674.400 ;
        RECT 73.950 673.950 76.050 674.400 ;
        RECT 165.000 673.950 169.050 674.400 ;
        RECT 211.950 673.950 214.050 677.400 ;
        RECT 214.950 677.400 232.050 678.600 ;
        RECT 214.950 676.950 217.050 677.400 ;
        RECT 229.950 676.800 232.050 677.400 ;
        RECT 256.950 676.800 259.050 678.900 ;
        RECT 290.400 678.750 291.600 682.950 ;
        RECT 311.400 679.050 312.600 682.950 ;
        RECT 319.950 681.600 322.050 682.950 ;
        RECT 314.400 681.000 322.050 681.600 ;
        RECT 314.400 680.400 321.450 681.000 ;
        RECT 289.950 676.650 292.050 678.750 ;
        RECT 310.950 676.950 313.050 679.050 ;
        RECT 235.950 675.600 238.050 676.050 ;
        RECT 256.950 675.600 259.050 676.050 ;
        RECT 235.950 674.400 259.050 675.600 ;
        RECT 235.950 673.950 238.050 674.400 ;
        RECT 256.950 673.950 259.050 674.400 ;
        RECT 295.950 675.600 298.050 676.050 ;
        RECT 314.400 675.600 315.600 680.400 ;
        RECT 316.950 678.600 319.050 679.050 ;
        RECT 323.400 678.600 324.600 682.950 ;
        RECT 346.950 681.600 349.050 685.050 ;
        RECT 355.950 684.600 358.050 685.050 ;
        RECT 373.950 684.600 376.050 685.050 ;
        RECT 355.950 683.400 376.050 684.600 ;
        RECT 355.950 682.950 358.050 683.400 ;
        RECT 373.950 682.950 376.050 683.400 ;
        RECT 397.950 684.600 402.000 685.050 ;
        RECT 409.950 684.600 412.050 685.050 ;
        RECT 421.950 684.600 424.050 685.050 ;
        RECT 397.950 682.950 402.600 684.600 ;
        RECT 409.950 683.400 424.050 684.600 ;
        RECT 409.950 682.950 412.050 683.400 ;
        RECT 421.950 682.950 424.050 683.400 ;
        RECT 433.950 682.950 436.050 685.050 ;
        RECT 469.950 684.600 472.050 685.200 ;
        RECT 475.950 684.750 478.050 685.050 ;
        RECT 484.950 684.750 487.050 685.200 ;
        RECT 469.950 683.400 474.600 684.600 ;
        RECT 469.950 683.100 472.050 683.400 ;
        RECT 338.400 681.000 349.050 681.600 ;
        RECT 401.400 681.600 402.600 682.950 ;
        RECT 338.400 680.400 348.600 681.000 ;
        RECT 401.400 680.400 408.600 681.600 ;
        RECT 316.950 677.400 324.600 678.600 ;
        RECT 331.950 678.600 334.050 678.750 ;
        RECT 338.400 678.600 339.600 680.400 ;
        RECT 331.950 677.400 339.600 678.600 ;
        RECT 340.950 678.600 343.050 679.050 ;
        RECT 349.950 678.600 352.050 678.750 ;
        RECT 340.950 677.400 352.050 678.600 ;
        RECT 407.400 678.600 408.600 680.400 ;
        RECT 424.950 678.600 427.050 679.050 ;
        RECT 434.400 678.750 435.600 682.950 ;
        RECT 473.400 682.050 474.600 683.400 ;
        RECT 475.950 683.550 487.050 684.750 ;
        RECT 475.950 682.950 478.050 683.550 ;
        RECT 484.950 683.100 487.050 683.550 ;
        RECT 517.950 682.950 520.050 685.050 ;
        RECT 523.950 684.600 526.050 684.900 ;
        RECT 532.950 684.600 535.050 685.950 ;
        RECT 523.950 684.000 535.050 684.600 ;
        RECT 536.400 685.950 541.050 687.600 ;
        RECT 565.950 687.600 568.050 688.050 ;
        RECT 571.950 687.600 574.050 688.050 ;
        RECT 622.950 687.600 625.050 688.050 ;
        RECT 718.950 687.600 721.050 688.050 ;
        RECT 736.950 687.600 739.050 688.050 ;
        RECT 565.950 686.400 597.600 687.600 ;
        RECT 565.950 685.950 568.050 686.400 ;
        RECT 571.950 685.950 574.050 686.400 ;
        RECT 523.950 683.400 534.450 684.000 ;
        RECT 473.400 681.900 477.000 682.050 ;
        RECT 473.400 680.400 478.050 681.900 ;
        RECT 474.000 679.950 478.050 680.400 ;
        RECT 475.950 679.800 478.050 679.950 ;
        RECT 407.400 677.400 427.050 678.600 ;
        RECT 316.950 676.950 319.050 677.400 ;
        RECT 331.950 676.650 334.050 677.400 ;
        RECT 340.950 676.950 343.050 677.400 ;
        RECT 349.950 676.650 352.050 677.400 ;
        RECT 424.950 676.950 427.050 677.400 ;
        RECT 433.950 678.600 436.050 678.750 ;
        RECT 448.950 678.600 451.050 678.750 ;
        RECT 433.950 677.400 451.050 678.600 ;
        RECT 433.950 676.650 436.050 677.400 ;
        RECT 448.950 676.650 451.050 677.400 ;
        RECT 460.950 678.600 463.050 679.050 ;
        RECT 472.950 678.600 475.050 679.050 ;
        RECT 460.950 677.400 475.050 678.600 ;
        RECT 460.950 676.950 463.050 677.400 ;
        RECT 472.950 676.950 475.050 677.400 ;
        RECT 487.950 678.600 490.050 678.900 ;
        RECT 496.950 678.600 499.050 679.050 ;
        RECT 487.950 677.400 499.050 678.600 ;
        RECT 518.400 678.600 519.600 682.950 ;
        RECT 523.950 682.800 526.050 683.400 ;
        RECT 520.950 678.600 523.050 678.750 ;
        RECT 518.400 677.400 523.050 678.600 ;
        RECT 487.950 676.800 490.050 677.400 ;
        RECT 496.950 676.950 499.050 677.400 ;
        RECT 520.950 676.650 523.050 677.400 ;
        RECT 524.400 676.050 525.600 682.800 ;
        RECT 536.400 679.050 537.600 685.950 ;
        RECT 538.950 685.800 541.050 685.950 ;
        RECT 596.400 685.050 597.600 686.400 ;
        RECT 622.950 686.400 669.600 687.600 ;
        RECT 622.950 685.950 625.050 686.400 ;
        RECT 562.950 681.600 565.050 685.050 ;
        RECT 595.950 684.600 600.000 685.050 ;
        RECT 604.950 684.600 607.050 685.050 ;
        RECT 613.950 684.600 616.050 685.050 ;
        RECT 652.950 684.600 655.050 685.200 ;
        RECT 595.950 682.950 600.600 684.600 ;
        RECT 604.950 683.400 616.050 684.600 ;
        RECT 604.950 682.950 607.050 683.400 ;
        RECT 613.950 682.950 616.050 683.400 ;
        RECT 632.400 683.400 655.050 684.600 ;
        RECT 557.400 681.000 565.050 681.600 ;
        RECT 557.400 680.400 564.600 681.000 ;
        RECT 535.950 676.950 538.050 679.050 ;
        RECT 541.950 678.600 544.050 678.750 ;
        RECT 550.950 678.600 553.050 679.050 ;
        RECT 557.400 678.900 558.600 680.400 ;
        RECT 599.400 679.050 600.600 682.950 ;
        RECT 541.950 677.400 553.050 678.600 ;
        RECT 541.950 676.650 544.050 677.400 ;
        RECT 550.950 676.950 553.050 677.400 ;
        RECT 556.950 676.800 559.050 678.900 ;
        RECT 565.950 678.300 568.050 678.750 ;
        RECT 574.950 678.300 577.050 678.750 ;
        RECT 565.950 677.100 577.050 678.300 ;
        RECT 565.950 676.650 568.050 677.100 ;
        RECT 574.950 676.650 577.050 677.100 ;
        RECT 598.950 676.950 601.050 679.050 ;
        RECT 604.950 678.600 607.050 679.050 ;
        RECT 632.400 678.600 633.600 683.400 ;
        RECT 652.950 683.100 655.050 683.400 ;
        RECT 658.950 683.100 661.050 685.200 ;
        RECT 668.400 685.050 669.600 686.400 ;
        RECT 698.400 686.400 739.050 687.600 ;
        RECT 698.400 685.050 699.600 686.400 ;
        RECT 718.950 685.950 721.050 686.400 ;
        RECT 736.950 685.950 739.050 686.400 ;
        RECT 668.400 683.400 673.050 685.050 ;
        RECT 604.950 677.400 633.600 678.600 ;
        RECT 604.950 676.950 607.050 677.400 ;
        RECT 295.950 674.400 315.600 675.600 ;
        RECT 364.950 675.600 367.050 676.050 ;
        RECT 385.950 675.600 388.050 676.050 ;
        RECT 364.950 674.400 388.050 675.600 ;
        RECT 295.950 673.950 298.050 674.400 ;
        RECT 364.950 673.950 367.050 674.400 ;
        RECT 385.950 673.950 388.050 674.400 ;
        RECT 475.950 675.600 478.050 676.050 ;
        RECT 481.950 675.600 484.050 676.050 ;
        RECT 522.000 675.600 525.600 676.050 ;
        RECT 475.950 674.400 484.050 675.600 ;
        RECT 475.950 673.950 478.050 674.400 ;
        RECT 481.950 673.950 484.050 674.400 ;
        RECT 520.950 674.400 525.600 675.600 ;
        RECT 559.950 675.600 562.050 676.050 ;
        RECT 571.950 675.600 574.050 676.050 ;
        RECT 559.950 674.400 574.050 675.600 ;
        RECT 520.950 673.950 525.000 674.400 ;
        RECT 559.950 673.950 562.050 674.400 ;
        RECT 571.950 673.950 574.050 674.400 ;
        RECT 601.950 675.600 604.050 676.050 ;
        RECT 610.950 675.600 613.050 676.050 ;
        RECT 601.950 674.400 613.050 675.600 ;
        RECT 659.400 675.600 660.600 683.100 ;
        RECT 669.000 682.950 673.050 683.400 ;
        RECT 697.950 682.950 700.050 685.050 ;
        RECT 703.950 684.600 706.050 685.050 ;
        RECT 715.950 684.600 718.050 685.050 ;
        RECT 703.950 683.400 718.050 684.600 ;
        RECT 703.950 682.950 706.050 683.400 ;
        RECT 715.950 682.950 718.050 683.400 ;
        RECT 748.950 684.600 751.050 685.200 ;
        RECT 763.950 684.600 766.050 685.200 ;
        RECT 784.950 684.600 787.050 685.200 ;
        RECT 748.950 683.400 787.050 684.600 ;
        RECT 748.950 683.100 751.050 683.400 ;
        RECT 763.950 683.100 766.050 683.400 ;
        RECT 784.950 683.100 787.050 683.400 ;
        RECT 805.950 684.600 810.000 685.050 ;
        RECT 835.950 684.600 838.050 685.050 ;
        RECT 853.950 684.600 856.050 685.050 ;
        RECT 805.950 682.950 810.600 684.600 ;
        RECT 835.950 683.400 856.050 684.600 ;
        RECT 835.950 682.950 838.050 683.400 ;
        RECT 853.950 682.950 856.050 683.400 ;
        RECT 698.400 679.050 699.600 682.950 ;
        RECT 809.400 679.050 810.600 682.950 ;
        RECT 694.950 677.400 699.600 679.050 ;
        RECT 793.950 678.450 796.050 678.900 ;
        RECT 802.950 678.450 805.050 678.900 ;
        RECT 694.950 676.950 699.000 677.400 ;
        RECT 793.950 677.250 805.050 678.450 ;
        RECT 793.950 676.800 796.050 677.250 ;
        RECT 802.950 676.800 805.050 677.250 ;
        RECT 808.950 676.950 811.050 679.050 ;
        RECT 829.950 678.600 832.050 679.050 ;
        RECT 835.950 678.600 838.050 678.750 ;
        RECT 829.950 678.300 838.050 678.600 ;
        RECT 856.950 678.300 859.050 678.750 ;
        RECT 829.950 677.400 859.050 678.300 ;
        RECT 829.950 676.950 832.050 677.400 ;
        RECT 835.950 677.100 859.050 677.400 ;
        RECT 835.950 676.650 838.050 677.100 ;
        RECT 856.950 676.650 859.050 677.100 ;
        RECT 670.950 675.600 673.050 675.900 ;
        RECT 659.400 674.400 673.050 675.600 ;
        RECT 601.950 673.950 604.050 674.400 ;
        RECT 610.950 673.950 613.050 674.400 ;
        RECT 520.950 673.500 523.050 673.950 ;
        RECT 670.950 673.800 673.050 674.400 ;
        RECT 712.950 675.600 715.050 676.050 ;
        RECT 718.950 675.600 721.050 676.050 ;
        RECT 712.950 674.400 721.050 675.600 ;
        RECT 712.950 673.950 715.050 674.400 ;
        RECT 718.950 673.950 721.050 674.400 ;
        RECT 757.950 675.600 760.050 676.050 ;
        RECT 766.950 675.600 769.050 676.050 ;
        RECT 757.950 674.400 769.050 675.600 ;
        RECT 757.950 673.950 760.050 674.400 ;
        RECT 766.950 673.950 769.050 674.400 ;
        RECT 121.950 672.600 124.050 673.050 ;
        RECT 145.950 672.600 148.050 673.050 ;
        RECT 154.950 672.600 157.050 673.050 ;
        RECT 121.950 671.400 157.050 672.600 ;
        RECT 121.950 670.950 124.050 671.400 ;
        RECT 145.950 670.950 148.050 671.400 ;
        RECT 154.950 670.950 157.050 671.400 ;
        RECT 193.950 672.600 196.050 673.050 ;
        RECT 220.950 672.600 223.050 673.050 ;
        RECT 193.950 671.400 223.050 672.600 ;
        RECT 193.950 670.950 196.050 671.400 ;
        RECT 220.950 670.950 223.050 671.400 ;
        RECT 298.950 672.600 301.050 673.050 ;
        RECT 307.950 672.600 310.050 673.050 ;
        RECT 331.950 672.600 334.050 673.050 ;
        RECT 298.950 671.400 334.050 672.600 ;
        RECT 298.950 670.950 301.050 671.400 ;
        RECT 307.950 670.950 310.050 671.400 ;
        RECT 331.950 670.950 334.050 671.400 ;
        RECT 391.950 672.600 394.050 673.050 ;
        RECT 406.950 672.600 409.050 673.050 ;
        RECT 418.950 672.600 421.050 673.050 ;
        RECT 391.950 671.400 421.050 672.600 ;
        RECT 391.950 670.950 394.050 671.400 ;
        RECT 406.950 670.950 409.050 671.400 ;
        RECT 418.950 670.950 421.050 671.400 ;
        RECT 451.950 672.600 454.050 673.050 ;
        RECT 493.950 672.600 496.050 673.050 ;
        RECT 451.950 671.400 496.050 672.600 ;
        RECT 451.950 670.950 454.050 671.400 ;
        RECT 493.950 670.950 496.050 671.400 ;
        RECT 535.950 672.600 538.050 673.050 ;
        RECT 550.950 672.600 553.050 673.050 ;
        RECT 535.950 671.400 553.050 672.600 ;
        RECT 535.950 670.950 538.050 671.400 ;
        RECT 550.950 670.950 553.050 671.400 ;
        RECT 628.950 672.600 631.050 673.050 ;
        RECT 640.950 672.600 643.050 673.050 ;
        RECT 628.950 671.400 643.050 672.600 ;
        RECT 628.950 670.950 631.050 671.400 ;
        RECT 640.950 670.950 643.050 671.400 ;
        RECT 655.950 672.600 658.050 673.050 ;
        RECT 700.950 672.600 703.050 673.050 ;
        RECT 721.950 672.600 724.050 673.050 ;
        RECT 655.950 671.400 724.050 672.600 ;
        RECT 655.950 670.950 658.050 671.400 ;
        RECT 700.950 670.950 703.050 671.400 ;
        RECT 721.950 670.950 724.050 671.400 ;
        RECT 814.950 672.600 817.050 673.050 ;
        RECT 820.950 672.600 823.050 673.050 ;
        RECT 841.950 672.600 844.050 673.050 ;
        RECT 814.950 671.400 844.050 672.600 ;
        RECT 814.950 670.950 817.050 671.400 ;
        RECT 820.950 670.950 823.050 671.400 ;
        RECT 841.950 670.950 844.050 671.400 ;
        RECT 19.950 669.600 22.050 670.050 ;
        RECT 58.950 669.600 61.050 670.050 ;
        RECT 19.950 668.400 61.050 669.600 ;
        RECT 19.950 667.950 22.050 668.400 ;
        RECT 58.950 667.950 61.050 668.400 ;
        RECT 115.950 669.600 118.050 670.050 ;
        RECT 127.950 669.600 130.050 670.050 ;
        RECT 115.950 668.400 130.050 669.600 ;
        RECT 115.950 667.950 118.050 668.400 ;
        RECT 127.950 667.950 130.050 668.400 ;
        RECT 184.950 669.600 187.050 670.050 ;
        RECT 217.950 669.600 220.050 670.050 ;
        RECT 184.950 668.400 220.050 669.600 ;
        RECT 184.950 667.950 187.050 668.400 ;
        RECT 217.950 667.950 220.050 668.400 ;
        RECT 238.950 669.600 241.050 670.050 ;
        RECT 295.950 669.600 298.050 670.050 ;
        RECT 238.950 668.400 298.050 669.600 ;
        RECT 238.950 667.950 241.050 668.400 ;
        RECT 295.950 667.950 298.050 668.400 ;
        RECT 370.950 669.600 373.050 670.050 ;
        RECT 379.950 669.600 382.050 670.050 ;
        RECT 370.950 668.400 382.050 669.600 ;
        RECT 370.950 667.950 373.050 668.400 ;
        RECT 379.950 667.950 382.050 668.400 ;
        RECT 421.950 669.600 424.050 670.050 ;
        RECT 466.950 669.600 469.050 670.050 ;
        RECT 421.950 668.400 469.050 669.600 ;
        RECT 421.950 667.950 424.050 668.400 ;
        RECT 466.950 667.950 469.050 668.400 ;
        RECT 514.950 669.600 517.050 670.050 ;
        RECT 526.950 669.600 529.050 670.050 ;
        RECT 514.950 668.400 529.050 669.600 ;
        RECT 514.950 667.950 517.050 668.400 ;
        RECT 526.950 667.950 529.050 668.400 ;
        RECT 712.950 669.600 715.050 670.050 ;
        RECT 751.950 669.600 754.050 670.050 ;
        RECT 760.950 669.600 763.050 670.050 ;
        RECT 712.950 668.400 763.050 669.600 ;
        RECT 712.950 667.950 715.050 668.400 ;
        RECT 751.950 667.950 754.050 668.400 ;
        RECT 760.950 667.950 763.050 668.400 ;
        RECT 766.950 669.600 769.050 670.050 ;
        RECT 784.950 669.600 787.050 670.050 ;
        RECT 766.950 668.400 787.050 669.600 ;
        RECT 766.950 667.950 769.050 668.400 ;
        RECT 784.950 667.950 787.050 668.400 ;
        RECT 46.950 666.600 49.050 667.050 ;
        RECT 79.950 666.600 82.050 667.050 ;
        RECT 106.950 666.600 109.050 667.050 ;
        RECT 46.950 665.400 109.050 666.600 ;
        RECT 46.950 664.950 49.050 665.400 ;
        RECT 79.950 664.950 82.050 665.400 ;
        RECT 106.950 664.950 109.050 665.400 ;
        RECT 223.950 666.600 226.050 667.050 ;
        RECT 289.950 666.600 292.050 667.050 ;
        RECT 223.950 665.400 292.050 666.600 ;
        RECT 223.950 664.950 226.050 665.400 ;
        RECT 289.950 664.950 292.050 665.400 ;
        RECT 325.950 666.600 328.050 667.050 ;
        RECT 331.950 666.600 334.050 667.050 ;
        RECT 325.950 665.400 334.050 666.600 ;
        RECT 325.950 664.950 328.050 665.400 ;
        RECT 331.950 664.950 334.050 665.400 ;
        RECT 397.950 666.600 400.050 667.050 ;
        RECT 415.950 666.600 418.050 667.050 ;
        RECT 448.950 666.600 451.050 667.050 ;
        RECT 397.950 665.400 451.050 666.600 ;
        RECT 397.950 664.950 400.050 665.400 ;
        RECT 415.950 664.950 418.050 665.400 ;
        RECT 448.950 664.950 451.050 665.400 ;
        RECT 538.950 666.600 541.050 667.050 ;
        RECT 547.950 666.600 550.050 667.050 ;
        RECT 538.950 665.400 550.050 666.600 ;
        RECT 538.950 664.950 541.050 665.400 ;
        RECT 547.950 664.950 550.050 665.400 ;
        RECT 604.950 666.600 607.050 667.050 ;
        RECT 655.950 666.600 658.050 667.050 ;
        RECT 604.950 665.400 658.050 666.600 ;
        RECT 604.950 664.950 607.050 665.400 ;
        RECT 655.950 664.950 658.050 665.400 ;
        RECT 736.950 666.600 739.050 667.050 ;
        RECT 781.950 666.600 784.050 667.050 ;
        RECT 736.950 665.400 784.050 666.600 ;
        RECT 736.950 664.950 739.050 665.400 ;
        RECT 781.950 664.950 784.050 665.400 ;
        RECT 163.950 663.600 166.050 664.050 ;
        RECT 175.950 663.600 178.050 664.050 ;
        RECT 163.950 662.400 178.050 663.600 ;
        RECT 163.950 661.950 166.050 662.400 ;
        RECT 175.950 661.950 178.050 662.400 ;
        RECT 202.950 663.600 205.050 664.050 ;
        RECT 214.950 663.600 217.050 664.050 ;
        RECT 202.950 662.400 217.050 663.600 ;
        RECT 202.950 661.950 205.050 662.400 ;
        RECT 214.950 661.950 217.050 662.400 ;
        RECT 229.950 663.600 232.050 664.050 ;
        RECT 241.950 663.600 244.050 664.050 ;
        RECT 229.950 662.400 244.050 663.600 ;
        RECT 229.950 661.950 232.050 662.400 ;
        RECT 241.950 661.950 244.050 662.400 ;
        RECT 364.950 663.600 367.050 664.050 ;
        RECT 370.950 663.600 373.050 664.050 ;
        RECT 364.950 662.400 373.050 663.600 ;
        RECT 364.950 661.950 367.050 662.400 ;
        RECT 370.950 661.950 373.050 662.400 ;
        RECT 376.950 663.600 379.050 664.050 ;
        RECT 454.950 663.600 457.050 664.050 ;
        RECT 376.950 662.400 457.050 663.600 ;
        RECT 376.950 661.950 379.050 662.400 ;
        RECT 454.950 661.950 457.050 662.400 ;
        RECT 463.950 663.600 466.050 664.050 ;
        RECT 502.950 663.600 505.050 664.050 ;
        RECT 463.950 662.400 505.050 663.600 ;
        RECT 463.950 661.950 466.050 662.400 ;
        RECT 502.950 661.950 505.050 662.400 ;
        RECT 574.950 663.600 577.050 664.050 ;
        RECT 631.950 663.600 634.050 664.050 ;
        RECT 646.950 663.600 649.050 664.050 ;
        RECT 691.950 663.600 694.050 664.050 ;
        RECT 574.950 662.400 694.050 663.600 ;
        RECT 574.950 661.950 577.050 662.400 ;
        RECT 631.950 661.950 634.050 662.400 ;
        RECT 646.950 661.950 649.050 662.400 ;
        RECT 691.950 661.950 694.050 662.400 ;
        RECT 796.950 663.600 799.050 664.050 ;
        RECT 841.950 663.600 844.050 664.050 ;
        RECT 796.950 662.400 844.050 663.600 ;
        RECT 796.950 661.950 799.050 662.400 ;
        RECT 841.950 661.950 844.050 662.400 ;
        RECT 139.950 660.600 142.050 661.050 ;
        RECT 148.950 660.600 151.050 661.050 ;
        RECT 139.950 659.400 151.050 660.600 ;
        RECT 139.950 658.950 142.050 659.400 ;
        RECT 148.950 658.950 151.050 659.400 ;
        RECT 208.950 660.600 211.050 661.050 ;
        RECT 238.950 660.600 241.050 661.050 ;
        RECT 208.950 659.400 241.050 660.600 ;
        RECT 208.950 658.950 211.050 659.400 ;
        RECT 238.950 658.950 241.050 659.400 ;
        RECT 259.950 660.600 262.050 661.050 ;
        RECT 322.950 660.600 325.050 661.050 ;
        RECT 355.950 660.600 358.050 661.050 ;
        RECT 259.950 659.400 285.600 660.600 ;
        RECT 259.950 658.950 262.050 659.400 ;
        RECT 13.950 657.600 16.050 658.050 ;
        RECT 34.950 657.600 37.050 658.050 ;
        RECT 43.950 657.600 46.050 658.050 ;
        RECT 13.950 656.400 46.050 657.600 ;
        RECT 13.950 655.950 16.050 656.400 ;
        RECT 34.950 655.950 37.050 656.400 ;
        RECT 43.950 655.950 46.050 656.400 ;
        RECT 64.950 657.600 67.050 658.050 ;
        RECT 76.950 657.600 79.050 658.050 ;
        RECT 88.950 657.600 91.050 658.050 ;
        RECT 97.950 657.600 100.050 658.050 ;
        RECT 64.950 656.400 100.050 657.600 ;
        RECT 64.950 655.950 67.050 656.400 ;
        RECT 76.950 655.950 79.050 656.400 ;
        RECT 88.950 655.950 91.050 656.400 ;
        RECT 97.950 655.950 100.050 656.400 ;
        RECT 190.950 657.600 193.050 658.050 ;
        RECT 196.950 657.600 199.050 658.050 ;
        RECT 190.950 656.400 199.050 657.600 ;
        RECT 190.950 655.950 193.050 656.400 ;
        RECT 196.950 655.950 199.050 656.400 ;
        RECT 220.950 657.600 223.050 658.050 ;
        RECT 265.950 657.600 268.050 658.050 ;
        RECT 277.950 657.600 280.050 658.050 ;
        RECT 220.950 656.400 258.600 657.600 ;
        RECT 220.950 655.950 223.050 656.400 ;
        RECT 55.950 654.600 58.050 655.050 ;
        RECT 47.400 653.400 58.050 654.600 ;
        RECT 13.950 650.100 16.050 652.200 ;
        RECT 19.950 651.600 22.050 652.050 ;
        RECT 28.950 651.600 31.050 652.200 ;
        RECT 19.950 650.400 31.050 651.600 ;
        RECT 14.400 642.600 15.600 650.100 ;
        RECT 19.950 649.950 22.050 650.400 ;
        RECT 28.950 650.100 31.050 650.400 ;
        RECT 47.400 645.900 48.600 653.400 ;
        RECT 55.950 652.950 58.050 653.400 ;
        RECT 205.950 652.950 208.050 655.050 ;
        RECT 49.950 651.600 52.050 652.200 ;
        RECT 49.950 650.400 57.600 651.600 ;
        RECT 49.950 650.100 52.050 650.400 ;
        RECT 56.400 646.050 57.600 650.400 ;
        RECT 61.950 648.600 64.050 652.050 ;
        RECT 67.950 650.250 70.050 652.350 ;
        RECT 73.950 651.600 76.050 652.350 ;
        RECT 100.950 651.600 103.050 651.900 ;
        RECT 73.950 650.400 103.050 651.600 ;
        RECT 73.950 650.250 76.050 650.400 ;
        RECT 61.950 648.000 66.600 648.600 ;
        RECT 62.400 647.400 66.600 648.000 ;
        RECT 31.950 645.600 34.050 645.900 ;
        RECT 46.950 645.600 49.050 645.900 ;
        RECT 31.950 644.400 49.050 645.600 ;
        RECT 31.950 643.800 34.050 644.400 ;
        RECT 46.950 643.800 49.050 644.400 ;
        RECT 55.950 643.950 58.050 646.050 ;
        RECT 52.950 642.600 55.050 643.050 ;
        RECT 14.400 641.400 55.050 642.600 ;
        RECT 65.400 642.600 66.600 647.400 ;
        RECT 68.400 645.600 69.600 650.250 ;
        RECT 100.950 649.800 103.050 650.400 ;
        RECT 106.950 649.950 109.050 652.050 ;
        RECT 112.950 650.250 115.050 652.350 ;
        RECT 130.950 651.900 133.050 652.350 ;
        RECT 136.950 651.900 139.050 652.350 ;
        RECT 130.950 650.700 139.050 651.900 ;
        RECT 130.950 650.250 133.050 650.700 ;
        RECT 136.950 650.250 139.050 650.700 ;
        RECT 107.400 646.050 108.600 649.950 ;
        RECT 91.950 645.600 94.050 646.050 ;
        RECT 68.400 644.400 94.050 645.600 ;
        RECT 91.950 643.950 94.050 644.400 ;
        RECT 106.950 643.950 109.050 646.050 ;
        RECT 113.400 645.600 114.600 650.250 ;
        RECT 142.950 649.950 145.050 652.050 ;
        RECT 163.950 650.250 166.050 652.350 ;
        RECT 169.950 651.600 174.000 652.050 ;
        RECT 143.400 646.050 144.600 649.950 ;
        RECT 164.400 646.050 165.600 650.250 ;
        RECT 169.950 649.950 174.600 651.600 ;
        RECT 184.950 650.100 187.050 652.200 ;
        RECT 196.950 651.600 199.050 652.350 ;
        RECT 194.400 650.400 199.050 651.600 ;
        RECT 173.400 648.600 174.600 649.950 ;
        RECT 173.400 648.000 180.600 648.600 ;
        RECT 173.400 647.400 181.050 648.000 ;
        RECT 127.950 645.600 130.050 646.050 ;
        RECT 113.400 644.400 130.050 645.600 ;
        RECT 127.950 643.950 130.050 644.400 ;
        RECT 142.950 643.950 145.050 646.050 ;
        RECT 163.950 643.950 166.050 646.050 ;
        RECT 178.950 643.950 181.050 647.400 ;
        RECT 70.950 642.600 73.050 643.050 ;
        RECT 85.950 642.600 88.050 643.050 ;
        RECT 65.400 641.400 88.050 642.600 ;
        RECT 92.400 642.600 93.600 643.950 ;
        RECT 109.950 642.600 112.050 643.050 ;
        RECT 92.400 641.400 112.050 642.600 ;
        RECT 52.950 640.950 55.050 641.400 ;
        RECT 70.950 640.950 73.050 641.400 ;
        RECT 85.950 640.950 88.050 641.400 ;
        RECT 109.950 640.950 112.050 641.400 ;
        RECT 139.950 642.600 142.050 643.050 ;
        RECT 148.950 642.600 151.050 643.050 ;
        RECT 139.950 641.400 151.050 642.600 ;
        RECT 185.400 642.600 186.600 650.100 ;
        RECT 194.400 646.050 195.600 650.400 ;
        RECT 196.950 650.250 199.050 650.400 ;
        RECT 206.400 646.050 207.600 652.950 ;
        RECT 211.950 651.750 214.050 652.200 ;
        RECT 235.950 651.750 238.050 652.200 ;
        RECT 211.950 650.550 238.050 651.750 ;
        RECT 211.950 650.100 214.050 650.550 ;
        RECT 235.950 650.100 238.050 650.550 ;
        RECT 244.950 651.600 247.050 652.050 ;
        RECT 253.950 651.600 256.050 652.350 ;
        RECT 244.950 650.400 256.050 651.600 ;
        RECT 236.400 648.600 237.600 650.100 ;
        RECT 244.950 649.950 247.050 650.400 ;
        RECT 253.950 650.250 256.050 650.400 ;
        RECT 257.400 648.600 258.600 656.400 ;
        RECT 265.950 656.400 280.050 657.600 ;
        RECT 284.400 657.600 285.600 659.400 ;
        RECT 322.950 659.400 358.050 660.600 ;
        RECT 322.950 658.950 325.050 659.400 ;
        RECT 355.950 658.950 358.050 659.400 ;
        RECT 445.950 660.600 448.050 661.050 ;
        RECT 592.950 660.600 595.050 661.050 ;
        RECT 604.950 660.600 607.050 661.050 ;
        RECT 445.950 659.400 519.600 660.600 ;
        RECT 445.950 658.950 448.050 659.400 ;
        RECT 518.400 658.050 519.600 659.400 ;
        RECT 592.950 659.400 607.050 660.600 ;
        RECT 592.950 658.950 595.050 659.400 ;
        RECT 604.950 658.950 607.050 659.400 ;
        RECT 610.950 660.600 613.050 661.050 ;
        RECT 628.950 660.600 631.050 661.050 ;
        RECT 610.950 659.400 631.050 660.600 ;
        RECT 610.950 658.950 613.050 659.400 ;
        RECT 628.950 658.950 631.050 659.400 ;
        RECT 706.950 660.600 709.050 661.050 ;
        RECT 763.950 660.600 766.050 661.050 ;
        RECT 772.950 660.600 775.050 661.050 ;
        RECT 706.950 659.400 775.050 660.600 ;
        RECT 706.950 658.950 709.050 659.400 ;
        RECT 763.950 658.950 766.050 659.400 ;
        RECT 772.950 658.950 775.050 659.400 ;
        RECT 826.950 660.600 829.050 661.050 ;
        RECT 835.950 660.600 838.050 661.050 ;
        RECT 826.950 659.400 838.050 660.600 ;
        RECT 826.950 658.950 829.050 659.400 ;
        RECT 835.950 658.950 838.050 659.400 ;
        RECT 325.950 657.600 328.050 658.050 ;
        RECT 284.400 656.400 328.050 657.600 ;
        RECT 265.950 655.950 268.050 656.400 ;
        RECT 277.950 655.950 280.050 656.400 ;
        RECT 325.950 655.950 328.050 656.400 ;
        RECT 364.950 657.600 367.050 658.050 ;
        RECT 388.950 657.600 391.050 658.050 ;
        RECT 364.950 656.400 391.050 657.600 ;
        RECT 364.950 655.950 367.050 656.400 ;
        RECT 388.950 655.950 391.050 656.400 ;
        RECT 424.950 657.600 427.050 658.050 ;
        RECT 442.950 657.600 445.050 658.050 ;
        RECT 424.950 656.400 445.050 657.600 ;
        RECT 424.950 655.950 427.050 656.400 ;
        RECT 442.950 655.950 445.050 656.400 ;
        RECT 484.950 657.600 487.050 658.050 ;
        RECT 502.950 657.600 505.050 658.050 ;
        RECT 484.950 656.400 505.050 657.600 ;
        RECT 484.950 655.950 487.050 656.400 ;
        RECT 502.950 655.950 505.050 656.400 ;
        RECT 517.950 657.600 520.050 658.050 ;
        RECT 529.950 657.600 532.050 658.050 ;
        RECT 517.950 656.400 532.050 657.600 ;
        RECT 517.950 655.950 520.050 656.400 ;
        RECT 529.950 655.950 532.050 656.400 ;
        RECT 598.950 657.600 601.050 658.050 ;
        RECT 727.950 657.600 730.050 658.050 ;
        RECT 742.800 657.600 744.900 658.050 ;
        RECT 598.950 656.400 630.600 657.600 ;
        RECT 598.950 655.950 601.050 656.400 ;
        RECT 328.950 654.600 331.050 655.050 ;
        RECT 337.800 654.600 339.900 655.050 ;
        RECT 328.950 653.400 339.900 654.600 ;
        RECT 328.950 652.950 331.050 653.400 ;
        RECT 337.800 652.950 339.900 653.400 ;
        RECT 340.950 654.600 343.050 655.050 ;
        RECT 361.950 654.600 364.050 655.050 ;
        RECT 340.950 653.400 364.050 654.600 ;
        RECT 340.950 652.950 343.050 653.400 ;
        RECT 361.950 652.950 364.050 653.400 ;
        RECT 448.950 654.600 451.050 655.050 ;
        RECT 499.950 654.600 502.050 655.050 ;
        RECT 604.950 654.600 607.050 655.050 ;
        RECT 613.950 654.600 616.050 655.050 ;
        RECT 448.950 653.400 495.600 654.600 ;
        RECT 448.950 652.950 451.050 653.400 ;
        RECT 298.950 651.600 301.050 652.350 ;
        RECT 307.800 651.600 309.900 652.050 ;
        RECT 298.950 650.400 309.900 651.600 ;
        RECT 298.950 650.250 301.050 650.400 ;
        RECT 307.800 649.950 309.900 650.400 ;
        RECT 310.950 651.600 313.050 652.050 ;
        RECT 325.950 651.600 328.050 652.050 ;
        RECT 343.950 651.900 346.050 652.350 ;
        RECT 349.950 651.900 352.050 652.350 ;
        RECT 310.950 650.400 324.600 651.600 ;
        RECT 310.950 649.950 313.050 650.400 ;
        RECT 236.400 648.000 249.600 648.600 ;
        RECT 236.400 647.400 250.050 648.000 ;
        RECT 257.400 647.400 264.600 648.600 ;
        RECT 193.950 643.950 196.050 646.050 ;
        RECT 205.950 643.950 208.050 646.050 ;
        RECT 247.950 643.950 250.050 647.400 ;
        RECT 263.400 645.600 264.600 647.400 ;
        RECT 323.400 646.050 324.600 650.400 ;
        RECT 325.950 650.400 342.600 651.600 ;
        RECT 325.950 649.950 328.050 650.400 ;
        RECT 341.400 648.600 342.600 650.400 ;
        RECT 343.950 650.700 352.050 651.900 ;
        RECT 343.950 650.250 346.050 650.700 ;
        RECT 349.950 650.250 352.050 650.700 ;
        RECT 355.950 651.600 358.050 652.050 ;
        RECT 364.950 651.600 367.050 652.200 ;
        RECT 355.950 650.400 367.050 651.600 ;
        RECT 355.950 649.950 358.050 650.400 ;
        RECT 364.950 650.100 367.050 650.400 ;
        RECT 388.950 650.250 391.050 652.350 ;
        RECT 406.950 651.600 409.050 652.200 ;
        RECT 427.950 651.600 430.050 652.050 ;
        RECT 395.400 650.400 409.050 651.600 ;
        RECT 341.400 647.400 387.600 648.600 ;
        RECT 268.950 645.600 271.050 646.050 ;
        RECT 263.400 644.400 271.050 645.600 ;
        RECT 268.950 643.950 271.050 644.400 ;
        RECT 307.950 645.450 310.050 645.900 ;
        RECT 313.950 645.450 316.050 645.900 ;
        RECT 307.950 644.250 316.050 645.450 ;
        RECT 323.400 644.400 328.050 646.050 ;
        RECT 307.950 643.800 310.050 644.250 ;
        RECT 313.950 643.800 316.050 644.250 ;
        RECT 324.000 643.950 328.050 644.400 ;
        RECT 346.950 645.450 349.050 645.900 ;
        RECT 373.950 645.450 376.050 645.900 ;
        RECT 346.950 644.250 376.050 645.450 ;
        RECT 346.950 643.800 349.050 644.250 ;
        RECT 373.950 643.800 376.050 644.250 ;
        RECT 202.950 642.600 205.050 643.050 ;
        RECT 185.400 641.400 205.050 642.600 ;
        RECT 139.950 640.950 142.050 641.400 ;
        RECT 148.950 640.950 151.050 641.400 ;
        RECT 202.950 640.950 205.050 641.400 ;
        RECT 274.950 642.600 277.050 643.050 ;
        RECT 301.950 642.600 304.050 643.050 ;
        RECT 274.950 641.400 304.050 642.600 ;
        RECT 386.400 642.600 387.600 647.400 ;
        RECT 389.400 646.050 390.600 650.250 ;
        RECT 395.400 646.050 396.600 650.400 ;
        RECT 406.950 650.100 409.050 650.400 ;
        RECT 410.400 650.400 430.050 651.600 ;
        RECT 388.950 643.950 391.050 646.050 ;
        RECT 394.950 643.950 397.050 646.050 ;
        RECT 410.400 645.900 411.600 650.400 ;
        RECT 427.950 649.950 430.050 650.400 ;
        RECT 463.950 651.600 466.050 652.350 ;
        RECT 494.400 651.600 495.600 653.400 ;
        RECT 499.950 653.400 546.600 654.600 ;
        RECT 499.950 652.950 502.050 653.400 ;
        RECT 538.950 651.600 541.050 652.050 ;
        RECT 463.950 650.400 486.600 651.600 ;
        RECT 494.400 650.400 541.050 651.600 ;
        RECT 463.950 650.250 466.050 650.400 ;
        RECT 451.950 648.600 454.050 649.050 ;
        RECT 422.400 648.000 454.050 648.600 ;
        RECT 421.950 647.400 454.050 648.000 ;
        RECT 485.400 648.600 486.600 650.400 ;
        RECT 538.950 649.950 541.050 650.400 ;
        RECT 545.400 648.600 546.600 653.400 ;
        RECT 604.950 653.400 616.050 654.600 ;
        RECT 629.400 654.600 630.600 656.400 ;
        RECT 727.950 656.400 744.900 657.600 ;
        RECT 727.950 655.950 730.050 656.400 ;
        RECT 742.800 655.950 744.900 656.400 ;
        RECT 745.950 657.600 748.050 658.050 ;
        RECT 751.950 657.600 754.050 658.050 ;
        RECT 745.950 656.400 754.050 657.600 ;
        RECT 745.950 655.950 748.050 656.400 ;
        RECT 751.950 655.950 754.050 656.400 ;
        RECT 643.950 654.600 646.050 655.050 ;
        RECT 629.400 653.400 646.050 654.600 ;
        RECT 604.950 652.950 607.050 653.400 ;
        RECT 613.950 652.950 616.050 653.400 ;
        RECT 643.950 652.950 646.050 653.400 ;
        RECT 649.950 654.600 652.050 655.050 ;
        RECT 664.950 654.600 667.050 655.050 ;
        RECT 765.000 654.600 769.050 655.050 ;
        RECT 805.800 654.600 807.900 655.050 ;
        RECT 649.950 653.400 667.050 654.600 ;
        RECT 649.950 652.950 652.050 653.400 ;
        RECT 664.950 652.950 667.050 653.400 ;
        RECT 764.400 652.950 769.050 654.600 ;
        RECT 797.400 653.400 807.900 654.600 ;
        RECT 577.950 651.600 580.050 652.050 ;
        RECT 572.400 650.400 580.050 651.600 ;
        RECT 572.400 648.600 573.600 650.400 ;
        RECT 577.950 649.950 580.050 650.400 ;
        RECT 583.950 651.600 586.050 652.050 ;
        RECT 616.950 651.600 619.050 651.900 ;
        RECT 685.950 651.600 688.050 652.350 ;
        RECT 583.950 650.400 619.050 651.600 ;
        RECT 583.950 649.950 586.050 650.400 ;
        RECT 616.950 649.800 619.050 650.400 ;
        RECT 668.400 650.400 688.050 651.600 ;
        RECT 661.950 648.600 664.050 649.050 ;
        RECT 668.400 648.600 669.600 650.400 ;
        RECT 685.950 650.250 688.050 650.400 ;
        RECT 706.950 650.250 709.050 652.350 ;
        RECT 485.400 648.000 489.600 648.600 ;
        RECT 533.400 648.000 546.600 648.600 ;
        RECT 566.400 648.000 621.600 648.600 ;
        RECT 485.400 647.400 490.050 648.000 ;
        RECT 409.950 643.800 412.050 645.900 ;
        RECT 421.950 643.950 424.050 647.400 ;
        RECT 451.950 646.950 454.050 647.400 ;
        RECT 487.950 643.950 490.050 647.400 ;
        RECT 532.950 647.400 546.600 648.000 ;
        RECT 565.950 647.400 621.600 648.000 ;
        RECT 511.950 645.600 514.050 646.050 ;
        RECT 526.950 645.600 529.050 646.050 ;
        RECT 511.950 644.400 529.050 645.600 ;
        RECT 511.950 643.950 514.050 644.400 ;
        RECT 526.950 643.950 529.050 644.400 ;
        RECT 532.950 643.950 535.050 647.400 ;
        RECT 565.950 643.950 568.050 647.400 ;
        RECT 586.950 645.600 589.050 646.050 ;
        RECT 601.950 645.600 604.050 646.050 ;
        RECT 610.950 645.600 613.050 646.050 ;
        RECT 586.950 644.400 613.050 645.600 ;
        RECT 586.950 643.950 589.050 644.400 ;
        RECT 601.950 643.950 604.050 644.400 ;
        RECT 610.950 643.950 613.050 644.400 ;
        RECT 403.950 642.600 406.050 643.050 ;
        RECT 386.400 641.400 406.050 642.600 ;
        RECT 274.950 640.950 277.050 641.400 ;
        RECT 301.950 640.950 304.050 641.400 ;
        RECT 403.950 640.950 406.050 641.400 ;
        RECT 436.950 642.600 439.050 643.050 ;
        RECT 493.950 642.600 496.050 643.050 ;
        RECT 436.950 641.400 496.050 642.600 ;
        RECT 436.950 640.950 439.050 641.400 ;
        RECT 493.950 640.950 496.050 641.400 ;
        RECT 508.950 642.600 511.050 643.050 ;
        RECT 541.950 642.600 544.050 643.050 ;
        RECT 556.950 642.600 559.050 643.050 ;
        RECT 508.950 641.400 528.600 642.600 ;
        RECT 508.950 640.950 511.050 641.400 ;
        RECT 10.950 639.600 13.050 640.050 ;
        RECT 25.950 639.600 28.050 640.050 ;
        RECT 10.950 638.400 28.050 639.600 ;
        RECT 10.950 637.950 13.050 638.400 ;
        RECT 25.950 637.950 28.050 638.400 ;
        RECT 211.950 639.600 214.050 640.050 ;
        RECT 250.950 639.600 253.050 640.050 ;
        RECT 256.950 639.600 259.050 639.900 ;
        RECT 211.950 638.400 259.050 639.600 ;
        RECT 211.950 637.950 214.050 638.400 ;
        RECT 250.950 637.950 253.050 638.400 ;
        RECT 256.950 637.800 259.050 638.400 ;
        RECT 277.950 639.600 280.050 640.050 ;
        RECT 310.950 639.600 313.050 640.050 ;
        RECT 277.950 638.400 313.050 639.600 ;
        RECT 277.950 637.950 280.050 638.400 ;
        RECT 310.950 637.950 313.050 638.400 ;
        RECT 466.950 639.600 469.050 640.050 ;
        RECT 475.950 639.600 478.050 640.050 ;
        RECT 466.950 638.400 478.050 639.600 ;
        RECT 466.950 637.950 469.050 638.400 ;
        RECT 475.950 637.950 478.050 638.400 ;
        RECT 505.950 639.600 508.050 640.050 ;
        RECT 523.950 639.600 526.050 640.050 ;
        RECT 505.950 638.400 526.050 639.600 ;
        RECT 527.400 639.600 528.600 641.400 ;
        RECT 541.950 641.400 559.050 642.600 ;
        RECT 620.400 642.600 621.600 647.400 ;
        RECT 661.950 647.400 669.600 648.600 ;
        RECT 661.950 646.950 664.050 647.400 ;
        RECT 685.950 645.600 688.050 646.050 ;
        RECT 707.400 645.600 708.600 650.250 ;
        RECT 730.950 650.100 733.050 652.200 ;
        RECT 748.950 651.600 751.050 652.350 ;
        RECT 754.800 651.600 756.900 652.050 ;
        RECT 748.950 650.400 756.900 651.600 ;
        RECT 748.950 650.250 751.050 650.400 ;
        RECT 721.950 648.600 724.050 649.050 ;
        RECT 731.400 648.600 732.600 650.100 ;
        RECT 754.800 649.950 756.900 650.400 ;
        RECT 757.950 649.950 760.050 652.050 ;
        RECT 721.950 647.400 732.600 648.600 ;
        RECT 721.950 646.950 724.050 647.400 ;
        RECT 758.400 646.050 759.600 649.950 ;
        RECT 764.400 646.050 765.600 652.950 ;
        RECT 769.950 651.600 772.050 652.350 ;
        RECT 797.400 652.050 798.600 653.400 ;
        RECT 805.800 652.950 807.900 653.400 ;
        RECT 775.950 651.600 778.050 652.050 ;
        RECT 769.950 650.400 778.050 651.600 ;
        RECT 769.950 650.250 772.050 650.400 ;
        RECT 775.950 649.950 778.050 650.400 ;
        RECT 793.950 650.400 798.600 652.050 ;
        RECT 808.950 651.600 811.050 655.050 ;
        RECT 817.950 654.600 820.050 655.050 ;
        RECT 806.400 651.000 811.050 651.600 ;
        RECT 812.400 653.400 820.050 654.600 ;
        RECT 806.400 650.400 810.600 651.000 ;
        RECT 793.950 649.950 798.000 650.400 ;
        RECT 806.400 646.050 807.600 650.400 ;
        RECT 812.400 646.050 813.600 653.400 ;
        RECT 817.950 652.950 820.050 653.400 ;
        RECT 826.950 654.600 829.050 655.050 ;
        RECT 832.950 654.600 835.050 655.050 ;
        RECT 826.950 653.400 835.050 654.600 ;
        RECT 826.950 652.950 829.050 653.400 ;
        RECT 832.950 652.950 835.050 653.400 ;
        RECT 829.950 651.600 832.050 652.050 ;
        RECT 818.400 650.400 832.050 651.600 ;
        RECT 818.400 646.050 819.600 650.400 ;
        RECT 829.950 649.950 832.050 650.400 ;
        RECT 835.950 651.600 838.050 652.050 ;
        RECT 847.950 651.600 850.050 652.350 ;
        RECT 853.950 651.600 856.050 652.050 ;
        RECT 835.950 650.400 843.450 651.600 ;
        RECT 835.950 649.950 838.050 650.400 ;
        RECT 842.250 646.050 843.450 650.400 ;
        RECT 847.950 650.400 856.050 651.600 ;
        RECT 847.950 650.250 850.050 650.400 ;
        RECT 853.950 649.950 856.050 650.400 ;
        RECT 685.950 644.400 708.600 645.600 ;
        RECT 745.950 645.600 748.050 646.050 ;
        RECT 751.950 645.600 754.050 646.050 ;
        RECT 745.950 644.400 754.050 645.600 ;
        RECT 685.950 643.950 688.050 644.400 ;
        RECT 745.950 643.950 748.050 644.400 ;
        RECT 751.950 643.950 754.050 644.400 ;
        RECT 757.950 643.950 760.050 646.050 ;
        RECT 763.950 643.950 766.050 646.050 ;
        RECT 775.950 645.600 778.050 646.050 ;
        RECT 787.950 645.600 790.050 646.050 ;
        RECT 775.950 644.400 790.050 645.600 ;
        RECT 775.950 643.950 778.050 644.400 ;
        RECT 787.950 643.950 790.050 644.400 ;
        RECT 805.950 643.950 808.050 646.050 ;
        RECT 811.950 643.950 814.050 646.050 ;
        RECT 817.950 643.950 820.050 646.050 ;
        RECT 841.800 643.950 843.900 646.050 ;
        RECT 844.950 645.600 847.050 646.050 ;
        RECT 859.950 645.600 862.050 646.050 ;
        RECT 844.950 644.400 862.050 645.600 ;
        RECT 844.950 643.950 847.050 644.400 ;
        RECT 859.950 643.950 862.050 644.400 ;
        RECT 628.950 642.600 631.050 643.050 ;
        RECT 620.400 641.400 631.050 642.600 ;
        RECT 541.950 640.950 544.050 641.400 ;
        RECT 556.950 640.950 559.050 641.400 ;
        RECT 628.950 640.950 631.050 641.400 ;
        RECT 655.950 642.600 658.050 643.050 ;
        RECT 667.950 642.600 670.050 643.050 ;
        RECT 655.950 641.400 670.050 642.600 ;
        RECT 655.950 640.950 658.050 641.400 ;
        RECT 667.950 640.950 670.050 641.400 ;
        RECT 538.950 639.600 541.050 640.050 ;
        RECT 527.400 638.400 541.050 639.600 ;
        RECT 505.950 637.950 508.050 638.400 ;
        RECT 523.950 637.950 526.050 638.400 ;
        RECT 538.950 637.950 541.050 638.400 ;
        RECT 559.950 639.600 562.050 640.050 ;
        RECT 586.950 639.600 589.050 640.050 ;
        RECT 559.950 638.400 589.050 639.600 ;
        RECT 559.950 637.950 562.050 638.400 ;
        RECT 586.950 637.950 589.050 638.400 ;
        RECT 631.950 639.600 634.050 640.050 ;
        RECT 721.950 639.600 724.050 640.050 ;
        RECT 739.950 639.600 742.050 640.050 ;
        RECT 631.950 638.400 742.050 639.600 ;
        RECT 631.950 637.950 634.050 638.400 ;
        RECT 721.950 637.950 724.050 638.400 ;
        RECT 739.950 637.950 742.050 638.400 ;
        RECT 787.950 639.600 790.050 640.050 ;
        RECT 808.950 639.600 811.050 640.050 ;
        RECT 838.950 639.600 841.050 640.050 ;
        RECT 787.950 638.400 841.050 639.600 ;
        RECT 787.950 637.950 790.050 638.400 ;
        RECT 808.950 637.950 811.050 638.400 ;
        RECT 838.950 637.950 841.050 638.400 ;
        RECT 52.950 636.600 55.050 637.050 ;
        RECT 61.950 636.600 64.050 637.050 ;
        RECT 163.950 636.600 166.050 637.050 ;
        RECT 52.950 635.400 166.050 636.600 ;
        RECT 52.950 634.950 55.050 635.400 ;
        RECT 61.950 634.950 64.050 635.400 ;
        RECT 163.950 634.950 166.050 635.400 ;
        RECT 181.950 636.600 184.050 637.050 ;
        RECT 205.950 636.600 208.050 637.050 ;
        RECT 220.950 636.600 223.050 637.050 ;
        RECT 181.950 635.400 223.050 636.600 ;
        RECT 181.950 634.950 184.050 635.400 ;
        RECT 205.950 634.950 208.050 635.400 ;
        RECT 220.950 634.950 223.050 635.400 ;
        RECT 247.950 636.600 250.050 637.050 ;
        RECT 268.800 636.600 270.900 637.050 ;
        RECT 247.950 635.400 270.900 636.600 ;
        RECT 247.950 634.950 250.050 635.400 ;
        RECT 268.800 634.950 270.900 635.400 ;
        RECT 271.950 636.600 274.050 637.050 ;
        RECT 316.950 636.600 319.050 637.050 ;
        RECT 271.950 635.400 319.050 636.600 ;
        RECT 271.950 634.950 274.050 635.400 ;
        RECT 316.950 634.950 319.050 635.400 ;
        RECT 370.950 636.600 373.050 637.050 ;
        RECT 379.950 636.600 382.050 637.050 ;
        RECT 370.950 635.400 382.050 636.600 ;
        RECT 370.950 634.950 373.050 635.400 ;
        RECT 379.950 634.950 382.050 635.400 ;
        RECT 466.950 636.600 469.050 636.900 ;
        RECT 481.800 636.600 483.900 637.050 ;
        RECT 466.950 635.400 483.900 636.600 ;
        RECT 466.950 634.800 469.050 635.400 ;
        RECT 481.800 634.950 483.900 635.400 ;
        RECT 553.950 636.600 556.050 637.050 ;
        RECT 574.950 636.600 577.050 637.050 ;
        RECT 553.950 635.400 577.050 636.600 ;
        RECT 553.950 634.950 556.050 635.400 ;
        RECT 574.950 634.950 577.050 635.400 ;
        RECT 652.950 636.600 655.050 637.050 ;
        RECT 661.950 636.600 664.050 637.050 ;
        RECT 709.950 636.600 712.050 637.050 ;
        RECT 652.950 635.400 712.050 636.600 ;
        RECT 652.950 634.950 655.050 635.400 ;
        RECT 661.950 634.950 664.050 635.400 ;
        RECT 709.950 634.950 712.050 635.400 ;
        RECT 754.950 636.600 757.050 637.050 ;
        RECT 784.950 636.600 787.050 636.900 ;
        RECT 754.950 635.400 787.050 636.600 ;
        RECT 754.950 634.950 757.050 635.400 ;
        RECT 784.950 634.800 787.050 635.400 ;
        RECT 799.950 636.600 802.050 637.050 ;
        RECT 823.950 636.600 826.050 637.050 ;
        RECT 799.950 635.400 826.050 636.600 ;
        RECT 799.950 634.950 802.050 635.400 ;
        RECT 823.950 634.950 826.050 635.400 ;
        RECT 64.950 633.600 67.050 634.050 ;
        RECT 76.950 633.600 79.050 634.050 ;
        RECT 64.950 632.400 79.050 633.600 ;
        RECT 64.950 631.950 67.050 632.400 ;
        RECT 76.950 631.950 79.050 632.400 ;
        RECT 175.950 633.600 178.050 634.050 ;
        RECT 199.950 633.600 202.050 634.050 ;
        RECT 175.950 632.400 202.050 633.600 ;
        RECT 175.950 631.950 178.050 632.400 ;
        RECT 199.950 631.950 202.050 632.400 ;
        RECT 208.950 633.600 211.050 634.050 ;
        RECT 277.800 633.600 279.900 634.050 ;
        RECT 208.950 632.400 279.900 633.600 ;
        RECT 208.950 631.950 211.050 632.400 ;
        RECT 277.800 631.950 279.900 632.400 ;
        RECT 280.950 633.600 283.050 634.050 ;
        RECT 307.950 633.600 310.050 634.050 ;
        RECT 280.950 632.400 310.050 633.600 ;
        RECT 280.950 631.950 283.050 632.400 ;
        RECT 307.950 631.950 310.050 632.400 ;
        RECT 385.950 633.600 388.050 634.050 ;
        RECT 433.950 633.600 436.050 634.050 ;
        RECT 385.950 632.400 436.050 633.600 ;
        RECT 385.950 631.950 388.050 632.400 ;
        RECT 433.950 631.950 436.050 632.400 ;
        RECT 445.950 633.600 448.050 634.050 ;
        RECT 514.950 633.600 517.050 634.050 ;
        RECT 445.950 632.400 517.050 633.600 ;
        RECT 445.950 631.950 448.050 632.400 ;
        RECT 514.950 631.950 517.050 632.400 ;
        RECT 523.950 633.600 526.050 634.050 ;
        RECT 592.950 633.600 595.050 634.050 ;
        RECT 523.950 632.400 595.050 633.600 ;
        RECT 523.950 631.950 526.050 632.400 ;
        RECT 592.950 631.950 595.050 632.400 ;
        RECT 667.950 633.600 670.050 634.050 ;
        RECT 688.950 633.600 691.050 634.050 ;
        RECT 703.950 633.600 706.050 634.050 ;
        RECT 667.950 632.400 706.050 633.600 ;
        RECT 667.950 631.950 670.050 632.400 ;
        RECT 688.950 631.950 691.050 632.400 ;
        RECT 703.950 631.950 706.050 632.400 ;
        RECT 727.950 633.600 730.050 634.050 ;
        RECT 760.950 633.600 763.050 634.050 ;
        RECT 727.950 632.400 763.050 633.600 ;
        RECT 727.950 631.950 730.050 632.400 ;
        RECT 760.950 631.950 763.050 632.400 ;
        RECT 118.950 630.600 121.050 631.050 ;
        RECT 133.950 630.600 136.050 631.050 ;
        RECT 187.950 630.600 190.050 631.050 ;
        RECT 118.950 629.400 190.050 630.600 ;
        RECT 118.950 628.950 121.050 629.400 ;
        RECT 133.950 628.950 136.050 629.400 ;
        RECT 187.950 628.950 190.050 629.400 ;
        RECT 199.950 630.600 202.050 630.900 ;
        RECT 292.950 630.600 295.050 631.050 ;
        RECT 199.950 629.400 295.050 630.600 ;
        RECT 199.950 628.800 202.050 629.400 ;
        RECT 292.950 628.950 295.050 629.400 ;
        RECT 319.950 630.600 322.050 631.050 ;
        RECT 367.950 630.600 370.050 631.050 ;
        RECT 319.950 629.400 370.050 630.600 ;
        RECT 319.950 628.950 322.050 629.400 ;
        RECT 367.950 628.950 370.050 629.400 ;
        RECT 517.950 630.600 520.050 631.050 ;
        RECT 529.950 630.600 532.050 631.050 ;
        RECT 571.950 630.600 574.050 631.050 ;
        RECT 769.950 630.600 772.050 631.050 ;
        RECT 517.950 629.400 574.050 630.600 ;
        RECT 517.950 628.950 520.050 629.400 ;
        RECT 529.950 628.950 532.050 629.400 ;
        RECT 571.950 628.950 574.050 629.400 ;
        RECT 620.400 629.400 772.050 630.600 ;
        RECT 190.950 627.600 193.050 628.050 ;
        RECT 202.950 627.600 205.050 628.050 ;
        RECT 190.950 626.400 205.050 627.600 ;
        RECT 190.950 625.950 193.050 626.400 ;
        RECT 202.950 625.950 205.050 626.400 ;
        RECT 229.950 627.600 232.050 628.050 ;
        RECT 262.950 627.600 265.050 628.050 ;
        RECT 229.950 626.400 265.050 627.600 ;
        RECT 229.950 625.950 232.050 626.400 ;
        RECT 262.950 625.950 265.050 626.400 ;
        RECT 268.950 627.600 271.050 628.050 ;
        RECT 304.950 627.600 307.050 628.050 ;
        RECT 268.950 626.400 307.050 627.600 ;
        RECT 268.950 625.950 271.050 626.400 ;
        RECT 304.950 625.950 307.050 626.400 ;
        RECT 382.950 627.600 385.050 628.050 ;
        RECT 400.950 627.600 403.050 628.050 ;
        RECT 499.950 627.600 502.050 628.050 ;
        RECT 382.950 626.400 393.600 627.600 ;
        RECT 382.950 625.950 385.050 626.400 ;
        RECT 392.400 625.050 393.600 626.400 ;
        RECT 400.950 626.400 502.050 627.600 ;
        RECT 400.950 625.950 403.050 626.400 ;
        RECT 499.950 625.950 502.050 626.400 ;
        RECT 529.950 627.600 532.050 627.900 ;
        RECT 541.950 627.600 544.050 628.050 ;
        RECT 529.950 626.400 544.050 627.600 ;
        RECT 529.950 625.800 532.050 626.400 ;
        RECT 541.950 625.950 544.050 626.400 ;
        RECT 580.950 627.600 583.050 628.050 ;
        RECT 595.950 627.600 598.050 628.050 ;
        RECT 620.400 627.600 621.600 629.400 ;
        RECT 769.950 628.950 772.050 629.400 ;
        RECT 580.950 626.400 594.600 627.600 ;
        RECT 580.950 625.950 583.050 626.400 ;
        RECT 160.950 624.600 163.050 625.050 ;
        RECT 274.950 624.600 277.050 625.050 ;
        RECT 160.950 623.400 277.050 624.600 ;
        RECT 160.950 622.950 163.050 623.400 ;
        RECT 274.950 622.950 277.050 623.400 ;
        RECT 316.950 624.600 319.050 625.050 ;
        RECT 331.950 624.600 334.050 625.050 ;
        RECT 316.950 623.400 334.050 624.600 ;
        RECT 316.950 622.950 319.050 623.400 ;
        RECT 331.950 622.950 334.050 623.400 ;
        RECT 349.950 624.600 352.050 625.050 ;
        RECT 379.950 624.600 382.050 625.050 ;
        RECT 349.950 623.400 382.050 624.600 ;
        RECT 349.950 622.950 352.050 623.400 ;
        RECT 379.950 622.950 382.050 623.400 ;
        RECT 391.950 624.600 394.050 625.050 ;
        RECT 436.950 624.600 439.050 625.050 ;
        RECT 391.950 623.400 439.050 624.600 ;
        RECT 391.950 622.950 394.050 623.400 ;
        RECT 436.950 622.950 439.050 623.400 ;
        RECT 550.950 624.600 553.050 625.050 ;
        RECT 577.950 624.600 580.050 625.050 ;
        RECT 550.950 623.400 580.050 624.600 ;
        RECT 593.400 624.600 594.600 626.400 ;
        RECT 595.950 626.400 621.600 627.600 ;
        RECT 802.950 627.600 805.050 628.050 ;
        RECT 838.950 627.600 841.050 628.050 ;
        RECT 853.950 627.600 856.050 628.050 ;
        RECT 802.950 626.400 856.050 627.600 ;
        RECT 595.950 625.950 598.050 626.400 ;
        RECT 802.950 625.950 805.050 626.400 ;
        RECT 838.950 625.950 841.050 626.400 ;
        RECT 853.950 625.950 856.050 626.400 ;
        RECT 598.950 624.600 601.050 625.050 ;
        RECT 613.950 624.600 616.050 625.050 ;
        RECT 593.400 623.400 616.050 624.600 ;
        RECT 550.950 622.950 553.050 623.400 ;
        RECT 577.950 622.950 580.050 623.400 ;
        RECT 598.950 622.950 601.050 623.400 ;
        RECT 613.950 622.950 616.050 623.400 ;
        RECT 628.950 624.600 631.050 625.050 ;
        RECT 649.950 624.600 652.050 625.050 ;
        RECT 628.950 623.400 652.050 624.600 ;
        RECT 628.950 622.950 631.050 623.400 ;
        RECT 649.950 622.950 652.050 623.400 ;
        RECT 25.950 621.600 28.050 622.050 ;
        RECT 70.950 621.600 73.050 622.050 ;
        RECT 25.950 620.400 73.050 621.600 ;
        RECT 25.950 619.950 28.050 620.400 ;
        RECT 70.950 619.950 73.050 620.400 ;
        RECT 103.950 621.600 106.050 622.050 ;
        RECT 127.950 621.600 130.050 622.050 ;
        RECT 103.950 620.400 130.050 621.600 ;
        RECT 103.950 619.950 106.050 620.400 ;
        RECT 127.950 619.950 130.050 620.400 ;
        RECT 169.950 621.600 172.050 622.050 ;
        RECT 208.950 621.600 211.050 622.050 ;
        RECT 241.950 621.600 244.050 622.050 ;
        RECT 169.950 620.400 211.050 621.600 ;
        RECT 169.950 619.950 172.050 620.400 ;
        RECT 208.950 619.950 211.050 620.400 ;
        RECT 218.400 620.400 244.050 621.600 ;
        RECT 1.950 618.600 4.050 619.050 ;
        RECT 91.950 618.600 94.050 619.050 ;
        RECT 1.950 617.400 94.050 618.600 ;
        RECT 1.950 616.950 4.050 617.400 ;
        RECT 91.950 616.950 94.050 617.400 ;
        RECT 106.950 618.600 109.050 619.050 ;
        RECT 121.950 618.600 124.050 619.050 ;
        RECT 136.950 618.600 139.050 619.050 ;
        RECT 106.950 617.400 139.050 618.600 ;
        RECT 106.950 616.950 109.050 617.400 ;
        RECT 121.950 616.950 124.050 617.400 ;
        RECT 136.950 616.950 139.050 617.400 ;
        RECT 154.950 618.600 157.050 619.050 ;
        RECT 172.950 618.600 175.050 619.050 ;
        RECT 154.950 617.400 175.050 618.600 ;
        RECT 154.950 616.950 157.050 617.400 ;
        RECT 172.950 616.950 175.050 617.400 ;
        RECT 193.950 618.600 196.050 619.050 ;
        RECT 218.400 618.600 219.600 620.400 ;
        RECT 241.950 619.950 244.050 620.400 ;
        RECT 274.950 621.600 277.050 621.900 ;
        RECT 289.800 621.600 291.900 622.050 ;
        RECT 274.950 620.400 291.900 621.600 ;
        RECT 274.950 619.800 277.050 620.400 ;
        RECT 289.800 619.950 291.900 620.400 ;
        RECT 292.950 621.600 295.050 622.050 ;
        RECT 307.950 621.600 310.050 622.050 ;
        RECT 346.950 621.600 349.050 622.050 ;
        RECT 292.950 620.400 306.600 621.600 ;
        RECT 292.950 619.950 295.050 620.400 ;
        RECT 193.950 617.400 219.600 618.600 ;
        RECT 238.950 618.600 241.050 619.050 ;
        RECT 265.950 618.600 268.050 619.050 ;
        RECT 238.950 617.400 268.050 618.600 ;
        RECT 305.400 618.600 306.600 620.400 ;
        RECT 307.950 620.400 349.050 621.600 ;
        RECT 307.950 619.950 310.050 620.400 ;
        RECT 346.950 619.950 349.050 620.400 ;
        RECT 355.950 621.600 358.050 622.050 ;
        RECT 376.950 621.600 379.050 622.050 ;
        RECT 355.950 620.400 379.050 621.600 ;
        RECT 355.950 619.950 358.050 620.400 ;
        RECT 376.950 619.950 379.050 620.400 ;
        RECT 397.950 621.600 400.050 622.050 ;
        RECT 439.950 621.600 442.050 622.050 ;
        RECT 397.950 620.400 442.050 621.600 ;
        RECT 397.950 619.950 400.050 620.400 ;
        RECT 439.950 619.950 442.050 620.400 ;
        RECT 526.950 621.600 529.050 622.050 ;
        RECT 544.950 621.600 547.050 622.050 ;
        RECT 751.950 621.600 754.050 622.050 ;
        RECT 772.950 621.600 775.050 622.050 ;
        RECT 526.950 620.400 549.600 621.600 ;
        RECT 526.950 619.950 529.050 620.400 ;
        RECT 544.950 619.950 547.050 620.400 ;
        RECT 322.950 618.600 325.050 619.050 ;
        RECT 305.400 617.400 325.050 618.600 ;
        RECT 193.950 616.950 196.050 617.400 ;
        RECT 238.950 616.950 241.050 617.400 ;
        RECT 265.950 616.950 268.050 617.400 ;
        RECT 322.950 616.950 325.050 617.400 ;
        RECT 382.950 618.600 385.050 619.050 ;
        RECT 475.950 618.600 478.050 619.050 ;
        RECT 487.950 618.600 490.050 619.050 ;
        RECT 532.950 618.600 535.050 619.050 ;
        RECT 382.950 617.400 490.050 618.600 ;
        RECT 382.950 616.950 385.050 617.400 ;
        RECT 475.950 616.950 478.050 617.400 ;
        RECT 487.950 616.950 490.050 617.400 ;
        RECT 491.400 617.400 516.600 618.600 ;
        RECT 130.950 615.600 133.050 616.050 ;
        RECT 169.950 615.600 172.050 616.050 ;
        RECT 130.950 614.400 172.050 615.600 ;
        RECT 130.950 613.950 133.050 614.400 ;
        RECT 169.950 613.950 172.050 614.400 ;
        RECT 187.950 615.600 190.050 616.050 ;
        RECT 223.950 615.600 226.050 616.050 ;
        RECT 187.950 614.400 226.050 615.600 ;
        RECT 187.950 613.950 190.050 614.400 ;
        RECT 223.950 613.950 226.050 614.400 ;
        RECT 250.950 615.600 253.050 616.050 ;
        RECT 286.950 615.600 289.050 616.050 ;
        RECT 250.950 614.400 289.050 615.600 ;
        RECT 250.950 613.950 253.050 614.400 ;
        RECT 286.950 613.950 289.050 614.400 ;
        RECT 301.950 615.600 304.050 616.050 ;
        RECT 349.950 615.600 352.050 616.050 ;
        RECT 301.950 614.400 352.050 615.600 ;
        RECT 301.950 613.950 304.050 614.400 ;
        RECT 349.950 613.950 352.050 614.400 ;
        RECT 358.950 615.600 361.050 616.050 ;
        RECT 376.950 615.600 379.050 616.050 ;
        RECT 358.950 614.400 379.050 615.600 ;
        RECT 358.950 613.950 361.050 614.400 ;
        RECT 376.950 613.950 379.050 614.400 ;
        RECT 391.950 615.600 394.050 616.050 ;
        RECT 491.400 615.600 492.600 617.400 ;
        RECT 391.950 614.400 492.600 615.600 ;
        RECT 515.400 615.600 516.600 617.400 ;
        RECT 521.400 617.400 535.050 618.600 ;
        RECT 521.400 615.600 522.600 617.400 ;
        RECT 532.950 616.950 535.050 617.400 ;
        RECT 538.950 618.600 541.050 619.050 ;
        RECT 544.950 618.600 547.050 618.900 ;
        RECT 538.950 617.400 547.050 618.600 ;
        RECT 548.400 618.600 549.600 620.400 ;
        RECT 751.950 620.400 775.050 621.600 ;
        RECT 751.950 619.950 754.050 620.400 ;
        RECT 772.950 619.950 775.050 620.400 ;
        RECT 784.950 621.600 787.050 622.050 ;
        RECT 832.950 621.600 835.050 622.050 ;
        RECT 784.950 620.400 835.050 621.600 ;
        RECT 784.950 619.950 787.050 620.400 ;
        RECT 832.950 619.950 835.050 620.400 ;
        RECT 559.800 618.600 561.900 619.050 ;
        RECT 548.400 617.400 561.900 618.600 ;
        RECT 538.950 616.950 541.050 617.400 ;
        RECT 544.950 616.800 547.050 617.400 ;
        RECT 559.800 616.950 561.900 617.400 ;
        RECT 562.950 618.600 565.050 619.050 ;
        RECT 619.950 618.600 622.050 619.050 ;
        RECT 664.950 618.600 667.050 619.050 ;
        RECT 679.950 618.600 682.050 619.050 ;
        RECT 691.950 618.600 694.050 619.050 ;
        RECT 562.950 617.400 582.600 618.600 ;
        RECT 562.950 616.950 565.050 617.400 ;
        RECT 515.400 614.400 522.600 615.600 ;
        RECT 535.950 615.600 538.050 616.050 ;
        RECT 562.950 615.600 565.050 615.900 ;
        RECT 535.950 614.400 565.050 615.600 ;
        RECT 581.400 615.600 582.600 617.400 ;
        RECT 619.950 617.400 694.050 618.600 ;
        RECT 619.950 616.950 622.050 617.400 ;
        RECT 664.950 616.950 667.050 617.400 ;
        RECT 679.950 616.950 682.050 617.400 ;
        RECT 691.950 616.950 694.050 617.400 ;
        RECT 697.950 618.600 700.050 619.050 ;
        RECT 712.950 618.600 715.050 619.050 ;
        RECT 697.950 617.400 715.050 618.600 ;
        RECT 697.950 616.950 700.050 617.400 ;
        RECT 712.950 616.950 715.050 617.400 ;
        RECT 607.950 615.600 610.050 616.050 ;
        RECT 751.950 615.600 754.050 616.050 ;
        RECT 581.400 614.400 610.050 615.600 ;
        RECT 391.950 613.950 394.050 614.400 ;
        RECT 535.950 613.950 538.050 614.400 ;
        RECT 562.950 613.800 565.050 614.400 ;
        RECT 607.950 613.950 610.050 614.400 ;
        RECT 614.400 614.400 754.050 615.600 ;
        RECT 76.950 612.600 79.050 613.050 ;
        RECT 82.950 612.600 85.050 613.050 ;
        RECT 76.950 611.400 85.050 612.600 ;
        RECT 76.950 610.950 79.050 611.400 ;
        RECT 82.950 610.950 85.050 611.400 ;
        RECT 109.950 612.600 112.050 613.050 ;
        RECT 163.950 612.600 166.050 613.050 ;
        RECT 109.950 611.400 166.050 612.600 ;
        RECT 109.950 610.950 112.050 611.400 ;
        RECT 163.950 610.950 166.050 611.400 ;
        RECT 19.950 609.600 22.050 610.050 ;
        RECT 28.950 609.600 31.050 610.050 ;
        RECT 17.400 608.400 31.050 609.600 ;
        RECT 17.400 600.750 18.600 608.400 ;
        RECT 19.950 607.950 22.050 608.400 ;
        RECT 28.950 607.950 31.050 608.400 ;
        RECT 55.950 609.600 58.050 610.050 ;
        RECT 77.400 609.600 78.600 610.950 ;
        RECT 55.950 608.400 78.600 609.600 ;
        RECT 85.950 609.600 88.050 609.900 ;
        RECT 91.950 609.600 94.050 610.050 ;
        RECT 85.950 608.400 94.050 609.600 ;
        RECT 55.950 607.950 58.050 608.400 ;
        RECT 85.950 607.800 88.050 608.400 ;
        RECT 91.950 607.950 94.050 608.400 ;
        RECT 148.950 609.600 151.050 610.050 ;
        RECT 160.950 609.600 163.050 610.050 ;
        RECT 148.950 608.400 163.050 609.600 ;
        RECT 148.950 607.950 151.050 608.400 ;
        RECT 160.950 607.950 163.050 608.400 ;
        RECT 166.950 609.600 169.050 610.050 ;
        RECT 196.950 609.600 199.050 610.050 ;
        RECT 208.950 609.600 211.050 610.050 ;
        RECT 166.950 608.400 211.050 609.600 ;
        RECT 166.950 607.950 169.050 608.400 ;
        RECT 196.950 607.950 199.050 608.400 ;
        RECT 208.950 607.950 211.050 608.400 ;
        RECT 244.950 609.600 247.050 610.050 ;
        RECT 250.950 609.600 253.050 610.050 ;
        RECT 244.950 608.400 253.050 609.600 ;
        RECT 244.950 607.950 247.050 608.400 ;
        RECT 250.950 607.950 253.050 608.400 ;
        RECT 256.950 609.600 259.050 610.050 ;
        RECT 277.950 609.600 280.050 613.050 ;
        RECT 328.950 612.600 331.050 613.050 ;
        RECT 346.950 612.600 349.050 613.050 ;
        RECT 328.950 611.400 349.050 612.600 ;
        RECT 328.950 610.950 331.050 611.400 ;
        RECT 346.950 610.950 349.050 611.400 ;
        RECT 355.950 612.600 358.050 613.050 ;
        RECT 385.950 612.600 388.050 613.050 ;
        RECT 355.950 611.400 388.050 612.600 ;
        RECT 355.950 610.950 358.050 611.400 ;
        RECT 385.950 610.950 388.050 611.400 ;
        RECT 436.950 612.600 439.050 613.050 ;
        RECT 442.950 612.600 445.050 613.050 ;
        RECT 436.950 611.400 445.050 612.600 ;
        RECT 436.950 610.950 439.050 611.400 ;
        RECT 442.950 610.950 445.050 611.400 ;
        RECT 469.950 612.600 472.050 613.050 ;
        RECT 511.950 612.600 514.050 613.050 ;
        RECT 469.950 611.400 514.050 612.600 ;
        RECT 469.950 610.950 472.050 611.400 ;
        RECT 511.950 610.950 514.050 611.400 ;
        RECT 256.950 609.000 280.050 609.600 ;
        RECT 322.950 609.600 325.050 610.050 ;
        RECT 352.950 609.600 355.050 610.050 ;
        RECT 256.950 608.400 279.600 609.000 ;
        RECT 322.950 608.400 355.050 609.600 ;
        RECT 256.950 607.950 259.050 608.400 ;
        RECT 322.950 607.950 325.050 608.400 ;
        RECT 19.950 604.800 22.050 606.900 ;
        RECT 34.950 606.600 37.050 607.050 ;
        RECT 43.950 606.600 46.050 607.050 ;
        RECT 51.000 606.600 55.050 607.050 ;
        RECT 34.950 605.400 46.050 606.600 ;
        RECT 34.950 604.950 37.050 605.400 ;
        RECT 43.950 604.950 46.050 605.400 ;
        RECT 50.400 604.950 55.050 606.600 ;
        RECT 58.950 604.950 61.050 607.050 ;
        RECT 79.950 606.600 82.050 607.050 ;
        RECT 65.400 605.400 82.050 606.600 ;
        RECT 16.950 598.650 19.050 600.750 ;
        RECT 20.400 600.600 21.600 604.800 ;
        RECT 50.400 601.050 51.600 604.950 ;
        RECT 31.950 600.600 34.050 600.750 ;
        RECT 20.400 599.400 34.050 600.600 ;
        RECT 31.950 598.650 34.050 599.400 ;
        RECT 49.950 598.950 52.050 601.050 ;
        RECT 59.400 600.750 60.600 604.950 ;
        RECT 65.400 601.050 66.600 605.400 ;
        RECT 79.950 604.950 82.050 605.400 ;
        RECT 94.950 603.600 97.050 607.050 ;
        RECT 100.950 606.600 103.050 607.050 ;
        RECT 106.950 606.600 109.050 607.050 ;
        RECT 126.000 606.600 130.050 607.050 ;
        RECT 100.950 605.400 109.050 606.600 ;
        RECT 100.950 604.950 103.050 605.400 ;
        RECT 106.950 604.950 109.050 605.400 ;
        RECT 125.400 604.950 130.050 606.600 ;
        RECT 142.950 604.950 145.050 607.050 ;
        RECT 163.950 604.950 166.050 607.050 ;
        RECT 199.950 606.600 202.050 607.050 ;
        RECT 191.400 605.400 202.050 606.600 ;
        RECT 109.950 603.600 112.050 604.050 ;
        RECT 94.950 603.000 112.050 603.600 ;
        RECT 95.400 602.400 112.050 603.000 ;
        RECT 109.950 601.950 112.050 602.400 ;
        RECT 58.950 598.650 61.050 600.750 ;
        RECT 64.950 598.950 67.050 601.050 ;
        RECT 125.400 600.900 126.600 604.950 ;
        RECT 124.950 600.600 127.050 600.900 ;
        RECT 133.950 600.600 136.050 600.900 ;
        RECT 124.950 599.400 136.050 600.600 ;
        RECT 124.950 598.800 127.050 599.400 ;
        RECT 133.950 598.800 136.050 599.400 ;
        RECT 143.400 598.050 144.600 604.950 ;
        RECT 164.400 600.600 165.600 604.950 ;
        RECT 191.400 601.050 192.600 605.400 ;
        RECT 199.950 604.950 202.050 605.400 ;
        RECT 214.950 606.600 217.050 607.050 ;
        RECT 232.950 606.600 235.050 607.200 ;
        RECT 214.950 605.400 235.050 606.600 ;
        RECT 214.950 604.950 217.050 605.400 ;
        RECT 232.950 605.100 235.050 605.400 ;
        RECT 247.950 603.600 250.050 607.050 ;
        RECT 268.950 605.100 271.050 607.200 ;
        RECT 292.950 606.600 295.050 607.050 ;
        RECT 292.950 605.400 315.600 606.600 ;
        RECT 247.950 603.000 255.600 603.600 ;
        RECT 248.400 602.400 255.600 603.000 ;
        RECT 181.950 600.600 184.050 600.750 ;
        RECT 164.400 599.400 184.050 600.600 ;
        RECT 181.950 598.650 184.050 599.400 ;
        RECT 190.950 598.950 193.050 601.050 ;
        RECT 217.950 600.600 220.050 600.750 ;
        RECT 244.950 600.600 247.050 601.050 ;
        RECT 254.400 600.750 255.600 602.400 ;
        RECT 217.950 599.400 247.050 600.600 ;
        RECT 217.950 598.650 220.050 599.400 ;
        RECT 244.950 598.950 247.050 599.400 ;
        RECT 253.950 598.650 256.050 600.750 ;
        RECT 259.950 600.600 262.050 601.050 ;
        RECT 269.400 600.600 270.600 605.100 ;
        RECT 292.950 604.950 295.050 605.400 ;
        RECT 314.400 600.900 315.600 605.400 ;
        RECT 259.950 599.400 270.600 600.600 ;
        RECT 289.950 600.300 292.050 600.750 ;
        RECT 304.950 600.300 307.050 600.750 ;
        RECT 259.950 598.950 262.050 599.400 ;
        RECT 289.950 599.100 307.050 600.300 ;
        RECT 289.950 598.650 292.050 599.100 ;
        RECT 304.950 598.650 307.050 599.100 ;
        RECT 313.950 598.800 316.050 600.900 ;
        RECT 322.950 600.600 325.050 601.050 ;
        RECT 332.400 600.600 333.600 608.400 ;
        RECT 352.950 607.950 355.050 608.400 ;
        RECT 388.950 609.600 391.050 610.050 ;
        RECT 394.950 609.600 397.050 610.050 ;
        RECT 388.950 608.400 397.050 609.600 ;
        RECT 388.950 607.950 391.050 608.400 ;
        RECT 394.950 607.950 397.050 608.400 ;
        RECT 412.950 609.600 415.050 610.050 ;
        RECT 412.950 608.400 420.600 609.600 ;
        RECT 412.950 607.950 415.050 608.400 ;
        RECT 334.950 604.950 337.050 607.050 ;
        RECT 322.950 599.400 333.600 600.600 ;
        RECT 335.400 600.600 336.600 604.950 ;
        RECT 340.950 603.600 343.050 607.050 ;
        RECT 358.950 606.750 361.050 607.200 ;
        RECT 367.950 606.750 370.050 607.200 ;
        RECT 358.950 605.550 370.050 606.750 ;
        RECT 358.950 605.100 361.050 605.550 ;
        RECT 367.950 605.100 370.050 605.550 ;
        RECT 382.950 603.600 385.050 607.050 ;
        RECT 400.950 606.600 403.050 607.200 ;
        RECT 400.950 605.400 417.600 606.600 ;
        RECT 400.950 605.100 403.050 605.400 ;
        RECT 340.950 603.000 345.600 603.600 ;
        RECT 382.950 603.000 390.600 603.600 ;
        RECT 341.400 602.400 345.600 603.000 ;
        RECT 383.400 602.400 390.600 603.000 ;
        RECT 344.400 600.600 345.600 602.400 ;
        RECT 385.950 600.600 388.050 601.050 ;
        RECT 335.400 599.400 342.600 600.600 ;
        RECT 344.400 599.400 388.050 600.600 ;
        RECT 389.400 600.600 390.600 602.400 ;
        RECT 389.400 600.000 414.600 600.600 ;
        RECT 389.400 599.400 415.050 600.000 ;
        RECT 322.950 598.950 325.050 599.400 ;
        RECT 31.950 597.600 34.050 598.050 ;
        RECT 52.950 597.600 55.050 598.050 ;
        RECT 31.950 596.400 55.050 597.600 ;
        RECT 31.950 595.950 34.050 596.400 ;
        RECT 52.950 595.950 55.050 596.400 ;
        RECT 58.950 597.600 61.050 598.050 ;
        RECT 73.950 597.600 76.050 598.050 ;
        RECT 58.950 596.400 76.050 597.600 ;
        RECT 58.950 595.950 61.050 596.400 ;
        RECT 73.950 595.950 76.050 596.400 ;
        RECT 94.950 597.600 97.050 598.050 ;
        RECT 106.950 597.600 109.050 598.050 ;
        RECT 115.950 597.600 118.050 598.050 ;
        RECT 94.950 596.400 118.050 597.600 ;
        RECT 94.950 595.950 97.050 596.400 ;
        RECT 106.950 595.950 109.050 596.400 ;
        RECT 115.950 595.950 118.050 596.400 ;
        RECT 142.950 595.950 145.050 598.050 ;
        RECT 331.950 597.600 334.050 598.050 ;
        RECT 337.950 597.600 340.050 598.050 ;
        RECT 331.950 596.400 340.050 597.600 ;
        RECT 341.400 597.600 342.600 599.400 ;
        RECT 385.950 598.950 388.050 599.400 ;
        RECT 355.950 597.600 358.050 598.050 ;
        RECT 341.400 596.400 358.050 597.600 ;
        RECT 331.950 595.950 334.050 596.400 ;
        RECT 337.950 595.950 340.050 596.400 ;
        RECT 355.950 595.950 358.050 596.400 ;
        RECT 403.950 597.600 406.050 598.050 ;
        RECT 409.800 597.600 411.900 598.050 ;
        RECT 403.950 596.400 411.900 597.600 ;
        RECT 403.950 595.950 406.050 596.400 ;
        RECT 409.800 595.950 411.900 596.400 ;
        RECT 412.950 595.950 415.050 599.400 ;
        RECT 100.950 594.600 103.050 595.050 ;
        RECT 145.950 594.600 148.050 595.050 ;
        RECT 178.950 594.600 181.050 595.050 ;
        RECT 100.950 593.400 114.600 594.600 ;
        RECT 100.950 592.950 103.050 593.400 ;
        RECT 113.400 591.600 114.600 593.400 ;
        RECT 145.950 593.400 181.050 594.600 ;
        RECT 145.950 592.950 148.050 593.400 ;
        RECT 178.950 592.950 181.050 593.400 ;
        RECT 319.950 594.600 322.050 595.050 ;
        RECT 397.950 594.600 400.050 595.050 ;
        RECT 416.400 594.600 417.600 605.400 ;
        RECT 419.400 598.050 420.600 608.400 ;
        RECT 529.950 607.950 532.050 610.050 ;
        RECT 532.950 609.600 535.050 613.050 ;
        RECT 544.950 612.600 547.050 613.050 ;
        RECT 556.950 612.600 559.050 613.050 ;
        RECT 544.950 611.400 559.050 612.600 ;
        RECT 544.950 610.950 547.050 611.400 ;
        RECT 556.950 610.950 559.050 611.400 ;
        RECT 580.950 612.600 583.050 613.050 ;
        RECT 614.400 612.600 615.600 614.400 ;
        RECT 751.950 613.950 754.050 614.400 ;
        RECT 763.950 615.600 766.050 616.050 ;
        RECT 790.950 615.600 793.050 616.050 ;
        RECT 763.950 614.400 793.050 615.600 ;
        RECT 763.950 613.950 766.050 614.400 ;
        RECT 790.950 613.950 793.050 614.400 ;
        RECT 580.950 611.400 615.600 612.600 ;
        RECT 673.950 612.600 676.050 613.050 ;
        RECT 685.950 612.600 688.050 613.050 ;
        RECT 673.950 611.400 688.050 612.600 ;
        RECT 580.950 610.950 583.050 611.400 ;
        RECT 673.950 610.950 676.050 611.400 ;
        RECT 685.950 610.950 688.050 611.400 ;
        RECT 805.950 612.600 808.050 613.050 ;
        RECT 823.950 612.600 826.050 613.050 ;
        RECT 805.950 611.400 826.050 612.600 ;
        RECT 805.950 610.950 808.050 611.400 ;
        RECT 823.950 610.950 826.050 611.400 ;
        RECT 571.950 609.600 574.050 610.050 ;
        RECT 595.950 609.600 598.050 610.050 ;
        RECT 532.950 609.000 537.600 609.600 ;
        RECT 533.400 608.400 537.600 609.000 ;
        RECT 439.950 606.600 442.050 607.050 ;
        RECT 460.950 606.600 463.050 607.050 ;
        RECT 439.950 605.400 447.600 606.600 ;
        RECT 439.950 604.950 442.050 605.400 ;
        RECT 446.400 601.050 447.600 605.400 ;
        RECT 452.400 605.400 463.050 606.600 ;
        RECT 452.400 601.050 453.600 605.400 ;
        RECT 460.950 604.950 463.050 605.400 ;
        RECT 466.950 604.950 469.050 607.050 ;
        RECT 481.950 606.600 484.050 607.050 ;
        RECT 499.950 606.600 502.050 606.900 ;
        RECT 523.950 606.600 526.050 607.050 ;
        RECT 481.950 605.400 502.050 606.600 ;
        RECT 481.950 604.950 484.050 605.400 ;
        RECT 445.950 598.950 448.050 601.050 ;
        RECT 451.950 598.950 454.050 601.050 ;
        RECT 457.950 600.600 460.050 600.900 ;
        RECT 467.400 600.600 468.600 604.950 ;
        RECT 499.950 603.600 502.050 605.400 ;
        RECT 515.400 605.400 526.050 606.600 ;
        RECT 499.950 603.000 510.600 603.600 ;
        RECT 500.400 602.400 511.050 603.000 ;
        RECT 457.950 599.400 468.600 600.600 ;
        RECT 469.950 600.600 472.050 601.050 ;
        RECT 478.950 600.600 481.050 600.750 ;
        RECT 469.950 599.400 481.050 600.600 ;
        RECT 457.950 598.800 460.050 599.400 ;
        RECT 469.950 598.950 472.050 599.400 ;
        RECT 478.950 598.650 481.050 599.400 ;
        RECT 508.950 598.950 511.050 602.400 ;
        RECT 515.400 600.900 516.600 605.400 ;
        RECT 523.950 604.950 526.050 605.400 ;
        RECT 514.950 598.800 517.050 600.900 ;
        RECT 530.400 600.600 531.600 607.950 ;
        RECT 536.400 606.600 537.600 608.400 ;
        RECT 571.950 608.400 598.050 609.600 ;
        RECT 571.950 607.950 574.050 608.400 ;
        RECT 595.950 607.950 598.050 608.400 ;
        RECT 697.950 609.600 700.050 610.050 ;
        RECT 718.950 609.600 721.050 610.050 ;
        RECT 697.950 608.400 721.050 609.600 ;
        RECT 697.950 607.950 700.050 608.400 ;
        RECT 718.950 607.950 721.050 608.400 ;
        RECT 742.950 609.600 745.050 610.050 ;
        RECT 760.950 609.600 763.050 610.050 ;
        RECT 742.950 608.400 763.050 609.600 ;
        RECT 742.950 607.950 745.050 608.400 ;
        RECT 760.950 607.950 763.050 608.400 ;
        RECT 796.950 609.600 799.050 610.050 ;
        RECT 811.950 609.600 814.050 610.050 ;
        RECT 856.950 609.600 859.050 610.050 ;
        RECT 862.950 609.600 865.050 610.050 ;
        RECT 796.950 608.400 816.600 609.600 ;
        RECT 796.950 607.950 799.050 608.400 ;
        RECT 811.950 607.950 814.050 608.400 ;
        RECT 574.950 606.600 577.050 607.050 ;
        RECT 536.400 605.400 540.600 606.600 ;
        RECT 539.400 600.600 540.600 605.400 ;
        RECT 574.950 605.400 594.600 606.600 ;
        RECT 574.950 604.950 577.050 605.400 ;
        RECT 593.400 604.050 594.600 605.400 ;
        RECT 598.950 604.950 601.050 607.050 ;
        RECT 607.950 606.600 610.050 607.050 ;
        RECT 607.950 605.400 615.600 606.600 ;
        RECT 607.950 604.950 610.050 605.400 ;
        RECT 593.400 602.400 598.050 604.050 ;
        RECT 594.000 601.950 598.050 602.400 ;
        RECT 547.950 600.600 550.050 601.050 ;
        RECT 599.400 600.600 600.600 604.950 ;
        RECT 614.400 601.050 615.600 605.400 ;
        RECT 619.950 604.950 622.050 607.050 ;
        RECT 628.950 606.750 631.050 607.200 ;
        RECT 637.950 606.750 640.050 607.200 ;
        RECT 628.950 605.550 640.050 606.750 ;
        RECT 628.950 605.100 631.050 605.550 ;
        RECT 637.950 605.100 640.050 605.550 ;
        RECT 643.950 605.100 646.050 607.200 ;
        RECT 652.950 606.750 655.050 607.200 ;
        RECT 658.950 606.750 661.050 607.200 ;
        RECT 652.950 605.550 661.050 606.750 ;
        RECT 652.950 605.100 655.050 605.550 ;
        RECT 658.950 605.100 661.050 605.550 ;
        RECT 530.400 600.000 534.600 600.600 ;
        RECT 530.400 599.400 535.050 600.000 ;
        RECT 539.400 599.400 550.050 600.600 ;
        RECT 418.950 595.950 421.050 598.050 ;
        RECT 532.950 595.950 535.050 599.400 ;
        RECT 547.950 598.950 550.050 599.400 ;
        RECT 587.400 599.400 600.600 600.600 ;
        RECT 556.950 597.600 559.050 598.050 ;
        RECT 571.950 597.600 574.050 598.050 ;
        RECT 556.950 596.400 574.050 597.600 ;
        RECT 556.950 595.950 559.050 596.400 ;
        RECT 571.950 595.950 574.050 596.400 ;
        RECT 580.950 597.600 583.050 598.050 ;
        RECT 587.400 597.600 588.600 599.400 ;
        RECT 613.950 598.950 616.050 601.050 ;
        RECT 580.950 596.400 588.600 597.600 ;
        RECT 604.950 597.600 607.050 598.050 ;
        RECT 620.400 597.600 621.600 604.950 ;
        RECT 644.400 600.600 645.600 605.100 ;
        RECT 673.950 604.950 676.050 607.050 ;
        RECT 703.950 606.600 706.050 607.050 ;
        RECT 724.950 606.600 727.050 607.050 ;
        RECT 733.950 606.600 736.050 607.050 ;
        RECT 703.950 605.400 736.050 606.600 ;
        RECT 703.950 604.950 706.050 605.400 ;
        RECT 724.950 604.950 727.050 605.400 ;
        RECT 733.950 604.950 736.050 605.400 ;
        RECT 778.950 604.950 781.050 607.050 ;
        RECT 674.400 601.050 675.600 604.950 ;
        RECT 661.950 600.600 664.050 600.900 ;
        RECT 644.400 599.400 664.050 600.600 ;
        RECT 661.950 598.800 664.050 599.400 ;
        RECT 673.950 598.950 676.050 601.050 ;
        RECT 700.950 600.300 703.050 600.750 ;
        RECT 712.950 600.300 715.050 600.750 ;
        RECT 700.950 599.100 715.050 600.300 ;
        RECT 779.400 600.600 780.600 604.950 ;
        RECT 815.400 603.600 816.600 608.400 ;
        RECT 856.950 608.400 865.050 609.600 ;
        RECT 856.950 607.950 859.050 608.400 ;
        RECT 862.950 607.950 865.050 608.400 ;
        RECT 832.950 605.100 835.050 607.200 ;
        RECT 815.400 603.000 822.600 603.600 ;
        RECT 815.400 602.400 823.050 603.000 ;
        RECT 799.950 600.600 802.050 600.750 ;
        RECT 779.400 599.400 802.050 600.600 ;
        RECT 700.950 598.650 703.050 599.100 ;
        RECT 712.950 598.650 715.050 599.100 ;
        RECT 799.950 598.650 802.050 599.400 ;
        RECT 820.950 598.950 823.050 602.400 ;
        RECT 604.950 596.400 621.600 597.600 ;
        RECT 640.950 597.600 643.050 598.050 ;
        RECT 655.950 597.600 658.050 598.050 ;
        RECT 640.950 596.400 658.050 597.600 ;
        RECT 580.950 595.950 583.050 596.400 ;
        RECT 604.950 595.950 607.050 596.400 ;
        RECT 640.950 595.950 643.050 596.400 ;
        RECT 655.950 595.950 658.050 596.400 ;
        RECT 685.950 597.600 688.050 598.050 ;
        RECT 691.950 597.600 694.050 598.050 ;
        RECT 685.950 596.400 694.050 597.600 ;
        RECT 713.400 597.600 714.600 598.650 ;
        RECT 833.400 598.050 834.600 605.100 ;
        RECT 838.950 604.950 841.050 607.050 ;
        RECT 839.400 601.050 840.600 604.950 ;
        RECT 838.950 598.950 841.050 601.050 ;
        RECT 721.950 597.600 724.050 598.050 ;
        RECT 713.400 596.400 724.050 597.600 ;
        RECT 685.950 595.950 688.050 596.400 ;
        RECT 691.950 595.950 694.050 596.400 ;
        RECT 721.950 595.950 724.050 596.400 ;
        RECT 769.950 597.600 772.050 598.050 ;
        RECT 817.950 597.600 820.050 598.050 ;
        RECT 769.950 596.400 820.050 597.600 ;
        RECT 769.950 595.950 772.050 596.400 ;
        RECT 817.950 595.950 820.050 596.400 ;
        RECT 832.950 595.950 835.050 598.050 ;
        RECT 319.950 593.400 327.600 594.600 ;
        RECT 319.950 592.950 322.050 593.400 ;
        RECT 133.950 591.600 136.050 592.050 ;
        RECT 113.400 590.400 136.050 591.600 ;
        RECT 133.950 589.950 136.050 590.400 ;
        RECT 139.950 591.600 142.050 592.050 ;
        RECT 148.950 591.600 151.050 592.050 ;
        RECT 139.950 590.400 151.050 591.600 ;
        RECT 139.950 589.950 142.050 590.400 ;
        RECT 148.950 589.950 151.050 590.400 ;
        RECT 244.950 591.600 247.050 592.050 ;
        RECT 259.800 591.600 261.900 592.050 ;
        RECT 244.950 590.400 261.900 591.600 ;
        RECT 244.950 589.950 247.050 590.400 ;
        RECT 259.800 589.950 261.900 590.400 ;
        RECT 262.950 591.600 265.050 592.050 ;
        RECT 268.950 591.600 271.050 592.050 ;
        RECT 262.950 590.400 271.050 591.600 ;
        RECT 262.950 589.950 265.050 590.400 ;
        RECT 268.950 589.950 271.050 590.400 ;
        RECT 277.950 591.600 280.050 592.050 ;
        RECT 295.950 591.600 298.050 592.050 ;
        RECT 277.950 590.400 298.050 591.600 ;
        RECT 326.400 591.600 327.600 593.400 ;
        RECT 397.950 593.400 417.600 594.600 ;
        RECT 469.950 594.600 472.050 595.050 ;
        RECT 490.950 594.600 493.050 595.050 ;
        RECT 469.950 593.400 493.050 594.600 ;
        RECT 397.950 592.950 400.050 593.400 ;
        RECT 469.950 592.950 472.050 593.400 ;
        RECT 490.950 592.950 493.050 593.400 ;
        RECT 496.950 594.600 499.050 595.050 ;
        RECT 544.950 594.600 547.050 595.050 ;
        RECT 496.950 593.400 547.050 594.600 ;
        RECT 496.950 592.950 499.050 593.400 ;
        RECT 544.950 592.950 547.050 593.400 ;
        RECT 601.950 594.600 604.050 595.050 ;
        RECT 628.950 594.600 631.050 595.050 ;
        RECT 601.950 593.400 631.050 594.600 ;
        RECT 601.950 592.950 604.050 593.400 ;
        RECT 628.950 592.950 631.050 593.400 ;
        RECT 667.950 594.600 670.050 595.050 ;
        RECT 676.950 594.600 679.050 595.050 ;
        RECT 667.950 593.400 679.050 594.600 ;
        RECT 667.950 592.950 670.050 593.400 ;
        RECT 676.950 592.950 679.050 593.400 ;
        RECT 772.950 594.600 775.050 595.050 ;
        RECT 811.950 594.600 814.050 595.050 ;
        RECT 772.950 593.400 814.050 594.600 ;
        RECT 772.950 592.950 775.050 593.400 ;
        RECT 811.950 592.950 814.050 593.400 ;
        RECT 835.950 594.600 838.050 595.050 ;
        RECT 853.950 594.600 856.050 595.050 ;
        RECT 862.950 594.600 865.050 595.050 ;
        RECT 835.950 593.400 865.050 594.600 ;
        RECT 835.950 592.950 838.050 593.400 ;
        RECT 853.950 592.950 856.050 593.400 ;
        RECT 862.950 592.950 865.050 593.400 ;
        RECT 355.950 591.600 358.050 592.050 ;
        RECT 326.400 590.400 358.050 591.600 ;
        RECT 277.950 589.950 280.050 590.400 ;
        RECT 295.950 589.950 298.050 590.400 ;
        RECT 355.950 589.950 358.050 590.400 ;
        RECT 379.950 591.600 382.050 592.050 ;
        RECT 394.950 591.600 397.050 592.050 ;
        RECT 379.950 590.400 397.050 591.600 ;
        RECT 379.950 589.950 382.050 590.400 ;
        RECT 394.950 589.950 397.050 590.400 ;
        RECT 430.950 591.600 433.050 592.050 ;
        RECT 472.950 591.600 475.050 592.050 ;
        RECT 511.800 591.600 513.900 592.050 ;
        RECT 430.950 590.400 513.900 591.600 ;
        RECT 430.950 589.950 433.050 590.400 ;
        RECT 472.950 589.950 475.050 590.400 ;
        RECT 511.800 589.950 513.900 590.400 ;
        RECT 514.950 591.600 517.050 592.050 ;
        RECT 520.950 591.600 523.050 592.050 ;
        RECT 514.950 590.400 523.050 591.600 ;
        RECT 514.950 589.950 517.050 590.400 ;
        RECT 520.950 589.950 523.050 590.400 ;
        RECT 526.950 591.600 529.050 592.050 ;
        RECT 586.950 591.600 589.050 592.050 ;
        RECT 526.950 590.400 589.050 591.600 ;
        RECT 526.950 589.950 529.050 590.400 ;
        RECT 586.950 589.950 589.050 590.400 ;
        RECT 592.950 591.600 595.050 592.050 ;
        RECT 688.950 591.600 691.050 592.050 ;
        RECT 592.950 590.400 691.050 591.600 ;
        RECT 592.950 589.950 595.050 590.400 ;
        RECT 688.950 589.950 691.050 590.400 ;
        RECT 694.950 591.600 697.050 592.050 ;
        RECT 847.950 591.600 850.050 592.050 ;
        RECT 694.950 590.400 850.050 591.600 ;
        RECT 694.950 589.950 697.050 590.400 ;
        RECT 847.950 589.950 850.050 590.400 ;
        RECT 31.950 588.600 34.050 589.050 ;
        RECT 82.950 588.600 85.050 589.050 ;
        RECT 109.950 588.600 112.050 589.050 ;
        RECT 31.950 587.400 112.050 588.600 ;
        RECT 31.950 586.950 34.050 587.400 ;
        RECT 82.950 586.950 85.050 587.400 ;
        RECT 109.950 586.950 112.050 587.400 ;
        RECT 157.950 588.600 160.050 589.050 ;
        RECT 166.950 588.600 169.050 589.050 ;
        RECT 157.950 587.400 169.050 588.600 ;
        RECT 157.950 586.950 160.050 587.400 ;
        RECT 166.950 586.950 169.050 587.400 ;
        RECT 178.950 588.600 181.050 589.050 ;
        RECT 220.950 588.600 223.050 589.050 ;
        RECT 229.950 588.600 232.050 589.050 ;
        RECT 178.950 587.400 232.050 588.600 ;
        RECT 178.950 586.950 181.050 587.400 ;
        RECT 220.950 586.950 223.050 587.400 ;
        RECT 229.950 586.950 232.050 587.400 ;
        RECT 241.950 588.600 244.050 589.050 ;
        RECT 262.950 588.600 265.050 588.900 ;
        RECT 241.950 587.400 265.050 588.600 ;
        RECT 241.950 586.950 244.050 587.400 ;
        RECT 262.950 586.800 265.050 587.400 ;
        RECT 307.950 588.600 310.050 589.050 ;
        RECT 355.950 588.600 358.050 588.900 ;
        RECT 307.950 587.400 358.050 588.600 ;
        RECT 307.950 586.950 310.050 587.400 ;
        RECT 355.950 586.800 358.050 587.400 ;
        RECT 364.950 588.600 367.050 589.050 ;
        RECT 409.800 588.600 411.900 589.050 ;
        RECT 364.950 587.400 411.900 588.600 ;
        RECT 364.950 586.950 367.050 587.400 ;
        RECT 409.800 586.950 411.900 587.400 ;
        RECT 412.950 588.600 415.050 589.050 ;
        RECT 418.950 588.600 421.050 589.050 ;
        RECT 412.950 587.400 421.050 588.600 ;
        RECT 412.950 586.950 415.050 587.400 ;
        RECT 418.950 586.950 421.050 587.400 ;
        RECT 463.950 588.600 466.050 589.050 ;
        RECT 472.950 588.600 475.050 588.900 ;
        RECT 463.950 587.400 475.050 588.600 ;
        RECT 463.950 586.950 466.050 587.400 ;
        RECT 472.950 586.800 475.050 587.400 ;
        RECT 508.950 588.600 511.050 589.050 ;
        RECT 521.400 588.600 522.600 589.950 ;
        RECT 529.950 588.600 532.050 589.050 ;
        RECT 508.950 587.400 532.050 588.600 ;
        RECT 508.950 586.950 511.050 587.400 ;
        RECT 529.950 586.950 532.050 587.400 ;
        RECT 538.950 588.600 541.050 589.050 ;
        RECT 577.950 588.600 580.050 589.050 ;
        RECT 538.950 587.400 580.050 588.600 ;
        RECT 538.950 586.950 541.050 587.400 ;
        RECT 577.950 586.950 580.050 587.400 ;
        RECT 613.950 588.600 616.050 589.050 ;
        RECT 658.950 588.600 661.050 589.050 ;
        RECT 757.950 588.600 760.050 589.050 ;
        RECT 613.950 587.400 661.050 588.600 ;
        RECT 613.950 586.950 616.050 587.400 ;
        RECT 658.950 586.950 661.050 587.400 ;
        RECT 746.400 587.400 760.050 588.600 ;
        RECT 746.400 586.050 747.600 587.400 ;
        RECT 757.950 586.950 760.050 587.400 ;
        RECT 10.950 585.600 13.050 586.050 ;
        RECT 19.950 585.600 22.050 586.050 ;
        RECT 10.950 584.400 22.050 585.600 ;
        RECT 10.950 583.950 13.050 584.400 ;
        RECT 19.950 583.950 22.050 584.400 ;
        RECT 55.950 585.600 58.050 586.050 ;
        RECT 67.950 585.600 70.050 586.050 ;
        RECT 121.950 585.600 124.050 586.050 ;
        RECT 55.950 584.400 124.050 585.600 ;
        RECT 55.950 583.950 58.050 584.400 ;
        RECT 67.950 583.950 70.050 584.400 ;
        RECT 121.950 583.950 124.050 584.400 ;
        RECT 139.950 585.600 142.050 586.050 ;
        RECT 163.950 585.600 166.050 586.050 ;
        RECT 139.950 584.400 166.050 585.600 ;
        RECT 139.950 583.950 142.050 584.400 ;
        RECT 163.950 583.950 166.050 584.400 ;
        RECT 265.950 585.600 268.050 586.050 ;
        RECT 274.950 585.600 277.050 586.050 ;
        RECT 319.950 585.600 322.050 586.050 ;
        RECT 265.950 584.400 322.050 585.600 ;
        RECT 265.950 583.950 268.050 584.400 ;
        RECT 274.950 583.950 277.050 584.400 ;
        RECT 319.950 583.950 322.050 584.400 ;
        RECT 445.950 585.600 448.050 586.050 ;
        RECT 466.950 585.600 469.050 586.050 ;
        RECT 445.950 584.400 469.050 585.600 ;
        RECT 445.950 583.950 448.050 584.400 ;
        RECT 466.950 583.950 469.050 584.400 ;
        RECT 532.950 585.600 535.050 586.050 ;
        RECT 547.950 585.600 550.050 586.050 ;
        RECT 532.950 584.400 550.050 585.600 ;
        RECT 532.950 583.950 535.050 584.400 ;
        RECT 547.950 583.950 550.050 584.400 ;
        RECT 595.950 585.600 598.050 586.050 ;
        RECT 604.950 585.600 607.050 586.050 ;
        RECT 595.950 584.400 607.050 585.600 ;
        RECT 595.950 583.950 598.050 584.400 ;
        RECT 604.950 583.950 607.050 584.400 ;
        RECT 619.950 585.600 622.050 586.050 ;
        RECT 634.950 585.600 637.050 586.050 ;
        RECT 619.950 584.400 637.050 585.600 ;
        RECT 619.950 583.950 622.050 584.400 ;
        RECT 634.950 583.950 637.050 584.400 ;
        RECT 706.950 585.600 709.050 586.050 ;
        RECT 712.950 585.600 715.050 586.050 ;
        RECT 706.950 584.400 715.050 585.600 ;
        RECT 706.950 583.950 709.050 584.400 ;
        RECT 712.950 583.950 715.050 584.400 ;
        RECT 727.950 585.600 730.050 586.050 ;
        RECT 745.950 585.600 748.050 586.050 ;
        RECT 727.950 584.400 748.050 585.600 ;
        RECT 727.950 583.950 730.050 584.400 ;
        RECT 745.950 583.950 748.050 584.400 ;
        RECT 829.950 585.600 832.050 586.050 ;
        RECT 862.950 585.600 865.050 586.050 ;
        RECT 829.950 584.400 865.050 585.600 ;
        RECT 829.950 583.950 832.050 584.400 ;
        RECT 862.950 583.950 865.050 584.400 ;
        RECT 136.950 582.600 139.050 583.050 ;
        RECT 145.950 582.600 148.050 583.050 ;
        RECT 136.950 581.400 148.050 582.600 ;
        RECT 136.950 580.950 139.050 581.400 ;
        RECT 145.950 580.950 148.050 581.400 ;
        RECT 154.950 582.600 157.050 583.050 ;
        RECT 163.950 582.600 166.050 582.900 ;
        RECT 154.950 581.400 166.050 582.600 ;
        RECT 154.950 580.950 157.050 581.400 ;
        RECT 163.950 580.800 166.050 581.400 ;
        RECT 190.950 582.600 193.050 583.050 ;
        RECT 211.950 582.600 214.050 583.050 ;
        RECT 190.950 581.400 214.050 582.600 ;
        RECT 190.950 580.950 193.050 581.400 ;
        RECT 211.950 580.950 214.050 581.400 ;
        RECT 346.950 582.600 349.050 583.050 ;
        RECT 373.950 582.600 376.050 583.050 ;
        RECT 346.950 581.400 376.050 582.600 ;
        RECT 346.950 580.950 349.050 581.400 ;
        RECT 373.950 580.950 376.050 581.400 ;
        RECT 391.950 582.600 394.050 583.050 ;
        RECT 415.950 582.600 418.050 583.050 ;
        RECT 391.950 581.400 418.050 582.600 ;
        RECT 391.950 580.950 394.050 581.400 ;
        RECT 415.950 580.950 418.050 581.400 ;
        RECT 451.950 582.600 454.050 583.050 ;
        RECT 526.950 582.600 529.050 583.050 ;
        RECT 451.950 581.400 529.050 582.600 ;
        RECT 451.950 580.950 454.050 581.400 ;
        RECT 526.950 580.950 529.050 581.400 ;
        RECT 535.950 582.600 538.050 583.050 ;
        RECT 574.950 582.600 577.050 583.050 ;
        RECT 535.950 581.400 577.050 582.600 ;
        RECT 535.950 580.950 538.050 581.400 ;
        RECT 574.950 580.950 577.050 581.400 ;
        RECT 592.950 582.600 595.050 583.050 ;
        RECT 610.950 582.600 613.050 583.050 ;
        RECT 652.950 582.600 655.050 583.050 ;
        RECT 664.950 582.600 667.050 583.050 ;
        RECT 592.950 581.400 606.600 582.600 ;
        RECT 592.950 580.950 595.050 581.400 ;
        RECT 1.950 579.600 4.050 580.050 ;
        RECT 13.950 579.600 16.050 580.050 ;
        RECT 1.950 578.400 16.050 579.600 ;
        RECT 1.950 577.950 4.050 578.400 ;
        RECT 13.950 577.950 16.050 578.400 ;
        RECT 49.950 579.600 52.050 580.050 ;
        RECT 61.950 579.600 64.050 580.050 ;
        RECT 49.950 578.400 64.050 579.600 ;
        RECT 49.950 577.950 52.050 578.400 ;
        RECT 61.950 577.950 64.050 578.400 ;
        RECT 85.950 579.600 88.050 580.050 ;
        RECT 97.950 579.600 100.050 580.050 ;
        RECT 85.950 578.400 100.050 579.600 ;
        RECT 85.950 577.950 88.050 578.400 ;
        RECT 97.950 577.950 100.050 578.400 ;
        RECT 184.950 579.600 187.050 580.050 ;
        RECT 238.950 579.600 241.050 580.050 ;
        RECT 244.950 579.600 247.050 580.050 ;
        RECT 184.950 578.400 198.600 579.600 ;
        RECT 184.950 577.950 187.050 578.400 ;
        RECT 197.400 577.050 198.600 578.400 ;
        RECT 238.950 578.400 247.050 579.600 ;
        RECT 238.950 577.950 241.050 578.400 ;
        RECT 244.950 577.950 247.050 578.400 ;
        RECT 271.950 579.600 274.050 580.050 ;
        RECT 280.950 579.600 283.050 580.050 ;
        RECT 271.950 578.400 283.050 579.600 ;
        RECT 271.950 577.950 274.050 578.400 ;
        RECT 280.950 577.950 283.050 578.400 ;
        RECT 319.950 579.600 322.050 580.050 ;
        RECT 325.950 579.600 328.050 580.050 ;
        RECT 366.000 579.600 370.050 580.050 ;
        RECT 319.950 578.400 328.050 579.600 ;
        RECT 319.950 577.950 322.050 578.400 ;
        RECT 325.950 577.950 328.050 578.400 ;
        RECT 365.400 577.950 370.050 579.600 ;
        RECT 385.950 579.600 388.050 580.050 ;
        RECT 505.950 579.600 508.050 580.050 ;
        RECT 517.950 579.600 520.050 580.050 ;
        RECT 385.950 578.400 399.600 579.600 ;
        RECT 385.950 577.950 388.050 578.400 ;
        RECT 4.950 576.600 7.050 577.050 ;
        RECT 25.950 576.600 28.050 577.050 ;
        RECT 4.950 575.400 28.050 576.600 ;
        RECT 4.950 574.950 7.050 575.400 ;
        RECT 25.950 574.950 28.050 575.400 ;
        RECT 115.950 576.600 118.050 577.050 ;
        RECT 130.950 576.600 133.050 577.050 ;
        RECT 151.800 576.600 153.900 576.900 ;
        RECT 156.000 576.600 160.050 577.050 ;
        RECT 115.950 575.400 153.900 576.600 ;
        RECT 115.950 574.950 118.050 575.400 ;
        RECT 130.950 574.950 133.050 575.400 ;
        RECT 151.800 574.800 153.900 575.400 ;
        RECT 155.400 574.950 160.050 576.600 ;
        RECT 172.950 574.950 175.050 577.050 ;
        RECT 193.800 576.000 195.900 577.050 ;
        RECT 196.950 576.600 199.050 577.050 ;
        RECT 208.950 576.600 211.050 577.050 ;
        RECT 193.800 574.950 196.050 576.000 ;
        RECT 196.950 575.400 211.050 576.600 ;
        RECT 196.950 574.950 199.050 575.400 ;
        RECT 208.950 574.950 211.050 575.400 ;
        RECT 214.950 576.600 217.050 577.050 ;
        RECT 223.950 576.600 226.050 577.050 ;
        RECT 214.950 575.400 226.050 576.600 ;
        RECT 214.950 574.950 217.050 575.400 ;
        RECT 223.950 574.950 226.050 575.400 ;
        RECT 325.950 576.600 328.050 576.900 ;
        RECT 325.950 575.400 357.600 576.600 ;
        RECT 19.950 573.600 24.000 574.050 ;
        RECT 49.950 573.600 52.050 574.200 ;
        RECT 64.950 573.600 69.000 574.050 ;
        RECT 73.950 573.900 76.050 574.350 ;
        RECT 79.950 573.900 82.050 574.350 ;
        RECT 73.950 573.600 82.050 573.900 ;
        RECT 88.950 573.600 91.050 574.350 ;
        RECT 19.950 571.950 24.600 573.600 ;
        RECT 49.950 572.400 57.600 573.600 ;
        RECT 49.950 572.100 52.050 572.400 ;
        RECT 23.400 568.050 24.600 571.950 ;
        RECT 4.950 567.600 7.050 568.050 ;
        RECT 10.950 567.600 13.050 567.900 ;
        RECT 4.950 566.400 13.050 567.600 ;
        RECT 4.950 565.950 7.050 566.400 ;
        RECT 10.950 565.800 13.050 566.400 ;
        RECT 22.950 565.950 25.050 568.050 ;
        RECT 28.950 567.600 31.050 568.050 ;
        RECT 37.950 567.600 40.050 568.050 ;
        RECT 52.950 567.600 55.050 567.900 ;
        RECT 28.950 566.400 55.050 567.600 ;
        RECT 28.950 565.950 31.050 566.400 ;
        RECT 37.950 565.950 40.050 566.400 ;
        RECT 52.950 565.800 55.050 566.400 ;
        RECT 56.400 565.050 57.600 572.400 ;
        RECT 64.950 571.950 69.600 573.600 ;
        RECT 73.950 572.700 91.050 573.600 ;
        RECT 73.950 572.250 76.050 572.700 ;
        RECT 79.950 572.400 91.050 572.700 ;
        RECT 79.950 572.250 82.050 572.400 ;
        RECT 88.950 572.250 91.050 572.400 ;
        RECT 94.950 572.250 97.050 574.350 ;
        RECT 100.950 573.750 103.050 574.200 ;
        RECT 106.950 573.750 109.050 574.200 ;
        RECT 100.950 572.550 109.050 573.750 ;
        RECT 68.400 568.050 69.600 571.950 ;
        RECT 95.400 570.600 96.600 572.250 ;
        RECT 100.950 572.100 103.050 572.550 ;
        RECT 106.950 572.100 109.050 572.550 ;
        RECT 112.950 572.100 115.050 574.200 ;
        RECT 113.400 570.600 114.600 572.100 ;
        RECT 142.950 570.600 145.050 571.050 ;
        RECT 95.400 570.000 99.600 570.600 ;
        RECT 95.400 569.400 100.050 570.000 ;
        RECT 113.400 569.400 145.050 570.600 ;
        RECT 67.950 565.950 70.050 568.050 ;
        RECT 97.950 565.950 100.050 569.400 ;
        RECT 109.950 567.450 112.050 567.900 ;
        RECT 121.950 567.450 124.050 567.900 ;
        RECT 109.950 566.250 124.050 567.450 ;
        RECT 109.950 565.800 112.050 566.250 ;
        RECT 121.950 565.800 124.050 566.250 ;
        RECT 133.950 565.950 136.050 569.400 ;
        RECT 142.950 568.950 145.050 569.400 ;
        RECT 155.400 568.050 156.600 574.950 ;
        RECT 169.950 573.600 172.050 574.050 ;
        RECT 161.400 572.400 172.050 573.600 ;
        RECT 161.400 568.050 162.600 572.400 ;
        RECT 169.950 571.950 172.050 572.400 ;
        RECT 173.400 568.050 174.600 574.950 ;
        RECT 183.000 573.600 187.050 574.050 ;
        RECT 182.400 571.950 187.050 573.600 ;
        RECT 193.950 573.600 196.050 574.950 ;
        RECT 325.950 574.800 328.050 575.400 ;
        RECT 193.950 573.000 201.450 573.600 ;
        RECT 194.400 572.400 201.450 573.000 ;
        RECT 182.400 568.050 183.600 571.950 ;
        RECT 200.250 568.050 201.450 572.400 ;
        RECT 202.950 571.950 205.050 574.050 ;
        RECT 219.000 573.600 223.050 574.050 ;
        RECT 232.950 573.600 235.050 574.350 ;
        RECT 244.800 573.600 246.900 574.050 ;
        RECT 218.400 571.950 223.050 573.600 ;
        RECT 227.400 572.400 235.050 573.600 ;
        RECT 203.400 568.050 204.600 571.950 ;
        RECT 154.950 565.950 157.050 568.050 ;
        RECT 160.950 565.950 163.050 568.050 ;
        RECT 172.950 565.950 175.050 568.050 ;
        RECT 181.950 565.950 184.050 568.050 ;
        RECT 199.800 565.950 201.900 568.050 ;
        RECT 202.950 565.950 205.050 568.050 ;
        RECT 218.400 567.900 219.600 571.950 ;
        RECT 227.400 567.900 228.600 572.400 ;
        RECT 232.950 572.250 235.050 572.400 ;
        RECT 236.400 572.400 246.900 573.600 ;
        RECT 236.400 570.600 237.600 572.400 ;
        RECT 244.800 571.950 246.900 572.400 ;
        RECT 247.950 573.600 252.000 574.050 ;
        RECT 247.950 571.950 252.600 573.600 ;
        RECT 253.950 572.250 256.050 574.350 ;
        RECT 258.000 573.600 262.050 574.050 ;
        RECT 233.400 570.000 237.600 570.600 ;
        RECT 232.950 569.400 237.600 570.000 ;
        RECT 217.950 565.800 220.050 567.900 ;
        RECT 226.950 565.800 229.050 567.900 ;
        RECT 232.950 565.950 235.050 569.400 ;
        RECT 251.400 568.050 252.600 571.950 ;
        RECT 250.950 565.950 253.050 568.050 ;
        RECT 55.950 562.950 58.050 565.050 ;
        RECT 70.950 564.600 73.050 565.050 ;
        RECT 85.950 564.600 88.050 565.050 ;
        RECT 70.950 563.400 88.050 564.600 ;
        RECT 70.950 562.950 73.050 563.400 ;
        RECT 85.950 562.950 88.050 563.400 ;
        RECT 103.950 564.600 106.050 565.050 ;
        RECT 127.950 564.600 130.050 565.050 ;
        RECT 142.950 564.600 145.050 565.050 ;
        RECT 103.950 563.400 145.050 564.600 ;
        RECT 103.950 562.950 106.050 563.400 ;
        RECT 127.950 562.950 130.050 563.400 ;
        RECT 142.950 562.950 145.050 563.400 ;
        RECT 238.950 564.600 241.050 565.050 ;
        RECT 254.400 564.600 255.600 572.250 ;
        RECT 238.950 563.400 255.600 564.600 ;
        RECT 257.400 571.950 262.050 573.600 ;
        RECT 301.950 573.600 306.000 574.050 ;
        RECT 301.950 571.950 306.600 573.600 ;
        RECT 322.800 573.000 324.900 574.050 ;
        RECT 322.800 571.950 325.050 573.000 ;
        RECT 325.950 571.950 328.050 574.050 ;
        RECT 343.950 573.600 346.050 574.050 ;
        RECT 352.950 573.600 355.050 574.350 ;
        RECT 343.950 572.400 355.050 573.600 ;
        RECT 343.950 571.950 346.050 572.400 ;
        RECT 352.950 572.250 355.050 572.400 ;
        RECT 238.950 562.950 241.050 563.400 ;
        RECT 1.950 561.600 4.050 562.050 ;
        RECT 46.950 561.600 49.050 562.050 ;
        RECT 100.950 561.600 103.050 562.050 ;
        RECT 1.950 560.400 103.050 561.600 ;
        RECT 1.950 559.950 4.050 560.400 ;
        RECT 46.950 559.950 49.050 560.400 ;
        RECT 100.950 559.950 103.050 560.400 ;
        RECT 163.950 561.600 166.050 562.050 ;
        RECT 187.950 561.600 190.050 561.900 ;
        RECT 163.950 560.400 190.050 561.600 ;
        RECT 163.950 559.950 166.050 560.400 ;
        RECT 187.950 559.800 190.050 560.400 ;
        RECT 208.950 561.600 211.050 562.050 ;
        RECT 223.950 561.600 226.050 562.050 ;
        RECT 235.950 561.600 238.050 562.050 ;
        RECT 208.950 560.400 238.050 561.600 ;
        RECT 208.950 559.950 211.050 560.400 ;
        RECT 223.950 559.950 226.050 560.400 ;
        RECT 235.950 559.950 238.050 560.400 ;
        RECT 241.950 561.600 244.050 562.050 ;
        RECT 257.400 561.600 258.600 571.950 ;
        RECT 305.400 570.600 306.600 571.950 ;
        RECT 322.950 570.600 325.050 571.950 ;
        RECT 275.400 570.000 306.600 570.600 ;
        RECT 274.950 569.400 306.600 570.000 ;
        RECT 259.950 567.600 262.050 568.050 ;
        RECT 274.950 567.600 277.050 569.400 ;
        RECT 305.400 568.050 306.600 569.400 ;
        RECT 320.400 570.000 325.050 570.600 ;
        RECT 320.400 569.400 324.450 570.000 ;
        RECT 259.950 566.400 277.050 567.600 ;
        RECT 259.950 565.950 262.050 566.400 ;
        RECT 274.950 565.950 277.050 566.400 ;
        RECT 304.950 565.950 307.050 568.050 ;
        RECT 286.950 564.600 289.050 565.050 ;
        RECT 320.400 564.600 321.600 569.400 ;
        RECT 326.400 568.050 327.600 571.950 ;
        RECT 356.400 568.050 357.600 575.400 ;
        RECT 365.400 568.050 366.600 577.950 ;
        RECT 370.950 574.950 373.050 577.050 ;
        RECT 398.400 576.600 399.600 578.400 ;
        RECT 505.950 578.400 520.050 579.600 ;
        RECT 505.950 577.950 508.050 578.400 ;
        RECT 517.950 577.950 520.050 578.400 ;
        RECT 529.950 579.600 532.050 580.050 ;
        RECT 550.950 579.600 553.050 580.050 ;
        RECT 529.950 578.400 553.050 579.600 ;
        RECT 529.950 577.950 532.050 578.400 ;
        RECT 550.950 577.950 553.050 578.400 ;
        RECT 586.950 579.600 589.050 580.050 ;
        RECT 595.950 579.600 598.050 580.050 ;
        RECT 586.950 578.400 598.050 579.600 ;
        RECT 605.400 579.600 606.600 581.400 ;
        RECT 610.950 581.400 667.050 582.600 ;
        RECT 610.950 580.950 613.050 581.400 ;
        RECT 652.950 580.950 655.050 581.400 ;
        RECT 664.950 580.950 667.050 581.400 ;
        RECT 691.950 582.600 694.050 583.050 ;
        RECT 748.950 582.600 751.050 583.050 ;
        RECT 691.950 581.400 751.050 582.600 ;
        RECT 691.950 580.950 694.050 581.400 ;
        RECT 748.950 580.950 751.050 581.400 ;
        RECT 718.950 579.600 721.050 580.050 ;
        RECT 733.950 579.600 736.050 580.050 ;
        RECT 605.400 578.400 615.600 579.600 ;
        RECT 586.950 577.950 589.050 578.400 ;
        RECT 595.950 577.950 598.050 578.400 ;
        RECT 403.950 576.600 406.050 577.050 ;
        RECT 398.400 575.400 406.050 576.600 ;
        RECT 403.950 574.950 406.050 575.400 ;
        RECT 538.950 576.600 543.000 577.050 ;
        RECT 601.950 576.600 604.050 577.050 ;
        RECT 538.950 574.950 543.600 576.600 ;
        RECT 322.950 566.400 327.600 568.050 ;
        RECT 334.950 567.600 337.050 567.900 ;
        RECT 349.950 567.600 352.050 568.050 ;
        RECT 334.950 566.400 352.050 567.600 ;
        RECT 322.950 565.950 327.000 566.400 ;
        RECT 334.950 565.800 337.050 566.400 ;
        RECT 349.950 565.950 352.050 566.400 ;
        RECT 355.950 565.950 358.050 568.050 ;
        RECT 364.950 565.950 367.050 568.050 ;
        RECT 371.400 567.600 372.600 574.950 ;
        RECT 373.950 573.900 376.050 574.350 ;
        RECT 394.950 573.900 397.050 574.350 ;
        RECT 373.950 572.700 397.050 573.900 ;
        RECT 373.950 572.250 376.050 572.700 ;
        RECT 394.950 572.250 397.050 572.700 ;
        RECT 409.950 571.950 412.050 574.050 ;
        RECT 424.950 572.100 427.050 574.200 ;
        RECT 481.950 573.600 484.050 574.350 ;
        RECT 505.950 573.600 508.050 574.200 ;
        RECT 514.800 573.600 516.900 574.050 ;
        RECT 481.950 572.400 498.600 573.600 ;
        RECT 481.950 572.250 484.050 572.400 ;
        RECT 410.400 568.050 411.600 571.950 ;
        RECT 425.400 570.600 426.600 572.100 ;
        RECT 425.400 569.400 429.600 570.600 ;
        RECT 379.950 567.600 382.050 568.050 ;
        RECT 371.400 566.400 382.050 567.600 ;
        RECT 379.950 565.950 382.050 566.400 ;
        RECT 388.950 567.600 391.050 567.900 ;
        RECT 394.950 567.600 397.050 568.050 ;
        RECT 388.950 566.400 397.050 567.600 ;
        RECT 388.950 565.800 391.050 566.400 ;
        RECT 394.950 565.950 397.050 566.400 ;
        RECT 409.950 565.950 412.050 568.050 ;
        RECT 428.400 567.600 429.600 569.400 ;
        RECT 497.400 567.900 498.600 572.400 ;
        RECT 505.950 572.400 516.900 573.600 ;
        RECT 505.950 572.100 508.050 572.400 ;
        RECT 445.950 567.600 448.050 567.900 ;
        RECT 428.400 566.400 448.050 567.600 ;
        RECT 445.950 565.800 448.050 566.400 ;
        RECT 496.950 565.800 499.050 567.900 ;
        RECT 506.400 567.600 507.600 572.100 ;
        RECT 514.800 571.950 516.900 572.400 ;
        RECT 517.950 573.600 520.050 574.350 ;
        RECT 517.950 572.400 528.600 573.600 ;
        RECT 517.950 572.250 520.050 572.400 ;
        RECT 527.400 568.050 528.600 572.400 ;
        RECT 529.950 572.100 532.050 574.200 ;
        RECT 535.950 572.100 538.050 574.200 ;
        RECT 500.400 566.400 507.600 567.600 ;
        RECT 286.950 563.400 321.600 564.600 ;
        RECT 343.950 564.600 346.050 565.050 ;
        RECT 370.950 564.600 373.050 565.050 ;
        RECT 343.950 563.400 373.050 564.600 ;
        RECT 286.950 562.950 289.050 563.400 ;
        RECT 343.950 562.950 346.050 563.400 ;
        RECT 370.950 562.950 373.050 563.400 ;
        RECT 241.950 560.400 258.600 561.600 ;
        RECT 307.950 561.600 310.050 562.050 ;
        RECT 322.950 561.600 325.050 562.050 ;
        RECT 307.950 560.400 325.050 561.600 ;
        RECT 241.950 559.950 244.050 560.400 ;
        RECT 307.950 559.950 310.050 560.400 ;
        RECT 322.950 559.950 325.050 560.400 ;
        RECT 382.950 561.600 385.050 562.050 ;
        RECT 415.950 561.600 418.050 562.050 ;
        RECT 382.950 560.400 418.050 561.600 ;
        RECT 382.950 559.950 385.050 560.400 ;
        RECT 415.950 559.950 418.050 560.400 ;
        RECT 445.950 561.600 448.050 562.050 ;
        RECT 454.950 561.600 457.050 562.050 ;
        RECT 445.950 560.400 457.050 561.600 ;
        RECT 445.950 559.950 448.050 560.400 ;
        RECT 454.950 559.950 457.050 560.400 ;
        RECT 484.950 561.600 487.050 562.050 ;
        RECT 500.400 561.600 501.600 566.400 ;
        RECT 526.950 565.950 529.050 568.050 ;
        RECT 523.950 564.600 526.050 565.050 ;
        RECT 530.400 564.600 531.600 572.100 ;
        RECT 536.400 570.600 537.600 572.100 ;
        RECT 542.400 570.600 543.600 574.950 ;
        RECT 593.400 575.400 604.050 576.600 ;
        RECT 547.950 573.600 552.000 574.050 ;
        RECT 568.950 573.600 571.050 574.200 ;
        RECT 547.950 571.950 552.600 573.600 ;
        RECT 536.400 569.400 543.600 570.600 ;
        RECT 551.400 568.050 552.600 571.950 ;
        RECT 563.400 572.400 571.050 573.600 ;
        RECT 563.400 568.050 564.600 572.400 ;
        RECT 568.950 572.100 571.050 572.400 ;
        RECT 574.950 573.600 577.050 574.200 ;
        RECT 593.400 573.600 594.600 575.400 ;
        RECT 601.950 574.950 604.050 575.400 ;
        RECT 604.950 573.600 607.050 574.200 ;
        RECT 574.950 572.400 594.600 573.600 ;
        RECT 596.250 572.400 607.050 573.600 ;
        RECT 574.950 572.100 577.050 572.400 ;
        RECT 590.400 568.050 591.600 572.400 ;
        RECT 596.250 568.050 597.450 572.400 ;
        RECT 604.950 572.100 607.050 572.400 ;
        RECT 538.950 567.450 541.050 567.900 ;
        RECT 544.950 567.450 547.050 567.900 ;
        RECT 538.950 566.250 547.050 567.450 ;
        RECT 538.950 565.800 541.050 566.250 ;
        RECT 544.950 565.800 547.050 566.250 ;
        RECT 550.950 565.950 553.050 568.050 ;
        RECT 559.950 566.400 564.600 568.050 ;
        RECT 571.950 567.600 574.050 567.900 ;
        RECT 580.950 567.600 583.050 567.900 ;
        RECT 571.950 566.400 583.050 567.600 ;
        RECT 559.950 565.950 564.000 566.400 ;
        RECT 571.950 565.800 574.050 566.400 ;
        RECT 580.950 565.800 583.050 566.400 ;
        RECT 589.950 565.950 592.050 568.050 ;
        RECT 595.800 565.950 597.900 568.050 ;
        RECT 614.400 567.900 615.600 578.400 ;
        RECT 718.950 578.400 736.050 579.600 ;
        RECT 718.950 577.950 721.050 578.400 ;
        RECT 733.950 577.950 736.050 578.400 ;
        RECT 775.950 579.600 778.050 580.050 ;
        RECT 802.950 579.600 805.050 580.050 ;
        RECT 775.950 578.400 805.050 579.600 ;
        RECT 775.950 577.950 778.050 578.400 ;
        RECT 802.950 577.950 805.050 578.400 ;
        RECT 829.950 579.600 832.050 580.050 ;
        RECT 841.950 579.600 844.050 580.050 ;
        RECT 829.950 578.400 844.050 579.600 ;
        RECT 829.950 577.950 832.050 578.400 ;
        RECT 841.950 577.950 844.050 578.400 ;
        RECT 646.950 576.600 649.050 577.200 ;
        RECT 635.400 575.400 649.050 576.600 ;
        RECT 622.950 570.600 625.050 570.900 ;
        RECT 635.400 570.600 636.600 575.400 ;
        RECT 646.950 575.100 649.050 575.400 ;
        RECT 682.950 576.600 685.050 577.050 ;
        RECT 691.950 576.600 694.050 577.050 ;
        RECT 682.950 575.400 694.050 576.600 ;
        RECT 682.950 574.950 685.050 575.400 ;
        RECT 691.950 574.950 694.050 575.400 ;
        RECT 712.950 576.600 715.050 577.050 ;
        RECT 739.950 576.600 742.050 577.050 ;
        RECT 772.950 576.600 775.050 577.050 ;
        RECT 781.950 576.600 784.050 577.050 ;
        RECT 712.950 575.400 744.600 576.600 ;
        RECT 712.950 574.950 715.050 575.400 ;
        RECT 739.950 574.950 742.050 575.400 ;
        RECT 646.800 571.950 648.900 574.050 ;
        RECT 649.950 573.600 652.050 574.050 ;
        RECT 658.950 573.600 661.050 573.900 ;
        RECT 649.950 572.400 661.050 573.600 ;
        RECT 649.950 571.950 652.050 572.400 ;
        RECT 622.950 569.400 636.600 570.600 ;
        RECT 647.400 570.600 648.600 571.950 ;
        RECT 658.950 571.800 661.050 572.400 ;
        RECT 676.950 571.950 679.050 574.050 ;
        RECT 697.950 573.600 700.050 574.050 ;
        RECT 706.950 573.600 709.050 574.200 ;
        RECT 697.950 572.400 709.050 573.600 ;
        RECT 697.950 571.950 700.050 572.400 ;
        RECT 706.950 572.100 709.050 572.400 ;
        RECT 647.400 570.000 651.600 570.600 ;
        RECT 647.400 569.400 652.050 570.000 ;
        RECT 622.950 568.800 625.050 569.400 ;
        RECT 598.950 567.450 601.050 567.900 ;
        RECT 607.950 567.450 610.050 567.900 ;
        RECT 598.950 566.250 610.050 567.450 ;
        RECT 598.950 565.800 601.050 566.250 ;
        RECT 607.950 565.800 610.050 566.250 ;
        RECT 613.950 567.600 616.050 567.900 ;
        RECT 637.950 567.600 640.050 568.050 ;
        RECT 613.950 566.400 640.050 567.600 ;
        RECT 613.950 565.800 616.050 566.400 ;
        RECT 637.950 565.950 640.050 566.400 ;
        RECT 649.950 565.950 652.050 569.400 ;
        RECT 677.400 568.050 678.600 571.950 ;
        RECT 743.400 568.050 744.600 575.400 ;
        RECT 772.950 575.400 784.050 576.600 ;
        RECT 772.950 574.950 775.050 575.400 ;
        RECT 781.950 574.950 784.050 575.400 ;
        RECT 811.950 576.600 814.050 577.050 ;
        RECT 823.950 576.600 826.050 577.050 ;
        RECT 811.950 575.400 826.050 576.600 ;
        RECT 811.950 574.950 814.050 575.400 ;
        RECT 823.950 574.950 826.050 575.400 ;
        RECT 751.950 571.950 754.050 574.050 ;
        RECT 787.950 573.600 790.050 574.200 ;
        RECT 785.400 572.400 790.050 573.600 ;
        RECT 752.400 568.050 753.600 571.950 ;
        RECT 785.400 568.050 786.600 572.400 ;
        RECT 787.950 572.100 790.050 572.400 ;
        RECT 793.950 573.600 796.050 574.050 ;
        RECT 793.950 572.400 807.600 573.600 ;
        RECT 793.950 571.950 796.050 572.400 ;
        RECT 806.400 568.050 807.600 572.400 ;
        RECT 820.950 571.950 823.050 574.050 ;
        RECT 841.950 573.600 844.050 574.350 ;
        RECT 850.950 573.600 853.050 574.050 ;
        RECT 841.950 572.400 853.050 573.600 ;
        RECT 841.950 572.250 844.050 572.400 ;
        RECT 850.950 571.950 853.050 572.400 ;
        RECT 821.400 568.050 822.600 571.950 ;
        RECT 676.950 565.950 679.050 568.050 ;
        RECT 688.950 567.600 691.050 567.900 ;
        RECT 703.950 567.600 706.050 567.900 ;
        RECT 688.950 566.400 706.050 567.600 ;
        RECT 688.950 565.800 691.050 566.400 ;
        RECT 703.950 565.800 706.050 566.400 ;
        RECT 709.950 567.600 712.050 567.900 ;
        RECT 724.950 567.600 727.050 567.900 ;
        RECT 709.950 566.400 727.050 567.600 ;
        RECT 709.950 565.800 712.050 566.400 ;
        RECT 724.950 565.800 727.050 566.400 ;
        RECT 742.950 565.950 745.050 568.050 ;
        RECT 751.950 565.950 754.050 568.050 ;
        RECT 784.950 565.950 787.050 568.050 ;
        RECT 805.950 565.950 808.050 568.050 ;
        RECT 820.950 565.950 823.050 568.050 ;
        RECT 523.950 563.400 531.600 564.600 ;
        RECT 652.950 564.600 655.050 565.050 ;
        RECT 670.950 564.600 673.050 565.050 ;
        RECT 652.950 563.400 673.050 564.600 ;
        RECT 523.950 562.950 526.050 563.400 ;
        RECT 652.950 562.950 655.050 563.400 ;
        RECT 670.950 562.950 673.050 563.400 ;
        RECT 484.950 560.400 501.600 561.600 ;
        RECT 520.950 561.600 523.050 562.050 ;
        RECT 526.950 561.600 529.050 562.050 ;
        RECT 532.950 561.600 535.050 562.050 ;
        RECT 520.950 560.400 535.050 561.600 ;
        RECT 484.950 559.950 487.050 560.400 ;
        RECT 520.950 559.950 523.050 560.400 ;
        RECT 526.950 559.950 529.050 560.400 ;
        RECT 532.950 559.950 535.050 560.400 ;
        RECT 598.950 561.600 601.050 562.050 ;
        RECT 619.950 561.600 622.050 562.050 ;
        RECT 598.950 560.400 622.050 561.600 ;
        RECT 598.950 559.950 601.050 560.400 ;
        RECT 619.950 559.950 622.050 560.400 ;
        RECT 637.950 561.600 640.050 562.050 ;
        RECT 643.950 561.600 646.050 562.050 ;
        RECT 637.950 560.400 646.050 561.600 ;
        RECT 637.950 559.950 640.050 560.400 ;
        RECT 643.950 559.950 646.050 560.400 ;
        RECT 697.950 561.600 700.050 562.050 ;
        RECT 757.950 561.600 760.050 562.050 ;
        RECT 697.950 560.400 760.050 561.600 ;
        RECT 697.950 559.950 700.050 560.400 ;
        RECT 757.950 559.950 760.050 560.400 ;
        RECT 766.950 561.600 769.050 562.050 ;
        RECT 787.950 561.600 790.050 562.050 ;
        RECT 790.950 561.600 793.050 562.050 ;
        RECT 766.950 560.400 793.050 561.600 ;
        RECT 766.950 559.950 769.050 560.400 ;
        RECT 787.950 559.950 790.050 560.400 ;
        RECT 790.950 559.950 793.050 560.400 ;
        RECT 805.950 561.600 808.050 562.050 ;
        RECT 835.950 561.600 838.050 562.050 ;
        RECT 805.950 560.400 838.050 561.600 ;
        RECT 805.950 559.950 808.050 560.400 ;
        RECT 835.950 559.950 838.050 560.400 ;
        RECT 61.950 558.600 64.050 559.050 ;
        RECT 76.950 558.600 79.050 559.050 ;
        RECT 91.950 558.600 94.050 559.050 ;
        RECT 61.950 557.400 94.050 558.600 ;
        RECT 61.950 556.950 64.050 557.400 ;
        RECT 76.950 556.950 79.050 557.400 ;
        RECT 91.950 556.950 94.050 557.400 ;
        RECT 103.950 558.600 106.050 559.050 ;
        RECT 121.950 558.600 124.050 559.050 ;
        RECT 103.950 557.400 124.050 558.600 ;
        RECT 103.950 556.950 106.050 557.400 ;
        RECT 121.950 556.950 124.050 557.400 ;
        RECT 184.950 558.600 187.050 559.050 ;
        RECT 199.950 558.600 202.050 559.050 ;
        RECT 184.950 557.400 202.050 558.600 ;
        RECT 184.950 556.950 187.050 557.400 ;
        RECT 199.950 556.950 202.050 557.400 ;
        RECT 379.950 558.600 382.050 559.050 ;
        RECT 406.950 558.600 409.050 559.050 ;
        RECT 379.950 557.400 409.050 558.600 ;
        RECT 379.950 556.950 382.050 557.400 ;
        RECT 406.950 556.950 409.050 557.400 ;
        RECT 502.950 558.600 505.050 559.050 ;
        RECT 511.950 558.600 514.050 559.050 ;
        RECT 559.950 558.600 562.050 559.050 ;
        RECT 502.950 557.400 562.050 558.600 ;
        RECT 502.950 556.950 505.050 557.400 ;
        RECT 511.950 556.950 514.050 557.400 ;
        RECT 559.950 556.950 562.050 557.400 ;
        RECT 631.950 558.600 634.050 559.050 ;
        RECT 664.950 558.600 667.050 559.050 ;
        RECT 631.950 557.400 667.050 558.600 ;
        RECT 631.950 556.950 634.050 557.400 ;
        RECT 664.950 556.950 667.050 557.400 ;
        RECT 718.950 558.600 721.050 559.050 ;
        RECT 748.950 558.600 751.050 559.050 ;
        RECT 718.950 557.400 751.050 558.600 ;
        RECT 718.950 556.950 721.050 557.400 ;
        RECT 748.950 556.950 751.050 557.400 ;
        RECT 799.950 558.600 802.050 559.050 ;
        RECT 850.950 558.600 853.050 559.050 ;
        RECT 799.950 557.400 853.050 558.600 ;
        RECT 799.950 556.950 802.050 557.400 ;
        RECT 850.950 556.950 853.050 557.400 ;
        RECT 169.950 555.600 172.050 556.050 ;
        RECT 211.950 555.600 214.050 556.050 ;
        RECT 169.950 554.400 214.050 555.600 ;
        RECT 169.950 553.950 172.050 554.400 ;
        RECT 211.950 553.950 214.050 554.400 ;
        RECT 313.950 555.600 316.050 556.050 ;
        RECT 334.950 555.600 337.050 556.050 ;
        RECT 382.950 555.600 385.050 556.050 ;
        RECT 313.950 554.400 337.050 555.600 ;
        RECT 313.950 553.950 316.050 554.400 ;
        RECT 334.950 553.950 337.050 554.400 ;
        RECT 338.400 554.400 385.050 555.600 ;
        RECT 31.950 552.600 34.050 553.050 ;
        RECT 97.950 552.600 100.050 553.050 ;
        RECT 115.950 552.600 118.050 553.050 ;
        RECT 31.950 551.400 118.050 552.600 ;
        RECT 31.950 550.950 34.050 551.400 ;
        RECT 97.950 550.950 100.050 551.400 ;
        RECT 115.950 550.950 118.050 551.400 ;
        RECT 124.950 552.600 127.050 553.050 ;
        RECT 175.950 552.600 178.050 553.050 ;
        RECT 124.950 551.400 178.050 552.600 ;
        RECT 124.950 550.950 127.050 551.400 ;
        RECT 175.950 550.950 178.050 551.400 ;
        RECT 199.950 552.600 202.050 553.050 ;
        RECT 211.950 552.600 214.050 552.900 ;
        RECT 259.950 552.600 262.050 553.050 ;
        RECT 199.950 551.400 262.050 552.600 ;
        RECT 199.950 550.950 202.050 551.400 ;
        RECT 211.950 550.800 214.050 551.400 ;
        RECT 259.950 550.950 262.050 551.400 ;
        RECT 268.950 552.600 271.050 553.050 ;
        RECT 286.950 552.600 289.050 553.050 ;
        RECT 268.950 551.400 289.050 552.600 ;
        RECT 268.950 550.950 271.050 551.400 ;
        RECT 286.950 550.950 289.050 551.400 ;
        RECT 331.950 552.600 334.050 553.050 ;
        RECT 338.400 552.600 339.600 554.400 ;
        RECT 382.950 553.950 385.050 554.400 ;
        RECT 400.950 555.600 403.050 556.050 ;
        RECT 421.950 555.600 424.050 556.050 ;
        RECT 400.950 554.400 424.050 555.600 ;
        RECT 400.950 553.950 403.050 554.400 ;
        RECT 421.950 553.950 424.050 554.400 ;
        RECT 589.950 555.600 592.050 556.050 ;
        RECT 634.950 555.600 637.050 556.050 ;
        RECT 589.950 554.400 637.050 555.600 ;
        RECT 589.950 553.950 592.050 554.400 ;
        RECT 634.950 553.950 637.050 554.400 ;
        RECT 331.950 551.400 339.600 552.600 ;
        RECT 349.950 552.600 352.050 553.050 ;
        RECT 373.950 552.600 376.050 553.050 ;
        RECT 349.950 551.400 376.050 552.600 ;
        RECT 331.950 550.950 334.050 551.400 ;
        RECT 349.950 550.950 352.050 551.400 ;
        RECT 373.950 550.950 376.050 551.400 ;
        RECT 403.950 552.600 406.050 553.050 ;
        RECT 412.950 552.600 415.050 553.050 ;
        RECT 403.950 551.400 415.050 552.600 ;
        RECT 403.950 550.950 406.050 551.400 ;
        RECT 412.950 550.950 415.050 551.400 ;
        RECT 604.950 552.600 607.050 553.050 ;
        RECT 631.950 552.600 634.050 553.050 ;
        RECT 604.950 551.400 634.050 552.600 ;
        RECT 604.950 550.950 607.050 551.400 ;
        RECT 631.950 550.950 634.050 551.400 ;
        RECT 727.950 552.600 730.050 553.050 ;
        RECT 757.950 552.600 760.050 553.050 ;
        RECT 727.950 551.400 760.050 552.600 ;
        RECT 727.950 550.950 730.050 551.400 ;
        RECT 757.950 550.950 760.050 551.400 ;
        RECT 40.950 549.600 43.050 550.050 ;
        RECT 64.950 549.600 67.050 550.050 ;
        RECT 40.950 548.400 67.050 549.600 ;
        RECT 40.950 547.950 43.050 548.400 ;
        RECT 64.950 547.950 67.050 548.400 ;
        RECT 118.950 549.600 121.050 550.050 ;
        RECT 190.950 549.600 193.050 550.050 ;
        RECT 118.950 548.400 193.050 549.600 ;
        RECT 118.950 547.950 121.050 548.400 ;
        RECT 190.950 547.950 193.050 548.400 ;
        RECT 262.950 549.600 265.050 550.050 ;
        RECT 295.950 549.600 298.050 550.050 ;
        RECT 343.950 549.600 346.050 550.050 ;
        RECT 361.950 549.600 364.050 550.050 ;
        RECT 262.950 548.400 273.600 549.600 ;
        RECT 262.950 547.950 265.050 548.400 ;
        RECT 85.950 546.600 88.050 547.050 ;
        RECT 115.950 546.600 118.050 547.050 ;
        RECT 85.950 545.400 118.050 546.600 ;
        RECT 85.950 544.950 88.050 545.400 ;
        RECT 115.950 544.950 118.050 545.400 ;
        RECT 139.950 546.600 142.050 547.050 ;
        RECT 160.800 546.600 162.900 547.050 ;
        RECT 139.950 545.400 162.900 546.600 ;
        RECT 139.950 544.950 142.050 545.400 ;
        RECT 160.800 544.950 162.900 545.400 ;
        RECT 163.950 546.600 166.050 547.050 ;
        RECT 175.950 546.600 178.050 547.050 ;
        RECT 163.950 545.400 178.050 546.600 ;
        RECT 163.950 544.950 166.050 545.400 ;
        RECT 175.950 544.950 178.050 545.400 ;
        RECT 193.950 546.600 196.050 547.050 ;
        RECT 268.950 546.600 271.050 547.050 ;
        RECT 193.950 545.400 271.050 546.600 ;
        RECT 272.400 546.600 273.600 548.400 ;
        RECT 295.950 548.400 364.050 549.600 ;
        RECT 295.950 547.950 298.050 548.400 ;
        RECT 343.950 547.950 346.050 548.400 ;
        RECT 361.950 547.950 364.050 548.400 ;
        RECT 385.950 549.600 388.050 550.050 ;
        RECT 409.950 549.600 412.050 550.050 ;
        RECT 445.950 549.600 448.050 550.050 ;
        RECT 385.950 548.400 412.050 549.600 ;
        RECT 385.950 547.950 388.050 548.400 ;
        RECT 409.950 547.950 412.050 548.400 ;
        RECT 416.400 548.400 448.050 549.600 ;
        RECT 298.950 546.600 301.050 547.050 ;
        RECT 319.950 546.600 322.050 547.050 ;
        RECT 272.400 545.400 322.050 546.600 ;
        RECT 193.950 544.950 196.050 545.400 ;
        RECT 268.950 544.950 271.050 545.400 ;
        RECT 298.950 544.950 301.050 545.400 ;
        RECT 319.950 544.950 322.050 545.400 ;
        RECT 346.950 546.600 349.050 547.050 ;
        RECT 367.950 546.600 370.050 547.050 ;
        RECT 346.950 545.400 370.050 546.600 ;
        RECT 346.950 544.950 349.050 545.400 ;
        RECT 367.950 544.950 370.050 545.400 ;
        RECT 373.950 546.600 376.050 547.050 ;
        RECT 397.950 546.600 400.050 547.050 ;
        RECT 373.950 545.400 400.050 546.600 ;
        RECT 373.950 544.950 376.050 545.400 ;
        RECT 397.950 544.950 400.050 545.400 ;
        RECT 406.950 546.600 409.050 547.050 ;
        RECT 416.400 546.600 417.600 548.400 ;
        RECT 445.950 547.950 448.050 548.400 ;
        RECT 457.950 549.600 460.050 550.050 ;
        RECT 475.950 549.600 478.050 550.050 ;
        RECT 487.950 549.600 490.050 550.050 ;
        RECT 457.950 548.400 465.600 549.600 ;
        RECT 457.950 547.950 460.050 548.400 ;
        RECT 406.950 545.400 417.600 546.600 ;
        RECT 464.400 546.600 465.600 548.400 ;
        RECT 475.950 548.400 490.050 549.600 ;
        RECT 475.950 547.950 478.050 548.400 ;
        RECT 487.950 547.950 490.050 548.400 ;
        RECT 550.950 549.600 553.050 550.050 ;
        RECT 577.950 549.600 580.050 550.050 ;
        RECT 550.950 548.400 580.050 549.600 ;
        RECT 550.950 547.950 553.050 548.400 ;
        RECT 577.950 547.950 580.050 548.400 ;
        RECT 607.950 549.600 610.050 550.050 ;
        RECT 664.950 549.600 667.050 550.050 ;
        RECT 838.950 549.600 841.050 550.050 ;
        RECT 607.950 548.400 667.050 549.600 ;
        RECT 607.950 547.950 610.050 548.400 ;
        RECT 664.950 547.950 667.050 548.400 ;
        RECT 785.400 548.400 841.050 549.600 ;
        RECT 508.950 546.600 511.050 547.050 ;
        RECT 523.950 546.600 526.050 547.050 ;
        RECT 464.400 545.400 526.050 546.600 ;
        RECT 406.950 544.950 409.050 545.400 ;
        RECT 508.950 544.950 511.050 545.400 ;
        RECT 523.950 544.950 526.050 545.400 ;
        RECT 625.950 546.600 628.050 547.050 ;
        RECT 676.950 546.600 679.050 547.050 ;
        RECT 625.950 545.400 679.050 546.600 ;
        RECT 625.950 544.950 628.050 545.400 ;
        RECT 676.950 544.950 679.050 545.400 ;
        RECT 733.950 546.600 736.050 547.050 ;
        RECT 785.400 546.600 786.600 548.400 ;
        RECT 838.950 547.950 841.050 548.400 ;
        RECT 733.950 545.400 786.600 546.600 ;
        RECT 733.950 544.950 736.050 545.400 ;
        RECT 121.950 543.600 124.050 544.050 ;
        RECT 163.950 543.600 166.050 543.900 ;
        RECT 121.950 542.400 166.050 543.600 ;
        RECT 121.950 541.950 124.050 542.400 ;
        RECT 163.950 541.800 166.050 542.400 ;
        RECT 190.950 543.600 193.050 544.050 ;
        RECT 202.950 543.600 205.050 544.050 ;
        RECT 190.950 542.400 205.050 543.600 ;
        RECT 190.950 541.950 193.050 542.400 ;
        RECT 202.950 541.950 205.050 542.400 ;
        RECT 295.950 543.600 298.050 544.050 ;
        RECT 349.950 543.600 352.050 544.050 ;
        RECT 295.950 542.400 352.050 543.600 ;
        RECT 295.950 541.950 298.050 542.400 ;
        RECT 349.950 541.950 352.050 542.400 ;
        RECT 460.950 543.600 463.050 544.050 ;
        RECT 472.950 543.600 475.050 544.050 ;
        RECT 460.950 542.400 475.050 543.600 ;
        RECT 460.950 541.950 463.050 542.400 ;
        RECT 472.950 541.950 475.050 542.400 ;
        RECT 529.950 543.600 532.050 544.050 ;
        RECT 547.950 543.600 550.050 544.050 ;
        RECT 529.950 542.400 550.050 543.600 ;
        RECT 529.950 541.950 532.050 542.400 ;
        RECT 547.950 541.950 550.050 542.400 ;
        RECT 580.950 543.600 583.050 544.050 ;
        RECT 604.950 543.600 607.050 544.050 ;
        RECT 580.950 542.400 607.050 543.600 ;
        RECT 580.950 541.950 583.050 542.400 ;
        RECT 604.950 541.950 607.050 542.400 ;
        RECT 610.950 543.600 613.050 544.050 ;
        RECT 622.950 543.600 625.050 544.050 ;
        RECT 610.950 542.400 625.050 543.600 ;
        RECT 610.950 541.950 613.050 542.400 ;
        RECT 622.950 541.950 625.050 542.400 ;
        RECT 820.950 543.600 823.050 544.050 ;
        RECT 841.950 543.600 844.050 544.050 ;
        RECT 820.950 542.400 844.050 543.600 ;
        RECT 820.950 541.950 823.050 542.400 ;
        RECT 841.950 541.950 844.050 542.400 ;
        RECT 1.950 540.600 4.050 541.050 ;
        RECT 118.950 540.600 121.050 541.050 ;
        RECT 1.950 539.400 121.050 540.600 ;
        RECT 1.950 538.950 4.050 539.400 ;
        RECT 118.950 538.950 121.050 539.400 ;
        RECT 124.950 540.600 127.050 541.050 ;
        RECT 157.950 540.600 160.050 541.050 ;
        RECT 217.950 540.600 220.050 541.050 ;
        RECT 124.950 539.400 220.050 540.600 ;
        RECT 124.950 538.950 127.050 539.400 ;
        RECT 157.950 538.950 160.050 539.400 ;
        RECT 217.950 538.950 220.050 539.400 ;
        RECT 226.950 540.600 229.050 541.050 ;
        RECT 250.950 540.600 253.050 541.050 ;
        RECT 226.950 539.400 253.050 540.600 ;
        RECT 226.950 538.950 229.050 539.400 ;
        RECT 250.950 538.950 253.050 539.400 ;
        RECT 397.950 540.600 400.050 541.050 ;
        RECT 427.950 540.600 430.050 541.050 ;
        RECT 397.950 539.400 430.050 540.600 ;
        RECT 397.950 538.950 400.050 539.400 ;
        RECT 427.950 538.950 430.050 539.400 ;
        RECT 463.950 540.600 466.050 541.050 ;
        RECT 559.950 540.600 562.050 541.050 ;
        RECT 463.950 539.400 562.050 540.600 ;
        RECT 463.950 538.950 466.050 539.400 ;
        RECT 559.950 538.950 562.050 539.400 ;
        RECT 631.950 540.600 634.050 541.050 ;
        RECT 727.950 540.600 730.050 541.050 ;
        RECT 631.950 539.400 730.050 540.600 ;
        RECT 631.950 538.950 634.050 539.400 ;
        RECT 727.950 538.950 730.050 539.400 ;
        RECT 163.950 537.600 166.050 538.050 ;
        RECT 193.950 537.600 196.050 538.050 ;
        RECT 163.950 536.400 196.050 537.600 ;
        RECT 163.950 535.950 166.050 536.400 ;
        RECT 193.950 535.950 196.050 536.400 ;
        RECT 226.950 537.600 229.050 537.900 ;
        RECT 238.950 537.600 241.050 538.050 ;
        RECT 256.950 537.600 259.050 538.050 ;
        RECT 226.950 536.400 241.050 537.600 ;
        RECT 226.950 535.800 229.050 536.400 ;
        RECT 238.950 535.950 241.050 536.400 ;
        RECT 251.400 536.400 259.050 537.600 ;
        RECT 76.950 534.600 79.050 535.050 ;
        RECT 109.950 534.600 112.050 535.050 ;
        RECT 76.950 533.400 112.050 534.600 ;
        RECT 76.950 532.950 79.050 533.400 ;
        RECT 109.950 532.950 112.050 533.400 ;
        RECT 115.950 534.600 118.050 535.050 ;
        RECT 130.950 534.600 133.050 535.050 ;
        RECT 115.950 533.400 133.050 534.600 ;
        RECT 115.950 532.950 118.050 533.400 ;
        RECT 130.950 532.950 133.050 533.400 ;
        RECT 151.950 534.600 154.050 535.050 ;
        RECT 169.950 534.600 172.050 535.050 ;
        RECT 178.950 534.600 181.050 535.050 ;
        RECT 151.950 533.400 181.050 534.600 ;
        RECT 151.950 532.950 154.050 533.400 ;
        RECT 169.950 532.950 172.050 533.400 ;
        RECT 178.950 532.950 181.050 533.400 ;
        RECT 202.950 534.600 205.050 535.050 ;
        RECT 220.950 534.600 223.050 535.050 ;
        RECT 251.400 534.600 252.600 536.400 ;
        RECT 256.950 535.950 259.050 536.400 ;
        RECT 316.950 537.600 319.050 538.050 ;
        RECT 346.950 537.600 349.050 538.050 ;
        RECT 316.950 536.400 349.050 537.600 ;
        RECT 316.950 535.950 319.050 536.400 ;
        RECT 346.950 535.950 349.050 536.400 ;
        RECT 361.950 537.600 364.050 538.050 ;
        RECT 403.950 537.600 406.050 538.050 ;
        RECT 361.950 536.400 406.050 537.600 ;
        RECT 361.950 535.950 364.050 536.400 ;
        RECT 403.950 535.950 406.050 536.400 ;
        RECT 430.950 537.600 433.050 538.050 ;
        RECT 457.950 537.600 460.050 538.050 ;
        RECT 430.950 536.400 460.050 537.600 ;
        RECT 430.950 535.950 433.050 536.400 ;
        RECT 457.950 535.950 460.050 536.400 ;
        RECT 475.950 537.600 478.050 538.050 ;
        RECT 490.800 537.600 492.900 538.050 ;
        RECT 475.950 536.400 492.900 537.600 ;
        RECT 560.400 537.600 561.600 538.950 ;
        RECT 580.950 537.600 583.050 538.050 ;
        RECT 560.400 536.400 583.050 537.600 ;
        RECT 475.950 535.950 478.050 536.400 ;
        RECT 490.800 535.950 492.900 536.400 ;
        RECT 580.950 535.950 583.050 536.400 ;
        RECT 736.950 537.600 739.050 538.050 ;
        RECT 781.950 537.600 784.050 538.050 ;
        RECT 736.950 536.400 784.050 537.600 ;
        RECT 736.950 535.950 739.050 536.400 ;
        RECT 781.950 535.950 784.050 536.400 ;
        RECT 829.950 537.600 832.050 538.050 ;
        RECT 835.950 537.600 838.050 538.050 ;
        RECT 829.950 536.400 838.050 537.600 ;
        RECT 829.950 535.950 832.050 536.400 ;
        RECT 835.950 535.950 838.050 536.400 ;
        RECT 202.950 533.400 252.600 534.600 ;
        RECT 271.950 534.600 274.050 535.050 ;
        RECT 280.950 534.600 283.050 535.050 ;
        RECT 349.950 534.600 352.050 535.050 ;
        RECT 391.800 534.600 393.900 535.050 ;
        RECT 271.950 533.400 283.050 534.600 ;
        RECT 202.950 532.950 205.050 533.400 ;
        RECT 220.950 532.950 223.050 533.400 ;
        RECT 271.950 532.950 274.050 533.400 ;
        RECT 280.950 532.950 283.050 533.400 ;
        RECT 332.400 533.400 393.900 534.600 ;
        RECT 332.400 532.050 333.600 533.400 ;
        RECT 349.950 532.950 352.050 533.400 ;
        RECT 391.800 532.950 393.900 533.400 ;
        RECT 427.950 534.600 430.050 535.050 ;
        RECT 532.950 534.600 535.050 535.050 ;
        RECT 427.950 533.400 535.050 534.600 ;
        RECT 427.950 532.950 430.050 533.400 ;
        RECT 532.950 532.950 535.050 533.400 ;
        RECT 853.950 534.600 856.050 535.050 ;
        RECT 859.950 534.600 862.050 535.050 ;
        RECT 853.950 533.400 862.050 534.600 ;
        RECT 853.950 532.950 856.050 533.400 ;
        RECT 859.950 532.950 862.050 533.400 ;
        RECT 19.950 531.600 22.050 532.050 ;
        RECT 34.950 531.600 37.050 532.050 ;
        RECT 19.950 530.400 37.050 531.600 ;
        RECT 19.950 529.950 22.050 530.400 ;
        RECT 34.950 529.950 37.050 530.400 ;
        RECT 136.950 531.600 139.050 532.050 ;
        RECT 142.950 531.600 145.050 532.050 ;
        RECT 136.950 530.400 145.050 531.600 ;
        RECT 136.950 529.950 139.050 530.400 ;
        RECT 142.950 529.950 145.050 530.400 ;
        RECT 172.950 531.600 177.000 532.050 ;
        RECT 190.950 531.600 193.050 532.050 ;
        RECT 172.950 529.950 177.600 531.600 ;
        RECT 31.950 526.950 34.050 529.050 ;
        RECT 88.950 528.600 91.050 529.050 ;
        RECT 97.950 528.600 100.050 529.050 ;
        RECT 88.950 527.400 100.050 528.600 ;
        RECT 88.950 526.950 91.050 527.400 ;
        RECT 97.950 526.950 100.050 527.400 ;
        RECT 103.950 528.600 106.050 529.050 ;
        RECT 118.950 528.600 121.050 529.050 ;
        RECT 103.950 527.400 121.050 528.600 ;
        RECT 103.950 526.950 106.050 527.400 ;
        RECT 118.950 526.950 121.050 527.400 ;
        RECT 32.400 522.750 33.600 526.950 ;
        RECT 124.950 526.800 127.050 528.900 ;
        RECT 125.400 523.050 126.600 526.800 ;
        RECT 130.950 525.600 133.050 529.050 ;
        RECT 130.950 525.000 138.600 525.600 ;
        RECT 131.400 524.400 138.600 525.000 ;
        RECT 16.950 522.600 19.050 522.750 ;
        RECT 31.950 522.600 34.050 522.750 ;
        RECT 16.950 521.400 34.050 522.600 ;
        RECT 16.950 520.650 19.050 521.400 ;
        RECT 31.950 520.650 34.050 521.400 ;
        RECT 37.950 522.600 40.050 522.750 ;
        RECT 43.950 522.600 46.050 523.050 ;
        RECT 37.950 521.400 46.050 522.600 ;
        RECT 37.950 520.650 40.050 521.400 ;
        RECT 43.950 520.950 46.050 521.400 ;
        RECT 64.950 522.600 67.050 523.050 ;
        RECT 73.950 522.600 76.050 522.750 ;
        RECT 64.950 521.400 76.050 522.600 ;
        RECT 64.950 520.950 67.050 521.400 ;
        RECT 73.950 520.650 76.050 521.400 ;
        RECT 100.950 522.600 103.050 522.750 ;
        RECT 121.950 522.600 124.050 522.750 ;
        RECT 100.950 521.400 124.050 522.600 ;
        RECT 125.400 521.400 130.050 523.050 ;
        RECT 137.400 522.600 138.600 524.400 ;
        RECT 154.950 522.600 157.050 522.900 ;
        RECT 176.400 522.750 177.600 529.950 ;
        RECT 182.400 530.400 193.050 531.600 ;
        RECT 182.400 522.750 183.600 530.400 ;
        RECT 190.950 529.950 193.050 530.400 ;
        RECT 265.950 529.950 268.050 532.050 ;
        RECT 328.950 530.400 333.600 532.050 ;
        RECT 328.950 529.950 333.000 530.400 ;
        RECT 376.950 529.950 379.050 532.050 ;
        RECT 409.950 531.600 412.050 531.900 ;
        RECT 421.950 531.600 424.050 532.050 ;
        RECT 409.950 530.400 424.050 531.600 ;
        RECT 187.950 528.600 190.050 529.050 ;
        RECT 193.950 528.600 196.050 529.050 ;
        RECT 187.950 527.400 196.050 528.600 ;
        RECT 187.950 526.950 190.050 527.400 ;
        RECT 193.950 526.950 196.050 527.400 ;
        RECT 211.950 526.950 214.050 529.050 ;
        RECT 217.950 526.950 220.050 529.050 ;
        RECT 238.800 528.000 240.900 529.050 ;
        RECT 238.800 526.950 241.050 528.000 ;
        RECT 241.950 526.950 244.050 529.050 ;
        RECT 212.400 523.050 213.600 526.950 ;
        RECT 137.400 521.400 157.050 522.600 ;
        RECT 100.950 520.650 103.050 521.400 ;
        RECT 121.950 520.650 124.050 521.400 ;
        RECT 126.000 520.950 130.050 521.400 ;
        RECT 154.950 520.800 157.050 521.400 ;
        RECT 175.950 520.650 178.050 522.750 ;
        RECT 181.950 520.650 184.050 522.750 ;
        RECT 211.950 520.950 214.050 523.050 ;
        RECT 218.400 522.750 219.600 526.950 ;
        RECT 238.950 525.600 241.050 526.950 ;
        RECT 224.400 525.000 241.050 525.600 ;
        RECT 223.950 524.400 240.450 525.000 ;
        RECT 217.950 520.650 220.050 522.750 ;
        RECT 223.950 520.950 226.050 524.400 ;
        RECT 242.400 522.600 243.600 526.950 ;
        RECT 247.950 525.600 250.050 529.050 ;
        RECT 247.950 525.000 255.600 525.600 ;
        RECT 248.400 524.400 255.600 525.000 ;
        RECT 239.400 522.000 243.600 522.600 ;
        RECT 238.950 521.400 243.600 522.000 ;
        RECT 254.400 522.600 255.600 524.400 ;
        RECT 266.400 522.900 267.600 529.950 ;
        RECT 268.950 525.600 271.050 529.050 ;
        RECT 292.950 526.950 295.050 529.050 ;
        RECT 268.950 525.000 282.600 525.600 ;
        RECT 269.400 524.400 282.600 525.000 ;
        RECT 259.950 522.600 262.050 522.900 ;
        RECT 254.400 521.400 262.050 522.600 ;
        RECT 43.950 519.600 46.050 519.900 ;
        RECT 52.950 519.600 55.050 520.050 ;
        RECT 43.950 518.400 55.050 519.600 ;
        RECT 43.950 517.800 46.050 518.400 ;
        RECT 52.950 517.950 55.050 518.400 ;
        RECT 91.950 519.600 94.050 520.050 ;
        RECT 133.950 519.600 136.050 520.050 ;
        RECT 166.950 519.600 169.050 520.050 ;
        RECT 91.950 518.400 169.050 519.600 ;
        RECT 91.950 517.950 94.050 518.400 ;
        RECT 133.950 517.950 136.050 518.400 ;
        RECT 166.950 517.950 169.050 518.400 ;
        RECT 238.950 517.950 241.050 521.400 ;
        RECT 259.950 520.800 262.050 521.400 ;
        RECT 265.950 520.800 268.050 522.900 ;
        RECT 281.400 522.600 282.600 524.400 ;
        RECT 293.400 523.050 294.600 526.950 ;
        RECT 298.950 525.600 301.050 529.050 ;
        RECT 296.400 525.000 301.050 525.600 ;
        RECT 296.400 524.400 300.600 525.000 ;
        RECT 289.800 522.600 291.900 523.050 ;
        RECT 281.400 521.400 291.900 522.600 ;
        RECT 289.800 520.950 291.900 521.400 ;
        RECT 292.950 520.950 295.050 523.050 ;
        RECT 296.400 519.600 297.600 524.400 ;
        RECT 298.950 522.600 301.050 522.750 ;
        RECT 313.950 522.600 316.050 522.900 ;
        RECT 340.950 522.600 343.050 522.750 ;
        RECT 298.950 521.400 316.050 522.600 ;
        RECT 335.400 522.000 343.050 522.600 ;
        RECT 298.950 520.650 301.050 521.400 ;
        RECT 313.950 520.800 316.050 521.400 ;
        RECT 334.950 521.400 343.050 522.000 ;
        RECT 307.950 519.600 310.050 520.050 ;
        RECT 296.400 518.400 310.050 519.600 ;
        RECT 307.950 517.950 310.050 518.400 ;
        RECT 334.950 517.950 337.050 521.400 ;
        RECT 340.950 520.650 343.050 521.400 ;
        RECT 358.950 522.600 361.050 522.750 ;
        RECT 367.950 522.600 370.050 523.050 ;
        RECT 377.400 522.900 378.600 529.950 ;
        RECT 409.950 529.800 412.050 530.400 ;
        RECT 421.950 529.950 424.050 530.400 ;
        RECT 436.950 531.600 439.050 532.050 ;
        RECT 445.950 531.600 448.050 532.050 ;
        RECT 463.950 531.600 466.050 532.050 ;
        RECT 436.950 530.400 466.050 531.600 ;
        RECT 436.950 529.950 439.050 530.400 ;
        RECT 445.950 529.950 448.050 530.400 ;
        RECT 463.950 529.950 466.050 530.400 ;
        RECT 667.950 531.600 670.050 532.050 ;
        RECT 703.950 531.600 706.050 532.050 ;
        RECT 718.950 531.600 721.050 532.050 ;
        RECT 769.950 531.600 772.050 532.050 ;
        RECT 667.950 530.400 721.050 531.600 ;
        RECT 667.950 529.950 670.050 530.400 ;
        RECT 703.950 529.950 706.050 530.400 ;
        RECT 718.950 529.950 721.050 530.400 ;
        RECT 743.400 530.400 772.050 531.600 ;
        RECT 384.000 528.600 388.050 529.050 ;
        RECT 383.400 526.950 388.050 528.600 ;
        RECT 383.400 522.900 384.600 526.950 ;
        RECT 400.950 525.600 403.050 529.050 ;
        RECT 418.950 527.100 421.050 529.200 ;
        RECT 454.950 528.600 457.050 529.200 ;
        RECT 474.000 528.600 478.050 529.050 ;
        RECT 449.400 527.400 457.050 528.600 ;
        RECT 398.400 525.000 403.050 525.600 ;
        RECT 419.400 525.600 420.600 527.100 ;
        RECT 398.400 524.400 402.600 525.000 ;
        RECT 419.400 524.400 432.600 525.600 ;
        RECT 358.950 521.400 370.050 522.600 ;
        RECT 358.950 520.650 361.050 521.400 ;
        RECT 367.950 520.950 370.050 521.400 ;
        RECT 376.950 520.800 379.050 522.900 ;
        RECT 382.950 520.800 385.050 522.900 ;
        RECT 394.950 522.600 397.050 522.750 ;
        RECT 398.400 522.600 399.600 524.400 ;
        RECT 394.950 521.400 399.600 522.600 ;
        RECT 409.950 522.600 412.050 522.900 ;
        RECT 424.950 522.600 427.050 523.050 ;
        RECT 409.950 521.400 427.050 522.600 ;
        RECT 431.400 522.600 432.600 524.400 ;
        RECT 433.950 522.600 436.050 522.750 ;
        RECT 431.400 521.400 436.050 522.600 ;
        RECT 394.950 520.650 397.050 521.400 ;
        RECT 409.950 520.800 412.050 521.400 ;
        RECT 424.950 520.950 427.050 521.400 ;
        RECT 433.950 520.650 436.050 521.400 ;
        RECT 442.950 519.600 445.050 520.050 ;
        RECT 449.400 519.600 450.600 527.400 ;
        RECT 454.950 527.100 457.050 527.400 ;
        RECT 473.400 526.950 478.050 528.600 ;
        RECT 496.950 526.950 499.050 529.050 ;
        RECT 514.950 527.100 517.050 529.200 ;
        RECT 473.400 522.900 474.600 526.950 ;
        RECT 472.950 520.800 475.050 522.900 ;
        RECT 497.400 522.600 498.600 526.950 ;
        RECT 515.400 525.600 516.600 527.100 ;
        RECT 529.950 526.950 532.050 529.050 ;
        RECT 538.950 528.750 541.050 529.200 ;
        RECT 553.950 528.750 556.050 529.200 ;
        RECT 538.950 527.550 556.050 528.750 ;
        RECT 571.950 528.600 574.050 529.200 ;
        RECT 610.950 528.600 613.050 529.050 ;
        RECT 538.950 527.100 541.050 527.550 ;
        RECT 553.950 527.100 556.050 527.550 ;
        RECT 557.400 527.400 574.050 528.600 ;
        RECT 515.400 525.000 519.600 525.600 ;
        RECT 515.400 524.400 520.050 525.000 ;
        RECT 502.950 522.600 505.050 523.050 ;
        RECT 497.400 521.400 505.050 522.600 ;
        RECT 502.950 520.950 505.050 521.400 ;
        RECT 517.950 520.950 520.050 524.400 ;
        RECT 530.400 522.750 531.600 526.950 ;
        RECT 541.950 525.600 544.050 526.050 ;
        RECT 557.400 525.600 558.600 527.400 ;
        RECT 571.950 527.100 574.050 527.400 ;
        RECT 590.400 527.400 613.050 528.600 ;
        RECT 541.950 524.400 558.600 525.600 ;
        RECT 541.950 523.950 544.050 524.400 ;
        RECT 529.950 520.650 532.050 522.750 ;
        RECT 574.950 522.600 577.050 523.050 ;
        RECT 590.400 522.900 591.600 527.400 ;
        RECT 610.950 526.950 613.050 527.400 ;
        RECT 616.950 527.100 619.050 529.200 ;
        RECT 649.950 528.600 652.050 528.900 ;
        RECT 655.950 528.600 658.050 529.050 ;
        RECT 649.950 527.400 658.050 528.600 ;
        RECT 554.400 521.400 577.050 522.600 ;
        RECT 442.950 518.400 450.600 519.600 ;
        RECT 538.950 519.600 541.050 519.900 ;
        RECT 554.400 519.600 555.600 521.400 ;
        RECT 574.950 520.950 577.050 521.400 ;
        RECT 589.950 520.800 592.050 522.900 ;
        RECT 617.400 522.600 618.600 527.100 ;
        RECT 649.950 526.800 652.050 527.400 ;
        RECT 655.950 526.950 658.050 527.400 ;
        RECT 664.950 528.750 667.050 529.200 ;
        RECT 676.950 528.750 679.050 529.200 ;
        RECT 664.950 527.550 679.050 528.750 ;
        RECT 664.950 527.100 667.050 527.550 ;
        RECT 676.950 527.100 679.050 527.550 ;
        RECT 682.950 528.600 685.050 529.200 ;
        RECT 688.800 528.600 690.900 529.050 ;
        RECT 682.950 527.400 690.900 528.600 ;
        RECT 682.950 527.100 685.050 527.400 ;
        RECT 688.800 526.950 690.900 527.400 ;
        RECT 691.950 528.750 694.050 529.200 ;
        RECT 697.950 528.750 700.050 529.200 ;
        RECT 691.950 527.550 700.050 528.750 ;
        RECT 691.950 527.100 694.050 527.550 ;
        RECT 697.950 527.100 700.050 527.550 ;
        RECT 724.950 525.600 727.050 529.050 ;
        RECT 739.950 525.600 742.050 526.050 ;
        RECT 724.950 525.000 742.050 525.600 ;
        RECT 725.400 524.400 742.050 525.000 ;
        RECT 658.950 522.600 661.050 522.750 ;
        RECT 679.950 522.600 682.050 522.900 ;
        RECT 691.950 522.600 694.050 523.050 ;
        RECT 608.400 521.400 618.600 522.600 ;
        RECT 653.400 522.000 678.600 522.600 ;
        RECT 652.950 521.400 678.600 522.000 ;
        RECT 608.400 520.050 609.600 521.400 ;
        RECT 538.950 518.400 555.600 519.600 ;
        RECT 559.950 519.600 562.050 520.050 ;
        RECT 595.950 519.600 598.050 520.050 ;
        RECT 559.950 518.400 598.050 519.600 ;
        RECT 442.950 517.950 445.050 518.400 ;
        RECT 538.950 517.800 541.050 518.400 ;
        RECT 559.950 517.950 562.050 518.400 ;
        RECT 595.950 517.950 598.050 518.400 ;
        RECT 604.950 518.400 609.600 520.050 ;
        RECT 604.950 517.950 609.000 518.400 ;
        RECT 652.950 517.950 655.050 521.400 ;
        RECT 658.950 520.650 661.050 521.400 ;
        RECT 677.400 519.600 678.600 521.400 ;
        RECT 679.950 521.400 694.050 522.600 ;
        RECT 679.950 520.800 682.050 521.400 ;
        RECT 691.950 520.950 694.050 521.400 ;
        RECT 706.950 522.600 709.050 522.900 ;
        RECT 715.950 522.600 718.050 522.750 ;
        RECT 706.950 521.400 718.050 522.600 ;
        RECT 706.950 520.800 709.050 521.400 ;
        RECT 682.950 519.600 685.050 520.050 ;
        RECT 677.400 518.400 685.050 519.600 ;
        RECT 682.950 517.950 685.050 518.400 ;
        RECT 694.950 519.600 697.050 520.050 ;
        RECT 707.400 519.600 708.600 520.800 ;
        RECT 715.950 520.650 718.050 521.400 ;
        RECT 694.950 518.400 708.600 519.600 ;
        RECT 694.950 517.950 697.050 518.400 ;
        RECT 88.950 516.600 91.050 517.050 ;
        RECT 100.950 516.600 103.050 517.050 ;
        RECT 88.950 515.400 103.050 516.600 ;
        RECT 88.950 514.950 91.050 515.400 ;
        RECT 100.950 514.950 103.050 515.400 ;
        RECT 118.950 516.600 121.050 517.050 ;
        RECT 127.950 516.600 130.050 517.050 ;
        RECT 118.950 515.400 130.050 516.600 ;
        RECT 118.950 514.950 121.050 515.400 ;
        RECT 127.950 514.950 130.050 515.400 ;
        RECT 175.950 516.600 178.050 517.050 ;
        RECT 199.950 516.600 202.050 517.050 ;
        RECT 175.950 515.400 202.050 516.600 ;
        RECT 175.950 514.950 178.050 515.400 ;
        RECT 199.950 514.950 202.050 515.400 ;
        RECT 241.950 516.600 244.050 517.050 ;
        RECT 280.950 516.600 283.050 517.050 ;
        RECT 241.950 515.400 283.050 516.600 ;
        RECT 241.950 514.950 244.050 515.400 ;
        RECT 280.950 514.950 283.050 515.400 ;
        RECT 289.950 516.600 292.050 517.050 ;
        RECT 319.950 516.600 322.050 517.050 ;
        RECT 289.950 515.400 322.050 516.600 ;
        RECT 289.950 514.950 292.050 515.400 ;
        RECT 319.950 514.950 322.050 515.400 ;
        RECT 331.950 516.600 334.050 517.050 ;
        RECT 355.950 516.600 358.050 517.050 ;
        RECT 331.950 515.400 358.050 516.600 ;
        RECT 331.950 514.950 334.050 515.400 ;
        RECT 355.950 514.950 358.050 515.400 ;
        RECT 403.950 516.600 406.050 517.050 ;
        RECT 412.950 516.600 415.050 517.050 ;
        RECT 403.950 515.400 415.050 516.600 ;
        RECT 403.950 514.950 406.050 515.400 ;
        RECT 412.950 514.950 415.050 515.400 ;
        RECT 493.950 516.600 496.050 517.050 ;
        RECT 517.950 516.600 520.050 517.050 ;
        RECT 493.950 515.400 520.050 516.600 ;
        RECT 493.950 514.950 496.050 515.400 ;
        RECT 517.950 514.950 520.050 515.400 ;
        RECT 700.950 516.600 703.050 517.050 ;
        RECT 725.400 516.600 726.600 524.400 ;
        RECT 739.950 523.950 742.050 524.400 ;
        RECT 727.950 522.600 730.050 522.750 ;
        RECT 743.400 522.600 744.600 530.400 ;
        RECT 769.950 529.950 772.050 530.400 ;
        RECT 760.950 528.600 763.050 529.050 ;
        RECT 772.950 528.600 775.050 529.050 ;
        RECT 760.950 527.400 775.050 528.600 ;
        RECT 760.950 526.950 763.050 527.400 ;
        RECT 772.950 526.950 775.050 527.400 ;
        RECT 793.950 528.600 796.050 529.050 ;
        RECT 802.950 528.600 805.050 529.200 ;
        RECT 832.950 528.600 835.050 529.050 ;
        RECT 793.950 527.400 805.050 528.600 ;
        RECT 793.950 526.950 796.050 527.400 ;
        RECT 802.950 527.100 805.050 527.400 ;
        RECT 818.400 527.400 835.050 528.600 ;
        RECT 757.950 525.600 760.050 526.050 ;
        RECT 757.950 524.400 768.600 525.600 ;
        RECT 757.950 523.950 760.050 524.400 ;
        RECT 767.400 522.900 768.600 524.400 ;
        RECT 727.950 521.400 744.600 522.600 ;
        RECT 727.950 520.650 730.050 521.400 ;
        RECT 766.950 520.800 769.050 522.900 ;
        RECT 805.950 522.600 808.050 523.050 ;
        RECT 814.950 522.600 817.050 526.050 ;
        RECT 805.950 522.000 817.050 522.600 ;
        RECT 805.950 521.400 816.600 522.000 ;
        RECT 805.950 520.950 808.050 521.400 ;
        RECT 760.950 519.600 763.050 520.050 ;
        RECT 799.950 519.600 802.050 520.050 ;
        RECT 760.950 518.400 802.050 519.600 ;
        RECT 760.950 517.950 763.050 518.400 ;
        RECT 799.950 517.950 802.050 518.400 ;
        RECT 811.950 519.600 814.050 520.050 ;
        RECT 818.400 519.600 819.600 527.400 ;
        RECT 832.950 526.950 835.050 527.400 ;
        RECT 841.950 526.950 844.050 529.050 ;
        RECT 847.950 528.600 850.050 529.050 ;
        RECT 856.950 528.600 859.050 528.900 ;
        RECT 847.950 527.400 859.050 528.600 ;
        RECT 847.950 526.950 850.050 527.400 ;
        RECT 842.400 520.050 843.600 526.950 ;
        RECT 856.950 526.800 859.050 527.400 ;
        RECT 811.950 518.400 819.600 519.600 ;
        RECT 811.950 517.950 814.050 518.400 ;
        RECT 841.950 517.950 844.050 520.050 ;
        RECT 850.950 519.600 853.050 520.050 ;
        RECT 856.950 519.600 859.050 520.050 ;
        RECT 850.950 518.400 859.050 519.600 ;
        RECT 850.950 517.950 853.050 518.400 ;
        RECT 856.950 517.950 859.050 518.400 ;
        RECT 700.950 515.400 726.600 516.600 ;
        RECT 700.950 514.950 703.050 515.400 ;
        RECT 85.950 513.600 88.050 514.050 ;
        RECT 119.400 513.600 120.600 514.950 ;
        RECT 85.950 512.400 120.600 513.600 ;
        RECT 130.950 513.600 133.050 514.050 ;
        RECT 142.950 513.600 145.050 514.050 ;
        RECT 130.950 512.400 145.050 513.600 ;
        RECT 85.950 511.950 88.050 512.400 ;
        RECT 130.950 511.950 133.050 512.400 ;
        RECT 142.950 511.950 145.050 512.400 ;
        RECT 190.950 513.600 193.050 514.050 ;
        RECT 208.950 513.600 211.050 514.050 ;
        RECT 190.950 512.400 211.050 513.600 ;
        RECT 190.950 511.950 193.050 512.400 ;
        RECT 208.950 511.950 211.050 512.400 ;
        RECT 250.950 513.600 253.050 514.050 ;
        RECT 283.800 513.600 285.900 514.050 ;
        RECT 250.950 512.400 285.900 513.600 ;
        RECT 250.950 511.950 253.050 512.400 ;
        RECT 283.800 511.950 285.900 512.400 ;
        RECT 286.950 513.600 289.050 514.050 ;
        RECT 316.950 513.600 319.050 514.050 ;
        RECT 286.950 512.400 319.050 513.600 ;
        RECT 286.950 511.950 289.050 512.400 ;
        RECT 316.950 511.950 319.050 512.400 ;
        RECT 346.950 513.600 349.050 514.050 ;
        RECT 394.950 513.600 397.050 514.050 ;
        RECT 346.950 512.400 397.050 513.600 ;
        RECT 346.950 511.950 349.050 512.400 ;
        RECT 394.950 511.950 397.050 512.400 ;
        RECT 415.950 513.600 418.050 514.050 ;
        RECT 442.950 513.600 445.050 514.050 ;
        RECT 415.950 512.400 445.050 513.600 ;
        RECT 415.950 511.950 418.050 512.400 ;
        RECT 442.950 511.950 445.050 512.400 ;
        RECT 553.950 513.600 556.050 514.050 ;
        RECT 577.950 513.600 580.050 514.050 ;
        RECT 670.950 513.600 673.050 514.050 ;
        RECT 553.950 512.400 580.050 513.600 ;
        RECT 584.400 513.000 673.050 513.600 ;
        RECT 553.950 511.950 556.050 512.400 ;
        RECT 577.950 511.950 580.050 512.400 ;
        RECT 583.950 512.400 673.050 513.000 ;
        RECT 70.950 510.600 73.050 511.050 ;
        RECT 82.950 510.600 85.050 511.050 ;
        RECT 70.950 509.400 85.050 510.600 ;
        RECT 70.950 508.950 73.050 509.400 ;
        RECT 82.950 508.950 85.050 509.400 ;
        RECT 109.950 510.600 112.050 511.050 ;
        RECT 115.950 510.600 118.050 511.050 ;
        RECT 109.950 509.400 118.050 510.600 ;
        RECT 109.950 508.950 112.050 509.400 ;
        RECT 115.950 508.950 118.050 509.400 ;
        RECT 202.950 510.600 205.050 511.050 ;
        RECT 268.950 510.600 271.050 511.050 ;
        RECT 202.950 509.400 252.600 510.600 ;
        RECT 202.950 508.950 205.050 509.400 ;
        RECT 67.950 507.600 70.050 508.050 ;
        RECT 103.950 507.600 106.050 508.050 ;
        RECT 67.950 506.400 106.050 507.600 ;
        RECT 67.950 505.950 70.050 506.400 ;
        RECT 103.950 505.950 106.050 506.400 ;
        RECT 154.950 507.600 157.050 508.050 ;
        RECT 160.800 507.600 162.900 508.050 ;
        RECT 223.950 507.600 226.050 508.050 ;
        RECT 154.950 506.400 162.900 507.600 ;
        RECT 154.950 505.950 157.050 506.400 ;
        RECT 160.800 505.950 162.900 506.400 ;
        RECT 200.400 506.400 226.050 507.600 ;
        RECT 251.400 507.600 252.600 509.400 ;
        RECT 257.400 509.400 271.050 510.600 ;
        RECT 257.400 507.600 258.600 509.400 ;
        RECT 268.950 508.950 271.050 509.400 ;
        RECT 319.950 510.600 322.050 511.050 ;
        RECT 328.950 510.600 331.050 511.050 ;
        RECT 319.950 509.400 331.050 510.600 ;
        RECT 319.950 508.950 322.050 509.400 ;
        RECT 328.950 508.950 331.050 509.400 ;
        RECT 451.950 510.600 454.050 511.050 ;
        RECT 460.950 510.600 463.050 511.050 ;
        RECT 451.950 509.400 463.050 510.600 ;
        RECT 451.950 508.950 454.050 509.400 ;
        RECT 460.950 508.950 463.050 509.400 ;
        RECT 517.950 510.600 520.050 511.050 ;
        RECT 541.950 510.600 544.050 511.050 ;
        RECT 517.950 509.400 544.050 510.600 ;
        RECT 517.950 508.950 520.050 509.400 ;
        RECT 541.950 508.950 544.050 509.400 ;
        RECT 550.950 510.600 553.050 511.050 ;
        RECT 562.950 510.600 565.050 511.050 ;
        RECT 550.950 509.400 565.050 510.600 ;
        RECT 550.950 508.950 553.050 509.400 ;
        RECT 562.950 508.950 565.050 509.400 ;
        RECT 583.950 508.950 586.050 512.400 ;
        RECT 670.950 511.950 673.050 512.400 ;
        RECT 808.950 513.600 811.050 514.050 ;
        RECT 817.950 513.600 820.050 514.050 ;
        RECT 844.950 513.600 847.050 514.050 ;
        RECT 808.950 512.400 847.050 513.600 ;
        RECT 808.950 511.950 811.050 512.400 ;
        RECT 817.950 511.950 820.050 512.400 ;
        RECT 844.950 511.950 847.050 512.400 ;
        RECT 607.950 510.600 610.050 511.050 ;
        RECT 667.950 510.600 670.050 511.050 ;
        RECT 607.950 509.400 670.050 510.600 ;
        RECT 607.950 508.950 610.050 509.400 ;
        RECT 667.950 508.950 670.050 509.400 ;
        RECT 694.950 510.600 697.050 511.050 ;
        RECT 721.950 510.600 724.050 511.050 ;
        RECT 694.950 509.400 724.050 510.600 ;
        RECT 694.950 508.950 697.050 509.400 ;
        RECT 721.950 508.950 724.050 509.400 ;
        RECT 742.950 510.600 745.050 511.050 ;
        RECT 853.950 510.600 856.050 511.050 ;
        RECT 742.950 509.400 856.050 510.600 ;
        RECT 742.950 508.950 745.050 509.400 ;
        RECT 853.950 508.950 856.050 509.400 ;
        RECT 251.400 506.400 258.600 507.600 ;
        RECT 259.950 507.600 262.050 508.050 ;
        RECT 274.950 507.600 277.050 508.050 ;
        RECT 259.950 506.400 277.050 507.600 ;
        RECT 200.400 505.050 201.600 506.400 ;
        RECT 223.950 505.950 226.050 506.400 ;
        RECT 259.950 505.950 262.050 506.400 ;
        RECT 274.950 505.950 277.050 506.400 ;
        RECT 307.950 507.600 310.050 508.050 ;
        RECT 316.950 507.600 319.050 508.050 ;
        RECT 307.950 506.400 319.050 507.600 ;
        RECT 307.950 505.950 310.050 506.400 ;
        RECT 316.950 505.950 319.050 506.400 ;
        RECT 337.950 507.600 340.050 508.050 ;
        RECT 367.950 507.600 370.050 508.050 ;
        RECT 337.950 506.400 370.050 507.600 ;
        RECT 337.950 505.950 340.050 506.400 ;
        RECT 367.950 505.950 370.050 506.400 ;
        RECT 391.950 507.600 394.050 508.050 ;
        RECT 409.950 507.600 412.050 508.050 ;
        RECT 478.950 507.600 481.050 508.050 ;
        RECT 391.950 506.400 412.050 507.600 ;
        RECT 391.950 505.950 394.050 506.400 ;
        RECT 409.950 505.950 412.050 506.400 ;
        RECT 449.400 506.400 481.050 507.600 ;
        RECT 79.950 504.600 82.050 505.050 ;
        RECT 124.950 504.600 127.050 505.050 ;
        RECT 148.950 504.600 151.050 505.050 ;
        RECT 199.950 504.600 202.050 505.050 ;
        RECT 79.950 503.400 202.050 504.600 ;
        RECT 79.950 502.950 82.050 503.400 ;
        RECT 124.950 502.950 127.050 503.400 ;
        RECT 148.950 502.950 151.050 503.400 ;
        RECT 199.950 502.950 202.050 503.400 ;
        RECT 229.950 504.600 232.050 505.050 ;
        RECT 235.950 504.600 238.050 505.050 ;
        RECT 229.950 503.400 238.050 504.600 ;
        RECT 229.950 502.950 232.050 503.400 ;
        RECT 235.950 502.950 238.050 503.400 ;
        RECT 256.950 504.600 259.050 505.050 ;
        RECT 271.950 504.600 274.050 505.050 ;
        RECT 256.950 503.400 274.050 504.600 ;
        RECT 256.950 502.950 259.050 503.400 ;
        RECT 271.950 502.950 274.050 503.400 ;
        RECT 283.950 504.600 286.050 505.050 ;
        RECT 304.950 504.600 307.050 505.050 ;
        RECT 283.950 503.400 307.050 504.600 ;
        RECT 283.950 502.950 286.050 503.400 ;
        RECT 304.950 502.950 307.050 503.400 ;
        RECT 337.950 504.600 340.050 504.900 ;
        RECT 349.950 504.600 352.050 505.050 ;
        RECT 337.950 503.400 352.050 504.600 ;
        RECT 337.950 502.800 340.050 503.400 ;
        RECT 349.950 502.950 352.050 503.400 ;
        RECT 412.950 504.600 415.050 505.050 ;
        RECT 430.950 504.600 433.050 505.050 ;
        RECT 449.400 504.600 450.600 506.400 ;
        RECT 478.950 505.950 481.050 506.400 ;
        RECT 523.950 507.600 526.050 508.050 ;
        RECT 568.950 507.600 571.050 508.050 ;
        RECT 574.950 507.600 577.050 508.050 ;
        RECT 523.950 506.400 577.050 507.600 ;
        RECT 523.950 505.950 526.050 506.400 ;
        RECT 568.950 505.950 571.050 506.400 ;
        RECT 574.950 505.950 577.050 506.400 ;
        RECT 580.950 507.600 583.050 508.050 ;
        RECT 604.950 507.600 607.050 508.050 ;
        RECT 580.950 506.400 607.050 507.600 ;
        RECT 580.950 505.950 583.050 506.400 ;
        RECT 604.950 505.950 607.050 506.400 ;
        RECT 622.950 507.600 625.050 508.050 ;
        RECT 631.950 507.600 634.050 508.050 ;
        RECT 622.950 506.400 634.050 507.600 ;
        RECT 622.950 505.950 625.050 506.400 ;
        RECT 631.950 505.950 634.050 506.400 ;
        RECT 676.950 507.600 679.050 508.050 ;
        RECT 697.950 507.600 700.050 508.050 ;
        RECT 715.950 507.600 718.050 508.050 ;
        RECT 676.950 506.400 690.600 507.600 ;
        RECT 676.950 505.950 679.050 506.400 ;
        RECT 412.950 503.400 450.600 504.600 ;
        RECT 487.950 504.600 490.050 505.050 ;
        RECT 505.950 504.600 508.050 505.050 ;
        RECT 487.950 503.400 508.050 504.600 ;
        RECT 412.950 502.950 415.050 503.400 ;
        RECT 430.950 502.950 433.050 503.400 ;
        RECT 487.950 502.950 490.050 503.400 ;
        RECT 505.950 502.950 508.050 503.400 ;
        RECT 580.950 504.600 583.050 504.900 ;
        RECT 598.950 504.600 601.050 505.050 ;
        RECT 580.950 503.400 601.050 504.600 ;
        RECT 689.400 504.600 690.600 506.400 ;
        RECT 697.950 506.400 718.050 507.600 ;
        RECT 697.950 505.950 700.050 506.400 ;
        RECT 715.950 505.950 718.050 506.400 ;
        RECT 745.950 507.600 748.050 508.050 ;
        RECT 760.950 507.600 763.050 508.050 ;
        RECT 745.950 506.400 763.050 507.600 ;
        RECT 745.950 505.950 748.050 506.400 ;
        RECT 760.950 505.950 763.050 506.400 ;
        RECT 712.950 504.600 715.050 505.050 ;
        RECT 739.950 504.600 742.050 505.050 ;
        RECT 805.950 504.600 808.050 505.050 ;
        RECT 689.400 503.400 808.050 504.600 ;
        RECT 580.950 502.800 583.050 503.400 ;
        RECT 598.950 502.950 601.050 503.400 ;
        RECT 712.950 502.950 715.050 503.400 ;
        RECT 739.950 502.950 742.050 503.400 ;
        RECT 805.950 502.950 808.050 503.400 ;
        RECT 13.950 501.600 16.050 502.050 ;
        RECT 37.950 501.600 40.050 502.050 ;
        RECT 13.950 500.400 40.050 501.600 ;
        RECT 13.950 499.950 16.050 500.400 ;
        RECT 37.950 499.950 40.050 500.400 ;
        RECT 58.950 501.600 61.050 502.050 ;
        RECT 76.950 501.600 79.050 502.050 ;
        RECT 58.950 500.400 79.050 501.600 ;
        RECT 58.950 499.950 61.050 500.400 ;
        RECT 76.950 499.950 79.050 500.400 ;
        RECT 82.950 501.600 85.050 502.050 ;
        RECT 97.950 501.600 100.050 502.050 ;
        RECT 82.950 500.400 100.050 501.600 ;
        RECT 82.950 499.950 85.050 500.400 ;
        RECT 97.950 499.950 100.050 500.400 ;
        RECT 109.950 501.600 112.050 502.050 ;
        RECT 145.950 501.600 148.050 502.050 ;
        RECT 169.950 501.600 172.050 502.050 ;
        RECT 109.950 500.400 144.600 501.600 ;
        RECT 109.950 499.950 112.050 500.400 ;
        RECT 4.950 498.600 7.050 499.050 ;
        RECT 10.950 498.600 13.050 499.050 ;
        RECT 4.950 497.400 13.050 498.600 ;
        RECT 143.400 498.600 144.600 500.400 ;
        RECT 145.950 500.400 172.050 501.600 ;
        RECT 145.950 499.950 148.050 500.400 ;
        RECT 169.950 499.950 172.050 500.400 ;
        RECT 205.950 501.600 208.050 502.050 ;
        RECT 232.950 501.600 235.050 502.050 ;
        RECT 205.950 500.400 235.050 501.600 ;
        RECT 205.950 499.950 208.050 500.400 ;
        RECT 232.950 499.950 235.050 500.400 ;
        RECT 262.950 501.600 265.050 502.050 ;
        RECT 268.950 501.600 271.050 502.050 ;
        RECT 262.950 500.400 271.050 501.600 ;
        RECT 262.950 499.950 265.050 500.400 ;
        RECT 268.950 499.950 271.050 500.400 ;
        RECT 283.950 501.600 286.050 501.900 ;
        RECT 289.950 501.600 292.050 502.050 ;
        RECT 283.950 500.400 292.050 501.600 ;
        RECT 283.950 499.800 286.050 500.400 ;
        RECT 289.950 499.950 292.050 500.400 ;
        RECT 307.950 501.600 310.050 502.050 ;
        RECT 352.950 501.600 355.050 502.050 ;
        RECT 307.950 500.400 355.050 501.600 ;
        RECT 307.950 499.950 310.050 500.400 ;
        RECT 352.950 499.950 355.050 500.400 ;
        RECT 367.950 501.600 370.050 502.050 ;
        RECT 403.950 501.600 406.050 502.050 ;
        RECT 367.950 500.400 406.050 501.600 ;
        RECT 367.950 499.950 370.050 500.400 ;
        RECT 403.950 499.950 406.050 500.400 ;
        RECT 427.950 501.600 430.050 502.050 ;
        RECT 502.950 501.600 505.050 502.050 ;
        RECT 427.950 500.400 505.050 501.600 ;
        RECT 427.950 499.950 430.050 500.400 ;
        RECT 502.950 499.950 505.050 500.400 ;
        RECT 532.950 501.600 535.050 502.050 ;
        RECT 556.950 501.600 559.050 502.050 ;
        RECT 532.950 500.400 559.050 501.600 ;
        RECT 532.950 499.950 535.050 500.400 ;
        RECT 556.950 499.950 559.050 500.400 ;
        RECT 613.950 501.600 616.050 502.050 ;
        RECT 634.950 501.600 637.050 502.050 ;
        RECT 613.950 500.400 637.050 501.600 ;
        RECT 613.950 499.950 616.050 500.400 ;
        RECT 634.950 499.950 637.050 500.400 ;
        RECT 748.950 501.600 751.050 502.050 ;
        RECT 784.950 501.600 787.050 502.050 ;
        RECT 748.950 500.400 787.050 501.600 ;
        RECT 748.950 499.950 751.050 500.400 ;
        RECT 784.950 499.950 787.050 500.400 ;
        RECT 178.800 498.600 180.900 499.050 ;
        RECT 143.400 497.400 180.900 498.600 ;
        RECT 4.950 496.950 7.050 497.400 ;
        RECT 10.950 496.950 13.050 497.400 ;
        RECT 178.800 496.950 180.900 497.400 ;
        RECT 181.950 496.950 184.050 499.050 ;
        RECT 193.950 498.600 196.050 499.050 ;
        RECT 202.950 498.600 205.050 499.050 ;
        RECT 193.950 497.400 205.050 498.600 ;
        RECT 193.950 496.950 196.050 497.400 ;
        RECT 202.950 496.950 205.050 497.400 ;
        RECT 220.950 498.600 223.050 498.900 ;
        RECT 259.950 498.600 262.050 499.050 ;
        RECT 220.950 497.400 262.050 498.600 ;
        RECT 34.950 495.750 37.050 496.200 ;
        RECT 49.950 495.750 52.050 496.200 ;
        RECT 34.950 494.550 52.050 495.750 ;
        RECT 61.950 495.600 64.050 496.350 ;
        RECT 34.950 494.100 37.050 494.550 ;
        RECT 49.950 494.100 52.050 494.550 ;
        RECT 53.400 494.400 64.050 495.600 ;
        RECT 53.400 492.600 54.600 494.400 ;
        RECT 61.950 494.250 64.050 494.400 ;
        RECT 67.950 495.600 70.050 496.350 ;
        RECT 79.950 495.600 84.000 496.050 ;
        RECT 85.950 495.600 88.050 496.200 ;
        RECT 97.950 495.600 100.050 496.050 ;
        RECT 67.950 494.400 78.600 495.600 ;
        RECT 67.950 494.250 70.050 494.400 ;
        RECT 47.400 491.400 54.600 492.600 ;
        RECT 77.400 492.600 78.600 494.400 ;
        RECT 79.950 493.950 84.600 495.600 ;
        RECT 85.950 494.400 100.050 495.600 ;
        RECT 85.950 494.100 88.050 494.400 ;
        RECT 97.950 493.950 100.050 494.400 ;
        RECT 118.950 493.950 121.050 496.050 ;
        RECT 130.950 495.900 133.050 496.350 ;
        RECT 139.950 495.900 142.050 496.350 ;
        RECT 130.950 494.700 142.050 495.900 ;
        RECT 130.950 494.250 133.050 494.700 ;
        RECT 139.950 494.250 142.050 494.700 ;
        RECT 154.950 495.600 159.000 496.050 ;
        RECT 160.950 495.600 163.050 496.350 ;
        RECT 178.950 495.600 181.050 496.350 ;
        RECT 154.950 493.950 159.600 495.600 ;
        RECT 160.950 494.400 168.600 495.600 ;
        RECT 160.950 494.250 163.050 494.400 ;
        RECT 77.400 492.000 81.450 492.600 ;
        RECT 77.400 491.400 82.050 492.000 ;
        RECT 1.950 489.600 4.050 490.050 ;
        RECT 47.400 489.900 48.600 491.400 ;
        RECT 79.950 490.050 82.050 491.400 ;
        RECT 25.950 489.600 28.050 489.900 ;
        RECT 1.950 488.400 28.050 489.600 ;
        RECT 1.950 487.950 4.050 488.400 ;
        RECT 25.950 487.800 28.050 488.400 ;
        RECT 46.950 487.800 49.050 489.900 ;
        RECT 79.800 489.000 82.050 490.050 ;
        RECT 83.400 489.900 84.600 493.950 ;
        RECT 79.800 487.950 81.900 489.000 ;
        RECT 82.950 487.800 85.050 489.900 ;
        RECT 88.950 489.600 91.050 489.900 ;
        RECT 106.950 489.600 109.050 489.900 ;
        RECT 115.950 489.600 118.050 490.050 ;
        RECT 88.950 488.400 118.050 489.600 ;
        RECT 119.400 489.600 120.600 493.950 ;
        RECT 158.400 490.050 159.600 493.950 ;
        RECT 121.950 489.600 124.050 489.900 ;
        RECT 119.400 488.400 124.050 489.600 ;
        RECT 88.950 487.800 91.050 488.400 ;
        RECT 106.950 487.800 109.050 488.400 ;
        RECT 115.950 487.950 118.050 488.400 ;
        RECT 121.950 487.800 124.050 488.400 ;
        RECT 157.950 487.950 160.050 490.050 ;
        RECT 167.400 487.050 168.600 494.400 ;
        RECT 173.400 494.400 181.050 495.600 ;
        RECT 173.400 490.050 174.600 494.400 ;
        RECT 178.950 494.250 181.050 494.400 ;
        RECT 182.400 490.050 183.600 496.950 ;
        RECT 220.950 496.800 223.050 497.400 ;
        RECT 259.950 496.950 262.050 497.400 ;
        RECT 277.950 498.600 280.050 499.050 ;
        RECT 292.950 498.600 295.050 499.050 ;
        RECT 277.950 497.400 295.050 498.600 ;
        RECT 277.950 496.950 280.050 497.400 ;
        RECT 292.950 496.950 295.050 497.400 ;
        RECT 304.950 498.600 307.050 499.050 ;
        RECT 406.950 498.600 409.050 499.050 ;
        RECT 439.950 498.600 442.050 499.050 ;
        RECT 304.950 497.400 345.600 498.600 ;
        RECT 304.950 496.950 307.050 497.400 ;
        RECT 234.000 495.600 238.050 496.050 ;
        RECT 233.400 493.950 238.050 495.600 ;
        RECT 244.950 495.600 247.050 496.200 ;
        RECT 268.950 495.600 271.050 496.350 ;
        RECT 274.950 495.600 277.050 495.900 ;
        RECT 244.950 494.400 252.450 495.600 ;
        RECT 244.950 494.100 247.050 494.400 ;
        RECT 190.950 492.600 193.050 493.050 ;
        RECT 211.950 492.600 214.050 493.050 ;
        RECT 190.950 491.400 214.050 492.600 ;
        RECT 190.950 490.950 193.050 491.400 ;
        RECT 211.950 490.950 214.050 491.400 ;
        RECT 172.950 487.950 175.050 490.050 ;
        RECT 181.950 487.950 184.050 490.050 ;
        RECT 233.400 489.900 234.600 493.950 ;
        RECT 251.250 490.050 252.450 494.400 ;
        RECT 268.950 494.400 277.050 495.600 ;
        RECT 268.950 494.250 271.050 494.400 ;
        RECT 274.950 493.800 277.050 494.400 ;
        RECT 283.950 495.600 286.050 496.200 ;
        RECT 289.950 495.600 292.050 496.200 ;
        RECT 283.950 494.400 288.600 495.600 ;
        RECT 283.950 494.100 286.050 494.400 ;
        RECT 232.950 487.800 235.050 489.900 ;
        RECT 250.800 487.950 252.900 490.050 ;
        RECT 253.950 489.600 256.050 490.050 ;
        RECT 259.950 489.600 262.050 490.050 ;
        RECT 253.950 488.400 262.050 489.600 ;
        RECT 287.400 489.600 288.600 494.400 ;
        RECT 289.950 494.400 297.600 495.600 ;
        RECT 289.950 494.100 292.050 494.400 ;
        RECT 296.400 492.600 297.600 494.400 ;
        RECT 301.950 494.250 304.050 496.350 ;
        RECT 296.400 492.000 300.600 492.600 ;
        RECT 296.400 491.400 301.050 492.000 ;
        RECT 292.950 489.600 295.050 490.050 ;
        RECT 287.400 488.400 295.050 489.600 ;
        RECT 253.950 487.950 256.050 488.400 ;
        RECT 259.950 487.950 262.050 488.400 ;
        RECT 292.950 487.950 295.050 488.400 ;
        RECT 298.950 487.950 301.050 491.400 ;
        RECT 142.950 486.600 145.050 487.050 ;
        RECT 151.950 486.600 154.050 487.050 ;
        RECT 142.950 485.400 154.050 486.600 ;
        RECT 142.950 484.950 145.050 485.400 ;
        RECT 151.950 484.950 154.050 485.400 ;
        RECT 166.950 484.950 169.050 487.050 ;
        RECT 229.950 486.600 232.050 487.050 ;
        RECT 241.950 486.600 244.050 487.050 ;
        RECT 229.950 485.400 244.050 486.600 ;
        RECT 229.950 484.950 232.050 485.400 ;
        RECT 241.950 484.950 244.050 485.400 ;
        RECT 268.950 486.600 271.050 487.050 ;
        RECT 299.400 486.600 300.600 487.950 ;
        RECT 268.950 485.400 300.600 486.600 ;
        RECT 268.950 484.950 271.050 485.400 ;
        RECT 40.950 483.600 43.050 484.050 ;
        RECT 46.950 483.600 49.050 484.050 ;
        RECT 40.950 482.400 49.050 483.600 ;
        RECT 40.950 481.950 43.050 482.400 ;
        RECT 46.950 481.950 49.050 482.400 ;
        RECT 70.950 483.600 73.050 484.050 ;
        RECT 97.950 483.600 100.050 484.050 ;
        RECT 70.950 482.400 100.050 483.600 ;
        RECT 70.950 481.950 73.050 482.400 ;
        RECT 97.950 481.950 100.050 482.400 ;
        RECT 202.950 480.600 205.050 481.050 ;
        RECT 214.950 480.600 217.050 481.050 ;
        RECT 202.950 479.400 217.050 480.600 ;
        RECT 302.400 480.600 303.600 494.250 ;
        RECT 310.950 493.950 313.050 496.050 ;
        RECT 331.800 495.600 333.900 496.200 ;
        RECT 326.400 494.400 333.900 495.600 ;
        RECT 311.400 490.050 312.600 493.950 ;
        RECT 326.400 492.600 327.600 494.400 ;
        RECT 331.800 494.100 333.900 494.400 ;
        RECT 323.400 491.400 327.600 492.600 ;
        RECT 323.400 490.050 324.600 491.400 ;
        RECT 344.400 490.050 345.600 497.400 ;
        RECT 406.950 497.400 442.050 498.600 ;
        RECT 406.950 496.950 409.050 497.400 ;
        RECT 364.950 495.600 367.050 496.350 ;
        RECT 382.950 495.600 385.050 496.350 ;
        RECT 409.950 495.600 412.050 496.050 ;
        RECT 364.950 494.400 381.600 495.600 ;
        RECT 364.950 494.250 367.050 494.400 ;
        RECT 380.400 492.600 381.600 494.400 ;
        RECT 382.950 494.400 412.050 495.600 ;
        RECT 382.950 494.250 385.050 494.400 ;
        RECT 350.400 492.000 381.600 492.600 ;
        RECT 349.950 491.400 381.600 492.000 ;
        RECT 307.950 488.400 312.600 490.050 ;
        RECT 319.950 488.400 324.600 490.050 ;
        RECT 307.950 487.950 312.000 488.400 ;
        RECT 319.950 487.950 324.000 488.400 ;
        RECT 343.950 487.950 346.050 490.050 ;
        RECT 349.950 487.950 352.050 491.400 ;
        RECT 380.400 490.050 381.600 491.400 ;
        RECT 389.400 490.050 390.600 494.400 ;
        RECT 409.950 493.950 412.050 494.400 ;
        RECT 421.950 495.600 424.050 496.200 ;
        RECT 421.950 494.400 426.600 495.600 ;
        RECT 421.950 494.100 424.050 494.400 ;
        RECT 355.950 489.600 358.050 490.050 ;
        RECT 370.950 489.600 373.050 490.050 ;
        RECT 355.950 488.400 373.050 489.600 ;
        RECT 355.950 487.950 358.050 488.400 ;
        RECT 370.950 487.950 373.050 488.400 ;
        RECT 379.950 487.950 382.050 490.050 ;
        RECT 388.950 487.950 391.050 490.050 ;
        RECT 394.950 489.600 397.050 490.050 ;
        RECT 400.950 489.600 403.050 490.050 ;
        RECT 394.950 488.400 403.050 489.600 ;
        RECT 394.950 487.950 397.050 488.400 ;
        RECT 400.950 487.950 403.050 488.400 ;
        RECT 371.400 486.600 372.600 487.950 ;
        RECT 425.400 487.050 426.600 494.400 ;
        RECT 428.400 490.050 429.600 497.400 ;
        RECT 439.950 496.950 442.050 497.400 ;
        RECT 520.950 498.600 523.050 499.050 ;
        RECT 547.950 498.600 550.050 499.050 ;
        RECT 520.950 497.400 550.050 498.600 ;
        RECT 520.950 496.950 523.050 497.400 ;
        RECT 547.950 496.950 550.050 497.400 ;
        RECT 595.950 498.600 600.000 499.050 ;
        RECT 601.950 498.600 604.050 499.050 ;
        RECT 607.950 498.600 610.050 499.200 ;
        RECT 595.950 496.950 600.600 498.600 ;
        RECT 601.950 497.400 610.050 498.600 ;
        RECT 601.950 496.950 604.050 497.400 ;
        RECT 607.950 497.100 610.050 497.400 ;
        RECT 709.950 498.600 712.050 499.050 ;
        RECT 718.950 498.600 721.050 499.050 ;
        RECT 709.950 497.400 721.050 498.600 ;
        RECT 709.950 496.950 712.050 497.400 ;
        RECT 718.950 496.950 721.050 497.400 ;
        RECT 829.950 498.600 832.050 499.050 ;
        RECT 841.950 498.600 844.050 499.050 ;
        RECT 829.950 497.400 844.050 498.600 ;
        RECT 829.950 496.950 832.050 497.400 ;
        RECT 841.950 496.950 844.050 497.400 ;
        RECT 445.950 495.600 448.050 496.350 ;
        RECT 466.950 495.600 469.050 496.050 ;
        RECT 445.950 494.400 469.050 495.600 ;
        RECT 445.950 494.250 448.050 494.400 ;
        RECT 466.950 493.950 469.050 494.400 ;
        RECT 496.950 495.600 499.050 496.350 ;
        RECT 496.950 494.400 516.600 495.600 ;
        RECT 496.950 494.250 499.050 494.400 ;
        RECT 427.950 487.950 430.050 490.050 ;
        RECT 515.400 489.900 516.600 494.400 ;
        RECT 544.950 492.600 547.050 496.050 ;
        RECT 550.950 495.750 553.050 496.200 ;
        RECT 559.800 495.750 561.900 496.200 ;
        RECT 550.950 494.550 561.900 495.750 ;
        RECT 550.950 494.100 553.050 494.550 ;
        RECT 559.800 494.100 561.900 494.550 ;
        RECT 562.950 493.950 565.050 496.050 ;
        RECT 574.800 494.100 576.900 496.200 ;
        RECT 577.950 495.750 580.050 496.200 ;
        RECT 589.950 495.750 592.050 496.200 ;
        RECT 577.950 494.550 592.050 495.750 ;
        RECT 577.950 494.100 580.050 494.550 ;
        RECT 589.950 494.100 592.050 494.550 ;
        RECT 599.400 495.600 600.600 496.950 ;
        RECT 607.950 495.600 610.050 496.050 ;
        RECT 631.950 495.600 634.050 496.050 ;
        RECT 599.400 494.400 610.050 495.600 ;
        RECT 533.400 492.000 547.050 492.600 ;
        RECT 533.400 491.400 546.600 492.000 ;
        RECT 533.400 490.050 534.600 491.400 ;
        RECT 514.950 487.800 517.050 489.900 ;
        RECT 529.950 488.400 534.600 490.050 ;
        RECT 535.950 489.450 538.050 489.900 ;
        RECT 547.950 489.450 550.050 489.900 ;
        RECT 529.950 487.950 534.000 488.400 ;
        RECT 535.950 488.250 550.050 489.450 ;
        RECT 563.400 489.600 564.600 493.950 ;
        RECT 575.400 492.600 576.600 494.100 ;
        RECT 607.950 493.950 610.050 494.400 ;
        RECT 626.400 494.400 634.050 495.600 ;
        RECT 626.400 492.600 627.600 494.400 ;
        RECT 631.950 493.950 634.050 494.400 ;
        RECT 643.950 495.600 646.050 496.050 ;
        RECT 655.950 495.600 658.050 496.350 ;
        RECT 643.950 494.400 658.050 495.600 ;
        RECT 643.950 493.950 646.050 494.400 ;
        RECT 655.950 494.250 658.050 494.400 ;
        RECT 691.950 495.750 694.050 496.200 ;
        RECT 703.950 495.750 706.050 496.200 ;
        RECT 691.950 494.550 706.050 495.750 ;
        RECT 691.950 494.100 694.050 494.550 ;
        RECT 703.950 494.100 706.050 494.550 ;
        RECT 712.950 495.600 717.000 496.050 ;
        RECT 712.950 493.950 717.600 495.600 ;
        RECT 721.950 494.100 724.050 496.200 ;
        RECT 733.950 495.600 736.050 496.200 ;
        RECT 725.400 494.400 736.050 495.600 ;
        RECT 685.950 492.600 688.050 493.050 ;
        RECT 575.400 491.400 627.600 492.600 ;
        RECT 659.400 492.000 688.050 492.600 ;
        RECT 658.950 491.400 688.050 492.000 ;
        RECT 716.400 492.600 717.600 493.950 ;
        RECT 722.400 492.600 723.600 494.100 ;
        RECT 716.400 491.400 723.600 492.600 ;
        RECT 583.950 489.600 586.050 490.050 ;
        RECT 611.400 489.900 612.600 491.400 ;
        RECT 563.400 488.400 586.050 489.600 ;
        RECT 535.950 487.800 538.050 488.250 ;
        RECT 547.950 487.800 550.050 488.250 ;
        RECT 583.950 487.950 586.050 488.400 ;
        RECT 610.950 487.800 613.050 489.900 ;
        RECT 637.950 489.600 640.050 490.050 ;
        RECT 652.950 489.600 655.050 490.050 ;
        RECT 637.950 488.400 655.050 489.600 ;
        RECT 637.950 487.950 640.050 488.400 ;
        RECT 652.950 487.950 655.050 488.400 ;
        RECT 658.950 487.950 661.050 491.400 ;
        RECT 685.950 490.950 688.050 491.400 ;
        RECT 725.400 490.050 726.600 494.400 ;
        RECT 733.950 494.100 736.050 494.400 ;
        RECT 742.950 493.950 745.050 496.050 ;
        RECT 772.950 495.600 775.050 496.050 ;
        RECT 784.950 495.600 787.050 496.200 ;
        RECT 799.950 495.600 802.050 496.350 ;
        RECT 772.950 494.400 802.050 495.600 ;
        RECT 772.950 493.950 775.050 494.400 ;
        RECT 784.950 494.100 787.050 494.400 ;
        RECT 799.950 494.250 802.050 494.400 ;
        RECT 823.950 495.600 826.050 496.350 ;
        RECT 853.950 495.600 856.050 496.050 ;
        RECT 823.950 494.400 856.050 495.600 ;
        RECT 823.950 494.250 826.050 494.400 ;
        RECT 853.950 493.950 856.050 494.400 ;
        RECT 743.400 490.050 744.600 493.950 ;
        RECT 724.950 487.950 727.050 490.050 ;
        RECT 742.950 487.950 745.050 490.050 ;
        RECT 802.950 489.600 805.050 490.050 ;
        RECT 808.950 489.600 811.050 490.050 ;
        RECT 802.950 488.400 811.050 489.600 ;
        RECT 802.950 487.950 805.050 488.400 ;
        RECT 808.950 487.950 811.050 488.400 ;
        RECT 385.950 486.600 388.050 487.050 ;
        RECT 406.950 486.600 409.050 487.050 ;
        RECT 371.400 485.400 409.050 486.600 ;
        RECT 425.400 486.900 429.000 487.050 ;
        RECT 425.400 485.400 430.050 486.900 ;
        RECT 385.950 484.950 388.050 485.400 ;
        RECT 406.950 484.950 409.050 485.400 ;
        RECT 426.000 484.950 430.050 485.400 ;
        RECT 442.950 486.600 445.050 487.050 ;
        RECT 517.950 486.600 520.050 487.050 ;
        RECT 442.950 485.400 520.050 486.600 ;
        RECT 442.950 484.950 445.050 485.400 ;
        RECT 517.950 484.950 520.050 485.400 ;
        RECT 541.950 486.600 544.050 487.050 ;
        RECT 550.950 486.600 553.050 487.050 ;
        RECT 571.950 486.600 574.050 487.050 ;
        RECT 541.950 485.400 574.050 486.600 ;
        RECT 541.950 484.950 544.050 485.400 ;
        RECT 550.950 484.950 553.050 485.400 ;
        RECT 571.950 484.950 574.050 485.400 ;
        RECT 691.950 486.600 694.050 487.050 ;
        RECT 736.950 486.600 739.050 487.050 ;
        RECT 691.950 485.400 739.050 486.600 ;
        RECT 691.950 484.950 694.050 485.400 ;
        RECT 736.950 484.950 739.050 485.400 ;
        RECT 820.950 486.600 823.050 487.050 ;
        RECT 838.950 486.600 841.050 487.050 ;
        RECT 820.950 485.400 841.050 486.600 ;
        RECT 820.950 484.950 823.050 485.400 ;
        RECT 838.950 484.950 841.050 485.400 ;
        RECT 427.950 484.800 430.050 484.950 ;
        RECT 319.950 483.600 322.050 484.050 ;
        RECT 331.950 483.600 334.050 484.050 ;
        RECT 319.950 482.400 334.050 483.600 ;
        RECT 319.950 481.950 322.050 482.400 ;
        RECT 331.950 481.950 334.050 482.400 ;
        RECT 340.950 483.600 343.050 484.050 ;
        RECT 361.950 483.600 364.050 484.050 ;
        RECT 340.950 482.400 364.050 483.600 ;
        RECT 340.950 481.950 343.050 482.400 ;
        RECT 361.950 481.950 364.050 482.400 ;
        RECT 472.950 483.600 475.050 484.050 ;
        RECT 508.950 483.600 511.050 484.050 ;
        RECT 472.950 482.400 511.050 483.600 ;
        RECT 472.950 481.950 475.050 482.400 ;
        RECT 508.950 481.950 511.050 482.400 ;
        RECT 583.950 483.600 586.050 484.050 ;
        RECT 622.950 483.600 625.050 484.050 ;
        RECT 583.950 482.400 625.050 483.600 ;
        RECT 583.950 481.950 586.050 482.400 ;
        RECT 622.950 481.950 625.050 482.400 ;
        RECT 634.950 483.600 637.050 484.050 ;
        RECT 742.950 483.600 745.050 484.050 ;
        RECT 634.950 482.400 745.050 483.600 ;
        RECT 634.950 481.950 637.050 482.400 ;
        RECT 742.950 481.950 745.050 482.400 ;
        RECT 322.950 480.600 325.050 481.050 ;
        RECT 337.950 480.600 340.050 481.050 ;
        RECT 302.400 479.400 312.600 480.600 ;
        RECT 202.950 478.950 205.050 479.400 ;
        RECT 214.950 478.950 217.050 479.400 ;
        RECT 76.950 477.600 79.050 478.050 ;
        RECT 130.950 477.600 133.050 478.050 ;
        RECT 76.950 476.400 133.050 477.600 ;
        RECT 76.950 475.950 79.050 476.400 ;
        RECT 130.950 475.950 133.050 476.400 ;
        RECT 247.950 477.600 250.050 478.050 ;
        RECT 274.950 477.600 277.050 478.050 ;
        RECT 247.950 476.400 277.050 477.600 ;
        RECT 247.950 475.950 250.050 476.400 ;
        RECT 274.950 475.950 277.050 476.400 ;
        RECT 298.950 477.600 301.050 478.050 ;
        RECT 307.950 477.600 310.050 478.050 ;
        RECT 298.950 476.400 310.050 477.600 ;
        RECT 311.400 477.600 312.600 479.400 ;
        RECT 322.950 479.400 340.050 480.600 ;
        RECT 322.950 478.950 325.050 479.400 ;
        RECT 337.950 478.950 340.050 479.400 ;
        RECT 385.950 480.600 388.050 481.050 ;
        RECT 418.950 480.600 421.050 481.050 ;
        RECT 385.950 479.400 421.050 480.600 ;
        RECT 385.950 478.950 388.050 479.400 ;
        RECT 418.950 478.950 421.050 479.400 ;
        RECT 517.950 480.600 520.050 481.050 ;
        RECT 577.950 480.600 580.050 481.050 ;
        RECT 517.950 479.400 580.050 480.600 ;
        RECT 517.950 478.950 520.050 479.400 ;
        RECT 577.950 478.950 580.050 479.400 ;
        RECT 601.950 480.600 604.050 481.050 ;
        RECT 616.950 480.600 619.050 481.050 ;
        RECT 601.950 479.400 619.050 480.600 ;
        RECT 601.950 478.950 604.050 479.400 ;
        RECT 616.950 478.950 619.050 479.400 ;
        RECT 631.950 480.600 634.050 481.050 ;
        RECT 778.950 480.600 781.050 481.050 ;
        RECT 631.950 479.400 781.050 480.600 ;
        RECT 631.950 478.950 634.050 479.400 ;
        RECT 778.950 478.950 781.050 479.400 ;
        RECT 799.950 480.600 802.050 481.050 ;
        RECT 829.950 480.600 832.050 481.050 ;
        RECT 799.950 479.400 832.050 480.600 ;
        RECT 799.950 478.950 802.050 479.400 ;
        RECT 829.950 478.950 832.050 479.400 ;
        RECT 337.950 477.600 340.050 477.900 ;
        RECT 311.400 476.400 340.050 477.600 ;
        RECT 298.950 475.950 301.050 476.400 ;
        RECT 307.950 475.950 310.050 476.400 ;
        RECT 337.950 475.800 340.050 476.400 ;
        RECT 487.950 477.600 490.050 478.050 ;
        RECT 514.950 477.600 517.050 478.050 ;
        RECT 580.950 477.600 583.050 478.050 ;
        RECT 487.950 476.400 583.050 477.600 ;
        RECT 487.950 475.950 490.050 476.400 ;
        RECT 514.950 475.950 517.050 476.400 ;
        RECT 580.950 475.950 583.050 476.400 ;
        RECT 586.950 477.600 589.050 478.050 ;
        RECT 643.950 477.600 646.050 478.050 ;
        RECT 586.950 476.400 646.050 477.600 ;
        RECT 586.950 475.950 589.050 476.400 ;
        RECT 643.950 475.950 646.050 476.400 ;
        RECT 673.950 477.600 676.050 478.050 ;
        RECT 790.950 477.600 793.050 478.050 ;
        RECT 796.950 477.600 799.050 478.050 ;
        RECT 673.950 477.000 762.600 477.600 ;
        RECT 673.950 476.400 763.050 477.000 ;
        RECT 673.950 475.950 676.050 476.400 ;
        RECT 34.950 474.600 37.050 475.050 ;
        RECT 40.950 474.600 43.050 475.050 ;
        RECT 313.800 474.600 315.900 475.050 ;
        RECT 34.950 473.400 315.900 474.600 ;
        RECT 34.950 472.950 37.050 473.400 ;
        RECT 40.950 472.950 43.050 473.400 ;
        RECT 313.800 472.950 315.900 473.400 ;
        RECT 316.950 474.600 319.050 475.050 ;
        RECT 340.950 474.600 343.050 475.050 ;
        RECT 316.950 473.400 343.050 474.600 ;
        RECT 316.950 472.950 319.050 473.400 ;
        RECT 340.950 472.950 343.050 473.400 ;
        RECT 358.950 474.600 361.050 475.050 ;
        RECT 436.950 474.600 439.050 475.050 ;
        RECT 358.950 473.400 439.050 474.600 ;
        RECT 358.950 472.950 361.050 473.400 ;
        RECT 436.950 472.950 439.050 473.400 ;
        RECT 457.950 474.600 460.050 475.050 ;
        RECT 502.950 474.600 505.050 475.050 ;
        RECT 520.950 474.600 523.050 475.050 ;
        RECT 529.950 474.600 532.050 475.050 ;
        RECT 457.950 473.400 532.050 474.600 ;
        RECT 457.950 472.950 460.050 473.400 ;
        RECT 502.950 472.950 505.050 473.400 ;
        RECT 520.950 472.950 523.050 473.400 ;
        RECT 529.950 472.950 532.050 473.400 ;
        RECT 544.950 474.600 547.050 475.050 ;
        RECT 587.400 474.600 588.600 475.950 ;
        RECT 544.950 473.400 588.600 474.600 ;
        RECT 544.950 472.950 547.050 473.400 ;
        RECT 760.950 472.950 763.050 476.400 ;
        RECT 790.950 476.400 799.050 477.600 ;
        RECT 790.950 475.950 793.050 476.400 ;
        RECT 796.950 475.950 799.050 476.400 ;
        RECT 97.950 471.600 100.050 472.050 ;
        RECT 109.950 471.600 112.050 472.050 ;
        RECT 97.950 470.400 112.050 471.600 ;
        RECT 97.950 469.950 100.050 470.400 ;
        RECT 109.950 469.950 112.050 470.400 ;
        RECT 151.950 471.600 154.050 472.050 ;
        RECT 268.950 471.600 271.050 472.050 ;
        RECT 151.950 470.400 271.050 471.600 ;
        RECT 151.950 469.950 154.050 470.400 ;
        RECT 268.950 469.950 271.050 470.400 ;
        RECT 274.950 471.600 277.050 472.050 ;
        RECT 341.400 471.600 342.600 472.950 ;
        RECT 394.950 471.600 397.050 472.050 ;
        RECT 412.950 471.600 415.050 472.050 ;
        RECT 274.950 470.400 324.600 471.600 ;
        RECT 341.400 470.400 415.050 471.600 ;
        RECT 274.950 469.950 277.050 470.400 ;
        RECT 283.950 468.600 286.050 469.050 ;
        RECT 323.400 468.600 324.600 470.400 ;
        RECT 394.950 469.950 397.050 470.400 ;
        RECT 412.950 469.950 415.050 470.400 ;
        RECT 427.950 471.600 430.050 472.050 ;
        RECT 748.950 471.600 751.050 472.050 ;
        RECT 790.950 471.600 793.050 472.050 ;
        RECT 814.950 471.600 817.050 472.050 ;
        RECT 427.950 470.400 817.050 471.600 ;
        RECT 427.950 469.950 430.050 470.400 ;
        RECT 748.950 469.950 751.050 470.400 ;
        RECT 790.950 469.950 793.050 470.400 ;
        RECT 814.950 469.950 817.050 470.400 ;
        RECT 385.950 468.600 388.050 469.050 ;
        RECT 283.950 467.400 300.600 468.600 ;
        RECT 323.400 467.400 388.050 468.600 ;
        RECT 283.950 466.950 286.050 467.400 ;
        RECT 61.950 465.600 64.050 466.050 ;
        RECT 64.950 465.600 67.050 466.050 ;
        RECT 100.950 465.600 103.050 466.050 ;
        RECT 61.950 464.400 103.050 465.600 ;
        RECT 61.950 463.950 64.050 464.400 ;
        RECT 64.950 463.950 67.050 464.400 ;
        RECT 100.950 463.950 103.050 464.400 ;
        RECT 109.950 465.600 112.050 466.050 ;
        RECT 205.950 465.600 208.050 466.050 ;
        RECT 109.950 464.400 208.050 465.600 ;
        RECT 299.400 465.600 300.600 467.400 ;
        RECT 385.950 466.950 388.050 467.400 ;
        RECT 466.950 468.600 469.050 469.050 ;
        RECT 631.950 468.600 634.050 469.050 ;
        RECT 466.950 467.400 634.050 468.600 ;
        RECT 466.950 466.950 469.050 467.400 ;
        RECT 631.950 466.950 634.050 467.400 ;
        RECT 643.950 468.600 646.050 469.050 ;
        RECT 688.950 468.600 691.050 469.050 ;
        RECT 643.950 467.400 691.050 468.600 ;
        RECT 643.950 466.950 646.050 467.400 ;
        RECT 688.950 466.950 691.050 467.400 ;
        RECT 718.950 468.600 721.050 469.050 ;
        RECT 739.950 468.600 742.050 469.050 ;
        RECT 718.950 467.400 742.050 468.600 ;
        RECT 718.950 466.950 721.050 467.400 ;
        RECT 739.950 466.950 742.050 467.400 ;
        RECT 388.950 465.600 391.050 466.050 ;
        RECT 299.400 464.400 391.050 465.600 ;
        RECT 109.950 463.950 112.050 464.400 ;
        RECT 205.950 463.950 208.050 464.400 ;
        RECT 388.950 463.950 391.050 464.400 ;
        RECT 406.950 465.600 409.050 466.050 ;
        RECT 430.950 465.600 433.050 466.050 ;
        RECT 406.950 464.400 433.050 465.600 ;
        RECT 406.950 463.950 409.050 464.400 ;
        RECT 430.950 463.950 433.050 464.400 ;
        RECT 571.950 465.600 574.050 466.050 ;
        RECT 628.950 465.600 631.050 466.050 ;
        RECT 571.950 464.400 631.050 465.600 ;
        RECT 571.950 463.950 574.050 464.400 ;
        RECT 628.950 463.950 631.050 464.400 ;
        RECT 679.950 465.600 682.050 466.050 ;
        RECT 700.950 465.600 703.050 466.050 ;
        RECT 679.950 464.400 703.050 465.600 ;
        RECT 679.950 463.950 682.050 464.400 ;
        RECT 700.950 463.950 703.050 464.400 ;
        RECT 502.950 462.600 505.050 463.050 ;
        RECT 532.950 462.600 535.050 463.050 ;
        RECT 553.950 462.600 556.050 463.050 ;
        RECT 502.950 461.400 556.050 462.600 ;
        RECT 502.950 460.950 505.050 461.400 ;
        RECT 532.950 460.950 535.050 461.400 ;
        RECT 553.950 460.950 556.050 461.400 ;
        RECT 586.950 462.600 589.050 463.050 ;
        RECT 634.950 462.600 637.050 463.050 ;
        RECT 586.950 461.400 637.050 462.600 ;
        RECT 586.950 460.950 589.050 461.400 ;
        RECT 634.950 460.950 637.050 461.400 ;
        RECT 670.950 462.600 673.050 463.050 ;
        RECT 745.950 462.600 748.050 463.050 ;
        RECT 670.950 461.400 748.050 462.600 ;
        RECT 670.950 460.950 673.050 461.400 ;
        RECT 745.950 460.950 748.050 461.400 ;
        RECT 766.950 462.600 769.050 463.050 ;
        RECT 823.950 462.600 826.050 463.050 ;
        RECT 766.950 461.400 826.050 462.600 ;
        RECT 766.950 460.950 769.050 461.400 ;
        RECT 823.950 460.950 826.050 461.400 ;
        RECT 64.950 459.600 67.050 460.050 ;
        RECT 79.950 459.600 82.050 460.050 ;
        RECT 64.950 458.400 82.050 459.600 ;
        RECT 64.950 457.950 67.050 458.400 ;
        RECT 79.950 457.950 82.050 458.400 ;
        RECT 94.950 459.600 97.050 460.050 ;
        RECT 106.950 459.600 109.050 460.050 ;
        RECT 94.950 458.400 109.050 459.600 ;
        RECT 94.950 457.950 97.050 458.400 ;
        RECT 106.950 457.950 109.050 458.400 ;
        RECT 190.950 459.600 193.050 460.050 ;
        RECT 205.950 459.600 208.050 460.050 ;
        RECT 220.950 459.600 223.050 460.050 ;
        RECT 190.950 458.400 223.050 459.600 ;
        RECT 190.950 457.950 193.050 458.400 ;
        RECT 205.950 457.950 208.050 458.400 ;
        RECT 220.950 457.950 223.050 458.400 ;
        RECT 298.950 459.600 301.050 460.050 ;
        RECT 307.800 459.600 309.900 460.050 ;
        RECT 298.950 458.400 309.900 459.600 ;
        RECT 298.950 457.950 301.050 458.400 ;
        RECT 307.800 457.950 309.900 458.400 ;
        RECT 550.950 459.600 553.050 460.050 ;
        RECT 583.950 459.600 586.050 460.050 ;
        RECT 643.950 459.600 646.050 460.050 ;
        RECT 550.950 458.400 570.600 459.600 ;
        RECT 550.950 457.950 553.050 458.400 ;
        RECT 10.950 456.600 13.050 457.050 ;
        RECT 16.950 456.600 19.050 457.050 ;
        RECT 10.950 455.400 19.050 456.600 ;
        RECT 10.950 454.950 13.050 455.400 ;
        RECT 16.950 454.950 19.050 455.400 ;
        RECT 445.950 456.600 448.050 457.050 ;
        RECT 475.950 456.600 478.050 457.050 ;
        RECT 445.950 455.400 478.050 456.600 ;
        RECT 569.400 456.600 570.600 458.400 ;
        RECT 583.950 458.400 646.050 459.600 ;
        RECT 583.950 457.950 586.050 458.400 ;
        RECT 643.950 457.950 646.050 458.400 ;
        RECT 826.950 459.600 829.050 460.050 ;
        RECT 832.950 459.600 835.050 460.050 ;
        RECT 826.950 458.400 835.050 459.600 ;
        RECT 826.950 457.950 829.050 458.400 ;
        RECT 832.950 457.950 835.050 458.400 ;
        RECT 604.950 456.600 607.050 457.050 ;
        RECT 569.400 455.400 607.050 456.600 ;
        RECT 445.950 454.950 448.050 455.400 ;
        RECT 475.950 454.950 478.050 455.400 ;
        RECT 590.400 454.050 591.600 455.400 ;
        RECT 604.950 454.950 607.050 455.400 ;
        RECT 658.950 456.600 661.050 457.050 ;
        RECT 694.950 456.600 697.050 457.050 ;
        RECT 658.950 455.400 697.050 456.600 ;
        RECT 658.950 454.950 661.050 455.400 ;
        RECT 694.950 454.950 697.050 455.400 ;
        RECT 25.950 453.600 28.050 454.050 ;
        RECT 34.950 453.600 37.050 454.050 ;
        RECT 25.950 452.400 37.050 453.600 ;
        RECT 25.950 451.950 28.050 452.400 ;
        RECT 34.950 451.950 37.050 452.400 ;
        RECT 55.950 453.600 58.050 453.900 ;
        RECT 70.950 453.600 73.050 454.050 ;
        RECT 55.950 452.400 73.050 453.600 ;
        RECT 55.950 451.800 58.050 452.400 ;
        RECT 70.950 451.950 73.050 452.400 ;
        RECT 76.950 453.600 79.050 454.050 ;
        RECT 130.950 453.600 133.050 454.050 ;
        RECT 142.950 453.600 145.050 454.050 ;
        RECT 76.950 452.400 84.600 453.600 ;
        RECT 76.950 451.950 79.050 452.400 ;
        RECT 10.950 449.100 13.050 451.200 ;
        RECT 11.400 445.050 12.600 449.100 ;
        RECT 22.950 448.950 25.050 451.050 ;
        RECT 63.000 450.600 67.050 451.050 ;
        RECT 62.400 448.950 67.050 450.600 ;
        RECT 23.400 445.050 24.600 448.950 ;
        RECT 7.950 443.400 12.600 445.050 ;
        RECT 7.950 442.950 12.000 443.400 ;
        RECT 22.950 442.950 25.050 445.050 ;
        RECT 58.950 444.600 61.050 444.750 ;
        RECT 62.400 444.600 63.600 448.950 ;
        RECT 58.950 443.400 63.600 444.600 ;
        RECT 67.950 444.300 70.050 444.750 ;
        RECT 79.950 444.300 82.050 444.750 ;
        RECT 58.950 442.650 61.050 443.400 ;
        RECT 67.950 443.100 82.050 444.300 ;
        RECT 67.950 442.650 70.050 443.100 ;
        RECT 79.950 442.650 82.050 443.100 ;
        RECT 83.400 442.050 84.600 452.400 ;
        RECT 130.950 452.400 145.050 453.600 ;
        RECT 130.950 451.950 133.050 452.400 ;
        RECT 142.950 451.950 145.050 452.400 ;
        RECT 85.950 448.950 88.050 451.050 ;
        RECT 94.950 449.100 97.050 451.200 ;
        RECT 100.950 450.750 103.050 451.200 ;
        RECT 109.950 450.750 112.050 451.200 ;
        RECT 100.950 449.550 112.050 450.750 ;
        RECT 100.950 449.100 103.050 449.550 ;
        RECT 109.950 449.100 112.050 449.550 ;
        RECT 115.950 449.100 118.050 451.200 ;
        RECT 121.950 450.750 124.050 451.200 ;
        RECT 130.950 450.750 133.050 450.900 ;
        RECT 121.950 449.550 133.050 450.750 ;
        RECT 175.950 450.600 178.050 454.050 ;
        RECT 187.950 453.600 190.050 454.050 ;
        RECT 211.950 453.600 214.050 454.050 ;
        RECT 187.950 452.400 214.050 453.600 ;
        RECT 187.950 451.950 190.050 452.400 ;
        RECT 211.950 451.950 214.050 452.400 ;
        RECT 319.950 453.600 322.050 454.050 ;
        RECT 355.950 453.600 358.050 454.050 ;
        RECT 370.950 453.600 373.050 454.050 ;
        RECT 319.950 452.400 327.600 453.600 ;
        RECT 319.950 451.950 322.050 452.400 ;
        RECT 196.950 450.600 199.050 451.050 ;
        RECT 208.950 450.600 211.050 451.050 ;
        RECT 175.950 450.000 211.050 450.600 ;
        RECT 121.950 449.100 124.050 449.550 ;
        RECT 86.400 445.050 87.600 448.950 ;
        RECT 95.400 447.600 96.600 449.100 ;
        RECT 116.400 447.600 117.600 449.100 ;
        RECT 130.950 448.800 133.050 449.550 ;
        RECT 176.400 449.400 211.050 450.000 ;
        RECT 196.950 448.950 199.050 449.400 ;
        RECT 95.400 447.000 105.600 447.600 ;
        RECT 95.400 446.400 106.050 447.000 ;
        RECT 116.400 446.400 126.600 447.600 ;
        RECT 85.950 442.950 88.050 445.050 ;
        RECT 103.950 442.950 106.050 446.400 ;
        RECT 109.950 444.600 112.050 445.050 ;
        RECT 118.950 444.600 121.050 444.900 ;
        RECT 109.950 443.400 121.050 444.600 ;
        RECT 125.400 444.600 126.600 446.400 ;
        RECT 133.950 444.600 136.050 445.050 ;
        RECT 125.400 443.400 136.050 444.600 ;
        RECT 109.950 442.950 112.050 443.400 ;
        RECT 118.950 442.800 121.050 443.400 ;
        RECT 133.950 442.950 136.050 443.400 ;
        RECT 139.950 444.600 142.050 444.750 ;
        RECT 151.950 444.600 154.050 448.050 ;
        RECT 139.950 444.000 154.050 444.600 ;
        RECT 175.950 444.300 178.050 444.750 ;
        RECT 202.950 444.300 205.050 444.750 ;
        RECT 139.950 443.400 153.600 444.000 ;
        RECT 139.950 442.650 142.050 443.400 ;
        RECT 175.950 443.100 205.050 444.300 ;
        RECT 175.950 442.650 178.050 443.100 ;
        RECT 202.950 442.650 205.050 443.100 ;
        RECT 206.400 442.050 207.600 449.400 ;
        RECT 208.950 448.950 211.050 449.400 ;
        RECT 214.950 450.600 217.050 451.050 ;
        RECT 247.950 450.600 250.050 451.050 ;
        RECT 283.950 450.600 286.050 451.050 ;
        RECT 214.950 449.400 250.050 450.600 ;
        RECT 275.400 450.000 286.050 450.600 ;
        RECT 214.950 448.950 217.050 449.400 ;
        RECT 247.950 448.950 250.050 449.400 ;
        RECT 274.950 449.400 286.050 450.000 ;
        RECT 274.950 445.800 277.050 449.400 ;
        RECT 283.950 448.950 286.050 449.400 ;
        RECT 292.950 448.950 295.050 451.050 ;
        RECT 304.800 449.100 307.050 451.200 ;
        RECT 307.950 450.600 310.050 451.050 ;
        RECT 322.950 450.600 325.050 451.200 ;
        RECT 307.950 449.400 325.050 450.600 ;
        RECT 211.950 444.600 214.050 445.050 ;
        RECT 277.950 444.600 280.050 445.050 ;
        RECT 283.950 444.600 286.050 445.050 ;
        RECT 211.950 443.400 286.050 444.600 ;
        RECT 293.400 444.600 294.600 448.950 ;
        RECT 305.400 447.600 306.600 449.100 ;
        RECT 307.950 448.950 310.050 449.400 ;
        RECT 322.950 449.100 325.050 449.400 ;
        RECT 305.400 446.400 315.600 447.600 ;
        RECT 314.400 444.600 315.600 446.400 ;
        RECT 319.950 444.600 322.050 444.900 ;
        RECT 293.400 443.400 303.600 444.600 ;
        RECT 314.400 443.400 322.050 444.600 ;
        RECT 211.950 442.950 214.050 443.400 ;
        RECT 277.950 442.950 280.050 443.400 ;
        RECT 283.950 442.950 286.050 443.400 ;
        RECT 4.950 441.600 7.050 442.050 ;
        RECT 19.950 441.600 22.050 442.050 ;
        RECT 4.950 440.400 22.050 441.600 ;
        RECT 4.950 439.950 7.050 440.400 ;
        RECT 19.950 439.950 22.050 440.400 ;
        RECT 82.950 439.950 85.050 442.050 ;
        RECT 91.950 441.600 94.050 442.050 ;
        RECT 106.950 441.600 109.050 442.050 ;
        RECT 91.950 440.400 109.050 441.600 ;
        RECT 91.950 439.950 94.050 440.400 ;
        RECT 106.950 439.950 109.050 440.400 ;
        RECT 130.950 441.600 133.050 442.050 ;
        RECT 136.950 441.600 139.050 442.050 ;
        RECT 130.950 440.400 139.050 441.600 ;
        RECT 130.950 439.950 133.050 440.400 ;
        RECT 136.950 439.950 139.050 440.400 ;
        RECT 205.950 439.950 208.050 442.050 ;
        RECT 302.400 441.600 303.600 443.400 ;
        RECT 319.950 442.800 322.050 443.400 ;
        RECT 326.400 442.050 327.600 452.400 ;
        RECT 355.950 452.400 373.050 453.600 ;
        RECT 355.950 451.950 358.050 452.400 ;
        RECT 370.950 451.950 373.050 452.400 ;
        RECT 505.950 451.950 508.050 454.050 ;
        RECT 586.950 452.400 591.600 454.050 ;
        RECT 703.950 453.600 706.050 454.050 ;
        RECT 709.950 453.600 712.050 454.050 ;
        RECT 703.950 452.400 712.050 453.600 ;
        RECT 586.950 451.950 591.000 452.400 ;
        RECT 703.950 451.950 706.050 452.400 ;
        RECT 709.950 451.950 712.050 452.400 ;
        RECT 745.950 453.600 748.050 454.050 ;
        RECT 763.950 453.600 766.050 454.050 ;
        RECT 780.000 453.600 784.050 454.050 ;
        RECT 745.950 452.400 766.050 453.600 ;
        RECT 745.950 451.950 748.050 452.400 ;
        RECT 763.950 451.950 766.050 452.400 ;
        RECT 779.400 451.950 784.050 453.600 ;
        RECT 829.950 453.600 832.050 454.050 ;
        RECT 850.950 453.600 853.050 454.050 ;
        RECT 829.950 452.400 853.050 453.600 ;
        RECT 829.950 451.950 832.050 452.400 ;
        RECT 850.950 451.950 853.050 452.400 ;
        RECT 331.950 448.950 334.050 451.050 ;
        RECT 364.950 449.100 367.050 451.200 ;
        RECT 400.950 450.600 403.050 451.200 ;
        RECT 436.950 450.600 439.050 451.050 ;
        RECT 457.950 450.600 460.050 451.200 ;
        RECT 400.950 449.400 417.600 450.600 ;
        RECT 400.950 449.100 403.050 449.400 ;
        RECT 332.400 445.050 333.600 448.950 ;
        RECT 331.950 442.950 334.050 445.050 ;
        RECT 352.950 444.600 355.050 445.050 ;
        RECT 365.400 444.600 366.600 449.100 ;
        RECT 352.950 443.400 366.600 444.600 ;
        RECT 382.950 444.600 385.050 444.900 ;
        RECT 406.950 444.600 409.050 445.050 ;
        RECT 382.950 443.400 409.050 444.600 ;
        RECT 416.400 444.600 417.600 449.400 ;
        RECT 436.950 449.400 460.050 450.600 ;
        RECT 436.950 448.950 439.050 449.400 ;
        RECT 457.950 449.100 460.050 449.400 ;
        RECT 466.950 450.750 469.050 451.200 ;
        RECT 484.950 450.750 487.050 451.200 ;
        RECT 466.950 449.550 487.050 450.750 ;
        RECT 466.950 449.100 469.050 449.550 ;
        RECT 484.950 449.100 487.050 449.550 ;
        RECT 458.400 447.600 459.600 449.100 ;
        RECT 458.400 446.400 468.600 447.600 ;
        RECT 427.950 444.600 430.050 445.050 ;
        RECT 416.400 443.400 430.050 444.600 ;
        RECT 352.950 442.950 355.050 443.400 ;
        RECT 382.950 442.800 385.050 443.400 ;
        RECT 406.950 442.950 409.050 443.400 ;
        RECT 427.950 442.950 430.050 443.400 ;
        RECT 433.950 444.600 436.050 444.750 ;
        RECT 442.800 444.600 444.900 445.050 ;
        RECT 433.950 443.400 444.900 444.600 ;
        RECT 433.950 442.650 436.050 443.400 ;
        RECT 442.800 442.950 444.900 443.400 ;
        RECT 445.950 444.450 448.050 444.900 ;
        RECT 454.950 444.450 457.050 444.900 ;
        RECT 445.950 443.250 457.050 444.450 ;
        RECT 467.400 444.600 468.600 446.400 ;
        RECT 467.400 443.400 471.600 444.600 ;
        RECT 445.950 442.800 448.050 443.250 ;
        RECT 454.950 442.800 457.050 443.250 ;
        RECT 310.950 441.600 313.050 442.050 ;
        RECT 302.400 440.400 313.050 441.600 ;
        RECT 310.950 439.950 313.050 440.400 ;
        RECT 322.950 440.400 327.600 442.050 ;
        RECT 334.950 441.600 337.050 442.050 ;
        RECT 343.950 441.600 346.050 442.050 ;
        RECT 334.950 440.400 346.050 441.600 ;
        RECT 470.400 441.600 471.600 443.400 ;
        RECT 493.950 444.450 496.050 444.900 ;
        RECT 502.950 444.450 505.050 444.900 ;
        RECT 493.950 443.250 505.050 444.450 ;
        RECT 506.400 444.600 507.600 451.950 ;
        RECT 514.950 450.600 517.050 451.200 ;
        RECT 523.950 450.600 526.050 451.050 ;
        RECT 514.950 449.400 526.050 450.600 ;
        RECT 514.950 449.100 517.050 449.400 ;
        RECT 523.950 448.950 526.050 449.400 ;
        RECT 556.950 450.750 559.050 451.200 ;
        RECT 562.950 450.750 565.050 451.200 ;
        RECT 556.950 449.550 565.050 450.750 ;
        RECT 556.950 449.100 559.050 449.550 ;
        RECT 562.950 449.100 565.050 449.550 ;
        RECT 571.950 450.600 574.050 451.200 ;
        RECT 643.950 450.600 646.050 451.200 ;
        RECT 658.950 450.600 661.050 451.200 ;
        RECT 571.950 449.400 591.600 450.600 ;
        RECT 571.950 449.100 574.050 449.400 ;
        RECT 557.400 447.600 558.600 449.100 ;
        RECT 554.400 446.400 558.600 447.600 ;
        RECT 554.400 444.900 555.600 446.400 ;
        RECT 590.400 444.900 591.600 449.400 ;
        RECT 629.400 449.400 646.050 450.600 ;
        RECT 517.950 444.600 520.050 444.900 ;
        RECT 506.400 443.400 520.050 444.600 ;
        RECT 493.950 442.800 496.050 443.250 ;
        RECT 502.950 442.800 505.050 443.250 ;
        RECT 517.950 442.800 520.050 443.400 ;
        RECT 523.950 444.300 526.050 444.750 ;
        RECT 529.950 444.300 532.050 444.750 ;
        RECT 523.950 443.100 532.050 444.300 ;
        RECT 523.950 442.650 526.050 443.100 ;
        RECT 529.950 442.650 532.050 443.100 ;
        RECT 553.950 442.800 556.050 444.900 ;
        RECT 565.950 444.450 568.050 444.900 ;
        RECT 580.950 444.450 583.050 444.900 ;
        RECT 565.950 443.250 583.050 444.450 ;
        RECT 565.950 442.800 568.050 443.250 ;
        RECT 580.950 442.800 583.050 443.250 ;
        RECT 589.950 442.800 592.050 444.900 ;
        RECT 629.400 444.750 630.600 449.400 ;
        RECT 643.950 449.100 646.050 449.400 ;
        RECT 647.400 449.400 661.050 450.600 ;
        RECT 647.400 444.900 648.600 449.400 ;
        RECT 658.950 449.100 661.050 449.400 ;
        RECT 664.950 450.600 667.050 451.200 ;
        RECT 679.950 450.600 682.050 451.200 ;
        RECT 664.950 449.400 682.050 450.600 ;
        RECT 664.950 449.100 667.050 449.400 ;
        RECT 679.950 449.100 682.050 449.400 ;
        RECT 685.950 449.100 688.050 451.200 ;
        RECT 628.950 442.650 631.050 444.750 ;
        RECT 646.950 442.800 649.050 444.900 ;
        RECT 686.400 442.050 687.600 449.100 ;
        RECT 688.950 444.600 691.050 444.900 ;
        RECT 694.950 444.600 697.050 445.050 ;
        RECT 700.950 444.600 703.050 444.750 ;
        RECT 688.950 443.400 703.050 444.600 ;
        RECT 688.950 442.800 691.050 443.400 ;
        RECT 694.950 442.950 697.050 443.400 ;
        RECT 700.950 442.650 703.050 443.400 ;
        RECT 724.950 444.600 727.050 444.750 ;
        RECT 730.950 444.600 733.050 445.050 ;
        RECT 754.950 444.600 757.050 444.900 ;
        RECT 763.950 444.600 766.050 445.050 ;
        RECT 724.950 443.400 766.050 444.600 ;
        RECT 724.950 442.650 727.050 443.400 ;
        RECT 730.950 442.950 733.050 443.400 ;
        RECT 754.950 442.800 757.050 443.400 ;
        RECT 763.950 442.950 766.050 443.400 ;
        RECT 475.950 441.600 478.050 442.050 ;
        RECT 470.400 440.400 478.050 441.600 ;
        RECT 322.950 439.950 327.000 440.400 ;
        RECT 334.950 439.950 337.050 440.400 ;
        RECT 343.950 439.950 346.050 440.400 ;
        RECT 475.950 439.950 478.050 440.400 ;
        RECT 637.950 441.600 640.050 442.050 ;
        RECT 661.950 441.600 664.050 442.050 ;
        RECT 637.950 440.400 664.050 441.600 ;
        RECT 637.950 439.950 640.050 440.400 ;
        RECT 661.950 439.950 664.050 440.400 ;
        RECT 685.950 439.950 688.050 442.050 ;
        RECT 37.950 438.600 40.050 439.050 ;
        RECT 73.800 438.600 75.900 439.050 ;
        RECT 37.950 437.400 75.900 438.600 ;
        RECT 37.950 436.950 40.050 437.400 ;
        RECT 73.800 436.950 75.900 437.400 ;
        RECT 76.950 438.600 79.050 439.050 ;
        RECT 92.400 438.600 93.600 439.950 ;
        RECT 76.950 437.400 93.600 438.600 ;
        RECT 232.950 438.600 235.050 439.050 ;
        RECT 241.950 438.600 244.050 439.050 ;
        RECT 298.950 438.600 301.050 439.050 ;
        RECT 232.950 437.400 301.050 438.600 ;
        RECT 76.950 436.950 79.050 437.400 ;
        RECT 232.950 436.950 235.050 437.400 ;
        RECT 241.950 436.950 244.050 437.400 ;
        RECT 298.950 436.950 301.050 437.400 ;
        RECT 313.950 438.600 316.050 439.050 ;
        RECT 394.950 438.600 397.050 439.050 ;
        RECT 313.950 437.400 397.050 438.600 ;
        RECT 313.950 436.950 316.050 437.400 ;
        RECT 394.950 436.950 397.050 437.400 ;
        RECT 427.950 438.600 430.050 439.050 ;
        RECT 463.950 438.600 466.050 439.050 ;
        RECT 427.950 437.400 466.050 438.600 ;
        RECT 427.950 436.950 430.050 437.400 ;
        RECT 463.950 436.950 466.050 437.400 ;
        RECT 511.950 438.600 514.050 439.050 ;
        RECT 619.950 438.600 622.050 439.050 ;
        RECT 511.950 437.400 622.050 438.600 ;
        RECT 511.950 436.950 514.050 437.400 ;
        RECT 619.950 436.950 622.050 437.400 ;
        RECT 655.950 438.600 658.050 439.050 ;
        RECT 670.950 438.600 673.050 439.050 ;
        RECT 655.950 437.400 673.050 438.600 ;
        RECT 655.950 436.950 658.050 437.400 ;
        RECT 670.950 436.950 673.050 437.400 ;
        RECT 706.950 438.600 709.050 439.050 ;
        RECT 766.950 438.600 769.050 439.050 ;
        RECT 772.950 438.600 775.050 439.050 ;
        RECT 706.950 437.400 775.050 438.600 ;
        RECT 779.400 438.600 780.600 451.950 ;
        RECT 796.950 450.600 799.050 451.050 ;
        RECT 782.400 449.400 799.050 450.600 ;
        RECT 782.400 444.900 783.600 449.400 ;
        RECT 796.950 448.950 799.050 449.400 ;
        RECT 781.950 442.800 784.050 444.900 ;
        RECT 784.950 441.600 787.050 442.050 ;
        RECT 811.950 441.600 814.050 442.050 ;
        RECT 784.950 440.400 814.050 441.600 ;
        RECT 784.950 439.950 787.050 440.400 ;
        RECT 811.950 439.950 814.050 440.400 ;
        RECT 790.800 438.600 792.900 439.050 ;
        RECT 779.400 437.400 792.900 438.600 ;
        RECT 706.950 436.950 709.050 437.400 ;
        RECT 766.950 436.950 769.050 437.400 ;
        RECT 772.950 436.950 775.050 437.400 ;
        RECT 790.800 436.950 792.900 437.400 ;
        RECT 793.950 438.600 796.050 439.050 ;
        RECT 826.950 438.600 829.050 439.050 ;
        RECT 793.950 437.400 829.050 438.600 ;
        RECT 793.950 436.950 796.050 437.400 ;
        RECT 826.950 436.950 829.050 437.400 ;
        RECT 28.950 435.600 31.050 436.050 ;
        RECT 64.950 435.600 67.050 436.050 ;
        RECT 28.950 434.400 67.050 435.600 ;
        RECT 28.950 433.950 31.050 434.400 ;
        RECT 64.950 433.950 67.050 434.400 ;
        RECT 79.950 435.600 82.050 436.050 ;
        RECT 127.950 435.600 130.050 436.050 ;
        RECT 79.950 434.400 130.050 435.600 ;
        RECT 79.950 433.950 82.050 434.400 ;
        RECT 127.950 433.950 130.050 434.400 ;
        RECT 133.950 435.600 136.050 436.050 ;
        RECT 157.950 435.600 160.050 436.050 ;
        RECT 133.950 434.400 160.050 435.600 ;
        RECT 133.950 433.950 136.050 434.400 ;
        RECT 157.950 433.950 160.050 434.400 ;
        RECT 208.950 435.600 211.050 436.050 ;
        RECT 233.400 435.600 234.600 436.950 ;
        RECT 208.950 434.400 234.600 435.600 ;
        RECT 685.950 435.600 688.050 436.050 ;
        RECT 715.950 435.600 718.050 436.050 ;
        RECT 736.950 435.600 739.050 436.050 ;
        RECT 799.950 435.600 802.050 436.050 ;
        RECT 685.950 434.400 802.050 435.600 ;
        RECT 208.950 433.950 211.050 434.400 ;
        RECT 685.950 433.950 688.050 434.400 ;
        RECT 715.950 433.950 718.050 434.400 ;
        RECT 736.950 433.950 739.050 434.400 ;
        RECT 799.950 433.950 802.050 434.400 ;
        RECT 61.950 432.600 64.050 433.050 ;
        RECT 103.950 432.600 106.050 433.050 ;
        RECT 61.950 431.400 106.050 432.600 ;
        RECT 61.950 430.950 64.050 431.400 ;
        RECT 103.950 430.950 106.050 431.400 ;
        RECT 181.950 432.600 184.050 433.050 ;
        RECT 265.950 432.600 268.050 433.050 ;
        RECT 181.950 431.400 268.050 432.600 ;
        RECT 181.950 430.950 184.050 431.400 ;
        RECT 265.950 430.950 268.050 431.400 ;
        RECT 271.950 432.600 274.050 433.050 ;
        RECT 295.950 432.600 298.050 433.050 ;
        RECT 271.950 431.400 298.050 432.600 ;
        RECT 271.950 430.950 274.050 431.400 ;
        RECT 295.950 430.950 298.050 431.400 ;
        RECT 466.950 432.600 469.050 433.050 ;
        RECT 499.950 432.600 502.050 433.050 ;
        RECT 466.950 431.400 502.050 432.600 ;
        RECT 466.950 430.950 469.050 431.400 ;
        RECT 499.950 430.950 502.050 431.400 ;
        RECT 610.950 432.600 613.050 433.050 ;
        RECT 616.950 432.600 619.050 433.050 ;
        RECT 682.950 432.600 685.050 433.050 ;
        RECT 610.950 431.400 685.050 432.600 ;
        RECT 610.950 430.950 613.050 431.400 ;
        RECT 616.950 430.950 619.050 431.400 ;
        RECT 682.950 430.950 685.050 431.400 ;
        RECT 781.950 432.600 784.050 433.050 ;
        RECT 796.950 432.600 799.050 433.050 ;
        RECT 781.950 431.400 799.050 432.600 ;
        RECT 781.950 430.950 784.050 431.400 ;
        RECT 796.950 430.950 799.050 431.400 ;
        RECT 64.950 429.600 67.050 430.050 ;
        RECT 97.950 429.600 100.050 430.050 ;
        RECT 64.950 428.400 100.050 429.600 ;
        RECT 64.950 427.950 67.050 428.400 ;
        RECT 97.950 427.950 100.050 428.400 ;
        RECT 214.950 429.600 217.050 430.050 ;
        RECT 256.950 429.600 259.050 430.050 ;
        RECT 214.950 428.400 259.050 429.600 ;
        RECT 214.950 427.950 217.050 428.400 ;
        RECT 256.950 427.950 259.050 428.400 ;
        RECT 268.950 429.600 271.050 430.050 ;
        RECT 280.950 429.600 283.050 430.050 ;
        RECT 268.950 428.400 283.050 429.600 ;
        RECT 268.950 427.950 271.050 428.400 ;
        RECT 280.950 427.950 283.050 428.400 ;
        RECT 325.950 429.600 328.050 430.050 ;
        RECT 352.950 429.600 355.050 430.050 ;
        RECT 325.950 428.400 355.050 429.600 ;
        RECT 325.950 427.950 328.050 428.400 ;
        RECT 352.950 427.950 355.050 428.400 ;
        RECT 460.950 429.600 463.050 430.050 ;
        RECT 523.950 429.600 526.050 430.050 ;
        RECT 460.950 428.400 526.050 429.600 ;
        RECT 460.950 427.950 463.050 428.400 ;
        RECT 523.950 427.950 526.050 428.400 ;
        RECT 619.950 429.600 622.050 430.050 ;
        RECT 784.950 429.600 787.050 430.050 ;
        RECT 619.950 428.400 787.050 429.600 ;
        RECT 619.950 427.950 622.050 428.400 ;
        RECT 784.950 427.950 787.050 428.400 ;
        RECT 160.950 426.600 163.050 427.050 ;
        RECT 175.950 426.600 178.050 427.050 ;
        RECT 160.950 425.400 178.050 426.600 ;
        RECT 160.950 424.950 163.050 425.400 ;
        RECT 175.950 424.950 178.050 425.400 ;
        RECT 388.950 426.600 391.050 427.050 ;
        RECT 412.950 426.600 415.050 427.050 ;
        RECT 388.950 425.400 415.050 426.600 ;
        RECT 388.950 424.950 391.050 425.400 ;
        RECT 412.950 424.950 415.050 425.400 ;
        RECT 463.950 426.600 466.050 427.050 ;
        RECT 517.950 426.600 520.050 427.050 ;
        RECT 463.950 425.400 520.050 426.600 ;
        RECT 463.950 424.950 466.050 425.400 ;
        RECT 517.950 424.950 520.050 425.400 ;
        RECT 766.950 426.600 769.050 427.050 ;
        RECT 790.950 426.600 793.050 427.050 ;
        RECT 766.950 425.400 793.050 426.600 ;
        RECT 766.950 424.950 769.050 425.400 ;
        RECT 790.950 424.950 793.050 425.400 ;
        RECT 802.950 426.600 805.050 427.050 ;
        RECT 829.950 426.600 832.050 427.050 ;
        RECT 802.950 425.400 832.050 426.600 ;
        RECT 802.950 424.950 805.050 425.400 ;
        RECT 829.950 424.950 832.050 425.400 ;
        RECT 13.950 423.600 16.050 424.050 ;
        RECT 25.950 423.600 28.050 424.050 ;
        RECT 13.950 422.400 28.050 423.600 ;
        RECT 13.950 421.950 16.050 422.400 ;
        RECT 25.950 421.950 28.050 422.400 ;
        RECT 31.950 423.600 34.050 424.050 ;
        RECT 40.950 423.600 43.050 424.050 ;
        RECT 31.950 422.400 43.050 423.600 ;
        RECT 31.950 421.950 34.050 422.400 ;
        RECT 40.950 421.950 43.050 422.400 ;
        RECT 127.950 423.600 130.050 424.050 ;
        RECT 154.950 423.600 157.050 424.050 ;
        RECT 184.950 423.600 187.050 424.050 ;
        RECT 127.950 422.400 187.050 423.600 ;
        RECT 127.950 421.950 130.050 422.400 ;
        RECT 154.950 421.950 157.050 422.400 ;
        RECT 184.950 421.950 187.050 422.400 ;
        RECT 256.950 423.600 259.050 424.050 ;
        RECT 280.950 423.600 283.050 424.050 ;
        RECT 256.950 422.400 283.050 423.600 ;
        RECT 256.950 421.950 259.050 422.400 ;
        RECT 280.950 421.950 283.050 422.400 ;
        RECT 400.950 423.600 403.050 424.050 ;
        RECT 415.950 423.600 418.050 424.050 ;
        RECT 400.950 422.400 418.050 423.600 ;
        RECT 400.950 421.950 403.050 422.400 ;
        RECT 415.950 421.950 418.050 422.400 ;
        RECT 565.950 423.600 568.050 424.050 ;
        RECT 589.950 423.600 592.050 424.050 ;
        RECT 604.950 423.600 607.050 424.050 ;
        RECT 565.950 422.400 607.050 423.600 ;
        RECT 565.950 421.950 568.050 422.400 ;
        RECT 589.950 421.950 592.050 422.400 ;
        RECT 604.950 421.950 607.050 422.400 ;
        RECT 616.950 423.600 619.050 424.050 ;
        RECT 628.950 423.600 631.050 424.050 ;
        RECT 616.950 422.400 631.050 423.600 ;
        RECT 616.950 421.950 619.050 422.400 ;
        RECT 628.950 421.950 631.050 422.400 ;
        RECT 652.950 423.600 655.050 424.050 ;
        RECT 703.950 423.600 706.050 424.050 ;
        RECT 652.950 422.400 706.050 423.600 ;
        RECT 652.950 421.950 655.050 422.400 ;
        RECT 703.950 421.950 706.050 422.400 ;
        RECT 805.950 423.600 808.050 424.050 ;
        RECT 826.950 423.600 829.050 424.050 ;
        RECT 805.950 422.400 829.050 423.600 ;
        RECT 805.950 421.950 808.050 422.400 ;
        RECT 826.950 421.950 829.050 422.400 ;
        RECT 4.950 420.600 7.050 421.050 ;
        RECT 10.950 420.600 13.050 421.050 ;
        RECT 4.950 419.400 13.050 420.600 ;
        RECT 4.950 418.950 7.050 419.400 ;
        RECT 10.950 418.950 13.050 419.400 ;
        RECT 34.950 420.600 37.050 421.050 ;
        RECT 46.950 420.600 49.050 421.050 ;
        RECT 52.950 420.600 55.050 421.050 ;
        RECT 34.950 419.400 55.050 420.600 ;
        RECT 34.950 418.950 37.050 419.400 ;
        RECT 46.950 418.950 49.050 419.400 ;
        RECT 52.950 418.950 55.050 419.400 ;
        RECT 205.950 420.600 208.050 421.050 ;
        RECT 217.950 420.600 220.050 421.050 ;
        RECT 223.950 420.600 226.050 421.050 ;
        RECT 205.950 419.400 213.600 420.600 ;
        RECT 205.950 418.950 208.050 419.400 ;
        RECT 16.950 416.250 19.050 418.350 ;
        RECT 21.000 417.600 25.050 418.050 ;
        RECT 17.400 412.050 18.600 416.250 ;
        RECT 20.400 415.950 25.050 417.600 ;
        RECT 28.950 415.950 31.050 418.050 ;
        RECT 70.950 417.600 73.050 418.200 ;
        RECT 88.950 417.600 91.050 418.350 ;
        RECT 50.400 416.400 73.050 417.600 ;
        RECT 20.400 412.050 21.600 415.950 ;
        RECT 4.950 411.600 7.050 412.050 ;
        RECT 13.800 411.600 15.900 412.050 ;
        RECT 4.950 410.400 15.900 411.600 ;
        RECT 4.950 409.950 7.050 410.400 ;
        RECT 13.800 409.950 15.900 410.400 ;
        RECT 16.800 409.950 18.900 412.050 ;
        RECT 19.950 409.950 22.050 412.050 ;
        RECT 29.400 411.600 30.600 415.950 ;
        RECT 50.400 412.050 51.600 416.400 ;
        RECT 70.950 416.100 73.050 416.400 ;
        RECT 74.400 416.400 91.050 417.600 ;
        RECT 74.400 414.600 75.600 416.400 ;
        RECT 88.950 416.250 91.050 416.400 ;
        RECT 94.950 416.250 97.050 418.350 ;
        RECT 103.950 417.600 106.050 418.050 ;
        RECT 109.950 417.600 112.050 418.350 ;
        RECT 103.950 416.400 112.050 417.600 ;
        RECT 68.400 413.400 75.600 414.600 ;
        RECT 31.950 411.600 34.050 411.900 ;
        RECT 29.400 410.400 34.050 411.600 ;
        RECT 20.400 408.600 21.600 409.950 ;
        RECT 31.950 409.800 34.050 410.400 ;
        RECT 37.950 411.600 40.050 412.050 ;
        RECT 49.950 411.600 52.050 412.050 ;
        RECT 68.400 411.900 69.600 413.400 ;
        RECT 95.400 412.050 96.600 416.250 ;
        RECT 103.950 415.950 106.050 416.400 ;
        RECT 109.950 416.250 112.050 416.400 ;
        RECT 115.950 416.250 118.050 418.350 ;
        RECT 136.950 417.750 139.050 418.200 ;
        RECT 142.950 417.750 145.050 418.200 ;
        RECT 136.950 416.550 145.050 417.750 ;
        RECT 148.950 417.600 151.050 418.200 ;
        RECT 37.950 410.400 52.050 411.600 ;
        RECT 37.950 409.950 40.050 410.400 ;
        RECT 49.950 409.950 52.050 410.400 ;
        RECT 67.950 409.800 70.050 411.900 ;
        RECT 94.800 409.950 96.900 412.050 ;
        RECT 97.950 411.600 100.050 412.050 ;
        RECT 116.400 411.600 117.600 416.250 ;
        RECT 136.950 416.100 139.050 416.550 ;
        RECT 142.950 416.100 145.050 416.550 ;
        RECT 146.400 416.400 151.050 417.600 ;
        RECT 146.400 414.600 147.600 416.400 ;
        RECT 148.950 416.100 151.050 416.400 ;
        RECT 154.950 414.600 157.050 418.050 ;
        RECT 163.950 416.100 166.050 418.200 ;
        RECT 187.950 417.600 190.050 418.350 ;
        RECT 202.950 417.600 205.050 418.350 ;
        RECT 167.400 416.400 190.050 417.600 ;
        RECT 134.400 414.000 147.600 414.600 ;
        RECT 133.950 413.400 147.600 414.000 ;
        RECT 152.400 414.000 157.050 414.600 ;
        RECT 152.400 413.400 156.600 414.000 ;
        RECT 130.800 411.600 132.900 411.900 ;
        RECT 97.950 410.400 132.900 411.600 ;
        RECT 97.950 409.950 100.050 410.400 ;
        RECT 130.800 409.800 132.900 410.400 ;
        RECT 133.950 409.950 136.050 413.400 ;
        RECT 152.400 411.900 153.600 413.400 ;
        RECT 164.400 412.050 165.600 416.100 ;
        RECT 151.950 409.800 154.050 411.900 ;
        RECT 160.950 410.400 165.600 412.050 ;
        RECT 160.950 409.950 165.000 410.400 ;
        RECT 167.400 409.050 168.600 416.400 ;
        RECT 187.950 416.250 190.050 416.400 ;
        RECT 191.400 416.400 205.050 417.600 ;
        RECT 191.400 414.600 192.600 416.400 ;
        RECT 202.950 416.250 205.050 416.400 ;
        RECT 188.400 414.000 192.600 414.600 ;
        RECT 187.950 413.400 192.600 414.000 ;
        RECT 187.950 409.950 190.050 413.400 ;
        RECT 212.400 412.050 213.600 419.400 ;
        RECT 217.950 419.400 226.050 420.600 ;
        RECT 217.950 418.950 220.050 419.400 ;
        RECT 223.950 418.950 226.050 419.400 ;
        RECT 247.950 420.600 250.050 421.050 ;
        RECT 253.950 420.600 256.050 421.050 ;
        RECT 247.950 419.400 256.050 420.600 ;
        RECT 247.950 418.950 250.050 419.400 ;
        RECT 253.950 418.950 256.050 419.400 ;
        RECT 268.950 418.950 271.050 421.050 ;
        RECT 283.950 420.600 286.050 421.050 ;
        RECT 289.950 420.600 292.050 421.050 ;
        RECT 316.950 420.600 319.050 421.050 ;
        RECT 388.950 420.600 391.050 421.200 ;
        RECT 622.950 421.050 625.050 421.200 ;
        RECT 283.950 419.400 391.050 420.600 ;
        RECT 283.950 418.950 286.050 419.400 ;
        RECT 289.950 418.950 292.050 419.400 ;
        RECT 316.950 418.950 319.050 419.400 ;
        RECT 388.950 419.100 391.050 419.400 ;
        RECT 412.950 420.600 415.050 421.050 ;
        RECT 622.950 420.600 627.000 421.050 ;
        RECT 742.950 420.600 745.050 421.050 ;
        RECT 760.950 420.600 763.050 421.050 ;
        RECT 787.950 420.600 790.050 421.050 ;
        RECT 412.950 419.400 444.600 420.600 ;
        RECT 412.950 418.950 415.050 419.400 ;
        RECT 226.950 417.600 229.050 418.350 ;
        RECT 238.950 417.600 241.050 418.050 ;
        RECT 265.950 417.600 268.050 418.200 ;
        RECT 226.950 416.400 241.050 417.600 ;
        RECT 226.950 416.250 229.050 416.400 ;
        RECT 238.950 415.950 241.050 416.400 ;
        RECT 254.400 416.400 268.050 417.600 ;
        RECT 254.400 412.050 255.600 416.400 ;
        RECT 265.950 416.100 268.050 416.400 ;
        RECT 211.950 409.950 214.050 412.050 ;
        RECT 229.950 411.600 232.050 412.050 ;
        RECT 235.950 411.600 238.050 412.050 ;
        RECT 244.950 411.600 247.050 412.050 ;
        RECT 229.950 410.400 247.050 411.600 ;
        RECT 229.950 409.950 232.050 410.400 ;
        RECT 235.950 409.950 238.050 410.400 ;
        RECT 244.950 409.950 247.050 410.400 ;
        RECT 253.950 409.950 256.050 412.050 ;
        RECT 269.400 411.600 270.600 418.950 ;
        RECT 271.950 417.600 274.050 418.200 ;
        RECT 304.950 417.600 307.050 418.350 ;
        RECT 271.950 416.400 285.600 417.600 ;
        RECT 271.950 416.100 274.050 416.400 ;
        RECT 274.950 411.600 277.050 412.050 ;
        RECT 284.400 411.900 285.600 416.400 ;
        RECT 304.950 416.400 333.600 417.600 ;
        RECT 304.950 416.250 307.050 416.400 ;
        RECT 332.400 414.600 333.600 416.400 ;
        RECT 337.950 416.100 340.050 418.200 ;
        RECT 343.950 417.750 346.050 418.200 ;
        RECT 364.950 417.750 367.050 418.200 ;
        RECT 343.950 416.550 367.050 417.750 ;
        RECT 343.950 416.100 346.050 416.550 ;
        RECT 364.950 416.100 367.050 416.550 ;
        RECT 376.950 417.600 379.050 418.200 ;
        RECT 388.950 417.600 391.050 418.050 ;
        RECT 376.950 416.400 391.050 417.600 ;
        RECT 376.950 416.100 379.050 416.400 ;
        RECT 332.400 413.400 336.600 414.600 ;
        RECT 269.400 410.400 277.050 411.600 ;
        RECT 274.950 409.950 277.050 410.400 ;
        RECT 283.950 409.800 286.050 411.900 ;
        RECT 289.950 411.600 292.050 412.050 ;
        RECT 295.950 411.600 298.050 412.050 ;
        RECT 289.950 410.400 298.050 411.600 ;
        RECT 289.950 409.950 292.050 410.400 ;
        RECT 295.950 409.950 298.050 410.400 ;
        RECT 319.950 411.600 322.050 411.900 ;
        RECT 328.950 411.600 331.050 412.050 ;
        RECT 335.400 411.900 336.600 413.400 ;
        RECT 319.950 410.400 331.050 411.600 ;
        RECT 319.950 409.800 322.050 410.400 ;
        RECT 328.950 409.950 331.050 410.400 ;
        RECT 334.950 409.800 337.050 411.900 ;
        RECT 338.400 411.600 339.600 416.100 ;
        RECT 388.950 415.950 391.050 416.400 ;
        RECT 400.800 415.950 402.900 418.050 ;
        RECT 403.950 416.100 406.050 418.200 ;
        RECT 409.950 417.600 412.050 418.200 ;
        RECT 439.950 417.600 442.050 418.050 ;
        RECT 409.950 416.400 442.050 417.600 ;
        RECT 443.400 417.600 444.600 419.400 ;
        RECT 622.950 419.100 627.600 420.600 ;
        RECT 624.000 418.950 627.600 419.100 ;
        RECT 742.950 419.400 763.050 420.600 ;
        RECT 742.950 418.950 745.050 419.400 ;
        RECT 760.950 418.950 763.050 419.400 ;
        RECT 776.400 419.400 790.050 420.600 ;
        RECT 448.950 417.600 451.050 418.200 ;
        RECT 457.950 417.600 460.050 418.050 ;
        RECT 443.400 416.400 460.050 417.600 ;
        RECT 409.950 416.100 412.050 416.400 ;
        RECT 358.950 411.600 361.050 411.900 ;
        RECT 338.400 410.400 361.050 411.600 ;
        RECT 358.950 409.800 361.050 410.400 ;
        RECT 364.950 411.600 367.050 412.050 ;
        RECT 391.950 411.600 394.050 411.900 ;
        RECT 364.950 410.400 394.050 411.600 ;
        RECT 401.400 411.600 402.600 415.950 ;
        RECT 404.400 414.600 405.600 416.100 ;
        RECT 439.950 415.950 442.050 416.400 ;
        RECT 448.950 416.100 451.050 416.400 ;
        RECT 457.950 415.950 460.050 416.400 ;
        RECT 547.950 417.900 550.050 418.350 ;
        RECT 556.950 417.900 559.050 418.350 ;
        RECT 547.950 416.700 559.050 417.900 ;
        RECT 547.950 416.250 550.050 416.700 ;
        RECT 556.950 416.250 559.050 416.700 ;
        RECT 454.950 414.600 457.050 415.050 ;
        RECT 565.950 414.600 568.050 418.050 ;
        RECT 571.950 416.100 574.050 418.200 ;
        RECT 622.950 417.600 625.050 418.050 ;
        RECT 608.400 416.400 625.050 417.600 ;
        RECT 404.400 413.400 457.050 414.600 ;
        RECT 454.950 412.950 457.050 413.400 ;
        RECT 563.400 414.000 568.050 414.600 ;
        RECT 563.400 413.400 567.600 414.000 ;
        RECT 412.950 411.600 415.050 411.900 ;
        RECT 401.400 410.400 415.050 411.600 ;
        RECT 364.950 409.950 367.050 410.400 ;
        RECT 391.950 409.800 394.050 410.400 ;
        RECT 412.950 409.800 415.050 410.400 ;
        RECT 430.950 411.450 433.050 411.900 ;
        RECT 439.950 411.450 442.050 411.900 ;
        RECT 430.950 410.250 442.050 411.450 ;
        RECT 430.950 409.800 433.050 410.250 ;
        RECT 439.950 409.800 442.050 410.250 ;
        RECT 457.950 411.600 460.050 412.050 ;
        RECT 463.950 411.600 466.050 412.050 ;
        RECT 457.950 410.400 466.050 411.600 ;
        RECT 457.950 409.950 460.050 410.400 ;
        RECT 463.950 409.950 466.050 410.400 ;
        RECT 553.950 411.600 556.050 412.050 ;
        RECT 563.400 411.600 564.600 413.400 ;
        RECT 553.950 410.400 564.600 411.600 ;
        RECT 565.950 411.600 568.050 412.050 ;
        RECT 572.400 411.600 573.600 416.100 ;
        RECT 565.950 410.400 573.600 411.600 ;
        RECT 592.950 411.600 595.050 411.900 ;
        RECT 608.400 411.600 609.600 416.400 ;
        RECT 622.950 415.950 625.050 416.400 ;
        RECT 626.400 411.900 627.600 418.950 ;
        RECT 640.950 417.750 643.050 418.200 ;
        RECT 649.950 417.750 652.050 418.200 ;
        RECT 640.950 416.550 652.050 417.750 ;
        RECT 640.950 416.100 643.050 416.550 ;
        RECT 649.950 416.100 652.050 416.550 ;
        RECT 682.950 417.600 685.050 418.350 ;
        RECT 691.950 417.600 694.050 418.050 ;
        RECT 682.950 416.400 694.050 417.600 ;
        RECT 682.950 416.250 685.050 416.400 ;
        RECT 691.950 415.950 694.050 416.400 ;
        RECT 697.950 416.100 700.050 418.200 ;
        RECT 712.950 417.600 715.050 418.050 ;
        RECT 724.950 417.600 727.050 418.200 ;
        RECT 712.950 416.400 727.050 417.600 ;
        RECT 592.950 410.400 609.600 411.600 ;
        RECT 553.950 409.950 556.050 410.400 ;
        RECT 565.950 409.950 568.050 410.400 ;
        RECT 592.950 409.800 595.050 410.400 ;
        RECT 625.950 409.800 628.050 411.900 ;
        RECT 649.950 411.600 652.050 412.050 ;
        RECT 679.950 411.600 682.050 412.050 ;
        RECT 649.950 410.400 682.050 411.600 ;
        RECT 649.950 409.950 652.050 410.400 ;
        RECT 679.950 409.950 682.050 410.400 ;
        RECT 685.950 411.600 688.050 412.050 ;
        RECT 698.400 411.600 699.600 416.100 ;
        RECT 712.950 415.950 715.050 416.400 ;
        RECT 724.950 416.100 727.050 416.400 ;
        RECT 736.950 417.600 739.050 418.050 ;
        RECT 745.950 417.600 748.050 418.350 ;
        RECT 736.950 416.400 748.050 417.600 ;
        RECT 736.950 415.950 739.050 416.400 ;
        RECT 745.950 416.250 748.050 416.400 ;
        RECT 776.400 412.050 777.600 419.400 ;
        RECT 787.950 418.950 790.050 419.400 ;
        RECT 838.950 420.600 841.050 421.050 ;
        RECT 838.950 419.400 846.600 420.600 ;
        RECT 838.950 418.950 841.050 419.400 ;
        RECT 789.000 417.600 793.050 418.050 ;
        RECT 788.400 415.950 793.050 417.600 ;
        RECT 796.950 415.950 799.050 418.050 ;
        RECT 814.950 417.750 817.050 418.200 ;
        RECT 835.950 417.750 838.050 418.200 ;
        RECT 814.950 416.550 838.050 417.750 ;
        RECT 814.950 416.100 817.050 416.550 ;
        RECT 835.950 416.100 838.050 416.550 ;
        RECT 788.400 412.050 789.600 415.950 ;
        RECT 685.950 410.400 699.600 411.600 ;
        RECT 721.950 411.600 724.050 411.900 ;
        RECT 754.950 411.600 757.050 412.050 ;
        RECT 721.950 410.400 757.050 411.600 ;
        RECT 685.950 409.950 688.050 410.400 ;
        RECT 721.950 409.800 724.050 410.400 ;
        RECT 754.950 409.950 757.050 410.400 ;
        RECT 763.950 411.600 766.050 412.050 ;
        RECT 769.950 411.600 772.050 412.050 ;
        RECT 763.950 410.400 772.050 411.600 ;
        RECT 763.950 409.950 766.050 410.400 ;
        RECT 769.950 409.950 772.050 410.400 ;
        RECT 775.950 409.950 778.050 412.050 ;
        RECT 787.950 409.950 790.050 412.050 ;
        RECT 797.400 411.600 798.600 415.950 ;
        RECT 845.400 412.050 846.600 419.400 ;
        RECT 847.950 417.600 850.050 418.050 ;
        RECT 859.950 417.600 862.050 418.050 ;
        RECT 847.950 416.400 862.050 417.600 ;
        RECT 847.950 415.950 850.050 416.400 ;
        RECT 859.950 415.950 862.050 416.400 ;
        RECT 823.950 411.600 826.050 411.900 ;
        RECT 797.400 410.400 826.050 411.600 ;
        RECT 823.950 409.800 826.050 410.400 ;
        RECT 844.950 409.950 847.050 412.050 ;
        RECT 55.950 408.600 58.050 409.050 ;
        RECT 20.400 407.400 58.050 408.600 ;
        RECT 55.950 406.950 58.050 407.400 ;
        RECT 91.950 408.600 94.050 409.050 ;
        RECT 91.950 407.400 147.600 408.600 ;
        RECT 91.950 406.950 94.050 407.400 ;
        RECT 146.400 406.050 147.600 407.400 ;
        RECT 163.950 407.400 168.600 409.050 ;
        RECT 301.950 408.600 304.050 409.050 ;
        RECT 310.950 408.600 313.050 409.050 ;
        RECT 340.950 408.600 343.050 409.050 ;
        RECT 301.950 407.400 343.050 408.600 ;
        RECT 163.950 406.950 168.000 407.400 ;
        RECT 301.950 406.950 304.050 407.400 ;
        RECT 310.950 406.950 313.050 407.400 ;
        RECT 340.950 406.950 343.050 407.400 ;
        RECT 391.950 408.600 394.050 408.750 ;
        RECT 397.950 408.600 400.050 409.050 ;
        RECT 391.950 407.400 400.050 408.600 ;
        RECT 391.950 406.650 394.050 407.400 ;
        RECT 397.950 406.950 400.050 407.400 ;
        RECT 454.950 408.600 457.050 409.050 ;
        RECT 469.950 408.600 472.050 409.050 ;
        RECT 454.950 407.400 472.050 408.600 ;
        RECT 454.950 406.950 457.050 407.400 ;
        RECT 469.950 406.950 472.050 407.400 ;
        RECT 577.950 408.600 580.050 409.050 ;
        RECT 604.950 408.600 607.050 409.050 ;
        RECT 631.950 408.600 634.050 409.050 ;
        RECT 718.950 408.600 721.050 408.900 ;
        RECT 757.950 408.600 760.050 409.050 ;
        RECT 799.950 408.600 802.050 409.050 ;
        RECT 814.950 408.600 817.050 409.050 ;
        RECT 577.950 407.400 817.050 408.600 ;
        RECT 577.950 406.950 580.050 407.400 ;
        RECT 604.950 406.950 607.050 407.400 ;
        RECT 631.950 406.950 634.050 407.400 ;
        RECT 718.950 406.800 721.050 407.400 ;
        RECT 757.950 406.950 760.050 407.400 ;
        RECT 799.950 406.950 802.050 407.400 ;
        RECT 814.950 406.950 817.050 407.400 ;
        RECT 61.950 405.600 64.050 406.050 ;
        RECT 73.950 405.600 76.050 406.050 ;
        RECT 61.950 404.400 76.050 405.600 ;
        RECT 61.950 403.950 64.050 404.400 ;
        RECT 73.950 403.950 76.050 404.400 ;
        RECT 94.950 405.600 97.050 406.050 ;
        RECT 118.950 405.600 121.050 406.050 ;
        RECT 94.950 404.400 121.050 405.600 ;
        RECT 94.950 403.950 97.050 404.400 ;
        RECT 118.950 403.950 121.050 404.400 ;
        RECT 145.950 405.600 148.050 406.050 ;
        RECT 166.950 405.600 169.050 406.050 ;
        RECT 145.950 404.400 169.050 405.600 ;
        RECT 145.950 403.950 148.050 404.400 ;
        RECT 166.950 403.950 169.050 404.400 ;
        RECT 211.950 405.600 214.050 406.050 ;
        RECT 250.950 405.600 253.050 406.050 ;
        RECT 211.950 404.400 253.050 405.600 ;
        RECT 211.950 403.950 214.050 404.400 ;
        RECT 250.950 403.950 253.050 404.400 ;
        RECT 397.950 405.600 400.050 405.900 ;
        RECT 421.950 405.600 424.050 406.050 ;
        RECT 481.950 405.600 484.050 406.050 ;
        RECT 487.950 405.600 490.050 406.050 ;
        RECT 397.950 404.400 490.050 405.600 ;
        RECT 397.950 403.800 400.050 404.400 ;
        RECT 421.950 403.950 424.050 404.400 ;
        RECT 481.950 403.950 484.050 404.400 ;
        RECT 487.950 403.950 490.050 404.400 ;
        RECT 562.950 405.600 565.050 406.050 ;
        RECT 598.950 405.600 601.050 406.050 ;
        RECT 562.950 404.400 601.050 405.600 ;
        RECT 562.950 403.950 565.050 404.400 ;
        RECT 598.950 403.950 601.050 404.400 ;
        RECT 691.950 405.600 694.050 406.050 ;
        RECT 706.950 405.600 709.050 406.050 ;
        RECT 691.950 404.400 709.050 405.600 ;
        RECT 691.950 403.950 694.050 404.400 ;
        RECT 706.950 403.950 709.050 404.400 ;
        RECT 715.950 405.600 718.050 406.050 ;
        RECT 727.950 405.600 730.050 406.050 ;
        RECT 715.950 404.400 730.050 405.600 ;
        RECT 715.950 403.950 718.050 404.400 ;
        RECT 727.950 403.950 730.050 404.400 ;
        RECT 748.950 405.600 751.050 406.050 ;
        RECT 772.800 405.600 774.900 406.050 ;
        RECT 748.950 404.400 774.900 405.600 ;
        RECT 748.950 403.950 751.050 404.400 ;
        RECT 772.800 403.950 774.900 404.400 ;
        RECT 775.950 405.600 778.050 406.050 ;
        RECT 805.950 405.600 808.050 406.050 ;
        RECT 775.950 404.400 808.050 405.600 ;
        RECT 775.950 403.950 778.050 404.400 ;
        RECT 805.950 403.950 808.050 404.400 ;
        RECT 190.950 402.600 193.050 403.050 ;
        RECT 289.950 402.600 292.050 403.050 ;
        RECT 742.950 402.600 745.050 403.050 ;
        RECT 190.950 401.400 292.050 402.600 ;
        RECT 190.950 400.950 193.050 401.400 ;
        RECT 289.950 400.950 292.050 401.400 ;
        RECT 734.400 401.400 745.050 402.600 ;
        RECT 145.950 399.600 148.050 400.050 ;
        RECT 157.950 399.600 160.050 400.050 ;
        RECT 217.950 399.600 220.050 400.050 ;
        RECT 145.950 398.400 220.050 399.600 ;
        RECT 145.950 397.950 148.050 398.400 ;
        RECT 157.950 397.950 160.050 398.400 ;
        RECT 217.950 397.950 220.050 398.400 ;
        RECT 673.950 399.600 676.050 400.050 ;
        RECT 700.950 399.600 703.050 400.050 ;
        RECT 673.950 398.400 703.050 399.600 ;
        RECT 673.950 397.950 676.050 398.400 ;
        RECT 700.950 397.950 703.050 398.400 ;
        RECT 712.950 399.600 715.050 400.050 ;
        RECT 734.400 399.600 735.600 401.400 ;
        RECT 742.950 400.950 745.050 401.400 ;
        RECT 712.950 398.400 735.600 399.600 ;
        RECT 754.950 399.600 757.050 400.050 ;
        RECT 778.950 399.600 781.050 400.050 ;
        RECT 754.950 398.400 781.050 399.600 ;
        RECT 712.950 397.950 715.050 398.400 ;
        RECT 754.950 397.950 757.050 398.400 ;
        RECT 778.950 397.950 781.050 398.400 ;
        RECT 187.950 396.600 190.050 397.050 ;
        RECT 205.950 396.600 208.050 397.050 ;
        RECT 187.950 395.400 208.050 396.600 ;
        RECT 187.950 394.950 190.050 395.400 ;
        RECT 205.950 394.950 208.050 395.400 ;
        RECT 223.950 396.600 226.050 397.050 ;
        RECT 256.950 396.600 259.050 397.050 ;
        RECT 382.950 396.600 385.050 397.050 ;
        RECT 223.950 395.400 385.050 396.600 ;
        RECT 223.950 394.950 226.050 395.400 ;
        RECT 256.950 394.950 259.050 395.400 ;
        RECT 382.950 394.950 385.050 395.400 ;
        RECT 601.950 396.600 604.050 397.050 ;
        RECT 646.950 396.600 649.050 397.050 ;
        RECT 601.950 395.400 649.050 396.600 ;
        RECT 601.950 394.950 604.050 395.400 ;
        RECT 646.950 394.950 649.050 395.400 ;
        RECT 736.950 396.600 739.050 397.050 ;
        RECT 829.950 396.600 832.050 397.050 ;
        RECT 736.950 395.400 832.050 396.600 ;
        RECT 736.950 394.950 739.050 395.400 ;
        RECT 829.950 394.950 832.050 395.400 ;
        RECT 28.950 393.600 31.050 394.050 ;
        RECT 82.950 393.600 85.050 394.050 ;
        RECT 28.950 392.400 85.050 393.600 ;
        RECT 28.950 391.950 31.050 392.400 ;
        RECT 82.950 391.950 85.050 392.400 ;
        RECT 142.950 393.600 145.050 394.050 ;
        RECT 160.950 393.600 163.050 394.050 ;
        RECT 238.950 393.600 241.050 394.050 ;
        RECT 142.950 392.400 241.050 393.600 ;
        RECT 142.950 391.950 145.050 392.400 ;
        RECT 160.950 391.950 163.050 392.400 ;
        RECT 238.950 391.950 241.050 392.400 ;
        RECT 268.950 393.600 271.050 394.050 ;
        RECT 322.950 393.600 325.050 394.050 ;
        RECT 268.950 392.400 325.050 393.600 ;
        RECT 268.950 391.950 271.050 392.400 ;
        RECT 322.950 391.950 325.050 392.400 ;
        RECT 346.950 393.600 349.050 394.050 ;
        RECT 367.950 393.600 370.050 394.050 ;
        RECT 397.950 393.600 400.050 394.050 ;
        RECT 346.950 392.400 400.050 393.600 ;
        RECT 346.950 391.950 349.050 392.400 ;
        RECT 367.950 391.950 370.050 392.400 ;
        RECT 397.950 391.950 400.050 392.400 ;
        RECT 169.950 390.600 172.050 391.050 ;
        RECT 187.950 390.600 190.050 391.050 ;
        RECT 169.950 389.400 190.050 390.600 ;
        RECT 169.950 388.950 172.050 389.400 ;
        RECT 187.950 388.950 190.050 389.400 ;
        RECT 199.950 390.600 202.050 391.050 ;
        RECT 223.950 390.600 226.050 391.050 ;
        RECT 199.950 389.400 226.050 390.600 ;
        RECT 199.950 388.950 202.050 389.400 ;
        RECT 223.950 388.950 226.050 389.400 ;
        RECT 319.950 390.600 322.050 391.050 ;
        RECT 406.950 390.600 409.050 391.050 ;
        RECT 838.950 390.600 841.050 391.050 ;
        RECT 319.950 389.400 409.050 390.600 ;
        RECT 319.950 388.950 322.050 389.400 ;
        RECT 406.950 388.950 409.050 389.400 ;
        RECT 815.400 389.400 841.050 390.600 ;
        RECT 112.950 387.600 115.050 388.050 ;
        RECT 145.950 387.600 148.050 388.050 ;
        RECT 112.950 386.400 148.050 387.600 ;
        RECT 112.950 385.950 115.050 386.400 ;
        RECT 145.950 385.950 148.050 386.400 ;
        RECT 175.950 387.600 178.050 388.050 ;
        RECT 484.950 387.600 487.050 388.050 ;
        RECT 175.950 386.400 487.050 387.600 ;
        RECT 175.950 385.950 178.050 386.400 ;
        RECT 484.950 385.950 487.050 386.400 ;
        RECT 541.950 387.600 544.050 388.050 ;
        RECT 640.950 387.600 643.050 388.050 ;
        RECT 664.950 387.600 667.050 388.050 ;
        RECT 670.950 387.600 673.050 388.050 ;
        RECT 541.950 386.400 673.050 387.600 ;
        RECT 541.950 385.950 544.050 386.400 ;
        RECT 640.950 385.950 643.050 386.400 ;
        RECT 664.950 385.950 667.050 386.400 ;
        RECT 670.950 385.950 673.050 386.400 ;
        RECT 685.950 387.600 688.050 388.050 ;
        RECT 815.400 387.600 816.600 389.400 ;
        RECT 838.950 388.950 841.050 389.400 ;
        RECT 685.950 386.400 816.600 387.600 ;
        RECT 685.950 385.950 688.050 386.400 ;
        RECT 4.950 384.600 7.050 385.050 ;
        RECT 25.950 384.600 28.050 385.050 ;
        RECT 4.950 383.400 28.050 384.600 ;
        RECT 4.950 382.950 7.050 383.400 ;
        RECT 25.950 382.950 28.050 383.400 ;
        RECT 661.950 384.600 664.050 385.050 ;
        RECT 682.950 384.600 685.050 385.050 ;
        RECT 823.950 384.600 826.050 385.050 ;
        RECT 661.950 383.400 685.050 384.600 ;
        RECT 812.400 384.000 826.050 384.600 ;
        RECT 661.950 382.950 664.050 383.400 ;
        RECT 682.950 382.950 685.050 383.400 ;
        RECT 811.950 383.400 826.050 384.000 ;
        RECT 235.950 381.600 238.050 382.050 ;
        RECT 253.950 381.600 256.050 382.050 ;
        RECT 235.950 380.400 256.050 381.600 ;
        RECT 235.950 379.950 238.050 380.400 ;
        RECT 253.950 379.950 256.050 380.400 ;
        RECT 274.950 381.600 277.050 382.050 ;
        RECT 286.950 381.600 289.050 382.050 ;
        RECT 274.950 380.400 289.050 381.600 ;
        RECT 274.950 379.950 277.050 380.400 ;
        RECT 286.950 379.950 289.050 380.400 ;
        RECT 610.950 381.600 613.050 382.050 ;
        RECT 616.950 381.600 619.050 382.050 ;
        RECT 610.950 380.400 619.050 381.600 ;
        RECT 610.950 379.950 613.050 380.400 ;
        RECT 616.950 379.950 619.050 380.400 ;
        RECT 766.950 381.600 769.050 382.050 ;
        RECT 787.950 381.600 790.050 382.050 ;
        RECT 766.950 380.400 790.050 381.600 ;
        RECT 766.950 379.950 769.050 380.400 ;
        RECT 787.950 379.950 790.050 380.400 ;
        RECT 811.950 379.950 814.050 383.400 ;
        RECT 823.950 382.950 826.050 383.400 ;
        RECT 40.950 378.600 43.050 379.050 ;
        RECT 61.950 378.600 64.050 379.050 ;
        RECT 40.950 377.400 64.050 378.600 ;
        RECT 40.950 376.950 43.050 377.400 ;
        RECT 61.950 376.950 64.050 377.400 ;
        RECT 97.950 378.600 100.050 379.050 ;
        RECT 112.950 378.600 115.050 379.050 ;
        RECT 133.950 378.600 136.050 379.050 ;
        RECT 97.950 377.400 136.050 378.600 ;
        RECT 97.950 376.950 100.050 377.400 ;
        RECT 112.950 376.950 115.050 377.400 ;
        RECT 133.950 376.950 136.050 377.400 ;
        RECT 169.950 378.600 172.050 379.050 ;
        RECT 178.950 378.600 181.050 379.050 ;
        RECT 169.950 377.400 181.050 378.600 ;
        RECT 169.950 376.950 172.050 377.400 ;
        RECT 178.950 376.950 181.050 377.400 ;
        RECT 193.950 378.600 196.050 379.050 ;
        RECT 217.950 378.600 220.050 379.050 ;
        RECT 193.950 377.400 220.050 378.600 ;
        RECT 193.950 376.950 196.050 377.400 ;
        RECT 217.950 376.950 220.050 377.400 ;
        RECT 232.950 378.600 235.050 379.050 ;
        RECT 271.950 378.600 274.050 379.050 ;
        RECT 232.950 377.400 274.050 378.600 ;
        RECT 232.950 376.950 235.050 377.400 ;
        RECT 271.950 376.950 274.050 377.400 ;
        RECT 328.950 378.600 331.050 379.050 ;
        RECT 343.950 378.600 346.050 379.050 ;
        RECT 376.950 378.600 379.050 379.050 ;
        RECT 328.950 377.400 379.050 378.600 ;
        RECT 328.950 376.950 331.050 377.400 ;
        RECT 343.950 376.950 346.050 377.400 ;
        RECT 376.950 376.950 379.050 377.400 ;
        RECT 508.950 378.600 511.050 379.050 ;
        RECT 529.950 378.600 532.050 379.050 ;
        RECT 508.950 377.400 532.050 378.600 ;
        RECT 508.950 376.950 511.050 377.400 ;
        RECT 529.950 376.950 532.050 377.400 ;
        RECT 598.950 378.600 601.050 379.050 ;
        RECT 625.950 378.600 628.050 379.050 ;
        RECT 598.950 377.400 628.050 378.600 ;
        RECT 598.950 376.950 601.050 377.400 ;
        RECT 625.950 376.950 628.050 377.400 ;
        RECT 643.950 378.600 646.050 379.050 ;
        RECT 655.950 378.600 658.050 379.050 ;
        RECT 643.950 377.400 658.050 378.600 ;
        RECT 643.950 376.950 646.050 377.400 ;
        RECT 655.950 376.950 658.050 377.400 ;
        RECT 664.950 378.600 667.050 379.050 ;
        RECT 703.950 378.600 706.050 379.050 ;
        RECT 814.950 378.600 817.050 379.050 ;
        RECT 832.950 378.600 835.050 379.050 ;
        RECT 853.950 378.600 856.050 379.050 ;
        RECT 664.950 377.400 774.600 378.600 ;
        RECT 664.950 376.950 667.050 377.400 ;
        RECT 703.950 376.950 706.050 377.400 ;
        RECT 773.400 376.050 774.600 377.400 ;
        RECT 814.950 377.400 856.050 378.600 ;
        RECT 814.950 376.950 817.050 377.400 ;
        RECT 832.950 376.950 835.050 377.400 ;
        RECT 853.950 376.950 856.050 377.400 ;
        RECT 136.950 375.600 139.050 376.050 ;
        RECT 166.950 375.600 169.050 376.050 ;
        RECT 136.950 374.400 169.050 375.600 ;
        RECT 136.950 373.950 139.050 374.400 ;
        RECT 166.950 373.950 169.050 374.400 ;
        RECT 220.950 375.600 223.050 376.050 ;
        RECT 241.950 375.600 244.050 376.050 ;
        RECT 220.950 374.400 244.050 375.600 ;
        RECT 220.950 373.950 223.050 374.400 ;
        RECT 241.950 373.950 244.050 374.400 ;
        RECT 280.950 375.600 283.050 376.050 ;
        RECT 298.950 375.600 301.050 376.050 ;
        RECT 340.950 375.600 343.050 376.050 ;
        RECT 370.950 375.600 373.050 376.050 ;
        RECT 400.950 375.600 403.050 376.050 ;
        RECT 496.950 375.600 499.050 376.050 ;
        RECT 280.950 374.400 403.050 375.600 ;
        RECT 280.950 373.950 283.050 374.400 ;
        RECT 298.950 373.950 301.050 374.400 ;
        RECT 340.950 373.950 343.050 374.400 ;
        RECT 370.950 373.950 373.050 374.400 ;
        RECT 400.950 373.950 403.050 374.400 ;
        RECT 470.400 374.400 499.050 375.600 ;
        RECT 12.000 372.600 16.050 373.050 ;
        RECT 11.400 370.950 16.050 372.600 ;
        RECT 19.950 372.600 22.050 373.050 ;
        RECT 28.950 372.600 31.050 373.050 ;
        RECT 19.950 371.400 31.050 372.600 ;
        RECT 19.950 370.950 22.050 371.400 ;
        RECT 28.950 370.950 31.050 371.400 ;
        RECT 43.800 370.950 45.900 373.050 ;
        RECT 46.950 371.100 49.050 373.200 ;
        RECT 55.950 372.600 58.050 373.200 ;
        RECT 64.950 372.600 67.050 373.050 ;
        RECT 55.950 371.400 67.050 372.600 ;
        RECT 55.950 371.100 58.050 371.400 ;
        RECT 11.400 367.050 12.600 370.950 ;
        RECT 44.400 367.050 45.600 370.950 ;
        RECT 47.400 369.600 48.600 371.100 ;
        RECT 64.950 370.950 67.050 371.400 ;
        RECT 91.950 372.600 94.050 373.050 ;
        RECT 118.950 372.600 121.050 373.050 ;
        RECT 133.950 372.600 136.050 373.200 ;
        RECT 174.000 372.600 178.050 373.050 ;
        RECT 91.950 371.400 136.050 372.600 ;
        RECT 91.950 370.950 94.050 371.400 ;
        RECT 118.950 370.950 121.050 371.400 ;
        RECT 133.950 371.100 136.050 371.400 ;
        RECT 173.400 370.950 178.050 372.600 ;
        RECT 181.950 372.600 184.050 373.050 ;
        RECT 181.950 371.400 192.600 372.600 ;
        RECT 181.950 370.950 184.050 371.400 ;
        RECT 47.400 368.400 51.600 369.600 ;
        RECT 7.950 365.400 12.600 367.050 ;
        RECT 16.950 366.600 19.050 366.750 ;
        RECT 31.950 366.600 34.050 366.750 ;
        RECT 16.950 365.400 34.050 366.600 ;
        RECT 7.950 364.950 12.000 365.400 ;
        RECT 16.950 364.650 19.050 365.400 ;
        RECT 31.950 364.650 34.050 365.400 ;
        RECT 43.950 364.950 46.050 367.050 ;
        RECT 50.400 366.600 51.600 368.400 ;
        RECT 173.400 367.050 174.600 370.950 ;
        RECT 50.400 365.400 54.600 366.600 ;
        RECT 53.400 364.050 54.600 365.400 ;
        RECT 94.950 366.300 97.050 366.750 ;
        RECT 103.950 366.600 106.050 366.750 ;
        RECT 115.950 366.600 118.050 366.750 ;
        RECT 103.950 366.300 118.050 366.600 ;
        RECT 94.950 365.400 118.050 366.300 ;
        RECT 94.950 365.100 106.050 365.400 ;
        RECT 94.950 364.650 97.050 365.100 ;
        RECT 103.950 364.650 106.050 365.100 ;
        RECT 115.950 364.650 118.050 365.400 ;
        RECT 136.950 366.450 139.050 366.900 ;
        RECT 157.950 366.450 160.050 366.900 ;
        RECT 136.950 365.250 160.050 366.450 ;
        RECT 136.950 364.800 139.050 365.250 ;
        RECT 157.950 364.800 160.050 365.250 ;
        RECT 172.950 364.950 175.050 367.050 ;
        RECT 184.950 366.600 187.050 367.050 ;
        RECT 191.400 366.900 192.600 371.400 ;
        RECT 202.950 371.100 205.050 373.200 ;
        RECT 211.950 372.750 214.050 373.200 ;
        RECT 232.950 372.750 235.050 373.200 ;
        RECT 211.950 371.550 235.050 372.750 ;
        RECT 211.950 371.100 214.050 371.550 ;
        RECT 232.950 371.100 235.050 371.550 ;
        RECT 250.950 372.600 253.050 373.050 ;
        RECT 256.950 372.600 259.050 373.050 ;
        RECT 250.950 371.400 259.050 372.600 ;
        RECT 203.400 367.050 204.600 371.100 ;
        RECT 250.950 370.950 253.050 371.400 ;
        RECT 256.950 370.950 259.050 371.400 ;
        RECT 265.950 372.600 268.050 373.200 ;
        RECT 291.000 372.600 295.050 373.050 ;
        RECT 307.950 372.600 310.050 373.200 ;
        RECT 265.950 371.400 276.600 372.600 ;
        RECT 265.950 371.100 268.050 371.400 ;
        RECT 275.400 367.050 276.600 371.400 ;
        RECT 290.400 370.950 295.050 372.600 ;
        RECT 302.400 371.400 310.050 372.600 ;
        RECT 190.950 366.600 193.050 366.900 ;
        RECT 184.950 365.400 193.050 366.600 ;
        RECT 184.950 364.950 187.050 365.400 ;
        RECT 190.950 364.800 193.050 365.400 ;
        RECT 199.950 365.400 204.600 367.050 ;
        RECT 229.950 366.450 232.050 366.900 ;
        RECT 244.950 366.600 247.050 366.900 ;
        RECT 253.800 366.600 255.900 367.050 ;
        RECT 244.950 366.450 255.900 366.600 ;
        RECT 229.950 365.400 255.900 366.450 ;
        RECT 199.950 364.950 204.000 365.400 ;
        RECT 229.950 365.250 247.050 365.400 ;
        RECT 229.950 364.800 232.050 365.250 ;
        RECT 244.950 364.800 247.050 365.250 ;
        RECT 253.800 364.950 255.900 365.400 ;
        RECT 256.950 366.450 259.050 366.900 ;
        RECT 262.950 366.450 265.050 366.900 ;
        RECT 256.950 365.250 265.050 366.450 ;
        RECT 256.950 364.800 259.050 365.250 ;
        RECT 262.950 364.800 265.050 365.250 ;
        RECT 274.950 364.950 277.050 367.050 ;
        RECT 290.400 366.750 291.600 370.950 ;
        RECT 295.950 369.600 298.050 370.050 ;
        RECT 302.400 369.600 303.600 371.400 ;
        RECT 307.950 371.100 310.050 371.400 ;
        RECT 322.950 372.750 325.050 373.200 ;
        RECT 334.800 372.750 336.900 373.200 ;
        RECT 322.950 371.550 336.900 372.750 ;
        RECT 322.950 371.100 325.050 371.550 ;
        RECT 334.800 371.100 336.900 371.550 ;
        RECT 337.950 372.750 340.050 373.200 ;
        RECT 349.950 372.750 352.050 373.200 ;
        RECT 337.950 372.600 352.050 372.750 ;
        RECT 364.950 372.600 367.050 373.200 ;
        RECT 385.950 372.600 388.050 373.200 ;
        RECT 337.950 371.550 367.050 372.600 ;
        RECT 337.950 371.100 340.050 371.550 ;
        RECT 349.950 371.400 367.050 371.550 ;
        RECT 349.950 371.100 352.050 371.400 ;
        RECT 364.950 371.100 367.050 371.400 ;
        RECT 368.400 371.400 388.050 372.600 ;
        RECT 368.400 369.600 369.600 371.400 ;
        RECT 385.950 371.100 388.050 371.400 ;
        RECT 412.950 372.600 415.050 373.050 ;
        RECT 418.950 372.600 421.050 373.050 ;
        RECT 448.950 372.600 451.050 373.200 ;
        RECT 470.400 373.050 471.600 374.400 ;
        RECT 496.950 373.950 499.050 374.400 ;
        RECT 505.950 375.600 510.000 376.050 ;
        RECT 607.950 375.600 610.050 376.050 ;
        RECT 619.950 375.600 622.050 376.050 ;
        RECT 505.950 373.950 510.600 375.600 ;
        RECT 607.950 374.400 622.050 375.600 ;
        RECT 607.950 373.950 610.050 374.400 ;
        RECT 619.950 373.950 622.050 374.400 ;
        RECT 649.950 375.600 652.050 376.050 ;
        RECT 773.400 375.600 778.050 376.050 ;
        RECT 649.950 374.400 666.600 375.600 ;
        RECT 773.400 375.000 810.600 375.600 ;
        RECT 773.400 374.400 811.050 375.000 ;
        RECT 649.950 373.950 652.050 374.400 ;
        RECT 412.950 371.400 421.050 372.600 ;
        RECT 412.950 370.950 415.050 371.400 ;
        RECT 418.950 370.950 421.050 371.400 ;
        RECT 437.400 371.400 451.050 372.600 ;
        RECT 295.950 368.400 303.600 369.600 ;
        RECT 362.400 368.400 369.600 369.600 ;
        RECT 295.950 367.950 298.050 368.400 ;
        RECT 289.950 364.650 292.050 366.750 ;
        RECT 310.950 366.600 313.050 366.900 ;
        RECT 334.950 366.600 337.050 367.050 ;
        RECT 362.400 366.900 363.600 368.400 ;
        RECT 437.400 367.050 438.600 371.400 ;
        RECT 448.950 371.100 451.050 371.400 ;
        RECT 454.950 370.950 457.050 373.050 ;
        RECT 463.950 372.600 466.050 373.050 ;
        RECT 469.800 372.600 471.900 373.050 ;
        RECT 463.950 371.400 471.900 372.600 ;
        RECT 463.950 370.950 466.050 371.400 ;
        RECT 469.800 370.950 471.900 371.400 ;
        RECT 472.950 372.750 475.050 373.200 ;
        RECT 478.950 372.750 481.050 373.200 ;
        RECT 472.950 371.550 481.050 372.750 ;
        RECT 493.950 372.600 496.050 373.050 ;
        RECT 472.950 371.100 475.050 371.550 ;
        RECT 478.950 371.100 481.050 371.550 ;
        RECT 482.400 371.400 496.050 372.600 ;
        RECT 455.400 367.050 456.600 370.950 ;
        RECT 352.950 366.600 355.050 366.900 ;
        RECT 361.950 366.600 364.050 366.900 ;
        RECT 310.950 365.400 364.050 366.600 ;
        RECT 310.950 364.800 313.050 365.400 ;
        RECT 334.950 364.950 337.050 365.400 ;
        RECT 352.950 364.800 355.050 365.400 ;
        RECT 361.950 364.800 364.050 365.400 ;
        RECT 376.950 366.600 379.050 367.050 ;
        RECT 421.950 366.600 424.050 366.750 ;
        RECT 376.950 365.400 424.050 366.600 ;
        RECT 376.950 364.950 379.050 365.400 ;
        RECT 421.950 364.650 424.050 365.400 ;
        RECT 436.950 364.950 439.050 367.050 ;
        RECT 454.950 364.950 457.050 367.050 ;
        RECT 482.400 366.900 483.600 371.400 ;
        RECT 493.950 370.950 496.050 371.400 ;
        RECT 502.950 370.950 505.050 373.050 ;
        RECT 481.950 364.800 484.050 366.900 ;
        RECT 487.950 366.600 490.050 366.900 ;
        RECT 503.400 366.600 504.600 370.950 ;
        RECT 509.400 369.600 510.600 373.950 ;
        RECT 541.950 372.750 544.050 373.200 ;
        RECT 547.950 372.750 550.050 373.200 ;
        RECT 541.950 371.550 550.050 372.750 ;
        RECT 541.950 371.100 544.050 371.550 ;
        RECT 547.950 371.100 550.050 371.550 ;
        RECT 556.950 372.750 559.050 373.200 ;
        RECT 562.950 372.750 565.050 373.200 ;
        RECT 556.950 371.550 565.050 372.750 ;
        RECT 556.950 371.100 559.050 371.550 ;
        RECT 562.950 371.100 565.050 371.550 ;
        RECT 589.950 372.600 592.050 373.200 ;
        RECT 595.950 372.600 598.050 373.050 ;
        RECT 589.950 371.400 598.050 372.600 ;
        RECT 589.950 371.100 592.050 371.400 ;
        RECT 595.950 370.950 598.050 371.400 ;
        RECT 604.950 372.600 607.050 373.050 ;
        RECT 634.950 372.600 637.050 373.050 ;
        RECT 604.950 371.400 633.600 372.600 ;
        RECT 604.950 370.950 607.050 371.400 ;
        RECT 509.400 368.400 513.600 369.600 ;
        RECT 512.400 366.900 513.600 368.400 ;
        RECT 487.950 365.400 504.600 366.600 ;
        RECT 487.950 364.800 490.050 365.400 ;
        RECT 511.950 364.800 514.050 366.900 ;
        RECT 574.950 366.600 577.050 366.900 ;
        RECT 586.950 366.600 589.050 366.900 ;
        RECT 632.400 366.750 633.600 371.400 ;
        RECT 634.950 371.400 654.600 372.600 ;
        RECT 634.950 370.950 637.050 371.400 ;
        RECT 653.400 366.750 654.600 371.400 ;
        RECT 665.400 367.050 666.600 374.400 ;
        RECT 774.000 373.950 778.050 374.400 ;
        RECT 676.950 371.100 679.050 373.200 ;
        RECT 712.950 372.750 715.050 373.200 ;
        RECT 721.950 372.750 724.050 373.200 ;
        RECT 712.950 371.550 724.050 372.750 ;
        RECT 712.950 371.100 715.050 371.550 ;
        RECT 721.950 371.100 724.050 371.550 ;
        RECT 739.950 372.600 742.050 373.050 ;
        RECT 745.950 372.600 748.050 373.200 ;
        RECT 739.950 371.400 748.050 372.600 ;
        RECT 677.400 369.600 678.600 371.100 ;
        RECT 739.950 370.950 742.050 371.400 ;
        RECT 745.950 371.100 748.050 371.400 ;
        RECT 784.950 372.750 787.050 373.200 ;
        RECT 790.950 372.750 793.050 373.200 ;
        RECT 784.950 371.550 793.050 372.750 ;
        RECT 784.950 371.100 787.050 371.550 ;
        RECT 790.950 371.100 793.050 371.550 ;
        RECT 808.950 370.950 811.050 374.400 ;
        RECT 814.950 369.600 817.050 373.050 ;
        RECT 826.950 372.600 829.050 373.050 ;
        RECT 677.400 368.400 705.600 369.600 ;
        RECT 574.950 365.400 589.050 366.600 ;
        RECT 574.950 364.800 577.050 365.400 ;
        RECT 586.950 364.800 589.050 365.400 ;
        RECT 595.950 366.300 598.050 366.750 ;
        RECT 601.950 366.300 604.050 366.750 ;
        RECT 595.950 365.100 604.050 366.300 ;
        RECT 595.950 364.650 598.050 365.100 ;
        RECT 601.950 364.650 604.050 365.100 ;
        RECT 613.950 366.300 616.050 366.750 ;
        RECT 619.950 366.300 622.050 366.750 ;
        RECT 613.950 365.100 622.050 366.300 ;
        RECT 613.950 364.650 616.050 365.100 ;
        RECT 619.950 364.650 622.050 365.100 ;
        RECT 631.950 364.650 634.050 366.750 ;
        RECT 652.950 364.650 655.050 366.750 ;
        RECT 664.950 364.950 667.050 367.050 ;
        RECT 704.400 366.600 705.600 368.400 ;
        RECT 803.400 369.000 817.050 369.600 ;
        RECT 818.400 371.400 829.050 372.600 ;
        RECT 803.400 368.400 816.600 369.000 ;
        RECT 709.950 366.600 712.050 367.050 ;
        RECT 803.400 366.900 804.600 368.400 ;
        RECT 818.400 367.050 819.600 371.400 ;
        RECT 826.950 370.950 829.050 371.400 ;
        RECT 838.950 372.600 841.050 373.050 ;
        RECT 856.950 372.600 859.050 373.050 ;
        RECT 862.950 372.600 865.050 373.050 ;
        RECT 838.950 371.400 865.050 372.600 ;
        RECT 838.950 370.950 841.050 371.400 ;
        RECT 856.950 370.950 859.050 371.400 ;
        RECT 862.950 370.950 865.050 371.400 ;
        RECT 704.400 365.400 712.050 366.600 ;
        RECT 709.950 364.950 712.050 365.400 ;
        RECT 739.950 366.450 742.050 366.900 ;
        RECT 757.950 366.450 760.050 366.900 ;
        RECT 739.950 365.250 760.050 366.450 ;
        RECT 739.950 364.800 742.050 365.250 ;
        RECT 757.950 364.800 760.050 365.250 ;
        RECT 802.950 364.800 805.050 366.900 ;
        RECT 814.950 365.400 819.600 367.050 ;
        RECT 814.950 364.950 819.000 365.400 ;
        RECT 53.400 362.400 58.050 364.050 ;
        RECT 82.950 363.600 85.050 364.050 ;
        RECT 54.000 361.950 58.050 362.400 ;
        RECT 62.400 362.400 85.050 363.600 ;
        RECT 10.950 360.600 13.050 361.050 ;
        RECT 62.400 360.600 63.600 362.400 ;
        RECT 82.950 361.950 85.050 362.400 ;
        RECT 130.950 363.600 133.050 364.050 ;
        RECT 142.950 363.600 145.050 364.050 ;
        RECT 130.950 362.400 145.050 363.600 ;
        RECT 130.950 361.950 133.050 362.400 ;
        RECT 142.950 361.950 145.050 362.400 ;
        RECT 271.950 363.600 274.050 364.050 ;
        RECT 283.950 363.600 286.050 364.050 ;
        RECT 271.950 362.400 286.050 363.600 ;
        RECT 271.950 361.950 274.050 362.400 ;
        RECT 283.950 361.950 286.050 362.400 ;
        RECT 382.950 363.600 385.050 364.050 ;
        RECT 412.950 363.600 415.050 364.050 ;
        RECT 382.950 362.400 415.050 363.600 ;
        RECT 382.950 361.950 385.050 362.400 ;
        RECT 412.950 361.950 415.050 362.400 ;
        RECT 445.950 363.600 448.050 364.050 ;
        RECT 469.950 363.600 472.050 364.050 ;
        RECT 445.950 362.400 472.050 363.600 ;
        RECT 445.950 361.950 448.050 362.400 ;
        RECT 469.950 361.950 472.050 362.400 ;
        RECT 730.950 363.600 733.050 364.050 ;
        RECT 748.950 363.600 751.050 364.050 ;
        RECT 730.950 362.400 751.050 363.600 ;
        RECT 730.950 361.950 733.050 362.400 ;
        RECT 748.950 361.950 751.050 362.400 ;
        RECT 811.950 363.600 814.050 364.050 ;
        RECT 835.950 363.600 838.050 364.050 ;
        RECT 811.950 362.400 838.050 363.600 ;
        RECT 811.950 361.950 814.050 362.400 ;
        RECT 835.950 361.950 838.050 362.400 ;
        RECT 10.950 359.400 63.600 360.600 ;
        RECT 145.950 360.600 148.050 361.050 ;
        RECT 154.950 360.600 157.050 360.900 ;
        RECT 145.950 359.400 157.050 360.600 ;
        RECT 10.950 358.950 13.050 359.400 ;
        RECT 145.950 358.950 148.050 359.400 ;
        RECT 154.950 358.800 157.050 359.400 ;
        RECT 178.950 360.600 181.050 361.050 ;
        RECT 247.950 360.600 250.050 361.050 ;
        RECT 268.950 360.600 271.050 361.050 ;
        RECT 178.950 359.400 271.050 360.600 ;
        RECT 178.950 358.950 181.050 359.400 ;
        RECT 247.950 358.950 250.050 359.400 ;
        RECT 268.950 358.950 271.050 359.400 ;
        RECT 274.950 360.600 277.050 361.050 ;
        RECT 280.950 360.600 283.050 361.050 ;
        RECT 304.950 360.600 307.050 361.050 ;
        RECT 274.950 359.400 307.050 360.600 ;
        RECT 274.950 358.950 277.050 359.400 ;
        RECT 280.950 358.950 283.050 359.400 ;
        RECT 304.950 358.950 307.050 359.400 ;
        RECT 361.950 360.600 364.050 361.050 ;
        RECT 383.400 360.600 384.600 361.950 ;
        RECT 361.950 359.400 384.600 360.600 ;
        RECT 562.950 360.600 565.050 361.050 ;
        RECT 607.950 360.600 610.050 361.050 ;
        RECT 562.950 359.400 610.050 360.600 ;
        RECT 361.950 358.950 364.050 359.400 ;
        RECT 562.950 358.950 565.050 359.400 ;
        RECT 607.950 358.950 610.050 359.400 ;
        RECT 658.950 360.600 661.050 361.050 ;
        RECT 685.950 360.600 688.050 361.050 ;
        RECT 658.950 359.400 688.050 360.600 ;
        RECT 658.950 358.950 661.050 359.400 ;
        RECT 685.950 358.950 688.050 359.400 ;
        RECT 721.950 360.600 724.050 361.050 ;
        RECT 763.950 360.600 766.050 361.050 ;
        RECT 721.950 359.400 766.050 360.600 ;
        RECT 721.950 358.950 724.050 359.400 ;
        RECT 763.950 358.950 766.050 359.400 ;
        RECT 91.950 357.600 94.050 358.050 ;
        RECT 109.950 357.600 112.050 358.050 ;
        RECT 91.950 356.400 112.050 357.600 ;
        RECT 91.950 355.950 94.050 356.400 ;
        RECT 109.950 355.950 112.050 356.400 ;
        RECT 124.950 357.600 127.050 358.050 ;
        RECT 142.950 357.600 145.050 358.050 ;
        RECT 124.950 356.400 145.050 357.600 ;
        RECT 124.950 355.950 127.050 356.400 ;
        RECT 142.950 355.950 145.050 356.400 ;
        RECT 211.950 357.600 214.050 358.050 ;
        RECT 217.950 357.600 220.050 358.050 ;
        RECT 211.950 356.400 220.050 357.600 ;
        RECT 211.950 355.950 214.050 356.400 ;
        RECT 217.950 355.950 220.050 356.400 ;
        RECT 421.950 357.600 424.050 358.050 ;
        RECT 460.950 357.600 463.050 358.050 ;
        RECT 421.950 356.400 463.050 357.600 ;
        RECT 421.950 355.950 424.050 356.400 ;
        RECT 460.950 355.950 463.050 356.400 ;
        RECT 472.950 357.600 475.050 358.050 ;
        RECT 499.950 357.600 502.050 358.050 ;
        RECT 472.950 356.400 502.050 357.600 ;
        RECT 472.950 355.950 475.050 356.400 ;
        RECT 499.950 355.950 502.050 356.400 ;
        RECT 4.950 354.600 7.050 355.050 ;
        RECT 16.950 354.600 19.050 355.050 ;
        RECT 4.950 353.400 19.050 354.600 ;
        RECT 4.950 352.950 7.050 353.400 ;
        RECT 16.950 352.950 19.050 353.400 ;
        RECT 31.950 354.600 34.050 355.050 ;
        RECT 61.950 354.600 64.050 355.050 ;
        RECT 31.950 353.400 64.050 354.600 ;
        RECT 31.950 352.950 34.050 353.400 ;
        RECT 61.950 352.950 64.050 353.400 ;
        RECT 76.950 354.600 79.050 355.050 ;
        RECT 199.950 354.600 202.050 355.050 ;
        RECT 208.950 354.600 211.050 355.050 ;
        RECT 76.950 353.400 150.600 354.600 ;
        RECT 76.950 352.950 79.050 353.400 ;
        RECT 149.400 352.050 150.600 353.400 ;
        RECT 199.950 353.400 211.050 354.600 ;
        RECT 199.950 352.950 202.050 353.400 ;
        RECT 208.950 352.950 211.050 353.400 ;
        RECT 301.950 354.600 304.050 355.050 ;
        RECT 325.950 354.600 328.050 355.050 ;
        RECT 301.950 353.400 328.050 354.600 ;
        RECT 301.950 352.950 304.050 353.400 ;
        RECT 325.950 352.950 328.050 353.400 ;
        RECT 382.950 354.600 385.050 355.050 ;
        RECT 394.950 354.600 397.050 355.050 ;
        RECT 382.950 353.400 397.050 354.600 ;
        RECT 382.950 352.950 385.050 353.400 ;
        RECT 394.950 352.950 397.050 353.400 ;
        RECT 148.950 351.600 151.050 352.050 ;
        RECT 172.950 351.600 175.050 352.050 ;
        RECT 148.950 350.400 175.050 351.600 ;
        RECT 148.950 349.950 151.050 350.400 ;
        RECT 172.950 349.950 175.050 350.400 ;
        RECT 253.950 351.600 256.050 352.050 ;
        RECT 271.950 351.600 274.050 352.050 ;
        RECT 253.950 350.400 274.050 351.600 ;
        RECT 253.950 349.950 256.050 350.400 ;
        RECT 271.950 349.950 274.050 350.400 ;
        RECT 298.950 351.600 301.050 352.050 ;
        RECT 313.950 351.600 316.050 352.050 ;
        RECT 298.950 350.400 316.050 351.600 ;
        RECT 298.950 349.950 301.050 350.400 ;
        RECT 313.950 349.950 316.050 350.400 ;
        RECT 349.950 351.600 352.050 352.050 ;
        RECT 376.950 351.600 379.050 352.050 ;
        RECT 349.950 350.400 379.050 351.600 ;
        RECT 349.950 349.950 352.050 350.400 ;
        RECT 376.950 349.950 379.050 350.400 ;
        RECT 406.950 351.600 409.050 352.050 ;
        RECT 430.950 351.600 433.050 352.050 ;
        RECT 406.950 350.400 433.050 351.600 ;
        RECT 406.950 349.950 409.050 350.400 ;
        RECT 430.950 349.950 433.050 350.400 ;
        RECT 487.950 351.600 490.050 352.050 ;
        RECT 499.950 351.600 502.050 352.050 ;
        RECT 487.950 350.400 502.050 351.600 ;
        RECT 487.950 349.950 490.050 350.400 ;
        RECT 499.950 349.950 502.050 350.400 ;
        RECT 625.950 351.600 628.050 352.050 ;
        RECT 640.950 351.600 643.050 352.050 ;
        RECT 625.950 350.400 643.050 351.600 ;
        RECT 625.950 349.950 628.050 350.400 ;
        RECT 640.950 349.950 643.050 350.400 ;
        RECT 790.950 351.600 793.050 352.050 ;
        RECT 820.950 351.600 823.050 352.050 ;
        RECT 790.950 350.400 823.050 351.600 ;
        RECT 790.950 349.950 793.050 350.400 ;
        RECT 820.950 349.950 823.050 350.400 ;
        RECT 37.950 348.600 40.050 349.050 ;
        RECT 76.950 348.600 79.050 349.050 ;
        RECT 88.950 348.600 91.050 349.050 ;
        RECT 37.950 347.400 72.600 348.600 ;
        RECT 37.950 346.950 40.050 347.400 ;
        RECT 19.950 345.600 22.050 346.050 ;
        RECT 43.950 345.600 46.050 346.050 ;
        RECT 19.950 344.400 46.050 345.600 ;
        RECT 71.400 345.600 72.600 347.400 ;
        RECT 76.950 347.400 91.050 348.600 ;
        RECT 76.950 346.950 79.050 347.400 ;
        RECT 88.950 346.950 91.050 347.400 ;
        RECT 100.950 348.600 103.050 349.050 ;
        RECT 145.950 348.600 148.050 349.050 ;
        RECT 100.950 347.400 148.050 348.600 ;
        RECT 100.950 346.950 103.050 347.400 ;
        RECT 145.950 346.950 148.050 347.400 ;
        RECT 151.950 348.600 154.050 349.050 ;
        RECT 196.950 348.600 199.050 349.050 ;
        RECT 151.950 347.400 199.050 348.600 ;
        RECT 151.950 346.950 154.050 347.400 ;
        RECT 196.950 346.950 199.050 347.400 ;
        RECT 202.950 348.600 205.050 349.050 ;
        RECT 235.950 348.600 238.050 349.050 ;
        RECT 202.950 347.400 238.050 348.600 ;
        RECT 202.950 346.950 205.050 347.400 ;
        RECT 235.950 346.950 238.050 347.400 ;
        RECT 268.950 348.600 271.050 349.050 ;
        RECT 319.950 348.600 322.050 349.050 ;
        RECT 565.950 348.600 568.050 349.050 ;
        RECT 268.950 347.400 322.050 348.600 ;
        RECT 268.950 346.950 271.050 347.400 ;
        RECT 319.950 346.950 322.050 347.400 ;
        RECT 503.400 347.400 568.050 348.600 ;
        RECT 103.950 345.600 106.050 346.050 ;
        RECT 71.400 344.400 106.050 345.600 ;
        RECT 19.950 343.950 22.050 344.400 ;
        RECT 43.950 343.950 46.050 344.400 ;
        RECT 103.950 343.950 106.050 344.400 ;
        RECT 127.950 345.600 130.050 346.050 ;
        RECT 139.950 345.600 142.050 346.050 ;
        RECT 127.950 344.400 142.050 345.600 ;
        RECT 127.950 343.950 130.050 344.400 ;
        RECT 139.950 343.950 142.050 344.400 ;
        RECT 187.950 345.600 190.050 346.050 ;
        RECT 199.950 345.600 202.050 346.050 ;
        RECT 187.950 344.400 202.050 345.600 ;
        RECT 187.950 343.950 190.050 344.400 ;
        RECT 199.950 343.950 202.050 344.400 ;
        RECT 250.950 345.600 253.050 346.050 ;
        RECT 256.950 345.600 259.050 346.050 ;
        RECT 334.950 345.600 337.050 346.050 ;
        RECT 355.950 345.600 358.050 346.050 ;
        RECT 250.950 344.400 259.050 345.600 ;
        RECT 250.950 343.950 253.050 344.400 ;
        RECT 256.950 343.950 259.050 344.400 ;
        RECT 284.400 344.400 358.050 345.600 ;
        RECT 64.950 342.600 67.050 343.050 ;
        RECT 109.950 342.600 112.050 343.050 ;
        RECT 64.950 341.400 112.050 342.600 ;
        RECT 64.950 340.950 67.050 341.400 ;
        RECT 109.950 340.950 112.050 341.400 ;
        RECT 142.950 342.600 145.050 343.050 ;
        RECT 151.950 342.600 154.050 343.050 ;
        RECT 142.950 341.400 154.050 342.600 ;
        RECT 142.950 340.950 145.050 341.400 ;
        RECT 151.950 340.950 154.050 341.400 ;
        RECT 238.950 342.600 241.050 343.050 ;
        RECT 284.400 342.600 285.600 344.400 ;
        RECT 334.950 343.950 337.050 344.400 ;
        RECT 355.950 343.950 358.050 344.400 ;
        RECT 367.950 345.600 370.050 346.050 ;
        RECT 385.950 345.600 388.050 346.050 ;
        RECT 367.950 344.400 388.050 345.600 ;
        RECT 367.950 343.950 370.050 344.400 ;
        RECT 385.950 343.950 388.050 344.400 ;
        RECT 415.950 345.600 418.050 346.050 ;
        RECT 427.950 345.600 430.050 346.050 ;
        RECT 415.950 344.400 430.050 345.600 ;
        RECT 415.950 343.950 418.050 344.400 ;
        RECT 427.950 343.950 430.050 344.400 ;
        RECT 490.950 345.600 493.050 346.050 ;
        RECT 503.400 345.600 504.600 347.400 ;
        RECT 565.950 346.950 568.050 347.400 ;
        RECT 748.950 348.600 751.050 349.050 ;
        RECT 766.950 348.600 769.050 349.050 ;
        RECT 748.950 347.400 769.050 348.600 ;
        RECT 748.950 346.950 751.050 347.400 ;
        RECT 766.950 346.950 769.050 347.400 ;
        RECT 829.950 348.600 832.050 349.050 ;
        RECT 850.950 348.600 853.050 349.050 ;
        RECT 829.950 347.400 853.050 348.600 ;
        RECT 829.950 346.950 832.050 347.400 ;
        RECT 850.950 346.950 853.050 347.400 ;
        RECT 490.950 344.400 504.600 345.600 ;
        RECT 754.950 345.600 757.050 346.050 ;
        RECT 784.950 345.600 787.050 346.050 ;
        RECT 754.950 344.400 787.050 345.600 ;
        RECT 490.950 343.950 493.050 344.400 ;
        RECT 754.950 343.950 757.050 344.400 ;
        RECT 784.950 343.950 787.050 344.400 ;
        RECT 826.950 345.600 829.050 346.050 ;
        RECT 835.950 345.600 838.050 346.050 ;
        RECT 826.950 344.400 838.050 345.600 ;
        RECT 826.950 343.950 829.050 344.400 ;
        RECT 835.950 343.950 838.050 344.400 ;
        RECT 238.950 341.400 285.600 342.600 ;
        RECT 337.950 342.600 342.000 343.050 ;
        RECT 436.950 342.600 439.050 343.050 ;
        RECT 442.950 342.600 445.050 343.050 ;
        RECT 238.950 340.950 241.050 341.400 ;
        RECT 337.950 340.950 342.600 342.600 ;
        RECT 436.950 341.400 445.050 342.600 ;
        RECT 436.950 340.950 439.050 341.400 ;
        RECT 442.950 340.950 445.050 341.400 ;
        RECT 13.950 339.600 16.050 340.200 ;
        RECT 25.950 339.600 28.050 340.350 ;
        RECT 13.950 338.400 28.050 339.600 ;
        RECT 13.950 338.100 16.050 338.400 ;
        RECT 17.250 334.050 18.450 338.400 ;
        RECT 25.950 338.250 28.050 338.400 ;
        RECT 31.950 339.600 34.050 340.350 ;
        RECT 31.950 338.400 42.600 339.600 ;
        RECT 31.950 338.250 34.050 338.400 ;
        RECT 41.400 334.050 42.600 338.400 ;
        RECT 52.950 338.250 55.050 340.350 ;
        RECT 61.950 339.600 64.050 340.050 ;
        RECT 70.950 339.600 73.050 340.200 ;
        RECT 61.950 338.400 73.050 339.600 ;
        RECT 53.400 334.050 54.600 338.250 ;
        RECT 61.950 337.950 64.050 338.400 ;
        RECT 70.950 338.100 73.050 338.400 ;
        RECT 100.950 337.950 103.050 340.050 ;
        RECT 115.950 339.900 118.050 340.350 ;
        RECT 136.950 339.900 139.050 340.350 ;
        RECT 115.950 338.700 139.050 339.900 ;
        RECT 115.950 338.250 118.050 338.700 ;
        RECT 136.950 338.250 139.050 338.700 ;
        RECT 172.950 339.750 175.050 340.200 ;
        RECT 193.950 339.750 196.050 340.200 ;
        RECT 172.950 338.550 196.050 339.750 ;
        RECT 172.950 338.100 175.050 338.550 ;
        RECT 193.950 338.100 196.050 338.550 ;
        RECT 211.950 339.750 214.050 340.200 ;
        RECT 232.950 339.750 235.050 340.200 ;
        RECT 211.950 338.550 235.050 339.750 ;
        RECT 211.950 338.100 214.050 338.550 ;
        RECT 232.950 338.100 235.050 338.550 ;
        RECT 250.950 339.600 255.000 340.050 ;
        RECT 256.950 339.600 259.050 340.350 ;
        RECT 265.950 339.600 268.050 340.050 ;
        RECT 250.950 337.950 255.600 339.600 ;
        RECT 256.950 338.400 268.050 339.600 ;
        RECT 256.950 338.250 259.050 338.400 ;
        RECT 265.950 337.950 268.050 338.400 ;
        RECT 286.950 338.100 289.050 340.200 ;
        RECT 298.950 339.600 301.050 340.050 ;
        RECT 307.950 339.600 310.050 340.350 ;
        RECT 298.950 338.400 310.050 339.600 ;
        RECT 101.400 334.050 102.600 337.950 ;
        RECT 254.400 334.050 255.600 337.950 ;
        RECT 4.950 333.600 7.050 334.050 ;
        RECT 10.950 333.600 13.050 333.900 ;
        RECT 4.950 332.400 13.050 333.600 ;
        RECT 4.950 331.950 7.050 332.400 ;
        RECT 10.950 331.800 13.050 332.400 ;
        RECT 16.800 331.950 18.900 334.050 ;
        RECT 19.950 333.600 22.050 334.050 ;
        RECT 28.950 333.600 31.050 334.050 ;
        RECT 19.950 332.400 31.050 333.600 ;
        RECT 19.950 331.950 22.050 332.400 ;
        RECT 28.950 331.950 31.050 332.400 ;
        RECT 40.950 331.950 43.050 334.050 ;
        RECT 52.950 331.950 55.050 334.050 ;
        RECT 73.950 333.600 76.050 333.900 ;
        RECT 88.950 333.600 91.050 333.900 ;
        RECT 56.400 332.400 91.050 333.600 ;
        RECT 49.950 330.600 52.050 331.050 ;
        RECT 56.400 330.600 57.600 332.400 ;
        RECT 73.950 331.800 76.050 332.400 ;
        RECT 88.950 331.800 91.050 332.400 ;
        RECT 100.950 331.950 103.050 334.050 ;
        RECT 115.950 333.600 118.050 334.050 ;
        RECT 124.950 333.600 127.050 334.050 ;
        RECT 115.950 332.400 127.050 333.600 ;
        RECT 115.950 331.950 118.050 332.400 ;
        RECT 124.950 331.950 127.050 332.400 ;
        RECT 136.950 333.600 139.050 334.050 ;
        RECT 145.950 333.600 148.050 333.900 ;
        RECT 136.950 332.400 148.050 333.600 ;
        RECT 136.950 331.950 139.050 332.400 ;
        RECT 145.950 331.800 148.050 332.400 ;
        RECT 163.950 333.600 166.050 333.900 ;
        RECT 187.950 333.600 190.050 334.050 ;
        RECT 163.950 332.400 190.050 333.600 ;
        RECT 163.950 331.800 166.050 332.400 ;
        RECT 187.950 331.950 190.050 332.400 ;
        RECT 196.950 333.600 199.050 333.900 ;
        RECT 196.950 332.400 201.600 333.600 ;
        RECT 196.950 331.800 199.050 332.400 ;
        RECT 49.950 329.400 57.600 330.600 ;
        RECT 67.950 330.600 70.050 331.050 ;
        RECT 112.950 330.600 115.050 331.050 ;
        RECT 67.950 329.400 115.050 330.600 ;
        RECT 200.400 330.600 201.600 332.400 ;
        RECT 217.950 333.450 220.050 333.900 ;
        RECT 235.950 333.450 238.050 333.900 ;
        RECT 217.950 332.250 238.050 333.450 ;
        RECT 217.950 331.800 220.050 332.250 ;
        RECT 235.950 331.800 238.050 332.250 ;
        RECT 253.950 331.950 256.050 334.050 ;
        RECT 259.950 333.600 262.050 334.050 ;
        RECT 287.400 333.600 288.600 338.100 ;
        RECT 298.950 337.950 301.050 338.400 ;
        RECT 307.950 338.250 310.050 338.400 ;
        RECT 313.950 336.600 316.050 340.050 ;
        RECT 322.950 339.600 325.050 340.350 ;
        RECT 331.950 339.600 334.050 340.050 ;
        RECT 322.950 338.400 334.050 339.600 ;
        RECT 322.950 338.250 325.050 338.400 ;
        RECT 331.950 337.950 334.050 338.400 ;
        RECT 313.950 336.000 318.600 336.600 ;
        RECT 314.400 335.400 319.050 336.000 ;
        RECT 259.950 332.400 288.600 333.600 ;
        RECT 289.950 333.600 292.050 333.900 ;
        RECT 304.950 333.600 307.050 334.050 ;
        RECT 289.950 332.400 307.050 333.600 ;
        RECT 259.950 331.950 262.050 332.400 ;
        RECT 289.950 331.800 292.050 332.400 ;
        RECT 304.950 331.950 307.050 332.400 ;
        RECT 316.950 331.950 319.050 335.400 ;
        RECT 341.400 333.900 342.600 340.950 ;
        RECT 366.000 339.600 370.050 340.050 ;
        RECT 382.950 339.600 385.050 340.050 ;
        RECT 391.950 339.600 394.050 340.200 ;
        RECT 365.400 337.950 370.050 339.600 ;
        RECT 371.400 338.400 385.050 339.600 ;
        RECT 340.950 331.800 343.050 333.900 ;
        RECT 358.950 333.600 361.050 333.900 ;
        RECT 365.400 333.600 366.600 337.950 ;
        RECT 371.400 336.600 372.600 338.400 ;
        RECT 382.950 337.950 385.050 338.400 ;
        RECT 389.400 338.400 394.050 339.600 ;
        RECT 385.950 336.600 388.050 337.050 ;
        RECT 368.400 336.000 372.600 336.600 ;
        RECT 358.950 332.400 366.600 333.600 ;
        RECT 367.950 335.400 372.600 336.000 ;
        RECT 374.400 335.400 388.050 336.600 ;
        RECT 358.950 331.800 361.050 332.400 ;
        RECT 367.950 331.950 370.050 335.400 ;
        RECT 374.400 333.900 375.600 335.400 ;
        RECT 385.950 334.950 388.050 335.400 ;
        RECT 389.400 334.050 390.600 338.400 ;
        RECT 391.950 338.100 394.050 338.400 ;
        RECT 421.950 338.100 424.050 340.200 ;
        RECT 430.950 339.600 433.050 340.050 ;
        RECT 490.950 339.600 493.050 340.200 ;
        RECT 430.950 338.400 493.050 339.600 ;
        RECT 422.400 334.050 423.600 338.100 ;
        RECT 430.950 337.950 433.050 338.400 ;
        RECT 490.950 338.100 493.050 338.400 ;
        RECT 499.950 338.100 502.050 340.200 ;
        RECT 505.950 339.600 508.050 340.200 ;
        RECT 511.950 339.600 514.050 343.050 ;
        RECT 601.950 342.600 604.050 343.050 ;
        RECT 634.950 342.600 637.050 343.050 ;
        RECT 640.950 342.600 643.050 343.050 ;
        RECT 601.950 341.400 643.050 342.600 ;
        RECT 601.950 340.950 604.050 341.400 ;
        RECT 634.950 340.950 637.050 341.400 ;
        RECT 640.950 340.950 643.050 341.400 ;
        RECT 697.950 342.600 700.050 343.050 ;
        RECT 733.950 342.600 736.050 343.050 ;
        RECT 760.950 342.600 763.050 343.050 ;
        RECT 697.950 341.400 763.050 342.600 ;
        RECT 697.950 340.950 700.050 341.400 ;
        RECT 733.950 340.950 736.050 341.400 ;
        RECT 760.950 340.950 763.050 341.400 ;
        RECT 847.950 340.950 850.050 343.050 ;
        RECT 853.950 340.950 856.050 343.050 ;
        RECT 505.950 339.000 514.050 339.600 ;
        RECT 514.950 339.600 517.050 340.050 ;
        RECT 526.950 339.600 529.050 340.350 ;
        RECT 505.950 338.400 513.600 339.000 ;
        RECT 514.950 338.400 529.050 339.600 ;
        RECT 505.950 338.100 508.050 338.400 ;
        RECT 500.400 336.600 501.600 338.100 ;
        RECT 514.950 337.950 517.050 338.400 ;
        RECT 526.950 338.250 529.050 338.400 ;
        RECT 535.950 338.100 538.050 340.200 ;
        RECT 580.950 339.750 583.050 340.200 ;
        RECT 589.950 339.750 592.050 340.200 ;
        RECT 580.950 338.550 592.050 339.750 ;
        RECT 580.950 338.100 583.050 338.550 ;
        RECT 589.950 338.100 592.050 338.550 ;
        RECT 643.950 339.600 646.050 339.900 ;
        RECT 652.950 339.600 655.050 340.350 ;
        RECT 667.950 339.600 670.050 340.200 ;
        RECT 643.950 338.400 655.050 339.600 ;
        RECT 500.400 335.400 519.600 336.600 ;
        RECT 373.950 331.800 376.050 333.900 ;
        RECT 388.950 331.950 391.050 334.050 ;
        RECT 403.950 333.450 406.050 333.900 ;
        RECT 412.950 333.450 415.050 333.900 ;
        RECT 403.950 332.250 415.050 333.450 ;
        RECT 422.400 332.400 426.900 334.050 ;
        RECT 403.950 331.800 406.050 332.250 ;
        RECT 412.950 331.800 415.050 332.250 ;
        RECT 423.000 331.950 426.900 332.400 ;
        RECT 427.950 333.600 430.050 334.050 ;
        RECT 460.950 333.600 463.050 333.900 ;
        RECT 427.950 332.400 463.050 333.600 ;
        RECT 427.950 331.950 430.050 332.400 ;
        RECT 460.950 331.800 463.050 332.400 ;
        RECT 508.950 333.450 511.050 333.900 ;
        RECT 514.950 333.450 517.050 333.900 ;
        RECT 508.950 332.250 517.050 333.450 ;
        RECT 518.400 333.600 519.600 335.400 ;
        RECT 523.950 333.600 526.050 334.050 ;
        RECT 518.400 332.400 526.050 333.600 ;
        RECT 508.950 331.800 511.050 332.250 ;
        RECT 514.950 331.800 517.050 332.250 ;
        RECT 523.950 331.950 526.050 332.400 ;
        RECT 529.950 333.600 532.050 334.050 ;
        RECT 536.400 333.600 537.600 338.100 ;
        RECT 643.950 337.800 646.050 338.400 ;
        RECT 652.950 338.250 655.050 338.400 ;
        RECT 656.400 338.400 670.050 339.600 ;
        RECT 656.400 336.600 657.600 338.400 ;
        RECT 667.950 338.100 670.050 338.400 ;
        RECT 691.950 338.250 694.050 340.350 ;
        RECT 724.950 339.600 727.050 340.050 ;
        RECT 742.950 339.600 745.050 340.200 ;
        RECT 724.950 338.400 745.050 339.600 ;
        RECT 650.400 336.000 657.600 336.600 ;
        RECT 649.950 335.400 657.600 336.000 ;
        RECT 692.400 336.600 693.600 338.250 ;
        RECT 724.950 337.950 727.050 338.400 ;
        RECT 742.950 338.100 745.050 338.400 ;
        RECT 772.950 339.750 775.050 340.200 ;
        RECT 778.950 339.750 781.050 340.200 ;
        RECT 772.950 338.550 781.050 339.750 ;
        RECT 772.950 338.100 775.050 338.550 ;
        RECT 778.950 338.100 781.050 338.550 ;
        RECT 796.950 338.100 799.050 340.200 ;
        RECT 820.950 339.750 823.050 340.200 ;
        RECT 829.950 339.750 832.050 340.200 ;
        RECT 820.950 338.550 832.050 339.750 ;
        RECT 843.000 339.600 847.050 340.050 ;
        RECT 820.950 338.100 823.050 338.550 ;
        RECT 829.950 338.100 832.050 338.550 ;
        RECT 700.950 336.600 703.050 337.050 ;
        RECT 692.400 335.400 703.050 336.600 ;
        RECT 797.400 336.600 798.600 338.100 ;
        RECT 842.400 337.950 847.050 339.600 ;
        RECT 797.400 336.000 816.600 336.600 ;
        RECT 797.400 335.400 817.050 336.000 ;
        RECT 562.950 333.600 565.050 333.900 ;
        RECT 529.950 332.400 537.600 333.600 ;
        RECT 551.400 332.400 565.050 333.600 ;
        RECT 529.950 331.950 532.050 332.400 ;
        RECT 211.950 330.600 214.050 331.050 ;
        RECT 223.950 330.600 226.050 331.050 ;
        RECT 200.400 329.400 226.050 330.600 ;
        RECT 49.950 328.950 52.050 329.400 ;
        RECT 67.950 328.950 70.050 329.400 ;
        RECT 112.950 328.950 115.050 329.400 ;
        RECT 211.950 328.950 214.050 329.400 ;
        RECT 223.950 328.950 226.050 329.400 ;
        RECT 379.950 330.600 382.050 331.050 ;
        RECT 385.950 330.600 388.050 331.050 ;
        RECT 379.950 329.400 388.050 330.600 ;
        RECT 379.950 328.950 382.050 329.400 ;
        RECT 385.950 328.950 388.050 329.400 ;
        RECT 418.950 330.600 421.050 331.050 ;
        RECT 433.950 330.600 436.050 331.050 ;
        RECT 418.950 329.400 436.050 330.600 ;
        RECT 418.950 328.950 421.050 329.400 ;
        RECT 433.950 328.950 436.050 329.400 ;
        RECT 532.950 330.600 535.050 331.050 ;
        RECT 551.400 330.600 552.600 332.400 ;
        RECT 562.950 331.800 565.050 332.400 ;
        RECT 577.950 333.600 580.050 333.900 ;
        RECT 598.950 333.600 601.050 333.900 ;
        RECT 577.950 332.400 601.050 333.600 ;
        RECT 577.950 331.800 580.050 332.400 ;
        RECT 598.950 331.800 601.050 332.400 ;
        RECT 649.950 331.950 652.050 335.400 ;
        RECT 700.950 334.950 703.050 335.400 ;
        RECT 655.950 333.600 658.050 334.050 ;
        RECT 664.950 333.600 667.050 333.900 ;
        RECT 655.950 332.400 667.050 333.600 ;
        RECT 655.950 331.950 658.050 332.400 ;
        RECT 664.950 331.800 667.050 332.400 ;
        RECT 673.950 333.600 676.050 333.900 ;
        RECT 685.950 333.600 688.050 334.050 ;
        RECT 673.950 332.400 688.050 333.600 ;
        RECT 673.950 331.800 676.050 332.400 ;
        RECT 685.950 331.950 688.050 332.400 ;
        RECT 703.950 333.450 706.050 333.900 ;
        RECT 709.950 333.450 712.050 333.900 ;
        RECT 703.950 332.250 712.050 333.450 ;
        RECT 703.950 331.800 706.050 332.250 ;
        RECT 709.950 331.800 712.050 332.250 ;
        RECT 715.950 333.600 718.050 333.900 ;
        RECT 724.950 333.600 727.050 333.900 ;
        RECT 715.950 333.450 727.050 333.600 ;
        RECT 730.950 333.450 733.050 333.900 ;
        RECT 715.950 332.400 733.050 333.450 ;
        RECT 715.950 331.800 718.050 332.400 ;
        RECT 724.950 332.250 733.050 332.400 ;
        RECT 724.950 331.800 727.050 332.250 ;
        RECT 730.950 331.800 733.050 332.250 ;
        RECT 763.950 333.600 766.050 333.900 ;
        RECT 772.950 333.600 775.050 334.050 ;
        RECT 763.950 332.400 775.050 333.600 ;
        RECT 763.950 331.800 766.050 332.400 ;
        RECT 772.950 331.950 775.050 332.400 ;
        RECT 814.950 331.950 817.050 335.400 ;
        RECT 842.400 334.050 843.600 337.950 ;
        RECT 841.950 331.950 844.050 334.050 ;
        RECT 848.400 331.050 849.600 340.950 ;
        RECT 854.400 334.050 855.600 340.950 ;
        RECT 853.950 331.950 856.050 334.050 ;
        RECT 532.950 329.400 552.600 330.600 ;
        RECT 562.950 330.600 565.050 331.050 ;
        RECT 607.950 330.600 610.050 331.050 ;
        RECT 562.950 329.400 610.050 330.600 ;
        RECT 532.950 328.950 535.050 329.400 ;
        RECT 562.950 328.950 565.050 329.400 ;
        RECT 607.950 328.950 610.050 329.400 ;
        RECT 745.950 330.600 748.050 331.050 ;
        RECT 754.950 330.600 757.050 331.050 ;
        RECT 745.950 329.400 757.050 330.600 ;
        RECT 848.400 329.400 853.050 331.050 ;
        RECT 745.950 328.950 748.050 329.400 ;
        RECT 754.950 328.950 757.050 329.400 ;
        RECT 849.000 328.950 853.050 329.400 ;
        RECT 106.950 327.600 109.050 328.050 ;
        RECT 139.950 327.600 142.050 328.050 ;
        RECT 106.950 326.400 142.050 327.600 ;
        RECT 106.950 325.950 109.050 326.400 ;
        RECT 139.950 325.950 142.050 326.400 ;
        RECT 151.950 327.600 154.050 328.050 ;
        RECT 208.950 327.600 211.050 328.050 ;
        RECT 151.950 326.400 211.050 327.600 ;
        RECT 151.950 325.950 154.050 326.400 ;
        RECT 208.950 325.950 211.050 326.400 ;
        RECT 241.950 327.600 244.050 328.050 ;
        RECT 265.950 327.600 268.050 328.050 ;
        RECT 319.950 327.600 322.050 328.050 ;
        RECT 241.950 326.400 322.050 327.600 ;
        RECT 241.950 325.950 244.050 326.400 ;
        RECT 265.950 325.950 268.050 326.400 ;
        RECT 319.950 325.950 322.050 326.400 ;
        RECT 517.950 327.600 520.050 328.050 ;
        RECT 553.950 327.600 556.050 328.050 ;
        RECT 517.950 326.400 556.050 327.600 ;
        RECT 517.950 325.950 520.050 326.400 ;
        RECT 553.950 325.950 556.050 326.400 ;
        RECT 589.950 327.600 592.050 328.050 ;
        RECT 616.950 327.600 619.050 328.050 ;
        RECT 589.950 326.400 619.050 327.600 ;
        RECT 589.950 325.950 592.050 326.400 ;
        RECT 616.950 325.950 619.050 326.400 ;
        RECT 664.950 327.600 667.050 328.050 ;
        RECT 679.950 327.600 682.050 328.050 ;
        RECT 664.950 326.400 682.050 327.600 ;
        RECT 664.950 325.950 667.050 326.400 ;
        RECT 679.950 325.950 682.050 326.400 ;
        RECT 790.950 327.600 793.050 328.050 ;
        RECT 832.950 327.600 835.050 328.050 ;
        RECT 790.950 326.400 835.050 327.600 ;
        RECT 790.950 325.950 793.050 326.400 ;
        RECT 832.950 325.950 835.050 326.400 ;
        RECT 82.950 324.600 85.050 325.050 ;
        RECT 130.950 324.600 133.050 325.050 ;
        RECT 82.950 323.400 133.050 324.600 ;
        RECT 82.950 322.950 85.050 323.400 ;
        RECT 130.950 322.950 133.050 323.400 ;
        RECT 145.950 324.600 148.050 325.050 ;
        RECT 217.950 324.600 220.050 325.050 ;
        RECT 145.950 323.400 220.050 324.600 ;
        RECT 145.950 322.950 148.050 323.400 ;
        RECT 217.950 322.950 220.050 323.400 ;
        RECT 331.950 324.600 334.050 325.050 ;
        RECT 502.950 324.600 505.050 325.050 ;
        RECT 331.950 323.400 505.050 324.600 ;
        RECT 331.950 322.950 334.050 323.400 ;
        RECT 502.950 322.950 505.050 323.400 ;
        RECT 640.950 324.600 643.050 325.050 ;
        RECT 655.950 324.600 658.050 325.050 ;
        RECT 640.950 323.400 658.050 324.600 ;
        RECT 640.950 322.950 643.050 323.400 ;
        RECT 655.950 322.950 658.050 323.400 ;
        RECT 115.950 321.600 118.050 322.050 ;
        RECT 172.950 321.600 175.050 322.050 ;
        RECT 115.950 320.400 175.050 321.600 ;
        RECT 115.950 319.950 118.050 320.400 ;
        RECT 172.950 319.950 175.050 320.400 ;
        RECT 271.950 321.600 274.050 322.050 ;
        RECT 292.950 321.600 295.050 322.050 ;
        RECT 271.950 320.400 295.050 321.600 ;
        RECT 271.950 319.950 274.050 320.400 ;
        RECT 292.950 319.950 295.050 320.400 ;
        RECT 298.950 321.600 301.050 322.050 ;
        RECT 325.950 321.600 328.050 322.050 ;
        RECT 298.950 320.400 328.050 321.600 ;
        RECT 298.950 319.950 301.050 320.400 ;
        RECT 325.950 319.950 328.050 320.400 ;
        RECT 397.950 321.600 400.050 322.050 ;
        RECT 454.950 321.600 457.050 322.050 ;
        RECT 757.950 321.600 760.050 322.050 ;
        RECT 769.950 321.600 772.050 322.050 ;
        RECT 817.950 321.600 820.050 322.050 ;
        RECT 397.950 320.400 501.600 321.600 ;
        RECT 397.950 319.950 400.050 320.400 ;
        RECT 454.950 319.950 457.050 320.400 ;
        RECT 500.400 318.600 501.600 320.400 ;
        RECT 757.950 320.400 820.050 321.600 ;
        RECT 757.950 319.950 760.050 320.400 ;
        RECT 769.950 319.950 772.050 320.400 ;
        RECT 817.950 319.950 820.050 320.400 ;
        RECT 514.950 318.600 517.050 319.050 ;
        RECT 500.400 317.400 517.050 318.600 ;
        RECT 514.950 316.950 517.050 317.400 ;
        RECT 643.950 318.600 646.050 319.050 ;
        RECT 700.950 318.600 703.050 319.050 ;
        RECT 721.950 318.600 724.050 319.050 ;
        RECT 805.950 318.600 808.050 319.050 ;
        RECT 643.950 317.400 808.050 318.600 ;
        RECT 643.950 316.950 646.050 317.400 ;
        RECT 700.950 316.950 703.050 317.400 ;
        RECT 721.950 316.950 724.050 317.400 ;
        RECT 805.950 316.950 808.050 317.400 ;
        RECT 814.950 318.600 817.050 319.050 ;
        RECT 847.950 318.600 850.050 319.050 ;
        RECT 814.950 317.400 850.050 318.600 ;
        RECT 814.950 316.950 817.050 317.400 ;
        RECT 847.950 316.950 850.050 317.400 ;
        RECT 280.950 315.600 283.050 316.050 ;
        RECT 310.950 315.600 313.050 316.050 ;
        RECT 280.950 314.400 313.050 315.600 ;
        RECT 280.950 313.950 283.050 314.400 ;
        RECT 310.950 313.950 313.050 314.400 ;
        RECT 592.950 315.600 595.050 316.050 ;
        RECT 613.950 315.600 616.050 316.050 ;
        RECT 592.950 314.400 616.050 315.600 ;
        RECT 592.950 313.950 595.050 314.400 ;
        RECT 613.950 313.950 616.050 314.400 ;
        RECT 781.950 315.600 784.050 316.050 ;
        RECT 796.950 315.600 799.050 316.050 ;
        RECT 781.950 314.400 799.050 315.600 ;
        RECT 781.950 313.950 784.050 314.400 ;
        RECT 796.950 313.950 799.050 314.400 ;
        RECT 37.950 312.600 40.050 313.050 ;
        RECT 52.950 312.600 55.050 313.050 ;
        RECT 37.950 311.400 55.050 312.600 ;
        RECT 37.950 310.950 40.050 311.400 ;
        RECT 52.950 310.950 55.050 311.400 ;
        RECT 400.950 312.600 403.050 313.050 ;
        RECT 424.950 312.600 427.050 313.050 ;
        RECT 484.950 312.600 487.050 313.050 ;
        RECT 568.950 312.600 571.050 313.050 ;
        RECT 400.950 311.400 571.050 312.600 ;
        RECT 400.950 310.950 403.050 311.400 ;
        RECT 424.950 310.950 427.050 311.400 ;
        RECT 484.950 310.950 487.050 311.400 ;
        RECT 568.950 310.950 571.050 311.400 ;
        RECT 28.950 309.600 31.050 310.050 ;
        RECT 67.950 309.600 70.050 310.050 ;
        RECT 28.950 308.400 70.050 309.600 ;
        RECT 28.950 307.950 31.050 308.400 ;
        RECT 67.950 307.950 70.050 308.400 ;
        RECT 79.950 309.600 82.050 310.050 ;
        RECT 151.950 309.600 154.050 310.050 ;
        RECT 79.950 308.400 154.050 309.600 ;
        RECT 79.950 307.950 82.050 308.400 ;
        RECT 151.950 307.950 154.050 308.400 ;
        RECT 199.950 309.600 202.050 310.050 ;
        RECT 250.950 309.600 253.050 310.050 ;
        RECT 199.950 308.400 253.050 309.600 ;
        RECT 199.950 307.950 202.050 308.400 ;
        RECT 250.950 307.950 253.050 308.400 ;
        RECT 472.950 309.600 475.050 310.050 ;
        RECT 532.950 309.600 535.050 310.050 ;
        RECT 472.950 308.400 535.050 309.600 ;
        RECT 472.950 307.950 475.050 308.400 ;
        RECT 532.950 307.950 535.050 308.400 ;
        RECT 604.950 309.600 607.050 310.050 ;
        RECT 793.950 309.600 796.050 310.050 ;
        RECT 814.950 309.600 817.050 310.050 ;
        RECT 604.950 309.000 681.600 309.600 ;
        RECT 604.950 308.400 682.050 309.000 ;
        RECT 604.950 307.950 607.050 308.400 ;
        RECT 10.950 306.600 13.050 307.050 ;
        RECT 16.950 306.600 19.050 307.050 ;
        RECT 10.950 305.400 19.050 306.600 ;
        RECT 10.950 304.950 13.050 305.400 ;
        RECT 16.950 304.950 19.050 305.400 ;
        RECT 148.950 306.600 151.050 307.050 ;
        RECT 169.950 306.600 172.050 307.050 ;
        RECT 148.950 305.400 172.050 306.600 ;
        RECT 148.950 304.950 151.050 305.400 ;
        RECT 169.950 304.950 172.050 305.400 ;
        RECT 193.950 306.600 196.050 307.050 ;
        RECT 265.950 306.600 268.050 307.050 ;
        RECT 193.950 305.400 268.050 306.600 ;
        RECT 193.950 304.950 196.050 305.400 ;
        RECT 265.950 304.950 268.050 305.400 ;
        RECT 277.950 306.600 280.050 307.050 ;
        RECT 301.950 306.600 304.050 307.050 ;
        RECT 277.950 305.400 304.050 306.600 ;
        RECT 277.950 304.950 280.050 305.400 ;
        RECT 301.950 304.950 304.050 305.400 ;
        RECT 547.950 306.600 550.050 307.050 ;
        RECT 598.950 306.600 601.050 307.050 ;
        RECT 547.950 305.400 601.050 306.600 ;
        RECT 547.950 304.950 550.050 305.400 ;
        RECT 598.950 304.950 601.050 305.400 ;
        RECT 679.950 304.950 682.050 308.400 ;
        RECT 793.950 308.400 817.050 309.600 ;
        RECT 793.950 307.950 796.050 308.400 ;
        RECT 814.950 307.950 817.050 308.400 ;
        RECT 697.950 306.600 700.050 307.050 ;
        RECT 751.950 306.600 754.050 307.050 ;
        RECT 697.950 305.400 754.050 306.600 ;
        RECT 697.950 304.950 700.050 305.400 ;
        RECT 751.950 304.950 754.050 305.400 ;
        RECT 4.950 303.600 7.050 304.050 ;
        RECT 34.950 303.600 37.050 304.050 ;
        RECT 4.950 302.400 37.050 303.600 ;
        RECT 4.950 301.950 7.050 302.400 ;
        RECT 34.950 301.950 37.050 302.400 ;
        RECT 76.950 303.600 79.050 304.050 ;
        RECT 118.950 303.600 121.050 304.050 ;
        RECT 430.950 303.600 433.050 304.050 ;
        RECT 460.950 303.600 463.050 304.050 ;
        RECT 76.950 302.400 372.600 303.600 ;
        RECT 76.950 301.950 79.050 302.400 ;
        RECT 118.950 301.950 121.050 302.400 ;
        RECT 371.400 301.050 372.600 302.400 ;
        RECT 430.950 302.400 463.050 303.600 ;
        RECT 430.950 301.950 433.050 302.400 ;
        RECT 460.950 301.950 463.050 302.400 ;
        RECT 529.950 303.600 532.050 304.050 ;
        RECT 535.950 303.600 538.050 304.050 ;
        RECT 529.950 302.400 538.050 303.600 ;
        RECT 529.950 301.950 532.050 302.400 ;
        RECT 535.950 301.950 538.050 302.400 ;
        RECT 640.950 303.600 643.050 304.050 ;
        RECT 646.950 303.600 649.050 304.050 ;
        RECT 640.950 302.400 649.050 303.600 ;
        RECT 640.950 301.950 643.050 302.400 ;
        RECT 646.950 301.950 649.050 302.400 ;
        RECT 691.950 303.600 694.050 304.050 ;
        RECT 739.950 303.600 742.050 304.050 ;
        RECT 691.950 302.400 742.050 303.600 ;
        RECT 691.950 301.950 694.050 302.400 ;
        RECT 739.950 301.950 742.050 302.400 ;
        RECT 802.950 303.600 805.050 304.050 ;
        RECT 811.950 303.600 814.050 304.050 ;
        RECT 802.950 302.400 814.050 303.600 ;
        RECT 802.950 301.950 805.050 302.400 ;
        RECT 811.950 301.950 814.050 302.400 ;
        RECT 256.950 300.600 259.050 301.050 ;
        RECT 286.950 300.600 289.050 301.050 ;
        RECT 256.950 299.400 289.050 300.600 ;
        RECT 256.950 298.950 259.050 299.400 ;
        RECT 286.950 298.950 289.050 299.400 ;
        RECT 370.950 300.600 373.050 301.050 ;
        RECT 388.950 300.600 391.050 301.050 ;
        RECT 370.950 299.400 391.050 300.600 ;
        RECT 370.950 298.950 373.050 299.400 ;
        RECT 388.950 298.950 391.050 299.400 ;
        RECT 574.950 300.600 577.050 301.050 ;
        RECT 592.950 300.600 595.050 301.050 ;
        RECT 574.950 299.400 595.050 300.600 ;
        RECT 574.950 298.950 577.050 299.400 ;
        RECT 592.950 298.950 595.050 299.400 ;
        RECT 727.950 300.600 730.050 301.050 ;
        RECT 793.950 300.600 796.050 301.050 ;
        RECT 727.950 299.400 796.050 300.600 ;
        RECT 727.950 298.950 730.050 299.400 ;
        RECT 793.950 298.950 796.050 299.400 ;
        RECT 838.950 300.600 841.050 301.050 ;
        RECT 859.950 300.600 862.050 301.050 ;
        RECT 838.950 299.400 862.050 300.600 ;
        RECT 838.950 298.950 841.050 299.400 ;
        RECT 859.950 298.950 862.050 299.400 ;
        RECT 223.950 297.600 226.050 298.050 ;
        RECT 316.950 297.600 319.050 298.050 ;
        RECT 223.950 296.400 319.050 297.600 ;
        RECT 223.950 295.950 226.050 296.400 ;
        RECT 316.950 295.950 319.050 296.400 ;
        RECT 355.950 297.600 358.050 298.050 ;
        RECT 361.950 297.600 364.050 298.050 ;
        RECT 418.950 297.600 421.050 298.050 ;
        RECT 355.950 296.400 364.050 297.600 ;
        RECT 355.950 295.950 358.050 296.400 ;
        RECT 361.950 295.950 364.050 296.400 ;
        RECT 383.400 296.400 421.050 297.600 ;
        RECT 16.950 294.600 19.050 295.050 ;
        RECT 28.950 294.600 31.050 295.050 ;
        RECT 16.950 293.400 31.050 294.600 ;
        RECT 16.950 292.950 19.050 293.400 ;
        RECT 28.950 292.950 31.050 293.400 ;
        RECT 37.950 292.950 40.050 295.050 ;
        RECT 46.950 294.750 49.050 295.200 ;
        RECT 58.950 294.750 61.050 295.050 ;
        RECT 64.950 294.750 67.050 295.200 ;
        RECT 46.950 293.550 67.050 294.750 ;
        RECT 75.000 294.600 79.050 295.050 ;
        RECT 46.950 293.100 49.050 293.550 ;
        RECT 58.950 292.950 61.050 293.550 ;
        RECT 64.950 293.100 67.050 293.550 ;
        RECT 74.400 292.950 79.050 294.600 ;
        RECT 82.950 293.100 85.050 295.200 ;
        RECT 91.950 294.750 94.050 295.200 ;
        RECT 97.950 294.750 100.050 295.200 ;
        RECT 91.950 293.550 100.050 294.750 ;
        RECT 91.950 293.100 94.050 293.550 ;
        RECT 97.950 293.100 100.050 293.550 ;
        RECT 4.950 288.600 7.050 289.050 ;
        RECT 38.400 288.750 39.600 292.950 ;
        RECT 74.400 288.900 75.600 292.950 ;
        RECT 13.950 288.600 16.050 288.750 ;
        RECT 4.950 287.400 16.050 288.600 ;
        RECT 4.950 286.950 7.050 287.400 ;
        RECT 13.950 286.650 16.050 287.400 ;
        RECT 37.950 286.650 40.050 288.750 ;
        RECT 73.950 286.800 76.050 288.900 ;
        RECT 58.950 285.600 61.050 286.050 ;
        RECT 64.950 285.600 67.050 286.050 ;
        RECT 83.400 285.600 84.600 293.100 ;
        RECT 124.950 292.950 127.050 295.050 ;
        RECT 130.950 294.600 133.050 295.050 ;
        RECT 136.950 294.600 139.050 295.050 ;
        RECT 130.950 293.400 139.050 294.600 ;
        RECT 130.950 292.950 133.050 293.400 ;
        RECT 136.950 292.950 139.050 293.400 ;
        RECT 142.950 293.100 145.050 295.200 ;
        RECT 172.950 294.750 175.050 295.200 ;
        RECT 184.950 294.750 187.050 295.200 ;
        RECT 172.950 293.550 187.050 294.750 ;
        RECT 172.950 293.100 175.050 293.550 ;
        RECT 184.950 293.100 187.050 293.550 ;
        RECT 125.400 289.050 126.600 292.950 ;
        RECT 121.950 287.400 126.600 289.050 ;
        RECT 127.950 288.600 130.050 288.750 ;
        RECT 143.400 288.600 144.600 293.100 ;
        RECT 202.950 291.600 205.050 295.050 ;
        RECT 226.950 294.600 229.050 295.050 ;
        RECT 253.950 294.600 256.050 295.050 ;
        RECT 226.950 293.400 256.050 294.600 ;
        RECT 226.950 292.950 229.050 293.400 ;
        RECT 253.950 292.950 256.050 293.400 ;
        RECT 274.950 294.600 277.050 295.050 ;
        RECT 306.000 294.600 310.050 295.050 ;
        RECT 274.950 293.400 282.600 294.600 ;
        RECT 274.950 292.950 277.050 293.400 ;
        RECT 202.950 291.000 207.600 291.600 ;
        RECT 203.400 290.400 207.600 291.000 ;
        RECT 127.950 287.400 144.600 288.600 ;
        RECT 160.950 288.600 163.050 288.900 ;
        RECT 169.950 288.600 172.050 289.050 ;
        RECT 160.950 287.400 172.050 288.600 ;
        RECT 121.950 286.950 126.000 287.400 ;
        RECT 127.950 286.650 130.050 287.400 ;
        RECT 160.950 286.800 163.050 287.400 ;
        RECT 169.950 286.950 172.050 287.400 ;
        RECT 187.950 288.600 190.050 288.900 ;
        RECT 202.950 288.600 205.050 288.750 ;
        RECT 187.950 287.400 205.050 288.600 ;
        RECT 206.400 288.600 207.600 290.400 ;
        RECT 281.400 289.050 282.600 293.400 ;
        RECT 305.400 292.950 310.050 294.600 ;
        RECT 313.950 294.600 316.050 295.050 ;
        RECT 322.950 294.600 325.050 295.200 ;
        RECT 383.400 295.050 384.600 296.400 ;
        RECT 418.950 295.950 421.050 296.400 ;
        RECT 433.950 297.600 438.000 298.050 ;
        RECT 523.950 297.600 526.050 298.050 ;
        RECT 544.950 297.600 547.050 298.050 ;
        RECT 568.950 297.600 571.050 298.050 ;
        RECT 433.950 295.950 438.600 297.600 ;
        RECT 523.950 296.400 571.050 297.600 ;
        RECT 523.950 295.950 526.050 296.400 ;
        RECT 544.950 295.950 547.050 296.400 ;
        RECT 568.950 295.950 571.050 296.400 ;
        RECT 625.950 297.600 628.050 298.050 ;
        RECT 631.950 297.600 634.050 298.050 ;
        RECT 646.950 297.600 649.050 298.050 ;
        RECT 625.950 296.400 649.050 297.600 ;
        RECT 625.950 295.950 628.050 296.400 ;
        RECT 631.950 295.950 634.050 296.400 ;
        RECT 646.950 295.950 649.050 296.400 ;
        RECT 670.950 297.600 673.050 298.050 ;
        RECT 697.950 297.600 700.050 298.050 ;
        RECT 670.950 296.400 700.050 297.600 ;
        RECT 670.950 295.950 673.050 296.400 ;
        RECT 697.950 295.950 700.050 296.400 ;
        RECT 751.950 297.600 754.050 298.050 ;
        RECT 778.950 297.600 781.050 298.050 ;
        RECT 790.950 297.600 793.050 298.050 ;
        RECT 751.950 296.400 793.050 297.600 ;
        RECT 751.950 295.950 754.050 296.400 ;
        RECT 778.950 295.950 781.050 296.400 ;
        RECT 790.950 295.950 793.050 296.400 ;
        RECT 808.950 297.600 813.000 298.050 ;
        RECT 808.950 295.950 813.600 297.600 ;
        RECT 313.950 293.400 325.050 294.600 ;
        RECT 313.950 292.950 316.050 293.400 ;
        RECT 322.950 293.100 325.050 293.400 ;
        RECT 337.950 292.950 340.050 295.050 ;
        RECT 346.950 292.950 349.050 295.050 ;
        RECT 352.950 294.600 355.050 295.050 ;
        RECT 367.950 294.600 370.050 295.050 ;
        RECT 376.950 294.600 379.050 295.050 ;
        RECT 352.950 293.400 379.050 294.600 ;
        RECT 352.950 292.950 355.050 293.400 ;
        RECT 367.950 292.950 370.050 293.400 ;
        RECT 376.950 292.950 379.050 293.400 ;
        RECT 382.950 292.950 385.050 295.050 ;
        RECT 388.950 294.600 391.050 295.050 ;
        RECT 394.950 294.600 397.050 295.050 ;
        RECT 388.950 293.400 397.050 294.600 ;
        RECT 388.950 292.950 391.050 293.400 ;
        RECT 394.950 292.950 397.050 293.400 ;
        RECT 403.950 292.950 406.050 295.050 ;
        RECT 412.950 293.100 415.050 295.200 ;
        RECT 423.000 294.600 427.050 295.050 ;
        RECT 220.950 288.600 223.050 288.750 ;
        RECT 206.400 287.400 223.050 288.600 ;
        RECT 187.950 286.800 190.050 287.400 ;
        RECT 202.950 286.650 205.050 287.400 ;
        RECT 220.950 286.650 223.050 287.400 ;
        RECT 268.950 288.300 271.050 288.750 ;
        RECT 274.950 288.300 277.050 288.750 ;
        RECT 268.950 287.100 277.050 288.300 ;
        RECT 268.950 286.650 271.050 287.100 ;
        RECT 274.950 286.650 277.050 287.100 ;
        RECT 280.950 286.950 283.050 289.050 ;
        RECT 58.950 284.400 84.600 285.600 ;
        RECT 91.950 285.600 94.050 286.050 ;
        RECT 115.950 285.600 118.050 286.050 ;
        RECT 91.950 284.400 118.050 285.600 ;
        RECT 58.950 283.950 61.050 284.400 ;
        RECT 64.950 283.950 67.050 284.400 ;
        RECT 91.950 283.950 94.050 284.400 ;
        RECT 115.950 283.950 118.050 284.400 ;
        RECT 172.950 285.600 175.050 286.050 ;
        RECT 184.950 285.600 187.050 286.050 ;
        RECT 172.950 284.400 187.050 285.600 ;
        RECT 172.950 283.950 175.050 284.400 ;
        RECT 184.950 283.950 187.050 284.400 ;
        RECT 283.950 285.600 286.050 286.050 ;
        RECT 305.400 285.600 306.600 292.950 ;
        RECT 338.400 289.050 339.600 292.950 ;
        RECT 347.400 289.050 348.600 292.950 ;
        RECT 334.950 287.400 339.600 289.050 ;
        RECT 334.950 286.950 339.000 287.400 ;
        RECT 346.950 286.950 349.050 289.050 ;
        RECT 352.950 288.600 355.050 289.050 ;
        RECT 358.950 288.600 361.050 288.900 ;
        RECT 352.950 287.400 361.050 288.600 ;
        RECT 352.950 286.950 355.050 287.400 ;
        RECT 358.950 286.800 361.050 287.400 ;
        RECT 364.950 288.600 367.050 288.900 ;
        RECT 383.400 288.600 384.600 292.950 ;
        RECT 364.950 287.400 384.600 288.600 ;
        RECT 397.950 288.600 400.050 288.750 ;
        RECT 404.400 288.600 405.600 292.950 ;
        RECT 397.950 287.400 405.600 288.600 ;
        RECT 364.950 286.800 367.050 287.400 ;
        RECT 397.950 286.650 400.050 287.400 ;
        RECT 413.400 286.050 414.600 293.100 ;
        RECT 422.400 292.950 427.050 294.600 ;
        RECT 430.950 292.950 433.050 295.050 ;
        RECT 422.400 288.900 423.600 292.950 ;
        RECT 431.400 289.050 432.600 292.950 ;
        RECT 437.400 289.050 438.600 295.950 ;
        RECT 478.950 294.600 481.050 295.050 ;
        RECT 484.950 294.600 487.050 295.050 ;
        RECT 478.950 293.400 487.050 294.600 ;
        RECT 478.950 292.950 481.050 293.400 ;
        RECT 484.950 292.950 487.050 293.400 ;
        RECT 490.950 294.600 493.050 295.050 ;
        RECT 496.950 294.600 499.050 295.050 ;
        RECT 490.950 293.400 499.050 294.600 ;
        RECT 490.950 292.950 493.050 293.400 ;
        RECT 496.950 292.950 499.050 293.400 ;
        RECT 547.800 292.950 549.900 295.050 ;
        RECT 550.950 294.600 553.050 295.050 ;
        RECT 565.950 294.750 568.050 295.200 ;
        RECT 583.950 294.750 586.050 295.200 ;
        RECT 550.950 293.400 558.600 294.600 ;
        RECT 550.950 292.950 553.050 293.400 ;
        RECT 421.950 286.800 424.050 288.900 ;
        RECT 430.950 286.950 433.050 289.050 ;
        RECT 437.400 287.400 442.050 289.050 ;
        RECT 548.250 288.750 549.450 292.950 ;
        RECT 557.400 288.900 558.600 293.400 ;
        RECT 565.950 293.550 586.050 294.750 ;
        RECT 619.950 294.600 622.050 295.200 ;
        RECT 565.950 293.100 568.050 293.550 ;
        RECT 583.950 293.100 586.050 293.550 ;
        RECT 608.400 293.400 622.050 294.600 ;
        RECT 438.000 286.950 442.050 287.400 ;
        RECT 478.950 288.300 481.050 288.750 ;
        RECT 484.950 288.300 487.050 288.750 ;
        RECT 478.950 287.100 487.050 288.300 ;
        RECT 478.950 286.650 481.050 287.100 ;
        RECT 484.950 286.650 487.050 287.100 ;
        RECT 547.800 286.650 549.900 288.750 ;
        RECT 556.950 288.600 559.050 288.900 ;
        RECT 571.950 288.600 574.050 289.050 ;
        RECT 556.950 287.400 574.050 288.600 ;
        RECT 556.950 286.800 559.050 287.400 ;
        RECT 571.950 286.950 574.050 287.400 ;
        RECT 592.950 288.600 595.050 289.050 ;
        RECT 608.400 288.900 609.600 293.400 ;
        RECT 619.950 293.100 622.050 293.400 ;
        RECT 694.950 294.600 699.000 295.050 ;
        RECT 700.950 294.600 703.050 295.200 ;
        RECT 706.950 294.600 709.050 295.050 ;
        RECT 694.950 292.950 699.600 294.600 ;
        RECT 700.950 293.400 709.050 294.600 ;
        RECT 700.950 293.100 703.050 293.400 ;
        RECT 706.950 292.950 709.050 293.400 ;
        RECT 715.950 293.100 718.050 295.200 ;
        RECT 744.000 294.600 748.050 295.050 ;
        RECT 698.400 288.900 699.600 292.950 ;
        RECT 601.950 288.600 604.050 288.900 ;
        RECT 592.950 287.400 604.050 288.600 ;
        RECT 592.950 286.950 595.050 287.400 ;
        RECT 601.950 286.800 604.050 287.400 ;
        RECT 607.950 286.800 610.050 288.900 ;
        RECT 697.950 286.800 700.050 288.900 ;
        RECT 706.950 288.450 709.050 288.900 ;
        RECT 712.950 288.450 715.050 288.900 ;
        RECT 706.950 287.250 715.050 288.450 ;
        RECT 716.400 288.600 717.600 293.100 ;
        RECT 743.400 292.950 748.050 294.600 ;
        RECT 743.400 288.900 744.600 292.950 ;
        RECT 796.950 291.600 799.050 295.050 ;
        RECT 805.950 294.600 810.000 295.050 ;
        RECT 805.950 292.950 810.600 294.600 ;
        RECT 796.950 291.000 801.600 291.600 ;
        RECT 797.400 290.400 802.050 291.000 ;
        RECT 716.400 287.400 720.600 288.600 ;
        RECT 706.950 286.800 709.050 287.250 ;
        RECT 712.950 286.800 715.050 287.250 ;
        RECT 719.400 286.050 720.600 287.400 ;
        RECT 742.950 286.800 745.050 288.900 ;
        RECT 769.950 288.450 772.050 288.900 ;
        RECT 775.950 288.450 778.050 288.900 ;
        RECT 769.950 287.250 778.050 288.450 ;
        RECT 769.950 286.800 772.050 287.250 ;
        RECT 775.950 286.800 778.050 287.250 ;
        RECT 799.950 286.950 802.050 290.400 ;
        RECT 809.400 288.900 810.600 292.950 ;
        RECT 812.400 291.600 813.600 295.950 ;
        RECT 817.950 293.100 820.050 295.200 ;
        RECT 812.400 290.400 816.600 291.600 ;
        RECT 808.950 286.800 811.050 288.900 ;
        RECT 815.400 286.050 816.600 290.400 ;
        RECT 818.400 289.050 819.600 293.100 ;
        RECT 818.400 287.400 823.050 289.050 ;
        RECT 819.000 286.950 823.050 287.400 ;
        RECT 829.950 288.450 832.050 288.900 ;
        RECT 841.950 288.600 844.050 288.900 ;
        RECT 862.950 288.600 865.050 289.050 ;
        RECT 841.950 288.450 865.050 288.600 ;
        RECT 829.950 287.400 865.050 288.450 ;
        RECT 829.950 287.250 844.050 287.400 ;
        RECT 829.950 286.800 832.050 287.250 ;
        RECT 841.950 286.800 844.050 287.250 ;
        RECT 862.950 286.950 865.050 287.400 ;
        RECT 283.950 284.400 306.600 285.600 ;
        RECT 283.950 283.950 286.050 284.400 ;
        RECT 412.950 283.950 415.050 286.050 ;
        RECT 442.950 285.600 445.050 286.050 ;
        RECT 451.950 285.600 454.050 286.050 ;
        RECT 442.950 284.400 454.050 285.600 ;
        RECT 719.400 284.400 724.050 286.050 ;
        RECT 442.950 283.950 445.050 284.400 ;
        RECT 451.950 283.950 454.050 284.400 ;
        RECT 720.000 283.950 724.050 284.400 ;
        RECT 742.950 285.600 745.050 286.050 ;
        RECT 754.950 285.600 757.050 286.050 ;
        RECT 742.950 284.400 757.050 285.600 ;
        RECT 742.950 283.950 745.050 284.400 ;
        RECT 754.950 283.950 757.050 284.400 ;
        RECT 781.950 285.600 784.050 286.050 ;
        RECT 781.950 284.400 789.600 285.600 ;
        RECT 781.950 283.950 784.050 284.400 ;
        RECT 13.950 282.600 16.050 283.050 ;
        RECT 25.950 282.600 28.050 283.050 ;
        RECT 13.950 281.400 28.050 282.600 ;
        RECT 13.950 280.950 16.050 281.400 ;
        RECT 25.950 280.950 28.050 281.400 ;
        RECT 100.950 282.600 103.050 283.050 ;
        RECT 115.950 282.600 118.050 282.900 ;
        RECT 100.950 281.400 118.050 282.600 ;
        RECT 100.950 280.950 103.050 281.400 ;
        RECT 115.950 280.800 118.050 281.400 ;
        RECT 274.950 282.600 277.050 283.050 ;
        RECT 289.950 282.600 292.050 283.050 ;
        RECT 274.950 281.400 292.050 282.600 ;
        RECT 274.950 280.950 277.050 281.400 ;
        RECT 289.950 280.950 292.050 281.400 ;
        RECT 415.950 282.600 418.050 283.050 ;
        RECT 430.950 282.600 433.050 283.050 ;
        RECT 415.950 281.400 433.050 282.600 ;
        RECT 415.950 280.950 418.050 281.400 ;
        RECT 430.950 280.950 433.050 281.400 ;
        RECT 568.950 282.600 571.050 283.050 ;
        RECT 607.950 282.600 610.050 283.050 ;
        RECT 568.950 281.400 610.050 282.600 ;
        RECT 568.950 280.950 571.050 281.400 ;
        RECT 607.950 280.950 610.050 281.400 ;
        RECT 661.950 282.600 664.050 283.050 ;
        RECT 667.950 282.600 670.050 283.050 ;
        RECT 727.950 282.600 730.050 283.050 ;
        RECT 661.950 281.400 670.050 282.600 ;
        RECT 661.950 280.950 664.050 281.400 ;
        RECT 667.950 280.950 670.050 281.400 ;
        RECT 719.400 281.400 730.050 282.600 ;
        RECT 788.400 282.600 789.600 284.400 ;
        RECT 811.950 284.400 816.600 286.050 ;
        RECT 811.950 283.950 816.000 284.400 ;
        RECT 805.950 282.600 808.050 283.050 ;
        RECT 788.400 281.400 808.050 282.600 ;
        RECT 97.950 279.600 100.050 280.050 ;
        RECT 145.950 279.600 148.050 280.050 ;
        RECT 97.950 278.400 148.050 279.600 ;
        RECT 97.950 277.950 100.050 278.400 ;
        RECT 145.950 277.950 148.050 278.400 ;
        RECT 181.950 279.600 184.050 280.050 ;
        RECT 193.950 279.600 196.050 280.050 ;
        RECT 337.950 279.600 340.050 280.050 ;
        RECT 181.950 278.400 196.050 279.600 ;
        RECT 181.950 277.950 184.050 278.400 ;
        RECT 193.950 277.950 196.050 278.400 ;
        RECT 266.400 278.400 288.600 279.600 ;
        RECT 266.400 277.050 267.600 278.400 ;
        RECT 241.950 276.600 244.050 277.050 ;
        RECT 265.950 276.600 268.050 277.050 ;
        RECT 241.950 275.400 268.050 276.600 ;
        RECT 287.400 276.600 288.600 278.400 ;
        RECT 293.400 278.400 340.050 279.600 ;
        RECT 293.400 276.600 294.600 278.400 ;
        RECT 337.950 277.950 340.050 278.400 ;
        RECT 364.950 279.600 367.050 280.050 ;
        RECT 439.950 279.600 442.050 280.050 ;
        RECT 364.950 278.400 442.050 279.600 ;
        RECT 364.950 277.950 367.050 278.400 ;
        RECT 439.950 277.950 442.050 278.400 ;
        RECT 484.950 279.600 487.050 280.050 ;
        RECT 598.950 279.600 601.050 280.050 ;
        RECT 484.950 278.400 601.050 279.600 ;
        RECT 484.950 277.950 487.050 278.400 ;
        RECT 598.950 277.950 601.050 278.400 ;
        RECT 661.950 279.600 664.050 279.900 ;
        RECT 719.400 279.600 720.600 281.400 ;
        RECT 727.950 280.950 730.050 281.400 ;
        RECT 805.950 280.950 808.050 281.400 ;
        RECT 661.950 278.400 720.600 279.600 ;
        RECT 754.950 279.600 757.050 280.050 ;
        RECT 814.950 279.600 817.050 280.050 ;
        RECT 754.950 278.400 817.050 279.600 ;
        RECT 661.950 277.800 664.050 278.400 ;
        RECT 754.950 277.950 757.050 278.400 ;
        RECT 814.950 277.950 817.050 278.400 ;
        RECT 287.400 275.400 294.600 276.600 ;
        RECT 436.950 276.600 439.050 277.050 ;
        RECT 451.950 276.600 454.050 277.050 ;
        RECT 436.950 275.400 454.050 276.600 ;
        RECT 241.950 274.950 244.050 275.400 ;
        RECT 265.950 274.950 268.050 275.400 ;
        RECT 436.950 274.950 439.050 275.400 ;
        RECT 451.950 274.950 454.050 275.400 ;
        RECT 556.950 276.600 559.050 277.050 ;
        RECT 565.950 276.600 568.050 277.050 ;
        RECT 556.950 275.400 568.050 276.600 ;
        RECT 556.950 274.950 559.050 275.400 ;
        RECT 565.950 274.950 568.050 275.400 ;
        RECT 760.950 276.600 763.050 277.050 ;
        RECT 778.950 276.600 781.050 277.050 ;
        RECT 760.950 275.400 781.050 276.600 ;
        RECT 760.950 274.950 763.050 275.400 ;
        RECT 778.950 274.950 781.050 275.400 ;
        RECT 55.950 273.600 58.050 274.050 ;
        RECT 61.950 273.600 64.050 274.050 ;
        RECT 55.950 272.400 64.050 273.600 ;
        RECT 55.950 271.950 58.050 272.400 ;
        RECT 61.950 271.950 64.050 272.400 ;
        RECT 112.950 273.600 115.050 274.050 ;
        RECT 136.950 273.600 139.050 274.050 ;
        RECT 112.950 272.400 139.050 273.600 ;
        RECT 112.950 271.950 115.050 272.400 ;
        RECT 136.950 271.950 139.050 272.400 ;
        RECT 202.950 273.600 205.050 274.050 ;
        RECT 211.950 273.600 214.050 274.050 ;
        RECT 232.950 273.600 235.050 274.050 ;
        RECT 244.950 273.600 247.050 274.050 ;
        RECT 202.950 272.400 247.050 273.600 ;
        RECT 202.950 271.950 205.050 272.400 ;
        RECT 211.950 271.950 214.050 272.400 ;
        RECT 232.950 271.950 235.050 272.400 ;
        RECT 244.950 271.950 247.050 272.400 ;
        RECT 262.950 273.600 265.050 274.050 ;
        RECT 286.950 273.600 289.050 274.050 ;
        RECT 262.950 272.400 289.050 273.600 ;
        RECT 262.950 271.950 265.050 272.400 ;
        RECT 286.950 271.950 289.050 272.400 ;
        RECT 304.950 273.600 307.050 274.050 ;
        RECT 427.950 273.600 430.050 274.050 ;
        RECT 496.950 273.600 499.050 274.050 ;
        RECT 625.950 273.600 628.050 274.050 ;
        RECT 649.950 273.600 652.050 274.050 ;
        RECT 304.950 272.400 426.600 273.600 ;
        RECT 304.950 271.950 307.050 272.400 ;
        RECT 325.950 270.600 328.050 271.050 ;
        RECT 334.950 270.600 337.050 271.050 ;
        RECT 325.950 269.400 337.050 270.600 ;
        RECT 425.400 270.600 426.600 272.400 ;
        RECT 427.950 272.400 652.050 273.600 ;
        RECT 427.950 271.950 430.050 272.400 ;
        RECT 496.950 271.950 499.050 272.400 ;
        RECT 625.950 271.950 628.050 272.400 ;
        RECT 649.950 271.950 652.050 272.400 ;
        RECT 820.950 271.950 823.050 274.050 ;
        RECT 673.950 270.600 676.050 271.050 ;
        RECT 425.400 269.400 676.050 270.600 ;
        RECT 325.950 268.950 328.050 269.400 ;
        RECT 334.950 268.950 337.050 269.400 ;
        RECT 673.950 268.950 676.050 269.400 ;
        RECT 736.950 270.600 739.050 271.050 ;
        RECT 775.950 270.600 778.050 271.050 ;
        RECT 736.950 269.400 778.050 270.600 ;
        RECT 736.950 268.950 739.050 269.400 ;
        RECT 775.950 268.950 778.050 269.400 ;
        RECT 136.950 267.600 139.050 268.050 ;
        RECT 178.800 267.600 180.900 268.050 ;
        RECT 136.950 266.400 180.900 267.600 ;
        RECT 136.950 265.950 139.050 266.400 ;
        RECT 178.800 265.950 180.900 266.400 ;
        RECT 181.950 267.600 184.050 268.050 ;
        RECT 196.950 267.600 199.050 268.050 ;
        RECT 181.950 266.400 199.050 267.600 ;
        RECT 181.950 265.950 184.050 266.400 ;
        RECT 196.950 265.950 199.050 266.400 ;
        RECT 214.950 267.600 217.050 268.050 ;
        RECT 256.950 267.600 259.050 268.050 ;
        RECT 214.950 266.400 259.050 267.600 ;
        RECT 214.950 265.950 217.050 266.400 ;
        RECT 256.950 265.950 259.050 266.400 ;
        RECT 277.950 267.600 280.050 268.050 ;
        RECT 301.950 267.600 304.050 268.050 ;
        RECT 277.950 266.400 304.050 267.600 ;
        RECT 277.950 265.950 280.050 266.400 ;
        RECT 301.950 265.950 304.050 266.400 ;
        RECT 373.950 267.600 376.050 268.050 ;
        RECT 379.800 267.600 381.900 268.050 ;
        RECT 373.950 266.400 381.900 267.600 ;
        RECT 373.950 265.950 376.050 266.400 ;
        RECT 379.800 265.950 381.900 266.400 ;
        RECT 382.950 267.600 385.050 268.050 ;
        RECT 418.950 267.600 421.050 268.050 ;
        RECT 382.950 266.400 421.050 267.600 ;
        RECT 382.950 265.950 385.050 266.400 ;
        RECT 418.950 265.950 421.050 266.400 ;
        RECT 439.950 267.600 442.050 268.050 ;
        RECT 451.950 267.600 454.050 268.050 ;
        RECT 439.950 266.400 454.050 267.600 ;
        RECT 439.950 265.950 442.050 266.400 ;
        RECT 451.950 265.950 454.050 266.400 ;
        RECT 463.950 267.600 466.050 268.050 ;
        RECT 556.950 267.600 559.050 268.050 ;
        RECT 463.950 266.400 559.050 267.600 ;
        RECT 463.950 265.950 466.050 266.400 ;
        RECT 556.950 265.950 559.050 266.400 ;
        RECT 679.950 267.600 682.050 268.050 ;
        RECT 697.950 267.600 700.050 268.050 ;
        RECT 679.950 266.400 700.050 267.600 ;
        RECT 679.950 265.950 682.050 266.400 ;
        RECT 697.950 265.950 700.050 266.400 ;
        RECT 4.950 261.750 7.050 262.200 ;
        RECT 16.950 261.750 19.050 262.200 ;
        RECT 4.950 260.550 19.050 261.750 ;
        RECT 4.950 260.100 7.050 260.550 ;
        RECT 16.950 260.100 19.050 260.550 ;
        RECT 34.950 259.950 37.050 262.050 ;
        RECT 67.950 261.750 70.050 262.200 ;
        RECT 73.950 261.750 76.050 262.200 ;
        RECT 67.950 260.550 76.050 261.750 ;
        RECT 67.950 260.100 70.050 260.550 ;
        RECT 73.950 260.100 76.050 260.550 ;
        RECT 82.950 261.600 85.050 262.350 ;
        RECT 88.950 261.600 91.050 265.050 ;
        RECT 109.950 264.600 112.050 265.050 ;
        RECT 121.950 264.600 124.050 265.050 ;
        RECT 151.950 264.600 154.050 265.050 ;
        RECT 109.950 263.400 154.050 264.600 ;
        RECT 109.950 262.950 112.050 263.400 ;
        RECT 121.950 262.950 124.050 263.400 ;
        RECT 151.950 262.950 154.050 263.400 ;
        RECT 238.950 264.600 241.050 265.050 ;
        RECT 262.950 264.600 265.050 265.050 ;
        RECT 238.950 263.400 265.050 264.600 ;
        RECT 238.950 262.950 241.050 263.400 ;
        RECT 262.950 262.950 265.050 263.400 ;
        RECT 292.950 264.600 295.050 265.050 ;
        RECT 316.950 264.600 319.050 265.050 ;
        RECT 292.950 263.400 319.050 264.600 ;
        RECT 292.950 262.950 295.050 263.400 ;
        RECT 316.950 262.950 319.050 263.400 ;
        RECT 328.950 264.600 331.050 265.050 ;
        RECT 367.950 264.600 370.050 265.050 ;
        RECT 427.950 264.600 430.050 265.050 ;
        RECT 328.950 263.400 430.050 264.600 ;
        RECT 328.950 262.950 331.050 263.400 ;
        RECT 367.950 262.950 370.050 263.400 ;
        RECT 427.950 262.950 430.050 263.400 ;
        RECT 475.950 264.600 478.050 265.050 ;
        RECT 496.950 264.600 499.050 265.050 ;
        RECT 475.950 263.400 499.050 264.600 ;
        RECT 475.950 262.950 478.050 263.400 ;
        RECT 496.950 262.950 499.050 263.400 ;
        RECT 673.950 264.600 676.050 265.050 ;
        RECT 715.950 264.600 718.050 265.050 ;
        RECT 751.950 264.600 754.050 265.050 ;
        RECT 769.950 264.600 772.050 265.050 ;
        RECT 673.950 263.400 744.450 264.600 ;
        RECT 673.950 262.950 676.050 263.400 ;
        RECT 715.950 262.950 718.050 263.400 ;
        RECT 82.950 261.000 91.050 261.600 ;
        RECT 94.950 261.750 97.050 262.200 ;
        RECT 103.950 261.750 106.050 262.200 ;
        RECT 82.950 260.400 90.600 261.000 ;
        RECT 94.950 260.550 106.050 261.750 ;
        RECT 82.950 260.250 85.050 260.400 ;
        RECT 94.950 260.100 97.050 260.550 ;
        RECT 103.950 260.100 106.050 260.550 ;
        RECT 118.950 261.600 121.050 262.050 ;
        RECT 148.950 261.600 151.050 262.050 ;
        RECT 172.950 261.600 175.050 262.200 ;
        RECT 118.950 260.400 151.050 261.600 ;
        RECT 118.950 259.950 121.050 260.400 ;
        RECT 148.950 259.950 151.050 260.400 ;
        RECT 164.400 260.400 175.050 261.600 ;
        RECT 22.950 255.600 25.050 255.900 ;
        RECT 35.400 255.600 36.600 259.950 ;
        RECT 136.950 258.600 139.050 259.050 ;
        RECT 136.950 258.000 159.600 258.600 ;
        RECT 136.950 257.400 160.050 258.000 ;
        RECT 136.950 256.950 139.050 257.400 ;
        RECT 22.950 254.400 36.600 255.600 ;
        RECT 49.950 255.600 52.050 255.900 ;
        RECT 94.950 255.600 97.050 256.050 ;
        RECT 49.950 254.400 97.050 255.600 ;
        RECT 22.950 253.800 25.050 254.400 ;
        RECT 49.950 253.800 52.050 254.400 ;
        RECT 94.950 253.950 97.050 254.400 ;
        RECT 106.950 255.450 109.050 255.900 ;
        RECT 115.950 255.450 118.050 255.900 ;
        RECT 106.950 254.250 118.050 255.450 ;
        RECT 106.950 253.800 109.050 254.250 ;
        RECT 115.950 253.800 118.050 254.250 ;
        RECT 157.950 253.950 160.050 257.400 ;
        RECT 164.400 256.050 165.600 260.400 ;
        RECT 172.950 260.100 175.050 260.400 ;
        RECT 184.950 261.750 187.050 262.200 ;
        RECT 190.950 261.750 193.050 262.200 ;
        RECT 184.950 260.550 193.050 261.750 ;
        RECT 307.950 261.600 310.050 262.200 ;
        RECT 312.000 261.600 316.050 262.050 ;
        RECT 355.950 261.600 358.050 262.050 ;
        RECT 184.950 260.100 187.050 260.550 ;
        RECT 190.950 260.100 193.050 260.550 ;
        RECT 281.400 260.400 310.050 261.600 ;
        RECT 281.400 256.050 282.600 260.400 ;
        RECT 307.950 260.100 310.050 260.400 ;
        RECT 311.400 259.950 316.050 261.600 ;
        RECT 332.400 260.400 358.050 261.600 ;
        RECT 163.950 253.950 166.050 256.050 ;
        RECT 175.950 255.600 178.050 255.900 ;
        RECT 184.950 255.600 187.050 256.050 ;
        RECT 175.950 254.400 187.050 255.600 ;
        RECT 175.950 253.800 178.050 254.400 ;
        RECT 184.950 253.950 187.050 254.400 ;
        RECT 193.950 255.600 196.050 255.900 ;
        RECT 259.950 255.600 262.050 256.050 ;
        RECT 193.950 254.400 262.050 255.600 ;
        RECT 193.950 253.800 196.050 254.400 ;
        RECT 259.950 253.950 262.050 254.400 ;
        RECT 268.950 255.600 271.050 256.050 ;
        RECT 274.950 255.600 277.050 256.050 ;
        RECT 268.950 254.400 277.050 255.600 ;
        RECT 268.950 253.950 271.050 254.400 ;
        RECT 274.950 253.950 277.050 254.400 ;
        RECT 280.950 253.950 283.050 256.050 ;
        RECT 295.950 255.600 298.050 256.050 ;
        RECT 311.400 255.600 312.600 259.950 ;
        RECT 332.400 256.050 333.600 260.400 ;
        RECT 355.950 259.950 358.050 260.400 ;
        RECT 373.950 261.600 376.050 262.050 ;
        RECT 373.950 260.400 384.600 261.600 ;
        RECT 373.950 259.950 376.050 260.400 ;
        RECT 383.400 256.050 384.600 260.400 ;
        RECT 388.950 258.600 391.050 262.050 ;
        RECT 418.950 261.600 421.050 262.050 ;
        RECT 445.950 261.750 448.050 262.200 ;
        RECT 460.950 261.750 463.050 262.200 ;
        RECT 418.950 260.400 426.600 261.600 ;
        RECT 418.950 259.950 421.050 260.400 ;
        RECT 425.400 258.600 426.600 260.400 ;
        RECT 445.950 260.550 463.050 261.750 ;
        RECT 472.950 261.600 475.050 262.350 ;
        RECT 445.950 260.100 448.050 260.550 ;
        RECT 460.950 260.100 463.050 260.550 ;
        RECT 464.400 260.400 475.050 261.600 ;
        RECT 464.400 258.600 465.600 260.400 ;
        RECT 472.950 260.250 475.050 260.400 ;
        RECT 499.950 261.750 502.050 262.200 ;
        RECT 508.950 261.750 511.050 262.200 ;
        RECT 499.950 261.600 511.050 261.750 ;
        RECT 523.950 261.600 526.050 262.350 ;
        RECT 499.950 260.550 526.050 261.600 ;
        RECT 499.950 260.100 502.050 260.550 ;
        RECT 508.950 260.400 526.050 260.550 ;
        RECT 508.950 260.100 511.050 260.400 ;
        RECT 523.950 260.250 526.050 260.400 ;
        RECT 529.950 261.900 532.050 262.350 ;
        RECT 535.950 261.900 538.050 262.350 ;
        RECT 529.950 260.700 538.050 261.900 ;
        RECT 529.950 260.250 532.050 260.700 ;
        RECT 535.950 260.250 538.050 260.700 ;
        RECT 559.950 261.750 562.050 262.200 ;
        RECT 568.950 261.750 571.050 262.200 ;
        RECT 559.950 260.550 571.050 261.750 ;
        RECT 598.950 261.600 601.050 262.200 ;
        RECT 559.950 260.100 562.050 260.550 ;
        RECT 568.950 260.100 571.050 260.550 ;
        RECT 590.400 260.400 601.050 261.600 ;
        RECT 388.950 258.000 393.600 258.600 ;
        RECT 389.400 257.400 393.600 258.000 ;
        RECT 425.400 257.400 450.600 258.600 ;
        RECT 392.400 256.050 393.600 257.400 ;
        RECT 295.950 254.400 312.600 255.600 ;
        RECT 316.950 255.600 319.050 256.050 ;
        RECT 322.950 255.600 325.050 256.050 ;
        RECT 316.950 254.400 325.050 255.600 ;
        RECT 295.950 253.950 298.050 254.400 ;
        RECT 316.950 253.950 319.050 254.400 ;
        RECT 322.950 253.950 325.050 254.400 ;
        RECT 331.950 253.950 334.050 256.050 ;
        RECT 361.950 255.600 364.050 255.900 ;
        RECT 376.950 255.600 379.050 256.050 ;
        RECT 361.950 254.400 379.050 255.600 ;
        RECT 361.950 253.800 364.050 254.400 ;
        RECT 376.950 253.950 379.050 254.400 ;
        RECT 382.950 253.950 385.050 256.050 ;
        RECT 392.400 254.400 397.050 256.050 ;
        RECT 449.400 255.900 450.600 257.400 ;
        RECT 455.400 257.400 465.600 258.600 ;
        RECT 455.400 255.900 456.600 257.400 ;
        RECT 590.400 256.050 591.600 260.400 ;
        RECT 598.950 260.100 601.050 260.400 ;
        RECT 604.950 261.750 607.050 262.200 ;
        RECT 616.950 261.750 619.050 262.200 ;
        RECT 604.950 260.550 619.050 261.750 ;
        RECT 604.950 260.100 607.050 260.550 ;
        RECT 616.950 260.100 619.050 260.550 ;
        RECT 625.950 261.600 628.050 262.200 ;
        RECT 658.950 261.600 661.050 262.200 ;
        RECT 694.950 261.600 697.050 262.200 ;
        RECT 625.950 260.400 661.050 261.600 ;
        RECT 625.950 260.100 628.050 260.400 ;
        RECT 658.950 260.100 661.050 260.400 ;
        RECT 689.400 260.400 697.050 261.600 ;
        RECT 689.400 256.050 690.600 260.400 ;
        RECT 694.950 260.100 697.050 260.400 ;
        RECT 700.950 261.750 703.050 262.200 ;
        RECT 706.950 261.750 709.050 262.050 ;
        RECT 700.950 261.600 709.050 261.750 ;
        RECT 727.950 261.600 730.050 262.200 ;
        RECT 700.950 260.550 730.050 261.600 ;
        RECT 700.950 260.100 703.050 260.550 ;
        RECT 706.950 260.400 730.050 260.550 ;
        RECT 706.950 259.950 709.050 260.400 ;
        RECT 727.950 260.100 730.050 260.400 ;
        RECT 733.950 260.100 736.050 262.200 ;
        RECT 734.400 256.050 735.600 260.100 ;
        RECT 743.250 256.050 744.450 263.400 ;
        RECT 751.950 263.400 772.050 264.600 ;
        RECT 751.950 262.950 754.050 263.400 ;
        RECT 769.950 262.950 772.050 263.400 ;
        RECT 802.950 264.600 805.050 265.050 ;
        RECT 802.950 263.400 810.600 264.600 ;
        RECT 802.950 262.950 805.050 263.400 ;
        RECT 745.950 260.250 748.050 262.350 ;
        RECT 757.950 261.750 760.050 262.200 ;
        RECT 763.950 261.750 766.050 262.200 ;
        RECT 757.950 260.550 766.050 261.750 ;
        RECT 746.400 256.050 747.600 260.250 ;
        RECT 757.950 260.100 760.050 260.550 ;
        RECT 763.950 260.100 766.050 260.550 ;
        RECT 769.950 261.600 772.050 262.200 ;
        RECT 787.950 261.600 790.050 262.200 ;
        RECT 769.950 260.400 783.600 261.600 ;
        RECT 769.950 260.100 772.050 260.400 ;
        RECT 393.000 253.950 397.050 254.400 ;
        RECT 448.950 253.800 451.050 255.900 ;
        RECT 454.950 253.800 457.050 255.900 ;
        RECT 541.950 255.450 544.050 255.900 ;
        RECT 556.950 255.450 559.050 255.900 ;
        RECT 541.950 254.250 559.050 255.450 ;
        RECT 541.950 253.800 544.050 254.250 ;
        RECT 556.950 253.800 559.050 254.250 ;
        RECT 589.950 253.950 592.050 256.050 ;
        RECT 622.950 255.600 625.050 255.900 ;
        RECT 605.400 254.400 625.050 255.600 ;
        RECT 605.400 253.050 606.600 254.400 ;
        RECT 622.950 253.800 625.050 254.400 ;
        RECT 631.950 255.450 634.050 255.900 ;
        RECT 646.950 255.450 649.050 255.900 ;
        RECT 631.950 254.250 649.050 255.450 ;
        RECT 631.950 253.800 634.050 254.250 ;
        RECT 646.950 253.800 649.050 254.250 ;
        RECT 688.950 253.950 691.050 256.050 ;
        RECT 697.950 255.600 700.050 255.900 ;
        RECT 712.950 255.600 715.050 255.900 ;
        RECT 721.950 255.600 724.050 256.050 ;
        RECT 697.950 254.400 724.050 255.600 ;
        RECT 734.400 254.400 739.050 256.050 ;
        RECT 697.950 253.800 700.050 254.400 ;
        RECT 712.950 253.800 715.050 254.400 ;
        RECT 721.950 253.950 724.050 254.400 ;
        RECT 735.000 253.950 739.050 254.400 ;
        RECT 742.800 253.950 744.900 256.050 ;
        RECT 745.950 253.950 748.050 256.050 ;
        RECT 766.950 255.600 769.050 255.900 ;
        RECT 775.950 255.600 778.050 256.050 ;
        RECT 766.950 254.400 778.050 255.600 ;
        RECT 782.400 255.600 783.600 260.400 ;
        RECT 787.950 260.400 798.600 261.600 ;
        RECT 787.950 260.100 790.050 260.400 ;
        RECT 797.400 256.050 798.600 260.400 ;
        RECT 809.400 256.050 810.600 263.400 ;
        RECT 811.950 261.600 816.000 262.050 ;
        RECT 811.950 259.950 816.600 261.600 ;
        RECT 790.950 255.600 793.050 255.900 ;
        RECT 782.400 254.400 793.050 255.600 ;
        RECT 766.950 253.800 769.050 254.400 ;
        RECT 775.950 253.950 778.050 254.400 ;
        RECT 790.950 253.800 793.050 254.400 ;
        RECT 796.950 253.950 799.050 256.050 ;
        RECT 808.950 253.950 811.050 256.050 ;
        RECT 815.400 255.900 816.600 259.950 ;
        RECT 821.400 256.050 822.600 271.950 ;
        RECT 826.950 267.600 829.050 268.050 ;
        RECT 847.950 267.600 850.050 268.050 ;
        RECT 826.950 266.400 850.050 267.600 ;
        RECT 826.950 265.950 829.050 266.400 ;
        RECT 847.950 265.950 850.050 266.400 ;
        RECT 826.950 259.950 829.050 262.050 ;
        RECT 841.950 261.750 844.050 262.200 ;
        RECT 850.950 261.750 853.050 262.200 ;
        RECT 841.950 260.550 853.050 261.750 ;
        RECT 841.950 260.100 844.050 260.550 ;
        RECT 850.950 260.100 853.050 260.550 ;
        RECT 827.400 256.050 828.600 259.950 ;
        RECT 814.950 253.800 817.050 255.900 ;
        RECT 820.950 253.950 823.050 256.050 ;
        RECT 826.950 253.950 829.050 256.050 ;
        RECT 475.950 252.600 478.050 253.050 ;
        RECT 499.950 252.600 502.050 253.050 ;
        RECT 475.950 251.400 502.050 252.600 ;
        RECT 475.950 250.950 478.050 251.400 ;
        RECT 499.950 250.950 502.050 251.400 ;
        RECT 601.950 251.400 606.600 253.050 ;
        RECT 778.950 252.600 781.050 253.050 ;
        RECT 784.950 252.600 787.050 253.050 ;
        RECT 778.950 251.400 787.050 252.600 ;
        RECT 601.950 250.950 606.000 251.400 ;
        RECT 778.950 250.950 781.050 251.400 ;
        RECT 784.950 250.950 787.050 251.400 ;
        RECT 823.950 252.600 826.050 253.050 ;
        RECT 832.950 252.600 835.050 253.050 ;
        RECT 823.950 251.400 835.050 252.600 ;
        RECT 823.950 250.950 826.050 251.400 ;
        RECT 832.950 250.950 835.050 251.400 ;
        RECT 31.950 249.600 34.050 250.050 ;
        RECT 40.950 249.600 43.050 250.050 ;
        RECT 58.950 249.600 61.050 250.050 ;
        RECT 121.950 249.600 124.050 250.050 ;
        RECT 31.950 248.400 124.050 249.600 ;
        RECT 31.950 247.950 34.050 248.400 ;
        RECT 40.950 247.950 43.050 248.400 ;
        RECT 58.950 247.950 61.050 248.400 ;
        RECT 121.950 247.950 124.050 248.400 ;
        RECT 151.950 249.600 154.050 250.050 ;
        RECT 199.950 249.600 202.050 250.050 ;
        RECT 151.950 248.400 202.050 249.600 ;
        RECT 151.950 247.950 154.050 248.400 ;
        RECT 199.950 247.950 202.050 248.400 ;
        RECT 217.950 249.600 220.050 250.050 ;
        RECT 331.950 249.600 334.050 250.050 ;
        RECT 217.950 248.400 334.050 249.600 ;
        RECT 217.950 247.950 220.050 248.400 ;
        RECT 331.950 247.950 334.050 248.400 ;
        RECT 433.950 249.600 436.050 250.050 ;
        RECT 460.950 249.600 463.050 250.050 ;
        RECT 469.950 249.600 472.050 250.050 ;
        RECT 433.950 248.400 472.050 249.600 ;
        RECT 433.950 247.950 436.050 248.400 ;
        RECT 460.950 247.950 463.050 248.400 ;
        RECT 469.950 247.950 472.050 248.400 ;
        RECT 481.950 249.600 484.050 250.050 ;
        RECT 529.950 249.600 532.050 250.050 ;
        RECT 550.950 249.600 553.050 250.050 ;
        RECT 481.950 248.400 495.600 249.600 ;
        RECT 481.950 247.950 484.050 248.400 ;
        RECT 85.950 246.600 88.050 247.050 ;
        RECT 94.950 246.600 97.050 247.050 ;
        RECT 152.400 246.600 153.600 247.950 ;
        RECT 85.950 245.400 153.600 246.600 ;
        RECT 202.950 246.600 205.050 247.050 ;
        RECT 259.950 246.600 262.050 247.050 ;
        RECT 403.950 246.600 406.050 247.050 ;
        RECT 448.950 246.600 451.050 247.050 ;
        RECT 202.950 245.400 451.050 246.600 ;
        RECT 494.400 246.600 495.600 248.400 ;
        RECT 529.950 248.400 553.050 249.600 ;
        RECT 529.950 247.950 532.050 248.400 ;
        RECT 550.950 247.950 553.050 248.400 ;
        RECT 616.950 249.600 619.050 250.050 ;
        RECT 640.950 249.600 643.050 250.050 ;
        RECT 616.950 248.400 643.050 249.600 ;
        RECT 616.950 247.950 619.050 248.400 ;
        RECT 640.950 247.950 643.050 248.400 ;
        RECT 664.950 249.600 667.050 250.050 ;
        RECT 676.950 249.600 679.050 250.050 ;
        RECT 664.950 248.400 679.050 249.600 ;
        RECT 664.950 247.950 667.050 248.400 ;
        RECT 676.950 247.950 679.050 248.400 ;
        RECT 757.950 249.600 760.050 250.050 ;
        RECT 805.950 249.600 808.050 250.050 ;
        RECT 757.950 248.400 808.050 249.600 ;
        RECT 757.950 247.950 760.050 248.400 ;
        RECT 805.950 247.950 808.050 248.400 ;
        RECT 811.950 249.600 814.050 250.050 ;
        RECT 820.950 249.600 823.050 250.050 ;
        RECT 811.950 248.400 823.050 249.600 ;
        RECT 811.950 247.950 814.050 248.400 ;
        RECT 820.950 247.950 823.050 248.400 ;
        RECT 499.950 246.600 502.050 247.050 ;
        RECT 494.400 245.400 502.050 246.600 ;
        RECT 85.950 244.950 88.050 245.400 ;
        RECT 94.950 244.950 97.050 245.400 ;
        RECT 202.950 244.950 205.050 245.400 ;
        RECT 259.950 244.950 262.050 245.400 ;
        RECT 403.950 244.950 406.050 245.400 ;
        RECT 448.950 244.950 451.050 245.400 ;
        RECT 499.950 244.950 502.050 245.400 ;
        RECT 526.950 246.600 529.050 247.050 ;
        RECT 580.950 246.600 583.050 247.050 ;
        RECT 526.950 245.400 583.050 246.600 ;
        RECT 526.950 244.950 529.050 245.400 ;
        RECT 580.950 244.950 583.050 245.400 ;
        RECT 601.950 246.600 604.050 247.050 ;
        RECT 607.950 246.600 610.050 247.050 ;
        RECT 601.950 245.400 610.050 246.600 ;
        RECT 601.950 244.950 604.050 245.400 ;
        RECT 607.950 244.950 610.050 245.400 ;
        RECT 691.950 246.600 694.050 247.050 ;
        RECT 709.950 246.600 712.050 247.050 ;
        RECT 691.950 245.400 712.050 246.600 ;
        RECT 691.950 244.950 694.050 245.400 ;
        RECT 709.950 244.950 712.050 245.400 ;
        RECT 730.950 246.600 733.050 247.050 ;
        RECT 745.950 246.600 748.050 247.050 ;
        RECT 730.950 245.400 748.050 246.600 ;
        RECT 730.950 244.950 733.050 245.400 ;
        RECT 745.950 244.950 748.050 245.400 ;
        RECT 223.950 243.600 226.050 244.050 ;
        RECT 238.950 243.600 241.050 244.050 ;
        RECT 223.950 242.400 241.050 243.600 ;
        RECT 223.950 241.950 226.050 242.400 ;
        RECT 238.950 241.950 241.050 242.400 ;
        RECT 247.950 243.600 250.050 244.050 ;
        RECT 277.950 243.600 280.050 244.050 ;
        RECT 289.950 243.600 292.050 244.050 ;
        RECT 247.950 242.400 292.050 243.600 ;
        RECT 247.950 241.950 250.050 242.400 ;
        RECT 277.950 241.950 280.050 242.400 ;
        RECT 289.950 241.950 292.050 242.400 ;
        RECT 322.950 243.600 325.050 244.050 ;
        RECT 397.950 243.600 400.050 244.050 ;
        RECT 433.950 243.600 436.050 244.050 ;
        RECT 322.950 242.400 436.050 243.600 ;
        RECT 322.950 241.950 325.050 242.400 ;
        RECT 397.950 241.950 400.050 242.400 ;
        RECT 433.950 241.950 436.050 242.400 ;
        RECT 439.950 243.600 442.050 244.050 ;
        RECT 490.950 243.600 493.050 244.050 ;
        RECT 439.950 242.400 493.050 243.600 ;
        RECT 439.950 241.950 442.050 242.400 ;
        RECT 490.950 241.950 493.050 242.400 ;
        RECT 793.950 243.600 796.050 244.050 ;
        RECT 826.950 243.600 829.050 244.050 ;
        RECT 793.950 242.400 829.050 243.600 ;
        RECT 793.950 241.950 796.050 242.400 ;
        RECT 826.950 241.950 829.050 242.400 ;
        RECT 205.950 240.600 208.050 241.050 ;
        RECT 214.950 240.600 217.050 241.050 ;
        RECT 205.950 239.400 217.050 240.600 ;
        RECT 205.950 238.950 208.050 239.400 ;
        RECT 214.950 238.950 217.050 239.400 ;
        RECT 226.950 240.600 229.050 241.050 ;
        RECT 295.950 240.600 298.050 241.050 ;
        RECT 226.950 239.400 298.050 240.600 ;
        RECT 226.950 238.950 229.050 239.400 ;
        RECT 295.950 238.950 298.050 239.400 ;
        RECT 544.950 240.600 547.050 241.050 ;
        RECT 559.950 240.600 562.050 241.050 ;
        RECT 583.950 240.600 586.050 241.050 ;
        RECT 544.950 239.400 586.050 240.600 ;
        RECT 544.950 238.950 547.050 239.400 ;
        RECT 559.950 238.950 562.050 239.400 ;
        RECT 583.950 238.950 586.050 239.400 ;
        RECT 751.950 240.600 754.050 241.050 ;
        RECT 829.950 240.600 832.050 241.050 ;
        RECT 751.950 239.400 832.050 240.600 ;
        RECT 751.950 238.950 754.050 239.400 ;
        RECT 829.950 238.950 832.050 239.400 ;
        RECT 340.950 237.600 343.050 238.050 ;
        RECT 358.950 237.600 361.050 238.050 ;
        RECT 499.950 237.600 502.050 238.050 ;
        RECT 340.950 236.400 502.050 237.600 ;
        RECT 340.950 235.950 343.050 236.400 ;
        RECT 358.950 235.950 361.050 236.400 ;
        RECT 499.950 235.950 502.050 236.400 ;
        RECT 199.950 234.600 202.050 235.050 ;
        RECT 226.950 234.600 229.050 235.050 ;
        RECT 199.950 233.400 229.050 234.600 ;
        RECT 199.950 232.950 202.050 233.400 ;
        RECT 226.950 232.950 229.050 233.400 ;
        RECT 292.950 234.600 295.050 235.050 ;
        RECT 304.950 234.600 307.050 235.050 ;
        RECT 322.950 234.600 325.050 235.050 ;
        RECT 292.950 233.400 325.050 234.600 ;
        RECT 292.950 232.950 295.050 233.400 ;
        RECT 304.950 232.950 307.050 233.400 ;
        RECT 322.950 232.950 325.050 233.400 ;
        RECT 337.950 234.600 340.050 235.050 ;
        RECT 352.950 234.600 355.050 235.050 ;
        RECT 337.950 233.400 355.050 234.600 ;
        RECT 337.950 232.950 340.050 233.400 ;
        RECT 352.950 232.950 355.050 233.400 ;
        RECT 649.950 234.600 652.050 235.050 ;
        RECT 739.950 234.600 742.050 235.050 ;
        RECT 649.950 233.400 742.050 234.600 ;
        RECT 649.950 232.950 652.050 233.400 ;
        RECT 739.950 232.950 742.050 233.400 ;
        RECT 757.950 234.600 760.050 235.050 ;
        RECT 790.950 234.600 793.050 235.050 ;
        RECT 757.950 233.400 793.050 234.600 ;
        RECT 757.950 232.950 760.050 233.400 ;
        RECT 790.950 232.950 793.050 233.400 ;
        RECT 106.950 231.600 109.050 232.050 ;
        RECT 163.950 231.600 166.050 232.050 ;
        RECT 106.950 230.400 166.050 231.600 ;
        RECT 106.950 229.950 109.050 230.400 ;
        RECT 163.950 229.950 166.050 230.400 ;
        RECT 175.950 231.600 178.050 232.050 ;
        RECT 190.950 231.600 193.050 232.050 ;
        RECT 175.950 230.400 193.050 231.600 ;
        RECT 175.950 229.950 178.050 230.400 ;
        RECT 190.950 229.950 193.050 230.400 ;
        RECT 196.950 231.600 199.050 232.050 ;
        RECT 361.950 231.600 364.050 232.050 ;
        RECT 196.950 230.400 364.050 231.600 ;
        RECT 196.950 229.950 199.050 230.400 ;
        RECT 361.950 229.950 364.050 230.400 ;
        RECT 367.950 231.600 370.050 232.050 ;
        RECT 376.950 231.600 379.050 232.050 ;
        RECT 367.950 230.400 379.050 231.600 ;
        RECT 367.950 229.950 370.050 230.400 ;
        RECT 376.950 229.950 379.050 230.400 ;
        RECT 391.950 231.600 394.050 232.050 ;
        RECT 445.950 231.600 448.050 232.050 ;
        RECT 391.950 230.400 448.050 231.600 ;
        RECT 391.950 229.950 394.050 230.400 ;
        RECT 445.950 229.950 448.050 230.400 ;
        RECT 574.950 231.600 577.050 232.050 ;
        RECT 586.950 231.600 589.050 232.050 ;
        RECT 574.950 230.400 589.050 231.600 ;
        RECT 574.950 229.950 577.050 230.400 ;
        RECT 586.950 229.950 589.050 230.400 ;
        RECT 736.950 231.600 739.050 232.050 ;
        RECT 766.950 231.600 769.050 232.050 ;
        RECT 736.950 230.400 769.050 231.600 ;
        RECT 736.950 229.950 739.050 230.400 ;
        RECT 766.950 229.950 769.050 230.400 ;
        RECT 820.950 231.600 823.050 232.050 ;
        RECT 826.950 231.600 829.050 232.050 ;
        RECT 856.950 231.600 859.050 232.050 ;
        RECT 820.950 230.400 859.050 231.600 ;
        RECT 820.950 229.950 823.050 230.400 ;
        RECT 826.950 229.950 829.050 230.400 ;
        RECT 856.950 229.950 859.050 230.400 ;
        RECT 121.950 228.600 124.050 229.050 ;
        RECT 127.950 228.600 130.050 229.050 ;
        RECT 121.950 227.400 130.050 228.600 ;
        RECT 121.950 226.950 124.050 227.400 ;
        RECT 127.950 226.950 130.050 227.400 ;
        RECT 271.950 228.600 274.050 229.050 ;
        RECT 301.950 228.600 304.050 229.050 ;
        RECT 271.950 227.400 304.050 228.600 ;
        RECT 271.950 226.950 274.050 227.400 ;
        RECT 301.950 226.950 304.050 227.400 ;
        RECT 322.950 228.600 325.050 229.050 ;
        RECT 343.950 228.600 346.050 229.050 ;
        RECT 322.950 227.400 346.050 228.600 ;
        RECT 322.950 226.950 325.050 227.400 ;
        RECT 343.950 226.950 346.050 227.400 ;
        RECT 472.950 228.600 475.050 229.050 ;
        RECT 496.950 228.600 499.050 229.050 ;
        RECT 532.950 228.600 535.050 229.050 ;
        RECT 472.950 227.400 535.050 228.600 ;
        RECT 472.950 226.950 475.050 227.400 ;
        RECT 496.950 226.950 499.050 227.400 ;
        RECT 532.950 226.950 535.050 227.400 ;
        RECT 613.950 228.600 616.050 229.050 ;
        RECT 637.950 228.600 640.050 229.050 ;
        RECT 613.950 227.400 640.050 228.600 ;
        RECT 613.950 226.950 616.050 227.400 ;
        RECT 637.950 226.950 640.050 227.400 ;
        RECT 67.950 225.600 70.050 226.050 ;
        RECT 190.950 225.600 193.050 226.050 ;
        RECT 67.950 224.400 193.050 225.600 ;
        RECT 67.950 223.950 70.050 224.400 ;
        RECT 190.950 223.950 193.050 224.400 ;
        RECT 316.950 225.600 319.050 226.050 ;
        RECT 334.950 225.600 337.050 226.050 ;
        RECT 316.950 224.400 337.050 225.600 ;
        RECT 316.950 223.950 319.050 224.400 ;
        RECT 334.950 223.950 337.050 224.400 ;
        RECT 355.950 225.600 358.050 226.050 ;
        RECT 391.950 225.600 394.050 226.050 ;
        RECT 355.950 224.400 394.050 225.600 ;
        RECT 355.950 223.950 358.050 224.400 ;
        RECT 391.950 223.950 394.050 224.400 ;
        RECT 418.950 225.600 421.050 226.050 ;
        RECT 514.950 225.600 517.050 226.050 ;
        RECT 418.950 224.400 517.050 225.600 ;
        RECT 418.950 223.950 421.050 224.400 ;
        RECT 514.950 223.950 517.050 224.400 ;
        RECT 556.950 225.600 559.050 226.050 ;
        RECT 610.950 225.600 613.050 226.050 ;
        RECT 556.950 224.400 613.050 225.600 ;
        RECT 556.950 223.950 559.050 224.400 ;
        RECT 610.950 223.950 613.050 224.400 ;
        RECT 667.950 225.600 670.050 226.050 ;
        RECT 751.950 225.600 754.050 226.050 ;
        RECT 667.950 224.400 754.050 225.600 ;
        RECT 667.950 223.950 670.050 224.400 ;
        RECT 751.950 223.950 754.050 224.400 ;
        RECT 790.950 225.600 793.050 226.050 ;
        RECT 796.950 225.600 799.050 226.050 ;
        RECT 790.950 224.400 799.050 225.600 ;
        RECT 790.950 223.950 793.050 224.400 ;
        RECT 796.950 223.950 799.050 224.400 ;
        RECT 814.950 225.600 817.050 226.050 ;
        RECT 850.950 225.600 853.050 226.050 ;
        RECT 814.950 224.400 853.050 225.600 ;
        RECT 814.950 223.950 817.050 224.400 ;
        RECT 850.950 223.950 853.050 224.400 ;
        RECT 121.950 222.600 124.050 223.050 ;
        RECT 145.950 222.600 148.050 223.050 ;
        RECT 121.950 221.400 148.050 222.600 ;
        RECT 121.950 220.950 124.050 221.400 ;
        RECT 145.950 220.950 148.050 221.400 ;
        RECT 232.950 222.600 235.050 223.050 ;
        RECT 241.950 222.600 244.050 223.050 ;
        RECT 232.950 221.400 244.050 222.600 ;
        RECT 232.950 220.950 235.050 221.400 ;
        RECT 241.950 220.950 244.050 221.400 ;
        RECT 298.950 222.600 301.050 223.050 ;
        RECT 343.950 222.600 346.050 223.050 ;
        RECT 298.950 221.400 346.050 222.600 ;
        RECT 298.950 220.950 301.050 221.400 ;
        RECT 343.950 220.950 346.050 221.400 ;
        RECT 406.950 222.600 409.050 223.050 ;
        RECT 424.950 222.600 427.050 223.050 ;
        RECT 406.950 221.400 427.050 222.600 ;
        RECT 406.950 220.950 409.050 221.400 ;
        RECT 424.950 220.950 427.050 221.400 ;
        RECT 193.950 219.600 196.050 220.050 ;
        RECT 211.950 219.600 214.050 220.050 ;
        RECT 340.950 219.600 343.050 220.050 ;
        RECT 193.950 218.400 214.050 219.600 ;
        RECT 193.950 217.950 196.050 218.400 ;
        RECT 211.950 217.950 214.050 218.400 ;
        RECT 329.400 218.400 343.050 219.600 ;
        RECT 22.950 216.600 25.050 217.200 ;
        RECT 46.950 216.600 49.050 217.050 ;
        RECT 22.950 215.400 49.050 216.600 ;
        RECT 22.950 215.100 25.050 215.400 ;
        RECT 46.950 214.950 49.050 215.400 ;
        RECT 85.950 216.600 88.050 217.200 ;
        RECT 105.000 216.600 109.050 217.050 ;
        RECT 139.950 216.600 142.050 217.200 ;
        RECT 190.950 216.600 193.050 217.200 ;
        RECT 85.950 215.400 90.600 216.600 ;
        RECT 85.950 215.100 88.050 215.400 ;
        RECT 89.400 211.050 90.600 215.400 ;
        RECT 104.400 214.950 109.050 216.600 ;
        RECT 119.400 215.400 142.050 216.600 ;
        RECT 70.950 210.600 73.050 210.900 ;
        RECT 76.950 210.600 79.050 211.050 ;
        RECT 82.950 210.600 85.050 210.900 ;
        RECT 70.950 209.400 85.050 210.600 ;
        RECT 70.950 208.800 73.050 209.400 ;
        RECT 76.950 208.950 79.050 209.400 ;
        RECT 82.950 208.800 85.050 209.400 ;
        RECT 88.950 208.950 91.050 211.050 ;
        RECT 104.400 210.900 105.600 214.950 ;
        RECT 119.400 210.900 120.600 215.400 ;
        RECT 139.950 215.100 142.050 215.400 ;
        RECT 179.400 215.400 193.050 216.600 ;
        RECT 179.400 210.900 180.600 215.400 ;
        RECT 190.950 215.100 193.050 215.400 ;
        RECT 235.950 216.600 238.050 217.050 ;
        RECT 250.950 216.600 253.050 217.200 ;
        RECT 235.950 215.400 253.050 216.600 ;
        RECT 235.950 214.950 238.050 215.400 ;
        RECT 250.950 215.100 253.050 215.400 ;
        RECT 310.950 215.100 313.050 217.200 ;
        RECT 321.000 216.600 324.900 217.050 ;
        RECT 251.400 211.050 252.600 215.100 ;
        RECT 103.950 208.800 106.050 210.900 ;
        RECT 118.950 208.800 121.050 210.900 ;
        RECT 178.950 208.800 181.050 210.900 ;
        RECT 251.400 209.400 256.050 211.050 ;
        RECT 252.000 208.950 256.050 209.400 ;
        RECT 295.950 210.600 298.050 210.750 ;
        RECT 311.400 210.600 312.600 215.100 ;
        RECT 320.400 214.950 324.900 216.600 ;
        RECT 325.950 216.600 328.050 217.200 ;
        RECT 329.400 216.600 330.600 218.400 ;
        RECT 340.950 217.950 343.050 218.400 ;
        RECT 370.950 219.600 373.050 220.050 ;
        RECT 379.950 219.600 382.050 220.050 ;
        RECT 370.950 218.400 382.050 219.600 ;
        RECT 370.950 217.950 373.050 218.400 ;
        RECT 379.950 217.950 382.050 218.400 ;
        RECT 354.000 216.600 358.050 217.050 ;
        RECT 325.950 215.400 330.600 216.600 ;
        RECT 325.950 215.100 328.050 215.400 ;
        RECT 353.400 214.950 358.050 216.600 ;
        RECT 373.950 214.950 376.050 217.050 ;
        RECT 409.950 216.600 412.050 220.050 ;
        RECT 568.950 219.600 571.050 220.050 ;
        RECT 622.950 219.600 625.050 220.050 ;
        RECT 568.950 218.400 625.050 219.600 ;
        RECT 568.950 217.950 571.050 218.400 ;
        RECT 622.950 217.950 625.050 218.400 ;
        RECT 706.950 219.600 709.050 220.050 ;
        RECT 832.950 219.600 835.050 220.050 ;
        RECT 847.950 219.600 850.050 220.050 ;
        RECT 706.950 218.400 717.600 219.600 ;
        RECT 706.950 217.950 709.050 218.400 ;
        RECT 418.950 216.600 421.050 217.050 ;
        RECT 454.950 216.600 457.050 217.200 ;
        RECT 407.400 216.000 412.050 216.600 ;
        RECT 407.400 215.400 411.600 216.000 ;
        RECT 413.400 215.400 421.050 216.600 ;
        RECT 320.400 210.900 321.600 214.950 ;
        RECT 353.400 210.900 354.600 214.950 ;
        RECT 374.400 211.050 375.600 214.950 ;
        RECT 407.400 213.600 408.600 215.400 ;
        RECT 413.400 213.600 414.600 215.400 ;
        RECT 418.950 214.950 421.050 215.400 ;
        RECT 437.400 215.400 457.050 216.600 ;
        RECT 404.400 212.400 408.600 213.600 ;
        RECT 410.400 212.400 414.600 213.600 ;
        RECT 295.950 209.400 312.600 210.600 ;
        RECT 295.950 208.650 298.050 209.400 ;
        RECT 319.950 208.800 322.050 210.900 ;
        RECT 352.950 208.800 355.050 210.900 ;
        RECT 373.950 208.950 376.050 211.050 ;
        RECT 404.400 210.900 405.600 212.400 ;
        RECT 410.400 210.900 411.600 212.400 ;
        RECT 388.950 210.450 391.050 210.900 ;
        RECT 397.950 210.450 400.050 210.900 ;
        RECT 388.950 209.250 400.050 210.450 ;
        RECT 388.950 208.800 391.050 209.250 ;
        RECT 397.950 208.800 400.050 209.250 ;
        RECT 403.950 208.800 406.050 210.900 ;
        RECT 409.950 208.800 412.050 210.900 ;
        RECT 427.950 210.600 430.050 210.750 ;
        RECT 437.400 210.600 438.600 215.400 ;
        RECT 454.950 215.100 457.050 215.400 ;
        RECT 490.950 216.600 493.050 217.050 ;
        RECT 499.950 216.600 502.050 217.050 ;
        RECT 490.950 215.400 502.050 216.600 ;
        RECT 490.950 214.950 493.050 215.400 ;
        RECT 499.950 214.950 502.050 215.400 ;
        RECT 505.950 216.600 508.050 217.050 ;
        RECT 511.950 216.600 514.050 217.050 ;
        RECT 505.950 215.400 514.050 216.600 ;
        RECT 505.950 214.950 508.050 215.400 ;
        RECT 511.950 214.950 514.050 215.400 ;
        RECT 517.950 216.600 520.050 217.050 ;
        RECT 538.950 216.600 541.050 217.200 ;
        RECT 517.950 215.400 541.050 216.600 ;
        RECT 517.950 214.950 520.050 215.400 ;
        RECT 538.950 215.100 541.050 215.400 ;
        RECT 544.950 214.950 547.050 217.050 ;
        RECT 550.950 214.950 553.050 217.050 ;
        RECT 559.950 216.750 562.050 217.200 ;
        RECT 568.950 216.750 571.050 217.200 ;
        RECT 559.950 215.550 571.050 216.750 ;
        RECT 559.950 215.100 562.050 215.550 ;
        RECT 568.950 215.100 571.050 215.550 ;
        RECT 577.950 215.100 580.050 217.200 ;
        RECT 631.950 215.100 634.050 217.200 ;
        RECT 660.000 216.600 664.050 217.050 ;
        RECT 682.950 216.600 685.050 217.200 ;
        RECT 427.950 209.400 438.600 210.600 ;
        RECT 520.950 210.600 523.050 210.750 ;
        RECT 529.950 210.600 532.050 211.050 ;
        RECT 520.950 209.400 532.050 210.600 ;
        RECT 427.950 208.650 430.050 209.400 ;
        RECT 520.950 208.650 523.050 209.400 ;
        RECT 529.950 208.950 532.050 209.400 ;
        RECT 541.950 210.600 544.050 210.900 ;
        RECT 545.400 210.600 546.600 214.950 ;
        RECT 551.400 211.050 552.600 214.950 ;
        RECT 541.950 209.400 546.600 210.600 ;
        RECT 547.950 209.400 552.600 211.050 ;
        RECT 559.950 210.600 562.050 210.750 ;
        RECT 578.400 210.600 579.600 215.100 ;
        RECT 632.400 211.050 633.600 215.100 ;
        RECT 659.400 214.950 664.050 216.600 ;
        RECT 674.400 215.400 685.050 216.600 ;
        RECT 659.400 211.050 660.600 214.950 ;
        RECT 674.400 213.600 675.600 215.400 ;
        RECT 682.950 215.100 685.050 215.400 ;
        RECT 697.950 216.600 700.050 217.050 ;
        RECT 703.950 216.600 706.050 217.050 ;
        RECT 697.950 215.400 706.050 216.600 ;
        RECT 697.950 214.950 700.050 215.400 ;
        RECT 703.950 214.950 706.050 215.400 ;
        RECT 709.950 213.600 712.050 217.050 ;
        RECT 665.400 212.400 675.600 213.600 ;
        RECT 704.400 213.000 712.050 213.600 ;
        RECT 704.400 212.400 711.600 213.000 ;
        RECT 559.950 209.400 579.600 210.600 ;
        RECT 595.950 210.600 598.050 210.900 ;
        RECT 607.950 210.600 610.050 210.900 ;
        RECT 595.950 209.400 610.050 210.600 ;
        RECT 632.400 209.400 637.050 211.050 ;
        RECT 541.950 208.800 544.050 209.400 ;
        RECT 547.950 208.950 552.000 209.400 ;
        RECT 559.950 208.650 562.050 209.400 ;
        RECT 595.950 208.800 598.050 209.400 ;
        RECT 607.950 208.800 610.050 209.400 ;
        RECT 633.000 208.950 637.050 209.400 ;
        RECT 658.950 208.950 661.050 211.050 ;
        RECT 665.400 210.750 666.600 212.400 ;
        RECT 664.950 208.650 667.050 210.750 ;
        RECT 670.950 210.600 673.050 211.050 ;
        RECT 676.950 210.600 679.050 211.050 ;
        RECT 670.950 209.400 679.050 210.600 ;
        RECT 670.950 208.950 673.050 209.400 ;
        RECT 676.950 208.950 679.050 209.400 ;
        RECT 694.950 210.600 697.050 211.050 ;
        RECT 704.400 210.600 705.600 212.400 ;
        RECT 694.950 209.400 705.600 210.600 ;
        RECT 706.950 210.600 709.050 210.750 ;
        RECT 716.400 210.600 717.600 218.400 ;
        RECT 832.950 218.400 850.050 219.600 ;
        RECT 832.950 217.950 835.050 218.400 ;
        RECT 847.950 217.950 850.050 218.400 ;
        RECT 781.950 216.600 784.050 217.200 ;
        RECT 799.950 216.600 802.050 217.200 ;
        RECT 770.400 215.400 784.050 216.600 ;
        RECT 770.400 210.900 771.600 215.400 ;
        RECT 781.950 215.100 784.050 215.400 ;
        RECT 785.400 215.400 802.050 216.600 ;
        RECT 785.400 210.900 786.600 215.400 ;
        RECT 799.950 215.100 802.050 215.400 ;
        RECT 811.950 214.950 814.050 217.050 ;
        RECT 838.950 216.750 841.050 217.200 ;
        RECT 856.950 216.750 859.050 217.200 ;
        RECT 838.950 215.550 859.050 216.750 ;
        RECT 838.950 215.100 841.050 215.550 ;
        RECT 856.950 215.100 859.050 215.550 ;
        RECT 706.950 209.400 717.600 210.600 ;
        RECT 739.950 210.450 742.050 210.900 ;
        RECT 745.950 210.450 748.050 210.900 ;
        RECT 694.950 208.950 697.050 209.400 ;
        RECT 706.950 208.650 709.050 209.400 ;
        RECT 739.950 209.250 748.050 210.450 ;
        RECT 739.950 208.800 742.050 209.250 ;
        RECT 745.950 208.800 748.050 209.250 ;
        RECT 769.950 208.800 772.050 210.900 ;
        RECT 784.950 208.800 787.050 210.900 ;
        RECT 802.950 210.600 805.050 210.900 ;
        RECT 812.400 210.600 813.600 214.950 ;
        RECT 817.950 210.600 820.050 210.750 ;
        RECT 802.950 209.400 820.050 210.600 ;
        RECT 802.950 208.800 805.050 209.400 ;
        RECT 817.950 208.650 820.050 209.400 ;
        RECT 841.950 210.450 844.050 210.900 ;
        RECT 853.950 210.450 856.050 210.900 ;
        RECT 841.950 209.250 856.050 210.450 ;
        RECT 841.950 208.800 844.050 209.250 ;
        RECT 853.950 208.800 856.050 209.250 ;
        RECT 49.950 207.600 52.050 208.050 ;
        RECT 61.950 207.600 64.050 208.050 ;
        RECT 49.950 206.400 64.050 207.600 ;
        RECT 49.950 205.950 52.050 206.400 ;
        RECT 61.950 205.950 64.050 206.400 ;
        RECT 223.950 207.600 226.050 208.050 ;
        RECT 256.950 207.600 259.050 208.050 ;
        RECT 292.950 207.600 295.050 208.050 ;
        RECT 223.950 206.400 295.050 207.600 ;
        RECT 223.950 205.950 226.050 206.400 ;
        RECT 256.950 205.950 259.050 206.400 ;
        RECT 292.950 205.950 295.050 206.400 ;
        RECT 499.950 207.600 502.050 208.050 ;
        RECT 514.950 207.600 517.050 208.050 ;
        RECT 535.950 207.600 538.050 208.050 ;
        RECT 553.950 207.600 556.050 208.050 ;
        RECT 499.950 206.400 556.050 207.600 ;
        RECT 499.950 205.950 502.050 206.400 ;
        RECT 514.950 205.950 517.050 206.400 ;
        RECT 535.950 205.950 538.050 206.400 ;
        RECT 553.950 205.950 556.050 206.400 ;
        RECT 649.950 207.600 652.050 208.050 ;
        RECT 655.950 207.600 658.050 208.050 ;
        RECT 649.950 206.400 658.050 207.600 ;
        RECT 649.950 205.950 652.050 206.400 ;
        RECT 655.950 205.950 658.050 206.400 ;
        RECT 679.950 207.600 682.050 208.050 ;
        RECT 691.950 207.600 694.050 208.050 ;
        RECT 679.950 206.400 694.050 207.600 ;
        RECT 679.950 205.950 682.050 206.400 ;
        RECT 691.950 205.950 694.050 206.400 ;
        RECT 403.950 204.600 406.050 205.050 ;
        RECT 433.950 204.600 436.050 205.050 ;
        RECT 403.950 203.400 436.050 204.600 ;
        RECT 403.950 202.950 406.050 203.400 ;
        RECT 433.950 202.950 436.050 203.400 ;
        RECT 607.950 204.600 610.050 205.050 ;
        RECT 697.950 204.600 700.050 205.050 ;
        RECT 607.950 203.400 700.050 204.600 ;
        RECT 607.950 202.950 610.050 203.400 ;
        RECT 697.950 202.950 700.050 203.400 ;
        RECT 778.950 204.600 781.050 205.050 ;
        RECT 808.950 204.600 811.050 205.050 ;
        RECT 778.950 203.400 811.050 204.600 ;
        RECT 778.950 202.950 781.050 203.400 ;
        RECT 808.950 202.950 811.050 203.400 ;
        RECT 91.950 201.600 94.050 202.050 ;
        RECT 112.950 201.600 115.050 202.050 ;
        RECT 307.950 201.600 310.050 202.050 ;
        RECT 340.950 201.600 343.050 202.050 ;
        RECT 91.950 200.400 132.600 201.600 ;
        RECT 91.950 199.950 94.050 200.400 ;
        RECT 112.950 199.950 115.050 200.400 ;
        RECT 7.950 198.600 10.050 199.050 ;
        RECT 16.950 198.600 19.050 199.050 ;
        RECT 7.950 197.400 19.050 198.600 ;
        RECT 131.400 198.600 132.600 200.400 ;
        RECT 307.950 200.400 343.050 201.600 ;
        RECT 307.950 199.950 310.050 200.400 ;
        RECT 340.950 199.950 343.050 200.400 ;
        RECT 355.950 201.600 358.050 202.050 ;
        RECT 379.950 201.600 382.050 202.050 ;
        RECT 355.950 200.400 382.050 201.600 ;
        RECT 355.950 199.950 358.050 200.400 ;
        RECT 379.950 199.950 382.050 200.400 ;
        RECT 421.950 201.600 424.050 202.050 ;
        RECT 430.950 201.600 433.050 202.050 ;
        RECT 505.950 201.600 508.050 202.050 ;
        RECT 421.950 200.400 508.050 201.600 ;
        RECT 421.950 199.950 424.050 200.400 ;
        RECT 430.950 199.950 433.050 200.400 ;
        RECT 505.950 199.950 508.050 200.400 ;
        RECT 553.950 201.600 556.050 202.050 ;
        RECT 559.950 201.600 562.050 202.050 ;
        RECT 553.950 200.400 562.050 201.600 ;
        RECT 553.950 199.950 556.050 200.400 ;
        RECT 559.950 199.950 562.050 200.400 ;
        RECT 604.950 201.600 607.050 202.050 ;
        RECT 637.950 201.600 640.050 202.050 ;
        RECT 604.950 200.400 640.050 201.600 ;
        RECT 604.950 199.950 607.050 200.400 ;
        RECT 637.950 199.950 640.050 200.400 ;
        RECT 181.950 198.600 184.050 199.050 ;
        RECT 131.400 197.400 184.050 198.600 ;
        RECT 7.950 196.950 10.050 197.400 ;
        RECT 16.950 196.950 19.050 197.400 ;
        RECT 181.950 196.950 184.050 197.400 ;
        RECT 373.950 198.600 376.050 199.050 ;
        RECT 382.950 198.600 385.050 199.050 ;
        RECT 373.950 197.400 385.050 198.600 ;
        RECT 373.950 196.950 376.050 197.400 ;
        RECT 382.950 196.950 385.050 197.400 ;
        RECT 589.950 198.600 592.050 199.050 ;
        RECT 763.950 198.600 766.050 199.050 ;
        RECT 589.950 197.400 766.050 198.600 ;
        RECT 589.950 196.950 592.050 197.400 ;
        RECT 763.950 196.950 766.050 197.400 ;
        RECT 793.950 198.600 796.050 199.050 ;
        RECT 814.950 198.600 817.050 199.050 ;
        RECT 793.950 197.400 817.050 198.600 ;
        RECT 793.950 196.950 796.050 197.400 ;
        RECT 814.950 196.950 817.050 197.400 ;
        RECT 127.950 195.600 130.050 196.050 ;
        RECT 214.950 195.600 217.050 196.050 ;
        RECT 127.950 194.400 217.050 195.600 ;
        RECT 127.950 193.950 130.050 194.400 ;
        RECT 214.950 193.950 217.050 194.400 ;
        RECT 232.950 195.600 235.050 196.050 ;
        RECT 325.950 195.600 328.050 196.050 ;
        RECT 232.950 194.400 328.050 195.600 ;
        RECT 232.950 193.950 235.050 194.400 ;
        RECT 325.950 193.950 328.050 194.400 ;
        RECT 343.950 195.600 346.050 196.050 ;
        RECT 352.950 195.600 355.050 196.050 ;
        RECT 421.950 195.600 424.050 196.050 ;
        RECT 343.950 194.400 355.050 195.600 ;
        RECT 343.950 193.950 346.050 194.400 ;
        RECT 352.950 193.950 355.050 194.400 ;
        RECT 356.400 194.400 424.050 195.600 ;
        RECT 13.950 192.600 16.050 193.050 ;
        RECT 28.950 192.600 31.050 193.050 ;
        RECT 13.950 191.400 31.050 192.600 ;
        RECT 13.950 190.950 16.050 191.400 ;
        RECT 28.950 190.950 31.050 191.400 ;
        RECT 88.950 192.600 91.050 193.050 ;
        RECT 124.950 192.600 127.050 193.050 ;
        RECT 139.950 192.600 142.050 193.050 ;
        RECT 88.950 191.400 142.050 192.600 ;
        RECT 88.950 190.950 91.050 191.400 ;
        RECT 124.950 190.950 127.050 191.400 ;
        RECT 139.950 190.950 142.050 191.400 ;
        RECT 148.950 192.600 151.050 193.050 ;
        RECT 160.950 192.600 163.050 193.050 ;
        RECT 148.950 191.400 163.050 192.600 ;
        RECT 148.950 190.950 151.050 191.400 ;
        RECT 160.950 190.950 163.050 191.400 ;
        RECT 184.950 192.600 187.050 193.050 ;
        RECT 205.950 192.600 208.050 193.050 ;
        RECT 184.950 191.400 208.050 192.600 ;
        RECT 184.950 190.950 187.050 191.400 ;
        RECT 205.950 190.950 208.050 191.400 ;
        RECT 235.950 192.600 238.050 193.050 ;
        RECT 277.950 192.600 280.050 193.050 ;
        RECT 304.950 192.600 307.050 193.050 ;
        RECT 235.950 191.400 307.050 192.600 ;
        RECT 235.950 190.950 238.050 191.400 ;
        RECT 277.950 190.950 280.050 191.400 ;
        RECT 304.950 190.950 307.050 191.400 ;
        RECT 331.950 192.600 334.050 193.050 ;
        RECT 356.400 192.600 357.600 194.400 ;
        RECT 421.950 193.950 424.050 194.400 ;
        RECT 676.950 195.600 679.050 196.050 ;
        RECT 685.950 195.600 688.050 196.050 ;
        RECT 676.950 194.400 688.050 195.600 ;
        RECT 676.950 193.950 679.050 194.400 ;
        RECT 685.950 193.950 688.050 194.400 ;
        RECT 826.950 195.600 829.050 196.050 ;
        RECT 838.950 195.600 841.050 196.050 ;
        RECT 826.950 194.400 841.050 195.600 ;
        RECT 826.950 193.950 829.050 194.400 ;
        RECT 838.950 193.950 841.050 194.400 ;
        RECT 331.950 191.400 357.600 192.600 ;
        RECT 544.950 192.600 547.050 193.050 ;
        RECT 553.950 192.600 556.050 193.050 ;
        RECT 568.950 192.600 571.050 193.050 ;
        RECT 544.950 191.400 571.050 192.600 ;
        RECT 331.950 190.950 334.050 191.400 ;
        RECT 544.950 190.950 547.050 191.400 ;
        RECT 553.950 190.950 556.050 191.400 ;
        RECT 568.950 190.950 571.050 191.400 ;
        RECT 577.950 192.600 580.050 193.050 ;
        RECT 613.950 192.600 616.050 193.050 ;
        RECT 628.950 192.600 631.050 193.050 ;
        RECT 577.950 191.400 631.050 192.600 ;
        RECT 577.950 190.950 580.050 191.400 ;
        RECT 613.950 190.950 616.050 191.400 ;
        RECT 628.950 190.950 631.050 191.400 ;
        RECT 697.950 192.600 700.050 193.050 ;
        RECT 706.950 192.600 709.050 193.050 ;
        RECT 697.950 191.400 709.050 192.600 ;
        RECT 697.950 190.950 700.050 191.400 ;
        RECT 706.950 190.950 709.050 191.400 ;
        RECT 238.950 189.600 241.050 190.050 ;
        RECT 283.950 189.600 286.050 190.050 ;
        RECT 20.400 189.000 66.600 189.600 ;
        RECT 19.950 188.400 66.600 189.000 ;
        RECT 19.950 184.950 22.050 188.400 ;
        RECT 65.400 187.050 66.600 188.400 ;
        RECT 238.950 188.400 286.050 189.600 ;
        RECT 238.950 187.950 241.050 188.400 ;
        RECT 283.950 187.950 286.050 188.400 ;
        RECT 370.950 189.600 373.050 190.050 ;
        RECT 376.950 189.600 379.050 190.050 ;
        RECT 370.950 188.400 379.050 189.600 ;
        RECT 370.950 187.950 373.050 188.400 ;
        RECT 376.950 187.950 379.050 188.400 ;
        RECT 394.950 189.600 397.050 190.050 ;
        RECT 730.950 189.600 733.050 190.050 ;
        RECT 745.950 189.600 748.050 190.050 ;
        RECT 394.950 188.400 429.600 189.600 ;
        RECT 394.950 187.950 397.050 188.400 ;
        RECT 64.950 186.600 67.050 187.050 ;
        RECT 76.950 186.600 79.050 187.050 ;
        RECT 64.950 185.400 79.050 186.600 ;
        RECT 64.950 184.950 67.050 185.400 ;
        RECT 76.950 184.950 79.050 185.400 ;
        RECT 85.950 186.600 88.050 187.050 ;
        RECT 94.950 186.600 97.050 187.050 ;
        RECT 85.950 185.400 97.050 186.600 ;
        RECT 85.950 184.950 88.050 185.400 ;
        RECT 94.950 184.950 97.050 185.400 ;
        RECT 106.950 186.600 109.050 187.050 ;
        RECT 112.950 186.600 115.050 187.050 ;
        RECT 133.950 186.600 136.050 187.050 ;
        RECT 106.950 185.400 136.050 186.600 ;
        RECT 106.950 184.950 109.050 185.400 ;
        RECT 112.950 184.950 115.050 185.400 ;
        RECT 133.950 184.950 136.050 185.400 ;
        RECT 148.950 186.600 151.050 187.050 ;
        RECT 172.950 186.600 175.050 187.050 ;
        RECT 187.950 186.600 190.050 187.050 ;
        RECT 148.950 185.400 190.050 186.600 ;
        RECT 148.950 184.950 151.050 185.400 ;
        RECT 172.950 184.950 175.050 185.400 ;
        RECT 187.950 184.950 190.050 185.400 ;
        RECT 196.950 186.600 199.050 187.050 ;
        RECT 202.950 186.600 205.050 187.050 ;
        RECT 196.950 185.400 205.050 186.600 ;
        RECT 196.950 184.950 199.050 185.400 ;
        RECT 202.950 184.950 205.050 185.400 ;
        RECT 208.950 186.600 211.050 187.050 ;
        RECT 217.950 186.600 220.050 187.050 ;
        RECT 208.950 185.400 220.050 186.600 ;
        RECT 208.950 184.950 211.050 185.400 ;
        RECT 217.950 184.950 220.050 185.400 ;
        RECT 256.950 186.600 259.050 187.050 ;
        RECT 307.950 186.600 310.050 187.050 ;
        RECT 256.950 185.400 310.050 186.600 ;
        RECT 428.400 186.600 429.600 188.400 ;
        RECT 730.950 188.400 748.050 189.600 ;
        RECT 730.950 187.950 733.050 188.400 ;
        RECT 745.950 187.950 748.050 188.400 ;
        RECT 751.950 189.600 754.050 190.050 ;
        RECT 760.950 189.600 763.050 190.050 ;
        RECT 766.950 189.600 769.050 190.050 ;
        RECT 751.950 188.400 769.050 189.600 ;
        RECT 751.950 187.950 754.050 188.400 ;
        RECT 760.950 187.950 763.050 188.400 ;
        RECT 766.950 187.950 769.050 188.400 ;
        RECT 775.950 189.600 778.050 190.050 ;
        RECT 793.950 189.600 796.050 190.050 ;
        RECT 775.950 188.400 796.050 189.600 ;
        RECT 775.950 187.950 778.050 188.400 ;
        RECT 793.950 187.950 796.050 188.400 ;
        RECT 439.950 186.600 442.050 187.050 ;
        RECT 428.400 185.400 442.050 186.600 ;
        RECT 256.950 184.950 259.050 185.400 ;
        RECT 307.950 184.950 310.050 185.400 ;
        RECT 439.950 184.950 442.050 185.400 ;
        RECT 448.950 186.600 451.050 187.050 ;
        RECT 475.950 186.600 478.050 187.050 ;
        RECT 448.950 185.400 478.050 186.600 ;
        RECT 448.950 184.950 451.050 185.400 ;
        RECT 475.950 184.950 478.050 185.400 ;
        RECT 655.950 186.600 658.050 187.050 ;
        RECT 700.950 186.600 703.050 187.050 ;
        RECT 655.950 185.400 703.050 186.600 ;
        RECT 655.950 184.950 658.050 185.400 ;
        RECT 700.950 184.950 703.050 185.400 ;
        RECT 7.950 182.100 10.050 184.200 ;
        RECT 31.950 183.750 34.050 184.200 ;
        RECT 97.950 183.750 100.050 184.200 ;
        RECT 31.950 182.550 100.050 183.750 ;
        RECT 124.950 183.600 127.050 184.050 ;
        RECT 31.950 182.100 34.050 182.550 ;
        RECT 97.950 182.100 100.050 182.550 ;
        RECT 116.400 182.400 127.050 183.600 ;
        RECT 8.400 178.050 9.600 182.100 ;
        RECT 4.950 176.400 9.600 178.050 ;
        RECT 31.950 177.600 34.050 178.050 ;
        RECT 116.400 177.900 117.600 182.400 ;
        RECT 124.950 181.950 127.050 182.400 ;
        RECT 193.950 183.600 196.050 184.050 ;
        RECT 213.000 183.600 217.050 184.050 ;
        RECT 193.950 182.400 207.600 183.600 ;
        RECT 193.950 181.950 196.050 182.400 ;
        RECT 206.400 178.050 207.600 182.400 ;
        RECT 212.400 181.950 217.050 183.600 ;
        RECT 220.950 183.600 223.050 184.050 ;
        RECT 229.950 183.600 232.050 184.200 ;
        RECT 238.950 183.600 241.050 184.050 ;
        RECT 220.950 182.400 232.050 183.600 ;
        RECT 220.950 181.950 223.050 182.400 ;
        RECT 229.950 182.100 232.050 182.400 ;
        RECT 233.400 182.400 241.050 183.600 ;
        RECT 212.400 178.050 213.600 181.950 ;
        RECT 233.400 180.600 234.600 182.400 ;
        RECT 238.950 181.950 241.050 182.400 ;
        RECT 268.950 182.100 271.050 184.200 ;
        RECT 277.950 183.600 280.050 184.050 ;
        RECT 295.950 183.600 298.050 184.050 ;
        RECT 304.950 183.600 307.050 184.200 ;
        RECT 277.950 182.400 288.600 183.600 ;
        RECT 256.950 180.600 259.050 181.050 ;
        RECT 227.400 179.400 234.600 180.600 ;
        RECT 242.400 179.400 259.050 180.600 ;
        RECT 37.950 177.600 40.050 177.900 ;
        RECT 31.950 176.400 40.050 177.600 ;
        RECT 4.950 175.950 9.000 176.400 ;
        RECT 31.950 175.950 34.050 176.400 ;
        RECT 37.950 175.800 40.050 176.400 ;
        RECT 79.950 177.600 82.050 177.900 ;
        RECT 94.950 177.600 97.050 177.900 ;
        RECT 79.950 177.450 97.050 177.600 ;
        RECT 106.950 177.450 109.050 177.900 ;
        RECT 79.950 176.400 109.050 177.450 ;
        RECT 79.950 175.800 82.050 176.400 ;
        RECT 94.950 176.250 109.050 176.400 ;
        RECT 94.950 175.800 97.050 176.250 ;
        RECT 106.950 175.800 109.050 176.250 ;
        RECT 115.950 175.800 118.050 177.900 ;
        RECT 121.950 177.450 124.050 177.900 ;
        RECT 127.950 177.450 130.050 177.900 ;
        RECT 121.950 176.250 130.050 177.450 ;
        RECT 121.950 175.800 124.050 176.250 ;
        RECT 127.950 175.800 130.050 176.250 ;
        RECT 136.950 177.600 139.050 177.900 ;
        RECT 148.950 177.600 151.050 178.050 ;
        RECT 136.950 176.400 151.050 177.600 ;
        RECT 136.950 175.800 139.050 176.400 ;
        RECT 148.950 175.950 151.050 176.400 ;
        RECT 181.950 177.600 184.050 178.050 ;
        RECT 190.950 177.600 193.050 177.900 ;
        RECT 181.950 176.400 193.050 177.600 ;
        RECT 181.950 175.950 184.050 176.400 ;
        RECT 190.950 175.800 193.050 176.400 ;
        RECT 205.950 175.950 208.050 178.050 ;
        RECT 211.950 175.950 214.050 178.050 ;
        RECT 227.400 177.900 228.600 179.400 ;
        RECT 242.400 177.900 243.600 179.400 ;
        RECT 256.950 178.950 259.050 179.400 ;
        RECT 226.950 175.800 229.050 177.900 ;
        RECT 241.950 175.800 244.050 177.900 ;
        RECT 269.400 177.600 270.600 182.100 ;
        RECT 277.950 181.950 280.050 182.400 ;
        RECT 287.400 178.050 288.600 182.400 ;
        RECT 295.950 182.400 307.050 183.600 ;
        RECT 295.950 181.950 298.050 182.400 ;
        RECT 304.950 182.100 307.050 182.400 ;
        RECT 310.950 182.100 313.050 184.200 ;
        RECT 352.950 183.750 355.050 184.200 ;
        RECT 364.950 183.750 367.050 184.200 ;
        RECT 352.950 182.550 367.050 183.750 ;
        RECT 352.950 182.100 355.050 182.550 ;
        RECT 364.950 182.100 367.050 182.550 ;
        RECT 376.950 183.750 379.050 184.200 ;
        RECT 391.950 183.750 394.050 184.200 ;
        RECT 376.950 182.550 394.050 183.750 ;
        RECT 376.950 182.100 379.050 182.550 ;
        RECT 391.950 182.100 394.050 182.550 ;
        RECT 311.400 178.050 312.600 182.100 ;
        RECT 397.950 181.950 400.050 184.050 ;
        RECT 403.950 182.100 406.050 184.200 ;
        RECT 409.950 183.600 412.050 184.200 ;
        RECT 418.950 183.600 421.050 184.200 ;
        RECT 409.950 182.400 421.050 183.600 ;
        RECT 409.950 182.100 412.050 182.400 ;
        RECT 418.950 182.100 421.050 182.400 ;
        RECT 424.950 182.100 427.050 184.200 ;
        RECT 505.950 183.600 508.050 184.350 ;
        RECT 529.950 183.600 532.050 184.050 ;
        RECT 505.950 182.400 532.050 183.600 ;
        RECT 505.950 182.250 508.050 182.400 ;
        RECT 280.950 177.600 283.050 178.050 ;
        RECT 269.400 176.400 283.050 177.600 ;
        RECT 280.950 175.950 283.050 176.400 ;
        RECT 286.950 175.950 289.050 178.050 ;
        RECT 292.950 177.600 295.050 178.050 ;
        RECT 301.950 177.600 304.050 177.900 ;
        RECT 292.950 176.400 304.050 177.600 ;
        RECT 311.400 176.400 316.050 178.050 ;
        RECT 292.950 175.950 295.050 176.400 ;
        RECT 301.950 175.800 304.050 176.400 ;
        RECT 312.000 175.950 316.050 176.400 ;
        RECT 319.950 177.600 322.050 178.050 ;
        RECT 328.950 177.600 331.050 177.900 ;
        RECT 379.950 177.600 382.050 177.900 ;
        RECT 319.950 176.400 382.050 177.600 ;
        RECT 398.400 177.600 399.600 181.950 ;
        RECT 400.950 177.600 403.050 177.900 ;
        RECT 398.400 176.400 403.050 177.600 ;
        RECT 319.950 175.950 322.050 176.400 ;
        RECT 328.950 175.800 331.050 176.400 ;
        RECT 379.950 175.800 382.050 176.400 ;
        RECT 400.950 175.800 403.050 176.400 ;
        RECT 64.950 174.600 67.050 175.050 ;
        RECT 85.950 174.600 88.050 175.050 ;
        RECT 121.950 174.600 124.050 174.750 ;
        RECT 64.950 173.400 124.050 174.600 ;
        RECT 64.950 172.950 67.050 173.400 ;
        RECT 85.950 172.950 88.050 173.400 ;
        RECT 121.950 172.650 124.050 173.400 ;
        RECT 217.950 174.600 220.050 175.050 ;
        RECT 232.950 174.600 235.050 175.050 ;
        RECT 217.950 173.400 235.050 174.600 ;
        RECT 217.950 172.950 220.050 173.400 ;
        RECT 232.950 172.950 235.050 173.400 ;
        RECT 316.950 174.600 319.050 175.050 ;
        RECT 346.950 174.600 349.050 175.050 ;
        RECT 316.950 173.400 349.050 174.600 ;
        RECT 316.950 172.950 319.050 173.400 ;
        RECT 346.950 172.950 349.050 173.400 ;
        RECT 385.950 174.600 388.050 175.050 ;
        RECT 404.400 174.600 405.600 182.100 ;
        RECT 425.400 178.050 426.600 182.100 ;
        RECT 529.950 181.950 532.050 182.400 ;
        RECT 559.950 183.750 562.050 184.200 ;
        RECT 577.950 183.750 580.050 184.200 ;
        RECT 559.950 182.550 580.050 183.750 ;
        RECT 559.950 182.100 562.050 182.550 ;
        RECT 577.950 182.100 580.050 182.550 ;
        RECT 601.950 183.600 604.050 184.050 ;
        RECT 613.950 183.600 616.050 184.350 ;
        RECT 601.950 182.400 616.050 183.600 ;
        RECT 601.950 181.950 604.050 182.400 ;
        RECT 613.950 182.250 616.050 182.400 ;
        RECT 628.950 183.600 631.050 184.350 ;
        RECT 649.950 183.600 652.050 184.200 ;
        RECT 628.950 182.400 652.050 183.600 ;
        RECT 628.950 182.250 631.050 182.400 ;
        RECT 425.400 176.400 430.050 178.050 ;
        RECT 426.000 175.950 430.050 176.400 ;
        RECT 478.950 177.600 481.050 178.050 ;
        RECT 490.950 177.600 493.050 177.900 ;
        RECT 478.950 177.450 493.050 177.600 ;
        RECT 508.950 177.450 511.050 178.050 ;
        RECT 514.950 177.450 517.050 177.900 ;
        RECT 478.950 176.400 517.050 177.450 ;
        RECT 478.950 175.950 481.050 176.400 ;
        RECT 490.950 176.250 517.050 176.400 ;
        RECT 490.950 175.800 493.050 176.250 ;
        RECT 508.950 175.950 511.050 176.250 ;
        RECT 514.950 175.800 517.050 176.250 ;
        RECT 568.950 177.600 571.050 178.050 ;
        RECT 610.950 177.600 613.050 178.050 ;
        RECT 568.950 176.400 613.050 177.600 ;
        RECT 568.950 175.950 571.050 176.400 ;
        RECT 610.950 175.950 613.050 176.400 ;
        RECT 622.950 177.600 625.050 178.050 ;
        RECT 629.400 177.600 630.600 182.250 ;
        RECT 649.950 182.100 652.050 182.400 ;
        RECT 658.950 181.950 661.050 184.050 ;
        RECT 676.950 183.600 681.000 184.050 ;
        RECT 715.950 183.600 718.050 184.050 ;
        RECT 724.950 183.600 727.050 184.200 ;
        RECT 676.950 181.950 681.600 183.600 ;
        RECT 715.950 182.400 727.050 183.600 ;
        RECT 727.950 183.600 730.050 187.050 ;
        RECT 781.950 186.600 784.050 187.050 ;
        RECT 790.950 186.600 793.050 187.050 ;
        RECT 781.950 185.400 793.050 186.600 ;
        RECT 781.950 184.950 784.050 185.400 ;
        RECT 790.950 184.950 793.050 185.400 ;
        RECT 757.950 183.600 762.000 184.050 ;
        RECT 727.950 183.000 735.600 183.600 ;
        RECT 728.400 182.400 735.600 183.000 ;
        RECT 715.950 181.950 718.050 182.400 ;
        RECT 724.950 182.100 727.050 182.400 ;
        RECT 659.400 178.050 660.600 181.950 ;
        RECT 622.950 176.400 630.600 177.600 ;
        RECT 631.950 177.600 634.050 178.050 ;
        RECT 652.950 177.600 655.050 177.900 ;
        RECT 631.950 176.400 655.050 177.600 ;
        RECT 622.950 175.950 625.050 176.400 ;
        RECT 631.950 175.950 634.050 176.400 ;
        RECT 652.950 175.800 655.050 176.400 ;
        RECT 658.950 175.950 661.050 178.050 ;
        RECT 680.400 177.900 681.600 181.950 ;
        RECT 734.400 178.050 735.600 182.400 ;
        RECT 757.950 181.950 762.600 183.600 ;
        RECT 761.400 178.050 762.600 181.950 ;
        RECT 763.950 180.600 766.050 184.050 ;
        RECT 778.950 183.750 781.050 184.200 ;
        RECT 787.950 183.750 790.050 184.200 ;
        RECT 778.950 182.550 790.050 183.750 ;
        RECT 778.950 182.100 781.050 182.550 ;
        RECT 787.950 182.100 790.050 182.550 ;
        RECT 826.950 183.600 829.050 184.200 ;
        RECT 838.950 183.600 841.050 184.200 ;
        RECT 826.950 182.400 841.050 183.600 ;
        RECT 826.950 182.100 829.050 182.400 ;
        RECT 838.950 182.100 841.050 182.400 ;
        RECT 817.950 180.600 820.050 181.050 ;
        RECT 763.950 180.000 820.050 180.600 ;
        RECT 764.400 179.400 820.050 180.000 ;
        RECT 817.950 178.950 820.050 179.400 ;
        RECT 679.950 175.800 682.050 177.900 ;
        RECT 715.950 177.450 718.050 177.900 ;
        RECT 721.950 177.450 724.050 177.900 ;
        RECT 715.950 176.250 724.050 177.450 ;
        RECT 715.950 175.800 718.050 176.250 ;
        RECT 721.950 175.800 724.050 176.250 ;
        RECT 733.950 175.950 736.050 178.050 ;
        RECT 748.950 177.600 751.050 177.900 ;
        RECT 760.950 177.600 763.050 178.050 ;
        RECT 748.950 176.400 763.050 177.600 ;
        RECT 748.950 175.800 751.050 176.400 ;
        RECT 760.950 175.950 763.050 176.400 ;
        RECT 385.950 173.400 405.600 174.600 ;
        RECT 421.950 174.600 424.050 175.050 ;
        RECT 448.950 174.600 451.050 175.050 ;
        RECT 472.950 174.600 475.050 175.050 ;
        RECT 421.950 173.400 475.050 174.600 ;
        RECT 385.950 172.950 388.050 173.400 ;
        RECT 421.950 172.950 424.050 173.400 ;
        RECT 448.950 172.950 451.050 173.400 ;
        RECT 472.950 172.950 475.050 173.400 ;
        RECT 547.950 174.600 550.050 175.050 ;
        RECT 553.950 174.600 556.050 175.050 ;
        RECT 742.950 174.600 745.050 175.050 ;
        RECT 775.950 174.600 778.050 175.050 ;
        RECT 547.950 173.400 556.050 174.600 ;
        RECT 547.950 172.950 550.050 173.400 ;
        RECT 553.950 172.950 556.050 173.400 ;
        RECT 710.400 173.400 778.050 174.600 ;
        RECT 710.400 172.050 711.600 173.400 ;
        RECT 742.950 172.950 745.050 173.400 ;
        RECT 775.950 172.950 778.050 173.400 ;
        RECT 787.950 174.600 790.050 175.050 ;
        RECT 814.950 174.600 817.050 175.050 ;
        RECT 787.950 173.400 817.050 174.600 ;
        RECT 787.950 172.950 790.050 173.400 ;
        RECT 814.950 172.950 817.050 173.400 ;
        RECT 100.950 171.600 103.050 172.050 ;
        RECT 118.950 171.600 121.050 172.050 ;
        RECT 100.950 170.400 121.050 171.600 ;
        RECT 100.950 169.950 103.050 170.400 ;
        RECT 118.950 169.950 121.050 170.400 ;
        RECT 136.950 171.600 139.050 172.050 ;
        RECT 145.950 171.600 148.050 172.050 ;
        RECT 136.950 170.400 148.050 171.600 ;
        RECT 136.950 169.950 139.050 170.400 ;
        RECT 145.950 169.950 148.050 170.400 ;
        RECT 220.950 171.600 223.050 172.050 ;
        RECT 229.950 171.600 232.050 172.050 ;
        RECT 220.950 170.400 232.050 171.600 ;
        RECT 220.950 169.950 223.050 170.400 ;
        RECT 229.950 169.950 232.050 170.400 ;
        RECT 235.950 171.600 238.050 172.050 ;
        RECT 250.950 171.600 253.050 172.050 ;
        RECT 235.950 170.400 253.050 171.600 ;
        RECT 235.950 169.950 238.050 170.400 ;
        RECT 250.950 169.950 253.050 170.400 ;
        RECT 286.950 171.600 289.050 172.050 ;
        RECT 310.950 171.600 313.050 172.050 ;
        RECT 286.950 170.400 313.050 171.600 ;
        RECT 286.950 169.950 289.050 170.400 ;
        RECT 310.950 169.950 313.050 170.400 ;
        RECT 391.950 171.600 394.050 172.050 ;
        RECT 403.950 171.600 406.050 172.050 ;
        RECT 391.950 170.400 406.050 171.600 ;
        RECT 391.950 169.950 394.050 170.400 ;
        RECT 403.950 169.950 406.050 170.400 ;
        RECT 616.950 171.600 619.050 172.050 ;
        RECT 694.950 171.600 697.050 172.050 ;
        RECT 709.950 171.600 712.050 172.050 ;
        RECT 616.950 170.400 712.050 171.600 ;
        RECT 616.950 169.950 619.050 170.400 ;
        RECT 694.950 169.950 697.050 170.400 ;
        RECT 709.950 169.950 712.050 170.400 ;
        RECT 727.950 171.600 730.050 172.050 ;
        RECT 736.950 171.600 739.050 172.050 ;
        RECT 727.950 170.400 739.050 171.600 ;
        RECT 727.950 169.950 730.050 170.400 ;
        RECT 736.950 169.950 739.050 170.400 ;
        RECT 745.950 171.600 748.050 171.900 ;
        RECT 769.950 171.600 772.050 172.050 ;
        RECT 745.950 170.400 772.050 171.600 ;
        RECT 745.950 169.800 748.050 170.400 ;
        RECT 769.950 169.950 772.050 170.400 ;
        RECT 790.950 171.600 793.050 172.050 ;
        RECT 799.950 171.600 802.050 172.050 ;
        RECT 790.950 170.400 802.050 171.600 ;
        RECT 790.950 169.950 793.050 170.400 ;
        RECT 799.950 169.950 802.050 170.400 ;
        RECT 280.950 168.600 283.050 169.050 ;
        RECT 394.950 168.600 397.050 169.050 ;
        RECT 280.950 167.400 397.050 168.600 ;
        RECT 280.950 166.950 283.050 167.400 ;
        RECT 394.950 166.950 397.050 167.400 ;
        RECT 778.950 168.600 781.050 169.050 ;
        RECT 808.950 168.600 811.050 169.050 ;
        RECT 778.950 167.400 811.050 168.600 ;
        RECT 778.950 166.950 781.050 167.400 ;
        RECT 808.950 166.950 811.050 167.400 ;
        RECT 49.950 165.600 52.050 166.050 ;
        RECT 154.950 165.600 157.050 166.050 ;
        RECT 49.950 164.400 157.050 165.600 ;
        RECT 49.950 163.950 52.050 164.400 ;
        RECT 154.950 163.950 157.050 164.400 ;
        RECT 295.950 165.600 298.050 166.050 ;
        RECT 322.950 165.600 325.050 166.050 ;
        RECT 295.950 164.400 325.050 165.600 ;
        RECT 295.950 163.950 298.050 164.400 ;
        RECT 322.950 163.950 325.050 164.400 ;
        RECT 334.950 165.600 337.050 166.050 ;
        RECT 400.950 165.600 403.050 166.050 ;
        RECT 436.950 165.600 439.050 166.050 ;
        RECT 484.950 165.600 487.050 166.050 ;
        RECT 334.950 164.400 393.600 165.600 ;
        RECT 334.950 163.950 337.050 164.400 ;
        RECT 10.950 162.600 13.050 163.050 ;
        RECT 22.950 162.600 25.050 163.050 ;
        RECT 28.950 162.600 31.050 163.050 ;
        RECT 10.950 161.400 31.050 162.600 ;
        RECT 10.950 160.950 13.050 161.400 ;
        RECT 22.950 160.950 25.050 161.400 ;
        RECT 28.950 160.950 31.050 161.400 ;
        RECT 319.950 162.600 322.050 163.050 ;
        RECT 334.950 162.600 337.050 162.900 ;
        RECT 361.950 162.600 364.050 163.050 ;
        RECT 319.950 161.400 364.050 162.600 ;
        RECT 392.400 162.600 393.600 164.400 ;
        RECT 400.950 164.400 439.050 165.600 ;
        RECT 400.950 163.950 403.050 164.400 ;
        RECT 436.950 163.950 439.050 164.400 ;
        RECT 473.400 164.400 487.050 165.600 ;
        RECT 473.400 162.600 474.600 164.400 ;
        RECT 484.950 163.950 487.050 164.400 ;
        RECT 502.950 165.600 505.050 166.050 ;
        RECT 556.950 165.600 559.050 166.050 ;
        RECT 502.950 164.400 559.050 165.600 ;
        RECT 502.950 163.950 505.050 164.400 ;
        RECT 556.950 163.950 559.050 164.400 ;
        RECT 595.950 165.600 598.050 166.050 ;
        RECT 691.950 165.600 694.050 166.050 ;
        RECT 595.950 164.400 694.050 165.600 ;
        RECT 595.950 163.950 598.050 164.400 ;
        RECT 691.950 163.950 694.050 164.400 ;
        RECT 697.950 165.600 700.050 166.050 ;
        RECT 772.950 165.600 775.050 166.050 ;
        RECT 697.950 164.400 775.050 165.600 ;
        RECT 697.950 163.950 700.050 164.400 ;
        RECT 772.950 163.950 775.050 164.400 ;
        RECT 392.400 161.400 474.600 162.600 ;
        RECT 793.950 162.600 796.050 163.050 ;
        RECT 841.950 162.600 844.050 163.050 ;
        RECT 793.950 161.400 844.050 162.600 ;
        RECT 319.950 160.950 322.050 161.400 ;
        RECT 334.950 160.800 337.050 161.400 ;
        RECT 361.950 160.950 364.050 161.400 ;
        RECT 793.950 160.950 796.050 161.400 ;
        RECT 841.950 160.950 844.050 161.400 ;
        RECT 388.950 159.600 391.050 160.050 ;
        RECT 478.950 159.600 481.050 160.050 ;
        RECT 388.950 158.400 481.050 159.600 ;
        RECT 388.950 157.950 391.050 158.400 ;
        RECT 478.950 157.950 481.050 158.400 ;
        RECT 691.950 159.600 694.050 160.050 ;
        RECT 736.950 159.600 739.050 160.050 ;
        RECT 790.950 159.600 793.050 160.050 ;
        RECT 691.950 158.400 793.050 159.600 ;
        RECT 691.950 157.950 694.050 158.400 ;
        RECT 736.950 157.950 739.050 158.400 ;
        RECT 790.950 157.950 793.050 158.400 ;
        RECT 115.950 156.600 118.050 157.050 ;
        RECT 160.950 156.600 163.050 157.050 ;
        RECT 115.950 155.400 163.050 156.600 ;
        RECT 115.950 154.950 118.050 155.400 ;
        RECT 160.950 154.950 163.050 155.400 ;
        RECT 340.950 156.600 343.050 157.050 ;
        RECT 511.950 156.600 514.050 157.050 ;
        RECT 340.950 155.400 514.050 156.600 ;
        RECT 340.950 154.950 343.050 155.400 ;
        RECT 511.950 154.950 514.050 155.400 ;
        RECT 532.950 156.600 535.050 157.050 ;
        RECT 640.950 156.600 643.050 157.050 ;
        RECT 532.950 155.400 643.050 156.600 ;
        RECT 532.950 154.950 535.050 155.400 ;
        RECT 640.950 154.950 643.050 155.400 ;
        RECT 688.950 156.600 691.050 157.050 ;
        RECT 709.950 156.600 712.050 157.050 ;
        RECT 688.950 155.400 712.050 156.600 ;
        RECT 688.950 154.950 691.050 155.400 ;
        RECT 709.950 154.950 712.050 155.400 ;
        RECT 346.950 153.600 349.050 154.050 ;
        RECT 421.950 153.600 424.050 154.050 ;
        RECT 346.950 152.400 424.050 153.600 ;
        RECT 346.950 151.950 349.050 152.400 ;
        RECT 421.950 151.950 424.050 152.400 ;
        RECT 733.950 153.600 736.050 154.050 ;
        RECT 766.950 153.600 769.050 154.050 ;
        RECT 733.950 152.400 769.050 153.600 ;
        RECT 733.950 151.950 736.050 152.400 ;
        RECT 766.950 151.950 769.050 152.400 ;
        RECT 130.950 150.600 133.050 151.050 ;
        RECT 232.950 150.600 235.050 151.050 ;
        RECT 130.950 149.400 235.050 150.600 ;
        RECT 130.950 148.950 133.050 149.400 ;
        RECT 232.950 148.950 235.050 149.400 ;
        RECT 475.950 150.600 478.050 151.050 ;
        RECT 517.950 150.600 520.050 151.050 ;
        RECT 475.950 149.400 520.050 150.600 ;
        RECT 475.950 148.950 478.050 149.400 ;
        RECT 517.950 148.950 520.050 149.400 ;
        RECT 562.950 150.600 565.050 151.050 ;
        RECT 586.950 150.600 589.050 151.050 ;
        RECT 562.950 149.400 589.050 150.600 ;
        RECT 562.950 148.950 565.050 149.400 ;
        RECT 586.950 148.950 589.050 149.400 ;
        RECT 604.950 150.600 607.050 151.050 ;
        RECT 613.950 150.600 616.050 151.050 ;
        RECT 604.950 149.400 616.050 150.600 ;
        RECT 604.950 148.950 607.050 149.400 ;
        RECT 613.950 148.950 616.050 149.400 ;
        RECT 817.950 150.600 820.050 151.050 ;
        RECT 859.950 150.600 862.050 151.050 ;
        RECT 817.950 149.400 862.050 150.600 ;
        RECT 817.950 148.950 820.050 149.400 ;
        RECT 859.950 148.950 862.050 149.400 ;
        RECT 223.950 147.600 226.050 148.050 ;
        RECT 241.950 147.600 244.050 148.050 ;
        RECT 223.950 146.400 244.050 147.600 ;
        RECT 223.950 145.950 226.050 146.400 ;
        RECT 241.950 145.950 244.050 146.400 ;
        RECT 247.950 147.600 250.050 148.050 ;
        RECT 286.950 147.600 289.050 148.050 ;
        RECT 247.950 146.400 289.050 147.600 ;
        RECT 247.950 145.950 250.050 146.400 ;
        RECT 286.950 145.950 289.050 146.400 ;
        RECT 352.950 147.600 355.050 148.050 ;
        RECT 358.800 147.600 360.900 148.050 ;
        RECT 352.950 146.400 360.900 147.600 ;
        RECT 352.950 145.950 355.050 146.400 ;
        RECT 358.800 145.950 360.900 146.400 ;
        RECT 361.950 147.600 364.050 148.050 ;
        RECT 400.950 147.600 403.050 148.050 ;
        RECT 361.950 146.400 403.050 147.600 ;
        RECT 361.950 145.950 364.050 146.400 ;
        RECT 400.950 145.950 403.050 146.400 ;
        RECT 442.950 147.600 445.050 148.050 ;
        RECT 532.950 147.600 535.050 148.050 ;
        RECT 442.950 146.400 535.050 147.600 ;
        RECT 442.950 145.950 445.050 146.400 ;
        RECT 532.950 145.950 535.050 146.400 ;
        RECT 670.950 147.600 673.050 148.050 ;
        RECT 676.950 147.600 679.050 148.050 ;
        RECT 697.950 147.600 700.050 148.050 ;
        RECT 670.950 146.400 700.050 147.600 ;
        RECT 670.950 145.950 673.050 146.400 ;
        RECT 676.950 145.950 679.050 146.400 ;
        RECT 697.950 145.950 700.050 146.400 ;
        RECT 790.950 147.600 793.050 148.050 ;
        RECT 790.950 147.000 849.600 147.600 ;
        RECT 790.950 146.400 850.050 147.000 ;
        RECT 790.950 145.950 793.050 146.400 ;
        RECT 49.950 144.600 52.050 145.050 ;
        RECT 91.950 144.600 94.050 145.050 ;
        RECT 103.950 144.600 106.050 145.050 ;
        RECT 49.950 143.400 87.600 144.600 ;
        RECT 49.950 142.950 52.050 143.400 ;
        RECT 13.950 141.600 16.050 142.050 ;
        RECT 40.950 141.600 43.050 142.050 ;
        RECT 13.950 140.400 43.050 141.600 ;
        RECT 86.400 141.600 87.600 143.400 ;
        RECT 91.950 143.400 106.050 144.600 ;
        RECT 91.950 142.950 94.050 143.400 ;
        RECT 103.950 142.950 106.050 143.400 ;
        RECT 151.950 144.600 154.050 145.050 ;
        RECT 208.950 144.600 211.050 145.050 ;
        RECT 151.950 143.400 211.050 144.600 ;
        RECT 151.950 142.950 154.050 143.400 ;
        RECT 208.950 142.950 211.050 143.400 ;
        RECT 220.950 144.600 223.050 145.050 ;
        RECT 307.950 144.600 310.050 145.050 ;
        RECT 349.950 144.600 352.050 145.050 ;
        RECT 406.950 144.600 409.050 145.050 ;
        RECT 424.950 144.600 427.050 145.050 ;
        RECT 220.950 143.400 427.050 144.600 ;
        RECT 220.950 142.950 223.050 143.400 ;
        RECT 307.950 142.950 310.050 143.400 ;
        RECT 349.950 142.950 352.050 143.400 ;
        RECT 406.950 142.950 409.050 143.400 ;
        RECT 424.950 142.950 427.050 143.400 ;
        RECT 508.950 144.600 511.050 145.050 ;
        RECT 520.950 144.600 523.050 145.050 ;
        RECT 529.950 144.600 532.050 145.050 ;
        RECT 508.950 143.400 523.050 144.600 ;
        RECT 508.950 142.950 511.050 143.400 ;
        RECT 520.950 142.950 523.050 143.400 ;
        RECT 524.400 143.400 532.050 144.600 ;
        RECT 169.950 141.600 172.050 142.050 ;
        RECT 86.400 140.400 117.600 141.600 ;
        RECT 13.950 139.950 16.050 140.400 ;
        RECT 40.950 139.950 43.050 140.400 ;
        RECT 31.950 138.600 34.050 139.200 ;
        RECT 31.950 137.400 45.600 138.600 ;
        RECT 31.950 137.100 34.050 137.400 ;
        RECT 4.950 132.600 7.050 133.050 ;
        RECT 10.950 132.600 13.050 132.900 ;
        RECT 4.950 131.400 13.050 132.600 ;
        RECT 44.400 132.600 45.600 137.400 ;
        RECT 55.950 135.600 58.050 139.050 ;
        RECT 64.950 138.600 67.050 139.200 ;
        RECT 70.950 138.600 73.050 139.050 ;
        RECT 64.950 137.400 73.050 138.600 ;
        RECT 64.950 137.100 67.050 137.400 ;
        RECT 70.950 136.950 73.050 137.400 ;
        RECT 79.950 138.750 82.050 139.200 ;
        RECT 97.950 138.750 100.050 139.200 ;
        RECT 79.950 137.550 100.050 138.750 ;
        RECT 79.950 137.100 82.050 137.550 ;
        RECT 97.950 137.100 100.050 137.550 ;
        RECT 116.400 136.050 117.600 140.400 ;
        RECT 158.400 140.400 172.050 141.600 ;
        RECT 121.950 138.600 124.050 139.050 ;
        RECT 139.950 138.750 142.050 139.200 ;
        RECT 145.950 138.750 148.050 139.200 ;
        RECT 121.950 137.400 129.600 138.600 ;
        RECT 121.950 136.950 124.050 137.400 ;
        RECT 96.000 135.600 100.050 136.050 ;
        RECT 53.400 135.000 58.050 135.600 ;
        RECT 53.400 134.400 57.600 135.000 ;
        RECT 46.950 132.600 49.050 132.900 ;
        RECT 44.400 131.400 49.050 132.600 ;
        RECT 4.950 130.950 7.050 131.400 ;
        RECT 10.950 130.800 13.050 131.400 ;
        RECT 46.950 130.800 49.050 131.400 ;
        RECT 53.400 130.050 54.600 134.400 ;
        RECT 95.400 133.950 100.050 135.600 ;
        RECT 115.950 133.950 118.050 136.050 ;
        RECT 128.400 135.600 129.600 137.400 ;
        RECT 139.950 137.550 148.050 138.750 ;
        RECT 139.950 137.100 142.050 137.550 ;
        RECT 145.950 137.100 148.050 137.550 ;
        RECT 158.400 135.600 159.600 140.400 ;
        RECT 169.950 139.950 172.050 140.400 ;
        RECT 223.950 139.950 226.050 142.050 ;
        RECT 256.950 141.600 259.050 142.050 ;
        RECT 262.950 141.600 265.050 142.050 ;
        RECT 256.950 140.400 265.050 141.600 ;
        RECT 256.950 139.950 259.050 140.400 ;
        RECT 262.950 139.950 265.050 140.400 ;
        RECT 268.950 141.600 271.050 142.050 ;
        RECT 274.950 141.600 277.050 142.050 ;
        RECT 268.950 140.400 277.050 141.600 ;
        RECT 268.950 139.950 271.050 140.400 ;
        RECT 274.950 139.950 277.050 140.400 ;
        RECT 286.950 141.600 289.050 142.050 ;
        RECT 292.950 141.600 295.050 142.050 ;
        RECT 286.950 140.400 295.050 141.600 ;
        RECT 286.950 139.950 289.050 140.400 ;
        RECT 292.950 139.950 295.050 140.400 ;
        RECT 445.950 141.600 448.050 142.050 ;
        RECT 478.950 141.600 481.050 142.050 ;
        RECT 445.950 140.400 481.050 141.600 ;
        RECT 445.950 139.950 448.050 140.400 ;
        RECT 478.950 139.950 481.050 140.400 ;
        RECT 490.950 141.600 493.050 142.050 ;
        RECT 505.950 141.600 508.050 142.050 ;
        RECT 524.400 141.600 525.600 143.400 ;
        RECT 529.950 142.950 532.050 143.400 ;
        RECT 535.950 144.600 538.050 145.050 ;
        RECT 550.950 144.600 553.050 145.050 ;
        RECT 535.950 143.400 553.050 144.600 ;
        RECT 535.950 142.950 538.050 143.400 ;
        RECT 550.950 142.950 553.050 143.400 ;
        RECT 583.950 144.600 586.050 145.050 ;
        RECT 607.950 144.600 610.050 145.050 ;
        RECT 583.950 143.400 610.050 144.600 ;
        RECT 583.950 142.950 586.050 143.400 ;
        RECT 607.950 142.950 610.050 143.400 ;
        RECT 646.950 144.600 649.050 145.050 ;
        RECT 667.950 144.600 670.050 145.050 ;
        RECT 646.950 143.400 670.050 144.600 ;
        RECT 646.950 142.950 649.050 143.400 ;
        RECT 667.950 142.950 670.050 143.400 ;
        RECT 682.950 144.600 685.050 145.050 ;
        RECT 691.950 144.600 694.050 145.050 ;
        RECT 682.950 143.400 694.050 144.600 ;
        RECT 682.950 142.950 685.050 143.400 ;
        RECT 691.950 142.950 694.050 143.400 ;
        RECT 847.950 142.950 850.050 146.400 ;
        RECT 490.950 140.400 504.600 141.600 ;
        RECT 490.950 139.950 493.050 140.400 ;
        RECT 160.950 137.100 163.050 139.200 ;
        RECT 193.950 138.600 196.050 139.050 ;
        RECT 199.950 138.600 202.050 139.050 ;
        RECT 193.950 137.400 202.050 138.600 ;
        RECT 128.400 134.400 144.600 135.600 ;
        RECT 55.950 132.450 58.050 132.900 ;
        RECT 76.950 132.450 79.050 132.900 ;
        RECT 95.400 132.600 96.600 133.950 ;
        RECT 143.400 132.900 144.600 134.400 ;
        RECT 152.400 134.400 159.600 135.600 ;
        RECT 55.950 131.250 79.050 132.450 ;
        RECT 80.400 132.000 96.600 132.600 ;
        RECT 55.950 130.800 58.050 131.250 ;
        RECT 76.950 130.800 79.050 131.250 ;
        RECT 79.950 131.400 96.600 132.000 ;
        RECT 22.950 129.600 25.050 130.050 ;
        RECT 28.950 129.600 31.050 130.050 ;
        RECT 22.950 128.400 31.050 129.600 ;
        RECT 22.950 127.950 25.050 128.400 ;
        RECT 28.950 127.950 31.050 128.400 ;
        RECT 52.950 127.950 55.050 130.050 ;
        RECT 79.950 127.950 82.050 131.400 ;
        RECT 142.950 130.800 145.050 132.900 ;
        RECT 148.950 132.600 151.050 132.900 ;
        RECT 152.400 132.600 153.600 134.400 ;
        RECT 161.400 133.050 162.600 137.100 ;
        RECT 193.950 136.950 196.050 137.400 ;
        RECT 199.950 136.950 202.050 137.400 ;
        RECT 205.950 138.600 208.050 139.050 ;
        RECT 211.950 138.600 214.050 139.050 ;
        RECT 205.950 137.400 214.050 138.600 ;
        RECT 205.950 136.950 208.050 137.400 ;
        RECT 211.950 136.950 214.050 137.400 ;
        RECT 148.950 131.400 153.600 132.600 ;
        RECT 157.950 131.400 162.600 133.050 ;
        RECT 224.400 132.900 225.600 139.950 ;
        RECT 226.950 137.100 229.050 139.200 ;
        RECT 187.950 132.450 190.050 132.900 ;
        RECT 193.950 132.450 196.050 132.900 ;
        RECT 148.950 130.800 151.050 131.400 ;
        RECT 157.950 130.950 162.000 131.400 ;
        RECT 187.950 131.250 196.050 132.450 ;
        RECT 187.950 130.800 190.050 131.250 ;
        RECT 193.950 130.800 196.050 131.250 ;
        RECT 202.950 132.600 205.050 132.750 ;
        RECT 202.950 132.000 210.600 132.600 ;
        RECT 202.950 131.400 211.050 132.000 ;
        RECT 202.950 130.650 205.050 131.400 ;
        RECT 106.950 129.600 109.050 130.050 ;
        RECT 133.950 129.600 136.050 130.050 ;
        RECT 106.950 128.400 136.050 129.600 ;
        RECT 106.950 127.950 109.050 128.400 ;
        RECT 133.950 127.950 136.050 128.400 ;
        RECT 208.950 127.950 211.050 131.400 ;
        RECT 223.950 130.800 226.050 132.900 ;
        RECT 220.950 129.600 223.050 130.050 ;
        RECT 227.400 129.600 228.600 137.100 ;
        RECT 259.950 136.950 262.050 139.050 ;
        RECT 277.950 137.100 280.050 139.200 ;
        RECT 260.400 133.050 261.600 136.950 ;
        RECT 278.400 133.050 279.600 137.100 ;
        RECT 289.950 136.950 292.050 139.050 ;
        RECT 290.400 133.050 291.600 136.950 ;
        RECT 346.950 135.600 349.050 139.050 ;
        RECT 373.950 138.600 376.050 139.050 ;
        RECT 379.800 138.600 381.900 139.200 ;
        RECT 373.950 137.400 381.900 138.600 ;
        RECT 373.950 136.950 376.050 137.400 ;
        RECT 379.800 137.100 381.900 137.400 ;
        RECT 382.950 138.600 387.000 139.050 ;
        RECT 400.950 138.600 403.050 139.200 ;
        RECT 409.950 138.600 412.050 139.050 ;
        RECT 382.950 136.950 387.600 138.600 ;
        RECT 400.950 137.400 412.050 138.600 ;
        RECT 400.950 137.100 403.050 137.400 ;
        RECT 409.950 136.950 412.050 137.400 ;
        RECT 433.950 136.950 436.050 139.050 ;
        RECT 439.950 138.600 442.050 139.050 ;
        RECT 454.950 138.750 457.050 139.200 ;
        RECT 460.950 138.750 463.050 139.200 ;
        RECT 439.950 137.400 447.600 138.600 ;
        RECT 439.950 136.950 442.050 137.400 ;
        RECT 346.950 135.000 372.600 135.600 ;
        RECT 347.400 134.400 372.600 135.000 ;
        RECT 259.950 130.950 262.050 133.050 ;
        RECT 274.950 131.400 279.600 133.050 ;
        RECT 274.950 130.950 279.000 131.400 ;
        RECT 289.950 130.950 292.050 133.050 ;
        RECT 304.950 132.450 307.050 132.900 ;
        RECT 310.950 132.450 313.050 132.900 ;
        RECT 304.950 131.250 313.050 132.450 ;
        RECT 304.950 130.800 307.050 131.250 ;
        RECT 310.950 130.800 313.050 131.250 ;
        RECT 352.950 132.450 355.050 133.050 ;
        RECT 367.950 132.450 370.050 132.900 ;
        RECT 352.950 131.250 370.050 132.450 ;
        RECT 371.400 132.600 372.600 134.400 ;
        RECT 386.400 133.050 387.600 136.950 ;
        RECT 434.400 133.050 435.600 136.950 ;
        RECT 382.950 132.600 385.050 133.050 ;
        RECT 371.400 131.400 385.050 132.600 ;
        RECT 386.400 131.400 391.050 133.050 ;
        RECT 352.950 130.950 355.050 131.250 ;
        RECT 367.950 130.800 370.050 131.250 ;
        RECT 382.950 130.950 385.050 131.400 ;
        RECT 387.000 130.950 391.050 131.400 ;
        RECT 430.950 131.400 435.600 133.050 ;
        RECT 446.400 132.600 447.600 137.400 ;
        RECT 454.950 137.550 463.050 138.750 ;
        RECT 454.950 137.100 457.050 137.550 ;
        RECT 460.950 137.100 463.050 137.550 ;
        RECT 496.950 135.600 499.050 139.050 ;
        RECT 485.400 135.000 499.050 135.600 ;
        RECT 484.950 134.400 498.600 135.000 ;
        RECT 463.950 132.600 466.050 133.050 ;
        RECT 446.400 131.400 466.050 132.600 ;
        RECT 430.950 130.950 435.000 131.400 ;
        RECT 463.950 130.950 466.050 131.400 ;
        RECT 484.950 130.950 487.050 134.400 ;
        RECT 503.400 132.900 504.600 140.400 ;
        RECT 505.950 140.400 525.600 141.600 ;
        RECT 601.950 141.600 604.050 142.050 ;
        RECT 631.950 141.600 634.050 142.050 ;
        RECT 601.950 140.400 634.050 141.600 ;
        RECT 505.950 139.950 508.050 140.400 ;
        RECT 601.950 139.950 604.050 140.400 ;
        RECT 631.950 139.950 634.050 140.400 ;
        RECT 751.950 141.600 754.050 142.050 ;
        RECT 757.950 141.600 760.050 142.050 ;
        RECT 787.950 141.600 790.050 142.050 ;
        RECT 751.950 140.400 790.050 141.600 ;
        RECT 751.950 139.950 754.050 140.400 ;
        RECT 757.950 139.950 760.050 140.400 ;
        RECT 787.950 139.950 790.050 140.400 ;
        RECT 811.950 141.600 814.050 142.050 ;
        RECT 829.950 141.600 832.050 142.050 ;
        RECT 811.950 140.400 832.050 141.600 ;
        RECT 811.950 139.950 814.050 140.400 ;
        RECT 829.950 139.950 832.050 140.400 ;
        RECT 517.950 138.600 520.050 139.050 ;
        RECT 529.950 138.750 532.050 139.200 ;
        RECT 535.950 138.750 538.050 139.200 ;
        RECT 517.950 137.400 528.600 138.600 ;
        RECT 517.950 136.950 520.050 137.400 ;
        RECT 527.400 135.600 528.600 137.400 ;
        RECT 529.950 137.550 538.050 138.750 ;
        RECT 529.950 137.100 532.050 137.550 ;
        RECT 535.950 137.100 538.050 137.550 ;
        RECT 550.950 136.950 553.050 139.050 ;
        RECT 568.950 137.100 571.050 139.200 ;
        RECT 588.000 138.600 592.050 139.050 ;
        RECT 527.400 134.400 549.600 135.600 ;
        RECT 502.950 130.800 505.050 132.900 ;
        RECT 517.950 132.600 520.050 133.050 ;
        RECT 548.400 132.900 549.600 134.400 ;
        RECT 547.950 132.600 550.050 132.900 ;
        RECT 517.950 131.400 550.050 132.600 ;
        RECT 551.400 132.600 552.600 136.950 ;
        RECT 569.400 133.050 570.600 137.100 ;
        RECT 587.400 136.950 592.050 138.600 ;
        RECT 595.950 138.600 600.000 139.050 ;
        RECT 595.950 136.950 600.600 138.600 ;
        RECT 667.950 137.100 670.050 139.200 ;
        RECT 565.950 132.600 568.050 132.900 ;
        RECT 551.400 131.400 568.050 132.600 ;
        RECT 569.400 131.400 574.050 133.050 ;
        RECT 587.400 132.900 588.600 136.950 ;
        RECT 599.400 132.900 600.600 136.950 ;
        RECT 668.400 133.050 669.600 137.100 ;
        RECT 676.950 136.950 679.050 139.050 ;
        RECT 682.950 138.600 685.050 139.200 ;
        RECT 691.950 138.600 696.000 139.050 ;
        RECT 718.950 138.750 721.050 139.200 ;
        RECT 724.950 138.750 727.050 139.200 ;
        RECT 682.950 137.400 687.600 138.600 ;
        RECT 682.950 137.100 685.050 137.400 ;
        RECT 677.400 133.050 678.600 136.950 ;
        RECT 686.400 133.050 687.600 137.400 ;
        RECT 691.950 136.950 696.600 138.600 ;
        RECT 718.950 137.550 727.050 138.750 ;
        RECT 718.950 137.100 721.050 137.550 ;
        RECT 724.950 137.100 727.050 137.550 ;
        RECT 772.950 138.750 775.050 139.200 ;
        RECT 778.950 138.750 781.050 139.200 ;
        RECT 772.950 137.550 781.050 138.750 ;
        RECT 772.950 137.100 775.050 137.550 ;
        RECT 778.950 137.100 781.050 137.550 ;
        RECT 796.950 138.750 799.050 139.200 ;
        RECT 805.950 138.750 808.050 139.200 ;
        RECT 796.950 138.600 808.050 138.750 ;
        RECT 817.950 138.600 822.000 139.050 ;
        RECT 832.950 138.750 835.050 139.200 ;
        RECT 838.950 138.750 841.050 139.200 ;
        RECT 796.950 137.550 816.600 138.600 ;
        RECT 796.950 137.100 799.050 137.550 ;
        RECT 805.950 137.400 816.600 137.550 ;
        RECT 805.950 137.100 808.050 137.400 ;
        RECT 695.400 135.600 696.600 136.950 ;
        RECT 695.400 134.400 711.600 135.600 ;
        RECT 517.950 130.950 520.050 131.400 ;
        RECT 547.950 130.800 550.050 131.400 ;
        RECT 565.950 130.800 568.050 131.400 ;
        RECT 570.000 130.950 574.050 131.400 ;
        RECT 586.950 130.800 589.050 132.900 ;
        RECT 598.950 130.800 601.050 132.900 ;
        RECT 631.950 132.600 634.050 133.050 ;
        RECT 664.950 132.600 667.050 132.900 ;
        RECT 631.950 131.400 667.050 132.600 ;
        RECT 668.400 131.400 673.050 133.050 ;
        RECT 631.950 130.950 634.050 131.400 ;
        RECT 664.950 130.800 667.050 131.400 ;
        RECT 669.000 130.950 673.050 131.400 ;
        RECT 676.950 130.950 679.050 133.050 ;
        RECT 685.950 130.950 688.050 133.050 ;
        RECT 691.950 132.600 694.050 133.050 ;
        RECT 703.950 132.600 706.050 133.050 ;
        RECT 691.950 131.400 706.050 132.600 ;
        RECT 710.400 132.600 711.600 134.400 ;
        RECT 815.400 133.050 816.600 137.400 ;
        RECT 817.950 136.950 822.600 138.600 ;
        RECT 832.950 137.550 841.050 138.750 ;
        RECT 832.950 137.100 835.050 137.550 ;
        RECT 838.950 137.100 841.050 137.550 ;
        RECT 847.950 137.100 850.050 139.200 ;
        RECT 721.950 132.600 724.050 133.050 ;
        RECT 710.400 131.400 724.050 132.600 ;
        RECT 691.950 130.950 694.050 131.400 ;
        RECT 703.950 130.950 706.050 131.400 ;
        RECT 721.950 130.950 724.050 131.400 ;
        RECT 778.950 132.600 781.050 133.050 ;
        RECT 790.950 132.600 793.050 132.750 ;
        RECT 778.950 131.400 793.050 132.600 ;
        RECT 778.950 130.950 781.050 131.400 ;
        RECT 790.950 130.650 793.050 131.400 ;
        RECT 814.950 130.950 817.050 133.050 ;
        RECT 821.400 132.900 822.600 136.950 ;
        RECT 848.400 135.600 849.600 137.100 ;
        RECT 848.400 135.000 852.600 135.600 ;
        RECT 848.400 134.400 853.050 135.000 ;
        RECT 820.950 130.800 823.050 132.900 ;
        RECT 850.950 130.950 853.050 134.400 ;
        RECT 220.950 128.400 228.600 129.600 ;
        RECT 265.950 129.600 268.050 130.050 ;
        RECT 292.950 129.600 295.050 130.050 ;
        RECT 265.950 128.400 295.050 129.600 ;
        RECT 220.950 127.950 223.050 128.400 ;
        RECT 265.950 127.950 268.050 128.400 ;
        RECT 292.950 127.950 295.050 128.400 ;
        RECT 472.950 129.600 475.050 130.050 ;
        RECT 493.950 129.600 496.050 130.050 ;
        RECT 472.950 128.400 496.050 129.600 ;
        RECT 472.950 127.950 475.050 128.400 ;
        RECT 493.950 127.950 496.050 128.400 ;
        RECT 508.950 129.600 511.050 130.050 ;
        RECT 514.950 129.600 517.050 130.050 ;
        RECT 508.950 128.400 517.050 129.600 ;
        RECT 508.950 127.950 511.050 128.400 ;
        RECT 514.950 127.950 517.050 128.400 ;
        RECT 547.950 129.600 550.050 130.050 ;
        RECT 595.950 129.600 598.050 130.050 ;
        RECT 547.950 128.400 598.050 129.600 ;
        RECT 547.950 127.950 550.050 128.400 ;
        RECT 595.950 127.950 598.050 128.400 ;
        RECT 625.950 129.600 628.050 130.050 ;
        RECT 634.950 129.600 637.050 130.050 ;
        RECT 625.950 128.400 637.050 129.600 ;
        RECT 625.950 127.950 628.050 128.400 ;
        RECT 634.950 127.950 637.050 128.400 ;
        RECT 673.950 129.600 676.050 130.050 ;
        RECT 682.950 129.600 685.050 130.050 ;
        RECT 673.950 128.400 685.050 129.600 ;
        RECT 673.950 127.950 676.050 128.400 ;
        RECT 682.950 127.950 685.050 128.400 ;
        RECT 739.950 129.600 742.050 130.050 ;
        RECT 745.950 129.600 748.050 130.050 ;
        RECT 739.950 128.400 748.050 129.600 ;
        RECT 739.950 127.950 742.050 128.400 ;
        RECT 745.950 127.950 748.050 128.400 ;
        RECT 751.950 129.600 754.050 130.050 ;
        RECT 757.950 129.600 760.050 130.050 ;
        RECT 763.950 129.600 766.050 130.050 ;
        RECT 787.950 129.600 790.050 130.050 ;
        RECT 751.950 128.400 766.050 129.600 ;
        RECT 751.950 127.950 754.050 128.400 ;
        RECT 757.950 127.950 760.050 128.400 ;
        RECT 763.950 127.950 766.050 128.400 ;
        RECT 767.400 128.400 790.050 129.600 ;
        RECT 82.950 126.600 85.050 127.050 ;
        RECT 133.950 126.600 136.050 126.900 ;
        RECT 217.950 126.600 220.050 127.050 ;
        RECT 232.950 126.600 235.050 127.050 ;
        RECT 82.950 125.400 136.050 126.600 ;
        RECT 82.950 124.950 85.050 125.400 ;
        RECT 133.950 124.800 136.050 125.400 ;
        RECT 143.400 125.400 201.600 126.600 ;
        RECT 4.950 123.600 7.050 124.050 ;
        RECT 16.950 123.600 19.050 124.050 ;
        RECT 4.950 122.400 19.050 123.600 ;
        RECT 4.950 121.950 7.050 122.400 ;
        RECT 16.950 121.950 19.050 122.400 ;
        RECT 46.950 123.600 49.050 124.050 ;
        RECT 61.950 123.600 64.050 124.050 ;
        RECT 46.950 122.400 64.050 123.600 ;
        RECT 46.950 121.950 49.050 122.400 ;
        RECT 61.950 121.950 64.050 122.400 ;
        RECT 127.950 123.600 130.050 124.050 ;
        RECT 143.400 123.600 144.600 125.400 ;
        RECT 127.950 122.400 144.600 123.600 ;
        RECT 200.400 123.600 201.600 125.400 ;
        RECT 217.950 125.400 235.050 126.600 ;
        RECT 217.950 124.950 220.050 125.400 ;
        RECT 232.950 124.950 235.050 125.400 ;
        RECT 256.950 126.600 259.050 127.050 ;
        RECT 310.950 126.600 313.050 127.050 ;
        RECT 343.950 126.600 346.050 127.050 ;
        RECT 256.950 125.400 300.600 126.600 ;
        RECT 256.950 124.950 259.050 125.400 ;
        RECT 220.950 123.600 223.050 124.050 ;
        RECT 200.400 122.400 223.050 123.600 ;
        RECT 127.950 121.950 130.050 122.400 ;
        RECT 220.950 121.950 223.050 122.400 ;
        RECT 250.950 123.600 253.050 124.050 ;
        RECT 256.950 123.600 259.050 123.900 ;
        RECT 250.950 122.400 259.050 123.600 ;
        RECT 299.400 123.600 300.600 125.400 ;
        RECT 310.950 125.400 346.050 126.600 ;
        RECT 310.950 124.950 313.050 125.400 ;
        RECT 343.950 124.950 346.050 125.400 ;
        RECT 373.950 126.600 376.050 127.050 ;
        RECT 388.950 126.600 391.050 127.050 ;
        RECT 373.950 125.400 391.050 126.600 ;
        RECT 373.950 124.950 376.050 125.400 ;
        RECT 388.950 124.950 391.050 125.400 ;
        RECT 463.950 126.600 466.050 127.050 ;
        RECT 487.950 126.600 490.050 127.050 ;
        RECT 463.950 125.400 490.050 126.600 ;
        RECT 463.950 124.950 466.050 125.400 ;
        RECT 487.950 124.950 490.050 125.400 ;
        RECT 628.950 126.600 631.050 127.050 ;
        RECT 649.950 126.600 652.050 127.050 ;
        RECT 661.950 126.600 664.050 127.050 ;
        RECT 685.950 126.600 688.050 127.050 ;
        RECT 628.950 125.400 688.050 126.600 ;
        RECT 628.950 124.950 631.050 125.400 ;
        RECT 649.950 124.950 652.050 125.400 ;
        RECT 661.950 124.950 664.050 125.400 ;
        RECT 685.950 124.950 688.050 125.400 ;
        RECT 721.950 126.600 724.050 127.050 ;
        RECT 767.400 126.600 768.600 128.400 ;
        RECT 787.950 127.950 790.050 128.400 ;
        RECT 793.950 129.600 796.050 130.050 ;
        RECT 808.950 129.600 811.050 130.050 ;
        RECT 793.950 128.400 811.050 129.600 ;
        RECT 793.950 127.950 796.050 128.400 ;
        RECT 808.950 127.950 811.050 128.400 ;
        RECT 856.950 126.600 859.050 127.050 ;
        RECT 721.950 125.400 768.600 126.600 ;
        RECT 803.400 125.400 859.050 126.600 ;
        RECT 721.950 124.950 724.050 125.400 ;
        RECT 307.950 123.600 310.050 124.050 ;
        RECT 299.400 122.400 310.050 123.600 ;
        RECT 250.950 121.950 253.050 122.400 ;
        RECT 256.950 121.800 259.050 122.400 ;
        RECT 307.950 121.950 310.050 122.400 ;
        RECT 313.950 123.600 316.050 124.050 ;
        RECT 319.950 123.600 322.050 124.050 ;
        RECT 313.950 122.400 322.050 123.600 ;
        RECT 313.950 121.950 316.050 122.400 ;
        RECT 319.950 121.950 322.050 122.400 ;
        RECT 355.950 123.600 358.050 124.050 ;
        RECT 400.950 123.600 403.050 124.050 ;
        RECT 355.950 122.400 403.050 123.600 ;
        RECT 355.950 121.950 358.050 122.400 ;
        RECT 400.950 121.950 403.050 122.400 ;
        RECT 409.950 123.600 412.050 124.050 ;
        RECT 454.950 123.600 457.050 124.050 ;
        RECT 409.950 122.400 457.050 123.600 ;
        RECT 409.950 121.950 412.050 122.400 ;
        RECT 454.950 121.950 457.050 122.400 ;
        RECT 787.950 123.600 790.050 124.050 ;
        RECT 803.400 123.600 804.600 125.400 ;
        RECT 856.950 124.950 859.050 125.400 ;
        RECT 787.950 122.400 804.600 123.600 ;
        RECT 805.950 123.600 808.050 124.050 ;
        RECT 829.950 123.600 832.050 124.050 ;
        RECT 805.950 122.400 832.050 123.600 ;
        RECT 787.950 121.950 790.050 122.400 ;
        RECT 805.950 121.950 808.050 122.400 ;
        RECT 829.950 121.950 832.050 122.400 ;
        RECT 40.950 120.600 43.050 121.050 ;
        RECT 55.950 120.600 58.050 121.050 ;
        RECT 40.950 119.400 58.050 120.600 ;
        RECT 40.950 118.950 43.050 119.400 ;
        RECT 55.950 118.950 58.050 119.400 ;
        RECT 70.950 120.600 73.050 121.050 ;
        RECT 88.950 120.600 91.050 121.050 ;
        RECT 70.950 119.400 91.050 120.600 ;
        RECT 70.950 118.950 73.050 119.400 ;
        RECT 88.950 118.950 91.050 119.400 ;
        RECT 193.950 120.600 196.050 121.050 ;
        RECT 292.950 120.600 295.050 121.050 ;
        RECT 193.950 119.400 295.050 120.600 ;
        RECT 193.950 118.950 196.050 119.400 ;
        RECT 292.950 118.950 295.050 119.400 ;
        RECT 370.950 120.600 373.050 121.050 ;
        RECT 385.950 120.600 388.050 121.050 ;
        RECT 370.950 119.400 388.050 120.600 ;
        RECT 370.950 118.950 373.050 119.400 ;
        RECT 385.950 118.950 388.050 119.400 ;
        RECT 427.950 120.600 430.050 121.050 ;
        RECT 448.950 120.600 451.050 121.050 ;
        RECT 427.950 119.400 451.050 120.600 ;
        RECT 427.950 118.950 430.050 119.400 ;
        RECT 448.950 118.950 451.050 119.400 ;
        RECT 478.950 120.600 481.050 121.050 ;
        RECT 547.950 120.600 550.050 121.050 ;
        RECT 571.950 120.600 574.050 121.050 ;
        RECT 670.950 120.600 673.050 121.050 ;
        RECT 679.950 120.600 682.050 121.050 ;
        RECT 478.950 119.400 682.050 120.600 ;
        RECT 478.950 118.950 481.050 119.400 ;
        RECT 547.950 118.950 550.050 119.400 ;
        RECT 571.950 118.950 574.050 119.400 ;
        RECT 670.950 118.950 673.050 119.400 ;
        RECT 679.950 118.950 682.050 119.400 ;
        RECT 757.950 120.600 760.050 121.050 ;
        RECT 769.950 120.600 772.050 121.050 ;
        RECT 757.950 119.400 772.050 120.600 ;
        RECT 757.950 118.950 760.050 119.400 ;
        RECT 769.950 118.950 772.050 119.400 ;
        RECT 133.950 117.600 136.050 118.050 ;
        RECT 178.950 117.600 181.050 118.050 ;
        RECT 133.950 116.400 181.050 117.600 ;
        RECT 133.950 115.950 136.050 116.400 ;
        RECT 178.950 115.950 181.050 116.400 ;
        RECT 238.950 117.600 241.050 118.050 ;
        RECT 244.950 117.600 247.050 118.050 ;
        RECT 238.950 116.400 247.050 117.600 ;
        RECT 238.950 115.950 241.050 116.400 ;
        RECT 244.950 115.950 247.050 116.400 ;
        RECT 271.950 117.600 276.000 118.050 ;
        RECT 283.950 117.600 286.050 118.050 ;
        RECT 289.950 117.600 292.050 118.050 ;
        RECT 271.950 115.950 276.600 117.600 ;
        RECT 283.950 116.400 292.050 117.600 ;
        RECT 283.950 115.950 286.050 116.400 ;
        RECT 289.950 115.950 292.050 116.400 ;
        RECT 307.950 117.600 310.050 118.050 ;
        RECT 340.950 117.600 343.050 118.050 ;
        RECT 307.950 116.400 343.050 117.600 ;
        RECT 307.950 115.950 310.050 116.400 ;
        RECT 340.950 115.950 343.050 116.400 ;
        RECT 382.950 117.600 385.050 118.050 ;
        RECT 403.950 117.600 406.050 118.050 ;
        RECT 382.950 116.400 406.050 117.600 ;
        RECT 382.950 115.950 385.050 116.400 ;
        RECT 403.950 115.950 406.050 116.400 ;
        RECT 493.950 117.600 496.050 118.050 ;
        RECT 520.950 117.600 523.050 118.050 ;
        RECT 493.950 116.400 523.050 117.600 ;
        RECT 493.950 115.950 496.050 116.400 ;
        RECT 520.950 115.950 523.050 116.400 ;
        RECT 574.950 117.600 577.050 118.050 ;
        RECT 580.950 117.600 583.050 118.050 ;
        RECT 574.950 116.400 583.050 117.600 ;
        RECT 574.950 115.950 577.050 116.400 ;
        RECT 580.950 115.950 583.050 116.400 ;
        RECT 685.950 117.600 688.050 118.050 ;
        RECT 694.950 117.600 697.050 118.050 ;
        RECT 685.950 116.400 697.050 117.600 ;
        RECT 685.950 115.950 688.050 116.400 ;
        RECT 694.950 115.950 697.050 116.400 ;
        RECT 16.950 114.600 19.050 115.050 ;
        RECT 76.950 114.600 79.050 115.050 ;
        RECT 85.950 114.600 88.050 115.050 ;
        RECT 16.950 113.400 88.050 114.600 ;
        RECT 16.950 112.950 19.050 113.400 ;
        RECT 76.950 112.950 79.050 113.400 ;
        RECT 85.950 112.950 88.050 113.400 ;
        RECT 91.950 114.600 94.050 115.050 ;
        RECT 100.950 114.600 103.050 115.050 ;
        RECT 91.950 113.400 103.050 114.600 ;
        RECT 91.950 112.950 94.050 113.400 ;
        RECT 100.950 112.950 103.050 113.400 ;
        RECT 157.950 114.600 160.050 115.050 ;
        RECT 163.950 114.600 166.050 115.050 ;
        RECT 157.950 113.400 166.050 114.600 ;
        RECT 275.400 114.600 276.600 115.950 ;
        RECT 349.950 114.600 352.050 115.050 ;
        RECT 394.950 114.600 397.050 115.050 ;
        RECT 275.400 113.400 330.600 114.600 ;
        RECT 157.950 112.950 160.050 113.400 ;
        RECT 163.950 112.950 166.050 113.400 ;
        RECT 329.400 112.050 330.600 113.400 ;
        RECT 349.950 113.400 397.050 114.600 ;
        RECT 349.950 112.950 352.050 113.400 ;
        RECT 394.950 112.950 397.050 113.400 ;
        RECT 412.950 114.600 415.050 115.050 ;
        RECT 421.950 114.600 424.050 115.050 ;
        RECT 460.950 114.600 463.050 115.050 ;
        RECT 412.950 113.400 463.050 114.600 ;
        RECT 412.950 112.950 415.050 113.400 ;
        RECT 421.950 112.950 424.050 113.400 ;
        RECT 460.950 112.950 463.050 113.400 ;
        RECT 544.950 114.600 547.050 115.050 ;
        RECT 559.950 114.600 562.050 115.050 ;
        RECT 565.950 114.600 568.050 115.050 ;
        RECT 571.950 114.600 574.050 115.050 ;
        RECT 619.950 114.600 622.050 115.050 ;
        RECT 658.950 114.600 661.050 115.050 ;
        RECT 682.950 114.600 685.050 115.050 ;
        RECT 802.950 114.600 805.050 115.050 ;
        RECT 544.950 113.400 805.050 114.600 ;
        RECT 544.950 112.950 547.050 113.400 ;
        RECT 559.950 112.950 562.050 113.400 ;
        RECT 565.950 112.950 568.050 113.400 ;
        RECT 571.950 112.950 574.050 113.400 ;
        RECT 619.950 112.950 622.050 113.400 ;
        RECT 658.950 112.950 661.050 113.400 ;
        RECT 682.950 112.950 685.050 113.400 ;
        RECT 802.950 112.950 805.050 113.400 ;
        RECT 34.950 111.600 37.050 112.050 ;
        RECT 43.950 111.600 46.050 112.050 ;
        RECT 34.950 110.400 46.050 111.600 ;
        RECT 34.950 109.950 37.050 110.400 ;
        RECT 43.950 109.950 46.050 110.400 ;
        RECT 70.950 111.600 73.050 112.050 ;
        RECT 79.950 111.600 82.050 112.050 ;
        RECT 70.950 110.400 82.050 111.600 ;
        RECT 70.950 109.950 73.050 110.400 ;
        RECT 79.950 109.950 82.050 110.400 ;
        RECT 166.950 111.600 169.050 112.050 ;
        RECT 187.950 111.600 190.050 112.050 ;
        RECT 211.950 111.600 214.050 112.050 ;
        RECT 235.950 111.600 238.050 112.050 ;
        RECT 271.950 111.600 274.050 112.050 ;
        RECT 166.950 110.400 180.600 111.600 ;
        RECT 166.950 109.950 169.050 110.400 ;
        RECT 97.950 108.600 100.050 108.900 ;
        RECT 179.400 108.600 180.600 110.400 ;
        RECT 187.950 110.400 274.050 111.600 ;
        RECT 187.950 109.950 190.050 110.400 ;
        RECT 211.950 109.950 214.050 110.400 ;
        RECT 235.950 109.950 238.050 110.400 ;
        RECT 271.950 109.950 274.050 110.400 ;
        RECT 328.950 111.600 331.050 112.050 ;
        RECT 376.950 111.600 379.050 112.050 ;
        RECT 430.950 111.600 433.050 112.050 ;
        RECT 328.950 110.400 433.050 111.600 ;
        RECT 328.950 109.950 331.050 110.400 ;
        RECT 376.950 109.950 379.050 110.400 ;
        RECT 430.950 109.950 433.050 110.400 ;
        RECT 436.950 109.950 439.050 112.050 ;
        RECT 607.950 111.600 610.050 112.050 ;
        RECT 613.950 111.600 616.050 112.050 ;
        RECT 607.950 110.400 616.050 111.600 ;
        RECT 607.950 109.950 610.050 110.400 ;
        RECT 613.950 109.950 616.050 110.400 ;
        RECT 628.950 111.600 631.050 112.050 ;
        RECT 649.950 111.600 652.050 112.050 ;
        RECT 628.950 110.400 652.050 111.600 ;
        RECT 628.950 109.950 631.050 110.400 ;
        RECT 649.950 109.950 652.050 110.400 ;
        RECT 667.950 111.600 670.050 112.050 ;
        RECT 676.950 111.600 679.050 112.050 ;
        RECT 667.950 110.400 679.050 111.600 ;
        RECT 667.950 109.950 670.050 110.400 ;
        RECT 676.950 109.950 679.050 110.400 ;
        RECT 697.950 111.600 700.050 112.050 ;
        RECT 760.950 111.600 763.050 112.050 ;
        RECT 697.950 110.400 763.050 111.600 ;
        RECT 697.950 109.950 700.050 110.400 ;
        RECT 760.950 109.950 763.050 110.400 ;
        RECT 193.950 108.600 196.050 109.050 ;
        RECT 97.950 107.400 174.600 108.600 ;
        RECT 179.400 107.400 196.050 108.600 ;
        RECT 97.950 106.800 100.050 107.400 ;
        RECT 34.950 104.100 37.050 106.200 ;
        RECT 46.950 105.600 49.050 106.050 ;
        RECT 52.950 105.600 55.050 106.200 ;
        RECT 46.950 104.400 55.050 105.600 ;
        RECT 7.950 102.600 10.050 103.050 ;
        RECT 35.400 102.600 36.600 104.100 ;
        RECT 46.950 103.950 49.050 104.400 ;
        RECT 52.950 104.100 55.050 104.400 ;
        RECT 58.950 105.600 61.050 106.200 ;
        RECT 58.950 104.400 63.600 105.600 ;
        RECT 58.950 104.100 61.050 104.400 ;
        RECT 7.950 101.400 36.600 102.600 ;
        RECT 7.950 100.950 10.050 101.400 ;
        RECT 62.400 100.050 63.600 104.400 ;
        RECT 173.400 102.600 174.600 107.400 ;
        RECT 193.950 106.950 196.050 107.400 ;
        RECT 292.950 108.600 295.050 109.050 ;
        RECT 337.950 108.600 340.050 109.050 ;
        RECT 292.950 107.400 340.050 108.600 ;
        RECT 292.950 106.950 295.050 107.400 ;
        RECT 337.950 106.950 340.050 107.400 ;
        RECT 175.950 105.750 178.050 106.200 ;
        RECT 181.950 105.750 184.050 106.200 ;
        RECT 175.950 104.550 184.050 105.750 ;
        RECT 175.950 104.100 178.050 104.550 ;
        RECT 181.950 104.100 184.050 104.550 ;
        RECT 202.950 105.600 205.050 106.050 ;
        RECT 211.950 105.600 214.050 106.350 ;
        RECT 202.950 104.400 214.050 105.600 ;
        RECT 202.950 103.950 205.050 104.400 ;
        RECT 211.950 104.250 214.050 104.400 ;
        RECT 238.950 105.600 243.000 106.050 ;
        RECT 238.950 103.950 243.600 105.600 ;
        RECT 295.950 104.100 298.050 106.200 ;
        RECT 355.950 105.600 358.050 109.050 ;
        RECT 409.950 108.600 412.050 109.050 ;
        RECT 386.400 107.400 412.050 108.600 ;
        RECT 361.950 105.600 364.050 106.200 ;
        RECT 355.950 105.000 364.050 105.600 ;
        RECT 356.400 104.400 364.050 105.000 ;
        RECT 361.950 104.100 364.050 104.400 ;
        RECT 367.950 105.600 370.050 106.200 ;
        RECT 386.400 105.600 387.600 107.400 ;
        RECT 409.950 106.950 412.050 107.400 ;
        RECT 418.950 105.900 421.050 106.350 ;
        RECT 424.950 105.900 427.050 106.350 ;
        RECT 367.950 104.400 393.600 105.600 ;
        RECT 367.950 104.100 370.050 104.400 ;
        RECT 235.950 102.600 238.050 103.050 ;
        RECT 173.400 101.400 180.600 102.600 ;
        RECT 215.400 102.000 238.050 102.600 ;
        RECT 25.950 99.600 28.050 99.900 ;
        RECT 17.400 98.400 28.050 99.600 ;
        RECT 17.400 94.050 18.600 98.400 ;
        RECT 25.950 97.800 28.050 98.400 ;
        RECT 37.950 99.450 40.050 99.900 ;
        RECT 46.950 99.450 49.050 99.900 ;
        RECT 37.950 98.250 49.050 99.450 ;
        RECT 37.950 97.800 40.050 98.250 ;
        RECT 46.950 97.800 49.050 98.250 ;
        RECT 61.950 97.950 64.050 100.050 ;
        RECT 67.950 99.600 70.050 100.050 ;
        RECT 73.950 99.600 76.050 100.050 ;
        RECT 67.950 98.400 76.050 99.600 ;
        RECT 67.950 97.950 70.050 98.400 ;
        RECT 73.950 97.950 76.050 98.400 ;
        RECT 79.950 99.600 82.050 100.050 ;
        RECT 106.950 99.600 109.050 99.900 ;
        RECT 79.950 98.400 109.050 99.600 ;
        RECT 79.950 97.950 82.050 98.400 ;
        RECT 106.950 97.800 109.050 98.400 ;
        RECT 127.950 99.600 130.050 100.050 ;
        RECT 139.950 99.600 142.050 100.050 ;
        RECT 127.950 98.400 142.050 99.600 ;
        RECT 127.950 97.950 130.050 98.400 ;
        RECT 139.950 97.950 142.050 98.400 ;
        RECT 157.950 99.450 160.050 99.900 ;
        RECT 166.950 99.450 169.050 99.900 ;
        RECT 157.950 98.250 169.050 99.450 ;
        RECT 179.400 99.600 180.600 101.400 ;
        RECT 214.950 101.400 238.050 102.000 ;
        RECT 190.950 99.600 193.050 99.900 ;
        RECT 179.400 98.400 193.050 99.600 ;
        RECT 157.950 97.800 160.050 98.250 ;
        RECT 166.950 97.800 169.050 98.250 ;
        RECT 190.950 97.800 193.050 98.400 ;
        RECT 196.950 99.450 199.050 99.900 ;
        RECT 202.950 99.450 205.050 99.900 ;
        RECT 196.950 98.250 205.050 99.450 ;
        RECT 196.950 97.800 199.050 98.250 ;
        RECT 202.950 97.800 205.050 98.250 ;
        RECT 214.950 97.950 217.050 101.400 ;
        RECT 235.950 100.950 238.050 101.400 ;
        RECT 242.400 99.900 243.600 103.950 ;
        RECT 241.950 97.800 244.050 99.900 ;
        RECT 268.950 99.600 271.050 99.900 ;
        RECT 280.950 99.600 283.050 100.050 ;
        RECT 268.950 98.400 283.050 99.600 ;
        RECT 268.950 97.800 271.050 98.400 ;
        RECT 280.950 97.950 283.050 98.400 ;
        RECT 286.950 99.600 289.050 100.050 ;
        RECT 296.400 99.600 297.600 104.100 ;
        RECT 392.400 100.050 393.600 104.400 ;
        RECT 418.950 104.700 427.050 105.900 ;
        RECT 418.950 104.250 421.050 104.700 ;
        RECT 424.950 104.250 427.050 104.700 ;
        RECT 437.400 105.600 438.600 109.950 ;
        RECT 439.950 108.600 442.050 109.050 ;
        RECT 445.950 108.600 448.050 109.050 ;
        RECT 439.950 107.400 448.050 108.600 ;
        RECT 439.950 106.950 442.050 107.400 ;
        RECT 445.950 106.950 448.050 107.400 ;
        RECT 463.950 108.600 466.050 109.050 ;
        RECT 493.950 108.600 496.050 109.050 ;
        RECT 463.950 107.400 496.050 108.600 ;
        RECT 463.950 106.950 466.050 107.400 ;
        RECT 493.950 106.950 496.050 107.400 ;
        RECT 547.950 106.950 550.050 109.050 ;
        RECT 556.950 108.600 559.050 109.050 ;
        RECT 592.950 108.600 595.050 109.050 ;
        RECT 688.950 108.600 691.050 109.050 ;
        RECT 703.950 108.600 706.050 109.050 ;
        RECT 775.950 108.600 778.050 109.050 ;
        RECT 556.950 107.400 595.050 108.600 ;
        RECT 556.950 106.950 559.050 107.400 ;
        RECT 592.950 106.950 595.050 107.400 ;
        RECT 602.400 107.400 778.050 108.600 ;
        RECT 478.950 105.600 481.050 106.050 ;
        RECT 437.400 104.400 441.600 105.600 ;
        RECT 286.950 98.400 297.600 99.600 ;
        RECT 307.950 99.450 310.050 99.900 ;
        RECT 313.950 99.450 316.050 99.900 ;
        RECT 286.950 97.950 289.050 98.400 ;
        RECT 307.950 98.250 316.050 99.450 ;
        RECT 307.950 97.800 310.050 98.250 ;
        RECT 313.950 97.800 316.050 98.250 ;
        RECT 337.950 99.600 340.050 99.900 ;
        RECT 373.950 99.600 376.050 100.050 ;
        RECT 379.950 99.600 382.050 99.900 ;
        RECT 337.950 98.400 382.050 99.600 ;
        RECT 337.950 97.800 340.050 98.400 ;
        RECT 373.950 97.950 376.050 98.400 ;
        RECT 379.950 97.800 382.050 98.400 ;
        RECT 391.950 97.950 394.050 100.050 ;
        RECT 412.950 99.600 415.050 100.050 ;
        RECT 421.950 99.600 424.050 100.050 ;
        RECT 440.400 99.900 441.600 104.400 ;
        RECT 461.400 104.400 481.050 105.600 ;
        RECT 461.400 102.600 462.600 104.400 ;
        RECT 478.950 103.950 481.050 104.400 ;
        RECT 514.950 103.950 517.050 106.050 ;
        RECT 529.950 105.750 532.050 106.200 ;
        RECT 535.950 105.750 538.050 106.200 ;
        RECT 529.950 104.550 538.050 105.750 ;
        RECT 529.950 104.100 532.050 104.550 ;
        RECT 535.950 104.100 538.050 104.550 ;
        RECT 458.400 101.400 462.600 102.600 ;
        RECT 458.400 99.900 459.600 101.400 ;
        RECT 515.400 100.050 516.600 103.950 ;
        RECT 548.400 102.600 549.600 106.950 ;
        RECT 550.950 104.250 553.050 106.350 ;
        RECT 574.950 105.600 577.050 106.050 ;
        RECT 569.400 104.400 577.050 105.600 ;
        RECT 545.400 102.000 549.600 102.600 ;
        RECT 544.950 101.400 549.600 102.000 ;
        RECT 412.950 98.400 424.050 99.600 ;
        RECT 412.950 97.950 415.050 98.400 ;
        RECT 421.950 97.950 424.050 98.400 ;
        RECT 439.950 97.800 442.050 99.900 ;
        RECT 457.950 97.800 460.050 99.900 ;
        RECT 475.950 99.600 478.050 99.900 ;
        RECT 464.400 98.400 478.050 99.600 ;
        RECT 464.400 97.050 465.600 98.400 ;
        RECT 475.950 97.800 478.050 98.400 ;
        RECT 481.950 99.450 484.050 99.900 ;
        RECT 502.950 99.450 505.050 99.900 ;
        RECT 481.950 98.250 505.050 99.450 ;
        RECT 481.950 97.800 484.050 98.250 ;
        RECT 502.950 97.800 505.050 98.250 ;
        RECT 514.950 97.950 517.050 100.050 ;
        RECT 544.950 97.950 547.050 101.400 ;
        RECT 551.400 100.050 552.600 104.250 ;
        RECT 569.400 102.600 570.600 104.400 ;
        RECT 574.950 103.950 577.050 104.400 ;
        RECT 580.950 105.600 583.050 106.350 ;
        RECT 589.950 105.600 592.050 106.050 ;
        RECT 580.950 104.400 592.050 105.600 ;
        RECT 580.950 104.250 583.050 104.400 ;
        RECT 589.950 103.950 592.050 104.400 ;
        RECT 563.400 102.000 570.600 102.600 ;
        RECT 562.950 101.400 570.600 102.000 ;
        RECT 550.950 97.950 553.050 100.050 ;
        RECT 562.950 97.950 565.050 101.400 ;
        RECT 571.950 99.600 574.050 100.050 ;
        RECT 577.950 99.600 580.050 100.050 ;
        RECT 602.400 99.900 603.600 107.400 ;
        RECT 688.950 106.950 691.050 107.400 ;
        RECT 703.950 106.950 706.050 107.400 ;
        RECT 775.950 106.950 778.050 107.400 ;
        RECT 781.950 108.600 784.050 109.200 ;
        RECT 796.950 108.600 799.050 109.050 ;
        RECT 781.950 107.400 799.050 108.600 ;
        RECT 781.950 107.100 784.050 107.400 ;
        RECT 796.950 106.950 799.050 107.400 ;
        RECT 604.950 105.600 607.050 106.050 ;
        RECT 613.950 105.600 616.050 106.200 ;
        RECT 631.950 105.600 634.050 106.200 ;
        RECT 604.950 104.400 616.050 105.600 ;
        RECT 604.950 103.950 607.050 104.400 ;
        RECT 613.950 104.100 616.050 104.400 ;
        RECT 617.400 104.400 634.050 105.600 ;
        RECT 617.400 102.600 618.600 104.400 ;
        RECT 631.950 104.100 634.050 104.400 ;
        RECT 646.950 105.750 649.050 106.200 ;
        RECT 655.950 105.750 658.050 106.200 ;
        RECT 646.950 104.550 658.050 105.750 ;
        RECT 676.950 105.600 679.050 106.200 ;
        RECT 646.950 104.100 649.050 104.550 ;
        RECT 655.950 104.100 658.050 104.550 ;
        RECT 659.400 104.400 679.050 105.600 ;
        RECT 611.400 102.000 618.600 102.600 ;
        RECT 610.950 101.400 618.600 102.000 ;
        RECT 571.950 98.400 580.050 99.600 ;
        RECT 571.950 97.950 574.050 98.400 ;
        RECT 577.950 97.950 580.050 98.400 ;
        RECT 601.950 97.800 604.050 99.900 ;
        RECT 610.950 97.950 613.050 101.400 ;
        RECT 659.400 99.900 660.600 104.400 ;
        RECT 676.950 104.100 679.050 104.400 ;
        RECT 685.950 103.950 688.050 106.050 ;
        RECT 757.950 103.950 760.050 106.050 ;
        RECT 763.950 103.950 766.050 106.050 ;
        RECT 781.950 103.950 784.050 106.050 ;
        RECT 799.950 105.600 804.000 106.050 ;
        RECT 799.950 103.950 804.600 105.600 ;
        RECT 686.400 100.050 687.600 103.950 ;
        RECT 758.400 100.050 759.600 103.950 ;
        RECT 764.400 100.050 765.600 103.950 ;
        RECT 782.400 102.600 783.600 103.950 ;
        RECT 779.400 102.000 783.600 102.600 ;
        RECT 778.950 101.400 783.600 102.000 ;
        RECT 658.950 97.800 661.050 99.900 ;
        RECT 685.950 97.950 688.050 100.050 ;
        RECT 718.950 99.600 721.050 100.050 ;
        RECT 751.950 99.600 754.050 100.050 ;
        RECT 718.950 98.400 754.050 99.600 ;
        RECT 718.950 97.950 721.050 98.400 ;
        RECT 751.950 97.950 754.050 98.400 ;
        RECT 757.950 97.950 760.050 100.050 ;
        RECT 763.950 97.950 766.050 100.050 ;
        RECT 778.950 97.950 781.050 101.400 ;
        RECT 803.400 100.050 804.600 103.950 ;
        RECT 802.950 97.950 805.050 100.050 ;
        RECT 814.950 99.450 817.050 99.900 ;
        RECT 835.950 99.450 838.050 99.900 ;
        RECT 814.950 98.250 838.050 99.450 ;
        RECT 814.950 97.800 817.050 98.250 ;
        RECT 835.950 97.800 838.050 98.250 ;
        RECT 352.950 96.600 355.050 97.050 ;
        RECT 364.950 96.600 367.050 97.050 ;
        RECT 352.950 95.400 367.050 96.600 ;
        RECT 352.950 94.950 355.050 95.400 ;
        RECT 364.950 94.950 367.050 95.400 ;
        RECT 445.950 96.600 448.050 97.050 ;
        RECT 454.950 96.600 457.050 97.050 ;
        RECT 445.950 95.400 457.050 96.600 ;
        RECT 445.950 94.950 448.050 95.400 ;
        RECT 454.950 94.950 457.050 95.400 ;
        RECT 460.950 95.400 465.600 97.050 ;
        RECT 466.950 96.600 469.050 97.050 ;
        RECT 482.400 96.600 483.600 97.800 ;
        RECT 466.950 95.400 483.600 96.600 ;
        RECT 511.950 96.600 514.050 97.050 ;
        RECT 520.950 96.600 523.050 97.050 ;
        RECT 538.950 96.600 541.050 97.050 ;
        RECT 511.950 95.400 541.050 96.600 ;
        RECT 460.950 94.950 465.000 95.400 ;
        RECT 466.950 94.950 469.050 95.400 ;
        RECT 511.950 94.950 514.050 95.400 ;
        RECT 520.950 94.950 523.050 95.400 ;
        RECT 538.950 94.950 541.050 95.400 ;
        RECT 613.950 96.600 616.050 97.050 ;
        RECT 628.800 96.600 630.900 97.050 ;
        RECT 613.950 95.400 630.900 96.600 ;
        RECT 613.950 94.950 616.050 95.400 ;
        RECT 628.800 94.950 630.900 95.400 ;
        RECT 631.950 96.600 634.050 97.050 ;
        RECT 646.950 96.600 649.050 97.050 ;
        RECT 631.950 95.400 649.050 96.600 ;
        RECT 631.950 94.950 634.050 95.400 ;
        RECT 646.950 94.950 649.050 95.400 ;
        RECT 760.950 96.600 763.050 97.050 ;
        RECT 769.950 96.600 772.050 97.050 ;
        RECT 760.950 95.400 772.050 96.600 ;
        RECT 760.950 94.950 763.050 95.400 ;
        RECT 769.950 94.950 772.050 95.400 ;
        RECT 847.950 96.600 850.050 97.050 ;
        RECT 853.950 96.600 856.050 97.050 ;
        RECT 847.950 95.400 856.050 96.600 ;
        RECT 847.950 94.950 850.050 95.400 ;
        RECT 853.950 94.950 856.050 95.400 ;
        RECT 16.950 91.950 19.050 94.050 ;
        RECT 79.950 93.600 82.050 94.050 ;
        RECT 115.950 93.600 118.050 94.050 ;
        RECT 130.950 93.600 133.050 94.050 ;
        RECT 79.950 92.400 133.050 93.600 ;
        RECT 79.950 91.950 82.050 92.400 ;
        RECT 115.950 91.950 118.050 92.400 ;
        RECT 130.950 91.950 133.050 92.400 ;
        RECT 148.950 93.600 151.050 94.050 ;
        RECT 163.950 93.600 166.050 94.050 ;
        RECT 148.950 92.400 166.050 93.600 ;
        RECT 148.950 91.950 151.050 92.400 ;
        RECT 163.950 91.950 166.050 92.400 ;
        RECT 181.950 93.600 184.050 94.050 ;
        RECT 208.950 93.600 211.050 94.050 ;
        RECT 181.950 92.400 211.050 93.600 ;
        RECT 181.950 91.950 184.050 92.400 ;
        RECT 208.950 91.950 211.050 92.400 ;
        RECT 250.950 93.600 253.050 94.050 ;
        RECT 256.950 93.600 259.050 94.050 ;
        RECT 274.950 93.600 277.050 94.050 ;
        RECT 322.950 93.600 325.050 94.050 ;
        RECT 337.950 93.600 340.050 94.050 ;
        RECT 445.950 93.600 448.050 93.900 ;
        RECT 467.400 93.600 468.600 94.950 ;
        RECT 250.950 92.400 468.600 93.600 ;
        RECT 514.950 93.600 517.050 94.050 ;
        RECT 610.950 93.600 613.050 94.050 ;
        RECT 514.950 92.400 613.050 93.600 ;
        RECT 250.950 91.950 253.050 92.400 ;
        RECT 256.950 91.950 259.050 92.400 ;
        RECT 274.950 91.950 277.050 92.400 ;
        RECT 322.950 91.950 325.050 92.400 ;
        RECT 337.950 91.950 340.050 92.400 ;
        RECT 209.400 90.600 210.600 91.950 ;
        RECT 445.950 91.800 448.050 92.400 ;
        RECT 514.950 91.950 517.050 92.400 ;
        RECT 610.950 91.950 613.050 92.400 ;
        RECT 622.950 93.600 625.050 94.050 ;
        RECT 670.950 93.600 673.050 94.050 ;
        RECT 622.950 92.400 673.050 93.600 ;
        RECT 622.950 91.950 625.050 92.400 ;
        RECT 670.950 91.950 673.050 92.400 ;
        RECT 349.950 90.600 352.050 91.050 ;
        RECT 376.950 90.600 379.050 91.050 ;
        RECT 209.400 89.400 352.050 90.600 ;
        RECT 349.950 88.950 352.050 89.400 ;
        RECT 353.400 89.400 379.050 90.600 ;
        RECT 262.950 87.600 265.050 88.050 ;
        RECT 328.950 87.600 331.050 88.050 ;
        RECT 353.400 87.600 354.600 89.400 ;
        RECT 376.950 88.950 379.050 89.400 ;
        RECT 415.950 90.600 418.050 91.050 ;
        RECT 433.950 90.600 436.050 91.050 ;
        RECT 415.950 89.400 436.050 90.600 ;
        RECT 415.950 88.950 418.050 89.400 ;
        RECT 433.950 88.950 436.050 89.400 ;
        RECT 547.950 90.600 550.050 91.050 ;
        RECT 562.950 90.600 565.050 91.050 ;
        RECT 547.950 89.400 565.050 90.600 ;
        RECT 547.950 88.950 550.050 89.400 ;
        RECT 562.950 88.950 565.050 89.400 ;
        RECT 574.950 90.600 577.050 91.050 ;
        RECT 583.950 90.600 586.050 91.050 ;
        RECT 574.950 89.400 586.050 90.600 ;
        RECT 574.950 88.950 577.050 89.400 ;
        RECT 583.950 88.950 586.050 89.400 ;
        RECT 628.950 90.600 631.050 91.050 ;
        RECT 652.950 90.600 655.050 91.050 ;
        RECT 628.950 89.400 655.050 90.600 ;
        RECT 628.950 88.950 631.050 89.400 ;
        RECT 652.950 88.950 655.050 89.400 ;
        RECT 775.950 90.600 778.050 91.050 ;
        RECT 790.950 90.600 793.050 91.050 ;
        RECT 775.950 89.400 793.050 90.600 ;
        RECT 775.950 88.950 778.050 89.400 ;
        RECT 790.950 88.950 793.050 89.400 ;
        RECT 262.950 86.400 354.600 87.600 ;
        RECT 382.950 87.600 385.050 88.050 ;
        RECT 625.950 87.600 628.050 88.050 ;
        RECT 382.950 86.400 519.600 87.600 ;
        RECT 262.950 85.950 265.050 86.400 ;
        RECT 328.950 85.950 331.050 86.400 ;
        RECT 382.950 85.950 385.050 86.400 ;
        RECT 121.950 84.600 124.050 85.050 ;
        RECT 148.950 84.600 151.050 85.050 ;
        RECT 121.950 83.400 151.050 84.600 ;
        RECT 121.950 82.950 124.050 83.400 ;
        RECT 148.950 82.950 151.050 83.400 ;
        RECT 286.950 84.600 289.050 85.050 ;
        RECT 358.950 84.600 361.050 85.050 ;
        RECT 286.950 83.400 361.050 84.600 ;
        RECT 286.950 82.950 289.050 83.400 ;
        RECT 358.950 82.950 361.050 83.400 ;
        RECT 376.950 84.600 379.050 85.050 ;
        RECT 511.950 84.600 514.050 85.050 ;
        RECT 376.950 83.400 514.050 84.600 ;
        RECT 518.400 84.600 519.600 86.400 ;
        RECT 587.400 86.400 628.050 87.600 ;
        RECT 526.950 84.600 529.050 85.050 ;
        RECT 518.400 83.400 529.050 84.600 ;
        RECT 376.950 82.950 379.050 83.400 ;
        RECT 511.950 82.950 514.050 83.400 ;
        RECT 526.950 82.950 529.050 83.400 ;
        RECT 541.950 84.600 544.050 85.050 ;
        RECT 587.400 84.600 588.600 86.400 ;
        RECT 625.950 85.950 628.050 86.400 ;
        RECT 700.950 87.600 703.050 88.050 ;
        RECT 733.950 87.600 736.050 88.050 ;
        RECT 700.950 86.400 736.050 87.600 ;
        RECT 700.950 85.950 703.050 86.400 ;
        RECT 733.950 85.950 736.050 86.400 ;
        RECT 757.950 87.600 760.050 88.050 ;
        RECT 814.950 87.600 817.050 88.050 ;
        RECT 757.950 86.400 817.050 87.600 ;
        RECT 757.950 85.950 760.050 86.400 ;
        RECT 814.950 85.950 817.050 86.400 ;
        RECT 541.950 83.400 588.600 84.600 ;
        RECT 589.950 84.600 592.050 85.050 ;
        RECT 622.950 84.600 625.050 85.050 ;
        RECT 589.950 83.400 625.050 84.600 ;
        RECT 541.950 82.950 544.050 83.400 ;
        RECT 589.950 82.950 592.050 83.400 ;
        RECT 622.950 82.950 625.050 83.400 ;
        RECT 679.950 84.600 682.050 85.050 ;
        RECT 688.950 84.600 691.050 85.050 ;
        RECT 712.950 84.600 715.050 85.050 ;
        RECT 679.950 83.400 715.050 84.600 ;
        RECT 679.950 82.950 682.050 83.400 ;
        RECT 688.950 82.950 691.050 83.400 ;
        RECT 712.950 82.950 715.050 83.400 ;
        RECT 808.950 84.600 811.050 85.050 ;
        RECT 823.950 84.600 826.050 85.050 ;
        RECT 808.950 83.400 826.050 84.600 ;
        RECT 808.950 82.950 811.050 83.400 ;
        RECT 823.950 82.950 826.050 83.400 ;
        RECT 187.950 81.600 190.050 82.050 ;
        RECT 262.950 81.600 265.050 82.050 ;
        RECT 187.950 80.400 265.050 81.600 ;
        RECT 187.950 79.950 190.050 80.400 ;
        RECT 262.950 79.950 265.050 80.400 ;
        RECT 463.950 81.600 466.050 82.050 ;
        RECT 487.950 81.600 490.050 82.050 ;
        RECT 493.950 81.600 496.050 82.050 ;
        RECT 463.950 80.400 496.050 81.600 ;
        RECT 512.400 81.600 513.600 82.950 ;
        RECT 553.950 81.600 556.050 82.050 ;
        RECT 512.400 80.400 556.050 81.600 ;
        RECT 463.950 79.950 466.050 80.400 ;
        RECT 487.950 79.950 490.050 80.400 ;
        RECT 493.950 79.950 496.050 80.400 ;
        RECT 553.950 79.950 556.050 80.400 ;
        RECT 766.950 81.600 769.050 82.050 ;
        RECT 778.950 81.600 781.050 82.050 ;
        RECT 766.950 80.400 781.050 81.600 ;
        RECT 766.950 79.950 769.050 80.400 ;
        RECT 778.950 79.950 781.050 80.400 ;
        RECT 235.950 78.600 238.050 79.050 ;
        RECT 355.950 78.600 358.050 79.050 ;
        RECT 235.950 77.400 358.050 78.600 ;
        RECT 235.950 76.950 238.050 77.400 ;
        RECT 355.950 76.950 358.050 77.400 ;
        RECT 397.950 78.600 400.050 79.050 ;
        RECT 622.950 78.600 625.050 79.050 ;
        RECT 397.950 77.400 625.050 78.600 ;
        RECT 397.950 76.950 400.050 77.400 ;
        RECT 622.950 76.950 625.050 77.400 ;
        RECT 634.950 78.600 637.050 79.050 ;
        RECT 643.950 78.600 646.050 79.050 ;
        RECT 634.950 77.400 646.050 78.600 ;
        RECT 634.950 76.950 637.050 77.400 ;
        RECT 643.950 76.950 646.050 77.400 ;
        RECT 649.950 78.600 652.050 79.050 ;
        RECT 694.950 78.600 697.050 79.050 ;
        RECT 649.950 77.400 697.050 78.600 ;
        RECT 649.950 76.950 652.050 77.400 ;
        RECT 694.950 76.950 697.050 77.400 ;
        RECT 28.950 75.600 31.050 76.050 ;
        RECT 43.950 75.600 46.050 76.050 ;
        RECT 28.950 74.400 46.050 75.600 ;
        RECT 28.950 73.950 31.050 74.400 ;
        RECT 43.950 73.950 46.050 74.400 ;
        RECT 166.950 75.600 169.050 76.050 ;
        RECT 184.950 75.600 187.050 76.050 ;
        RECT 220.950 75.600 223.050 76.050 ;
        RECT 232.950 75.600 235.050 76.050 ;
        RECT 166.950 74.400 235.050 75.600 ;
        RECT 166.950 73.950 169.050 74.400 ;
        RECT 184.950 73.950 187.050 74.400 ;
        RECT 220.950 73.950 223.050 74.400 ;
        RECT 232.950 73.950 235.050 74.400 ;
        RECT 238.950 72.600 241.050 73.050 ;
        RECT 253.950 72.600 256.050 76.050 ;
        RECT 259.950 75.600 262.050 76.050 ;
        RECT 277.950 75.600 280.050 76.050 ;
        RECT 259.950 74.400 280.050 75.600 ;
        RECT 259.950 73.950 262.050 74.400 ;
        RECT 277.950 73.950 280.050 74.400 ;
        RECT 751.950 75.600 754.050 76.050 ;
        RECT 772.950 75.600 775.050 76.050 ;
        RECT 751.950 74.400 775.050 75.600 ;
        RECT 751.950 73.950 754.050 74.400 ;
        RECT 772.950 73.950 775.050 74.400 ;
        RECT 796.950 75.600 799.050 76.050 ;
        RECT 808.950 75.600 811.050 76.050 ;
        RECT 796.950 74.400 811.050 75.600 ;
        RECT 796.950 73.950 799.050 74.400 ;
        RECT 808.950 73.950 811.050 74.400 ;
        RECT 484.950 72.600 487.050 73.050 ;
        RECT 238.950 71.400 487.050 72.600 ;
        RECT 238.950 70.950 241.050 71.400 ;
        RECT 484.950 70.950 487.050 71.400 ;
        RECT 493.950 72.600 496.050 73.050 ;
        RECT 592.950 72.600 595.050 73.050 ;
        RECT 598.950 72.600 601.050 73.050 ;
        RECT 493.950 71.400 601.050 72.600 ;
        RECT 493.950 70.950 496.050 71.400 ;
        RECT 592.950 70.950 595.050 71.400 ;
        RECT 598.950 70.950 601.050 71.400 ;
        RECT 10.950 69.600 13.050 70.050 ;
        RECT 61.950 69.600 64.050 70.050 ;
        RECT 10.950 68.400 64.050 69.600 ;
        RECT 10.950 67.950 13.050 68.400 ;
        RECT 61.950 67.950 64.050 68.400 ;
        RECT 271.950 69.600 274.050 70.050 ;
        RECT 286.950 69.600 289.050 70.050 ;
        RECT 271.950 68.400 289.050 69.600 ;
        RECT 271.950 67.950 274.050 68.400 ;
        RECT 286.950 67.950 289.050 68.400 ;
        RECT 301.950 69.600 304.050 70.050 ;
        RECT 337.950 69.600 340.050 70.050 ;
        RECT 301.950 68.400 340.050 69.600 ;
        RECT 301.950 67.950 304.050 68.400 ;
        RECT 337.950 67.950 340.050 68.400 ;
        RECT 355.950 69.600 358.050 70.050 ;
        RECT 409.950 69.600 412.050 70.050 ;
        RECT 355.950 68.400 412.050 69.600 ;
        RECT 355.950 67.950 358.050 68.400 ;
        RECT 409.950 67.950 412.050 68.400 ;
        RECT 478.950 69.600 481.050 70.050 ;
        RECT 574.950 69.600 577.050 70.050 ;
        RECT 478.950 68.400 577.050 69.600 ;
        RECT 478.950 67.950 481.050 68.400 ;
        RECT 574.950 67.950 577.050 68.400 ;
        RECT 691.950 69.600 694.050 70.050 ;
        RECT 697.950 69.600 700.050 70.050 ;
        RECT 718.950 69.600 721.050 70.050 ;
        RECT 691.950 68.400 721.050 69.600 ;
        RECT 691.950 67.950 694.050 68.400 ;
        RECT 697.950 67.950 700.050 68.400 ;
        RECT 718.950 67.950 721.050 68.400 ;
        RECT 244.950 66.600 247.050 67.050 ;
        RECT 259.950 66.600 262.050 67.050 ;
        RECT 244.950 65.400 262.050 66.600 ;
        RECT 244.950 64.950 247.050 65.400 ;
        RECT 259.950 64.950 262.050 65.400 ;
        RECT 268.950 66.600 271.050 67.050 ;
        RECT 292.950 66.600 295.050 67.050 ;
        RECT 298.950 66.600 301.050 67.050 ;
        RECT 382.950 66.600 385.050 67.050 ;
        RECT 268.950 65.400 385.050 66.600 ;
        RECT 268.950 64.950 271.050 65.400 ;
        RECT 292.950 64.950 295.050 65.400 ;
        RECT 298.950 64.950 301.050 65.400 ;
        RECT 382.950 64.950 385.050 65.400 ;
        RECT 436.950 66.600 439.050 67.050 ;
        RECT 457.950 66.600 460.050 67.050 ;
        RECT 436.950 65.400 460.050 66.600 ;
        RECT 436.950 64.950 439.050 65.400 ;
        RECT 457.950 64.950 460.050 65.400 ;
        RECT 553.950 66.600 556.050 67.050 ;
        RECT 577.950 66.600 580.050 67.050 ;
        RECT 604.950 66.600 607.050 67.050 ;
        RECT 553.950 65.400 607.050 66.600 ;
        RECT 553.950 64.950 556.050 65.400 ;
        RECT 577.950 64.950 580.050 65.400 ;
        RECT 604.950 64.950 607.050 65.400 ;
        RECT 667.950 66.600 670.050 67.050 ;
        RECT 679.950 66.600 682.050 67.050 ;
        RECT 667.950 65.400 682.050 66.600 ;
        RECT 667.950 64.950 670.050 65.400 ;
        RECT 679.950 64.950 682.050 65.400 ;
        RECT 760.950 66.600 763.050 67.050 ;
        RECT 790.950 66.600 793.050 67.050 ;
        RECT 850.950 66.600 853.050 67.050 ;
        RECT 760.950 65.400 853.050 66.600 ;
        RECT 760.950 64.950 763.050 65.400 ;
        RECT 790.950 64.950 793.050 65.400 ;
        RECT 850.950 64.950 853.050 65.400 ;
        RECT 46.950 63.600 49.050 64.050 ;
        RECT 103.950 63.600 106.050 64.050 ;
        RECT 121.950 63.600 124.050 64.050 ;
        RECT 163.950 63.600 166.050 64.050 ;
        RECT 169.950 63.600 172.050 64.050 ;
        RECT 46.950 62.400 172.050 63.600 ;
        RECT 46.950 61.950 49.050 62.400 ;
        RECT 103.950 61.950 106.050 62.400 ;
        RECT 121.950 61.950 124.050 62.400 ;
        RECT 163.950 61.950 166.050 62.400 ;
        RECT 169.950 61.950 172.050 62.400 ;
        RECT 178.950 63.600 181.050 64.050 ;
        RECT 202.950 63.600 205.050 64.050 ;
        RECT 178.950 62.400 205.050 63.600 ;
        RECT 178.950 61.950 181.050 62.400 ;
        RECT 202.950 61.950 205.050 62.400 ;
        RECT 328.950 61.950 331.050 64.050 ;
        RECT 334.950 63.600 337.050 64.050 ;
        RECT 349.950 63.600 352.050 64.050 ;
        RECT 334.950 62.400 352.050 63.600 ;
        RECT 334.950 61.950 337.050 62.400 ;
        RECT 349.950 61.950 352.050 62.400 ;
        RECT 625.950 63.600 628.050 64.050 ;
        RECT 700.950 63.600 703.050 64.050 ;
        RECT 625.950 62.400 703.050 63.600 ;
        RECT 625.950 61.950 628.050 62.400 ;
        RECT 16.950 60.600 21.000 61.050 ;
        RECT 37.950 60.600 40.050 61.200 ;
        RECT 67.950 60.750 70.050 61.200 ;
        RECT 73.950 60.750 76.050 61.200 ;
        RECT 16.950 58.950 21.600 60.600 ;
        RECT 37.950 59.400 66.600 60.600 ;
        RECT 37.950 59.100 40.050 59.400 ;
        RECT 20.400 54.900 21.600 58.950 ;
        RECT 65.400 54.900 66.600 59.400 ;
        RECT 67.950 59.550 76.050 60.750 ;
        RECT 67.950 59.100 70.050 59.550 ;
        RECT 73.950 59.100 76.050 59.550 ;
        RECT 85.950 58.950 88.050 61.050 ;
        RECT 106.950 60.750 109.050 61.200 ;
        RECT 112.950 60.750 115.050 61.200 ;
        RECT 106.950 59.550 115.050 60.750 ;
        RECT 106.950 59.100 109.050 59.550 ;
        RECT 112.950 59.100 115.050 59.550 ;
        RECT 139.950 60.600 142.050 61.200 ;
        RECT 157.950 60.600 160.050 61.050 ;
        RECT 139.950 59.400 160.050 60.600 ;
        RECT 139.950 59.100 142.050 59.400 ;
        RECT 157.950 58.950 160.050 59.400 ;
        RECT 205.950 60.600 208.050 61.050 ;
        RECT 214.950 60.600 217.050 61.050 ;
        RECT 205.950 59.400 217.050 60.600 ;
        RECT 205.950 58.950 208.050 59.400 ;
        RECT 214.950 58.950 217.050 59.400 ;
        RECT 262.950 60.600 267.000 61.050 ;
        RECT 262.950 58.950 267.600 60.600 ;
        RECT 274.950 59.100 277.050 61.200 ;
        RECT 286.950 60.600 289.050 61.050 ;
        RECT 307.950 60.600 310.050 61.050 ;
        RECT 286.950 59.400 310.050 60.600 ;
        RECT 13.950 54.600 16.050 54.900 ;
        RECT 19.950 54.600 22.050 54.900 ;
        RECT 13.950 53.400 22.050 54.600 ;
        RECT 13.950 52.800 16.050 53.400 ;
        RECT 19.950 52.800 22.050 53.400 ;
        RECT 64.950 52.800 67.050 54.900 ;
        RECT 73.950 54.600 76.050 55.050 ;
        RECT 82.950 54.600 85.050 54.750 ;
        RECT 73.950 53.400 85.050 54.600 ;
        RECT 86.400 54.600 87.600 58.950 ;
        RECT 235.950 57.600 238.050 58.050 ;
        RECT 218.400 56.400 238.050 57.600 ;
        RECT 94.950 54.600 97.050 54.900 ;
        RECT 86.400 54.450 97.050 54.600 ;
        RECT 127.950 54.450 130.050 54.900 ;
        RECT 86.400 53.400 130.050 54.450 ;
        RECT 73.950 52.950 76.050 53.400 ;
        RECT 82.950 52.650 85.050 53.400 ;
        RECT 94.950 53.250 130.050 53.400 ;
        RECT 94.950 52.800 97.050 53.250 ;
        RECT 127.950 52.800 130.050 53.250 ;
        RECT 148.950 54.600 151.050 55.050 ;
        RECT 196.950 54.600 199.050 54.900 ;
        RECT 148.950 53.400 199.050 54.600 ;
        RECT 148.950 52.950 151.050 53.400 ;
        RECT 196.950 52.800 199.050 53.400 ;
        RECT 202.950 54.600 205.050 55.050 ;
        RECT 218.400 54.750 219.600 56.400 ;
        RECT 235.950 55.950 238.050 56.400 ;
        RECT 266.400 54.900 267.600 58.950 ;
        RECT 211.950 54.600 214.050 54.750 ;
        RECT 202.950 53.400 214.050 54.600 ;
        RECT 202.950 52.950 205.050 53.400 ;
        RECT 211.950 52.650 214.050 53.400 ;
        RECT 217.950 52.650 220.050 54.750 ;
        RECT 226.950 54.450 229.050 54.900 ;
        RECT 259.950 54.450 262.050 54.900 ;
        RECT 226.950 53.250 262.050 54.450 ;
        RECT 226.950 52.800 229.050 53.250 ;
        RECT 259.950 52.800 262.050 53.250 ;
        RECT 265.950 52.800 268.050 54.900 ;
        RECT 275.400 54.600 276.600 59.100 ;
        RECT 286.950 58.950 289.050 59.400 ;
        RECT 307.950 58.950 310.050 59.400 ;
        RECT 313.950 58.950 316.050 61.050 ;
        RECT 319.950 60.750 322.050 61.200 ;
        RECT 325.950 60.750 328.050 61.200 ;
        RECT 319.950 59.550 328.050 60.750 ;
        RECT 319.950 59.100 322.050 59.550 ;
        RECT 325.950 59.100 328.050 59.550 ;
        RECT 289.950 54.600 292.050 54.750 ;
        RECT 275.400 53.400 292.050 54.600 ;
        RECT 289.950 52.650 292.050 53.400 ;
        RECT 295.950 54.600 298.050 55.050 ;
        RECT 314.400 54.600 315.600 58.950 ;
        RECT 329.400 54.900 330.600 61.950 ;
        RECT 331.950 59.100 334.050 61.200 ;
        RECT 332.400 57.600 333.600 59.100 ;
        RECT 358.950 57.600 361.050 58.050 ;
        RECT 379.950 57.600 382.050 61.050 ;
        RECT 385.950 60.600 388.050 61.050 ;
        RECT 394.950 60.600 397.050 61.050 ;
        RECT 385.950 59.400 397.050 60.600 ;
        RECT 385.950 58.950 388.050 59.400 ;
        RECT 394.950 58.950 397.050 59.400 ;
        RECT 415.950 60.750 418.050 60.900 ;
        RECT 421.950 60.750 424.050 61.200 ;
        RECT 415.950 59.550 424.050 60.750 ;
        RECT 415.950 58.800 418.050 59.550 ;
        RECT 421.950 59.100 424.050 59.550 ;
        RECT 448.950 57.600 451.050 61.050 ;
        RECT 478.950 59.100 481.050 61.200 ;
        RECT 505.950 60.600 508.050 61.050 ;
        RECT 517.950 60.600 520.050 61.050 ;
        RECT 505.950 59.400 520.050 60.600 ;
        RECT 332.400 56.400 361.050 57.600 ;
        RECT 358.950 55.950 361.050 56.400 ;
        RECT 368.400 56.400 417.600 57.600 ;
        RECT 448.950 57.000 459.600 57.600 ;
        RECT 449.400 56.400 459.600 57.000 ;
        RECT 368.400 54.900 369.600 56.400 ;
        RECT 295.950 53.400 315.600 54.600 ;
        RECT 295.950 52.950 298.050 53.400 ;
        RECT 328.950 52.800 331.050 54.900 ;
        RECT 367.950 52.800 370.050 54.900 ;
        RECT 388.950 54.600 391.050 54.750 ;
        RECT 412.950 54.600 415.050 55.050 ;
        RECT 388.950 53.400 415.050 54.600 ;
        RECT 416.400 54.600 417.600 56.400 ;
        RECT 424.950 54.600 427.050 54.900 ;
        RECT 416.400 53.400 427.050 54.600 ;
        RECT 388.950 52.650 391.050 53.400 ;
        RECT 412.950 52.950 415.050 53.400 ;
        RECT 424.950 52.800 427.050 53.400 ;
        RECT 445.950 54.300 448.050 54.750 ;
        RECT 454.950 54.300 457.050 54.750 ;
        RECT 445.950 53.100 457.050 54.300 ;
        RECT 445.950 52.650 448.050 53.100 ;
        RECT 454.950 52.650 457.050 53.100 ;
        RECT 58.950 51.600 61.050 52.050 ;
        RECT 130.950 51.600 133.050 52.050 ;
        RECT 280.950 51.600 283.050 52.050 ;
        RECT 58.950 50.400 283.050 51.600 ;
        RECT 58.950 49.950 61.050 50.400 ;
        RECT 130.950 49.950 133.050 50.400 ;
        RECT 280.950 49.950 283.050 50.400 ;
        RECT 403.950 51.600 406.050 52.050 ;
        RECT 409.950 51.600 412.050 52.050 ;
        RECT 403.950 50.400 412.050 51.600 ;
        RECT 458.400 51.600 459.600 56.400 ;
        RECT 466.950 54.600 469.050 54.750 ;
        RECT 479.400 54.600 480.600 59.100 ;
        RECT 505.950 58.950 508.050 59.400 ;
        RECT 517.950 58.950 520.050 59.400 ;
        RECT 526.950 60.750 529.050 61.200 ;
        RECT 547.950 60.750 550.050 61.200 ;
        RECT 526.950 59.550 550.050 60.750 ;
        RECT 526.950 59.100 529.050 59.550 ;
        RECT 536.400 55.050 537.600 59.550 ;
        RECT 547.950 59.100 550.050 59.550 ;
        RECT 556.950 58.950 559.050 61.050 ;
        RECT 568.950 60.750 571.050 61.200 ;
        RECT 574.950 60.750 577.050 61.200 ;
        RECT 568.950 59.550 577.050 60.750 ;
        RECT 568.950 59.100 571.050 59.550 ;
        RECT 574.950 59.100 577.050 59.550 ;
        RECT 607.950 60.600 610.050 61.050 ;
        RECT 613.950 60.600 616.050 61.050 ;
        RECT 619.950 60.600 622.050 60.900 ;
        RECT 607.950 59.400 622.050 60.600 ;
        RECT 607.950 58.950 610.050 59.400 ;
        RECT 613.950 58.950 616.050 59.400 ;
        RECT 557.400 55.050 558.600 58.950 ;
        RECT 619.950 58.800 622.050 59.400 ;
        RECT 634.950 58.950 637.050 61.050 ;
        RECT 635.400 55.050 636.600 58.950 ;
        RECT 466.950 53.400 480.600 54.600 ;
        RECT 499.950 54.450 502.050 54.900 ;
        RECT 505.950 54.450 508.050 54.900 ;
        RECT 466.950 52.650 469.050 53.400 ;
        RECT 499.950 53.250 508.050 54.450 ;
        RECT 499.950 52.800 502.050 53.250 ;
        RECT 505.950 52.800 508.050 53.250 ;
        RECT 535.950 52.950 538.050 55.050 ;
        RECT 556.950 52.950 559.050 55.050 ;
        RECT 577.950 54.450 580.050 54.900 ;
        RECT 586.950 54.450 589.050 54.900 ;
        RECT 577.950 53.250 589.050 54.450 ;
        RECT 577.950 52.800 580.050 53.250 ;
        RECT 586.950 52.800 589.050 53.250 ;
        RECT 601.950 54.600 604.050 54.750 ;
        RECT 610.950 54.600 613.050 55.050 ;
        RECT 601.950 53.400 613.050 54.600 ;
        RECT 601.950 52.650 604.050 53.400 ;
        RECT 610.950 52.950 613.050 53.400 ;
        RECT 634.950 52.950 637.050 55.050 ;
        RECT 644.400 54.900 645.600 62.400 ;
        RECT 700.950 61.950 703.050 62.400 ;
        RECT 646.950 60.600 649.050 61.050 ;
        RECT 667.950 60.600 670.050 61.050 ;
        RECT 673.950 60.600 676.050 61.200 ;
        RECT 678.000 60.600 682.050 61.050 ;
        RECT 646.950 59.400 670.050 60.600 ;
        RECT 646.950 58.950 649.050 59.400 ;
        RECT 667.950 58.950 670.050 59.400 ;
        RECT 671.400 59.400 676.050 60.600 ;
        RECT 671.400 55.050 672.600 59.400 ;
        RECT 673.950 59.100 676.050 59.400 ;
        RECT 643.950 52.800 646.050 54.900 ;
        RECT 667.950 53.400 672.600 55.050 ;
        RECT 677.400 58.950 682.050 60.600 ;
        RECT 685.950 60.600 688.050 61.050 ;
        RECT 703.950 60.600 706.050 61.050 ;
        RECT 712.950 60.600 715.050 61.050 ;
        RECT 685.950 59.400 702.600 60.600 ;
        RECT 685.950 58.950 688.050 59.400 ;
        RECT 677.400 54.900 678.600 58.950 ;
        RECT 701.400 57.600 702.600 59.400 ;
        RECT 703.950 59.400 715.050 60.600 ;
        RECT 703.950 58.950 706.050 59.400 ;
        RECT 712.950 58.950 715.050 59.400 ;
        RECT 730.950 60.600 733.050 61.200 ;
        RECT 736.950 60.600 739.050 61.050 ;
        RECT 742.950 60.600 745.050 61.050 ;
        RECT 730.950 59.400 745.050 60.600 ;
        RECT 730.950 59.100 733.050 59.400 ;
        RECT 736.950 58.950 739.050 59.400 ;
        RECT 742.950 58.950 745.050 59.400 ;
        RECT 751.950 57.600 754.050 61.050 ;
        RECT 757.950 60.600 760.050 61.050 ;
        RECT 766.950 60.600 769.050 61.200 ;
        RECT 757.950 59.400 769.050 60.600 ;
        RECT 757.950 58.950 760.050 59.400 ;
        RECT 766.950 59.100 769.050 59.400 ;
        RECT 775.950 60.600 778.050 61.050 ;
        RECT 781.950 60.600 784.050 61.200 ;
        RECT 775.950 59.400 784.050 60.600 ;
        RECT 775.950 58.950 778.050 59.400 ;
        RECT 781.950 59.100 784.050 59.400 ;
        RECT 799.950 60.750 802.050 61.200 ;
        RECT 805.950 60.750 808.050 61.200 ;
        RECT 799.950 59.550 808.050 60.750 ;
        RECT 799.950 59.100 802.050 59.550 ;
        RECT 805.950 59.100 808.050 59.550 ;
        RECT 823.950 60.750 826.050 61.200 ;
        RECT 832.950 60.750 835.050 61.200 ;
        RECT 823.950 59.550 835.050 60.750 ;
        RECT 823.950 59.100 826.050 59.550 ;
        RECT 832.950 59.100 835.050 59.550 ;
        RECT 701.400 56.400 717.600 57.600 ;
        RECT 751.950 57.000 765.600 57.600 ;
        RECT 752.400 56.400 765.600 57.000 ;
        RECT 667.950 52.950 672.000 53.400 ;
        RECT 676.950 52.800 679.050 54.900 ;
        RECT 716.400 54.750 717.600 56.400 ;
        RECT 764.400 54.900 765.600 56.400 ;
        RECT 715.950 54.600 718.050 54.750 ;
        RECT 727.950 54.600 730.050 54.900 ;
        RECT 715.950 53.400 730.050 54.600 ;
        RECT 715.950 52.650 718.050 53.400 ;
        RECT 727.950 52.800 730.050 53.400 ;
        RECT 763.950 52.800 766.050 54.900 ;
        RECT 817.950 54.600 820.050 54.900 ;
        RECT 829.950 54.600 832.050 54.900 ;
        RECT 817.950 53.400 832.050 54.600 ;
        RECT 817.950 52.800 820.050 53.400 ;
        RECT 829.950 52.800 832.050 53.400 ;
        RECT 523.950 51.600 526.050 52.050 ;
        RECT 541.950 51.600 544.050 52.050 ;
        RECT 458.400 50.400 474.600 51.600 ;
        RECT 403.950 49.950 406.050 50.400 ;
        RECT 409.950 49.950 412.050 50.400 ;
        RECT 473.400 49.050 474.600 50.400 ;
        RECT 523.950 50.400 544.050 51.600 ;
        RECT 523.950 49.950 526.050 50.400 ;
        RECT 541.950 49.950 544.050 50.400 ;
        RECT 613.950 51.600 616.050 52.050 ;
        RECT 637.950 51.600 640.050 52.050 ;
        RECT 613.950 50.400 640.050 51.600 ;
        RECT 613.950 49.950 616.050 50.400 ;
        RECT 637.950 49.950 640.050 50.400 ;
        RECT 766.950 51.600 769.050 52.050 ;
        RECT 784.950 51.600 787.050 52.050 ;
        RECT 808.950 51.600 811.050 52.050 ;
        RECT 766.950 50.400 811.050 51.600 ;
        RECT 766.950 49.950 769.050 50.400 ;
        RECT 784.950 49.950 787.050 50.400 ;
        RECT 808.950 49.950 811.050 50.400 ;
        RECT 160.950 48.600 163.050 49.050 ;
        RECT 187.950 48.600 190.050 49.050 ;
        RECT 160.950 47.400 190.050 48.600 ;
        RECT 160.950 46.950 163.050 47.400 ;
        RECT 187.950 46.950 190.050 47.400 ;
        RECT 199.950 48.600 202.050 49.050 ;
        RECT 211.950 48.600 214.050 49.050 ;
        RECT 199.950 47.400 214.050 48.600 ;
        RECT 199.950 46.950 202.050 47.400 ;
        RECT 211.950 46.950 214.050 47.400 ;
        RECT 271.950 48.600 274.050 49.050 ;
        RECT 277.950 48.600 280.050 49.050 ;
        RECT 271.950 47.400 280.050 48.600 ;
        RECT 271.950 46.950 274.050 47.400 ;
        RECT 277.950 46.950 280.050 47.400 ;
        RECT 358.950 48.600 361.050 49.050 ;
        RECT 415.950 48.600 418.050 49.050 ;
        RECT 358.950 47.400 418.050 48.600 ;
        RECT 358.950 46.950 361.050 47.400 ;
        RECT 415.950 46.950 418.050 47.400 ;
        RECT 472.950 48.600 475.050 49.050 ;
        RECT 520.950 48.600 523.050 49.050 ;
        RECT 472.950 47.400 523.050 48.600 ;
        RECT 472.950 46.950 475.050 47.400 ;
        RECT 520.950 46.950 523.050 47.400 ;
        RECT 538.950 48.600 541.050 49.050 ;
        RECT 550.950 48.600 553.050 49.050 ;
        RECT 538.950 47.400 553.050 48.600 ;
        RECT 538.950 46.950 541.050 47.400 ;
        RECT 550.950 46.950 553.050 47.400 ;
        RECT 634.950 48.600 637.050 49.050 ;
        RECT 643.950 48.600 646.050 49.050 ;
        RECT 634.950 47.400 646.050 48.600 ;
        RECT 634.950 46.950 637.050 47.400 ;
        RECT 643.950 46.950 646.050 47.400 ;
        RECT 667.950 48.600 670.050 49.050 ;
        RECT 694.950 48.600 697.050 49.050 ;
        RECT 703.950 48.600 706.050 49.050 ;
        RECT 667.950 47.400 706.050 48.600 ;
        RECT 809.400 48.600 810.600 49.950 ;
        RECT 850.950 48.600 853.050 49.050 ;
        RECT 809.400 47.400 853.050 48.600 ;
        RECT 667.950 46.950 670.050 47.400 ;
        RECT 694.950 46.950 697.050 47.400 ;
        RECT 703.950 46.950 706.050 47.400 ;
        RECT 850.950 46.950 853.050 47.400 ;
        RECT 106.950 45.600 109.050 46.050 ;
        RECT 154.950 45.600 157.050 46.050 ;
        RECT 106.950 44.400 157.050 45.600 ;
        RECT 106.950 43.950 109.050 44.400 ;
        RECT 154.950 43.950 157.050 44.400 ;
        RECT 301.950 45.600 304.050 46.050 ;
        RECT 319.950 45.600 322.050 46.050 ;
        RECT 442.950 45.600 445.050 46.050 ;
        RECT 301.950 44.400 322.050 45.600 ;
        RECT 301.950 43.950 304.050 44.400 ;
        RECT 319.950 43.950 322.050 44.400 ;
        RECT 392.400 44.400 445.050 45.600 ;
        RECT 355.950 42.600 358.050 43.050 ;
        RECT 367.950 42.600 370.050 43.050 ;
        RECT 392.400 42.600 393.600 44.400 ;
        RECT 442.950 43.950 445.050 44.400 ;
        RECT 448.950 45.600 451.050 46.050 ;
        RECT 523.950 45.600 526.050 46.050 ;
        RECT 448.950 44.400 526.050 45.600 ;
        RECT 448.950 43.950 451.050 44.400 ;
        RECT 523.950 43.950 526.050 44.400 ;
        RECT 529.950 45.600 532.050 46.050 ;
        RECT 574.950 45.600 577.050 46.050 ;
        RECT 529.950 44.400 577.050 45.600 ;
        RECT 529.950 43.950 532.050 44.400 ;
        RECT 574.950 43.950 577.050 44.400 ;
        RECT 355.950 41.400 393.600 42.600 ;
        RECT 394.950 42.600 397.050 43.050 ;
        RECT 406.950 42.600 409.050 43.050 ;
        RECT 439.950 42.600 442.050 43.050 ;
        RECT 394.950 41.400 442.050 42.600 ;
        RECT 355.950 40.950 358.050 41.400 ;
        RECT 367.950 40.950 370.050 41.400 ;
        RECT 394.950 40.950 397.050 41.400 ;
        RECT 406.950 40.950 409.050 41.400 ;
        RECT 439.950 40.950 442.050 41.400 ;
        RECT 454.950 42.600 457.050 43.050 ;
        RECT 460.950 42.600 463.050 43.050 ;
        RECT 454.950 41.400 463.050 42.600 ;
        RECT 454.950 40.950 457.050 41.400 ;
        RECT 460.950 40.950 463.050 41.400 ;
        RECT 622.950 42.600 625.050 43.050 ;
        RECT 748.950 42.600 751.050 43.050 ;
        RECT 622.950 41.400 751.050 42.600 ;
        RECT 622.950 40.950 625.050 41.400 ;
        RECT 748.950 40.950 751.050 41.400 ;
        RECT 763.950 42.600 766.050 43.050 ;
        RECT 844.950 42.600 847.050 43.050 ;
        RECT 763.950 41.400 847.050 42.600 ;
        RECT 763.950 40.950 766.050 41.400 ;
        RECT 844.950 40.950 847.050 41.400 ;
        RECT 334.950 39.600 337.050 40.050 ;
        RECT 364.950 39.600 367.050 40.050 ;
        RECT 334.950 38.400 367.050 39.600 ;
        RECT 334.950 37.950 337.050 38.400 ;
        RECT 364.950 37.950 367.050 38.400 ;
        RECT 457.950 39.600 460.050 40.050 ;
        RECT 487.950 39.600 490.050 40.050 ;
        RECT 457.950 38.400 490.050 39.600 ;
        RECT 457.950 37.950 460.050 38.400 ;
        RECT 487.950 37.950 490.050 38.400 ;
        RECT 520.950 39.600 523.050 40.050 ;
        RECT 535.950 39.600 538.050 40.050 ;
        RECT 520.950 38.400 538.050 39.600 ;
        RECT 520.950 37.950 523.050 38.400 ;
        RECT 535.950 37.950 538.050 38.400 ;
        RECT 556.950 39.600 559.050 40.050 ;
        RECT 562.950 39.600 565.050 40.050 ;
        RECT 556.950 38.400 565.050 39.600 ;
        RECT 556.950 37.950 559.050 38.400 ;
        RECT 562.950 37.950 565.050 38.400 ;
        RECT 631.950 39.600 634.050 40.050 ;
        RECT 652.950 39.600 655.050 40.050 ;
        RECT 631.950 38.400 655.050 39.600 ;
        RECT 631.950 37.950 634.050 38.400 ;
        RECT 652.950 37.950 655.050 38.400 ;
        RECT 700.950 39.600 703.050 40.050 ;
        RECT 730.950 39.600 733.050 40.050 ;
        RECT 700.950 38.400 733.050 39.600 ;
        RECT 700.950 37.950 703.050 38.400 ;
        RECT 730.950 37.950 733.050 38.400 ;
        RECT 805.950 39.600 808.050 40.050 ;
        RECT 817.950 39.600 820.050 40.050 ;
        RECT 805.950 38.400 820.050 39.600 ;
        RECT 805.950 37.950 808.050 38.400 ;
        RECT 817.950 37.950 820.050 38.400 ;
        RECT 160.950 36.600 163.050 37.050 ;
        RECT 238.950 36.600 241.050 37.050 ;
        RECT 160.950 35.400 241.050 36.600 ;
        RECT 160.950 34.950 163.050 35.400 ;
        RECT 238.950 34.950 241.050 35.400 ;
        RECT 295.950 36.600 298.050 37.050 ;
        RECT 335.400 36.600 336.600 37.950 ;
        RECT 295.950 35.400 336.600 36.600 ;
        RECT 403.950 36.600 406.050 37.050 ;
        RECT 412.950 36.600 415.050 37.050 ;
        RECT 508.950 36.600 511.050 37.050 ;
        RECT 403.950 35.400 511.050 36.600 ;
        RECT 295.950 34.950 298.050 35.400 ;
        RECT 403.950 34.950 406.050 35.400 ;
        RECT 412.950 34.950 415.050 35.400 ;
        RECT 508.950 34.950 511.050 35.400 ;
        RECT 592.950 36.600 595.050 37.050 ;
        RECT 598.950 36.600 601.050 37.050 ;
        RECT 592.950 35.400 601.050 36.600 ;
        RECT 592.950 34.950 595.050 35.400 ;
        RECT 598.950 34.950 601.050 35.400 ;
        RECT 52.950 33.600 55.050 34.050 ;
        RECT 64.950 33.600 67.050 34.050 ;
        RECT 52.950 32.400 67.050 33.600 ;
        RECT 52.950 31.950 55.050 32.400 ;
        RECT 64.950 31.950 67.050 32.400 ;
        RECT 259.950 33.600 262.050 34.050 ;
        RECT 298.950 33.600 301.050 34.050 ;
        RECT 259.950 32.400 301.050 33.600 ;
        RECT 259.950 31.950 262.050 32.400 ;
        RECT 298.950 31.950 301.050 32.400 ;
        RECT 427.950 33.600 430.050 34.050 ;
        RECT 448.950 33.600 451.050 34.050 ;
        RECT 427.950 32.400 451.050 33.600 ;
        RECT 427.950 31.950 430.050 32.400 ;
        RECT 448.950 31.950 451.050 32.400 ;
        RECT 490.950 33.600 493.050 34.050 ;
        RECT 517.950 33.600 520.050 34.050 ;
        RECT 490.950 32.400 520.050 33.600 ;
        RECT 490.950 31.950 493.050 32.400 ;
        RECT 517.950 31.950 520.050 32.400 ;
        RECT 538.950 33.600 541.050 34.050 ;
        RECT 712.950 33.600 715.050 34.050 ;
        RECT 538.950 32.400 715.050 33.600 ;
        RECT 538.950 31.950 541.050 32.400 ;
        RECT 712.950 31.950 715.050 32.400 ;
        RECT 718.950 33.600 721.050 34.050 ;
        RECT 748.950 33.600 751.050 34.050 ;
        RECT 766.950 33.600 769.050 34.050 ;
        RECT 718.950 32.400 751.050 33.600 ;
        RECT 718.950 31.950 721.050 32.400 ;
        RECT 748.950 31.950 751.050 32.400 ;
        RECT 752.400 32.400 769.050 33.600 ;
        RECT 142.950 30.600 145.050 31.050 ;
        RECT 184.950 30.600 187.050 31.050 ;
        RECT 217.950 30.600 220.050 31.050 ;
        RECT 280.950 30.600 283.050 31.050 ;
        RECT 142.950 29.400 220.050 30.600 ;
        RECT 142.950 28.950 145.050 29.400 ;
        RECT 184.950 28.950 187.050 29.400 ;
        RECT 217.950 28.950 220.050 29.400 ;
        RECT 275.400 29.400 283.050 30.600 ;
        RECT 4.950 27.750 7.050 28.200 ;
        RECT 13.950 27.750 16.050 28.200 ;
        RECT 4.950 27.600 16.050 27.750 ;
        RECT 19.950 27.600 22.050 28.200 ;
        RECT 4.950 26.550 22.050 27.600 ;
        RECT 4.950 26.100 7.050 26.550 ;
        RECT 13.950 26.400 22.050 26.550 ;
        RECT 13.950 26.100 16.050 26.400 ;
        RECT 19.950 26.100 22.050 26.400 ;
        RECT 58.950 27.600 61.050 28.200 ;
        RECT 73.950 27.600 76.050 28.050 ;
        RECT 82.950 27.600 85.050 28.350 ;
        RECT 58.950 26.400 72.600 27.600 ;
        RECT 58.950 26.100 61.050 26.400 ;
        RECT 71.400 24.600 72.600 26.400 ;
        RECT 73.950 26.400 85.050 27.600 ;
        RECT 73.950 25.950 76.050 26.400 ;
        RECT 82.950 26.250 85.050 26.400 ;
        RECT 94.950 26.100 97.050 28.200 ;
        RECT 106.950 27.600 109.050 28.050 ;
        RECT 127.950 27.600 130.050 28.050 ;
        RECT 136.950 27.600 139.050 28.200 ;
        RECT 106.950 26.400 130.050 27.600 ;
        RECT 95.400 24.600 96.600 26.100 ;
        RECT 106.950 25.950 109.050 26.400 ;
        RECT 127.950 25.950 130.050 26.400 ;
        RECT 131.400 26.400 139.050 27.600 ;
        RECT 131.400 24.600 132.600 26.400 ;
        RECT 136.950 26.100 139.050 26.400 ;
        RECT 148.950 27.600 151.050 28.050 ;
        RECT 154.950 27.600 157.050 28.350 ;
        RECT 148.950 26.400 157.050 27.600 ;
        RECT 148.950 25.950 151.050 26.400 ;
        RECT 154.950 26.250 157.050 26.400 ;
        RECT 196.950 27.750 199.050 28.200 ;
        RECT 202.950 27.750 205.050 28.200 ;
        RECT 196.950 26.550 205.050 27.750 ;
        RECT 196.950 26.100 199.050 26.550 ;
        RECT 202.950 26.100 205.050 26.550 ;
        RECT 223.950 27.600 226.050 28.050 ;
        RECT 232.950 27.600 235.050 28.200 ;
        RECT 250.950 27.600 253.050 28.350 ;
        RECT 223.950 26.400 235.050 27.600 ;
        RECT 223.950 25.950 226.050 26.400 ;
        RECT 232.950 26.100 235.050 26.400 ;
        RECT 236.400 26.400 253.050 27.600 ;
        RECT 236.400 24.600 237.600 26.400 ;
        RECT 250.950 26.250 253.050 26.400 ;
        RECT 71.400 24.000 81.600 24.600 ;
        RECT 86.400 24.000 132.600 24.600 ;
        RECT 71.400 23.400 82.050 24.000 ;
        RECT 10.950 21.450 13.050 21.900 ;
        RECT 28.950 21.450 31.050 21.900 ;
        RECT 10.950 20.250 31.050 21.450 ;
        RECT 10.950 19.800 13.050 20.250 ;
        RECT 28.950 19.800 31.050 20.250 ;
        RECT 37.950 21.600 40.050 21.900 ;
        RECT 52.950 21.600 55.050 22.050 ;
        RECT 37.950 20.400 55.050 21.600 ;
        RECT 37.950 19.800 40.050 20.400 ;
        RECT 52.950 19.950 55.050 20.400 ;
        RECT 67.950 21.450 70.050 21.900 ;
        RECT 73.950 21.450 76.050 21.900 ;
        RECT 67.950 20.250 76.050 21.450 ;
        RECT 67.950 19.800 70.050 20.250 ;
        RECT 73.950 19.800 76.050 20.250 ;
        RECT 79.950 19.950 82.050 23.400 ;
        RECT 85.950 23.400 132.600 24.000 ;
        RECT 230.400 23.400 237.600 24.600 ;
        RECT 85.950 19.950 88.050 23.400 ;
        RECT 106.950 21.450 109.050 21.900 ;
        RECT 112.950 21.450 115.050 21.900 ;
        RECT 106.950 20.250 115.050 21.450 ;
        RECT 106.950 19.800 109.050 20.250 ;
        RECT 112.950 19.800 115.050 20.250 ;
        RECT 127.950 21.600 130.050 22.050 ;
        RECT 148.800 21.600 150.900 22.050 ;
        RECT 127.950 20.400 150.900 21.600 ;
        RECT 127.950 19.950 130.050 20.400 ;
        RECT 148.800 19.950 150.900 20.400 ;
        RECT 151.950 21.600 154.050 22.050 ;
        RECT 157.950 21.600 160.050 22.050 ;
        RECT 230.400 21.900 231.600 23.400 ;
        RECT 275.400 22.050 276.600 29.400 ;
        RECT 280.950 28.950 283.050 29.400 ;
        RECT 340.950 30.600 343.050 31.050 ;
        RECT 382.950 30.600 385.050 31.050 ;
        RECT 340.950 29.400 385.050 30.600 ;
        RECT 340.950 28.950 343.050 29.400 ;
        RECT 382.950 28.950 385.050 29.400 ;
        RECT 466.950 30.600 469.050 31.050 ;
        RECT 475.950 30.600 478.050 31.050 ;
        RECT 466.950 29.400 478.050 30.600 ;
        RECT 466.950 28.950 469.050 29.400 ;
        RECT 475.950 28.950 478.050 29.400 ;
        RECT 484.950 28.950 487.050 31.050 ;
        RECT 520.950 28.950 523.050 31.050 ;
        RECT 289.950 26.100 292.050 28.200 ;
        RECT 328.950 27.600 331.050 28.200 ;
        RECT 340.950 27.600 343.050 28.200 ;
        RECT 328.950 26.400 343.050 27.600 ;
        RECT 328.950 26.100 331.050 26.400 ;
        RECT 340.950 26.100 343.050 26.400 ;
        RECT 397.950 27.600 400.050 28.200 ;
        RECT 415.950 27.600 418.050 28.050 ;
        RECT 421.950 27.600 424.050 28.200 ;
        RECT 397.950 26.400 424.050 27.600 ;
        RECT 397.950 26.100 400.050 26.400 ;
        RECT 290.400 24.600 291.600 26.100 ;
        RECT 415.950 25.950 418.050 26.400 ;
        RECT 421.950 26.100 424.050 26.400 ;
        RECT 364.950 24.600 367.050 25.050 ;
        RECT 451.950 24.600 454.050 28.050 ;
        RECT 485.400 24.600 486.600 28.950 ;
        RECT 499.950 27.600 502.050 28.350 ;
        RECT 499.950 26.400 516.600 27.600 ;
        RECT 499.950 26.250 502.050 26.400 ;
        RECT 290.400 23.400 294.600 24.600 ;
        RECT 151.950 20.400 160.050 21.600 ;
        RECT 151.950 19.950 154.050 20.400 ;
        RECT 157.950 19.950 160.050 20.400 ;
        RECT 178.950 21.450 181.050 21.900 ;
        RECT 223.950 21.450 226.050 21.900 ;
        RECT 178.950 20.250 226.050 21.450 ;
        RECT 178.950 19.800 181.050 20.250 ;
        RECT 223.950 19.800 226.050 20.250 ;
        RECT 229.950 19.800 232.050 21.900 ;
        RECT 247.950 21.600 250.050 22.050 ;
        RECT 268.950 21.600 271.050 22.050 ;
        RECT 247.950 20.400 271.050 21.600 ;
        RECT 247.950 19.950 250.050 20.400 ;
        RECT 268.950 19.950 271.050 20.400 ;
        RECT 274.950 19.950 277.050 22.050 ;
        RECT 280.950 21.450 283.050 21.900 ;
        RECT 286.950 21.450 289.050 21.900 ;
        RECT 280.950 20.250 289.050 21.450 ;
        RECT 293.400 21.600 294.600 23.400 ;
        RECT 364.950 23.400 408.600 24.600 ;
        RECT 364.950 22.950 367.050 23.400 ;
        RECT 298.800 21.600 300.900 22.050 ;
        RECT 293.400 20.400 300.900 21.600 ;
        RECT 280.950 19.800 283.050 20.250 ;
        RECT 286.950 19.800 289.050 20.250 ;
        RECT 298.800 19.950 300.900 20.400 ;
        RECT 301.950 21.450 304.050 21.900 ;
        RECT 319.950 21.450 322.050 21.900 ;
        RECT 301.950 20.250 322.050 21.450 ;
        RECT 301.950 19.800 304.050 20.250 ;
        RECT 319.950 19.800 322.050 20.250 ;
        RECT 367.950 21.600 370.050 22.050 ;
        RECT 373.950 21.600 376.050 21.900 ;
        RECT 367.950 20.400 376.050 21.600 ;
        RECT 367.950 19.950 370.050 20.400 ;
        RECT 373.950 19.800 376.050 20.400 ;
        RECT 394.950 21.450 397.050 21.900 ;
        RECT 403.950 21.450 406.050 21.900 ;
        RECT 394.950 20.250 406.050 21.450 ;
        RECT 407.400 21.600 408.600 23.400 ;
        RECT 440.400 24.000 454.050 24.600 ;
        RECT 440.400 23.400 453.600 24.000 ;
        RECT 482.400 23.400 486.600 24.600 ;
        RECT 440.400 21.900 441.600 23.400 ;
        RECT 482.400 21.900 483.600 23.400 ;
        RECT 515.400 21.900 516.600 26.400 ;
        RECT 521.400 21.900 522.600 28.950 ;
        RECT 529.950 27.600 532.050 28.200 ;
        RECT 565.950 27.600 568.050 28.050 ;
        RECT 529.950 26.400 568.050 27.600 ;
        RECT 529.950 26.100 532.050 26.400 ;
        RECT 530.400 22.050 531.600 26.100 ;
        RECT 565.950 25.950 568.050 26.400 ;
        RECT 574.950 27.600 577.050 28.350 ;
        RECT 580.950 27.600 583.050 31.050 ;
        RECT 752.400 30.600 753.600 32.400 ;
        RECT 766.950 31.950 769.050 32.400 ;
        RECT 772.950 33.600 775.050 34.050 ;
        RECT 814.950 33.600 817.050 34.050 ;
        RECT 826.950 33.600 829.050 34.050 ;
        RECT 772.950 32.400 810.600 33.600 ;
        RECT 772.950 31.950 775.050 32.400 ;
        RECT 749.400 29.400 753.600 30.600 ;
        RECT 809.400 30.600 810.600 32.400 ;
        RECT 814.950 32.400 829.050 33.600 ;
        RECT 814.950 31.950 817.050 32.400 ;
        RECT 826.950 31.950 829.050 32.400 ;
        RECT 829.950 30.600 832.050 31.050 ;
        RECT 809.400 29.400 832.050 30.600 ;
        RECT 574.950 27.000 583.050 27.600 ;
        RECT 583.950 27.750 586.050 28.200 ;
        RECT 592.950 27.750 595.050 28.200 ;
        RECT 574.950 26.400 582.600 27.000 ;
        RECT 583.950 26.550 595.050 27.750 ;
        RECT 598.950 27.600 601.050 28.200 ;
        RECT 574.950 26.250 577.050 26.400 ;
        RECT 583.950 26.100 586.050 26.550 ;
        RECT 592.950 26.100 595.050 26.550 ;
        RECT 596.400 26.400 601.050 27.600 ;
        RECT 596.400 24.600 597.600 26.400 ;
        RECT 598.950 26.100 601.050 26.400 ;
        RECT 631.950 27.600 634.050 28.200 ;
        RECT 661.950 27.600 664.050 28.200 ;
        RECT 676.950 27.600 679.050 28.200 ;
        RECT 631.950 26.400 679.050 27.600 ;
        RECT 631.950 26.100 634.050 26.400 ;
        RECT 661.950 26.100 664.050 26.400 ;
        RECT 676.950 26.100 679.050 26.400 ;
        RECT 700.950 27.750 703.050 28.200 ;
        RECT 709.950 27.750 712.050 28.200 ;
        RECT 700.950 26.550 712.050 27.750 ;
        RECT 700.950 26.100 703.050 26.550 ;
        RECT 709.950 26.100 712.050 26.550 ;
        RECT 739.950 27.750 742.050 28.200 ;
        RECT 745.950 27.750 748.050 28.200 ;
        RECT 739.950 26.550 748.050 27.750 ;
        RECT 739.950 26.100 742.050 26.550 ;
        RECT 745.950 26.100 748.050 26.550 ;
        RECT 749.400 24.600 750.600 29.400 ;
        RECT 760.950 27.600 763.050 27.900 ;
        RECT 769.950 27.600 772.050 28.200 ;
        RECT 778.950 27.600 781.050 28.050 ;
        RECT 760.950 26.400 772.050 27.600 ;
        RECT 760.950 25.800 763.050 26.400 ;
        RECT 769.950 26.100 772.050 26.400 ;
        RECT 773.400 26.400 781.050 27.600 ;
        RECT 578.400 24.000 597.600 24.600 ;
        RECT 722.400 24.000 750.600 24.600 ;
        RECT 430.950 21.600 433.050 21.900 ;
        RECT 407.400 20.400 433.050 21.600 ;
        RECT 394.950 19.800 397.050 20.250 ;
        RECT 403.950 19.800 406.050 20.250 ;
        RECT 430.950 19.800 433.050 20.400 ;
        RECT 439.950 19.800 442.050 21.900 ;
        RECT 481.950 19.800 484.050 21.900 ;
        RECT 514.950 19.800 517.050 21.900 ;
        RECT 520.950 19.800 523.050 21.900 ;
        RECT 526.950 20.400 531.600 22.050 ;
        RECT 577.950 23.400 597.600 24.000 ;
        RECT 721.950 23.400 750.600 24.000 ;
        RECT 556.950 21.450 559.050 21.900 ;
        RECT 562.950 21.450 565.050 21.900 ;
        RECT 526.950 19.950 531.000 20.400 ;
        RECT 556.950 20.250 565.050 21.450 ;
        RECT 556.950 19.800 559.050 20.250 ;
        RECT 562.950 19.800 565.050 20.250 ;
        RECT 577.950 19.950 580.050 23.400 ;
        RECT 595.950 21.600 598.050 21.900 ;
        RECT 664.950 21.600 667.050 21.900 ;
        RECT 595.950 21.450 667.050 21.600 ;
        RECT 670.950 21.450 673.050 21.900 ;
        RECT 595.950 20.400 673.050 21.450 ;
        RECT 595.950 19.800 598.050 20.400 ;
        RECT 664.950 20.250 673.050 20.400 ;
        RECT 664.950 19.800 667.050 20.250 ;
        RECT 670.950 19.800 673.050 20.250 ;
        RECT 679.950 21.600 682.050 21.900 ;
        RECT 688.950 21.600 691.050 22.050 ;
        RECT 679.950 20.400 691.050 21.600 ;
        RECT 679.950 19.800 682.050 20.400 ;
        RECT 688.950 19.950 691.050 20.400 ;
        RECT 697.950 21.600 700.050 21.900 ;
        RECT 715.950 21.600 718.050 22.050 ;
        RECT 697.950 20.400 718.050 21.600 ;
        RECT 697.950 19.800 700.050 20.400 ;
        RECT 715.950 19.950 718.050 20.400 ;
        RECT 721.950 19.950 724.050 23.400 ;
        RECT 733.950 21.600 736.050 21.900 ;
        RECT 739.950 21.600 742.050 22.050 ;
        RECT 733.950 20.400 742.050 21.600 ;
        RECT 733.950 19.800 736.050 20.400 ;
        RECT 739.950 19.950 742.050 20.400 ;
        RECT 748.950 21.600 751.050 21.900 ;
        RECT 757.950 21.600 760.050 22.050 ;
        RECT 773.400 21.900 774.600 26.400 ;
        RECT 778.950 25.950 781.050 26.400 ;
        RECT 787.950 27.600 790.050 28.200 ;
        RECT 799.950 27.900 802.050 28.350 ;
        RECT 808.950 27.900 811.050 28.350 ;
        RECT 799.950 27.600 811.050 27.900 ;
        RECT 787.950 26.700 811.050 27.600 ;
        RECT 787.950 26.400 802.050 26.700 ;
        RECT 787.950 26.100 790.050 26.400 ;
        RECT 799.950 26.250 802.050 26.400 ;
        RECT 808.950 26.250 811.050 26.700 ;
        RECT 815.400 22.050 816.600 29.400 ;
        RECT 829.950 28.950 832.050 29.400 ;
        RECT 748.950 20.400 760.050 21.600 ;
        RECT 46.950 18.600 49.050 19.050 ;
        RECT 103.950 18.600 106.050 19.050 ;
        RECT 121.950 18.600 124.050 19.050 ;
        RECT 169.950 18.600 172.050 19.050 ;
        RECT 46.950 17.400 172.050 18.600 ;
        RECT 46.950 16.950 49.050 17.400 ;
        RECT 103.950 16.950 106.050 17.400 ;
        RECT 121.950 16.950 124.050 17.400 ;
        RECT 169.950 16.950 172.050 17.400 ;
        RECT 205.950 18.600 208.050 19.050 ;
        RECT 214.950 18.600 217.050 19.050 ;
        RECT 205.950 17.400 217.050 18.600 ;
        RECT 205.950 16.950 208.050 17.400 ;
        RECT 214.950 16.950 217.050 17.400 ;
        RECT 235.950 18.600 238.050 19.050 ;
        RECT 253.950 18.600 256.050 19.050 ;
        RECT 235.950 17.400 256.050 18.600 ;
        RECT 404.400 18.600 405.600 19.800 ;
        RECT 424.950 18.600 427.050 19.050 ;
        RECT 404.400 17.400 427.050 18.600 ;
        RECT 235.950 16.950 238.050 17.400 ;
        RECT 253.950 16.950 256.050 17.400 ;
        RECT 424.950 16.950 427.050 17.400 ;
        RECT 496.950 18.600 499.050 19.050 ;
        RECT 520.950 18.600 523.050 19.050 ;
        RECT 496.950 17.400 523.050 18.600 ;
        RECT 563.400 18.600 564.600 19.800 ;
        RECT 604.950 18.600 607.050 19.050 ;
        RECT 563.400 17.400 607.050 18.600 ;
        RECT 740.400 18.600 741.600 19.950 ;
        RECT 748.950 19.800 751.050 20.400 ;
        RECT 757.950 19.950 760.050 20.400 ;
        RECT 772.950 19.800 775.050 21.900 ;
        RECT 814.950 19.950 817.050 22.050 ;
        RECT 820.950 21.600 823.050 22.050 ;
        RECT 826.950 21.600 829.050 22.050 ;
        RECT 820.950 20.400 829.050 21.600 ;
        RECT 820.950 19.950 823.050 20.400 ;
        RECT 826.950 19.950 829.050 20.400 ;
        RECT 799.950 18.600 802.050 19.050 ;
        RECT 740.400 17.400 802.050 18.600 ;
        RECT 496.950 16.950 499.050 17.400 ;
        RECT 520.950 16.950 523.050 17.400 ;
        RECT 604.950 16.950 607.050 17.400 ;
        RECT 799.950 16.950 802.050 17.400 ;
        RECT 823.950 18.600 826.050 19.050 ;
        RECT 832.950 18.600 835.050 19.050 ;
        RECT 823.950 17.400 835.050 18.600 ;
        RECT 823.950 16.950 826.050 17.400 ;
        RECT 832.950 16.950 835.050 17.400 ;
        RECT 202.950 15.600 205.050 16.050 ;
        RECT 232.950 15.600 235.050 16.050 ;
        RECT 202.950 14.400 235.050 15.600 ;
        RECT 202.950 13.950 205.050 14.400 ;
        RECT 232.950 13.950 235.050 14.400 ;
        RECT 238.950 15.600 241.050 16.050 ;
        RECT 247.950 15.600 250.050 16.050 ;
        RECT 238.950 14.400 250.050 15.600 ;
        RECT 238.950 13.950 241.050 14.400 ;
        RECT 247.950 13.950 250.050 14.400 ;
        RECT 292.950 15.600 295.050 16.050 ;
        RECT 343.950 15.600 346.050 16.050 ;
        RECT 361.950 15.600 364.050 16.050 ;
        RECT 292.950 14.400 364.050 15.600 ;
        RECT 292.950 13.950 295.050 14.400 ;
        RECT 343.950 13.950 346.050 14.400 ;
        RECT 361.950 13.950 364.050 14.400 ;
        RECT 373.950 15.600 376.050 16.050 ;
        RECT 388.950 15.600 391.050 16.050 ;
        RECT 373.950 14.400 391.050 15.600 ;
        RECT 373.950 13.950 376.050 14.400 ;
        RECT 388.950 13.950 391.050 14.400 ;
        RECT 508.950 15.600 511.050 16.050 ;
        RECT 517.950 15.600 520.050 16.050 ;
        RECT 508.950 14.400 520.050 15.600 ;
        RECT 508.950 13.950 511.050 14.400 ;
        RECT 517.950 13.950 520.050 14.400 ;
        RECT 523.950 15.600 526.050 16.050 ;
        RECT 538.950 15.600 541.050 16.050 ;
        RECT 523.950 14.400 541.050 15.600 ;
        RECT 523.950 13.950 526.050 14.400 ;
        RECT 538.950 13.950 541.050 14.400 ;
        RECT 742.950 15.600 745.050 16.050 ;
        RECT 766.950 15.600 769.050 16.050 ;
        RECT 742.950 14.400 769.050 15.600 ;
        RECT 742.950 13.950 745.050 14.400 ;
        RECT 766.950 13.950 769.050 14.400 ;
        RECT 793.950 15.600 796.050 16.050 ;
        RECT 808.950 15.600 811.050 16.050 ;
        RECT 793.950 14.400 811.050 15.600 ;
        RECT 793.950 13.950 796.050 14.400 ;
        RECT 808.950 13.950 811.050 14.400 ;
        RECT 814.950 15.600 817.050 16.050 ;
        RECT 838.950 15.600 841.050 16.050 ;
        RECT 814.950 14.400 841.050 15.600 ;
        RECT 814.950 13.950 817.050 14.400 ;
        RECT 838.950 13.950 841.050 14.400 ;
        RECT 28.950 12.600 31.050 13.050 ;
        RECT 61.950 12.600 64.050 13.050 ;
        RECT 28.950 11.400 64.050 12.600 ;
        RECT 28.950 10.950 31.050 11.400 ;
        RECT 61.950 10.950 64.050 11.400 ;
        RECT 163.950 12.600 166.050 13.050 ;
        RECT 184.950 12.600 187.050 13.050 ;
        RECT 163.950 11.400 187.050 12.600 ;
        RECT 163.950 10.950 166.050 11.400 ;
        RECT 184.950 10.950 187.050 11.400 ;
        RECT 298.950 12.600 301.050 13.050 ;
        RECT 310.950 12.600 313.050 13.050 ;
        RECT 472.950 12.600 475.050 13.050 ;
        RECT 298.950 11.400 313.050 12.600 ;
        RECT 298.950 10.950 301.050 11.400 ;
        RECT 310.950 10.950 313.050 11.400 ;
        RECT 413.400 11.400 475.050 12.600 ;
        RECT 358.950 9.600 361.050 10.050 ;
        RECT 413.400 9.600 414.600 11.400 ;
        RECT 472.950 10.950 475.050 11.400 ;
        RECT 583.950 12.600 586.050 13.050 ;
        RECT 613.950 12.600 616.050 13.050 ;
        RECT 583.950 11.400 616.050 12.600 ;
        RECT 583.950 10.950 586.050 11.400 ;
        RECT 613.950 10.950 616.050 11.400 ;
        RECT 358.950 8.400 414.600 9.600 ;
        RECT 490.950 9.600 493.050 10.050 ;
        RECT 547.950 9.600 550.050 10.050 ;
        RECT 490.950 8.400 550.050 9.600 ;
        RECT 358.950 7.950 361.050 8.400 ;
        RECT 490.950 7.950 493.050 8.400 ;
        RECT 547.950 7.950 550.050 8.400 ;
        RECT 760.950 9.600 763.050 10.050 ;
        RECT 784.950 9.600 787.050 10.050 ;
        RECT 805.950 9.600 808.050 10.050 ;
        RECT 760.950 8.400 808.050 9.600 ;
        RECT 760.950 7.950 763.050 8.400 ;
        RECT 784.950 7.950 787.050 8.400 ;
        RECT 805.950 7.950 808.050 8.400 ;
        RECT 430.950 6.600 433.050 7.050 ;
        RECT 457.950 6.600 460.050 7.050 ;
        RECT 430.950 5.400 460.050 6.600 ;
        RECT 430.950 4.950 433.050 5.400 ;
        RECT 457.950 4.950 460.050 5.400 ;
  END
END fir_pe
END LIBRARY

