magic
tech scmos
magscale 1 6
timestamp 1719894952
<< checkpaint >>
rect 684 5132 1062 5136
rect -121 5130 1062 5132
rect -121 4932 1134 5130
rect -121 4930 1171 4932
rect -260 -320 1171 4930
rect -260 -321 13 -320
<< nwell >>
rect 31 4220 841 4552
rect 31 2260 841 3820
<< psubstratepdiff >>
rect 31 4680 841 5012
rect 31 0 841 1560
<< nsubstratendiff >>
rect 31 4220 841 4552
rect 31 2260 841 3820
<< metal1 >>
rect 7 4680 865 5012
rect 7 4220 865 4552
rect 7 2260 865 3820
rect 7 0 865 1560
<< metal2 >>
rect 7 4680 865 5012
rect 7 4220 865 4552
rect 7 2260 865 3820
rect 7 0 865 1560
<< metal3 >>
rect 31 4680 841 5012
rect 31 4220 841 4552
rect 31 2260 841 3820
rect 31 0 841 1560
use IOFILLER10  IOFILLER10_0 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/chip_top/pads_ETRI050
timestamp 1537935238
transform 1 0 7 0 1 0
box -7 0 207 5012
use IOFILLER10  IOFILLER10_1
timestamp 1537935238
transform 1 0 665 0 1 0
box -7 0 207 5012
use IOFILLER10  IOFILLER10_2
timestamp 1537935238
transform 1 0 171 0 1 0
box -7 0 207 5012
use IOFILLER10  IOFILLER10_3
timestamp 1537935238
transform 1 0 335 0 1 0
box -7 0 207 5012
use IOFILLER10  IOFILLER10_4
timestamp 1537935238
transform 1 0 501 0 1 0
box -7 0 207 5012
<< end >>
