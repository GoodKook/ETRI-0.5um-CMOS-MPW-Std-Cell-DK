magic
tech scmos
magscale 1 2
timestamp 1702316108
<< nwell >>
rect -13 154 253 272
rect 11 152 74 154
<< ntransistor >>
rect 25 14 29 54
rect 45 14 49 34
rect 55 14 59 34
rect 77 14 81 34
rect 87 14 91 34
rect 109 14 113 34
rect 149 14 153 34
rect 159 14 163 34
rect 183 14 187 34
rect 193 14 197 34
rect 215 14 219 54
<< ptransistor >>
rect 25 166 29 246
rect 45 206 49 246
rect 61 206 65 246
rect 81 206 85 246
rect 93 206 97 246
rect 113 206 117 246
rect 153 206 157 246
rect 163 206 167 246
rect 183 226 187 246
rect 193 226 197 246
rect 215 166 219 246
<< ndiffusion >>
rect 23 14 25 54
rect 29 14 31 54
rect 43 14 45 34
rect 49 14 55 34
rect 59 14 63 34
rect 75 14 77 34
rect 81 14 87 34
rect 91 14 93 34
rect 105 14 109 34
rect 113 14 115 34
rect 147 14 149 34
rect 153 14 159 34
rect 163 14 165 34
rect 177 14 183 34
rect 187 14 193 34
rect 197 14 199 34
rect 211 14 215 54
rect 219 14 221 54
<< pdiffusion >>
rect 23 166 25 246
rect 29 166 31 246
rect 43 206 45 246
rect 49 206 61 246
rect 65 206 67 246
rect 79 206 81 246
rect 85 206 93 246
rect 97 206 99 246
rect 111 206 113 246
rect 117 206 119 246
rect 151 206 153 246
rect 157 206 163 246
rect 167 206 169 246
rect 181 226 183 246
rect 187 226 193 246
rect 197 226 201 246
rect 213 166 215 246
rect 219 166 221 246
<< ndcontact >>
rect 11 14 23 54
rect 31 14 43 54
rect 63 14 75 34
rect 93 14 105 34
rect 115 14 127 34
rect 135 14 147 34
rect 165 14 177 34
rect 199 14 211 54
rect 221 14 233 54
<< pdcontact >>
rect 11 166 23 246
rect 31 166 43 246
rect 67 206 79 246
rect 99 206 111 246
rect 119 206 131 246
rect 139 206 151 246
rect 169 206 181 246
rect 201 166 213 246
rect 221 166 233 246
<< psubstratepcontact >>
rect -6 -6 246 6
<< nsubstratencontact >>
rect -6 254 246 266
<< polysilicon >>
rect 25 246 29 250
rect 45 246 49 250
rect 61 246 65 250
rect 81 246 85 250
rect 93 246 97 250
rect 113 246 117 250
rect 153 246 157 250
rect 163 246 167 250
rect 183 246 187 250
rect 193 246 197 250
rect 215 246 219 250
rect 25 117 29 166
rect 25 54 29 105
rect 45 34 49 206
rect 61 142 65 206
rect 81 162 85 206
rect 93 200 97 206
rect 85 150 88 162
rect 61 138 76 142
rect 72 90 76 138
rect 84 70 88 150
rect 55 66 88 70
rect 55 34 59 66
rect 93 52 97 188
rect 113 180 117 206
rect 153 204 157 206
rect 127 200 157 204
rect 77 34 81 46
rect 87 36 101 40
rect 87 34 91 36
rect 109 34 113 168
rect 125 40 129 188
rect 163 186 167 206
rect 183 186 187 226
rect 193 200 197 226
rect 193 196 199 200
rect 161 174 167 186
rect 141 49 145 66
rect 163 57 167 174
rect 195 135 199 196
rect 163 53 187 57
rect 141 44 163 49
rect 125 36 153 40
rect 149 34 153 36
rect 159 34 163 44
rect 183 34 187 53
rect 193 34 197 65
rect 215 54 219 166
rect 25 10 29 14
rect 45 10 49 14
rect 55 10 59 14
rect 77 10 81 14
rect 87 10 91 14
rect 109 10 113 14
rect 149 10 153 14
rect 159 10 163 14
rect 183 10 187 14
rect 193 10 197 14
rect 215 10 219 14
<< polycontact >>
rect 23 105 35 117
rect 93 188 105 200
rect 73 150 85 162
rect 49 118 61 130
rect 64 78 76 90
rect 69 46 81 58
rect 105 168 117 180
rect 125 188 137 200
rect 89 40 101 52
rect 149 174 161 186
rect 175 174 187 186
rect 137 66 149 78
rect 188 123 200 135
rect 203 83 215 95
rect 185 65 197 77
<< metal1 >>
rect -6 266 246 268
rect -6 252 246 254
rect 31 246 43 252
rect 99 246 111 252
rect 139 246 151 252
rect 201 246 213 252
rect 7 166 11 178
rect 53 206 67 212
rect 119 200 125 206
rect 105 194 125 200
rect 67 172 105 180
rect 123 176 149 182
rect 7 160 13 166
rect 123 162 129 176
rect 167 168 175 186
rect 7 152 73 160
rect 7 54 13 152
rect 85 156 129 162
rect 143 162 175 168
rect 23 123 37 137
rect 103 130 117 137
rect 23 117 35 123
rect 61 123 117 130
rect 27 86 35 105
rect 27 78 64 86
rect 143 78 149 162
rect 221 137 233 166
rect 203 135 233 137
rect 200 123 233 135
rect 181 83 203 90
rect 69 70 137 78
rect 69 58 76 70
rect 221 74 233 123
rect 197 65 233 74
rect 7 42 11 54
rect 221 54 233 65
rect 101 40 121 46
rect 63 34 75 38
rect 115 34 121 40
rect 165 34 167 48
rect 51 28 63 34
rect 31 8 43 14
rect 93 8 105 14
rect 135 8 143 14
rect 199 8 211 14
rect -6 6 246 8
rect -6 -8 246 -6
<< m2contact >>
rect 53 192 67 206
rect 167 192 181 206
rect 53 172 67 186
rect 167 82 181 96
rect 49 34 63 48
rect 167 34 181 48
<< metal2 >>
rect 53 186 67 192
rect 55 153 63 172
rect 51 145 63 153
rect 51 48 59 145
rect 167 96 175 192
rect 167 48 175 82
<< m1p >>
rect -6 252 246 268
rect 23 123 37 137
rect 103 123 117 137
rect 203 123 217 137
rect -6 -8 246 8
<< labels >>
rlabel nsubstratencontact 120 260 120 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 120 0 120 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 30 131 30 131 0 CLK
port 2 nsew clock input
rlabel metal1 110 131 110 131 0 D
port 1 nsew signal input
rlabel metal1 210 131 210 131 0 Q
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 240 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
