magic
tech scmos
magscale 1 6
timestamp 1555589239
<< checkpaint >>
rect -110 -116 374 288
<< ntransistor >>
rect 49 14 59 114
rect 101 14 111 114
rect 153 14 163 114
rect 205 14 215 114
<< ndiffusion >>
rect 12 94 49 114
rect 12 82 22 94
rect 34 82 49 94
rect 12 70 49 82
rect 12 58 22 70
rect 34 58 49 70
rect 12 46 49 58
rect 12 34 22 46
rect 34 34 49 46
rect 12 14 49 34
rect 59 94 101 114
rect 59 82 74 94
rect 86 82 101 94
rect 59 70 101 82
rect 59 58 74 70
rect 86 58 101 70
rect 59 46 101 58
rect 59 34 74 46
rect 86 34 101 46
rect 59 14 101 34
rect 111 94 153 114
rect 111 82 126 94
rect 138 82 153 94
rect 111 70 153 82
rect 111 58 126 70
rect 138 58 153 70
rect 111 46 153 58
rect 111 34 126 46
rect 138 34 153 46
rect 111 14 153 34
rect 163 94 205 114
rect 163 82 178 94
rect 190 82 205 94
rect 163 70 205 82
rect 163 58 178 70
rect 190 58 205 70
rect 163 46 205 58
rect 163 34 178 46
rect 190 34 205 46
rect 163 14 205 34
rect 215 94 252 114
rect 215 82 230 94
rect 242 82 252 94
rect 215 70 252 82
rect 215 58 230 70
rect 242 58 252 70
rect 215 46 252 58
rect 215 34 230 46
rect 242 34 252 46
rect 215 14 252 34
<< ndcontact >>
rect 22 82 34 94
rect 22 58 34 70
rect 22 34 34 46
rect 74 82 86 94
rect 74 58 86 70
rect 74 34 86 46
rect 126 82 138 94
rect 126 58 138 70
rect 126 34 138 46
rect 178 82 190 94
rect 178 58 190 70
rect 178 34 190 46
rect 230 82 242 94
rect 230 58 242 70
rect 230 34 242 46
<< polysilicon >>
rect 49 114 59 134
rect 101 114 111 134
rect 153 114 163 134
rect 205 114 215 134
rect 49 4 59 14
rect 101 4 111 14
rect 153 4 163 14
rect 205 4 215 14
<< metal1 >>
rect 10 94 46 116
rect 10 82 22 94
rect 34 82 46 94
rect 10 70 46 82
rect 10 58 22 70
rect 34 58 46 70
rect 10 46 46 58
rect 10 34 22 46
rect 34 34 46 46
rect 10 12 46 34
rect 62 94 98 116
rect 62 82 74 94
rect 86 82 98 94
rect 62 70 98 82
rect 62 58 74 70
rect 86 58 98 70
rect 62 46 98 58
rect 62 34 74 46
rect 86 34 98 46
rect 62 12 98 34
rect 114 94 150 116
rect 114 82 126 94
rect 138 82 150 94
rect 114 70 150 82
rect 114 58 126 70
rect 138 58 150 70
rect 114 46 150 58
rect 114 34 126 46
rect 138 34 150 46
rect 114 12 150 34
rect 166 94 202 116
rect 166 82 178 94
rect 190 82 202 94
rect 166 70 202 82
rect 166 58 178 70
rect 190 58 202 70
rect 166 46 202 58
rect 166 34 178 46
rect 190 34 202 46
rect 166 12 202 34
rect 218 94 254 116
rect 218 82 230 94
rect 242 82 254 94
rect 218 70 254 82
rect 218 58 230 70
rect 242 58 254 70
rect 218 46 254 58
rect 218 34 230 46
rect 242 34 254 46
rect 218 12 254 34
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_0
timestamp 1555589239
transform 1 0 36 0 1 132
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_1
timestamp 1555589239
transform 1 0 88 0 1 132
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_2
timestamp 1555589239
transform 1 0 140 0 1 132
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_3
timestamp 1555589239
transform 1 0 192 0 1 132
box 0 0 36 36
<< end >>
