magic
tech scmos
magscale 1 60
timestamp 1709379016
<< checkpaint >>
rect -11389 22164 33724 75102
rect -1602 16129 29816 22164
rect -1200 15800 22105 16129
rect -1200 -1200 21900 15800
<< metal1 >>
rect 0 16500 17000 17000
rect 0 500 500 16500
rect 700 16180 1100 16300
rect 700 16020 820 16180
rect 980 16020 1100 16180
rect 700 15900 1100 16020
rect 1500 16180 1900 16300
rect 1500 16020 1620 16180
rect 1780 16020 1900 16180
rect 1500 15900 1900 16020
rect 2300 16180 2700 16300
rect 2300 16020 2420 16180
rect 2580 16020 2700 16180
rect 2300 15900 2700 16020
rect 3100 16180 3500 16300
rect 3100 16020 3220 16180
rect 3380 16020 3500 16180
rect 3100 15900 3500 16020
rect 3900 16180 4300 16300
rect 3900 16020 4020 16180
rect 4180 16020 4300 16180
rect 3900 15900 4300 16020
rect 4700 16180 5100 16300
rect 4700 16020 4820 16180
rect 4980 16020 5100 16180
rect 4700 15900 5100 16020
rect 5500 16180 5900 16300
rect 5500 16020 5620 16180
rect 5780 16020 5900 16180
rect 5500 15900 5900 16020
rect 6300 16180 6700 16300
rect 6300 16020 6420 16180
rect 6580 16020 6700 16180
rect 6300 15900 6700 16020
rect 7100 16180 7500 16300
rect 7100 16020 7220 16180
rect 7380 16020 7500 16180
rect 7100 15900 7500 16020
rect 7900 16180 8300 16300
rect 7900 16020 8020 16180
rect 8180 16020 8300 16180
rect 7900 15900 8300 16020
rect 8700 16180 9100 16300
rect 8700 16020 8820 16180
rect 8980 16020 9100 16180
rect 8700 15900 9100 16020
rect 9500 16180 9900 16300
rect 9500 16020 9620 16180
rect 9780 16020 9900 16180
rect 9500 15900 9900 16020
rect 10300 16180 10700 16300
rect 10300 16020 10420 16180
rect 10580 16020 10700 16180
rect 10300 15900 10700 16020
rect 11100 16180 11500 16300
rect 11100 16020 11220 16180
rect 11380 16020 11500 16180
rect 11100 15900 11500 16020
rect 11900 16180 12300 16300
rect 11900 16020 12020 16180
rect 12180 16020 12300 16180
rect 11900 15900 12300 16020
rect 12700 16180 13100 16300
rect 12700 16020 12820 16180
rect 12980 16020 13100 16180
rect 12700 15900 13100 16020
rect 13500 16180 13900 16300
rect 13500 16020 13620 16180
rect 13780 16020 13900 16180
rect 13500 15900 13900 16020
rect 14300 16180 14700 16300
rect 14300 16020 14420 16180
rect 14580 16020 14700 16180
rect 14300 15900 14700 16020
rect 15100 16180 15500 16300
rect 15100 16020 15220 16180
rect 15380 16020 15500 16180
rect 15100 15900 15500 16020
rect 15900 16180 16300 16300
rect 15900 16020 16020 16180
rect 16180 16020 16300 16180
rect 15900 15900 16300 16020
rect 700 15380 1100 15500
rect 700 15220 820 15380
rect 980 15220 1100 15380
rect 700 15100 1100 15220
rect 1500 15380 1900 15500
rect 1500 15220 1620 15380
rect 1780 15220 1900 15380
rect 1500 15100 1900 15220
rect 2300 15380 2700 15500
rect 2300 15220 2420 15380
rect 2580 15220 2700 15380
rect 2300 15100 2700 15220
rect 3100 15380 3500 15500
rect 3100 15220 3220 15380
rect 3380 15220 3500 15380
rect 3100 15100 3500 15220
rect 3900 15380 4300 15500
rect 3900 15220 4020 15380
rect 4180 15220 4300 15380
rect 3900 15100 4300 15220
rect 4700 15380 5100 15500
rect 4700 15220 4820 15380
rect 4980 15220 5100 15380
rect 4700 15100 5100 15220
rect 5500 15380 5900 15500
rect 5500 15220 5620 15380
rect 5780 15220 5900 15380
rect 5500 15100 5900 15220
rect 6300 15380 6700 15500
rect 6300 15220 6420 15380
rect 6580 15220 6700 15380
rect 6300 15100 6700 15220
rect 7100 15380 7500 15500
rect 7100 15220 7220 15380
rect 7380 15220 7500 15380
rect 7100 15100 7500 15220
rect 7900 15380 8300 15500
rect 7900 15220 8020 15380
rect 8180 15220 8300 15380
rect 7900 15100 8300 15220
rect 8700 15380 9100 15500
rect 8700 15220 8820 15380
rect 8980 15220 9100 15380
rect 8700 15100 9100 15220
rect 9500 15380 9900 15500
rect 9500 15220 9620 15380
rect 9780 15220 9900 15380
rect 9500 15100 9900 15220
rect 10300 15380 10700 15500
rect 10300 15220 10420 15380
rect 10580 15220 10700 15380
rect 10300 15100 10700 15220
rect 11100 15380 11500 15500
rect 11100 15220 11220 15380
rect 11380 15220 11500 15380
rect 11100 15100 11500 15220
rect 11900 15380 12300 15500
rect 11900 15220 12020 15380
rect 12180 15220 12300 15380
rect 11900 15100 12300 15220
rect 12700 15380 13100 15500
rect 12700 15220 12820 15380
rect 12980 15220 13100 15380
rect 12700 15100 13100 15220
rect 13500 15380 13900 15500
rect 13500 15220 13620 15380
rect 13780 15220 13900 15380
rect 13500 15100 13900 15220
rect 14300 15380 14700 15500
rect 14300 15220 14420 15380
rect 14580 15220 14700 15380
rect 14300 15100 14700 15220
rect 15100 15380 15500 15500
rect 15100 15220 15220 15380
rect 15380 15220 15500 15380
rect 15100 15100 15500 15220
rect 15900 15380 16300 15500
rect 15900 15220 16020 15380
rect 16180 15220 16300 15380
rect 15900 15100 16300 15220
rect 700 14580 1100 14700
rect 700 14420 820 14580
rect 980 14420 1100 14580
rect 700 14300 1100 14420
rect 1500 14580 1900 14700
rect 1500 14420 1620 14580
rect 1780 14420 1900 14580
rect 1500 14300 1900 14420
rect 2300 14580 2700 14700
rect 2300 14420 2420 14580
rect 2580 14420 2700 14580
rect 2300 14300 2700 14420
rect 3100 14580 3500 14700
rect 3100 14420 3220 14580
rect 3380 14420 3500 14580
rect 3100 14300 3500 14420
rect 3900 14580 4300 14700
rect 3900 14420 4020 14580
rect 4180 14420 4300 14580
rect 3900 14300 4300 14420
rect 4700 14580 5100 14700
rect 4700 14420 4820 14580
rect 4980 14420 5100 14580
rect 4700 14300 5100 14420
rect 5500 14580 5900 14700
rect 5500 14420 5620 14580
rect 5780 14420 5900 14580
rect 5500 14300 5900 14420
rect 6300 14580 6700 14700
rect 6300 14420 6420 14580
rect 6580 14420 6700 14580
rect 6300 14300 6700 14420
rect 7100 14580 7500 14700
rect 7100 14420 7220 14580
rect 7380 14420 7500 14580
rect 7100 14300 7500 14420
rect 7900 14580 8300 14700
rect 7900 14420 8020 14580
rect 8180 14420 8300 14580
rect 7900 14300 8300 14420
rect 8700 14580 9100 14700
rect 8700 14420 8820 14580
rect 8980 14420 9100 14580
rect 8700 14300 9100 14420
rect 9500 14580 9900 14700
rect 9500 14420 9620 14580
rect 9780 14420 9900 14580
rect 9500 14300 9900 14420
rect 10300 14580 10700 14700
rect 10300 14420 10420 14580
rect 10580 14420 10700 14580
rect 10300 14300 10700 14420
rect 11100 14580 11500 14700
rect 11100 14420 11220 14580
rect 11380 14420 11500 14580
rect 11100 14300 11500 14420
rect 11900 14580 12300 14700
rect 11900 14420 12020 14580
rect 12180 14420 12300 14580
rect 11900 14300 12300 14420
rect 12700 14580 13100 14700
rect 12700 14420 12820 14580
rect 12980 14420 13100 14580
rect 12700 14300 13100 14420
rect 13500 14580 13900 14700
rect 13500 14420 13620 14580
rect 13780 14420 13900 14580
rect 13500 14300 13900 14420
rect 14300 14580 14700 14700
rect 14300 14420 14420 14580
rect 14580 14420 14700 14580
rect 14300 14300 14700 14420
rect 15100 14580 15500 14700
rect 15100 14420 15220 14580
rect 15380 14420 15500 14580
rect 15100 14300 15500 14420
rect 15900 14580 16300 14700
rect 15900 14420 16020 14580
rect 16180 14420 16300 14580
rect 15900 14300 16300 14420
rect 700 13780 1100 13900
rect 700 13620 820 13780
rect 980 13620 1100 13780
rect 700 13500 1100 13620
rect 1500 13780 1900 13900
rect 1500 13620 1620 13780
rect 1780 13620 1900 13780
rect 1500 13500 1900 13620
rect 2300 13780 2700 13900
rect 2300 13620 2420 13780
rect 2580 13620 2700 13780
rect 2300 13500 2700 13620
rect 3100 13780 3500 13900
rect 3100 13620 3220 13780
rect 3380 13620 3500 13780
rect 3100 13500 3500 13620
rect 3900 13780 4300 13900
rect 3900 13620 4020 13780
rect 4180 13620 4300 13780
rect 3900 13500 4300 13620
rect 4700 13780 5100 13900
rect 4700 13620 4820 13780
rect 4980 13620 5100 13780
rect 4700 13500 5100 13620
rect 5500 13780 5900 13900
rect 5500 13620 5620 13780
rect 5780 13620 5900 13780
rect 5500 13500 5900 13620
rect 6300 13780 6700 13900
rect 6300 13620 6420 13780
rect 6580 13620 6700 13780
rect 6300 13500 6700 13620
rect 7100 13780 7500 13900
rect 7100 13620 7220 13780
rect 7380 13620 7500 13780
rect 7100 13500 7500 13620
rect 7900 13780 8300 13900
rect 7900 13620 8020 13780
rect 8180 13620 8300 13780
rect 7900 13500 8300 13620
rect 8700 13780 9100 13900
rect 8700 13620 8820 13780
rect 8980 13620 9100 13780
rect 8700 13500 9100 13620
rect 9500 13780 9900 13900
rect 9500 13620 9620 13780
rect 9780 13620 9900 13780
rect 9500 13500 9900 13620
rect 10300 13780 10700 13900
rect 10300 13620 10420 13780
rect 10580 13620 10700 13780
rect 10300 13500 10700 13620
rect 11100 13780 11500 13900
rect 11100 13620 11220 13780
rect 11380 13620 11500 13780
rect 11100 13500 11500 13620
rect 11900 13780 12300 13900
rect 11900 13620 12020 13780
rect 12180 13620 12300 13780
rect 11900 13500 12300 13620
rect 12700 13780 13100 13900
rect 12700 13620 12820 13780
rect 12980 13620 13100 13780
rect 12700 13500 13100 13620
rect 13500 13780 13900 13900
rect 13500 13620 13620 13780
rect 13780 13620 13900 13780
rect 13500 13500 13900 13620
rect 14300 13780 14700 13900
rect 14300 13620 14420 13780
rect 14580 13620 14700 13780
rect 14300 13500 14700 13620
rect 15100 13780 15500 13900
rect 15100 13620 15220 13780
rect 15380 13620 15500 13780
rect 15100 13500 15500 13620
rect 15900 13780 16300 13900
rect 15900 13620 16020 13780
rect 16180 13620 16300 13780
rect 15900 13500 16300 13620
rect 700 12980 1100 13100
rect 700 12820 820 12980
rect 980 12820 1100 12980
rect 700 12700 1100 12820
rect 1500 12980 1900 13100
rect 1500 12820 1620 12980
rect 1780 12820 1900 12980
rect 1500 12700 1900 12820
rect 2300 12980 2700 13100
rect 2300 12820 2420 12980
rect 2580 12820 2700 12980
rect 2300 12700 2700 12820
rect 3100 12980 3500 13100
rect 3100 12820 3220 12980
rect 3380 12820 3500 12980
rect 3100 12700 3500 12820
rect 3900 12980 4300 13100
rect 3900 12820 4020 12980
rect 4180 12820 4300 12980
rect 3900 12700 4300 12820
rect 4700 12980 5100 13100
rect 4700 12820 4820 12980
rect 4980 12820 5100 12980
rect 4700 12700 5100 12820
rect 5500 12980 5900 13100
rect 5500 12820 5620 12980
rect 5780 12820 5900 12980
rect 5500 12700 5900 12820
rect 6300 12980 6700 13100
rect 6300 12820 6420 12980
rect 6580 12820 6700 12980
rect 6300 12700 6700 12820
rect 7100 12980 7500 13100
rect 7100 12820 7220 12980
rect 7380 12820 7500 12980
rect 7100 12700 7500 12820
rect 7900 12980 8300 13100
rect 7900 12820 8020 12980
rect 8180 12820 8300 12980
rect 7900 12700 8300 12820
rect 8700 12980 9100 13100
rect 8700 12820 8820 12980
rect 8980 12820 9100 12980
rect 8700 12700 9100 12820
rect 9500 12980 9900 13100
rect 9500 12820 9620 12980
rect 9780 12820 9900 12980
rect 9500 12700 9900 12820
rect 10300 12980 10700 13100
rect 10300 12820 10420 12980
rect 10580 12820 10700 12980
rect 10300 12700 10700 12820
rect 11100 12980 11500 13100
rect 11100 12820 11220 12980
rect 11380 12820 11500 12980
rect 11100 12700 11500 12820
rect 11900 12980 12300 13100
rect 11900 12820 12020 12980
rect 12180 12820 12300 12980
rect 11900 12700 12300 12820
rect 12700 12980 13100 13100
rect 12700 12820 12820 12980
rect 12980 12820 13100 12980
rect 12700 12700 13100 12820
rect 13500 12980 13900 13100
rect 13500 12820 13620 12980
rect 13780 12820 13900 12980
rect 13500 12700 13900 12820
rect 14300 12980 14700 13100
rect 14300 12820 14420 12980
rect 14580 12820 14700 12980
rect 14300 12700 14700 12820
rect 15100 12980 15500 13100
rect 15100 12820 15220 12980
rect 15380 12820 15500 12980
rect 15100 12700 15500 12820
rect 15900 12980 16300 13100
rect 15900 12820 16020 12980
rect 16180 12820 16300 12980
rect 15900 12700 16300 12820
rect 700 12180 1100 12300
rect 700 12020 820 12180
rect 980 12020 1100 12180
rect 700 11900 1100 12020
rect 1500 12180 1900 12300
rect 1500 12020 1620 12180
rect 1780 12020 1900 12180
rect 1500 11900 1900 12020
rect 2300 12180 2700 12300
rect 2300 12020 2420 12180
rect 2580 12020 2700 12180
rect 2300 11900 2700 12020
rect 3100 12180 3500 12300
rect 3100 12020 3220 12180
rect 3380 12020 3500 12180
rect 3100 11900 3500 12020
rect 3900 12180 4300 12300
rect 3900 12020 4020 12180
rect 4180 12020 4300 12180
rect 3900 11900 4300 12020
rect 4700 12180 5100 12300
rect 4700 12020 4820 12180
rect 4980 12020 5100 12180
rect 4700 11900 5100 12020
rect 5500 12180 5900 12300
rect 5500 12020 5620 12180
rect 5780 12020 5900 12180
rect 5500 11900 5900 12020
rect 6300 12180 6700 12300
rect 6300 12020 6420 12180
rect 6580 12020 6700 12180
rect 6300 11900 6700 12020
rect 7100 12180 7500 12300
rect 7100 12020 7220 12180
rect 7380 12020 7500 12180
rect 7100 11900 7500 12020
rect 7900 12180 8300 12300
rect 7900 12020 8020 12180
rect 8180 12020 8300 12180
rect 7900 11900 8300 12020
rect 8700 12180 9100 12300
rect 8700 12020 8820 12180
rect 8980 12020 9100 12180
rect 8700 11900 9100 12020
rect 9500 12180 9900 12300
rect 9500 12020 9620 12180
rect 9780 12020 9900 12180
rect 9500 11900 9900 12020
rect 10300 12180 10700 12300
rect 10300 12020 10420 12180
rect 10580 12020 10700 12180
rect 10300 11900 10700 12020
rect 11100 12180 11500 12300
rect 11100 12020 11220 12180
rect 11380 12020 11500 12180
rect 11100 11900 11500 12020
rect 11900 12180 12300 12300
rect 11900 12020 12020 12180
rect 12180 12020 12300 12180
rect 11900 11900 12300 12020
rect 12700 12180 13100 12300
rect 12700 12020 12820 12180
rect 12980 12020 13100 12180
rect 12700 11900 13100 12020
rect 13500 12180 13900 12300
rect 13500 12020 13620 12180
rect 13780 12020 13900 12180
rect 13500 11900 13900 12020
rect 14300 12180 14700 12300
rect 14300 12020 14420 12180
rect 14580 12020 14700 12180
rect 14300 11900 14700 12020
rect 15100 12180 15500 12300
rect 15100 12020 15220 12180
rect 15380 12020 15500 12180
rect 15100 11900 15500 12020
rect 15900 12180 16300 12300
rect 15900 12020 16020 12180
rect 16180 12020 16300 12180
rect 15900 11900 16300 12020
rect 700 11380 1100 11500
rect 700 11220 820 11380
rect 980 11220 1100 11380
rect 700 11100 1100 11220
rect 1500 11380 1900 11500
rect 1500 11220 1620 11380
rect 1780 11220 1900 11380
rect 1500 11100 1900 11220
rect 2300 11380 2700 11500
rect 2300 11220 2420 11380
rect 2580 11220 2700 11380
rect 2300 11100 2700 11220
rect 3100 11380 3500 11500
rect 3100 11220 3220 11380
rect 3380 11220 3500 11380
rect 3100 11100 3500 11220
rect 3900 11380 4300 11500
rect 3900 11220 4020 11380
rect 4180 11220 4300 11380
rect 3900 11100 4300 11220
rect 4700 11380 5100 11500
rect 4700 11220 4820 11380
rect 4980 11220 5100 11380
rect 4700 11100 5100 11220
rect 5500 11380 5900 11500
rect 5500 11220 5620 11380
rect 5780 11220 5900 11380
rect 5500 11100 5900 11220
rect 6300 11380 6700 11500
rect 6300 11220 6420 11380
rect 6580 11220 6700 11380
rect 6300 11100 6700 11220
rect 7100 11380 7500 11500
rect 7100 11220 7220 11380
rect 7380 11220 7500 11380
rect 7100 11100 7500 11220
rect 7900 11380 8300 11500
rect 7900 11220 8020 11380
rect 8180 11220 8300 11380
rect 7900 11100 8300 11220
rect 8700 11380 9100 11500
rect 8700 11220 8820 11380
rect 8980 11220 9100 11380
rect 8700 11100 9100 11220
rect 9500 11380 9900 11500
rect 9500 11220 9620 11380
rect 9780 11220 9900 11380
rect 9500 11100 9900 11220
rect 10300 11380 10700 11500
rect 10300 11220 10420 11380
rect 10580 11220 10700 11380
rect 10300 11100 10700 11220
rect 11100 11380 11500 11500
rect 11100 11220 11220 11380
rect 11380 11220 11500 11380
rect 11100 11100 11500 11220
rect 11900 11380 12300 11500
rect 11900 11220 12020 11380
rect 12180 11220 12300 11380
rect 11900 11100 12300 11220
rect 12700 11380 13100 11500
rect 12700 11220 12820 11380
rect 12980 11220 13100 11380
rect 12700 11100 13100 11220
rect 13500 11380 13900 11500
rect 13500 11220 13620 11380
rect 13780 11220 13900 11380
rect 13500 11100 13900 11220
rect 14300 11380 14700 11500
rect 14300 11220 14420 11380
rect 14580 11220 14700 11380
rect 14300 11100 14700 11220
rect 15100 11380 15500 11500
rect 15100 11220 15220 11380
rect 15380 11220 15500 11380
rect 15100 11100 15500 11220
rect 15900 11380 16300 11500
rect 15900 11220 16020 11380
rect 16180 11220 16300 11380
rect 15900 11100 16300 11220
rect 700 10580 1100 10700
rect 700 10420 820 10580
rect 980 10420 1100 10580
rect 700 10300 1100 10420
rect 1500 10580 1900 10700
rect 1500 10420 1620 10580
rect 1780 10420 1900 10580
rect 1500 10300 1900 10420
rect 2300 10580 2700 10700
rect 2300 10420 2420 10580
rect 2580 10420 2700 10580
rect 2300 10300 2700 10420
rect 3100 10580 3500 10700
rect 3100 10420 3220 10580
rect 3380 10420 3500 10580
rect 3100 10300 3500 10420
rect 3900 10580 4300 10700
rect 3900 10420 4020 10580
rect 4180 10420 4300 10580
rect 3900 10300 4300 10420
rect 4700 10580 5100 10700
rect 4700 10420 4820 10580
rect 4980 10420 5100 10580
rect 4700 10300 5100 10420
rect 5500 10580 5900 10700
rect 5500 10420 5620 10580
rect 5780 10420 5900 10580
rect 5500 10300 5900 10420
rect 6300 10580 6700 10700
rect 6300 10420 6420 10580
rect 6580 10420 6700 10580
rect 6300 10300 6700 10420
rect 7100 10580 7500 10700
rect 7100 10420 7220 10580
rect 7380 10420 7500 10580
rect 7100 10300 7500 10420
rect 7900 10580 8300 10700
rect 7900 10420 8020 10580
rect 8180 10420 8300 10580
rect 7900 10300 8300 10420
rect 8700 10580 9100 10700
rect 8700 10420 8820 10580
rect 8980 10420 9100 10580
rect 8700 10300 9100 10420
rect 9500 10580 9900 10700
rect 9500 10420 9620 10580
rect 9780 10420 9900 10580
rect 9500 10300 9900 10420
rect 10300 10580 10700 10700
rect 10300 10420 10420 10580
rect 10580 10420 10700 10580
rect 10300 10300 10700 10420
rect 11100 10580 11500 10700
rect 11100 10420 11220 10580
rect 11380 10420 11500 10580
rect 11100 10300 11500 10420
rect 11900 10580 12300 10700
rect 11900 10420 12020 10580
rect 12180 10420 12300 10580
rect 11900 10300 12300 10420
rect 12700 10580 13100 10700
rect 12700 10420 12820 10580
rect 12980 10420 13100 10580
rect 12700 10300 13100 10420
rect 13500 10580 13900 10700
rect 13500 10420 13620 10580
rect 13780 10420 13900 10580
rect 13500 10300 13900 10420
rect 14300 10580 14700 10700
rect 14300 10420 14420 10580
rect 14580 10420 14700 10580
rect 14300 10300 14700 10420
rect 15100 10580 15500 10700
rect 15100 10420 15220 10580
rect 15380 10420 15500 10580
rect 15100 10300 15500 10420
rect 15900 10580 16300 10700
rect 15900 10420 16020 10580
rect 16180 10420 16300 10580
rect 15900 10300 16300 10420
rect 700 9780 1100 9900
rect 700 9620 820 9780
rect 980 9620 1100 9780
rect 700 9500 1100 9620
rect 1500 9780 1900 9900
rect 1500 9620 1620 9780
rect 1780 9620 1900 9780
rect 1500 9500 1900 9620
rect 2300 9780 2700 9900
rect 2300 9620 2420 9780
rect 2580 9620 2700 9780
rect 2300 9500 2700 9620
rect 3100 9780 3500 9900
rect 3100 9620 3220 9780
rect 3380 9620 3500 9780
rect 3100 9500 3500 9620
rect 3900 9780 4300 9900
rect 3900 9620 4020 9780
rect 4180 9620 4300 9780
rect 3900 9500 4300 9620
rect 4700 9780 5100 9900
rect 4700 9620 4820 9780
rect 4980 9620 5100 9780
rect 4700 9500 5100 9620
rect 5500 9780 5900 9900
rect 5500 9620 5620 9780
rect 5780 9620 5900 9780
rect 5500 9500 5900 9620
rect 6300 9780 6700 9900
rect 6300 9620 6420 9780
rect 6580 9620 6700 9780
rect 6300 9500 6700 9620
rect 7100 9780 7500 9900
rect 7100 9620 7220 9780
rect 7380 9620 7500 9780
rect 7100 9500 7500 9620
rect 7900 9780 8300 9900
rect 7900 9620 8020 9780
rect 8180 9620 8300 9780
rect 7900 9500 8300 9620
rect 8700 9780 9100 9900
rect 8700 9620 8820 9780
rect 8980 9620 9100 9780
rect 8700 9500 9100 9620
rect 9500 9780 9900 9900
rect 9500 9620 9620 9780
rect 9780 9620 9900 9780
rect 9500 9500 9900 9620
rect 10300 9780 10700 9900
rect 10300 9620 10420 9780
rect 10580 9620 10700 9780
rect 10300 9500 10700 9620
rect 11100 9780 11500 9900
rect 11100 9620 11220 9780
rect 11380 9620 11500 9780
rect 11100 9500 11500 9620
rect 11900 9780 12300 9900
rect 11900 9620 12020 9780
rect 12180 9620 12300 9780
rect 11900 9500 12300 9620
rect 12700 9780 13100 9900
rect 12700 9620 12820 9780
rect 12980 9620 13100 9780
rect 12700 9500 13100 9620
rect 13500 9780 13900 9900
rect 13500 9620 13620 9780
rect 13780 9620 13900 9780
rect 13500 9500 13900 9620
rect 14300 9780 14700 9900
rect 14300 9620 14420 9780
rect 14580 9620 14700 9780
rect 14300 9500 14700 9620
rect 15100 9780 15500 9900
rect 15100 9620 15220 9780
rect 15380 9620 15500 9780
rect 15100 9500 15500 9620
rect 15900 9780 16300 9900
rect 15900 9620 16020 9780
rect 16180 9620 16300 9780
rect 15900 9500 16300 9620
rect 700 8980 1100 9100
rect 700 8820 820 8980
rect 980 8820 1100 8980
rect 700 8700 1100 8820
rect 1500 8980 1900 9100
rect 1500 8820 1620 8980
rect 1780 8820 1900 8980
rect 1500 8700 1900 8820
rect 2300 8980 2700 9100
rect 2300 8820 2420 8980
rect 2580 8820 2700 8980
rect 2300 8700 2700 8820
rect 3100 8980 3500 9100
rect 3100 8820 3220 8980
rect 3380 8820 3500 8980
rect 3100 8700 3500 8820
rect 3900 8980 4300 9100
rect 3900 8820 4020 8980
rect 4180 8820 4300 8980
rect 3900 8700 4300 8820
rect 4700 8980 5100 9100
rect 4700 8820 4820 8980
rect 4980 8820 5100 8980
rect 4700 8700 5100 8820
rect 5500 8980 5900 9100
rect 5500 8820 5620 8980
rect 5780 8820 5900 8980
rect 5500 8700 5900 8820
rect 6300 8980 6700 9100
rect 6300 8820 6420 8980
rect 6580 8820 6700 8980
rect 6300 8700 6700 8820
rect 7100 8980 7500 9100
rect 7100 8820 7220 8980
rect 7380 8820 7500 8980
rect 7100 8700 7500 8820
rect 7900 8980 8300 9100
rect 7900 8820 8020 8980
rect 8180 8820 8300 8980
rect 7900 8700 8300 8820
rect 8700 8980 9100 9100
rect 8700 8820 8820 8980
rect 8980 8820 9100 8980
rect 8700 8700 9100 8820
rect 9500 8980 9900 9100
rect 9500 8820 9620 8980
rect 9780 8820 9900 8980
rect 9500 8700 9900 8820
rect 10300 8980 10700 9100
rect 10300 8820 10420 8980
rect 10580 8820 10700 8980
rect 10300 8700 10700 8820
rect 11100 8980 11500 9100
rect 11100 8820 11220 8980
rect 11380 8820 11500 8980
rect 11100 8700 11500 8820
rect 11900 8980 12300 9100
rect 11900 8820 12020 8980
rect 12180 8820 12300 8980
rect 11900 8700 12300 8820
rect 12700 8980 13100 9100
rect 12700 8820 12820 8980
rect 12980 8820 13100 8980
rect 12700 8700 13100 8820
rect 13500 8980 13900 9100
rect 13500 8820 13620 8980
rect 13780 8820 13900 8980
rect 13500 8700 13900 8820
rect 14300 8980 14700 9100
rect 14300 8820 14420 8980
rect 14580 8820 14700 8980
rect 14300 8700 14700 8820
rect 15100 8980 15500 9100
rect 15100 8820 15220 8980
rect 15380 8820 15500 8980
rect 15100 8700 15500 8820
rect 15900 8980 16300 9100
rect 15900 8820 16020 8980
rect 16180 8820 16300 8980
rect 15900 8700 16300 8820
rect 700 8180 1100 8300
rect 700 8020 820 8180
rect 980 8020 1100 8180
rect 700 7900 1100 8020
rect 1500 8180 1900 8300
rect 1500 8020 1620 8180
rect 1780 8020 1900 8180
rect 1500 7900 1900 8020
rect 2300 8180 2700 8300
rect 2300 8020 2420 8180
rect 2580 8020 2700 8180
rect 2300 7900 2700 8020
rect 3100 8180 3500 8300
rect 3100 8020 3220 8180
rect 3380 8020 3500 8180
rect 3100 7900 3500 8020
rect 3900 8180 4300 8300
rect 3900 8020 4020 8180
rect 4180 8020 4300 8180
rect 3900 7900 4300 8020
rect 4700 8180 5100 8300
rect 4700 8020 4820 8180
rect 4980 8020 5100 8180
rect 4700 7900 5100 8020
rect 5500 8180 5900 8300
rect 5500 8020 5620 8180
rect 5780 8020 5900 8180
rect 5500 7900 5900 8020
rect 6300 8180 6700 8300
rect 6300 8020 6420 8180
rect 6580 8020 6700 8180
rect 6300 7900 6700 8020
rect 7100 8180 7500 8300
rect 7100 8020 7220 8180
rect 7380 8020 7500 8180
rect 7100 7900 7500 8020
rect 7900 8180 8300 8300
rect 7900 8020 8020 8180
rect 8180 8020 8300 8180
rect 7900 7900 8300 8020
rect 8700 8180 9100 8300
rect 8700 8020 8820 8180
rect 8980 8020 9100 8180
rect 8700 7900 9100 8020
rect 9500 8180 9900 8300
rect 9500 8020 9620 8180
rect 9780 8020 9900 8180
rect 9500 7900 9900 8020
rect 10300 8180 10700 8300
rect 10300 8020 10420 8180
rect 10580 8020 10700 8180
rect 10300 7900 10700 8020
rect 11100 8180 11500 8300
rect 11100 8020 11220 8180
rect 11380 8020 11500 8180
rect 11100 7900 11500 8020
rect 11900 8180 12300 8300
rect 11900 8020 12020 8180
rect 12180 8020 12300 8180
rect 11900 7900 12300 8020
rect 12700 8180 13100 8300
rect 12700 8020 12820 8180
rect 12980 8020 13100 8180
rect 12700 7900 13100 8020
rect 13500 8180 13900 8300
rect 13500 8020 13620 8180
rect 13780 8020 13900 8180
rect 13500 7900 13900 8020
rect 14300 8180 14700 8300
rect 14300 8020 14420 8180
rect 14580 8020 14700 8180
rect 14300 7900 14700 8020
rect 15100 8180 15500 8300
rect 15100 8020 15220 8180
rect 15380 8020 15500 8180
rect 15100 7900 15500 8020
rect 15900 8180 16300 8300
rect 15900 8020 16020 8180
rect 16180 8020 16300 8180
rect 15900 7900 16300 8020
rect 700 7380 1100 7500
rect 700 7220 820 7380
rect 980 7220 1100 7380
rect 700 7100 1100 7220
rect 1500 7380 1900 7500
rect 1500 7220 1620 7380
rect 1780 7220 1900 7380
rect 1500 7100 1900 7220
rect 2300 7380 2700 7500
rect 2300 7220 2420 7380
rect 2580 7220 2700 7380
rect 2300 7100 2700 7220
rect 3100 7380 3500 7500
rect 3100 7220 3220 7380
rect 3380 7220 3500 7380
rect 3100 7100 3500 7220
rect 3900 7380 4300 7500
rect 3900 7220 4020 7380
rect 4180 7220 4300 7380
rect 3900 7100 4300 7220
rect 4700 7380 5100 7500
rect 4700 7220 4820 7380
rect 4980 7220 5100 7380
rect 4700 7100 5100 7220
rect 5500 7380 5900 7500
rect 5500 7220 5620 7380
rect 5780 7220 5900 7380
rect 5500 7100 5900 7220
rect 6300 7380 6700 7500
rect 6300 7220 6420 7380
rect 6580 7220 6700 7380
rect 6300 7100 6700 7220
rect 7100 7380 7500 7500
rect 7100 7220 7220 7380
rect 7380 7220 7500 7380
rect 7100 7100 7500 7220
rect 7900 7380 8300 7500
rect 7900 7220 8020 7380
rect 8180 7220 8300 7380
rect 7900 7100 8300 7220
rect 8700 7380 9100 7500
rect 8700 7220 8820 7380
rect 8980 7220 9100 7380
rect 8700 7100 9100 7220
rect 9500 7380 9900 7500
rect 9500 7220 9620 7380
rect 9780 7220 9900 7380
rect 9500 7100 9900 7220
rect 10300 7380 10700 7500
rect 10300 7220 10420 7380
rect 10580 7220 10700 7380
rect 10300 7100 10700 7220
rect 11100 7380 11500 7500
rect 11100 7220 11220 7380
rect 11380 7220 11500 7380
rect 11100 7100 11500 7220
rect 11900 7380 12300 7500
rect 11900 7220 12020 7380
rect 12180 7220 12300 7380
rect 11900 7100 12300 7220
rect 12700 7380 13100 7500
rect 12700 7220 12820 7380
rect 12980 7220 13100 7380
rect 12700 7100 13100 7220
rect 13500 7380 13900 7500
rect 13500 7220 13620 7380
rect 13780 7220 13900 7380
rect 13500 7100 13900 7220
rect 14300 7380 14700 7500
rect 14300 7220 14420 7380
rect 14580 7220 14700 7380
rect 14300 7100 14700 7220
rect 15100 7380 15500 7500
rect 15100 7220 15220 7380
rect 15380 7220 15500 7380
rect 15100 7100 15500 7220
rect 15900 7380 16300 7500
rect 15900 7220 16020 7380
rect 16180 7220 16300 7380
rect 15900 7100 16300 7220
rect 700 6580 1100 6700
rect 700 6420 820 6580
rect 980 6420 1100 6580
rect 700 6300 1100 6420
rect 1500 6580 1900 6700
rect 1500 6420 1620 6580
rect 1780 6420 1900 6580
rect 1500 6300 1900 6420
rect 2300 6580 2700 6700
rect 2300 6420 2420 6580
rect 2580 6420 2700 6580
rect 2300 6300 2700 6420
rect 3100 6580 3500 6700
rect 3100 6420 3220 6580
rect 3380 6420 3500 6580
rect 3100 6300 3500 6420
rect 3900 6580 4300 6700
rect 3900 6420 4020 6580
rect 4180 6420 4300 6580
rect 3900 6300 4300 6420
rect 4700 6580 5100 6700
rect 4700 6420 4820 6580
rect 4980 6420 5100 6580
rect 4700 6300 5100 6420
rect 5500 6580 5900 6700
rect 5500 6420 5620 6580
rect 5780 6420 5900 6580
rect 5500 6300 5900 6420
rect 6300 6580 6700 6700
rect 6300 6420 6420 6580
rect 6580 6420 6700 6580
rect 6300 6300 6700 6420
rect 7100 6580 7500 6700
rect 7100 6420 7220 6580
rect 7380 6420 7500 6580
rect 7100 6300 7500 6420
rect 7900 6580 8300 6700
rect 7900 6420 8020 6580
rect 8180 6420 8300 6580
rect 7900 6300 8300 6420
rect 8700 6580 9100 6700
rect 8700 6420 8820 6580
rect 8980 6420 9100 6580
rect 8700 6300 9100 6420
rect 9500 6580 9900 6700
rect 9500 6420 9620 6580
rect 9780 6420 9900 6580
rect 9500 6300 9900 6420
rect 10300 6580 10700 6700
rect 10300 6420 10420 6580
rect 10580 6420 10700 6580
rect 10300 6300 10700 6420
rect 11100 6580 11500 6700
rect 11100 6420 11220 6580
rect 11380 6420 11500 6580
rect 11100 6300 11500 6420
rect 11900 6580 12300 6700
rect 11900 6420 12020 6580
rect 12180 6420 12300 6580
rect 11900 6300 12300 6420
rect 12700 6580 13100 6700
rect 12700 6420 12820 6580
rect 12980 6420 13100 6580
rect 12700 6300 13100 6420
rect 13500 6580 13900 6700
rect 13500 6420 13620 6580
rect 13780 6420 13900 6580
rect 13500 6300 13900 6420
rect 14300 6580 14700 6700
rect 14300 6420 14420 6580
rect 14580 6420 14700 6580
rect 14300 6300 14700 6420
rect 15100 6580 15500 6700
rect 15100 6420 15220 6580
rect 15380 6420 15500 6580
rect 15100 6300 15500 6420
rect 15900 6580 16300 6700
rect 15900 6420 16020 6580
rect 16180 6420 16300 6580
rect 15900 6300 16300 6420
rect 700 5780 1100 5900
rect 700 5620 820 5780
rect 980 5620 1100 5780
rect 700 5500 1100 5620
rect 1500 5780 1900 5900
rect 1500 5620 1620 5780
rect 1780 5620 1900 5780
rect 1500 5500 1900 5620
rect 2300 5780 2700 5900
rect 2300 5620 2420 5780
rect 2580 5620 2700 5780
rect 2300 5500 2700 5620
rect 3100 5780 3500 5900
rect 3100 5620 3220 5780
rect 3380 5620 3500 5780
rect 3100 5500 3500 5620
rect 3900 5780 4300 5900
rect 3900 5620 4020 5780
rect 4180 5620 4300 5780
rect 3900 5500 4300 5620
rect 4700 5780 5100 5900
rect 4700 5620 4820 5780
rect 4980 5620 5100 5780
rect 4700 5500 5100 5620
rect 5500 5780 5900 5900
rect 5500 5620 5620 5780
rect 5780 5620 5900 5780
rect 5500 5500 5900 5620
rect 6300 5780 6700 5900
rect 6300 5620 6420 5780
rect 6580 5620 6700 5780
rect 6300 5500 6700 5620
rect 7100 5780 7500 5900
rect 7100 5620 7220 5780
rect 7380 5620 7500 5780
rect 7100 5500 7500 5620
rect 7900 5780 8300 5900
rect 7900 5620 8020 5780
rect 8180 5620 8300 5780
rect 7900 5500 8300 5620
rect 8700 5780 9100 5900
rect 8700 5620 8820 5780
rect 8980 5620 9100 5780
rect 8700 5500 9100 5620
rect 9500 5780 9900 5900
rect 9500 5620 9620 5780
rect 9780 5620 9900 5780
rect 9500 5500 9900 5620
rect 10300 5780 10700 5900
rect 10300 5620 10420 5780
rect 10580 5620 10700 5780
rect 10300 5500 10700 5620
rect 11100 5780 11500 5900
rect 11100 5620 11220 5780
rect 11380 5620 11500 5780
rect 11100 5500 11500 5620
rect 11900 5780 12300 5900
rect 11900 5620 12020 5780
rect 12180 5620 12300 5780
rect 11900 5500 12300 5620
rect 12700 5780 13100 5900
rect 12700 5620 12820 5780
rect 12980 5620 13100 5780
rect 12700 5500 13100 5620
rect 13500 5780 13900 5900
rect 13500 5620 13620 5780
rect 13780 5620 13900 5780
rect 13500 5500 13900 5620
rect 14300 5780 14700 5900
rect 14300 5620 14420 5780
rect 14580 5620 14700 5780
rect 14300 5500 14700 5620
rect 15100 5780 15500 5900
rect 15100 5620 15220 5780
rect 15380 5620 15500 5780
rect 15100 5500 15500 5620
rect 15900 5780 16300 5900
rect 15900 5620 16020 5780
rect 16180 5620 16300 5780
rect 15900 5500 16300 5620
rect 700 4980 1100 5100
rect 700 4820 820 4980
rect 980 4820 1100 4980
rect 700 4700 1100 4820
rect 1500 4980 1900 5100
rect 1500 4820 1620 4980
rect 1780 4820 1900 4980
rect 1500 4700 1900 4820
rect 2300 4980 2700 5100
rect 2300 4820 2420 4980
rect 2580 4820 2700 4980
rect 2300 4700 2700 4820
rect 3100 4980 3500 5100
rect 3100 4820 3220 4980
rect 3380 4820 3500 4980
rect 3100 4700 3500 4820
rect 3900 4980 4300 5100
rect 3900 4820 4020 4980
rect 4180 4820 4300 4980
rect 3900 4700 4300 4820
rect 4700 4980 5100 5100
rect 4700 4820 4820 4980
rect 4980 4820 5100 4980
rect 4700 4700 5100 4820
rect 5500 4980 5900 5100
rect 5500 4820 5620 4980
rect 5780 4820 5900 4980
rect 5500 4700 5900 4820
rect 6300 4980 6700 5100
rect 6300 4820 6420 4980
rect 6580 4820 6700 4980
rect 6300 4700 6700 4820
rect 7100 4980 7500 5100
rect 7100 4820 7220 4980
rect 7380 4820 7500 4980
rect 7100 4700 7500 4820
rect 7900 4980 8300 5100
rect 7900 4820 8020 4980
rect 8180 4820 8300 4980
rect 7900 4700 8300 4820
rect 8700 4980 9100 5100
rect 8700 4820 8820 4980
rect 8980 4820 9100 4980
rect 8700 4700 9100 4820
rect 9500 4980 9900 5100
rect 9500 4820 9620 4980
rect 9780 4820 9900 4980
rect 9500 4700 9900 4820
rect 10300 4980 10700 5100
rect 10300 4820 10420 4980
rect 10580 4820 10700 4980
rect 10300 4700 10700 4820
rect 11100 4980 11500 5100
rect 11100 4820 11220 4980
rect 11380 4820 11500 4980
rect 11100 4700 11500 4820
rect 11900 4980 12300 5100
rect 11900 4820 12020 4980
rect 12180 4820 12300 4980
rect 11900 4700 12300 4820
rect 12700 4980 13100 5100
rect 12700 4820 12820 4980
rect 12980 4820 13100 4980
rect 12700 4700 13100 4820
rect 13500 4980 13900 5100
rect 13500 4820 13620 4980
rect 13780 4820 13900 4980
rect 13500 4700 13900 4820
rect 14300 4980 14700 5100
rect 14300 4820 14420 4980
rect 14580 4820 14700 4980
rect 14300 4700 14700 4820
rect 15100 4980 15500 5100
rect 15100 4820 15220 4980
rect 15380 4820 15500 4980
rect 15100 4700 15500 4820
rect 15900 4980 16300 5100
rect 15900 4820 16020 4980
rect 16180 4820 16300 4980
rect 15900 4700 16300 4820
rect 700 4180 1100 4300
rect 700 4020 820 4180
rect 980 4020 1100 4180
rect 700 3900 1100 4020
rect 1500 4180 1900 4300
rect 1500 4020 1620 4180
rect 1780 4020 1900 4180
rect 1500 3900 1900 4020
rect 2300 4180 2700 4300
rect 2300 4020 2420 4180
rect 2580 4020 2700 4180
rect 2300 3900 2700 4020
rect 3100 4180 3500 4300
rect 3100 4020 3220 4180
rect 3380 4020 3500 4180
rect 3100 3900 3500 4020
rect 3900 4180 4300 4300
rect 3900 4020 4020 4180
rect 4180 4020 4300 4180
rect 3900 3900 4300 4020
rect 4700 4180 5100 4300
rect 4700 4020 4820 4180
rect 4980 4020 5100 4180
rect 4700 3900 5100 4020
rect 5500 4180 5900 4300
rect 5500 4020 5620 4180
rect 5780 4020 5900 4180
rect 5500 3900 5900 4020
rect 6300 4180 6700 4300
rect 6300 4020 6420 4180
rect 6580 4020 6700 4180
rect 6300 3900 6700 4020
rect 7100 4180 7500 4300
rect 7100 4020 7220 4180
rect 7380 4020 7500 4180
rect 7100 3900 7500 4020
rect 7900 4180 8300 4300
rect 7900 4020 8020 4180
rect 8180 4020 8300 4180
rect 7900 3900 8300 4020
rect 8700 4180 9100 4300
rect 8700 4020 8820 4180
rect 8980 4020 9100 4180
rect 8700 3900 9100 4020
rect 9500 4180 9900 4300
rect 9500 4020 9620 4180
rect 9780 4020 9900 4180
rect 9500 3900 9900 4020
rect 10300 4180 10700 4300
rect 10300 4020 10420 4180
rect 10580 4020 10700 4180
rect 10300 3900 10700 4020
rect 11100 4180 11500 4300
rect 11100 4020 11220 4180
rect 11380 4020 11500 4180
rect 11100 3900 11500 4020
rect 11900 4180 12300 4300
rect 11900 4020 12020 4180
rect 12180 4020 12300 4180
rect 11900 3900 12300 4020
rect 12700 4180 13100 4300
rect 12700 4020 12820 4180
rect 12980 4020 13100 4180
rect 12700 3900 13100 4020
rect 13500 4180 13900 4300
rect 13500 4020 13620 4180
rect 13780 4020 13900 4180
rect 13500 3900 13900 4020
rect 14300 4180 14700 4300
rect 14300 4020 14420 4180
rect 14580 4020 14700 4180
rect 14300 3900 14700 4020
rect 15100 4180 15500 4300
rect 15100 4020 15220 4180
rect 15380 4020 15500 4180
rect 15100 3900 15500 4020
rect 15900 4180 16300 4300
rect 15900 4020 16020 4180
rect 16180 4020 16300 4180
rect 15900 3900 16300 4020
rect 700 3380 1100 3500
rect 700 3220 820 3380
rect 980 3220 1100 3380
rect 700 3100 1100 3220
rect 1500 3380 1900 3500
rect 1500 3220 1620 3380
rect 1780 3220 1900 3380
rect 1500 3100 1900 3220
rect 2300 3380 2700 3500
rect 2300 3220 2420 3380
rect 2580 3220 2700 3380
rect 2300 3100 2700 3220
rect 3100 3380 3500 3500
rect 3100 3220 3220 3380
rect 3380 3220 3500 3380
rect 3100 3100 3500 3220
rect 3900 3380 4300 3500
rect 3900 3220 4020 3380
rect 4180 3220 4300 3380
rect 3900 3100 4300 3220
rect 4700 3380 5100 3500
rect 4700 3220 4820 3380
rect 4980 3220 5100 3380
rect 4700 3100 5100 3220
rect 5500 3380 5900 3500
rect 5500 3220 5620 3380
rect 5780 3220 5900 3380
rect 5500 3100 5900 3220
rect 6300 3380 6700 3500
rect 6300 3220 6420 3380
rect 6580 3220 6700 3380
rect 6300 3100 6700 3220
rect 7100 3380 7500 3500
rect 7100 3220 7220 3380
rect 7380 3220 7500 3380
rect 7100 3100 7500 3220
rect 7900 3380 8300 3500
rect 7900 3220 8020 3380
rect 8180 3220 8300 3380
rect 7900 3100 8300 3220
rect 8700 3380 9100 3500
rect 8700 3220 8820 3380
rect 8980 3220 9100 3380
rect 8700 3100 9100 3220
rect 9500 3380 9900 3500
rect 9500 3220 9620 3380
rect 9780 3220 9900 3380
rect 9500 3100 9900 3220
rect 10300 3380 10700 3500
rect 10300 3220 10420 3380
rect 10580 3220 10700 3380
rect 10300 3100 10700 3220
rect 11100 3380 11500 3500
rect 11100 3220 11220 3380
rect 11380 3220 11500 3380
rect 11100 3100 11500 3220
rect 11900 3380 12300 3500
rect 11900 3220 12020 3380
rect 12180 3220 12300 3380
rect 11900 3100 12300 3220
rect 12700 3380 13100 3500
rect 12700 3220 12820 3380
rect 12980 3220 13100 3380
rect 12700 3100 13100 3220
rect 13500 3380 13900 3500
rect 13500 3220 13620 3380
rect 13780 3220 13900 3380
rect 13500 3100 13900 3220
rect 14300 3380 14700 3500
rect 14300 3220 14420 3380
rect 14580 3220 14700 3380
rect 14300 3100 14700 3220
rect 15100 3380 15500 3500
rect 15100 3220 15220 3380
rect 15380 3220 15500 3380
rect 15100 3100 15500 3220
rect 15900 3380 16300 3500
rect 15900 3220 16020 3380
rect 16180 3220 16300 3380
rect 15900 3100 16300 3220
rect 700 2580 1100 2700
rect 700 2420 820 2580
rect 980 2420 1100 2580
rect 700 2300 1100 2420
rect 1500 2580 1900 2700
rect 1500 2420 1620 2580
rect 1780 2420 1900 2580
rect 1500 2300 1900 2420
rect 2300 2580 2700 2700
rect 2300 2420 2420 2580
rect 2580 2420 2700 2580
rect 2300 2300 2700 2420
rect 3100 2580 3500 2700
rect 3100 2420 3220 2580
rect 3380 2420 3500 2580
rect 3100 2300 3500 2420
rect 3900 2580 4300 2700
rect 3900 2420 4020 2580
rect 4180 2420 4300 2580
rect 3900 2300 4300 2420
rect 4700 2580 5100 2700
rect 4700 2420 4820 2580
rect 4980 2420 5100 2580
rect 4700 2300 5100 2420
rect 5500 2580 5900 2700
rect 5500 2420 5620 2580
rect 5780 2420 5900 2580
rect 5500 2300 5900 2420
rect 6300 2580 6700 2700
rect 6300 2420 6420 2580
rect 6580 2420 6700 2580
rect 6300 2300 6700 2420
rect 7100 2580 7500 2700
rect 7100 2420 7220 2580
rect 7380 2420 7500 2580
rect 7100 2300 7500 2420
rect 7900 2580 8300 2700
rect 7900 2420 8020 2580
rect 8180 2420 8300 2580
rect 7900 2300 8300 2420
rect 8700 2580 9100 2700
rect 8700 2420 8820 2580
rect 8980 2420 9100 2580
rect 8700 2300 9100 2420
rect 9500 2580 9900 2700
rect 9500 2420 9620 2580
rect 9780 2420 9900 2580
rect 9500 2300 9900 2420
rect 10300 2580 10700 2700
rect 10300 2420 10420 2580
rect 10580 2420 10700 2580
rect 10300 2300 10700 2420
rect 11100 2580 11500 2700
rect 11100 2420 11220 2580
rect 11380 2420 11500 2580
rect 11100 2300 11500 2420
rect 11900 2580 12300 2700
rect 11900 2420 12020 2580
rect 12180 2420 12300 2580
rect 11900 2300 12300 2420
rect 12700 2580 13100 2700
rect 12700 2420 12820 2580
rect 12980 2420 13100 2580
rect 12700 2300 13100 2420
rect 13500 2580 13900 2700
rect 13500 2420 13620 2580
rect 13780 2420 13900 2580
rect 13500 2300 13900 2420
rect 14300 2580 14700 2700
rect 14300 2420 14420 2580
rect 14580 2420 14700 2580
rect 14300 2300 14700 2420
rect 15100 2580 15500 2700
rect 15100 2420 15220 2580
rect 15380 2420 15500 2580
rect 15100 2300 15500 2420
rect 15900 2580 16300 2700
rect 15900 2420 16020 2580
rect 16180 2420 16300 2580
rect 15900 2300 16300 2420
rect 700 1780 1100 1900
rect 700 1620 820 1780
rect 980 1620 1100 1780
rect 700 1500 1100 1620
rect 1500 1780 1900 1900
rect 1500 1620 1620 1780
rect 1780 1620 1900 1780
rect 1500 1500 1900 1620
rect 2300 1780 2700 1900
rect 2300 1620 2420 1780
rect 2580 1620 2700 1780
rect 2300 1500 2700 1620
rect 3100 1780 3500 1900
rect 3100 1620 3220 1780
rect 3380 1620 3500 1780
rect 3100 1500 3500 1620
rect 3900 1780 4300 1900
rect 3900 1620 4020 1780
rect 4180 1620 4300 1780
rect 3900 1500 4300 1620
rect 4700 1780 5100 1900
rect 4700 1620 4820 1780
rect 4980 1620 5100 1780
rect 4700 1500 5100 1620
rect 5500 1780 5900 1900
rect 5500 1620 5620 1780
rect 5780 1620 5900 1780
rect 5500 1500 5900 1620
rect 6300 1780 6700 1900
rect 6300 1620 6420 1780
rect 6580 1620 6700 1780
rect 6300 1500 6700 1620
rect 7100 1780 7500 1900
rect 7100 1620 7220 1780
rect 7380 1620 7500 1780
rect 7100 1500 7500 1620
rect 7900 1780 8300 1900
rect 7900 1620 8020 1780
rect 8180 1620 8300 1780
rect 7900 1500 8300 1620
rect 8700 1780 9100 1900
rect 8700 1620 8820 1780
rect 8980 1620 9100 1780
rect 8700 1500 9100 1620
rect 9500 1780 9900 1900
rect 9500 1620 9620 1780
rect 9780 1620 9900 1780
rect 9500 1500 9900 1620
rect 10300 1780 10700 1900
rect 10300 1620 10420 1780
rect 10580 1620 10700 1780
rect 10300 1500 10700 1620
rect 11100 1780 11500 1900
rect 11100 1620 11220 1780
rect 11380 1620 11500 1780
rect 11100 1500 11500 1620
rect 11900 1780 12300 1900
rect 11900 1620 12020 1780
rect 12180 1620 12300 1780
rect 11900 1500 12300 1620
rect 12700 1780 13100 1900
rect 12700 1620 12820 1780
rect 12980 1620 13100 1780
rect 12700 1500 13100 1620
rect 13500 1780 13900 1900
rect 13500 1620 13620 1780
rect 13780 1620 13900 1780
rect 13500 1500 13900 1620
rect 14300 1780 14700 1900
rect 14300 1620 14420 1780
rect 14580 1620 14700 1780
rect 14300 1500 14700 1620
rect 15100 1780 15500 1900
rect 15100 1620 15220 1780
rect 15380 1620 15500 1780
rect 15100 1500 15500 1620
rect 15900 1780 16300 1900
rect 15900 1620 16020 1780
rect 16180 1620 16300 1780
rect 15900 1500 16300 1620
rect 700 980 1100 1100
rect 700 820 820 980
rect 980 820 1100 980
rect 700 700 1100 820
rect 1500 980 1900 1100
rect 1500 820 1620 980
rect 1780 820 1900 980
rect 1500 700 1900 820
rect 2300 980 2700 1100
rect 2300 820 2420 980
rect 2580 820 2700 980
rect 2300 700 2700 820
rect 3100 980 3500 1100
rect 3100 820 3220 980
rect 3380 820 3500 980
rect 3100 700 3500 820
rect 3900 980 4300 1100
rect 3900 820 4020 980
rect 4180 820 4300 980
rect 3900 700 4300 820
rect 4700 980 5100 1100
rect 4700 820 4820 980
rect 4980 820 5100 980
rect 4700 700 5100 820
rect 5500 980 5900 1100
rect 5500 820 5620 980
rect 5780 820 5900 980
rect 5500 700 5900 820
rect 6300 980 6700 1100
rect 6300 820 6420 980
rect 6580 820 6700 980
rect 6300 700 6700 820
rect 7100 980 7500 1100
rect 7100 820 7220 980
rect 7380 820 7500 980
rect 7100 700 7500 820
rect 7900 980 8300 1100
rect 7900 820 8020 980
rect 8180 820 8300 980
rect 7900 700 8300 820
rect 8700 980 9100 1100
rect 8700 820 8820 980
rect 8980 820 9100 980
rect 8700 700 9100 820
rect 9500 980 9900 1100
rect 9500 820 9620 980
rect 9780 820 9900 980
rect 9500 700 9900 820
rect 10300 980 10700 1100
rect 10300 820 10420 980
rect 10580 820 10700 980
rect 10300 700 10700 820
rect 11100 980 11500 1100
rect 11100 820 11220 980
rect 11380 820 11500 980
rect 11100 700 11500 820
rect 11900 980 12300 1100
rect 11900 820 12020 980
rect 12180 820 12300 980
rect 11900 700 12300 820
rect 12700 980 13100 1100
rect 12700 820 12820 980
rect 12980 820 13100 980
rect 12700 700 13100 820
rect 13500 980 13900 1100
rect 13500 820 13620 980
rect 13780 820 13900 980
rect 13500 700 13900 820
rect 14300 980 14700 1100
rect 14300 820 14420 980
rect 14580 820 14700 980
rect 14300 700 14700 820
rect 15100 980 15500 1100
rect 15100 820 15220 980
rect 15380 820 15500 980
rect 15100 700 15500 820
rect 15900 980 16300 1100
rect 15900 820 16020 980
rect 16180 820 16300 980
rect 15900 700 16300 820
rect 16500 500 17000 16500
rect 0 0 17000 500
<< m2contact >>
rect 820 16020 980 16180
rect 1620 16020 1780 16180
rect 2420 16020 2580 16180
rect 3220 16020 3380 16180
rect 4020 16020 4180 16180
rect 4820 16020 4980 16180
rect 5620 16020 5780 16180
rect 6420 16020 6580 16180
rect 7220 16020 7380 16180
rect 8020 16020 8180 16180
rect 8820 16020 8980 16180
rect 9620 16020 9780 16180
rect 10420 16020 10580 16180
rect 11220 16020 11380 16180
rect 12020 16020 12180 16180
rect 12820 16020 12980 16180
rect 13620 16020 13780 16180
rect 14420 16020 14580 16180
rect 15220 16020 15380 16180
rect 16020 16020 16180 16180
rect 820 15220 980 15380
rect 1620 15220 1780 15380
rect 2420 15220 2580 15380
rect 3220 15220 3380 15380
rect 4020 15220 4180 15380
rect 4820 15220 4980 15380
rect 5620 15220 5780 15380
rect 6420 15220 6580 15380
rect 7220 15220 7380 15380
rect 8020 15220 8180 15380
rect 8820 15220 8980 15380
rect 9620 15220 9780 15380
rect 10420 15220 10580 15380
rect 11220 15220 11380 15380
rect 12020 15220 12180 15380
rect 12820 15220 12980 15380
rect 13620 15220 13780 15380
rect 14420 15220 14580 15380
rect 15220 15220 15380 15380
rect 16020 15220 16180 15380
rect 820 14420 980 14580
rect 1620 14420 1780 14580
rect 2420 14420 2580 14580
rect 3220 14420 3380 14580
rect 4020 14420 4180 14580
rect 4820 14420 4980 14580
rect 5620 14420 5780 14580
rect 6420 14420 6580 14580
rect 7220 14420 7380 14580
rect 8020 14420 8180 14580
rect 8820 14420 8980 14580
rect 9620 14420 9780 14580
rect 10420 14420 10580 14580
rect 11220 14420 11380 14580
rect 12020 14420 12180 14580
rect 12820 14420 12980 14580
rect 13620 14420 13780 14580
rect 14420 14420 14580 14580
rect 15220 14420 15380 14580
rect 16020 14420 16180 14580
rect 820 13620 980 13780
rect 1620 13620 1780 13780
rect 2420 13620 2580 13780
rect 3220 13620 3380 13780
rect 4020 13620 4180 13780
rect 4820 13620 4980 13780
rect 5620 13620 5780 13780
rect 6420 13620 6580 13780
rect 7220 13620 7380 13780
rect 8020 13620 8180 13780
rect 8820 13620 8980 13780
rect 9620 13620 9780 13780
rect 10420 13620 10580 13780
rect 11220 13620 11380 13780
rect 12020 13620 12180 13780
rect 12820 13620 12980 13780
rect 13620 13620 13780 13780
rect 14420 13620 14580 13780
rect 15220 13620 15380 13780
rect 16020 13620 16180 13780
rect 820 12820 980 12980
rect 1620 12820 1780 12980
rect 2420 12820 2580 12980
rect 3220 12820 3380 12980
rect 4020 12820 4180 12980
rect 4820 12820 4980 12980
rect 5620 12820 5780 12980
rect 6420 12820 6580 12980
rect 7220 12820 7380 12980
rect 8020 12820 8180 12980
rect 8820 12820 8980 12980
rect 9620 12820 9780 12980
rect 10420 12820 10580 12980
rect 11220 12820 11380 12980
rect 12020 12820 12180 12980
rect 12820 12820 12980 12980
rect 13620 12820 13780 12980
rect 14420 12820 14580 12980
rect 15220 12820 15380 12980
rect 16020 12820 16180 12980
rect 820 12020 980 12180
rect 1620 12020 1780 12180
rect 2420 12020 2580 12180
rect 3220 12020 3380 12180
rect 4020 12020 4180 12180
rect 4820 12020 4980 12180
rect 5620 12020 5780 12180
rect 6420 12020 6580 12180
rect 7220 12020 7380 12180
rect 8020 12020 8180 12180
rect 8820 12020 8980 12180
rect 9620 12020 9780 12180
rect 10420 12020 10580 12180
rect 11220 12020 11380 12180
rect 12020 12020 12180 12180
rect 12820 12020 12980 12180
rect 13620 12020 13780 12180
rect 14420 12020 14580 12180
rect 15220 12020 15380 12180
rect 16020 12020 16180 12180
rect 820 11220 980 11380
rect 1620 11220 1780 11380
rect 2420 11220 2580 11380
rect 3220 11220 3380 11380
rect 4020 11220 4180 11380
rect 4820 11220 4980 11380
rect 5620 11220 5780 11380
rect 6420 11220 6580 11380
rect 7220 11220 7380 11380
rect 8020 11220 8180 11380
rect 8820 11220 8980 11380
rect 9620 11220 9780 11380
rect 10420 11220 10580 11380
rect 11220 11220 11380 11380
rect 12020 11220 12180 11380
rect 12820 11220 12980 11380
rect 13620 11220 13780 11380
rect 14420 11220 14580 11380
rect 15220 11220 15380 11380
rect 16020 11220 16180 11380
rect 820 10420 980 10580
rect 1620 10420 1780 10580
rect 2420 10420 2580 10580
rect 3220 10420 3380 10580
rect 4020 10420 4180 10580
rect 4820 10420 4980 10580
rect 5620 10420 5780 10580
rect 6420 10420 6580 10580
rect 7220 10420 7380 10580
rect 8020 10420 8180 10580
rect 8820 10420 8980 10580
rect 9620 10420 9780 10580
rect 10420 10420 10580 10580
rect 11220 10420 11380 10580
rect 12020 10420 12180 10580
rect 12820 10420 12980 10580
rect 13620 10420 13780 10580
rect 14420 10420 14580 10580
rect 15220 10420 15380 10580
rect 16020 10420 16180 10580
rect 820 9620 980 9780
rect 1620 9620 1780 9780
rect 2420 9620 2580 9780
rect 3220 9620 3380 9780
rect 4020 9620 4180 9780
rect 4820 9620 4980 9780
rect 5620 9620 5780 9780
rect 6420 9620 6580 9780
rect 7220 9620 7380 9780
rect 8020 9620 8180 9780
rect 8820 9620 8980 9780
rect 9620 9620 9780 9780
rect 10420 9620 10580 9780
rect 11220 9620 11380 9780
rect 12020 9620 12180 9780
rect 12820 9620 12980 9780
rect 13620 9620 13780 9780
rect 14420 9620 14580 9780
rect 15220 9620 15380 9780
rect 16020 9620 16180 9780
rect 820 8820 980 8980
rect 1620 8820 1780 8980
rect 2420 8820 2580 8980
rect 3220 8820 3380 8980
rect 4020 8820 4180 8980
rect 4820 8820 4980 8980
rect 5620 8820 5780 8980
rect 6420 8820 6580 8980
rect 7220 8820 7380 8980
rect 8020 8820 8180 8980
rect 8820 8820 8980 8980
rect 9620 8820 9780 8980
rect 10420 8820 10580 8980
rect 11220 8820 11380 8980
rect 12020 8820 12180 8980
rect 12820 8820 12980 8980
rect 13620 8820 13780 8980
rect 14420 8820 14580 8980
rect 15220 8820 15380 8980
rect 16020 8820 16180 8980
rect 820 8020 980 8180
rect 1620 8020 1780 8180
rect 2420 8020 2580 8180
rect 3220 8020 3380 8180
rect 4020 8020 4180 8180
rect 4820 8020 4980 8180
rect 5620 8020 5780 8180
rect 6420 8020 6580 8180
rect 7220 8020 7380 8180
rect 8020 8020 8180 8180
rect 8820 8020 8980 8180
rect 9620 8020 9780 8180
rect 10420 8020 10580 8180
rect 11220 8020 11380 8180
rect 12020 8020 12180 8180
rect 12820 8020 12980 8180
rect 13620 8020 13780 8180
rect 14420 8020 14580 8180
rect 15220 8020 15380 8180
rect 16020 8020 16180 8180
rect 820 7220 980 7380
rect 1620 7220 1780 7380
rect 2420 7220 2580 7380
rect 3220 7220 3380 7380
rect 4020 7220 4180 7380
rect 4820 7220 4980 7380
rect 5620 7220 5780 7380
rect 6420 7220 6580 7380
rect 7220 7220 7380 7380
rect 8020 7220 8180 7380
rect 8820 7220 8980 7380
rect 9620 7220 9780 7380
rect 10420 7220 10580 7380
rect 11220 7220 11380 7380
rect 12020 7220 12180 7380
rect 12820 7220 12980 7380
rect 13620 7220 13780 7380
rect 14420 7220 14580 7380
rect 15220 7220 15380 7380
rect 16020 7220 16180 7380
rect 820 6420 980 6580
rect 1620 6420 1780 6580
rect 2420 6420 2580 6580
rect 3220 6420 3380 6580
rect 4020 6420 4180 6580
rect 4820 6420 4980 6580
rect 5620 6420 5780 6580
rect 6420 6420 6580 6580
rect 7220 6420 7380 6580
rect 8020 6420 8180 6580
rect 8820 6420 8980 6580
rect 9620 6420 9780 6580
rect 10420 6420 10580 6580
rect 11220 6420 11380 6580
rect 12020 6420 12180 6580
rect 12820 6420 12980 6580
rect 13620 6420 13780 6580
rect 14420 6420 14580 6580
rect 15220 6420 15380 6580
rect 16020 6420 16180 6580
rect 820 5620 980 5780
rect 1620 5620 1780 5780
rect 2420 5620 2580 5780
rect 3220 5620 3380 5780
rect 4020 5620 4180 5780
rect 4820 5620 4980 5780
rect 5620 5620 5780 5780
rect 6420 5620 6580 5780
rect 7220 5620 7380 5780
rect 8020 5620 8180 5780
rect 8820 5620 8980 5780
rect 9620 5620 9780 5780
rect 10420 5620 10580 5780
rect 11220 5620 11380 5780
rect 12020 5620 12180 5780
rect 12820 5620 12980 5780
rect 13620 5620 13780 5780
rect 14420 5620 14580 5780
rect 15220 5620 15380 5780
rect 16020 5620 16180 5780
rect 820 4820 980 4980
rect 1620 4820 1780 4980
rect 2420 4820 2580 4980
rect 3220 4820 3380 4980
rect 4020 4820 4180 4980
rect 4820 4820 4980 4980
rect 5620 4820 5780 4980
rect 6420 4820 6580 4980
rect 7220 4820 7380 4980
rect 8020 4820 8180 4980
rect 8820 4820 8980 4980
rect 9620 4820 9780 4980
rect 10420 4820 10580 4980
rect 11220 4820 11380 4980
rect 12020 4820 12180 4980
rect 12820 4820 12980 4980
rect 13620 4820 13780 4980
rect 14420 4820 14580 4980
rect 15220 4820 15380 4980
rect 16020 4820 16180 4980
rect 820 4020 980 4180
rect 1620 4020 1780 4180
rect 2420 4020 2580 4180
rect 3220 4020 3380 4180
rect 4020 4020 4180 4180
rect 4820 4020 4980 4180
rect 5620 4020 5780 4180
rect 6420 4020 6580 4180
rect 7220 4020 7380 4180
rect 8020 4020 8180 4180
rect 8820 4020 8980 4180
rect 9620 4020 9780 4180
rect 10420 4020 10580 4180
rect 11220 4020 11380 4180
rect 12020 4020 12180 4180
rect 12820 4020 12980 4180
rect 13620 4020 13780 4180
rect 14420 4020 14580 4180
rect 15220 4020 15380 4180
rect 16020 4020 16180 4180
rect 820 3220 980 3380
rect 1620 3220 1780 3380
rect 2420 3220 2580 3380
rect 3220 3220 3380 3380
rect 4020 3220 4180 3380
rect 4820 3220 4980 3380
rect 5620 3220 5780 3380
rect 6420 3220 6580 3380
rect 7220 3220 7380 3380
rect 8020 3220 8180 3380
rect 8820 3220 8980 3380
rect 9620 3220 9780 3380
rect 10420 3220 10580 3380
rect 11220 3220 11380 3380
rect 12020 3220 12180 3380
rect 12820 3220 12980 3380
rect 13620 3220 13780 3380
rect 14420 3220 14580 3380
rect 15220 3220 15380 3380
rect 16020 3220 16180 3380
rect 820 2420 980 2580
rect 1620 2420 1780 2580
rect 2420 2420 2580 2580
rect 3220 2420 3380 2580
rect 4020 2420 4180 2580
rect 4820 2420 4980 2580
rect 5620 2420 5780 2580
rect 6420 2420 6580 2580
rect 7220 2420 7380 2580
rect 8020 2420 8180 2580
rect 8820 2420 8980 2580
rect 9620 2420 9780 2580
rect 10420 2420 10580 2580
rect 11220 2420 11380 2580
rect 12020 2420 12180 2580
rect 12820 2420 12980 2580
rect 13620 2420 13780 2580
rect 14420 2420 14580 2580
rect 15220 2420 15380 2580
rect 16020 2420 16180 2580
rect 820 1620 980 1780
rect 1620 1620 1780 1780
rect 2420 1620 2580 1780
rect 3220 1620 3380 1780
rect 4020 1620 4180 1780
rect 4820 1620 4980 1780
rect 5620 1620 5780 1780
rect 6420 1620 6580 1780
rect 7220 1620 7380 1780
rect 8020 1620 8180 1780
rect 8820 1620 8980 1780
rect 9620 1620 9780 1780
rect 10420 1620 10580 1780
rect 11220 1620 11380 1780
rect 12020 1620 12180 1780
rect 12820 1620 12980 1780
rect 13620 1620 13780 1780
rect 14420 1620 14580 1780
rect 15220 1620 15380 1780
rect 16020 1620 16180 1780
rect 820 820 980 980
rect 1620 820 1780 980
rect 2420 820 2580 980
rect 3220 820 3380 980
rect 4020 820 4180 980
rect 4820 820 4980 980
rect 5620 820 5780 980
rect 6420 820 6580 980
rect 7220 820 7380 980
rect 8020 820 8180 980
rect 8820 820 8980 980
rect 9620 820 9780 980
rect 10420 820 10580 980
rect 11220 820 11380 980
rect 12020 820 12180 980
rect 12820 820 12980 980
rect 13620 820 13780 980
rect 14420 820 14580 980
rect 15220 820 15380 980
rect 16020 820 16180 980
<< metal2 >>
rect 0 16500 17000 17000
rect 0 500 500 16500
rect 700 16180 1100 16300
rect 700 16020 820 16180
rect 980 16020 1100 16180
rect 700 15900 1100 16020
rect 1500 16180 1900 16300
rect 1500 16020 1620 16180
rect 1780 16020 1900 16180
rect 1500 15900 1900 16020
rect 2300 16180 2700 16300
rect 2300 16020 2420 16180
rect 2580 16020 2700 16180
rect 2300 15900 2700 16020
rect 3100 16180 3500 16300
rect 3100 16020 3220 16180
rect 3380 16020 3500 16180
rect 3100 15900 3500 16020
rect 3900 16180 4300 16300
rect 3900 16020 4020 16180
rect 4180 16020 4300 16180
rect 3900 15900 4300 16020
rect 4700 16180 5100 16300
rect 4700 16020 4820 16180
rect 4980 16020 5100 16180
rect 4700 15900 5100 16020
rect 5500 16180 5900 16300
rect 5500 16020 5620 16180
rect 5780 16020 5900 16180
rect 5500 15900 5900 16020
rect 6300 16180 6700 16300
rect 6300 16020 6420 16180
rect 6580 16020 6700 16180
rect 6300 15900 6700 16020
rect 7100 16180 7500 16300
rect 7100 16020 7220 16180
rect 7380 16020 7500 16180
rect 7100 15900 7500 16020
rect 7900 16180 8300 16300
rect 7900 16020 8020 16180
rect 8180 16020 8300 16180
rect 7900 15900 8300 16020
rect 8700 16180 9100 16300
rect 8700 16020 8820 16180
rect 8980 16020 9100 16180
rect 8700 15900 9100 16020
rect 9500 16180 9900 16300
rect 9500 16020 9620 16180
rect 9780 16020 9900 16180
rect 9500 15900 9900 16020
rect 10300 16180 10700 16300
rect 10300 16020 10420 16180
rect 10580 16020 10700 16180
rect 10300 15900 10700 16020
rect 11100 16180 11500 16300
rect 11100 16020 11220 16180
rect 11380 16020 11500 16180
rect 11100 15900 11500 16020
rect 11900 16180 12300 16300
rect 11900 16020 12020 16180
rect 12180 16020 12300 16180
rect 11900 15900 12300 16020
rect 12700 16180 13100 16300
rect 12700 16020 12820 16180
rect 12980 16020 13100 16180
rect 12700 15900 13100 16020
rect 13500 16180 13900 16300
rect 13500 16020 13620 16180
rect 13780 16020 13900 16180
rect 13500 15900 13900 16020
rect 14300 16180 14700 16300
rect 14300 16020 14420 16180
rect 14580 16020 14700 16180
rect 14300 15900 14700 16020
rect 15100 16180 15500 16300
rect 15100 16020 15220 16180
rect 15380 16020 15500 16180
rect 15100 15900 15500 16020
rect 15900 16180 16300 16300
rect 15900 16020 16020 16180
rect 16180 16020 16300 16180
rect 15900 15900 16300 16020
rect 1100 15780 1500 15900
rect 1100 15620 1220 15780
rect 1380 15620 1500 15780
rect 1100 15500 1500 15620
rect 1900 15780 2300 15900
rect 1900 15620 2020 15780
rect 2180 15620 2300 15780
rect 1900 15500 2300 15620
rect 2700 15780 3100 15900
rect 2700 15620 2820 15780
rect 2980 15620 3100 15780
rect 2700 15500 3100 15620
rect 3500 15780 3900 15900
rect 3500 15620 3620 15780
rect 3780 15620 3900 15780
rect 3500 15500 3900 15620
rect 4300 15780 4700 15900
rect 4300 15620 4420 15780
rect 4580 15620 4700 15780
rect 4300 15500 4700 15620
rect 5100 15780 5500 15900
rect 5100 15620 5220 15780
rect 5380 15620 5500 15780
rect 5100 15500 5500 15620
rect 5900 15780 6300 15900
rect 5900 15620 6020 15780
rect 6180 15620 6300 15780
rect 5900 15500 6300 15620
rect 6700 15780 7100 15900
rect 6700 15620 6820 15780
rect 6980 15620 7100 15780
rect 6700 15500 7100 15620
rect 7500 15780 7900 15900
rect 7500 15620 7620 15780
rect 7780 15620 7900 15780
rect 7500 15500 7900 15620
rect 8300 15780 8700 15900
rect 8300 15620 8420 15780
rect 8580 15620 8700 15780
rect 8300 15500 8700 15620
rect 9100 15780 9500 15900
rect 9100 15620 9220 15780
rect 9380 15620 9500 15780
rect 9100 15500 9500 15620
rect 9900 15780 10300 15900
rect 9900 15620 10020 15780
rect 10180 15620 10300 15780
rect 9900 15500 10300 15620
rect 10700 15780 11100 15900
rect 10700 15620 10820 15780
rect 10980 15620 11100 15780
rect 10700 15500 11100 15620
rect 11500 15780 11900 15900
rect 11500 15620 11620 15780
rect 11780 15620 11900 15780
rect 11500 15500 11900 15620
rect 12300 15780 12700 15900
rect 12300 15620 12420 15780
rect 12580 15620 12700 15780
rect 12300 15500 12700 15620
rect 13100 15780 13500 15900
rect 13100 15620 13220 15780
rect 13380 15620 13500 15780
rect 13100 15500 13500 15620
rect 13900 15780 14300 15900
rect 13900 15620 14020 15780
rect 14180 15620 14300 15780
rect 13900 15500 14300 15620
rect 14700 15780 15100 15900
rect 14700 15620 14820 15780
rect 14980 15620 15100 15780
rect 14700 15500 15100 15620
rect 15500 15780 15900 15900
rect 15500 15620 15620 15780
rect 15780 15620 15900 15780
rect 15500 15500 15900 15620
rect 700 15380 1100 15500
rect 700 15220 820 15380
rect 980 15220 1100 15380
rect 700 15100 1100 15220
rect 1500 15380 1900 15500
rect 1500 15220 1620 15380
rect 1780 15220 1900 15380
rect 1500 15100 1900 15220
rect 2300 15380 2700 15500
rect 2300 15220 2420 15380
rect 2580 15220 2700 15380
rect 2300 15100 2700 15220
rect 3100 15380 3500 15500
rect 3100 15220 3220 15380
rect 3380 15220 3500 15380
rect 3100 15100 3500 15220
rect 3900 15380 4300 15500
rect 3900 15220 4020 15380
rect 4180 15220 4300 15380
rect 3900 15100 4300 15220
rect 4700 15380 5100 15500
rect 4700 15220 4820 15380
rect 4980 15220 5100 15380
rect 4700 15100 5100 15220
rect 5500 15380 5900 15500
rect 5500 15220 5620 15380
rect 5780 15220 5900 15380
rect 5500 15100 5900 15220
rect 6300 15380 6700 15500
rect 6300 15220 6420 15380
rect 6580 15220 6700 15380
rect 6300 15100 6700 15220
rect 7100 15380 7500 15500
rect 7100 15220 7220 15380
rect 7380 15220 7500 15380
rect 7100 15100 7500 15220
rect 7900 15380 8300 15500
rect 7900 15220 8020 15380
rect 8180 15220 8300 15380
rect 7900 15100 8300 15220
rect 8700 15380 9100 15500
rect 8700 15220 8820 15380
rect 8980 15220 9100 15380
rect 8700 15100 9100 15220
rect 9500 15380 9900 15500
rect 9500 15220 9620 15380
rect 9780 15220 9900 15380
rect 9500 15100 9900 15220
rect 10300 15380 10700 15500
rect 10300 15220 10420 15380
rect 10580 15220 10700 15380
rect 10300 15100 10700 15220
rect 11100 15380 11500 15500
rect 11100 15220 11220 15380
rect 11380 15220 11500 15380
rect 11100 15100 11500 15220
rect 11900 15380 12300 15500
rect 11900 15220 12020 15380
rect 12180 15220 12300 15380
rect 11900 15100 12300 15220
rect 12700 15380 13100 15500
rect 12700 15220 12820 15380
rect 12980 15220 13100 15380
rect 12700 15100 13100 15220
rect 13500 15380 13900 15500
rect 13500 15220 13620 15380
rect 13780 15220 13900 15380
rect 13500 15100 13900 15220
rect 14300 15380 14700 15500
rect 14300 15220 14420 15380
rect 14580 15220 14700 15380
rect 14300 15100 14700 15220
rect 15100 15380 15500 15500
rect 15100 15220 15220 15380
rect 15380 15220 15500 15380
rect 15100 15100 15500 15220
rect 15900 15380 16300 15500
rect 15900 15220 16020 15380
rect 16180 15220 16300 15380
rect 15900 15100 16300 15220
rect 1100 14980 1500 15100
rect 1100 14820 1220 14980
rect 1380 14820 1500 14980
rect 1100 14700 1500 14820
rect 1900 14980 2300 15100
rect 1900 14820 2020 14980
rect 2180 14820 2300 14980
rect 1900 14700 2300 14820
rect 2700 14980 3100 15100
rect 2700 14820 2820 14980
rect 2980 14820 3100 14980
rect 2700 14700 3100 14820
rect 3500 14980 3900 15100
rect 3500 14820 3620 14980
rect 3780 14820 3900 14980
rect 3500 14700 3900 14820
rect 4300 14980 4700 15100
rect 4300 14820 4420 14980
rect 4580 14820 4700 14980
rect 4300 14700 4700 14820
rect 5100 14980 5500 15100
rect 5100 14820 5220 14980
rect 5380 14820 5500 14980
rect 5100 14700 5500 14820
rect 5900 14980 6300 15100
rect 5900 14820 6020 14980
rect 6180 14820 6300 14980
rect 5900 14700 6300 14820
rect 6700 14980 7100 15100
rect 6700 14820 6820 14980
rect 6980 14820 7100 14980
rect 6700 14700 7100 14820
rect 7500 14980 7900 15100
rect 7500 14820 7620 14980
rect 7780 14820 7900 14980
rect 7500 14700 7900 14820
rect 8300 14980 8700 15100
rect 8300 14820 8420 14980
rect 8580 14820 8700 14980
rect 8300 14700 8700 14820
rect 9100 14980 9500 15100
rect 9100 14820 9220 14980
rect 9380 14820 9500 14980
rect 9100 14700 9500 14820
rect 9900 14980 10300 15100
rect 9900 14820 10020 14980
rect 10180 14820 10300 14980
rect 9900 14700 10300 14820
rect 10700 14980 11100 15100
rect 10700 14820 10820 14980
rect 10980 14820 11100 14980
rect 10700 14700 11100 14820
rect 11500 14980 11900 15100
rect 11500 14820 11620 14980
rect 11780 14820 11900 14980
rect 11500 14700 11900 14820
rect 12300 14980 12700 15100
rect 12300 14820 12420 14980
rect 12580 14820 12700 14980
rect 12300 14700 12700 14820
rect 13100 14980 13500 15100
rect 13100 14820 13220 14980
rect 13380 14820 13500 14980
rect 13100 14700 13500 14820
rect 13900 14980 14300 15100
rect 13900 14820 14020 14980
rect 14180 14820 14300 14980
rect 13900 14700 14300 14820
rect 14700 14980 15100 15100
rect 14700 14820 14820 14980
rect 14980 14820 15100 14980
rect 14700 14700 15100 14820
rect 15500 14980 15900 15100
rect 15500 14820 15620 14980
rect 15780 14820 15900 14980
rect 15500 14700 15900 14820
rect 700 14580 1100 14700
rect 700 14420 820 14580
rect 980 14420 1100 14580
rect 700 14300 1100 14420
rect 1500 14580 1900 14700
rect 1500 14420 1620 14580
rect 1780 14420 1900 14580
rect 1500 14300 1900 14420
rect 2300 14580 2700 14700
rect 2300 14420 2420 14580
rect 2580 14420 2700 14580
rect 2300 14300 2700 14420
rect 3100 14580 3500 14700
rect 3100 14420 3220 14580
rect 3380 14420 3500 14580
rect 3100 14300 3500 14420
rect 3900 14580 4300 14700
rect 3900 14420 4020 14580
rect 4180 14420 4300 14580
rect 3900 14300 4300 14420
rect 4700 14580 5100 14700
rect 4700 14420 4820 14580
rect 4980 14420 5100 14580
rect 4700 14300 5100 14420
rect 5500 14580 5900 14700
rect 5500 14420 5620 14580
rect 5780 14420 5900 14580
rect 5500 14300 5900 14420
rect 6300 14580 6700 14700
rect 6300 14420 6420 14580
rect 6580 14420 6700 14580
rect 6300 14300 6700 14420
rect 7100 14580 7500 14700
rect 7100 14420 7220 14580
rect 7380 14420 7500 14580
rect 7100 14300 7500 14420
rect 7900 14580 8300 14700
rect 7900 14420 8020 14580
rect 8180 14420 8300 14580
rect 7900 14300 8300 14420
rect 8700 14580 9100 14700
rect 8700 14420 8820 14580
rect 8980 14420 9100 14580
rect 8700 14300 9100 14420
rect 9500 14580 9900 14700
rect 9500 14420 9620 14580
rect 9780 14420 9900 14580
rect 9500 14300 9900 14420
rect 10300 14580 10700 14700
rect 10300 14420 10420 14580
rect 10580 14420 10700 14580
rect 10300 14300 10700 14420
rect 11100 14580 11500 14700
rect 11100 14420 11220 14580
rect 11380 14420 11500 14580
rect 11100 14300 11500 14420
rect 11900 14580 12300 14700
rect 11900 14420 12020 14580
rect 12180 14420 12300 14580
rect 11900 14300 12300 14420
rect 12700 14580 13100 14700
rect 12700 14420 12820 14580
rect 12980 14420 13100 14580
rect 12700 14300 13100 14420
rect 13500 14580 13900 14700
rect 13500 14420 13620 14580
rect 13780 14420 13900 14580
rect 13500 14300 13900 14420
rect 14300 14580 14700 14700
rect 14300 14420 14420 14580
rect 14580 14420 14700 14580
rect 14300 14300 14700 14420
rect 15100 14580 15500 14700
rect 15100 14420 15220 14580
rect 15380 14420 15500 14580
rect 15100 14300 15500 14420
rect 15900 14580 16300 14700
rect 15900 14420 16020 14580
rect 16180 14420 16300 14580
rect 15900 14300 16300 14420
rect 1100 14180 1500 14300
rect 1100 14020 1220 14180
rect 1380 14020 1500 14180
rect 1100 13900 1500 14020
rect 1900 14180 2300 14300
rect 1900 14020 2020 14180
rect 2180 14020 2300 14180
rect 1900 13900 2300 14020
rect 2700 14180 3100 14300
rect 2700 14020 2820 14180
rect 2980 14020 3100 14180
rect 2700 13900 3100 14020
rect 3500 14180 3900 14300
rect 3500 14020 3620 14180
rect 3780 14020 3900 14180
rect 3500 13900 3900 14020
rect 4300 14180 4700 14300
rect 4300 14020 4420 14180
rect 4580 14020 4700 14180
rect 4300 13900 4700 14020
rect 5100 14180 5500 14300
rect 5100 14020 5220 14180
rect 5380 14020 5500 14180
rect 5100 13900 5500 14020
rect 5900 14180 6300 14300
rect 5900 14020 6020 14180
rect 6180 14020 6300 14180
rect 5900 13900 6300 14020
rect 6700 14180 7100 14300
rect 6700 14020 6820 14180
rect 6980 14020 7100 14180
rect 6700 13900 7100 14020
rect 7500 14180 7900 14300
rect 7500 14020 7620 14180
rect 7780 14020 7900 14180
rect 7500 13900 7900 14020
rect 8300 14180 8700 14300
rect 8300 14020 8420 14180
rect 8580 14020 8700 14180
rect 8300 13900 8700 14020
rect 9100 14180 9500 14300
rect 9100 14020 9220 14180
rect 9380 14020 9500 14180
rect 9100 13900 9500 14020
rect 9900 14180 10300 14300
rect 9900 14020 10020 14180
rect 10180 14020 10300 14180
rect 9900 13900 10300 14020
rect 10700 14180 11100 14300
rect 10700 14020 10820 14180
rect 10980 14020 11100 14180
rect 10700 13900 11100 14020
rect 11500 14180 11900 14300
rect 11500 14020 11620 14180
rect 11780 14020 11900 14180
rect 11500 13900 11900 14020
rect 12300 14180 12700 14300
rect 12300 14020 12420 14180
rect 12580 14020 12700 14180
rect 12300 13900 12700 14020
rect 13100 14180 13500 14300
rect 13100 14020 13220 14180
rect 13380 14020 13500 14180
rect 13100 13900 13500 14020
rect 13900 14180 14300 14300
rect 13900 14020 14020 14180
rect 14180 14020 14300 14180
rect 13900 13900 14300 14020
rect 14700 14180 15100 14300
rect 14700 14020 14820 14180
rect 14980 14020 15100 14180
rect 14700 13900 15100 14020
rect 15500 14180 15900 14300
rect 15500 14020 15620 14180
rect 15780 14020 15900 14180
rect 15500 13900 15900 14020
rect 700 13780 1100 13900
rect 700 13620 820 13780
rect 980 13620 1100 13780
rect 700 13500 1100 13620
rect 1500 13780 1900 13900
rect 1500 13620 1620 13780
rect 1780 13620 1900 13780
rect 1500 13500 1900 13620
rect 2300 13780 2700 13900
rect 2300 13620 2420 13780
rect 2580 13620 2700 13780
rect 2300 13500 2700 13620
rect 3100 13780 3500 13900
rect 3100 13620 3220 13780
rect 3380 13620 3500 13780
rect 3100 13500 3500 13620
rect 3900 13780 4300 13900
rect 3900 13620 4020 13780
rect 4180 13620 4300 13780
rect 3900 13500 4300 13620
rect 4700 13780 5100 13900
rect 4700 13620 4820 13780
rect 4980 13620 5100 13780
rect 4700 13500 5100 13620
rect 5500 13780 5900 13900
rect 5500 13620 5620 13780
rect 5780 13620 5900 13780
rect 5500 13500 5900 13620
rect 6300 13780 6700 13900
rect 6300 13620 6420 13780
rect 6580 13620 6700 13780
rect 6300 13500 6700 13620
rect 7100 13780 7500 13900
rect 7100 13620 7220 13780
rect 7380 13620 7500 13780
rect 7100 13500 7500 13620
rect 7900 13780 8300 13900
rect 7900 13620 8020 13780
rect 8180 13620 8300 13780
rect 7900 13500 8300 13620
rect 8700 13780 9100 13900
rect 8700 13620 8820 13780
rect 8980 13620 9100 13780
rect 8700 13500 9100 13620
rect 9500 13780 9900 13900
rect 9500 13620 9620 13780
rect 9780 13620 9900 13780
rect 9500 13500 9900 13620
rect 10300 13780 10700 13900
rect 10300 13620 10420 13780
rect 10580 13620 10700 13780
rect 10300 13500 10700 13620
rect 11100 13780 11500 13900
rect 11100 13620 11220 13780
rect 11380 13620 11500 13780
rect 11100 13500 11500 13620
rect 11900 13780 12300 13900
rect 11900 13620 12020 13780
rect 12180 13620 12300 13780
rect 11900 13500 12300 13620
rect 12700 13780 13100 13900
rect 12700 13620 12820 13780
rect 12980 13620 13100 13780
rect 12700 13500 13100 13620
rect 13500 13780 13900 13900
rect 13500 13620 13620 13780
rect 13780 13620 13900 13780
rect 13500 13500 13900 13620
rect 14300 13780 14700 13900
rect 14300 13620 14420 13780
rect 14580 13620 14700 13780
rect 14300 13500 14700 13620
rect 15100 13780 15500 13900
rect 15100 13620 15220 13780
rect 15380 13620 15500 13780
rect 15100 13500 15500 13620
rect 15900 13780 16300 13900
rect 15900 13620 16020 13780
rect 16180 13620 16300 13780
rect 15900 13500 16300 13620
rect 1100 13380 1500 13500
rect 1100 13220 1220 13380
rect 1380 13220 1500 13380
rect 1100 13100 1500 13220
rect 1900 13380 2300 13500
rect 1900 13220 2020 13380
rect 2180 13220 2300 13380
rect 1900 13100 2300 13220
rect 2700 13380 3100 13500
rect 2700 13220 2820 13380
rect 2980 13220 3100 13380
rect 2700 13100 3100 13220
rect 3500 13380 3900 13500
rect 3500 13220 3620 13380
rect 3780 13220 3900 13380
rect 3500 13100 3900 13220
rect 4300 13380 4700 13500
rect 4300 13220 4420 13380
rect 4580 13220 4700 13380
rect 4300 13100 4700 13220
rect 5100 13380 5500 13500
rect 5100 13220 5220 13380
rect 5380 13220 5500 13380
rect 5100 13100 5500 13220
rect 5900 13380 6300 13500
rect 5900 13220 6020 13380
rect 6180 13220 6300 13380
rect 5900 13100 6300 13220
rect 6700 13380 7100 13500
rect 6700 13220 6820 13380
rect 6980 13220 7100 13380
rect 6700 13100 7100 13220
rect 7500 13380 7900 13500
rect 7500 13220 7620 13380
rect 7780 13220 7900 13380
rect 7500 13100 7900 13220
rect 8300 13380 8700 13500
rect 8300 13220 8420 13380
rect 8580 13220 8700 13380
rect 8300 13100 8700 13220
rect 9100 13380 9500 13500
rect 9100 13220 9220 13380
rect 9380 13220 9500 13380
rect 9100 13100 9500 13220
rect 9900 13380 10300 13500
rect 9900 13220 10020 13380
rect 10180 13220 10300 13380
rect 9900 13100 10300 13220
rect 10700 13380 11100 13500
rect 10700 13220 10820 13380
rect 10980 13220 11100 13380
rect 10700 13100 11100 13220
rect 11500 13380 11900 13500
rect 11500 13220 11620 13380
rect 11780 13220 11900 13380
rect 11500 13100 11900 13220
rect 12300 13380 12700 13500
rect 12300 13220 12420 13380
rect 12580 13220 12700 13380
rect 12300 13100 12700 13220
rect 13100 13380 13500 13500
rect 13100 13220 13220 13380
rect 13380 13220 13500 13380
rect 13100 13100 13500 13220
rect 13900 13380 14300 13500
rect 13900 13220 14020 13380
rect 14180 13220 14300 13380
rect 13900 13100 14300 13220
rect 14700 13380 15100 13500
rect 14700 13220 14820 13380
rect 14980 13220 15100 13380
rect 14700 13100 15100 13220
rect 15500 13380 15900 13500
rect 15500 13220 15620 13380
rect 15780 13220 15900 13380
rect 15500 13100 15900 13220
rect 700 12980 1100 13100
rect 700 12820 820 12980
rect 980 12820 1100 12980
rect 700 12700 1100 12820
rect 1500 12980 1900 13100
rect 1500 12820 1620 12980
rect 1780 12820 1900 12980
rect 1500 12700 1900 12820
rect 2300 12980 2700 13100
rect 2300 12820 2420 12980
rect 2580 12820 2700 12980
rect 2300 12700 2700 12820
rect 3100 12980 3500 13100
rect 3100 12820 3220 12980
rect 3380 12820 3500 12980
rect 3100 12700 3500 12820
rect 3900 12980 4300 13100
rect 3900 12820 4020 12980
rect 4180 12820 4300 12980
rect 3900 12700 4300 12820
rect 4700 12980 5100 13100
rect 4700 12820 4820 12980
rect 4980 12820 5100 12980
rect 4700 12700 5100 12820
rect 5500 12980 5900 13100
rect 5500 12820 5620 12980
rect 5780 12820 5900 12980
rect 5500 12700 5900 12820
rect 6300 12980 6700 13100
rect 6300 12820 6420 12980
rect 6580 12820 6700 12980
rect 6300 12700 6700 12820
rect 7100 12980 7500 13100
rect 7100 12820 7220 12980
rect 7380 12820 7500 12980
rect 7100 12700 7500 12820
rect 7900 12980 8300 13100
rect 7900 12820 8020 12980
rect 8180 12820 8300 12980
rect 7900 12700 8300 12820
rect 8700 12980 9100 13100
rect 8700 12820 8820 12980
rect 8980 12820 9100 12980
rect 8700 12700 9100 12820
rect 9500 12980 9900 13100
rect 9500 12820 9620 12980
rect 9780 12820 9900 12980
rect 9500 12700 9900 12820
rect 10300 12980 10700 13100
rect 10300 12820 10420 12980
rect 10580 12820 10700 12980
rect 10300 12700 10700 12820
rect 11100 12980 11500 13100
rect 11100 12820 11220 12980
rect 11380 12820 11500 12980
rect 11100 12700 11500 12820
rect 11900 12980 12300 13100
rect 11900 12820 12020 12980
rect 12180 12820 12300 12980
rect 11900 12700 12300 12820
rect 12700 12980 13100 13100
rect 12700 12820 12820 12980
rect 12980 12820 13100 12980
rect 12700 12700 13100 12820
rect 13500 12980 13900 13100
rect 13500 12820 13620 12980
rect 13780 12820 13900 12980
rect 13500 12700 13900 12820
rect 14300 12980 14700 13100
rect 14300 12820 14420 12980
rect 14580 12820 14700 12980
rect 14300 12700 14700 12820
rect 15100 12980 15500 13100
rect 15100 12820 15220 12980
rect 15380 12820 15500 12980
rect 15100 12700 15500 12820
rect 15900 12980 16300 13100
rect 15900 12820 16020 12980
rect 16180 12820 16300 12980
rect 15900 12700 16300 12820
rect 1100 12580 1500 12700
rect 1100 12420 1220 12580
rect 1380 12420 1500 12580
rect 1100 12300 1500 12420
rect 1900 12580 2300 12700
rect 1900 12420 2020 12580
rect 2180 12420 2300 12580
rect 1900 12300 2300 12420
rect 2700 12580 3100 12700
rect 2700 12420 2820 12580
rect 2980 12420 3100 12580
rect 2700 12300 3100 12420
rect 3500 12580 3900 12700
rect 3500 12420 3620 12580
rect 3780 12420 3900 12580
rect 3500 12300 3900 12420
rect 4300 12580 4700 12700
rect 4300 12420 4420 12580
rect 4580 12420 4700 12580
rect 4300 12300 4700 12420
rect 5100 12580 5500 12700
rect 5100 12420 5220 12580
rect 5380 12420 5500 12580
rect 5100 12300 5500 12420
rect 5900 12580 6300 12700
rect 5900 12420 6020 12580
rect 6180 12420 6300 12580
rect 5900 12300 6300 12420
rect 6700 12580 7100 12700
rect 6700 12420 6820 12580
rect 6980 12420 7100 12580
rect 6700 12300 7100 12420
rect 7500 12580 7900 12700
rect 7500 12420 7620 12580
rect 7780 12420 7900 12580
rect 7500 12300 7900 12420
rect 8300 12580 8700 12700
rect 8300 12420 8420 12580
rect 8580 12420 8700 12580
rect 8300 12300 8700 12420
rect 9100 12580 9500 12700
rect 9100 12420 9220 12580
rect 9380 12420 9500 12580
rect 9100 12300 9500 12420
rect 9900 12580 10300 12700
rect 9900 12420 10020 12580
rect 10180 12420 10300 12580
rect 9900 12300 10300 12420
rect 10700 12580 11100 12700
rect 10700 12420 10820 12580
rect 10980 12420 11100 12580
rect 10700 12300 11100 12420
rect 11500 12580 11900 12700
rect 11500 12420 11620 12580
rect 11780 12420 11900 12580
rect 11500 12300 11900 12420
rect 12300 12580 12700 12700
rect 12300 12420 12420 12580
rect 12580 12420 12700 12580
rect 12300 12300 12700 12420
rect 13100 12580 13500 12700
rect 13100 12420 13220 12580
rect 13380 12420 13500 12580
rect 13100 12300 13500 12420
rect 13900 12580 14300 12700
rect 13900 12420 14020 12580
rect 14180 12420 14300 12580
rect 13900 12300 14300 12420
rect 14700 12580 15100 12700
rect 14700 12420 14820 12580
rect 14980 12420 15100 12580
rect 14700 12300 15100 12420
rect 15500 12580 15900 12700
rect 15500 12420 15620 12580
rect 15780 12420 15900 12580
rect 15500 12300 15900 12420
rect 700 12180 1100 12300
rect 700 12020 820 12180
rect 980 12020 1100 12180
rect 700 11900 1100 12020
rect 1500 12180 1900 12300
rect 1500 12020 1620 12180
rect 1780 12020 1900 12180
rect 1500 11900 1900 12020
rect 2300 12180 2700 12300
rect 2300 12020 2420 12180
rect 2580 12020 2700 12180
rect 2300 11900 2700 12020
rect 3100 12180 3500 12300
rect 3100 12020 3220 12180
rect 3380 12020 3500 12180
rect 3100 11900 3500 12020
rect 3900 12180 4300 12300
rect 3900 12020 4020 12180
rect 4180 12020 4300 12180
rect 3900 11900 4300 12020
rect 4700 12180 5100 12300
rect 4700 12020 4820 12180
rect 4980 12020 5100 12180
rect 4700 11900 5100 12020
rect 5500 12180 5900 12300
rect 5500 12020 5620 12180
rect 5780 12020 5900 12180
rect 5500 11900 5900 12020
rect 6300 12180 6700 12300
rect 6300 12020 6420 12180
rect 6580 12020 6700 12180
rect 6300 11900 6700 12020
rect 7100 12180 7500 12300
rect 7100 12020 7220 12180
rect 7380 12020 7500 12180
rect 7100 11900 7500 12020
rect 7900 12180 8300 12300
rect 7900 12020 8020 12180
rect 8180 12020 8300 12180
rect 7900 11900 8300 12020
rect 8700 12180 9100 12300
rect 8700 12020 8820 12180
rect 8980 12020 9100 12180
rect 8700 11900 9100 12020
rect 9500 12180 9900 12300
rect 9500 12020 9620 12180
rect 9780 12020 9900 12180
rect 9500 11900 9900 12020
rect 10300 12180 10700 12300
rect 10300 12020 10420 12180
rect 10580 12020 10700 12180
rect 10300 11900 10700 12020
rect 11100 12180 11500 12300
rect 11100 12020 11220 12180
rect 11380 12020 11500 12180
rect 11100 11900 11500 12020
rect 11900 12180 12300 12300
rect 11900 12020 12020 12180
rect 12180 12020 12300 12180
rect 11900 11900 12300 12020
rect 12700 12180 13100 12300
rect 12700 12020 12820 12180
rect 12980 12020 13100 12180
rect 12700 11900 13100 12020
rect 13500 12180 13900 12300
rect 13500 12020 13620 12180
rect 13780 12020 13900 12180
rect 13500 11900 13900 12020
rect 14300 12180 14700 12300
rect 14300 12020 14420 12180
rect 14580 12020 14700 12180
rect 14300 11900 14700 12020
rect 15100 12180 15500 12300
rect 15100 12020 15220 12180
rect 15380 12020 15500 12180
rect 15100 11900 15500 12020
rect 15900 12180 16300 12300
rect 15900 12020 16020 12180
rect 16180 12020 16300 12180
rect 15900 11900 16300 12020
rect 1100 11780 1500 11900
rect 1100 11620 1220 11780
rect 1380 11620 1500 11780
rect 1100 11500 1500 11620
rect 1900 11780 2300 11900
rect 1900 11620 2020 11780
rect 2180 11620 2300 11780
rect 1900 11500 2300 11620
rect 2700 11780 3100 11900
rect 2700 11620 2820 11780
rect 2980 11620 3100 11780
rect 2700 11500 3100 11620
rect 3500 11780 3900 11900
rect 3500 11620 3620 11780
rect 3780 11620 3900 11780
rect 3500 11500 3900 11620
rect 4300 11780 4700 11900
rect 4300 11620 4420 11780
rect 4580 11620 4700 11780
rect 4300 11500 4700 11620
rect 5100 11780 5500 11900
rect 5100 11620 5220 11780
rect 5380 11620 5500 11780
rect 5100 11500 5500 11620
rect 5900 11780 6300 11900
rect 5900 11620 6020 11780
rect 6180 11620 6300 11780
rect 5900 11500 6300 11620
rect 6700 11780 7100 11900
rect 6700 11620 6820 11780
rect 6980 11620 7100 11780
rect 6700 11500 7100 11620
rect 7500 11780 7900 11900
rect 7500 11620 7620 11780
rect 7780 11620 7900 11780
rect 7500 11500 7900 11620
rect 8300 11780 8700 11900
rect 8300 11620 8420 11780
rect 8580 11620 8700 11780
rect 8300 11500 8700 11620
rect 9100 11780 9500 11900
rect 9100 11620 9220 11780
rect 9380 11620 9500 11780
rect 9100 11500 9500 11620
rect 9900 11780 10300 11900
rect 9900 11620 10020 11780
rect 10180 11620 10300 11780
rect 9900 11500 10300 11620
rect 10700 11780 11100 11900
rect 10700 11620 10820 11780
rect 10980 11620 11100 11780
rect 10700 11500 11100 11620
rect 11500 11780 11900 11900
rect 11500 11620 11620 11780
rect 11780 11620 11900 11780
rect 11500 11500 11900 11620
rect 12300 11780 12700 11900
rect 12300 11620 12420 11780
rect 12580 11620 12700 11780
rect 12300 11500 12700 11620
rect 13100 11780 13500 11900
rect 13100 11620 13220 11780
rect 13380 11620 13500 11780
rect 13100 11500 13500 11620
rect 13900 11780 14300 11900
rect 13900 11620 14020 11780
rect 14180 11620 14300 11780
rect 13900 11500 14300 11620
rect 14700 11780 15100 11900
rect 14700 11620 14820 11780
rect 14980 11620 15100 11780
rect 14700 11500 15100 11620
rect 15500 11780 15900 11900
rect 15500 11620 15620 11780
rect 15780 11620 15900 11780
rect 15500 11500 15900 11620
rect 700 11380 1100 11500
rect 700 11220 820 11380
rect 980 11220 1100 11380
rect 700 11100 1100 11220
rect 1500 11380 1900 11500
rect 1500 11220 1620 11380
rect 1780 11220 1900 11380
rect 1500 11100 1900 11220
rect 2300 11380 2700 11500
rect 2300 11220 2420 11380
rect 2580 11220 2700 11380
rect 2300 11100 2700 11220
rect 3100 11380 3500 11500
rect 3100 11220 3220 11380
rect 3380 11220 3500 11380
rect 3100 11100 3500 11220
rect 3900 11380 4300 11500
rect 3900 11220 4020 11380
rect 4180 11220 4300 11380
rect 3900 11100 4300 11220
rect 4700 11380 5100 11500
rect 4700 11220 4820 11380
rect 4980 11220 5100 11380
rect 4700 11100 5100 11220
rect 5500 11380 5900 11500
rect 5500 11220 5620 11380
rect 5780 11220 5900 11380
rect 5500 11100 5900 11220
rect 6300 11380 6700 11500
rect 6300 11220 6420 11380
rect 6580 11220 6700 11380
rect 6300 11100 6700 11220
rect 7100 11380 7500 11500
rect 7100 11220 7220 11380
rect 7380 11220 7500 11380
rect 7100 11100 7500 11220
rect 7900 11380 8300 11500
rect 7900 11220 8020 11380
rect 8180 11220 8300 11380
rect 7900 11100 8300 11220
rect 8700 11380 9100 11500
rect 8700 11220 8820 11380
rect 8980 11220 9100 11380
rect 8700 11100 9100 11220
rect 9500 11380 9900 11500
rect 9500 11220 9620 11380
rect 9780 11220 9900 11380
rect 9500 11100 9900 11220
rect 10300 11380 10700 11500
rect 10300 11220 10420 11380
rect 10580 11220 10700 11380
rect 10300 11100 10700 11220
rect 11100 11380 11500 11500
rect 11100 11220 11220 11380
rect 11380 11220 11500 11380
rect 11100 11100 11500 11220
rect 11900 11380 12300 11500
rect 11900 11220 12020 11380
rect 12180 11220 12300 11380
rect 11900 11100 12300 11220
rect 12700 11380 13100 11500
rect 12700 11220 12820 11380
rect 12980 11220 13100 11380
rect 12700 11100 13100 11220
rect 13500 11380 13900 11500
rect 13500 11220 13620 11380
rect 13780 11220 13900 11380
rect 13500 11100 13900 11220
rect 14300 11380 14700 11500
rect 14300 11220 14420 11380
rect 14580 11220 14700 11380
rect 14300 11100 14700 11220
rect 15100 11380 15500 11500
rect 15100 11220 15220 11380
rect 15380 11220 15500 11380
rect 15100 11100 15500 11220
rect 15900 11380 16300 11500
rect 15900 11220 16020 11380
rect 16180 11220 16300 11380
rect 15900 11100 16300 11220
rect 1100 10980 1500 11100
rect 1100 10820 1220 10980
rect 1380 10820 1500 10980
rect 1100 10700 1500 10820
rect 1900 10980 2300 11100
rect 1900 10820 2020 10980
rect 2180 10820 2300 10980
rect 1900 10700 2300 10820
rect 2700 10980 3100 11100
rect 2700 10820 2820 10980
rect 2980 10820 3100 10980
rect 2700 10700 3100 10820
rect 3500 10980 3900 11100
rect 3500 10820 3620 10980
rect 3780 10820 3900 10980
rect 3500 10700 3900 10820
rect 4300 10980 4700 11100
rect 4300 10820 4420 10980
rect 4580 10820 4700 10980
rect 4300 10700 4700 10820
rect 5100 10980 5500 11100
rect 5100 10820 5220 10980
rect 5380 10820 5500 10980
rect 5100 10700 5500 10820
rect 5900 10980 6300 11100
rect 5900 10820 6020 10980
rect 6180 10820 6300 10980
rect 5900 10700 6300 10820
rect 6700 10980 7100 11100
rect 6700 10820 6820 10980
rect 6980 10820 7100 10980
rect 6700 10700 7100 10820
rect 7500 10980 7900 11100
rect 7500 10820 7620 10980
rect 7780 10820 7900 10980
rect 7500 10700 7900 10820
rect 8300 10980 8700 11100
rect 8300 10820 8420 10980
rect 8580 10820 8700 10980
rect 8300 10700 8700 10820
rect 9100 10980 9500 11100
rect 9100 10820 9220 10980
rect 9380 10820 9500 10980
rect 9100 10700 9500 10820
rect 9900 10980 10300 11100
rect 9900 10820 10020 10980
rect 10180 10820 10300 10980
rect 9900 10700 10300 10820
rect 10700 10980 11100 11100
rect 10700 10820 10820 10980
rect 10980 10820 11100 10980
rect 10700 10700 11100 10820
rect 11500 10980 11900 11100
rect 11500 10820 11620 10980
rect 11780 10820 11900 10980
rect 11500 10700 11900 10820
rect 12300 10980 12700 11100
rect 12300 10820 12420 10980
rect 12580 10820 12700 10980
rect 12300 10700 12700 10820
rect 13100 10980 13500 11100
rect 13100 10820 13220 10980
rect 13380 10820 13500 10980
rect 13100 10700 13500 10820
rect 13900 10980 14300 11100
rect 13900 10820 14020 10980
rect 14180 10820 14300 10980
rect 13900 10700 14300 10820
rect 14700 10980 15100 11100
rect 14700 10820 14820 10980
rect 14980 10820 15100 10980
rect 14700 10700 15100 10820
rect 15500 10980 15900 11100
rect 15500 10820 15620 10980
rect 15780 10820 15900 10980
rect 15500 10700 15900 10820
rect 700 10580 1100 10700
rect 700 10420 820 10580
rect 980 10420 1100 10580
rect 700 10300 1100 10420
rect 1500 10580 1900 10700
rect 1500 10420 1620 10580
rect 1780 10420 1900 10580
rect 1500 10300 1900 10420
rect 2300 10580 2700 10700
rect 2300 10420 2420 10580
rect 2580 10420 2700 10580
rect 2300 10300 2700 10420
rect 3100 10580 3500 10700
rect 3100 10420 3220 10580
rect 3380 10420 3500 10580
rect 3100 10300 3500 10420
rect 3900 10580 4300 10700
rect 3900 10420 4020 10580
rect 4180 10420 4300 10580
rect 3900 10300 4300 10420
rect 4700 10580 5100 10700
rect 4700 10420 4820 10580
rect 4980 10420 5100 10580
rect 4700 10300 5100 10420
rect 5500 10580 5900 10700
rect 5500 10420 5620 10580
rect 5780 10420 5900 10580
rect 5500 10300 5900 10420
rect 6300 10580 6700 10700
rect 6300 10420 6420 10580
rect 6580 10420 6700 10580
rect 6300 10300 6700 10420
rect 7100 10580 7500 10700
rect 7100 10420 7220 10580
rect 7380 10420 7500 10580
rect 7100 10300 7500 10420
rect 7900 10580 8300 10700
rect 7900 10420 8020 10580
rect 8180 10420 8300 10580
rect 7900 10300 8300 10420
rect 8700 10580 9100 10700
rect 8700 10420 8820 10580
rect 8980 10420 9100 10580
rect 8700 10300 9100 10420
rect 9500 10580 9900 10700
rect 9500 10420 9620 10580
rect 9780 10420 9900 10580
rect 9500 10300 9900 10420
rect 10300 10580 10700 10700
rect 10300 10420 10420 10580
rect 10580 10420 10700 10580
rect 10300 10300 10700 10420
rect 11100 10580 11500 10700
rect 11100 10420 11220 10580
rect 11380 10420 11500 10580
rect 11100 10300 11500 10420
rect 11900 10580 12300 10700
rect 11900 10420 12020 10580
rect 12180 10420 12300 10580
rect 11900 10300 12300 10420
rect 12700 10580 13100 10700
rect 12700 10420 12820 10580
rect 12980 10420 13100 10580
rect 12700 10300 13100 10420
rect 13500 10580 13900 10700
rect 13500 10420 13620 10580
rect 13780 10420 13900 10580
rect 13500 10300 13900 10420
rect 14300 10580 14700 10700
rect 14300 10420 14420 10580
rect 14580 10420 14700 10580
rect 14300 10300 14700 10420
rect 15100 10580 15500 10700
rect 15100 10420 15220 10580
rect 15380 10420 15500 10580
rect 15100 10300 15500 10420
rect 15900 10580 16300 10700
rect 15900 10420 16020 10580
rect 16180 10420 16300 10580
rect 15900 10300 16300 10420
rect 1100 10180 1500 10300
rect 1100 10020 1220 10180
rect 1380 10020 1500 10180
rect 1100 9900 1500 10020
rect 1900 10180 2300 10300
rect 1900 10020 2020 10180
rect 2180 10020 2300 10180
rect 1900 9900 2300 10020
rect 2700 10180 3100 10300
rect 2700 10020 2820 10180
rect 2980 10020 3100 10180
rect 2700 9900 3100 10020
rect 3500 10180 3900 10300
rect 3500 10020 3620 10180
rect 3780 10020 3900 10180
rect 3500 9900 3900 10020
rect 4300 10180 4700 10300
rect 4300 10020 4420 10180
rect 4580 10020 4700 10180
rect 4300 9900 4700 10020
rect 5100 10180 5500 10300
rect 5100 10020 5220 10180
rect 5380 10020 5500 10180
rect 5100 9900 5500 10020
rect 5900 10180 6300 10300
rect 5900 10020 6020 10180
rect 6180 10020 6300 10180
rect 5900 9900 6300 10020
rect 6700 10180 7100 10300
rect 6700 10020 6820 10180
rect 6980 10020 7100 10180
rect 6700 9900 7100 10020
rect 7500 10180 7900 10300
rect 7500 10020 7620 10180
rect 7780 10020 7900 10180
rect 7500 9900 7900 10020
rect 8300 10180 8700 10300
rect 8300 10020 8420 10180
rect 8580 10020 8700 10180
rect 8300 9900 8700 10020
rect 9100 10180 9500 10300
rect 9100 10020 9220 10180
rect 9380 10020 9500 10180
rect 9100 9900 9500 10020
rect 9900 10180 10300 10300
rect 9900 10020 10020 10180
rect 10180 10020 10300 10180
rect 9900 9900 10300 10020
rect 10700 10180 11100 10300
rect 10700 10020 10820 10180
rect 10980 10020 11100 10180
rect 10700 9900 11100 10020
rect 11500 10180 11900 10300
rect 11500 10020 11620 10180
rect 11780 10020 11900 10180
rect 11500 9900 11900 10020
rect 12300 10180 12700 10300
rect 12300 10020 12420 10180
rect 12580 10020 12700 10180
rect 12300 9900 12700 10020
rect 13100 10180 13500 10300
rect 13100 10020 13220 10180
rect 13380 10020 13500 10180
rect 13100 9900 13500 10020
rect 13900 10180 14300 10300
rect 13900 10020 14020 10180
rect 14180 10020 14300 10180
rect 13900 9900 14300 10020
rect 14700 10180 15100 10300
rect 14700 10020 14820 10180
rect 14980 10020 15100 10180
rect 14700 9900 15100 10020
rect 15500 10180 15900 10300
rect 15500 10020 15620 10180
rect 15780 10020 15900 10180
rect 15500 9900 15900 10020
rect 700 9780 1100 9900
rect 700 9620 820 9780
rect 980 9620 1100 9780
rect 700 9500 1100 9620
rect 1500 9780 1900 9900
rect 1500 9620 1620 9780
rect 1780 9620 1900 9780
rect 1500 9500 1900 9620
rect 2300 9780 2700 9900
rect 2300 9620 2420 9780
rect 2580 9620 2700 9780
rect 2300 9500 2700 9620
rect 3100 9780 3500 9900
rect 3100 9620 3220 9780
rect 3380 9620 3500 9780
rect 3100 9500 3500 9620
rect 3900 9780 4300 9900
rect 3900 9620 4020 9780
rect 4180 9620 4300 9780
rect 3900 9500 4300 9620
rect 4700 9780 5100 9900
rect 4700 9620 4820 9780
rect 4980 9620 5100 9780
rect 4700 9500 5100 9620
rect 5500 9780 5900 9900
rect 5500 9620 5620 9780
rect 5780 9620 5900 9780
rect 5500 9500 5900 9620
rect 6300 9780 6700 9900
rect 6300 9620 6420 9780
rect 6580 9620 6700 9780
rect 6300 9500 6700 9620
rect 7100 9780 7500 9900
rect 7100 9620 7220 9780
rect 7380 9620 7500 9780
rect 7100 9500 7500 9620
rect 7900 9780 8300 9900
rect 7900 9620 8020 9780
rect 8180 9620 8300 9780
rect 7900 9500 8300 9620
rect 8700 9780 9100 9900
rect 8700 9620 8820 9780
rect 8980 9620 9100 9780
rect 8700 9500 9100 9620
rect 9500 9780 9900 9900
rect 9500 9620 9620 9780
rect 9780 9620 9900 9780
rect 9500 9500 9900 9620
rect 10300 9780 10700 9900
rect 10300 9620 10420 9780
rect 10580 9620 10700 9780
rect 10300 9500 10700 9620
rect 11100 9780 11500 9900
rect 11100 9620 11220 9780
rect 11380 9620 11500 9780
rect 11100 9500 11500 9620
rect 11900 9780 12300 9900
rect 11900 9620 12020 9780
rect 12180 9620 12300 9780
rect 11900 9500 12300 9620
rect 12700 9780 13100 9900
rect 12700 9620 12820 9780
rect 12980 9620 13100 9780
rect 12700 9500 13100 9620
rect 13500 9780 13900 9900
rect 13500 9620 13620 9780
rect 13780 9620 13900 9780
rect 13500 9500 13900 9620
rect 14300 9780 14700 9900
rect 14300 9620 14420 9780
rect 14580 9620 14700 9780
rect 14300 9500 14700 9620
rect 15100 9780 15500 9900
rect 15100 9620 15220 9780
rect 15380 9620 15500 9780
rect 15100 9500 15500 9620
rect 15900 9780 16300 9900
rect 15900 9620 16020 9780
rect 16180 9620 16300 9780
rect 15900 9500 16300 9620
rect 1100 9380 1500 9500
rect 1100 9220 1220 9380
rect 1380 9220 1500 9380
rect 1100 9100 1500 9220
rect 1900 9380 2300 9500
rect 1900 9220 2020 9380
rect 2180 9220 2300 9380
rect 1900 9100 2300 9220
rect 2700 9380 3100 9500
rect 2700 9220 2820 9380
rect 2980 9220 3100 9380
rect 2700 9100 3100 9220
rect 3500 9380 3900 9500
rect 3500 9220 3620 9380
rect 3780 9220 3900 9380
rect 3500 9100 3900 9220
rect 4300 9380 4700 9500
rect 4300 9220 4420 9380
rect 4580 9220 4700 9380
rect 4300 9100 4700 9220
rect 5100 9380 5500 9500
rect 5100 9220 5220 9380
rect 5380 9220 5500 9380
rect 5100 9100 5500 9220
rect 5900 9380 6300 9500
rect 5900 9220 6020 9380
rect 6180 9220 6300 9380
rect 5900 9100 6300 9220
rect 6700 9380 7100 9500
rect 6700 9220 6820 9380
rect 6980 9220 7100 9380
rect 6700 9100 7100 9220
rect 7500 9380 7900 9500
rect 7500 9220 7620 9380
rect 7780 9220 7900 9380
rect 7500 9100 7900 9220
rect 8300 9380 8700 9500
rect 8300 9220 8420 9380
rect 8580 9220 8700 9380
rect 8300 9100 8700 9220
rect 9100 9380 9500 9500
rect 9100 9220 9220 9380
rect 9380 9220 9500 9380
rect 9100 9100 9500 9220
rect 9900 9380 10300 9500
rect 9900 9220 10020 9380
rect 10180 9220 10300 9380
rect 9900 9100 10300 9220
rect 10700 9380 11100 9500
rect 10700 9220 10820 9380
rect 10980 9220 11100 9380
rect 10700 9100 11100 9220
rect 11500 9380 11900 9500
rect 11500 9220 11620 9380
rect 11780 9220 11900 9380
rect 11500 9100 11900 9220
rect 12300 9380 12700 9500
rect 12300 9220 12420 9380
rect 12580 9220 12700 9380
rect 12300 9100 12700 9220
rect 13100 9380 13500 9500
rect 13100 9220 13220 9380
rect 13380 9220 13500 9380
rect 13100 9100 13500 9220
rect 13900 9380 14300 9500
rect 13900 9220 14020 9380
rect 14180 9220 14300 9380
rect 13900 9100 14300 9220
rect 14700 9380 15100 9500
rect 14700 9220 14820 9380
rect 14980 9220 15100 9380
rect 14700 9100 15100 9220
rect 15500 9380 15900 9500
rect 15500 9220 15620 9380
rect 15780 9220 15900 9380
rect 15500 9100 15900 9220
rect 700 8980 1100 9100
rect 700 8820 820 8980
rect 980 8820 1100 8980
rect 700 8700 1100 8820
rect 1500 8980 1900 9100
rect 1500 8820 1620 8980
rect 1780 8820 1900 8980
rect 1500 8700 1900 8820
rect 2300 8980 2700 9100
rect 2300 8820 2420 8980
rect 2580 8820 2700 8980
rect 2300 8700 2700 8820
rect 3100 8980 3500 9100
rect 3100 8820 3220 8980
rect 3380 8820 3500 8980
rect 3100 8700 3500 8820
rect 3900 8980 4300 9100
rect 3900 8820 4020 8980
rect 4180 8820 4300 8980
rect 3900 8700 4300 8820
rect 4700 8980 5100 9100
rect 4700 8820 4820 8980
rect 4980 8820 5100 8980
rect 4700 8700 5100 8820
rect 5500 8980 5900 9100
rect 5500 8820 5620 8980
rect 5780 8820 5900 8980
rect 5500 8700 5900 8820
rect 6300 8980 6700 9100
rect 6300 8820 6420 8980
rect 6580 8820 6700 8980
rect 6300 8700 6700 8820
rect 7100 8980 7500 9100
rect 7100 8820 7220 8980
rect 7380 8820 7500 8980
rect 7100 8700 7500 8820
rect 7900 8980 8300 9100
rect 7900 8820 8020 8980
rect 8180 8820 8300 8980
rect 7900 8700 8300 8820
rect 8700 8980 9100 9100
rect 8700 8820 8820 8980
rect 8980 8820 9100 8980
rect 8700 8700 9100 8820
rect 9500 8980 9900 9100
rect 9500 8820 9620 8980
rect 9780 8820 9900 8980
rect 9500 8700 9900 8820
rect 10300 8980 10700 9100
rect 10300 8820 10420 8980
rect 10580 8820 10700 8980
rect 10300 8700 10700 8820
rect 11100 8980 11500 9100
rect 11100 8820 11220 8980
rect 11380 8820 11500 8980
rect 11100 8700 11500 8820
rect 11900 8980 12300 9100
rect 11900 8820 12020 8980
rect 12180 8820 12300 8980
rect 11900 8700 12300 8820
rect 12700 8980 13100 9100
rect 12700 8820 12820 8980
rect 12980 8820 13100 8980
rect 12700 8700 13100 8820
rect 13500 8980 13900 9100
rect 13500 8820 13620 8980
rect 13780 8820 13900 8980
rect 13500 8700 13900 8820
rect 14300 8980 14700 9100
rect 14300 8820 14420 8980
rect 14580 8820 14700 8980
rect 14300 8700 14700 8820
rect 15100 8980 15500 9100
rect 15100 8820 15220 8980
rect 15380 8820 15500 8980
rect 15100 8700 15500 8820
rect 15900 8980 16300 9100
rect 15900 8820 16020 8980
rect 16180 8820 16300 8980
rect 15900 8700 16300 8820
rect 1100 8580 1500 8700
rect 1100 8420 1220 8580
rect 1380 8420 1500 8580
rect 1100 8300 1500 8420
rect 1900 8580 2300 8700
rect 1900 8420 2020 8580
rect 2180 8420 2300 8580
rect 1900 8300 2300 8420
rect 2700 8580 3100 8700
rect 2700 8420 2820 8580
rect 2980 8420 3100 8580
rect 2700 8300 3100 8420
rect 3500 8580 3900 8700
rect 3500 8420 3620 8580
rect 3780 8420 3900 8580
rect 3500 8300 3900 8420
rect 4300 8580 4700 8700
rect 4300 8420 4420 8580
rect 4580 8420 4700 8580
rect 4300 8300 4700 8420
rect 5100 8580 5500 8700
rect 5100 8420 5220 8580
rect 5380 8420 5500 8580
rect 5100 8300 5500 8420
rect 5900 8580 6300 8700
rect 5900 8420 6020 8580
rect 6180 8420 6300 8580
rect 5900 8300 6300 8420
rect 6700 8580 7100 8700
rect 6700 8420 6820 8580
rect 6980 8420 7100 8580
rect 6700 8300 7100 8420
rect 7500 8580 7900 8700
rect 7500 8420 7620 8580
rect 7780 8420 7900 8580
rect 7500 8300 7900 8420
rect 8300 8580 8700 8700
rect 8300 8420 8420 8580
rect 8580 8420 8700 8580
rect 8300 8300 8700 8420
rect 9100 8580 9500 8700
rect 9100 8420 9220 8580
rect 9380 8420 9500 8580
rect 9100 8300 9500 8420
rect 9900 8580 10300 8700
rect 9900 8420 10020 8580
rect 10180 8420 10300 8580
rect 9900 8300 10300 8420
rect 10700 8580 11100 8700
rect 10700 8420 10820 8580
rect 10980 8420 11100 8580
rect 10700 8300 11100 8420
rect 11500 8580 11900 8700
rect 11500 8420 11620 8580
rect 11780 8420 11900 8580
rect 11500 8300 11900 8420
rect 12300 8580 12700 8700
rect 12300 8420 12420 8580
rect 12580 8420 12700 8580
rect 12300 8300 12700 8420
rect 13100 8580 13500 8700
rect 13100 8420 13220 8580
rect 13380 8420 13500 8580
rect 13100 8300 13500 8420
rect 13900 8580 14300 8700
rect 13900 8420 14020 8580
rect 14180 8420 14300 8580
rect 13900 8300 14300 8420
rect 14700 8580 15100 8700
rect 14700 8420 14820 8580
rect 14980 8420 15100 8580
rect 14700 8300 15100 8420
rect 15500 8580 15900 8700
rect 15500 8420 15620 8580
rect 15780 8420 15900 8580
rect 15500 8300 15900 8420
rect 700 8180 1100 8300
rect 700 8020 820 8180
rect 980 8020 1100 8180
rect 700 7900 1100 8020
rect 1500 8180 1900 8300
rect 1500 8020 1620 8180
rect 1780 8020 1900 8180
rect 1500 7900 1900 8020
rect 2300 8180 2700 8300
rect 2300 8020 2420 8180
rect 2580 8020 2700 8180
rect 2300 7900 2700 8020
rect 3100 8180 3500 8300
rect 3100 8020 3220 8180
rect 3380 8020 3500 8180
rect 3100 7900 3500 8020
rect 3900 8180 4300 8300
rect 3900 8020 4020 8180
rect 4180 8020 4300 8180
rect 3900 7900 4300 8020
rect 4700 8180 5100 8300
rect 4700 8020 4820 8180
rect 4980 8020 5100 8180
rect 4700 7900 5100 8020
rect 5500 8180 5900 8300
rect 5500 8020 5620 8180
rect 5780 8020 5900 8180
rect 5500 7900 5900 8020
rect 6300 8180 6700 8300
rect 6300 8020 6420 8180
rect 6580 8020 6700 8180
rect 6300 7900 6700 8020
rect 7100 8180 7500 8300
rect 7100 8020 7220 8180
rect 7380 8020 7500 8180
rect 7100 7900 7500 8020
rect 7900 8180 8300 8300
rect 7900 8020 8020 8180
rect 8180 8020 8300 8180
rect 7900 7900 8300 8020
rect 8700 8180 9100 8300
rect 8700 8020 8820 8180
rect 8980 8020 9100 8180
rect 8700 7900 9100 8020
rect 9500 8180 9900 8300
rect 9500 8020 9620 8180
rect 9780 8020 9900 8180
rect 9500 7900 9900 8020
rect 10300 8180 10700 8300
rect 10300 8020 10420 8180
rect 10580 8020 10700 8180
rect 10300 7900 10700 8020
rect 11100 8180 11500 8300
rect 11100 8020 11220 8180
rect 11380 8020 11500 8180
rect 11100 7900 11500 8020
rect 11900 8180 12300 8300
rect 11900 8020 12020 8180
rect 12180 8020 12300 8180
rect 11900 7900 12300 8020
rect 12700 8180 13100 8300
rect 12700 8020 12820 8180
rect 12980 8020 13100 8180
rect 12700 7900 13100 8020
rect 13500 8180 13900 8300
rect 13500 8020 13620 8180
rect 13780 8020 13900 8180
rect 13500 7900 13900 8020
rect 14300 8180 14700 8300
rect 14300 8020 14420 8180
rect 14580 8020 14700 8180
rect 14300 7900 14700 8020
rect 15100 8180 15500 8300
rect 15100 8020 15220 8180
rect 15380 8020 15500 8180
rect 15100 7900 15500 8020
rect 15900 8180 16300 8300
rect 15900 8020 16020 8180
rect 16180 8020 16300 8180
rect 15900 7900 16300 8020
rect 1100 7780 1500 7900
rect 1100 7620 1220 7780
rect 1380 7620 1500 7780
rect 1100 7500 1500 7620
rect 1900 7780 2300 7900
rect 1900 7620 2020 7780
rect 2180 7620 2300 7780
rect 1900 7500 2300 7620
rect 2700 7780 3100 7900
rect 2700 7620 2820 7780
rect 2980 7620 3100 7780
rect 2700 7500 3100 7620
rect 3500 7780 3900 7900
rect 3500 7620 3620 7780
rect 3780 7620 3900 7780
rect 3500 7500 3900 7620
rect 4300 7780 4700 7900
rect 4300 7620 4420 7780
rect 4580 7620 4700 7780
rect 4300 7500 4700 7620
rect 5100 7780 5500 7900
rect 5100 7620 5220 7780
rect 5380 7620 5500 7780
rect 5100 7500 5500 7620
rect 5900 7780 6300 7900
rect 5900 7620 6020 7780
rect 6180 7620 6300 7780
rect 5900 7500 6300 7620
rect 6700 7780 7100 7900
rect 6700 7620 6820 7780
rect 6980 7620 7100 7780
rect 6700 7500 7100 7620
rect 7500 7780 7900 7900
rect 7500 7620 7620 7780
rect 7780 7620 7900 7780
rect 7500 7500 7900 7620
rect 8300 7780 8700 7900
rect 8300 7620 8420 7780
rect 8580 7620 8700 7780
rect 8300 7500 8700 7620
rect 9100 7780 9500 7900
rect 9100 7620 9220 7780
rect 9380 7620 9500 7780
rect 9100 7500 9500 7620
rect 9900 7780 10300 7900
rect 9900 7620 10020 7780
rect 10180 7620 10300 7780
rect 9900 7500 10300 7620
rect 10700 7780 11100 7900
rect 10700 7620 10820 7780
rect 10980 7620 11100 7780
rect 10700 7500 11100 7620
rect 11500 7780 11900 7900
rect 11500 7620 11620 7780
rect 11780 7620 11900 7780
rect 11500 7500 11900 7620
rect 12300 7780 12700 7900
rect 12300 7620 12420 7780
rect 12580 7620 12700 7780
rect 12300 7500 12700 7620
rect 13100 7780 13500 7900
rect 13100 7620 13220 7780
rect 13380 7620 13500 7780
rect 13100 7500 13500 7620
rect 13900 7780 14300 7900
rect 13900 7620 14020 7780
rect 14180 7620 14300 7780
rect 13900 7500 14300 7620
rect 14700 7780 15100 7900
rect 14700 7620 14820 7780
rect 14980 7620 15100 7780
rect 14700 7500 15100 7620
rect 15500 7780 15900 7900
rect 15500 7620 15620 7780
rect 15780 7620 15900 7780
rect 15500 7500 15900 7620
rect 700 7380 1100 7500
rect 700 7220 820 7380
rect 980 7220 1100 7380
rect 700 7100 1100 7220
rect 1500 7380 1900 7500
rect 1500 7220 1620 7380
rect 1780 7220 1900 7380
rect 1500 7100 1900 7220
rect 2300 7380 2700 7500
rect 2300 7220 2420 7380
rect 2580 7220 2700 7380
rect 2300 7100 2700 7220
rect 3100 7380 3500 7500
rect 3100 7220 3220 7380
rect 3380 7220 3500 7380
rect 3100 7100 3500 7220
rect 3900 7380 4300 7500
rect 3900 7220 4020 7380
rect 4180 7220 4300 7380
rect 3900 7100 4300 7220
rect 4700 7380 5100 7500
rect 4700 7220 4820 7380
rect 4980 7220 5100 7380
rect 4700 7100 5100 7220
rect 5500 7380 5900 7500
rect 5500 7220 5620 7380
rect 5780 7220 5900 7380
rect 5500 7100 5900 7220
rect 6300 7380 6700 7500
rect 6300 7220 6420 7380
rect 6580 7220 6700 7380
rect 6300 7100 6700 7220
rect 7100 7380 7500 7500
rect 7100 7220 7220 7380
rect 7380 7220 7500 7380
rect 7100 7100 7500 7220
rect 7900 7380 8300 7500
rect 7900 7220 8020 7380
rect 8180 7220 8300 7380
rect 7900 7100 8300 7220
rect 8700 7380 9100 7500
rect 8700 7220 8820 7380
rect 8980 7220 9100 7380
rect 8700 7100 9100 7220
rect 9500 7380 9900 7500
rect 9500 7220 9620 7380
rect 9780 7220 9900 7380
rect 9500 7100 9900 7220
rect 10300 7380 10700 7500
rect 10300 7220 10420 7380
rect 10580 7220 10700 7380
rect 10300 7100 10700 7220
rect 11100 7380 11500 7500
rect 11100 7220 11220 7380
rect 11380 7220 11500 7380
rect 11100 7100 11500 7220
rect 11900 7380 12300 7500
rect 11900 7220 12020 7380
rect 12180 7220 12300 7380
rect 11900 7100 12300 7220
rect 12700 7380 13100 7500
rect 12700 7220 12820 7380
rect 12980 7220 13100 7380
rect 12700 7100 13100 7220
rect 13500 7380 13900 7500
rect 13500 7220 13620 7380
rect 13780 7220 13900 7380
rect 13500 7100 13900 7220
rect 14300 7380 14700 7500
rect 14300 7220 14420 7380
rect 14580 7220 14700 7380
rect 14300 7100 14700 7220
rect 15100 7380 15500 7500
rect 15100 7220 15220 7380
rect 15380 7220 15500 7380
rect 15100 7100 15500 7220
rect 15900 7380 16300 7500
rect 15900 7220 16020 7380
rect 16180 7220 16300 7380
rect 15900 7100 16300 7220
rect 1100 6980 1500 7100
rect 1100 6820 1220 6980
rect 1380 6820 1500 6980
rect 1100 6700 1500 6820
rect 1900 6980 2300 7100
rect 1900 6820 2020 6980
rect 2180 6820 2300 6980
rect 1900 6700 2300 6820
rect 2700 6980 3100 7100
rect 2700 6820 2820 6980
rect 2980 6820 3100 6980
rect 2700 6700 3100 6820
rect 3500 6980 3900 7100
rect 3500 6820 3620 6980
rect 3780 6820 3900 6980
rect 3500 6700 3900 6820
rect 4300 6980 4700 7100
rect 4300 6820 4420 6980
rect 4580 6820 4700 6980
rect 4300 6700 4700 6820
rect 5100 6980 5500 7100
rect 5100 6820 5220 6980
rect 5380 6820 5500 6980
rect 5100 6700 5500 6820
rect 5900 6980 6300 7100
rect 5900 6820 6020 6980
rect 6180 6820 6300 6980
rect 5900 6700 6300 6820
rect 6700 6980 7100 7100
rect 6700 6820 6820 6980
rect 6980 6820 7100 6980
rect 6700 6700 7100 6820
rect 7500 6980 7900 7100
rect 7500 6820 7620 6980
rect 7780 6820 7900 6980
rect 7500 6700 7900 6820
rect 8300 6980 8700 7100
rect 8300 6820 8420 6980
rect 8580 6820 8700 6980
rect 8300 6700 8700 6820
rect 9100 6980 9500 7100
rect 9100 6820 9220 6980
rect 9380 6820 9500 6980
rect 9100 6700 9500 6820
rect 9900 6980 10300 7100
rect 9900 6820 10020 6980
rect 10180 6820 10300 6980
rect 9900 6700 10300 6820
rect 10700 6980 11100 7100
rect 10700 6820 10820 6980
rect 10980 6820 11100 6980
rect 10700 6700 11100 6820
rect 11500 6980 11900 7100
rect 11500 6820 11620 6980
rect 11780 6820 11900 6980
rect 11500 6700 11900 6820
rect 12300 6980 12700 7100
rect 12300 6820 12420 6980
rect 12580 6820 12700 6980
rect 12300 6700 12700 6820
rect 13100 6980 13500 7100
rect 13100 6820 13220 6980
rect 13380 6820 13500 6980
rect 13100 6700 13500 6820
rect 13900 6980 14300 7100
rect 13900 6820 14020 6980
rect 14180 6820 14300 6980
rect 13900 6700 14300 6820
rect 14700 6980 15100 7100
rect 14700 6820 14820 6980
rect 14980 6820 15100 6980
rect 14700 6700 15100 6820
rect 15500 6980 15900 7100
rect 15500 6820 15620 6980
rect 15780 6820 15900 6980
rect 15500 6700 15900 6820
rect 700 6580 1100 6700
rect 700 6420 820 6580
rect 980 6420 1100 6580
rect 700 6300 1100 6420
rect 1500 6580 1900 6700
rect 1500 6420 1620 6580
rect 1780 6420 1900 6580
rect 1500 6300 1900 6420
rect 2300 6580 2700 6700
rect 2300 6420 2420 6580
rect 2580 6420 2700 6580
rect 2300 6300 2700 6420
rect 3100 6580 3500 6700
rect 3100 6420 3220 6580
rect 3380 6420 3500 6580
rect 3100 6300 3500 6420
rect 3900 6580 4300 6700
rect 3900 6420 4020 6580
rect 4180 6420 4300 6580
rect 3900 6300 4300 6420
rect 4700 6580 5100 6700
rect 4700 6420 4820 6580
rect 4980 6420 5100 6580
rect 4700 6300 5100 6420
rect 5500 6580 5900 6700
rect 5500 6420 5620 6580
rect 5780 6420 5900 6580
rect 5500 6300 5900 6420
rect 6300 6580 6700 6700
rect 6300 6420 6420 6580
rect 6580 6420 6700 6580
rect 6300 6300 6700 6420
rect 7100 6580 7500 6700
rect 7100 6420 7220 6580
rect 7380 6420 7500 6580
rect 7100 6300 7500 6420
rect 7900 6580 8300 6700
rect 7900 6420 8020 6580
rect 8180 6420 8300 6580
rect 7900 6300 8300 6420
rect 8700 6580 9100 6700
rect 8700 6420 8820 6580
rect 8980 6420 9100 6580
rect 8700 6300 9100 6420
rect 9500 6580 9900 6700
rect 9500 6420 9620 6580
rect 9780 6420 9900 6580
rect 9500 6300 9900 6420
rect 10300 6580 10700 6700
rect 10300 6420 10420 6580
rect 10580 6420 10700 6580
rect 10300 6300 10700 6420
rect 11100 6580 11500 6700
rect 11100 6420 11220 6580
rect 11380 6420 11500 6580
rect 11100 6300 11500 6420
rect 11900 6580 12300 6700
rect 11900 6420 12020 6580
rect 12180 6420 12300 6580
rect 11900 6300 12300 6420
rect 12700 6580 13100 6700
rect 12700 6420 12820 6580
rect 12980 6420 13100 6580
rect 12700 6300 13100 6420
rect 13500 6580 13900 6700
rect 13500 6420 13620 6580
rect 13780 6420 13900 6580
rect 13500 6300 13900 6420
rect 14300 6580 14700 6700
rect 14300 6420 14420 6580
rect 14580 6420 14700 6580
rect 14300 6300 14700 6420
rect 15100 6580 15500 6700
rect 15100 6420 15220 6580
rect 15380 6420 15500 6580
rect 15100 6300 15500 6420
rect 15900 6580 16300 6700
rect 15900 6420 16020 6580
rect 16180 6420 16300 6580
rect 15900 6300 16300 6420
rect 1100 6180 1500 6300
rect 1100 6020 1220 6180
rect 1380 6020 1500 6180
rect 1100 5900 1500 6020
rect 1900 6180 2300 6300
rect 1900 6020 2020 6180
rect 2180 6020 2300 6180
rect 1900 5900 2300 6020
rect 2700 6180 3100 6300
rect 2700 6020 2820 6180
rect 2980 6020 3100 6180
rect 2700 5900 3100 6020
rect 3500 6180 3900 6300
rect 3500 6020 3620 6180
rect 3780 6020 3900 6180
rect 3500 5900 3900 6020
rect 4300 6180 4700 6300
rect 4300 6020 4420 6180
rect 4580 6020 4700 6180
rect 4300 5900 4700 6020
rect 5100 6180 5500 6300
rect 5100 6020 5220 6180
rect 5380 6020 5500 6180
rect 5100 5900 5500 6020
rect 5900 6180 6300 6300
rect 5900 6020 6020 6180
rect 6180 6020 6300 6180
rect 5900 5900 6300 6020
rect 6700 6180 7100 6300
rect 6700 6020 6820 6180
rect 6980 6020 7100 6180
rect 6700 5900 7100 6020
rect 7500 6180 7900 6300
rect 7500 6020 7620 6180
rect 7780 6020 7900 6180
rect 7500 5900 7900 6020
rect 8300 6180 8700 6300
rect 8300 6020 8420 6180
rect 8580 6020 8700 6180
rect 8300 5900 8700 6020
rect 9100 6180 9500 6300
rect 9100 6020 9220 6180
rect 9380 6020 9500 6180
rect 9100 5900 9500 6020
rect 9900 6180 10300 6300
rect 9900 6020 10020 6180
rect 10180 6020 10300 6180
rect 9900 5900 10300 6020
rect 10700 6180 11100 6300
rect 10700 6020 10820 6180
rect 10980 6020 11100 6180
rect 10700 5900 11100 6020
rect 11500 6180 11900 6300
rect 11500 6020 11620 6180
rect 11780 6020 11900 6180
rect 11500 5900 11900 6020
rect 12300 6180 12700 6300
rect 12300 6020 12420 6180
rect 12580 6020 12700 6180
rect 12300 5900 12700 6020
rect 13100 6180 13500 6300
rect 13100 6020 13220 6180
rect 13380 6020 13500 6180
rect 13100 5900 13500 6020
rect 13900 6180 14300 6300
rect 13900 6020 14020 6180
rect 14180 6020 14300 6180
rect 13900 5900 14300 6020
rect 14700 6180 15100 6300
rect 14700 6020 14820 6180
rect 14980 6020 15100 6180
rect 14700 5900 15100 6020
rect 15500 6180 15900 6300
rect 15500 6020 15620 6180
rect 15780 6020 15900 6180
rect 15500 5900 15900 6020
rect 700 5780 1100 5900
rect 700 5620 820 5780
rect 980 5620 1100 5780
rect 700 5500 1100 5620
rect 1500 5780 1900 5900
rect 1500 5620 1620 5780
rect 1780 5620 1900 5780
rect 1500 5500 1900 5620
rect 2300 5780 2700 5900
rect 2300 5620 2420 5780
rect 2580 5620 2700 5780
rect 2300 5500 2700 5620
rect 3100 5780 3500 5900
rect 3100 5620 3220 5780
rect 3380 5620 3500 5780
rect 3100 5500 3500 5620
rect 3900 5780 4300 5900
rect 3900 5620 4020 5780
rect 4180 5620 4300 5780
rect 3900 5500 4300 5620
rect 4700 5780 5100 5900
rect 4700 5620 4820 5780
rect 4980 5620 5100 5780
rect 4700 5500 5100 5620
rect 5500 5780 5900 5900
rect 5500 5620 5620 5780
rect 5780 5620 5900 5780
rect 5500 5500 5900 5620
rect 6300 5780 6700 5900
rect 6300 5620 6420 5780
rect 6580 5620 6700 5780
rect 6300 5500 6700 5620
rect 7100 5780 7500 5900
rect 7100 5620 7220 5780
rect 7380 5620 7500 5780
rect 7100 5500 7500 5620
rect 7900 5780 8300 5900
rect 7900 5620 8020 5780
rect 8180 5620 8300 5780
rect 7900 5500 8300 5620
rect 8700 5780 9100 5900
rect 8700 5620 8820 5780
rect 8980 5620 9100 5780
rect 8700 5500 9100 5620
rect 9500 5780 9900 5900
rect 9500 5620 9620 5780
rect 9780 5620 9900 5780
rect 9500 5500 9900 5620
rect 10300 5780 10700 5900
rect 10300 5620 10420 5780
rect 10580 5620 10700 5780
rect 10300 5500 10700 5620
rect 11100 5780 11500 5900
rect 11100 5620 11220 5780
rect 11380 5620 11500 5780
rect 11100 5500 11500 5620
rect 11900 5780 12300 5900
rect 11900 5620 12020 5780
rect 12180 5620 12300 5780
rect 11900 5500 12300 5620
rect 12700 5780 13100 5900
rect 12700 5620 12820 5780
rect 12980 5620 13100 5780
rect 12700 5500 13100 5620
rect 13500 5780 13900 5900
rect 13500 5620 13620 5780
rect 13780 5620 13900 5780
rect 13500 5500 13900 5620
rect 14300 5780 14700 5900
rect 14300 5620 14420 5780
rect 14580 5620 14700 5780
rect 14300 5500 14700 5620
rect 15100 5780 15500 5900
rect 15100 5620 15220 5780
rect 15380 5620 15500 5780
rect 15100 5500 15500 5620
rect 15900 5780 16300 5900
rect 15900 5620 16020 5780
rect 16180 5620 16300 5780
rect 15900 5500 16300 5620
rect 1100 5380 1500 5500
rect 1100 5220 1220 5380
rect 1380 5220 1500 5380
rect 1100 5100 1500 5220
rect 1900 5380 2300 5500
rect 1900 5220 2020 5380
rect 2180 5220 2300 5380
rect 1900 5100 2300 5220
rect 2700 5380 3100 5500
rect 2700 5220 2820 5380
rect 2980 5220 3100 5380
rect 2700 5100 3100 5220
rect 3500 5380 3900 5500
rect 3500 5220 3620 5380
rect 3780 5220 3900 5380
rect 3500 5100 3900 5220
rect 4300 5380 4700 5500
rect 4300 5220 4420 5380
rect 4580 5220 4700 5380
rect 4300 5100 4700 5220
rect 5100 5380 5500 5500
rect 5100 5220 5220 5380
rect 5380 5220 5500 5380
rect 5100 5100 5500 5220
rect 5900 5380 6300 5500
rect 5900 5220 6020 5380
rect 6180 5220 6300 5380
rect 5900 5100 6300 5220
rect 6700 5380 7100 5500
rect 6700 5220 6820 5380
rect 6980 5220 7100 5380
rect 6700 5100 7100 5220
rect 7500 5380 7900 5500
rect 7500 5220 7620 5380
rect 7780 5220 7900 5380
rect 7500 5100 7900 5220
rect 8300 5380 8700 5500
rect 8300 5220 8420 5380
rect 8580 5220 8700 5380
rect 8300 5100 8700 5220
rect 9100 5380 9500 5500
rect 9100 5220 9220 5380
rect 9380 5220 9500 5380
rect 9100 5100 9500 5220
rect 9900 5380 10300 5500
rect 9900 5220 10020 5380
rect 10180 5220 10300 5380
rect 9900 5100 10300 5220
rect 10700 5380 11100 5500
rect 10700 5220 10820 5380
rect 10980 5220 11100 5380
rect 10700 5100 11100 5220
rect 11500 5380 11900 5500
rect 11500 5220 11620 5380
rect 11780 5220 11900 5380
rect 11500 5100 11900 5220
rect 12300 5380 12700 5500
rect 12300 5220 12420 5380
rect 12580 5220 12700 5380
rect 12300 5100 12700 5220
rect 13100 5380 13500 5500
rect 13100 5220 13220 5380
rect 13380 5220 13500 5380
rect 13100 5100 13500 5220
rect 13900 5380 14300 5500
rect 13900 5220 14020 5380
rect 14180 5220 14300 5380
rect 13900 5100 14300 5220
rect 14700 5380 15100 5500
rect 14700 5220 14820 5380
rect 14980 5220 15100 5380
rect 14700 5100 15100 5220
rect 15500 5380 15900 5500
rect 15500 5220 15620 5380
rect 15780 5220 15900 5380
rect 15500 5100 15900 5220
rect 700 4980 1100 5100
rect 700 4820 820 4980
rect 980 4820 1100 4980
rect 700 4700 1100 4820
rect 1500 4980 1900 5100
rect 1500 4820 1620 4980
rect 1780 4820 1900 4980
rect 1500 4700 1900 4820
rect 2300 4980 2700 5100
rect 2300 4820 2420 4980
rect 2580 4820 2700 4980
rect 2300 4700 2700 4820
rect 3100 4980 3500 5100
rect 3100 4820 3220 4980
rect 3380 4820 3500 4980
rect 3100 4700 3500 4820
rect 3900 4980 4300 5100
rect 3900 4820 4020 4980
rect 4180 4820 4300 4980
rect 3900 4700 4300 4820
rect 4700 4980 5100 5100
rect 4700 4820 4820 4980
rect 4980 4820 5100 4980
rect 4700 4700 5100 4820
rect 5500 4980 5900 5100
rect 5500 4820 5620 4980
rect 5780 4820 5900 4980
rect 5500 4700 5900 4820
rect 6300 4980 6700 5100
rect 6300 4820 6420 4980
rect 6580 4820 6700 4980
rect 6300 4700 6700 4820
rect 7100 4980 7500 5100
rect 7100 4820 7220 4980
rect 7380 4820 7500 4980
rect 7100 4700 7500 4820
rect 7900 4980 8300 5100
rect 7900 4820 8020 4980
rect 8180 4820 8300 4980
rect 7900 4700 8300 4820
rect 8700 4980 9100 5100
rect 8700 4820 8820 4980
rect 8980 4820 9100 4980
rect 8700 4700 9100 4820
rect 9500 4980 9900 5100
rect 9500 4820 9620 4980
rect 9780 4820 9900 4980
rect 9500 4700 9900 4820
rect 10300 4980 10700 5100
rect 10300 4820 10420 4980
rect 10580 4820 10700 4980
rect 10300 4700 10700 4820
rect 11100 4980 11500 5100
rect 11100 4820 11220 4980
rect 11380 4820 11500 4980
rect 11100 4700 11500 4820
rect 11900 4980 12300 5100
rect 11900 4820 12020 4980
rect 12180 4820 12300 4980
rect 11900 4700 12300 4820
rect 12700 4980 13100 5100
rect 12700 4820 12820 4980
rect 12980 4820 13100 4980
rect 12700 4700 13100 4820
rect 13500 4980 13900 5100
rect 13500 4820 13620 4980
rect 13780 4820 13900 4980
rect 13500 4700 13900 4820
rect 14300 4980 14700 5100
rect 14300 4820 14420 4980
rect 14580 4820 14700 4980
rect 14300 4700 14700 4820
rect 15100 4980 15500 5100
rect 15100 4820 15220 4980
rect 15380 4820 15500 4980
rect 15100 4700 15500 4820
rect 15900 4980 16300 5100
rect 15900 4820 16020 4980
rect 16180 4820 16300 4980
rect 15900 4700 16300 4820
rect 1100 4580 1500 4700
rect 1100 4420 1220 4580
rect 1380 4420 1500 4580
rect 1100 4300 1500 4420
rect 1900 4580 2300 4700
rect 1900 4420 2020 4580
rect 2180 4420 2300 4580
rect 1900 4300 2300 4420
rect 2700 4580 3100 4700
rect 2700 4420 2820 4580
rect 2980 4420 3100 4580
rect 2700 4300 3100 4420
rect 3500 4580 3900 4700
rect 3500 4420 3620 4580
rect 3780 4420 3900 4580
rect 3500 4300 3900 4420
rect 4300 4580 4700 4700
rect 4300 4420 4420 4580
rect 4580 4420 4700 4580
rect 4300 4300 4700 4420
rect 5100 4580 5500 4700
rect 5100 4420 5220 4580
rect 5380 4420 5500 4580
rect 5100 4300 5500 4420
rect 5900 4580 6300 4700
rect 5900 4420 6020 4580
rect 6180 4420 6300 4580
rect 5900 4300 6300 4420
rect 6700 4580 7100 4700
rect 6700 4420 6820 4580
rect 6980 4420 7100 4580
rect 6700 4300 7100 4420
rect 7500 4580 7900 4700
rect 7500 4420 7620 4580
rect 7780 4420 7900 4580
rect 7500 4300 7900 4420
rect 8300 4580 8700 4700
rect 8300 4420 8420 4580
rect 8580 4420 8700 4580
rect 8300 4300 8700 4420
rect 9100 4580 9500 4700
rect 9100 4420 9220 4580
rect 9380 4420 9500 4580
rect 9100 4300 9500 4420
rect 9900 4580 10300 4700
rect 9900 4420 10020 4580
rect 10180 4420 10300 4580
rect 9900 4300 10300 4420
rect 10700 4580 11100 4700
rect 10700 4420 10820 4580
rect 10980 4420 11100 4580
rect 10700 4300 11100 4420
rect 11500 4580 11900 4700
rect 11500 4420 11620 4580
rect 11780 4420 11900 4580
rect 11500 4300 11900 4420
rect 12300 4580 12700 4700
rect 12300 4420 12420 4580
rect 12580 4420 12700 4580
rect 12300 4300 12700 4420
rect 13100 4580 13500 4700
rect 13100 4420 13220 4580
rect 13380 4420 13500 4580
rect 13100 4300 13500 4420
rect 13900 4580 14300 4700
rect 13900 4420 14020 4580
rect 14180 4420 14300 4580
rect 13900 4300 14300 4420
rect 14700 4580 15100 4700
rect 14700 4420 14820 4580
rect 14980 4420 15100 4580
rect 14700 4300 15100 4420
rect 15500 4580 15900 4700
rect 15500 4420 15620 4580
rect 15780 4420 15900 4580
rect 15500 4300 15900 4420
rect 700 4180 1100 4300
rect 700 4020 820 4180
rect 980 4020 1100 4180
rect 700 3900 1100 4020
rect 1500 4180 1900 4300
rect 1500 4020 1620 4180
rect 1780 4020 1900 4180
rect 1500 3900 1900 4020
rect 2300 4180 2700 4300
rect 2300 4020 2420 4180
rect 2580 4020 2700 4180
rect 2300 3900 2700 4020
rect 3100 4180 3500 4300
rect 3100 4020 3220 4180
rect 3380 4020 3500 4180
rect 3100 3900 3500 4020
rect 3900 4180 4300 4300
rect 3900 4020 4020 4180
rect 4180 4020 4300 4180
rect 3900 3900 4300 4020
rect 4700 4180 5100 4300
rect 4700 4020 4820 4180
rect 4980 4020 5100 4180
rect 4700 3900 5100 4020
rect 5500 4180 5900 4300
rect 5500 4020 5620 4180
rect 5780 4020 5900 4180
rect 5500 3900 5900 4020
rect 6300 4180 6700 4300
rect 6300 4020 6420 4180
rect 6580 4020 6700 4180
rect 6300 3900 6700 4020
rect 7100 4180 7500 4300
rect 7100 4020 7220 4180
rect 7380 4020 7500 4180
rect 7100 3900 7500 4020
rect 7900 4180 8300 4300
rect 7900 4020 8020 4180
rect 8180 4020 8300 4180
rect 7900 3900 8300 4020
rect 8700 4180 9100 4300
rect 8700 4020 8820 4180
rect 8980 4020 9100 4180
rect 8700 3900 9100 4020
rect 9500 4180 9900 4300
rect 9500 4020 9620 4180
rect 9780 4020 9900 4180
rect 9500 3900 9900 4020
rect 10300 4180 10700 4300
rect 10300 4020 10420 4180
rect 10580 4020 10700 4180
rect 10300 3900 10700 4020
rect 11100 4180 11500 4300
rect 11100 4020 11220 4180
rect 11380 4020 11500 4180
rect 11100 3900 11500 4020
rect 11900 4180 12300 4300
rect 11900 4020 12020 4180
rect 12180 4020 12300 4180
rect 11900 3900 12300 4020
rect 12700 4180 13100 4300
rect 12700 4020 12820 4180
rect 12980 4020 13100 4180
rect 12700 3900 13100 4020
rect 13500 4180 13900 4300
rect 13500 4020 13620 4180
rect 13780 4020 13900 4180
rect 13500 3900 13900 4020
rect 14300 4180 14700 4300
rect 14300 4020 14420 4180
rect 14580 4020 14700 4180
rect 14300 3900 14700 4020
rect 15100 4180 15500 4300
rect 15100 4020 15220 4180
rect 15380 4020 15500 4180
rect 15100 3900 15500 4020
rect 15900 4180 16300 4300
rect 15900 4020 16020 4180
rect 16180 4020 16300 4180
rect 15900 3900 16300 4020
rect 1100 3780 1500 3900
rect 1100 3620 1220 3780
rect 1380 3620 1500 3780
rect 1100 3500 1500 3620
rect 1900 3780 2300 3900
rect 1900 3620 2020 3780
rect 2180 3620 2300 3780
rect 1900 3500 2300 3620
rect 2700 3780 3100 3900
rect 2700 3620 2820 3780
rect 2980 3620 3100 3780
rect 2700 3500 3100 3620
rect 3500 3780 3900 3900
rect 3500 3620 3620 3780
rect 3780 3620 3900 3780
rect 3500 3500 3900 3620
rect 4300 3780 4700 3900
rect 4300 3620 4420 3780
rect 4580 3620 4700 3780
rect 4300 3500 4700 3620
rect 5100 3780 5500 3900
rect 5100 3620 5220 3780
rect 5380 3620 5500 3780
rect 5100 3500 5500 3620
rect 5900 3780 6300 3900
rect 5900 3620 6020 3780
rect 6180 3620 6300 3780
rect 5900 3500 6300 3620
rect 6700 3780 7100 3900
rect 6700 3620 6820 3780
rect 6980 3620 7100 3780
rect 6700 3500 7100 3620
rect 7500 3780 7900 3900
rect 7500 3620 7620 3780
rect 7780 3620 7900 3780
rect 7500 3500 7900 3620
rect 8300 3780 8700 3900
rect 8300 3620 8420 3780
rect 8580 3620 8700 3780
rect 8300 3500 8700 3620
rect 9100 3780 9500 3900
rect 9100 3620 9220 3780
rect 9380 3620 9500 3780
rect 9100 3500 9500 3620
rect 9900 3780 10300 3900
rect 9900 3620 10020 3780
rect 10180 3620 10300 3780
rect 9900 3500 10300 3620
rect 10700 3780 11100 3900
rect 10700 3620 10820 3780
rect 10980 3620 11100 3780
rect 10700 3500 11100 3620
rect 11500 3780 11900 3900
rect 11500 3620 11620 3780
rect 11780 3620 11900 3780
rect 11500 3500 11900 3620
rect 12300 3780 12700 3900
rect 12300 3620 12420 3780
rect 12580 3620 12700 3780
rect 12300 3500 12700 3620
rect 13100 3780 13500 3900
rect 13100 3620 13220 3780
rect 13380 3620 13500 3780
rect 13100 3500 13500 3620
rect 13900 3780 14300 3900
rect 13900 3620 14020 3780
rect 14180 3620 14300 3780
rect 13900 3500 14300 3620
rect 14700 3780 15100 3900
rect 14700 3620 14820 3780
rect 14980 3620 15100 3780
rect 14700 3500 15100 3620
rect 15500 3780 15900 3900
rect 15500 3620 15620 3780
rect 15780 3620 15900 3780
rect 15500 3500 15900 3620
rect 700 3380 1100 3500
rect 700 3220 820 3380
rect 980 3220 1100 3380
rect 700 3100 1100 3220
rect 1500 3380 1900 3500
rect 1500 3220 1620 3380
rect 1780 3220 1900 3380
rect 1500 3100 1900 3220
rect 2300 3380 2700 3500
rect 2300 3220 2420 3380
rect 2580 3220 2700 3380
rect 2300 3100 2700 3220
rect 3100 3380 3500 3500
rect 3100 3220 3220 3380
rect 3380 3220 3500 3380
rect 3100 3100 3500 3220
rect 3900 3380 4300 3500
rect 3900 3220 4020 3380
rect 4180 3220 4300 3380
rect 3900 3100 4300 3220
rect 4700 3380 5100 3500
rect 4700 3220 4820 3380
rect 4980 3220 5100 3380
rect 4700 3100 5100 3220
rect 5500 3380 5900 3500
rect 5500 3220 5620 3380
rect 5780 3220 5900 3380
rect 5500 3100 5900 3220
rect 6300 3380 6700 3500
rect 6300 3220 6420 3380
rect 6580 3220 6700 3380
rect 6300 3100 6700 3220
rect 7100 3380 7500 3500
rect 7100 3220 7220 3380
rect 7380 3220 7500 3380
rect 7100 3100 7500 3220
rect 7900 3380 8300 3500
rect 7900 3220 8020 3380
rect 8180 3220 8300 3380
rect 7900 3100 8300 3220
rect 8700 3380 9100 3500
rect 8700 3220 8820 3380
rect 8980 3220 9100 3380
rect 8700 3100 9100 3220
rect 9500 3380 9900 3500
rect 9500 3220 9620 3380
rect 9780 3220 9900 3380
rect 9500 3100 9900 3220
rect 10300 3380 10700 3500
rect 10300 3220 10420 3380
rect 10580 3220 10700 3380
rect 10300 3100 10700 3220
rect 11100 3380 11500 3500
rect 11100 3220 11220 3380
rect 11380 3220 11500 3380
rect 11100 3100 11500 3220
rect 11900 3380 12300 3500
rect 11900 3220 12020 3380
rect 12180 3220 12300 3380
rect 11900 3100 12300 3220
rect 12700 3380 13100 3500
rect 12700 3220 12820 3380
rect 12980 3220 13100 3380
rect 12700 3100 13100 3220
rect 13500 3380 13900 3500
rect 13500 3220 13620 3380
rect 13780 3220 13900 3380
rect 13500 3100 13900 3220
rect 14300 3380 14700 3500
rect 14300 3220 14420 3380
rect 14580 3220 14700 3380
rect 14300 3100 14700 3220
rect 15100 3380 15500 3500
rect 15100 3220 15220 3380
rect 15380 3220 15500 3380
rect 15100 3100 15500 3220
rect 15900 3380 16300 3500
rect 15900 3220 16020 3380
rect 16180 3220 16300 3380
rect 15900 3100 16300 3220
rect 1100 2980 1500 3100
rect 1100 2820 1220 2980
rect 1380 2820 1500 2980
rect 1100 2700 1500 2820
rect 1900 2980 2300 3100
rect 1900 2820 2020 2980
rect 2180 2820 2300 2980
rect 1900 2700 2300 2820
rect 2700 2980 3100 3100
rect 2700 2820 2820 2980
rect 2980 2820 3100 2980
rect 2700 2700 3100 2820
rect 3500 2980 3900 3100
rect 3500 2820 3620 2980
rect 3780 2820 3900 2980
rect 3500 2700 3900 2820
rect 4300 2980 4700 3100
rect 4300 2820 4420 2980
rect 4580 2820 4700 2980
rect 4300 2700 4700 2820
rect 5100 2980 5500 3100
rect 5100 2820 5220 2980
rect 5380 2820 5500 2980
rect 5100 2700 5500 2820
rect 5900 2980 6300 3100
rect 5900 2820 6020 2980
rect 6180 2820 6300 2980
rect 5900 2700 6300 2820
rect 6700 2980 7100 3100
rect 6700 2820 6820 2980
rect 6980 2820 7100 2980
rect 6700 2700 7100 2820
rect 7500 2980 7900 3100
rect 7500 2820 7620 2980
rect 7780 2820 7900 2980
rect 7500 2700 7900 2820
rect 8300 2980 8700 3100
rect 8300 2820 8420 2980
rect 8580 2820 8700 2980
rect 8300 2700 8700 2820
rect 9100 2980 9500 3100
rect 9100 2820 9220 2980
rect 9380 2820 9500 2980
rect 9100 2700 9500 2820
rect 9900 2980 10300 3100
rect 9900 2820 10020 2980
rect 10180 2820 10300 2980
rect 9900 2700 10300 2820
rect 10700 2980 11100 3100
rect 10700 2820 10820 2980
rect 10980 2820 11100 2980
rect 10700 2700 11100 2820
rect 11500 2980 11900 3100
rect 11500 2820 11620 2980
rect 11780 2820 11900 2980
rect 11500 2700 11900 2820
rect 12300 2980 12700 3100
rect 12300 2820 12420 2980
rect 12580 2820 12700 2980
rect 12300 2700 12700 2820
rect 13100 2980 13500 3100
rect 13100 2820 13220 2980
rect 13380 2820 13500 2980
rect 13100 2700 13500 2820
rect 13900 2980 14300 3100
rect 13900 2820 14020 2980
rect 14180 2820 14300 2980
rect 13900 2700 14300 2820
rect 14700 2980 15100 3100
rect 14700 2820 14820 2980
rect 14980 2820 15100 2980
rect 14700 2700 15100 2820
rect 15500 2980 15900 3100
rect 15500 2820 15620 2980
rect 15780 2820 15900 2980
rect 15500 2700 15900 2820
rect 700 2580 1100 2700
rect 700 2420 820 2580
rect 980 2420 1100 2580
rect 700 2300 1100 2420
rect 1500 2580 1900 2700
rect 1500 2420 1620 2580
rect 1780 2420 1900 2580
rect 1500 2300 1900 2420
rect 2300 2580 2700 2700
rect 2300 2420 2420 2580
rect 2580 2420 2700 2580
rect 2300 2300 2700 2420
rect 3100 2580 3500 2700
rect 3100 2420 3220 2580
rect 3380 2420 3500 2580
rect 3100 2300 3500 2420
rect 3900 2580 4300 2700
rect 3900 2420 4020 2580
rect 4180 2420 4300 2580
rect 3900 2300 4300 2420
rect 4700 2580 5100 2700
rect 4700 2420 4820 2580
rect 4980 2420 5100 2580
rect 4700 2300 5100 2420
rect 5500 2580 5900 2700
rect 5500 2420 5620 2580
rect 5780 2420 5900 2580
rect 5500 2300 5900 2420
rect 6300 2580 6700 2700
rect 6300 2420 6420 2580
rect 6580 2420 6700 2580
rect 6300 2300 6700 2420
rect 7100 2580 7500 2700
rect 7100 2420 7220 2580
rect 7380 2420 7500 2580
rect 7100 2300 7500 2420
rect 7900 2580 8300 2700
rect 7900 2420 8020 2580
rect 8180 2420 8300 2580
rect 7900 2300 8300 2420
rect 8700 2580 9100 2700
rect 8700 2420 8820 2580
rect 8980 2420 9100 2580
rect 8700 2300 9100 2420
rect 9500 2580 9900 2700
rect 9500 2420 9620 2580
rect 9780 2420 9900 2580
rect 9500 2300 9900 2420
rect 10300 2580 10700 2700
rect 10300 2420 10420 2580
rect 10580 2420 10700 2580
rect 10300 2300 10700 2420
rect 11100 2580 11500 2700
rect 11100 2420 11220 2580
rect 11380 2420 11500 2580
rect 11100 2300 11500 2420
rect 11900 2580 12300 2700
rect 11900 2420 12020 2580
rect 12180 2420 12300 2580
rect 11900 2300 12300 2420
rect 12700 2580 13100 2700
rect 12700 2420 12820 2580
rect 12980 2420 13100 2580
rect 12700 2300 13100 2420
rect 13500 2580 13900 2700
rect 13500 2420 13620 2580
rect 13780 2420 13900 2580
rect 13500 2300 13900 2420
rect 14300 2580 14700 2700
rect 14300 2420 14420 2580
rect 14580 2420 14700 2580
rect 14300 2300 14700 2420
rect 15100 2580 15500 2700
rect 15100 2420 15220 2580
rect 15380 2420 15500 2580
rect 15100 2300 15500 2420
rect 15900 2580 16300 2700
rect 15900 2420 16020 2580
rect 16180 2420 16300 2580
rect 15900 2300 16300 2420
rect 1100 2180 1500 2300
rect 1100 2020 1220 2180
rect 1380 2020 1500 2180
rect 1100 1900 1500 2020
rect 1900 2180 2300 2300
rect 1900 2020 2020 2180
rect 2180 2020 2300 2180
rect 1900 1900 2300 2020
rect 2700 2180 3100 2300
rect 2700 2020 2820 2180
rect 2980 2020 3100 2180
rect 2700 1900 3100 2020
rect 3500 2180 3900 2300
rect 3500 2020 3620 2180
rect 3780 2020 3900 2180
rect 3500 1900 3900 2020
rect 4300 2180 4700 2300
rect 4300 2020 4420 2180
rect 4580 2020 4700 2180
rect 4300 1900 4700 2020
rect 5100 2180 5500 2300
rect 5100 2020 5220 2180
rect 5380 2020 5500 2180
rect 5100 1900 5500 2020
rect 5900 2180 6300 2300
rect 5900 2020 6020 2180
rect 6180 2020 6300 2180
rect 5900 1900 6300 2020
rect 6700 2180 7100 2300
rect 6700 2020 6820 2180
rect 6980 2020 7100 2180
rect 6700 1900 7100 2020
rect 7500 2180 7900 2300
rect 7500 2020 7620 2180
rect 7780 2020 7900 2180
rect 7500 1900 7900 2020
rect 8300 2180 8700 2300
rect 8300 2020 8420 2180
rect 8580 2020 8700 2180
rect 8300 1900 8700 2020
rect 9100 2180 9500 2300
rect 9100 2020 9220 2180
rect 9380 2020 9500 2180
rect 9100 1900 9500 2020
rect 9900 2180 10300 2300
rect 9900 2020 10020 2180
rect 10180 2020 10300 2180
rect 9900 1900 10300 2020
rect 10700 2180 11100 2300
rect 10700 2020 10820 2180
rect 10980 2020 11100 2180
rect 10700 1900 11100 2020
rect 11500 2180 11900 2300
rect 11500 2020 11620 2180
rect 11780 2020 11900 2180
rect 11500 1900 11900 2020
rect 12300 2180 12700 2300
rect 12300 2020 12420 2180
rect 12580 2020 12700 2180
rect 12300 1900 12700 2020
rect 13100 2180 13500 2300
rect 13100 2020 13220 2180
rect 13380 2020 13500 2180
rect 13100 1900 13500 2020
rect 13900 2180 14300 2300
rect 13900 2020 14020 2180
rect 14180 2020 14300 2180
rect 13900 1900 14300 2020
rect 14700 2180 15100 2300
rect 14700 2020 14820 2180
rect 14980 2020 15100 2180
rect 14700 1900 15100 2020
rect 15500 2180 15900 2300
rect 15500 2020 15620 2180
rect 15780 2020 15900 2180
rect 15500 1900 15900 2020
rect 700 1780 1100 1900
rect 700 1620 820 1780
rect 980 1620 1100 1780
rect 700 1500 1100 1620
rect 1500 1780 1900 1900
rect 1500 1620 1620 1780
rect 1780 1620 1900 1780
rect 1500 1500 1900 1620
rect 2300 1780 2700 1900
rect 2300 1620 2420 1780
rect 2580 1620 2700 1780
rect 2300 1500 2700 1620
rect 3100 1780 3500 1900
rect 3100 1620 3220 1780
rect 3380 1620 3500 1780
rect 3100 1500 3500 1620
rect 3900 1780 4300 1900
rect 3900 1620 4020 1780
rect 4180 1620 4300 1780
rect 3900 1500 4300 1620
rect 4700 1780 5100 1900
rect 4700 1620 4820 1780
rect 4980 1620 5100 1780
rect 4700 1500 5100 1620
rect 5500 1780 5900 1900
rect 5500 1620 5620 1780
rect 5780 1620 5900 1780
rect 5500 1500 5900 1620
rect 6300 1780 6700 1900
rect 6300 1620 6420 1780
rect 6580 1620 6700 1780
rect 6300 1500 6700 1620
rect 7100 1780 7500 1900
rect 7100 1620 7220 1780
rect 7380 1620 7500 1780
rect 7100 1500 7500 1620
rect 7900 1780 8300 1900
rect 7900 1620 8020 1780
rect 8180 1620 8300 1780
rect 7900 1500 8300 1620
rect 8700 1780 9100 1900
rect 8700 1620 8820 1780
rect 8980 1620 9100 1780
rect 8700 1500 9100 1620
rect 9500 1780 9900 1900
rect 9500 1620 9620 1780
rect 9780 1620 9900 1780
rect 9500 1500 9900 1620
rect 10300 1780 10700 1900
rect 10300 1620 10420 1780
rect 10580 1620 10700 1780
rect 10300 1500 10700 1620
rect 11100 1780 11500 1900
rect 11100 1620 11220 1780
rect 11380 1620 11500 1780
rect 11100 1500 11500 1620
rect 11900 1780 12300 1900
rect 11900 1620 12020 1780
rect 12180 1620 12300 1780
rect 11900 1500 12300 1620
rect 12700 1780 13100 1900
rect 12700 1620 12820 1780
rect 12980 1620 13100 1780
rect 12700 1500 13100 1620
rect 13500 1780 13900 1900
rect 13500 1620 13620 1780
rect 13780 1620 13900 1780
rect 13500 1500 13900 1620
rect 14300 1780 14700 1900
rect 14300 1620 14420 1780
rect 14580 1620 14700 1780
rect 14300 1500 14700 1620
rect 15100 1780 15500 1900
rect 15100 1620 15220 1780
rect 15380 1620 15500 1780
rect 15100 1500 15500 1620
rect 15900 1780 16300 1900
rect 15900 1620 16020 1780
rect 16180 1620 16300 1780
rect 15900 1500 16300 1620
rect 1100 1380 1500 1500
rect 1100 1220 1220 1380
rect 1380 1220 1500 1380
rect 1100 1100 1500 1220
rect 1900 1380 2300 1500
rect 1900 1220 2020 1380
rect 2180 1220 2300 1380
rect 1900 1100 2300 1220
rect 2700 1380 3100 1500
rect 2700 1220 2820 1380
rect 2980 1220 3100 1380
rect 2700 1100 3100 1220
rect 3500 1380 3900 1500
rect 3500 1220 3620 1380
rect 3780 1220 3900 1380
rect 3500 1100 3900 1220
rect 4300 1380 4700 1500
rect 4300 1220 4420 1380
rect 4580 1220 4700 1380
rect 4300 1100 4700 1220
rect 5100 1380 5500 1500
rect 5100 1220 5220 1380
rect 5380 1220 5500 1380
rect 5100 1100 5500 1220
rect 5900 1380 6300 1500
rect 5900 1220 6020 1380
rect 6180 1220 6300 1380
rect 5900 1100 6300 1220
rect 6700 1380 7100 1500
rect 6700 1220 6820 1380
rect 6980 1220 7100 1380
rect 6700 1100 7100 1220
rect 7500 1380 7900 1500
rect 7500 1220 7620 1380
rect 7780 1220 7900 1380
rect 7500 1100 7900 1220
rect 8300 1380 8700 1500
rect 8300 1220 8420 1380
rect 8580 1220 8700 1380
rect 8300 1100 8700 1220
rect 9100 1380 9500 1500
rect 9100 1220 9220 1380
rect 9380 1220 9500 1380
rect 9100 1100 9500 1220
rect 9900 1380 10300 1500
rect 9900 1220 10020 1380
rect 10180 1220 10300 1380
rect 9900 1100 10300 1220
rect 10700 1380 11100 1500
rect 10700 1220 10820 1380
rect 10980 1220 11100 1380
rect 10700 1100 11100 1220
rect 11500 1380 11900 1500
rect 11500 1220 11620 1380
rect 11780 1220 11900 1380
rect 11500 1100 11900 1220
rect 12300 1380 12700 1500
rect 12300 1220 12420 1380
rect 12580 1220 12700 1380
rect 12300 1100 12700 1220
rect 13100 1380 13500 1500
rect 13100 1220 13220 1380
rect 13380 1220 13500 1380
rect 13100 1100 13500 1220
rect 13900 1380 14300 1500
rect 13900 1220 14020 1380
rect 14180 1220 14300 1380
rect 13900 1100 14300 1220
rect 14700 1380 15100 1500
rect 14700 1220 14820 1380
rect 14980 1220 15100 1380
rect 14700 1100 15100 1220
rect 15500 1380 15900 1500
rect 15500 1220 15620 1380
rect 15780 1220 15900 1380
rect 15500 1100 15900 1220
rect 700 980 1100 1100
rect 700 820 820 980
rect 980 820 1100 980
rect 700 700 1100 820
rect 1500 980 1900 1100
rect 1500 820 1620 980
rect 1780 820 1900 980
rect 1500 700 1900 820
rect 2300 980 2700 1100
rect 2300 820 2420 980
rect 2580 820 2700 980
rect 2300 700 2700 820
rect 3100 980 3500 1100
rect 3100 820 3220 980
rect 3380 820 3500 980
rect 3100 700 3500 820
rect 3900 980 4300 1100
rect 3900 820 4020 980
rect 4180 820 4300 980
rect 3900 700 4300 820
rect 4700 980 5100 1100
rect 4700 820 4820 980
rect 4980 820 5100 980
rect 4700 700 5100 820
rect 5500 980 5900 1100
rect 5500 820 5620 980
rect 5780 820 5900 980
rect 5500 700 5900 820
rect 6300 980 6700 1100
rect 6300 820 6420 980
rect 6580 820 6700 980
rect 6300 700 6700 820
rect 7100 980 7500 1100
rect 7100 820 7220 980
rect 7380 820 7500 980
rect 7100 700 7500 820
rect 7900 980 8300 1100
rect 7900 820 8020 980
rect 8180 820 8300 980
rect 7900 700 8300 820
rect 8700 980 9100 1100
rect 8700 820 8820 980
rect 8980 820 9100 980
rect 8700 700 9100 820
rect 9500 980 9900 1100
rect 9500 820 9620 980
rect 9780 820 9900 980
rect 9500 700 9900 820
rect 10300 980 10700 1100
rect 10300 820 10420 980
rect 10580 820 10700 980
rect 10300 700 10700 820
rect 11100 980 11500 1100
rect 11100 820 11220 980
rect 11380 820 11500 980
rect 11100 700 11500 820
rect 11900 980 12300 1100
rect 11900 820 12020 980
rect 12180 820 12300 980
rect 11900 700 12300 820
rect 12700 980 13100 1100
rect 12700 820 12820 980
rect 12980 820 13100 980
rect 12700 700 13100 820
rect 13500 980 13900 1100
rect 13500 820 13620 980
rect 13780 820 13900 980
rect 13500 700 13900 820
rect 14300 980 14700 1100
rect 14300 820 14420 980
rect 14580 820 14700 980
rect 14300 700 14700 820
rect 15100 980 15500 1100
rect 15100 820 15220 980
rect 15380 820 15500 980
rect 15100 700 15500 820
rect 15900 980 16300 1100
rect 15900 820 16020 980
rect 16180 820 16300 980
rect 15900 700 16300 820
rect 16500 500 17000 16500
rect 0 0 17000 500
<< m3contact >>
rect 1220 15620 1380 15780
rect 2020 15620 2180 15780
rect 2820 15620 2980 15780
rect 3620 15620 3780 15780
rect 4420 15620 4580 15780
rect 5220 15620 5380 15780
rect 6020 15620 6180 15780
rect 6820 15620 6980 15780
rect 7620 15620 7780 15780
rect 8420 15620 8580 15780
rect 9220 15620 9380 15780
rect 10020 15620 10180 15780
rect 10820 15620 10980 15780
rect 11620 15620 11780 15780
rect 12420 15620 12580 15780
rect 13220 15620 13380 15780
rect 14020 15620 14180 15780
rect 14820 15620 14980 15780
rect 15620 15620 15780 15780
rect 1220 14820 1380 14980
rect 2020 14820 2180 14980
rect 2820 14820 2980 14980
rect 3620 14820 3780 14980
rect 4420 14820 4580 14980
rect 5220 14820 5380 14980
rect 6020 14820 6180 14980
rect 6820 14820 6980 14980
rect 7620 14820 7780 14980
rect 8420 14820 8580 14980
rect 9220 14820 9380 14980
rect 10020 14820 10180 14980
rect 10820 14820 10980 14980
rect 11620 14820 11780 14980
rect 12420 14820 12580 14980
rect 13220 14820 13380 14980
rect 14020 14820 14180 14980
rect 14820 14820 14980 14980
rect 15620 14820 15780 14980
rect 1220 14020 1380 14180
rect 2020 14020 2180 14180
rect 2820 14020 2980 14180
rect 3620 14020 3780 14180
rect 4420 14020 4580 14180
rect 5220 14020 5380 14180
rect 6020 14020 6180 14180
rect 6820 14020 6980 14180
rect 7620 14020 7780 14180
rect 8420 14020 8580 14180
rect 9220 14020 9380 14180
rect 10020 14020 10180 14180
rect 10820 14020 10980 14180
rect 11620 14020 11780 14180
rect 12420 14020 12580 14180
rect 13220 14020 13380 14180
rect 14020 14020 14180 14180
rect 14820 14020 14980 14180
rect 15620 14020 15780 14180
rect 1220 13220 1380 13380
rect 2020 13220 2180 13380
rect 2820 13220 2980 13380
rect 3620 13220 3780 13380
rect 4420 13220 4580 13380
rect 5220 13220 5380 13380
rect 6020 13220 6180 13380
rect 6820 13220 6980 13380
rect 7620 13220 7780 13380
rect 8420 13220 8580 13380
rect 9220 13220 9380 13380
rect 10020 13220 10180 13380
rect 10820 13220 10980 13380
rect 11620 13220 11780 13380
rect 12420 13220 12580 13380
rect 13220 13220 13380 13380
rect 14020 13220 14180 13380
rect 14820 13220 14980 13380
rect 15620 13220 15780 13380
rect 1220 12420 1380 12580
rect 2020 12420 2180 12580
rect 2820 12420 2980 12580
rect 3620 12420 3780 12580
rect 4420 12420 4580 12580
rect 5220 12420 5380 12580
rect 6020 12420 6180 12580
rect 6820 12420 6980 12580
rect 7620 12420 7780 12580
rect 8420 12420 8580 12580
rect 9220 12420 9380 12580
rect 10020 12420 10180 12580
rect 10820 12420 10980 12580
rect 11620 12420 11780 12580
rect 12420 12420 12580 12580
rect 13220 12420 13380 12580
rect 14020 12420 14180 12580
rect 14820 12420 14980 12580
rect 15620 12420 15780 12580
rect 1220 11620 1380 11780
rect 2020 11620 2180 11780
rect 2820 11620 2980 11780
rect 3620 11620 3780 11780
rect 4420 11620 4580 11780
rect 5220 11620 5380 11780
rect 6020 11620 6180 11780
rect 6820 11620 6980 11780
rect 7620 11620 7780 11780
rect 8420 11620 8580 11780
rect 9220 11620 9380 11780
rect 10020 11620 10180 11780
rect 10820 11620 10980 11780
rect 11620 11620 11780 11780
rect 12420 11620 12580 11780
rect 13220 11620 13380 11780
rect 14020 11620 14180 11780
rect 14820 11620 14980 11780
rect 15620 11620 15780 11780
rect 1220 10820 1380 10980
rect 2020 10820 2180 10980
rect 2820 10820 2980 10980
rect 3620 10820 3780 10980
rect 4420 10820 4580 10980
rect 5220 10820 5380 10980
rect 6020 10820 6180 10980
rect 6820 10820 6980 10980
rect 7620 10820 7780 10980
rect 8420 10820 8580 10980
rect 9220 10820 9380 10980
rect 10020 10820 10180 10980
rect 10820 10820 10980 10980
rect 11620 10820 11780 10980
rect 12420 10820 12580 10980
rect 13220 10820 13380 10980
rect 14020 10820 14180 10980
rect 14820 10820 14980 10980
rect 15620 10820 15780 10980
rect 1220 10020 1380 10180
rect 2020 10020 2180 10180
rect 2820 10020 2980 10180
rect 3620 10020 3780 10180
rect 4420 10020 4580 10180
rect 5220 10020 5380 10180
rect 6020 10020 6180 10180
rect 6820 10020 6980 10180
rect 7620 10020 7780 10180
rect 8420 10020 8580 10180
rect 9220 10020 9380 10180
rect 10020 10020 10180 10180
rect 10820 10020 10980 10180
rect 11620 10020 11780 10180
rect 12420 10020 12580 10180
rect 13220 10020 13380 10180
rect 14020 10020 14180 10180
rect 14820 10020 14980 10180
rect 15620 10020 15780 10180
rect 1220 9220 1380 9380
rect 2020 9220 2180 9380
rect 2820 9220 2980 9380
rect 3620 9220 3780 9380
rect 4420 9220 4580 9380
rect 5220 9220 5380 9380
rect 6020 9220 6180 9380
rect 6820 9220 6980 9380
rect 7620 9220 7780 9380
rect 8420 9220 8580 9380
rect 9220 9220 9380 9380
rect 10020 9220 10180 9380
rect 10820 9220 10980 9380
rect 11620 9220 11780 9380
rect 12420 9220 12580 9380
rect 13220 9220 13380 9380
rect 14020 9220 14180 9380
rect 14820 9220 14980 9380
rect 15620 9220 15780 9380
rect 1220 8420 1380 8580
rect 2020 8420 2180 8580
rect 2820 8420 2980 8580
rect 3620 8420 3780 8580
rect 4420 8420 4580 8580
rect 5220 8420 5380 8580
rect 6020 8420 6180 8580
rect 6820 8420 6980 8580
rect 7620 8420 7780 8580
rect 8420 8420 8580 8580
rect 9220 8420 9380 8580
rect 10020 8420 10180 8580
rect 10820 8420 10980 8580
rect 11620 8420 11780 8580
rect 12420 8420 12580 8580
rect 13220 8420 13380 8580
rect 14020 8420 14180 8580
rect 14820 8420 14980 8580
rect 15620 8420 15780 8580
rect 1220 7620 1380 7780
rect 2020 7620 2180 7780
rect 2820 7620 2980 7780
rect 3620 7620 3780 7780
rect 4420 7620 4580 7780
rect 5220 7620 5380 7780
rect 6020 7620 6180 7780
rect 6820 7620 6980 7780
rect 7620 7620 7780 7780
rect 8420 7620 8580 7780
rect 9220 7620 9380 7780
rect 10020 7620 10180 7780
rect 10820 7620 10980 7780
rect 11620 7620 11780 7780
rect 12420 7620 12580 7780
rect 13220 7620 13380 7780
rect 14020 7620 14180 7780
rect 14820 7620 14980 7780
rect 15620 7620 15780 7780
rect 1220 6820 1380 6980
rect 2020 6820 2180 6980
rect 2820 6820 2980 6980
rect 3620 6820 3780 6980
rect 4420 6820 4580 6980
rect 5220 6820 5380 6980
rect 6020 6820 6180 6980
rect 6820 6820 6980 6980
rect 7620 6820 7780 6980
rect 8420 6820 8580 6980
rect 9220 6820 9380 6980
rect 10020 6820 10180 6980
rect 10820 6820 10980 6980
rect 11620 6820 11780 6980
rect 12420 6820 12580 6980
rect 13220 6820 13380 6980
rect 14020 6820 14180 6980
rect 14820 6820 14980 6980
rect 15620 6820 15780 6980
rect 1220 6020 1380 6180
rect 2020 6020 2180 6180
rect 2820 6020 2980 6180
rect 3620 6020 3780 6180
rect 4420 6020 4580 6180
rect 5220 6020 5380 6180
rect 6020 6020 6180 6180
rect 6820 6020 6980 6180
rect 7620 6020 7780 6180
rect 8420 6020 8580 6180
rect 9220 6020 9380 6180
rect 10020 6020 10180 6180
rect 10820 6020 10980 6180
rect 11620 6020 11780 6180
rect 12420 6020 12580 6180
rect 13220 6020 13380 6180
rect 14020 6020 14180 6180
rect 14820 6020 14980 6180
rect 15620 6020 15780 6180
rect 1220 5220 1380 5380
rect 2020 5220 2180 5380
rect 2820 5220 2980 5380
rect 3620 5220 3780 5380
rect 4420 5220 4580 5380
rect 5220 5220 5380 5380
rect 6020 5220 6180 5380
rect 6820 5220 6980 5380
rect 7620 5220 7780 5380
rect 8420 5220 8580 5380
rect 9220 5220 9380 5380
rect 10020 5220 10180 5380
rect 10820 5220 10980 5380
rect 11620 5220 11780 5380
rect 12420 5220 12580 5380
rect 13220 5220 13380 5380
rect 14020 5220 14180 5380
rect 14820 5220 14980 5380
rect 15620 5220 15780 5380
rect 1220 4420 1380 4580
rect 2020 4420 2180 4580
rect 2820 4420 2980 4580
rect 3620 4420 3780 4580
rect 4420 4420 4580 4580
rect 5220 4420 5380 4580
rect 6020 4420 6180 4580
rect 6820 4420 6980 4580
rect 7620 4420 7780 4580
rect 8420 4420 8580 4580
rect 9220 4420 9380 4580
rect 10020 4420 10180 4580
rect 10820 4420 10980 4580
rect 11620 4420 11780 4580
rect 12420 4420 12580 4580
rect 13220 4420 13380 4580
rect 14020 4420 14180 4580
rect 14820 4420 14980 4580
rect 15620 4420 15780 4580
rect 1220 3620 1380 3780
rect 2020 3620 2180 3780
rect 2820 3620 2980 3780
rect 3620 3620 3780 3780
rect 4420 3620 4580 3780
rect 5220 3620 5380 3780
rect 6020 3620 6180 3780
rect 6820 3620 6980 3780
rect 7620 3620 7780 3780
rect 8420 3620 8580 3780
rect 9220 3620 9380 3780
rect 10020 3620 10180 3780
rect 10820 3620 10980 3780
rect 11620 3620 11780 3780
rect 12420 3620 12580 3780
rect 13220 3620 13380 3780
rect 14020 3620 14180 3780
rect 14820 3620 14980 3780
rect 15620 3620 15780 3780
rect 1220 2820 1380 2980
rect 2020 2820 2180 2980
rect 2820 2820 2980 2980
rect 3620 2820 3780 2980
rect 4420 2820 4580 2980
rect 5220 2820 5380 2980
rect 6020 2820 6180 2980
rect 6820 2820 6980 2980
rect 7620 2820 7780 2980
rect 8420 2820 8580 2980
rect 9220 2820 9380 2980
rect 10020 2820 10180 2980
rect 10820 2820 10980 2980
rect 11620 2820 11780 2980
rect 12420 2820 12580 2980
rect 13220 2820 13380 2980
rect 14020 2820 14180 2980
rect 14820 2820 14980 2980
rect 15620 2820 15780 2980
rect 1220 2020 1380 2180
rect 2020 2020 2180 2180
rect 2820 2020 2980 2180
rect 3620 2020 3780 2180
rect 4420 2020 4580 2180
rect 5220 2020 5380 2180
rect 6020 2020 6180 2180
rect 6820 2020 6980 2180
rect 7620 2020 7780 2180
rect 8420 2020 8580 2180
rect 9220 2020 9380 2180
rect 10020 2020 10180 2180
rect 10820 2020 10980 2180
rect 11620 2020 11780 2180
rect 12420 2020 12580 2180
rect 13220 2020 13380 2180
rect 14020 2020 14180 2180
rect 14820 2020 14980 2180
rect 15620 2020 15780 2180
rect 1220 1220 1380 1380
rect 2020 1220 2180 1380
rect 2820 1220 2980 1380
rect 3620 1220 3780 1380
rect 4420 1220 4580 1380
rect 5220 1220 5380 1380
rect 6020 1220 6180 1380
rect 6820 1220 6980 1380
rect 7620 1220 7780 1380
rect 8420 1220 8580 1380
rect 9220 1220 9380 1380
rect 10020 1220 10180 1380
rect 10820 1220 10980 1380
rect 11620 1220 11780 1380
rect 12420 1220 12580 1380
rect 13220 1220 13380 1380
rect 14020 1220 14180 1380
rect 14820 1220 14980 1380
rect 15620 1220 15780 1380
<< metal3 >>
rect 0 16500 17000 17000
rect 0 500 500 16500
rect 16500 500 17000 16500
rect 0 0 17000 500
<< pad >>
rect 500 15780 16500 16500
rect 500 15620 1220 15780
rect 1380 15620 2020 15780
rect 2180 15620 2820 15780
rect 2980 15620 3620 15780
rect 3780 15620 4420 15780
rect 4580 15620 5220 15780
rect 5380 15620 6020 15780
rect 6180 15620 6820 15780
rect 6980 15620 7620 15780
rect 7780 15620 8420 15780
rect 8580 15620 9220 15780
rect 9380 15620 10020 15780
rect 10180 15620 10820 15780
rect 10980 15620 11620 15780
rect 11780 15620 12420 15780
rect 12580 15620 13220 15780
rect 13380 15620 14020 15780
rect 14180 15620 14820 15780
rect 14980 15620 15620 15780
rect 15780 15620 16500 15780
rect 500 14980 16500 15620
rect 500 14820 1220 14980
rect 1380 14820 2020 14980
rect 2180 14820 2820 14980
rect 2980 14820 3620 14980
rect 3780 14820 4420 14980
rect 4580 14820 5220 14980
rect 5380 14820 6020 14980
rect 6180 14820 6820 14980
rect 6980 14820 7620 14980
rect 7780 14820 8420 14980
rect 8580 14820 9220 14980
rect 9380 14820 10020 14980
rect 10180 14820 10820 14980
rect 10980 14820 11620 14980
rect 11780 14820 12420 14980
rect 12580 14820 13220 14980
rect 13380 14820 14020 14980
rect 14180 14820 14820 14980
rect 14980 14820 15620 14980
rect 15780 14820 16500 14980
rect 500 14180 16500 14820
rect 500 14020 1220 14180
rect 1380 14020 2020 14180
rect 2180 14020 2820 14180
rect 2980 14020 3620 14180
rect 3780 14020 4420 14180
rect 4580 14020 5220 14180
rect 5380 14020 6020 14180
rect 6180 14020 6820 14180
rect 6980 14020 7620 14180
rect 7780 14020 8420 14180
rect 8580 14020 9220 14180
rect 9380 14020 10020 14180
rect 10180 14020 10820 14180
rect 10980 14020 11620 14180
rect 11780 14020 12420 14180
rect 12580 14020 13220 14180
rect 13380 14020 14020 14180
rect 14180 14020 14820 14180
rect 14980 14020 15620 14180
rect 15780 14020 16500 14180
rect 500 13380 16500 14020
rect 500 13220 1220 13380
rect 1380 13220 2020 13380
rect 2180 13220 2820 13380
rect 2980 13220 3620 13380
rect 3780 13220 4420 13380
rect 4580 13220 5220 13380
rect 5380 13220 6020 13380
rect 6180 13220 6820 13380
rect 6980 13220 7620 13380
rect 7780 13220 8420 13380
rect 8580 13220 9220 13380
rect 9380 13220 10020 13380
rect 10180 13220 10820 13380
rect 10980 13220 11620 13380
rect 11780 13220 12420 13380
rect 12580 13220 13220 13380
rect 13380 13220 14020 13380
rect 14180 13220 14820 13380
rect 14980 13220 15620 13380
rect 15780 13220 16500 13380
rect 500 12580 16500 13220
rect 500 12420 1220 12580
rect 1380 12420 2020 12580
rect 2180 12420 2820 12580
rect 2980 12420 3620 12580
rect 3780 12420 4420 12580
rect 4580 12420 5220 12580
rect 5380 12420 6020 12580
rect 6180 12420 6820 12580
rect 6980 12420 7620 12580
rect 7780 12420 8420 12580
rect 8580 12420 9220 12580
rect 9380 12420 10020 12580
rect 10180 12420 10820 12580
rect 10980 12420 11620 12580
rect 11780 12420 12420 12580
rect 12580 12420 13220 12580
rect 13380 12420 14020 12580
rect 14180 12420 14820 12580
rect 14980 12420 15620 12580
rect 15780 12420 16500 12580
rect 500 11780 16500 12420
rect 500 11620 1220 11780
rect 1380 11620 2020 11780
rect 2180 11620 2820 11780
rect 2980 11620 3620 11780
rect 3780 11620 4420 11780
rect 4580 11620 5220 11780
rect 5380 11620 6020 11780
rect 6180 11620 6820 11780
rect 6980 11620 7620 11780
rect 7780 11620 8420 11780
rect 8580 11620 9220 11780
rect 9380 11620 10020 11780
rect 10180 11620 10820 11780
rect 10980 11620 11620 11780
rect 11780 11620 12420 11780
rect 12580 11620 13220 11780
rect 13380 11620 14020 11780
rect 14180 11620 14820 11780
rect 14980 11620 15620 11780
rect 15780 11620 16500 11780
rect 500 10980 16500 11620
rect 500 10820 1220 10980
rect 1380 10820 2020 10980
rect 2180 10820 2820 10980
rect 2980 10820 3620 10980
rect 3780 10820 4420 10980
rect 4580 10820 5220 10980
rect 5380 10820 6020 10980
rect 6180 10820 6820 10980
rect 6980 10820 7620 10980
rect 7780 10820 8420 10980
rect 8580 10820 9220 10980
rect 9380 10820 10020 10980
rect 10180 10820 10820 10980
rect 10980 10820 11620 10980
rect 11780 10820 12420 10980
rect 12580 10820 13220 10980
rect 13380 10820 14020 10980
rect 14180 10820 14820 10980
rect 14980 10820 15620 10980
rect 15780 10820 16500 10980
rect 500 10180 16500 10820
rect 500 10020 1220 10180
rect 1380 10020 2020 10180
rect 2180 10020 2820 10180
rect 2980 10020 3620 10180
rect 3780 10020 4420 10180
rect 4580 10020 5220 10180
rect 5380 10020 6020 10180
rect 6180 10020 6820 10180
rect 6980 10020 7620 10180
rect 7780 10020 8420 10180
rect 8580 10020 9220 10180
rect 9380 10020 10020 10180
rect 10180 10020 10820 10180
rect 10980 10020 11620 10180
rect 11780 10020 12420 10180
rect 12580 10020 13220 10180
rect 13380 10020 14020 10180
rect 14180 10020 14820 10180
rect 14980 10020 15620 10180
rect 15780 10020 16500 10180
rect 500 9380 16500 10020
rect 500 9220 1220 9380
rect 1380 9220 2020 9380
rect 2180 9220 2820 9380
rect 2980 9220 3620 9380
rect 3780 9220 4420 9380
rect 4580 9220 5220 9380
rect 5380 9220 6020 9380
rect 6180 9220 6820 9380
rect 6980 9220 7620 9380
rect 7780 9220 8420 9380
rect 8580 9220 9220 9380
rect 9380 9220 10020 9380
rect 10180 9220 10820 9380
rect 10980 9220 11620 9380
rect 11780 9220 12420 9380
rect 12580 9220 13220 9380
rect 13380 9220 14020 9380
rect 14180 9220 14820 9380
rect 14980 9220 15620 9380
rect 15780 9220 16500 9380
rect 500 8580 16500 9220
rect 500 8420 1220 8580
rect 1380 8420 2020 8580
rect 2180 8420 2820 8580
rect 2980 8420 3620 8580
rect 3780 8420 4420 8580
rect 4580 8420 5220 8580
rect 5380 8420 6020 8580
rect 6180 8420 6820 8580
rect 6980 8420 7620 8580
rect 7780 8420 8420 8580
rect 8580 8420 9220 8580
rect 9380 8420 10020 8580
rect 10180 8420 10820 8580
rect 10980 8420 11620 8580
rect 11780 8420 12420 8580
rect 12580 8420 13220 8580
rect 13380 8420 14020 8580
rect 14180 8420 14820 8580
rect 14980 8420 15620 8580
rect 15780 8420 16500 8580
rect 500 7780 16500 8420
rect 500 7620 1220 7780
rect 1380 7620 2020 7780
rect 2180 7620 2820 7780
rect 2980 7620 3620 7780
rect 3780 7620 4420 7780
rect 4580 7620 5220 7780
rect 5380 7620 6020 7780
rect 6180 7620 6820 7780
rect 6980 7620 7620 7780
rect 7780 7620 8420 7780
rect 8580 7620 9220 7780
rect 9380 7620 10020 7780
rect 10180 7620 10820 7780
rect 10980 7620 11620 7780
rect 11780 7620 12420 7780
rect 12580 7620 13220 7780
rect 13380 7620 14020 7780
rect 14180 7620 14820 7780
rect 14980 7620 15620 7780
rect 15780 7620 16500 7780
rect 500 6980 16500 7620
rect 500 6820 1220 6980
rect 1380 6820 2020 6980
rect 2180 6820 2820 6980
rect 2980 6820 3620 6980
rect 3780 6820 4420 6980
rect 4580 6820 5220 6980
rect 5380 6820 6020 6980
rect 6180 6820 6820 6980
rect 6980 6820 7620 6980
rect 7780 6820 8420 6980
rect 8580 6820 9220 6980
rect 9380 6820 10020 6980
rect 10180 6820 10820 6980
rect 10980 6820 11620 6980
rect 11780 6820 12420 6980
rect 12580 6820 13220 6980
rect 13380 6820 14020 6980
rect 14180 6820 14820 6980
rect 14980 6820 15620 6980
rect 15780 6820 16500 6980
rect 500 6180 16500 6820
rect 500 6020 1220 6180
rect 1380 6020 2020 6180
rect 2180 6020 2820 6180
rect 2980 6020 3620 6180
rect 3780 6020 4420 6180
rect 4580 6020 5220 6180
rect 5380 6020 6020 6180
rect 6180 6020 6820 6180
rect 6980 6020 7620 6180
rect 7780 6020 8420 6180
rect 8580 6020 9220 6180
rect 9380 6020 10020 6180
rect 10180 6020 10820 6180
rect 10980 6020 11620 6180
rect 11780 6020 12420 6180
rect 12580 6020 13220 6180
rect 13380 6020 14020 6180
rect 14180 6020 14820 6180
rect 14980 6020 15620 6180
rect 15780 6020 16500 6180
rect 500 5380 16500 6020
rect 500 5220 1220 5380
rect 1380 5220 2020 5380
rect 2180 5220 2820 5380
rect 2980 5220 3620 5380
rect 3780 5220 4420 5380
rect 4580 5220 5220 5380
rect 5380 5220 6020 5380
rect 6180 5220 6820 5380
rect 6980 5220 7620 5380
rect 7780 5220 8420 5380
rect 8580 5220 9220 5380
rect 9380 5220 10020 5380
rect 10180 5220 10820 5380
rect 10980 5220 11620 5380
rect 11780 5220 12420 5380
rect 12580 5220 13220 5380
rect 13380 5220 14020 5380
rect 14180 5220 14820 5380
rect 14980 5220 15620 5380
rect 15780 5220 16500 5380
rect 500 4580 16500 5220
rect 500 4420 1220 4580
rect 1380 4420 2020 4580
rect 2180 4420 2820 4580
rect 2980 4420 3620 4580
rect 3780 4420 4420 4580
rect 4580 4420 5220 4580
rect 5380 4420 6020 4580
rect 6180 4420 6820 4580
rect 6980 4420 7620 4580
rect 7780 4420 8420 4580
rect 8580 4420 9220 4580
rect 9380 4420 10020 4580
rect 10180 4420 10820 4580
rect 10980 4420 11620 4580
rect 11780 4420 12420 4580
rect 12580 4420 13220 4580
rect 13380 4420 14020 4580
rect 14180 4420 14820 4580
rect 14980 4420 15620 4580
rect 15780 4420 16500 4580
rect 500 3780 16500 4420
rect 500 3620 1220 3780
rect 1380 3620 2020 3780
rect 2180 3620 2820 3780
rect 2980 3620 3620 3780
rect 3780 3620 4420 3780
rect 4580 3620 5220 3780
rect 5380 3620 6020 3780
rect 6180 3620 6820 3780
rect 6980 3620 7620 3780
rect 7780 3620 8420 3780
rect 8580 3620 9220 3780
rect 9380 3620 10020 3780
rect 10180 3620 10820 3780
rect 10980 3620 11620 3780
rect 11780 3620 12420 3780
rect 12580 3620 13220 3780
rect 13380 3620 14020 3780
rect 14180 3620 14820 3780
rect 14980 3620 15620 3780
rect 15780 3620 16500 3780
rect 500 2980 16500 3620
rect 500 2820 1220 2980
rect 1380 2820 2020 2980
rect 2180 2820 2820 2980
rect 2980 2820 3620 2980
rect 3780 2820 4420 2980
rect 4580 2820 5220 2980
rect 5380 2820 6020 2980
rect 6180 2820 6820 2980
rect 6980 2820 7620 2980
rect 7780 2820 8420 2980
rect 8580 2820 9220 2980
rect 9380 2820 10020 2980
rect 10180 2820 10820 2980
rect 10980 2820 11620 2980
rect 11780 2820 12420 2980
rect 12580 2820 13220 2980
rect 13380 2820 14020 2980
rect 14180 2820 14820 2980
rect 14980 2820 15620 2980
rect 15780 2820 16500 2980
rect 500 2180 16500 2820
rect 500 2020 1220 2180
rect 1380 2020 2020 2180
rect 2180 2020 2820 2180
rect 2980 2020 3620 2180
rect 3780 2020 4420 2180
rect 4580 2020 5220 2180
rect 5380 2020 6020 2180
rect 6180 2020 6820 2180
rect 6980 2020 7620 2180
rect 7780 2020 8420 2180
rect 8580 2020 9220 2180
rect 9380 2020 10020 2180
rect 10180 2020 10820 2180
rect 10980 2020 11620 2180
rect 11780 2020 12420 2180
rect 12580 2020 13220 2180
rect 13380 2020 14020 2180
rect 14180 2020 14820 2180
rect 14980 2020 15620 2180
rect 15780 2020 16500 2180
rect 500 1380 16500 2020
rect 500 1220 1220 1380
rect 1380 1220 2020 1380
rect 2180 1220 2820 1380
rect 2980 1220 3620 1380
rect 3780 1220 4420 1380
rect 4580 1220 5220 1380
rect 5380 1220 6020 1380
rect 6180 1220 6820 1380
rect 6980 1220 7620 1380
rect 7780 1220 8420 1380
rect 8580 1220 9220 1380
rect 9380 1220 10020 1380
rect 10180 1220 10820 1380
rect 10980 1220 11620 1380
rect 11780 1220 12420 1380
rect 12580 1220 13220 1380
rect 13380 1220 14020 1380
rect 14180 1220 14820 1380
rect 14980 1220 15620 1380
rect 15780 1220 16500 1380
rect 500 500 16500 1220
<< labels >>
flabel m3contact 8500 8500 8500 8500 0 FreeSans 10000 0 0 0 PIC_0.PAD
<< end >>
