* NGSPICE file created from BUFX2.ext - technology: scmos

.subckt BUFX2 A Y vdd gnd
M1000 gnd A a_4_12# gnd nfet w=3u l=0.6u
+  ad=4.95p pd=7.8u as=4.5p ps=9u
M1001 vdd A a_4_12# vdd pfet w=6u l=0.6u
+  ad=9.900001p pd=13.8u as=9p ps=15.000001u
M1002 Y a_4_12# vdd vdd pfet w=12u l=0.6u
+  ad=18p pd=27.000002u as=9.900001p ps=13.8u
M1003 Y a_4_12# gnd gnd nfet w=6u l=0.6u
+  ad=9p pd=15.000001u as=4.95p ps=7.8u
.ends

