magic
tech scmos
magscale 1 2
timestamp 1726555477
<< nwell >>
rect -12 154 152 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 48 14 52 54
rect 68 14 72 54
rect 78 14 82 54
rect 100 14 104 54
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 50 166 54 246
rect 70 166 74 246
rect 78 166 82 246
rect 100 166 104 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 48 40 54
rect 24 14 26 48
rect 38 14 40 48
rect 44 14 48 54
rect 52 50 68 54
rect 52 14 54 50
rect 66 14 68 50
rect 72 14 78 54
rect 82 48 100 54
rect 82 14 84 48
rect 96 14 100 48
rect 104 14 106 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 180 26 246
rect 38 180 40 246
rect 24 166 40 180
rect 44 166 50 246
rect 54 166 56 246
rect 68 166 70 246
rect 74 166 78 246
rect 82 180 84 246
rect 98 180 100 246
rect 82 166 100 180
rect 104 166 106 246
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 48
rect 54 14 66 50
rect 84 14 96 48
rect 106 14 118 54
<< pdcontact >>
rect 6 166 18 246
rect 26 180 38 246
rect 56 166 68 246
rect 84 180 98 246
rect 106 166 118 246
<< psubstratepcontact >>
rect -6 -6 146 6
<< nsubstratencontact >>
rect -6 254 146 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 50 246 54 250
rect 70 246 74 250
rect 78 246 82 250
rect 100 246 104 250
rect 20 102 24 166
rect 40 162 44 166
rect 16 90 24 102
rect 20 54 24 90
rect 30 158 44 162
rect 30 130 35 158
rect 50 150 54 166
rect 30 118 33 130
rect 30 62 35 118
rect 53 96 57 138
rect 70 116 74 166
rect 78 160 82 166
rect 100 160 104 166
rect 78 156 104 160
rect 53 92 72 96
rect 30 58 44 62
rect 40 54 44 58
rect 48 54 52 72
rect 68 54 72 92
rect 100 62 104 156
rect 78 58 104 62
rect 78 54 82 58
rect 100 54 104 58
rect 20 10 24 14
rect 40 10 44 14
rect 48 10 52 14
rect 68 10 72 14
rect 78 10 82 14
rect 100 10 104 14
<< polycontact >>
rect 4 90 16 102
rect 45 138 57 150
rect 33 118 45 130
rect 65 104 77 116
rect 44 72 56 84
rect 104 116 116 128
<< metal1 >>
rect -6 266 146 268
rect -6 252 146 254
rect 26 246 38 252
rect 84 246 98 252
rect 18 166 23 172
rect 6 163 23 166
rect 68 166 77 172
rect 23 152 57 158
rect 45 150 57 152
rect 69 136 77 166
rect 97 166 106 172
rect 97 163 118 166
rect 77 122 89 129
rect 33 104 43 118
rect 16 98 17 102
rect 65 98 77 104
rect 16 90 44 98
rect 58 90 77 98
rect 83 84 89 122
rect 64 78 89 84
rect 11 58 23 72
rect 11 54 18 58
rect 64 50 70 78
rect 97 58 117 65
rect 66 39 70 50
rect 106 54 117 58
rect 26 8 38 14
rect 84 8 96 14
rect -6 6 146 8
rect -6 -8 146 -6
<< m2contact >>
rect 23 158 37 172
rect 83 158 97 172
rect 63 122 77 136
rect 3 102 17 116
rect 43 104 57 118
rect 44 84 58 98
rect 103 102 117 116
rect 23 58 37 72
rect 83 58 97 72
<< metal2 >>
rect 6 116 14 134
rect 26 72 32 158
rect 66 136 74 154
rect 87 116 94 158
rect 57 110 94 116
rect 87 72 94 110
rect 106 86 114 102
<< m1p >>
rect -6 252 146 268
rect -6 -8 146 8
<< m2p >>
rect 66 138 74 154
rect 6 118 14 134
rect 106 86 114 100
<< labels >>
rlabel metal1 -6 252 126 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 126 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal2 10 130 10 130 1 A
port 1 n signal input
rlabel metal2 70 150 70 150 1 Y
port 3 n signal output
rlabel metal2 110 90 110 90 5 B
port 2 n signal input
<< properties >>
string FIXED_BBOX 0 0 140 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
