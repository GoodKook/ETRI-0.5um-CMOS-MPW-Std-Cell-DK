magic
tech scmos
magscale 1 2
timestamp 1727733069
<< nwell >>
rect -12 134 133 252
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
rect 80 14 84 54
<< ptransistor >>
rect 20 146 24 226
rect 40 146 44 226
rect 60 146 64 226
rect 80 146 84 226
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 26 54
rect 38 14 40 54
rect 44 14 46 54
rect 58 14 60 54
rect 64 14 66 54
rect 78 14 80 54
rect 84 14 86 54
<< pdiffusion >>
rect 18 146 20 226
rect 24 146 26 226
rect 38 146 40 226
rect 44 146 46 226
rect 58 146 60 226
rect 64 146 66 226
rect 78 146 80 226
rect 84 146 86 226
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 54
rect 46 14 58 54
rect 66 14 78 54
rect 86 14 98 54
<< pdcontact >>
rect 6 146 18 226
rect 26 146 38 226
rect 46 146 58 226
rect 66 146 78 226
rect 86 146 98 226
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 234 126 246
<< polysilicon >>
rect 20 226 24 230
rect 40 226 44 230
rect 60 226 64 230
rect 80 226 84 230
rect 20 142 24 146
rect 40 142 44 146
rect 60 142 64 146
rect 80 142 84 146
rect 20 138 84 142
rect 20 109 26 138
rect 20 97 24 109
rect 20 62 26 97
rect 20 58 84 62
rect 20 54 24 58
rect 40 54 44 58
rect 60 54 64 58
rect 80 54 84 58
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
rect 80 10 84 14
<< polycontact >>
rect 24 97 36 109
<< metal1 >>
rect -6 246 126 248
rect -6 232 126 234
rect 6 226 18 232
rect 46 226 58 232
rect 86 226 98 232
rect 26 140 38 146
rect 66 140 74 146
rect 26 134 74 140
rect 66 97 74 134
rect 23 83 37 97
rect 63 83 77 97
rect 66 68 74 83
rect 26 60 74 68
rect 26 54 34 60
rect 66 54 74 60
rect 6 8 18 14
rect 46 8 58 14
rect 86 8 98 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m1p >>
rect 23 83 37 97
rect 63 83 77 97
<< labels >>
rlabel metal1 -6 -8 126 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 63 83 77 97 0 Y
port 1 nsew signal output
rlabel metal1 23 83 37 97 0 A
port 0 nsew signal input
rlabel metal1 -6 232 126 248 0 vdd
port 2 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 120 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
