magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -56 -56 254 84
<< diffusion >>
rect 5 5 193 23
<< genericcontact >>
rect 12 11 18 17
rect 40 11 46 17
rect 68 11 74 17
rect 96 11 102 17
rect 124 11 130 17
rect 152 11 158 17
rect 180 11 186 17
<< metal1 >>
rect 4 4 194 24
<< end >>
