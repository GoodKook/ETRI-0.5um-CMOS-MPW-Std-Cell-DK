magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -60 -60 78 78
<< polysilicon >>
rect 1 15 17 17
rect 1 3 3 15
rect 15 3 17 15
rect 1 1 17 3
<< polycontact >>
rect 3 3 15 15
<< metal1 >>
rect 0 15 18 18
rect 0 3 3 15
rect 15 3 18 15
rect 0 0 18 3
<< end >>
