magic
tech scmos
magscale 1 2
timestamp 1727136778
<< error_p >>
rect 44 166 48 174
<< nwell >>
rect -13 154 153 272
<< ntransistor >>
rect 18 14 22 54
rect 58 14 62 54
rect 78 14 82 54
rect 98 14 102 54
rect 118 14 122 54
<< ptransistor >>
rect 18 166 22 246
rect 58 166 62 246
rect 78 166 82 246
rect 98 166 102 246
rect 118 166 122 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 24 54
rect 56 14 58 54
rect 62 26 64 54
rect 76 26 78 54
rect 62 14 78 26
rect 82 14 84 54
rect 96 14 98 54
rect 102 48 118 54
rect 102 14 104 48
rect 116 14 118 48
rect 122 14 124 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 24 246
rect 56 166 58 246
rect 62 234 78 246
rect 62 166 64 234
rect 76 166 78 234
rect 82 166 84 246
rect 96 166 98 246
rect 102 242 118 246
rect 102 180 104 242
rect 116 180 118 242
rect 102 166 118 180
rect 122 166 124 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 54
rect 44 14 56 54
rect 64 26 76 54
rect 84 14 96 54
rect 104 14 116 48
rect 124 14 136 54
<< pdcontact >>
rect 4 166 16 246
rect 24 166 36 246
rect 44 166 56 246
rect 64 166 76 234
rect 84 166 96 246
rect 104 180 116 242
rect 124 166 136 246
<< psubstratepcontact >>
rect -7 -6 147 6
<< nsubstratencontact >>
rect -7 254 147 266
<< polysilicon >>
rect 18 246 22 250
rect 58 246 62 250
rect 78 246 82 250
rect 98 246 102 250
rect 118 246 122 250
rect 18 103 22 166
rect 58 162 62 166
rect 78 162 82 166
rect 38 158 82 162
rect 98 162 102 166
rect 118 162 122 166
rect 98 158 122 162
rect 38 153 42 158
rect 18 62 22 91
rect 118 62 122 158
rect 18 58 82 62
rect 18 54 22 58
rect 58 54 62 58
rect 78 54 82 58
rect 98 58 122 62
rect 98 54 102 58
rect 118 54 122 58
rect 18 10 22 14
rect 58 10 62 14
rect 78 10 82 14
rect 98 10 102 14
rect 118 10 122 14
<< polycontact >>
rect 30 141 42 153
rect 10 91 22 103
rect 106 91 118 103
<< metal1 >>
rect -7 266 147 268
rect -7 252 147 254
rect 4 246 16 252
rect 56 240 84 246
rect 104 242 116 252
rect 96 166 124 174
rect 30 153 36 166
rect 30 54 36 141
rect 64 117 70 166
rect 64 54 70 103
rect 84 54 132 60
rect 56 14 84 20
rect 4 8 16 14
rect 104 8 116 14
rect -7 6 147 8
rect -7 -8 147 -6
<< m2contact >>
rect 6 103 20 117
rect 64 103 78 117
rect 104 103 118 117
<< metal2 >>
rect 6 117 14 134
rect 66 117 74 134
rect 106 117 114 134
<< m1p >>
rect -7 252 147 268
rect -7 -8 147 8
<< m2p >>
rect 6 117 14 134
rect 66 117 74 134
rect 106 117 114 134
<< labels >>
rlabel metal1 -7 252 147 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -7 -8 147 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal2 11 130 11 130 3 EN
port 2 n signal input
rlabel metal2 70 131 70 131 3 Y
port 3 n signal output
rlabel metal2 110 131 110 131 7 A
port 1 n signal input
<< properties >>
string FIXED_BBOX 0 0 140 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
