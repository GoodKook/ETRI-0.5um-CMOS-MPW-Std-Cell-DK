magic
tech scmos
magscale 1 3
timestamp 1725342160
<< genericcontact >>
rect 14 15 20 21
rect 1020 15 1026 21
<< metal1 >>
rect 8 8 26 28
rect 1014 8 1032 28
<< pseudo_rpoly2 >>
rect 8 8 1032 28
<< end >>
