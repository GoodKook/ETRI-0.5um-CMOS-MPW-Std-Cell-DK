magic
tech scmos
magscale 1 2
timestamp 1727840468
<< nwell >>
rect -14 134 132 252
<< ntransistor >>
rect 24 14 28 54
rect 32 14 36 54
rect 52 14 56 54
rect 60 14 64 54
<< ptransistor >>
rect 20 146 24 226
rect 40 146 44 226
rect 60 146 64 226
rect 80 146 84 226
<< ndiffusion >>
rect 22 14 24 54
rect 28 14 32 54
rect 36 14 38 54
rect 50 14 52 54
rect 56 14 60 54
rect 64 14 66 54
<< pdiffusion >>
rect 18 148 20 226
rect 6 146 20 148
rect 24 160 26 226
rect 38 160 40 226
rect 24 146 40 160
rect 44 148 46 226
rect 58 148 60 226
rect 44 146 60 148
rect 64 214 80 226
rect 64 146 66 214
rect 78 146 80 214
rect 84 146 86 226
<< ndcontact >>
rect 10 14 22 54
rect 38 14 50 54
rect 66 14 78 54
<< pdcontact >>
rect 6 148 18 226
rect 26 160 38 226
rect 46 148 58 226
rect 66 146 78 214
rect 86 146 98 226
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 234 126 246
<< polysilicon >>
rect 20 226 24 230
rect 40 226 44 230
rect 60 226 64 230
rect 80 226 84 230
rect 20 124 24 146
rect 40 124 44 146
rect 5 123 24 124
rect 17 118 24 123
rect 32 118 44 124
rect 11 69 17 111
rect 32 89 36 118
rect 60 89 64 146
rect 80 124 84 146
rect 80 123 90 124
rect 80 118 84 123
rect 60 77 63 89
rect 11 62 28 69
rect 24 54 28 62
rect 32 54 36 77
rect 60 75 64 77
rect 52 68 64 75
rect 52 54 56 68
rect 84 63 90 111
rect 60 59 90 63
rect 60 54 64 59
rect 24 10 28 14
rect 32 10 36 14
rect 52 10 56 14
rect 60 10 64 14
<< polycontact >>
rect 5 111 17 123
rect 84 111 96 123
rect 25 77 37 89
rect 63 77 75 89
<< metal1 >>
rect -6 246 126 248
rect -6 232 126 234
rect 26 226 38 232
rect 18 148 46 154
rect 58 220 86 226
rect 66 140 78 146
rect 51 134 78 140
rect 51 111 57 134
rect 43 54 50 97
rect 10 8 22 14
rect 66 8 78 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m2contact >>
rect 3 97 17 111
rect 23 89 37 103
rect 43 97 57 111
rect 63 89 77 103
rect 83 97 97 111
<< metal2 >>
rect 3 83 17 97
rect 23 103 37 117
rect 43 83 57 97
rect 63 103 77 117
rect 83 83 97 97
<< m2p >>
rect 23 103 37 117
rect 63 103 77 117
rect 3 83 17 97
rect 43 83 57 97
rect 83 83 97 97
<< labels >>
rlabel metal1 -6 -8 126 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 -6 232 126 248 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal2 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal2 23 103 37 117 0 B
port 1 nsew signal input
rlabel metal2 83 83 97 97 0 C
port 2 nsew signal input
rlabel metal2 63 103 77 117 0 D
port 3 nsew signal input
rlabel metal2 43 83 57 97 0 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
